.subckt dig22inv a o vccx vssx
.ends
.subckt ckt_dig_1 vi vo vccx vssx
xi0 vi vo vccx vssx dig22inv
.ends ckt_dig_1
.END
