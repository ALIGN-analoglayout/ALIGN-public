MACRO Switch_NMOS_B_nfin48_nf1_m1_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin48_nf1_m1_n12_X2_Y2 0 0 ;
  SIZE 0.8000 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.2960 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.8880 0.3400 2.1360 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 0.5160 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 1.2440 0.5960 1.2760 ;
    LAYER M2 ;
      RECT 0.2040 1.3280 0.5160 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.5160 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.2440 0.1760 1.2760 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER V2 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
  END
END Switch_NMOS_B_nfin48_nf1_m1_n12_X2_Y2
MACRO DP_NMOS_B_nfin48_n12_X4_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin48_n12_X4_Y1 0 0 ;
  SIZE 1.7600 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.5560 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 1.4760 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 1.3160 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 1.4760 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.9920 1.3160 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 1.4760 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.8880 1.2960 1.1280 ;
    LAYER M1 ;
      RECT 1.2640 1.3920 1.2960 1.6320 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.0480 1.4560 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.8880 1.4560 1.1280 ;
    LAYER M1 ;
      RECT 1.4240 1.3920 1.4560 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.3440 0.0680 1.3760 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.4240 0.1520 1.4560 0.1840 ;
    LAYER V1 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V1 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 1.2640 0.2360 1.2960 0.2680 ;
    LAYER V1 ;
      RECT 1.2640 0.9920 1.2960 1.0240 ;
    LAYER V1 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9920 0.6560 1.0240 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.4040 1.2960 0.4360 ;
    LAYER V0 ;
      RECT 1.2640 0.5300 1.2960 0.5620 ;
    LAYER V0 ;
      RECT 1.2640 0.6560 1.2960 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V0 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.4040 1.4560 0.4360 ;
    LAYER V0 ;
      RECT 1.4240 0.5300 1.4560 0.5620 ;
    LAYER V0 ;
      RECT 1.4240 0.6560 1.4560 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V0 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
  END
END DP_NMOS_B_nfin48_n12_X4_Y1
MACRO Switch_NMOS_nfin144_n12_X4_Y3
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin144_n12_X4_Y3 0 0 ;
  SIZE 1.1200 BY 4.2000 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 3.9000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 2.5560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.8880 0.5000 3.3120 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.4000 0.3360 3.1440 ;
    LAYER M1 ;
      RECT 0.3040 3.2400 0.3360 3.4800 ;
    LAYER M1 ;
      RECT 0.3040 3.7440 0.3360 3.9840 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.2240 2.4000 0.2560 3.1440 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.4000 0.4160 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.4000 0.4960 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 3.2400 0.4960 3.4800 ;
    LAYER M1 ;
      RECT 0.4640 3.7440 0.4960 3.9840 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 2.4000 0.5760 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.4000 0.6560 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 3.2400 0.6560 3.4800 ;
    LAYER M1 ;
      RECT 0.6240 3.7440 0.6560 3.9840 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.4000 0.7360 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.4000 0.8160 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 3.2400 0.8160 3.4800 ;
    LAYER M1 ;
      RECT 0.7840 3.7440 0.8160 3.9840 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.8640 2.4000 0.8960 3.1440 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.8360 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 0.8360 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.8360 2.1160 ;
    LAYER M2 ;
      RECT 0.2040 2.4200 0.9160 2.4520 ;
    LAYER M2 ;
      RECT 0.2840 3.8480 0.8360 3.8800 ;
    LAYER M2 ;
      RECT 0.2840 2.5040 0.8360 2.5360 ;
    LAYER M2 ;
      RECT 0.2840 3.2600 0.8360 3.2920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 2.4200 0.2560 2.4520 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 2.4200 0.4160 2.4520 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 2.4200 0.5760 2.4520 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 2.4200 0.7360 2.4520 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 2.4200 0.8960 2.4520 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.5040 0.6560 2.5360 ;
    LAYER V1 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V1 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.5040 0.8160 2.5360 ;
    LAYER V1 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V1 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER V1 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V1 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.5040 0.4960 2.5360 ;
    LAYER V1 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V1 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.4200 0.3360 2.4520 ;
    LAYER V2 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.3840 2.5040 0.4160 2.5360 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V2 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.7560 0.3360 2.7880 ;
    LAYER V0 ;
      RECT 0.3040 2.8820 0.3360 2.9140 ;
    LAYER V0 ;
      RECT 0.3040 3.0080 0.3360 3.0400 ;
    LAYER V0 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.2240 2.7560 0.2560 2.7880 ;
    LAYER V0 ;
      RECT 0.2240 2.8820 0.2560 2.9140 ;
    LAYER V0 ;
      RECT 0.2240 3.0080 0.2560 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.7560 0.4960 2.7880 ;
    LAYER V0 ;
      RECT 0.4640 2.8820 0.4960 2.9140 ;
    LAYER V0 ;
      RECT 0.4640 3.0080 0.4960 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.7560 0.6560 2.7880 ;
    LAYER V0 ;
      RECT 0.6240 2.8820 0.6560 2.9140 ;
    LAYER V0 ;
      RECT 0.6240 3.0080 0.6560 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.7560 0.8160 2.7880 ;
    LAYER V0 ;
      RECT 0.7840 2.8820 0.8160 2.9140 ;
    LAYER V0 ;
      RECT 0.7840 3.0080 0.8160 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
  END
END Switch_NMOS_nfin144_n12_X4_Y3
MACRO Switch_NMOS_B_nfin48_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin48_n12_X2_Y2 0 0 ;
  SIZE 0.8000 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.2960 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.8880 0.3400 2.1360 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 0.5160 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 1.2440 0.5960 1.2760 ;
    LAYER M2 ;
      RECT 0.2040 1.3280 0.5160 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.5160 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.2440 0.1760 1.2760 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER V2 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
  END
END Switch_NMOS_B_nfin48_n12_X2_Y2
MACRO Switch_NMOS_nfin72_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin72_n12_X3_Y2 0 0 ;
  SIZE 0.9600 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.1320 0.3400 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.8880 0.4200 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.6760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.6760 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.7560 1.2760 ;
    LAYER M2 ;
      RECT 0.2040 2.6720 0.6760 2.7040 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 0.6760 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.6760 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V2 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V2 ;
      RECT 0.2240 2.6720 0.2560 2.7040 ;
    LAYER V2 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V2 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V2 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V2 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
  END
END Switch_NMOS_nfin72_n12_X3_Y2
MACRO DP_NMOS_B_nfin192_n12_X8_Y2
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin192_n12_X8_Y2 0 0 ;
  SIZE 3.0400 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1800 0.0480 1.2200 1.2960 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2600 0.1320 1.3000 1.3800 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3400 0.2160 1.3800 1.4640 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4200 0.8880 1.4600 2.1360 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5000 0.9720 1.5400 2.2200 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 2.7560 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.5680 0.8160 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.2240 0.9760 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 2.0640 0.9760 2.3040 ;
    LAYER M1 ;
      RECT 0.9440 2.5680 0.9760 2.8080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.2240 1.1360 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 2.0640 1.1360 2.3040 ;
    LAYER M1 ;
      RECT 1.1040 2.5680 1.1360 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.8880 1.2960 1.1280 ;
    LAYER M1 ;
      RECT 1.2640 1.2240 1.2960 1.9680 ;
    LAYER M1 ;
      RECT 1.2640 2.0640 1.2960 2.3040 ;
    LAYER M1 ;
      RECT 1.2640 2.5680 1.2960 2.8080 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.4240 0.0480 1.4560 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.8880 1.4560 1.1280 ;
    LAYER M1 ;
      RECT 1.4240 1.2240 1.4560 1.9680 ;
    LAYER M1 ;
      RECT 1.4240 2.0640 1.4560 2.3040 ;
    LAYER M1 ;
      RECT 1.4240 2.5680 1.4560 2.8080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.2240 1.6160 1.9680 ;
    LAYER M1 ;
      RECT 1.5840 2.0640 1.6160 2.3040 ;
    LAYER M1 ;
      RECT 1.5840 2.5680 1.6160 2.8080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 1.2240 1.6960 1.9680 ;
    LAYER M1 ;
      RECT 1.7440 0.0480 1.7760 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.8880 1.7760 1.1280 ;
    LAYER M1 ;
      RECT 1.7440 1.2240 1.7760 1.9680 ;
    LAYER M1 ;
      RECT 1.7440 2.0640 1.7760 2.3040 ;
    LAYER M1 ;
      RECT 1.7440 2.5680 1.7760 2.8080 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.8240 1.2240 1.8560 1.9680 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.8880 1.9360 1.1280 ;
    LAYER M1 ;
      RECT 1.9040 1.2240 1.9360 1.9680 ;
    LAYER M1 ;
      RECT 1.9040 2.0640 1.9360 2.3040 ;
    LAYER M1 ;
      RECT 1.9040 2.5680 1.9360 2.8080 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 1.9840 1.2240 2.0160 1.9680 ;
    LAYER M1 ;
      RECT 2.0640 0.0480 2.0960 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.8880 2.0960 1.1280 ;
    LAYER M1 ;
      RECT 2.0640 1.2240 2.0960 1.9680 ;
    LAYER M1 ;
      RECT 2.0640 2.0640 2.0960 2.3040 ;
    LAYER M1 ;
      RECT 2.0640 2.5680 2.0960 2.8080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.1440 1.2240 2.1760 1.9680 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.2240 2.2560 1.9680 ;
    LAYER M1 ;
      RECT 2.2240 2.0640 2.2560 2.3040 ;
    LAYER M1 ;
      RECT 2.2240 2.5680 2.2560 2.8080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 1.2240 2.3360 1.9680 ;
    LAYER M1 ;
      RECT 2.3840 0.0480 2.4160 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.8880 2.4160 1.1280 ;
    LAYER M1 ;
      RECT 2.3840 1.2240 2.4160 1.9680 ;
    LAYER M1 ;
      RECT 2.3840 2.0640 2.4160 2.3040 ;
    LAYER M1 ;
      RECT 2.3840 2.5680 2.4160 2.8080 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER M1 ;
      RECT 2.4640 1.2240 2.4960 1.9680 ;
    LAYER M1 ;
      RECT 2.5440 0.0480 2.5760 0.7920 ;
    LAYER M1 ;
      RECT 2.5440 0.8880 2.5760 1.1280 ;
    LAYER M1 ;
      RECT 2.5440 1.2240 2.5760 1.9680 ;
    LAYER M1 ;
      RECT 2.5440 2.0640 2.5760 2.3040 ;
    LAYER M1 ;
      RECT 2.5440 2.5680 2.5760 2.8080 ;
    LAYER M1 ;
      RECT 2.6240 0.0480 2.6560 0.7920 ;
    LAYER M1 ;
      RECT 2.6240 1.2240 2.6560 1.9680 ;
    LAYER M1 ;
      RECT 2.7040 0.0480 2.7360 0.7920 ;
    LAYER M1 ;
      RECT 2.7040 0.8880 2.7360 1.1280 ;
    LAYER M1 ;
      RECT 2.7040 1.2240 2.7360 1.9680 ;
    LAYER M1 ;
      RECT 2.7040 2.0640 2.7360 2.3040 ;
    LAYER M1 ;
      RECT 2.7040 2.5680 2.7360 2.8080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER M1 ;
      RECT 2.7840 1.2240 2.8160 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 2.7560 0.1840 ;
    LAYER M2 ;
      RECT 0.4440 0.2360 2.5960 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 2.7560 0.9400 ;
    LAYER M2 ;
      RECT 0.4440 0.9920 2.5960 1.0240 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 2.8360 1.2760 ;
    LAYER M2 ;
      RECT 0.4440 1.3280 2.5960 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 1.4120 2.7560 1.4440 ;
    LAYER M2 ;
      RECT 0.4440 2.0840 2.5960 2.1160 ;
    LAYER M2 ;
      RECT 0.2840 2.1680 2.7560 2.2000 ;
    LAYER V1 ;
      RECT 2.6240 0.0680 2.6560 0.1000 ;
    LAYER V1 ;
      RECT 2.6240 1.2440 2.6560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 1.2440 2.8160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.3440 0.0680 1.3760 0.1000 ;
    LAYER V1 ;
      RECT 1.3440 1.2440 1.3760 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 1.2440 1.6960 1.2760 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 1.2440 1.8560 1.2760 ;
    LAYER V1 ;
      RECT 1.9840 0.0680 2.0160 0.1000 ;
    LAYER V1 ;
      RECT 1.9840 1.2440 2.0160 1.2760 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 1.2440 2.1760 1.2760 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 1.2440 2.3360 1.2760 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 1.2440 2.4960 1.2760 ;
    LAYER V1 ;
      RECT 2.7040 0.1520 2.7360 0.1840 ;
    LAYER V1 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V1 ;
      RECT 2.7040 1.4120 2.7360 1.4440 ;
    LAYER V1 ;
      RECT 2.7040 2.1680 2.7360 2.2000 ;
    LAYER V1 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4120 0.3360 1.4440 ;
    LAYER V1 ;
      RECT 0.3040 2.1680 0.3360 2.2000 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4120 0.8160 1.4440 ;
    LAYER V1 ;
      RECT 0.7840 2.1680 0.8160 2.2000 ;
    LAYER V1 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4120 0.9760 1.4440 ;
    LAYER V1 ;
      RECT 0.9440 2.1680 0.9760 2.2000 ;
    LAYER V1 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V1 ;
      RECT 1.4240 0.1520 1.4560 0.1840 ;
    LAYER V1 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V1 ;
      RECT 1.4240 1.4120 1.4560 1.4440 ;
    LAYER V1 ;
      RECT 1.4240 2.1680 1.4560 2.2000 ;
    LAYER V1 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V1 ;
      RECT 1.5840 0.1520 1.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4120 1.6160 1.4440 ;
    LAYER V1 ;
      RECT 1.5840 2.1680 1.6160 2.2000 ;
    LAYER V1 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V1 ;
      RECT 2.0640 0.1520 2.0960 0.1840 ;
    LAYER V1 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V1 ;
      RECT 2.0640 1.4120 2.0960 1.4440 ;
    LAYER V1 ;
      RECT 2.0640 2.1680 2.0960 2.2000 ;
    LAYER V1 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.2240 1.4120 2.2560 1.4440 ;
    LAYER V1 ;
      RECT 2.2240 2.1680 2.2560 2.2000 ;
    LAYER V1 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V1 ;
      RECT 2.5440 0.2360 2.5760 0.2680 ;
    LAYER V1 ;
      RECT 2.5440 0.9920 2.5760 1.0240 ;
    LAYER V1 ;
      RECT 2.5440 1.3280 2.5760 1.3600 ;
    LAYER V1 ;
      RECT 2.5440 2.0840 2.5760 2.1160 ;
    LAYER V1 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9920 0.6560 1.0240 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.3280 1.1360 1.3600 ;
    LAYER V1 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V1 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V1 ;
      RECT 1.2640 0.2360 1.2960 0.2680 ;
    LAYER V1 ;
      RECT 1.2640 0.9920 1.2960 1.0240 ;
    LAYER V1 ;
      RECT 1.2640 1.3280 1.2960 1.3600 ;
    LAYER V1 ;
      RECT 1.2640 2.0840 1.2960 2.1160 ;
    LAYER V1 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V1 ;
      RECT 1.7440 0.2360 1.7760 0.2680 ;
    LAYER V1 ;
      RECT 1.7440 0.9920 1.7760 1.0240 ;
    LAYER V1 ;
      RECT 1.7440 1.3280 1.7760 1.3600 ;
    LAYER V1 ;
      RECT 1.7440 2.0840 1.7760 2.1160 ;
    LAYER V1 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V1 ;
      RECT 1.9040 0.2360 1.9360 0.2680 ;
    LAYER V1 ;
      RECT 1.9040 0.9920 1.9360 1.0240 ;
    LAYER V1 ;
      RECT 1.9040 1.3280 1.9360 1.3600 ;
    LAYER V1 ;
      RECT 1.9040 2.0840 1.9360 2.1160 ;
    LAYER V1 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V1 ;
      RECT 2.3840 0.2360 2.4160 0.2680 ;
    LAYER V1 ;
      RECT 2.3840 0.9920 2.4160 1.0240 ;
    LAYER V1 ;
      RECT 2.3840 1.3280 2.4160 1.3600 ;
    LAYER V1 ;
      RECT 2.3840 2.0840 2.4160 2.1160 ;
    LAYER V1 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V2 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V2 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V2 ;
      RECT 1.2640 0.1520 1.2960 0.1840 ;
    LAYER V2 ;
      RECT 1.2640 1.3280 1.2960 1.3600 ;
    LAYER V2 ;
      RECT 1.3440 0.2360 1.3760 0.2680 ;
    LAYER V2 ;
      RECT 1.3440 1.4120 1.3760 1.4440 ;
    LAYER V2 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V2 ;
      RECT 1.4240 2.0840 1.4560 2.1160 ;
    LAYER V2 ;
      RECT 1.5040 0.9920 1.5360 1.0240 ;
    LAYER V2 ;
      RECT 1.5040 2.1680 1.5360 2.2000 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.5800 0.9760 1.6120 ;
    LAYER V0 ;
      RECT 0.9440 1.7060 0.9760 1.7380 ;
    LAYER V0 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.5800 1.1360 1.6120 ;
    LAYER V0 ;
      RECT 1.1040 1.7060 1.1360 1.7380 ;
    LAYER V0 ;
      RECT 1.1040 1.8320 1.1360 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.2640 0.4040 1.2960 0.4360 ;
    LAYER V0 ;
      RECT 1.2640 0.5300 1.2960 0.5620 ;
    LAYER V0 ;
      RECT 1.2640 0.6560 1.2960 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V0 ;
      RECT 1.2640 1.5800 1.2960 1.6120 ;
    LAYER V0 ;
      RECT 1.2640 1.7060 1.2960 1.7380 ;
    LAYER V0 ;
      RECT 1.2640 1.8320 1.2960 1.8640 ;
    LAYER V0 ;
      RECT 1.2640 2.0840 1.2960 2.1160 ;
    LAYER V0 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V0 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.4240 0.4040 1.4560 0.4360 ;
    LAYER V0 ;
      RECT 1.4240 0.5300 1.4560 0.5620 ;
    LAYER V0 ;
      RECT 1.4240 0.6560 1.4560 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V0 ;
      RECT 1.4240 1.5800 1.4560 1.6120 ;
    LAYER V0 ;
      RECT 1.4240 1.7060 1.4560 1.7380 ;
    LAYER V0 ;
      RECT 1.4240 1.8320 1.4560 1.8640 ;
    LAYER V0 ;
      RECT 1.4240 2.0840 1.4560 2.1160 ;
    LAYER V0 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V0 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.5800 1.6160 1.6120 ;
    LAYER V0 ;
      RECT 1.5840 1.7060 1.6160 1.7380 ;
    LAYER V0 ;
      RECT 1.5840 1.8320 1.6160 1.8640 ;
    LAYER V0 ;
      RECT 1.5840 2.0840 1.6160 2.1160 ;
    LAYER V0 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V0 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.7440 0.4040 1.7760 0.4360 ;
    LAYER V0 ;
      RECT 1.7440 0.5300 1.7760 0.5620 ;
    LAYER V0 ;
      RECT 1.7440 0.6560 1.7760 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.9080 1.7760 0.9400 ;
    LAYER V0 ;
      RECT 1.7440 1.5800 1.7760 1.6120 ;
    LAYER V0 ;
      RECT 1.7440 1.7060 1.7760 1.7380 ;
    LAYER V0 ;
      RECT 1.7440 1.8320 1.7760 1.8640 ;
    LAYER V0 ;
      RECT 1.7440 2.0840 1.7760 2.1160 ;
    LAYER V0 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V0 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.9040 0.4040 1.9360 0.4360 ;
    LAYER V0 ;
      RECT 1.9040 0.5300 1.9360 0.5620 ;
    LAYER V0 ;
      RECT 1.9040 0.6560 1.9360 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.9080 1.9360 0.9400 ;
    LAYER V0 ;
      RECT 1.9040 1.5800 1.9360 1.6120 ;
    LAYER V0 ;
      RECT 1.9040 1.7060 1.9360 1.7380 ;
    LAYER V0 ;
      RECT 1.9040 1.8320 1.9360 1.8640 ;
    LAYER V0 ;
      RECT 1.9040 2.0840 1.9360 2.1160 ;
    LAYER V0 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V0 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 1.5800 2.0160 1.6120 ;
    LAYER V0 ;
      RECT 1.9840 1.5800 2.0160 1.6120 ;
    LAYER V0 ;
      RECT 1.9840 1.7060 2.0160 1.7380 ;
    LAYER V0 ;
      RECT 1.9840 1.7060 2.0160 1.7380 ;
    LAYER V0 ;
      RECT 1.9840 1.8320 2.0160 1.8640 ;
    LAYER V0 ;
      RECT 1.9840 1.8320 2.0160 1.8640 ;
    LAYER V0 ;
      RECT 2.0640 0.4040 2.0960 0.4360 ;
    LAYER V0 ;
      RECT 2.0640 0.5300 2.0960 0.5620 ;
    LAYER V0 ;
      RECT 2.0640 0.6560 2.0960 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V0 ;
      RECT 2.0640 1.5800 2.0960 1.6120 ;
    LAYER V0 ;
      RECT 2.0640 1.7060 2.0960 1.7380 ;
    LAYER V0 ;
      RECT 2.0640 1.8320 2.0960 1.8640 ;
    LAYER V0 ;
      RECT 2.0640 2.0840 2.0960 2.1160 ;
    LAYER V0 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V0 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.5800 2.2560 1.6120 ;
    LAYER V0 ;
      RECT 2.2240 1.7060 2.2560 1.7380 ;
    LAYER V0 ;
      RECT 2.2240 1.8320 2.2560 1.8640 ;
    LAYER V0 ;
      RECT 2.2240 2.0840 2.2560 2.1160 ;
    LAYER V0 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V0 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 1.5800 2.3360 1.6120 ;
    LAYER V0 ;
      RECT 2.3040 1.5800 2.3360 1.6120 ;
    LAYER V0 ;
      RECT 2.3040 1.7060 2.3360 1.7380 ;
    LAYER V0 ;
      RECT 2.3040 1.7060 2.3360 1.7380 ;
    LAYER V0 ;
      RECT 2.3040 1.8320 2.3360 1.8640 ;
    LAYER V0 ;
      RECT 2.3040 1.8320 2.3360 1.8640 ;
    LAYER V0 ;
      RECT 2.3840 0.4040 2.4160 0.4360 ;
    LAYER V0 ;
      RECT 2.3840 0.5300 2.4160 0.5620 ;
    LAYER V0 ;
      RECT 2.3840 0.6560 2.4160 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.9080 2.4160 0.9400 ;
    LAYER V0 ;
      RECT 2.3840 1.5800 2.4160 1.6120 ;
    LAYER V0 ;
      RECT 2.3840 1.7060 2.4160 1.7380 ;
    LAYER V0 ;
      RECT 2.3840 1.8320 2.4160 1.8640 ;
    LAYER V0 ;
      RECT 2.3840 2.0840 2.4160 2.1160 ;
    LAYER V0 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V0 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.5440 0.4040 2.5760 0.4360 ;
    LAYER V0 ;
      RECT 2.5440 0.5300 2.5760 0.5620 ;
    LAYER V0 ;
      RECT 2.5440 0.6560 2.5760 0.6880 ;
    LAYER V0 ;
      RECT 2.5440 0.9080 2.5760 0.9400 ;
    LAYER V0 ;
      RECT 2.5440 1.5800 2.5760 1.6120 ;
    LAYER V0 ;
      RECT 2.5440 1.7060 2.5760 1.7380 ;
    LAYER V0 ;
      RECT 2.5440 1.8320 2.5760 1.8640 ;
    LAYER V0 ;
      RECT 2.5440 2.0840 2.5760 2.1160 ;
    LAYER V0 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V0 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 1.5800 2.6560 1.6120 ;
    LAYER V0 ;
      RECT 2.6240 1.5800 2.6560 1.6120 ;
    LAYER V0 ;
      RECT 2.6240 1.7060 2.6560 1.7380 ;
    LAYER V0 ;
      RECT 2.6240 1.7060 2.6560 1.7380 ;
    LAYER V0 ;
      RECT 2.6240 1.8320 2.6560 1.8640 ;
    LAYER V0 ;
      RECT 2.6240 1.8320 2.6560 1.8640 ;
    LAYER V0 ;
      RECT 2.7040 0.4040 2.7360 0.4360 ;
    LAYER V0 ;
      RECT 2.7040 0.5300 2.7360 0.5620 ;
    LAYER V0 ;
      RECT 2.7040 0.6560 2.7360 0.6880 ;
    LAYER V0 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V0 ;
      RECT 2.7040 1.5800 2.7360 1.6120 ;
    LAYER V0 ;
      RECT 2.7040 1.7060 2.7360 1.7380 ;
    LAYER V0 ;
      RECT 2.7040 1.8320 2.7360 1.8640 ;
    LAYER V0 ;
      RECT 2.7040 2.0840 2.7360 2.1160 ;
    LAYER V0 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V0 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.7840 1.5800 2.8160 1.6120 ;
    LAYER V0 ;
      RECT 2.7840 1.7060 2.8160 1.7380 ;
    LAYER V0 ;
      RECT 2.7840 1.8320 2.8160 1.8640 ;
  END
END DP_NMOS_B_nfin192_n12_X8_Y2
MACRO Switch_NMOS_B_nfin144_n12_X4_Y3
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin144_n12_X4_Y3 0 0 ;
  SIZE 1.1200 BY 4.2000 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 2.4720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 2.5560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.8880 0.5000 3.3120 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 3.8480 0.8360 3.8800 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.4000 0.3360 3.1440 ;
    LAYER M1 ;
      RECT 0.3040 3.2400 0.3360 3.4800 ;
    LAYER M1 ;
      RECT 0.3040 3.7440 0.3360 3.9840 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.2240 2.4000 0.2560 3.1440 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.4000 0.4160 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.4000 0.4960 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 3.2400 0.4960 3.4800 ;
    LAYER M1 ;
      RECT 0.4640 3.7440 0.4960 3.9840 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 2.4000 0.5760 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.4000 0.6560 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 3.2400 0.6560 3.4800 ;
    LAYER M1 ;
      RECT 0.6240 3.7440 0.6560 3.9840 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.4000 0.7360 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.4000 0.8160 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 3.2400 0.8160 3.4800 ;
    LAYER M1 ;
      RECT 0.7840 3.7440 0.8160 3.9840 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.8640 2.4000 0.8960 3.1440 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.8360 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 0.8360 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.8360 2.1160 ;
    LAYER M2 ;
      RECT 0.2040 2.4200 0.9160 2.4520 ;
    LAYER M2 ;
      RECT 0.2840 2.5040 0.8360 2.5360 ;
    LAYER M2 ;
      RECT 0.2840 3.2600 0.8360 3.2920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 2.4200 0.2560 2.4520 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 2.4200 0.4160 2.4520 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 2.4200 0.5760 2.4520 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 2.4200 0.7360 2.4520 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 2.4200 0.8960 2.4520 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.5040 0.6560 2.5360 ;
    LAYER V1 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V1 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.5040 0.8160 2.5360 ;
    LAYER V1 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V1 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER V1 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V1 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.5040 0.4960 2.5360 ;
    LAYER V1 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V1 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.4200 0.3360 2.4520 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.3840 2.5040 0.4160 2.5360 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V2 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.7560 0.3360 2.7880 ;
    LAYER V0 ;
      RECT 0.3040 2.8820 0.3360 2.9140 ;
    LAYER V0 ;
      RECT 0.3040 3.0080 0.3360 3.0400 ;
    LAYER V0 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.3040 3.8480 0.3360 3.8800 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.2240 2.7560 0.2560 2.7880 ;
    LAYER V0 ;
      RECT 0.2240 2.8820 0.2560 2.9140 ;
    LAYER V0 ;
      RECT 0.2240 3.0080 0.2560 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.7560 0.4960 2.7880 ;
    LAYER V0 ;
      RECT 0.4640 2.8820 0.4960 2.9140 ;
    LAYER V0 ;
      RECT 0.4640 3.0080 0.4960 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.4640 3.8480 0.4960 3.8800 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.7560 0.6560 2.7880 ;
    LAYER V0 ;
      RECT 0.6240 2.8820 0.6560 2.9140 ;
    LAYER V0 ;
      RECT 0.6240 3.0080 0.6560 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.6240 3.8480 0.6560 3.8800 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.7560 0.8160 2.7880 ;
    LAYER V0 ;
      RECT 0.7840 2.8820 0.8160 2.9140 ;
    LAYER V0 ;
      RECT 0.7840 3.0080 0.8160 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.7840 3.8480 0.8160 3.8800 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
  END
END Switch_NMOS_B_nfin144_n12_X4_Y3
MACRO SCM_NMOS_nfin72_nf1_m1_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin72_nf1_m1_n12_X3_Y2 0 0 ;
  SIZE 1.4400 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 2.7240 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 2.1360 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.2160 0.6600 1.4640 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.5680 0.8160 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.2240 0.9760 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 2.0640 0.9760 2.3040 ;
    LAYER M1 ;
      RECT 0.9440 2.5680 0.9760 2.8080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.2240 1.1360 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 2.0640 1.1360 2.3040 ;
    LAYER M1 ;
      RECT 1.1040 2.5680 1.1360 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 1.1560 0.9400 ;
    LAYER M2 ;
      RECT 0.4440 0.2360 1.1560 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.2360 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 2.6720 1.1560 2.7040 ;
    LAYER M2 ;
      RECT 0.4440 1.3280 1.1560 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 1.1560 2.1160 ;
    LAYER M2 ;
      RECT 0.2840 1.4120 0.9960 1.4440 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4120 0.6560 1.4440 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4120 0.9760 1.4440 ;
    LAYER V1 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V1 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4120 0.3360 1.4440 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.3280 1.1360 1.3600 ;
    LAYER V1 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V1 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.2440 0.4960 1.2760 ;
    LAYER V2 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.5440 0.1520 0.5760 0.1840 ;
    LAYER V2 ;
      RECT 0.5440 0.9080 0.5760 0.9400 ;
    LAYER V2 ;
      RECT 0.5440 1.3280 0.5760 1.3600 ;
    LAYER V2 ;
      RECT 0.5440 2.0840 0.5760 2.1160 ;
    LAYER V2 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V2 ;
      RECT 0.6240 1.4120 0.6560 1.4440 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.5800 0.9760 1.6120 ;
    LAYER V0 ;
      RECT 0.9440 1.7060 0.9760 1.7380 ;
    LAYER V0 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.5800 1.1360 1.6120 ;
    LAYER V0 ;
      RECT 1.1040 1.7060 1.1360 1.7380 ;
    LAYER V0 ;
      RECT 1.1040 1.8320 1.1360 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
  END
END SCM_NMOS_nfin72_nf1_m1_n12_X3_Y2
MACRO Switch_NMOS_B_nfin288_n12_X6_Y4
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin288_n12_X6_Y4 0 0 ;
  SIZE 1.4400 BY 5.3760 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 3.6480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 3.7320 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.8880 0.6600 4.4880 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 5.0240 1.1560 5.0560 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.4000 0.3360 3.1440 ;
    LAYER M1 ;
      RECT 0.3040 3.2400 0.3360 3.4800 ;
    LAYER M1 ;
      RECT 0.3040 3.5760 0.3360 4.3200 ;
    LAYER M1 ;
      RECT 0.3040 4.4160 0.3360 4.6560 ;
    LAYER M1 ;
      RECT 0.3040 4.9200 0.3360 5.1600 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.2240 2.4000 0.2560 3.1440 ;
    LAYER M1 ;
      RECT 0.2240 3.5760 0.2560 4.3200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.4000 0.4160 3.1440 ;
    LAYER M1 ;
      RECT 0.3840 3.5760 0.4160 4.3200 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.4000 0.4960 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 3.2400 0.4960 3.4800 ;
    LAYER M1 ;
      RECT 0.4640 3.5760 0.4960 4.3200 ;
    LAYER M1 ;
      RECT 0.4640 4.4160 0.4960 4.6560 ;
    LAYER M1 ;
      RECT 0.4640 4.9200 0.4960 5.1600 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 2.4000 0.5760 3.1440 ;
    LAYER M1 ;
      RECT 0.5440 3.5760 0.5760 4.3200 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.4000 0.6560 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 3.2400 0.6560 3.4800 ;
    LAYER M1 ;
      RECT 0.6240 3.5760 0.6560 4.3200 ;
    LAYER M1 ;
      RECT 0.6240 4.4160 0.6560 4.6560 ;
    LAYER M1 ;
      RECT 0.6240 4.9200 0.6560 5.1600 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.4000 0.7360 3.1440 ;
    LAYER M1 ;
      RECT 0.7040 3.5760 0.7360 4.3200 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.4000 0.8160 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 3.2400 0.8160 3.4800 ;
    LAYER M1 ;
      RECT 0.7840 3.5760 0.8160 4.3200 ;
    LAYER M1 ;
      RECT 0.7840 4.4160 0.8160 4.6560 ;
    LAYER M1 ;
      RECT 0.7840 4.9200 0.8160 5.1600 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.8640 2.4000 0.8960 3.1440 ;
    LAYER M1 ;
      RECT 0.8640 3.5760 0.8960 4.3200 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.2240 0.9760 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 2.0640 0.9760 2.3040 ;
    LAYER M1 ;
      RECT 0.9440 2.4000 0.9760 3.1440 ;
    LAYER M1 ;
      RECT 0.9440 3.2400 0.9760 3.4800 ;
    LAYER M1 ;
      RECT 0.9440 3.5760 0.9760 4.3200 ;
    LAYER M1 ;
      RECT 0.9440 4.4160 0.9760 4.6560 ;
    LAYER M1 ;
      RECT 0.9440 4.9200 0.9760 5.1600 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.4000 1.0560 3.1440 ;
    LAYER M1 ;
      RECT 1.0240 3.5760 1.0560 4.3200 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.2240 1.1360 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 2.0640 1.1360 2.3040 ;
    LAYER M1 ;
      RECT 1.1040 2.4000 1.1360 3.1440 ;
    LAYER M1 ;
      RECT 1.1040 3.2400 1.1360 3.4800 ;
    LAYER M1 ;
      RECT 1.1040 3.5760 1.1360 4.3200 ;
    LAYER M1 ;
      RECT 1.1040 4.4160 1.1360 4.6560 ;
    LAYER M1 ;
      RECT 1.1040 4.9200 1.1360 5.1600 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.1840 2.4000 1.2160 3.1440 ;
    LAYER M1 ;
      RECT 1.1840 3.5760 1.2160 4.3200 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 1.1560 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 1.1560 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.2360 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 1.1560 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 1.1560 2.1160 ;
    LAYER M2 ;
      RECT 0.2040 2.4200 1.2360 2.4520 ;
    LAYER M2 ;
      RECT 0.2840 2.5040 1.1560 2.5360 ;
    LAYER M2 ;
      RECT 0.2840 3.2600 1.1560 3.2920 ;
    LAYER M2 ;
      RECT 0.2040 3.5960 1.2360 3.6280 ;
    LAYER M2 ;
      RECT 0.2840 3.6800 1.1560 3.7120 ;
    LAYER M2 ;
      RECT 0.2840 4.4360 1.1560 4.4680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 2.4200 0.2560 2.4520 ;
    LAYER V1 ;
      RECT 0.2240 3.5960 0.2560 3.6280 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 2.4200 0.4160 2.4520 ;
    LAYER V1 ;
      RECT 0.3840 3.5960 0.4160 3.6280 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 2.4200 0.5760 2.4520 ;
    LAYER V1 ;
      RECT 0.5440 3.5960 0.5760 3.6280 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 2.4200 0.7360 2.4520 ;
    LAYER V1 ;
      RECT 0.7040 3.5960 0.7360 3.6280 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 2.4200 0.8960 2.4520 ;
    LAYER V1 ;
      RECT 0.8640 3.5960 0.8960 3.6280 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V1 ;
      RECT 1.0240 2.4200 1.0560 2.4520 ;
    LAYER V1 ;
      RECT 1.0240 3.5960 1.0560 3.6280 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 2.4200 1.2160 2.4520 ;
    LAYER V1 ;
      RECT 1.1840 3.5960 1.2160 3.6280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER V1 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V1 ;
      RECT 0.3040 3.6800 0.3360 3.7120 ;
    LAYER V1 ;
      RECT 0.3040 4.4360 0.3360 4.4680 ;
    LAYER V1 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.5040 0.4960 2.5360 ;
    LAYER V1 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V1 ;
      RECT 0.4640 3.6800 0.4960 3.7120 ;
    LAYER V1 ;
      RECT 0.4640 4.4360 0.4960 4.4680 ;
    LAYER V1 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.5040 0.6560 2.5360 ;
    LAYER V1 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V1 ;
      RECT 0.6240 3.6800 0.6560 3.7120 ;
    LAYER V1 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V1 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.5040 0.8160 2.5360 ;
    LAYER V1 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V1 ;
      RECT 0.7840 3.6800 0.8160 3.7120 ;
    LAYER V1 ;
      RECT 0.7840 4.4360 0.8160 4.4680 ;
    LAYER V1 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.3280 0.9760 1.3600 ;
    LAYER V1 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V1 ;
      RECT 0.9440 2.5040 0.9760 2.5360 ;
    LAYER V1 ;
      RECT 0.9440 3.2600 0.9760 3.2920 ;
    LAYER V1 ;
      RECT 0.9440 3.6800 0.9760 3.7120 ;
    LAYER V1 ;
      RECT 0.9440 4.4360 0.9760 4.4680 ;
    LAYER V1 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V1 ;
      RECT 1.1040 0.1520 1.1360 0.1840 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.3280 1.1360 1.3600 ;
    LAYER V1 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V1 ;
      RECT 1.1040 2.5040 1.1360 2.5360 ;
    LAYER V1 ;
      RECT 1.1040 3.2600 1.1360 3.2920 ;
    LAYER V1 ;
      RECT 1.1040 3.6800 1.1360 3.7120 ;
    LAYER V1 ;
      RECT 1.1040 4.4360 1.1360 4.4680 ;
    LAYER V1 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.2440 0.4960 1.2760 ;
    LAYER V2 ;
      RECT 0.4640 2.4200 0.4960 2.4520 ;
    LAYER V2 ;
      RECT 0.4640 3.5960 0.4960 3.6280 ;
    LAYER V2 ;
      RECT 0.5440 0.1520 0.5760 0.1840 ;
    LAYER V2 ;
      RECT 0.5440 1.3280 0.5760 1.3600 ;
    LAYER V2 ;
      RECT 0.5440 2.5040 0.5760 2.5360 ;
    LAYER V2 ;
      RECT 0.5440 3.6800 0.5760 3.7120 ;
    LAYER V2 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V2 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V2 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V2 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.7560 0.3360 2.7880 ;
    LAYER V0 ;
      RECT 0.3040 2.8820 0.3360 2.9140 ;
    LAYER V0 ;
      RECT 0.3040 3.0080 0.3360 3.0400 ;
    LAYER V0 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 3.9320 0.3360 3.9640 ;
    LAYER V0 ;
      RECT 0.3040 4.0580 0.3360 4.0900 ;
    LAYER V0 ;
      RECT 0.3040 4.1840 0.3360 4.2160 ;
    LAYER V0 ;
      RECT 0.3040 4.4360 0.3360 4.4680 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.2240 2.7560 0.2560 2.7880 ;
    LAYER V0 ;
      RECT 0.2240 2.8820 0.2560 2.9140 ;
    LAYER V0 ;
      RECT 0.2240 3.0080 0.2560 3.0400 ;
    LAYER V0 ;
      RECT 0.2240 3.9320 0.2560 3.9640 ;
    LAYER V0 ;
      RECT 0.2240 4.0580 0.2560 4.0900 ;
    LAYER V0 ;
      RECT 0.2240 4.1840 0.2560 4.2160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.9320 0.4160 3.9640 ;
    LAYER V0 ;
      RECT 0.3840 3.9320 0.4160 3.9640 ;
    LAYER V0 ;
      RECT 0.3840 4.0580 0.4160 4.0900 ;
    LAYER V0 ;
      RECT 0.3840 4.0580 0.4160 4.0900 ;
    LAYER V0 ;
      RECT 0.3840 4.1840 0.4160 4.2160 ;
    LAYER V0 ;
      RECT 0.3840 4.1840 0.4160 4.2160 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.7560 0.4960 2.7880 ;
    LAYER V0 ;
      RECT 0.4640 2.8820 0.4960 2.9140 ;
    LAYER V0 ;
      RECT 0.4640 3.0080 0.4960 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.4640 3.9320 0.4960 3.9640 ;
    LAYER V0 ;
      RECT 0.4640 4.0580 0.4960 4.0900 ;
    LAYER V0 ;
      RECT 0.4640 4.1840 0.4960 4.2160 ;
    LAYER V0 ;
      RECT 0.4640 4.4360 0.4960 4.4680 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.7560 0.6560 2.7880 ;
    LAYER V0 ;
      RECT 0.6240 2.8820 0.6560 2.9140 ;
    LAYER V0 ;
      RECT 0.6240 3.0080 0.6560 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V0 ;
      RECT 0.6240 3.9320 0.6560 3.9640 ;
    LAYER V0 ;
      RECT 0.6240 4.0580 0.6560 4.0900 ;
    LAYER V0 ;
      RECT 0.6240 4.1840 0.6560 4.2160 ;
    LAYER V0 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.9320 0.7360 3.9640 ;
    LAYER V0 ;
      RECT 0.7040 3.9320 0.7360 3.9640 ;
    LAYER V0 ;
      RECT 0.7040 4.0580 0.7360 4.0900 ;
    LAYER V0 ;
      RECT 0.7040 4.0580 0.7360 4.0900 ;
    LAYER V0 ;
      RECT 0.7040 4.1840 0.7360 4.2160 ;
    LAYER V0 ;
      RECT 0.7040 4.1840 0.7360 4.2160 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.7560 0.8160 2.7880 ;
    LAYER V0 ;
      RECT 0.7840 2.8820 0.8160 2.9140 ;
    LAYER V0 ;
      RECT 0.7840 3.0080 0.8160 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V0 ;
      RECT 0.7840 3.9320 0.8160 3.9640 ;
    LAYER V0 ;
      RECT 0.7840 4.0580 0.8160 4.0900 ;
    LAYER V0 ;
      RECT 0.7840 4.1840 0.8160 4.2160 ;
    LAYER V0 ;
      RECT 0.7840 4.4360 0.8160 4.4680 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.5800 0.9760 1.6120 ;
    LAYER V0 ;
      RECT 0.9440 1.7060 0.9760 1.7380 ;
    LAYER V0 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V0 ;
      RECT 0.9440 2.7560 0.9760 2.7880 ;
    LAYER V0 ;
      RECT 0.9440 2.8820 0.9760 2.9140 ;
    LAYER V0 ;
      RECT 0.9440 3.0080 0.9760 3.0400 ;
    LAYER V0 ;
      RECT 0.9440 3.2600 0.9760 3.2920 ;
    LAYER V0 ;
      RECT 0.9440 3.9320 0.9760 3.9640 ;
    LAYER V0 ;
      RECT 0.9440 4.0580 0.9760 4.0900 ;
    LAYER V0 ;
      RECT 0.9440 4.1840 0.9760 4.2160 ;
    LAYER V0 ;
      RECT 0.9440 4.4360 0.9760 4.4680 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.7560 1.0560 2.7880 ;
    LAYER V0 ;
      RECT 1.0240 2.7560 1.0560 2.7880 ;
    LAYER V0 ;
      RECT 1.0240 2.8820 1.0560 2.9140 ;
    LAYER V0 ;
      RECT 1.0240 2.8820 1.0560 2.9140 ;
    LAYER V0 ;
      RECT 1.0240 3.0080 1.0560 3.0400 ;
    LAYER V0 ;
      RECT 1.0240 3.0080 1.0560 3.0400 ;
    LAYER V0 ;
      RECT 1.0240 3.9320 1.0560 3.9640 ;
    LAYER V0 ;
      RECT 1.0240 3.9320 1.0560 3.9640 ;
    LAYER V0 ;
      RECT 1.0240 4.0580 1.0560 4.0900 ;
    LAYER V0 ;
      RECT 1.0240 4.0580 1.0560 4.0900 ;
    LAYER V0 ;
      RECT 1.0240 4.1840 1.0560 4.2160 ;
    LAYER V0 ;
      RECT 1.0240 4.1840 1.0560 4.2160 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.5800 1.1360 1.6120 ;
    LAYER V0 ;
      RECT 1.1040 1.7060 1.1360 1.7380 ;
    LAYER V0 ;
      RECT 1.1040 1.8320 1.1360 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V0 ;
      RECT 1.1040 2.7560 1.1360 2.7880 ;
    LAYER V0 ;
      RECT 1.1040 2.8820 1.1360 2.9140 ;
    LAYER V0 ;
      RECT 1.1040 3.0080 1.1360 3.0400 ;
    LAYER V0 ;
      RECT 1.1040 3.2600 1.1360 3.2920 ;
    LAYER V0 ;
      RECT 1.1040 3.9320 1.1360 3.9640 ;
    LAYER V0 ;
      RECT 1.1040 4.0580 1.1360 4.0900 ;
    LAYER V0 ;
      RECT 1.1040 4.1840 1.1360 4.2160 ;
    LAYER V0 ;
      RECT 1.1040 4.4360 1.1360 4.4680 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 2.7560 1.2160 2.7880 ;
    LAYER V0 ;
      RECT 1.1840 2.8820 1.2160 2.9140 ;
    LAYER V0 ;
      RECT 1.1840 3.0080 1.2160 3.0400 ;
    LAYER V0 ;
      RECT 1.1840 3.9320 1.2160 3.9640 ;
    LAYER V0 ;
      RECT 1.1840 4.0580 1.2160 4.0900 ;
    LAYER V0 ;
      RECT 1.1840 4.1840 1.2160 4.2160 ;
  END
END Switch_NMOS_B_nfin288_n12_X6_Y4
MACRO DP_NMOS_B_nfin96_n12_X8_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin96_n12_X8_Y1 0 0 ;
  SIZE 3.0400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.8360 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 2.7560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 2.5960 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 2.7560 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.9920 2.5960 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 2.7560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.8880 1.2960 1.1280 ;
    LAYER M1 ;
      RECT 1.2640 1.3920 1.2960 1.6320 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.0480 1.4560 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.8880 1.4560 1.1280 ;
    LAYER M1 ;
      RECT 1.4240 1.3920 1.4560 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.3920 1.6160 1.6320 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.0480 1.7760 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.8880 1.7760 1.1280 ;
    LAYER M1 ;
      RECT 1.7440 1.3920 1.7760 1.6320 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.8880 1.9360 1.1280 ;
    LAYER M1 ;
      RECT 1.9040 1.3920 1.9360 1.6320 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.0480 2.0960 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.8880 2.0960 1.1280 ;
    LAYER M1 ;
      RECT 2.0640 1.3920 2.0960 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.3920 2.2560 1.6320 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.0480 2.4160 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.8880 2.4160 1.1280 ;
    LAYER M1 ;
      RECT 2.3840 1.3920 2.4160 1.6320 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER M1 ;
      RECT 2.5440 0.0480 2.5760 0.7920 ;
    LAYER M1 ;
      RECT 2.5440 0.8880 2.5760 1.1280 ;
    LAYER M1 ;
      RECT 2.5440 1.3920 2.5760 1.6320 ;
    LAYER M1 ;
      RECT 2.6240 0.0480 2.6560 0.7920 ;
    LAYER M1 ;
      RECT 2.7040 0.0480 2.7360 0.7920 ;
    LAYER M1 ;
      RECT 2.7040 0.8880 2.7360 1.1280 ;
    LAYER M1 ;
      RECT 2.7040 1.3920 2.7360 1.6320 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER V1 ;
      RECT 2.6240 0.0680 2.6560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.3440 0.0680 1.3760 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.9840 0.0680 2.0160 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 2.7040 0.1520 2.7360 0.1840 ;
    LAYER V1 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V1 ;
      RECT 2.7040 1.4960 2.7360 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 1.4240 0.1520 1.4560 0.1840 ;
    LAYER V1 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V1 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V1 ;
      RECT 1.5840 0.1520 1.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V1 ;
      RECT 2.0640 0.1520 2.0960 0.1840 ;
    LAYER V1 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V1 ;
      RECT 2.0640 1.4960 2.0960 1.5280 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V1 ;
      RECT 2.5440 0.2360 2.5760 0.2680 ;
    LAYER V1 ;
      RECT 2.5440 0.9920 2.5760 1.0240 ;
    LAYER V1 ;
      RECT 2.5440 1.4960 2.5760 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9920 0.6560 1.0240 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V1 ;
      RECT 1.2640 0.2360 1.2960 0.2680 ;
    LAYER V1 ;
      RECT 1.2640 0.9920 1.2960 1.0240 ;
    LAYER V1 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V1 ;
      RECT 1.7440 0.2360 1.7760 0.2680 ;
    LAYER V1 ;
      RECT 1.7440 0.9920 1.7760 1.0240 ;
    LAYER V1 ;
      RECT 1.7440 1.4960 1.7760 1.5280 ;
    LAYER V1 ;
      RECT 1.9040 0.2360 1.9360 0.2680 ;
    LAYER V1 ;
      RECT 1.9040 0.9920 1.9360 1.0240 ;
    LAYER V1 ;
      RECT 1.9040 1.4960 1.9360 1.5280 ;
    LAYER V1 ;
      RECT 2.3840 0.2360 2.4160 0.2680 ;
    LAYER V1 ;
      RECT 2.3840 0.9920 2.4160 1.0240 ;
    LAYER V1 ;
      RECT 2.3840 1.4960 2.4160 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.4040 1.2960 0.4360 ;
    LAYER V0 ;
      RECT 1.2640 0.5300 1.2960 0.5620 ;
    LAYER V0 ;
      RECT 1.2640 0.6560 1.2960 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V0 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.4040 1.4560 0.4360 ;
    LAYER V0 ;
      RECT 1.4240 0.5300 1.4560 0.5620 ;
    LAYER V0 ;
      RECT 1.4240 0.6560 1.4560 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V0 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.4040 1.7760 0.4360 ;
    LAYER V0 ;
      RECT 1.7440 0.5300 1.7760 0.5620 ;
    LAYER V0 ;
      RECT 1.7440 0.6560 1.7760 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.9080 1.7760 0.9400 ;
    LAYER V0 ;
      RECT 1.7440 1.4960 1.7760 1.5280 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.4040 1.9360 0.4360 ;
    LAYER V0 ;
      RECT 1.9040 0.5300 1.9360 0.5620 ;
    LAYER V0 ;
      RECT 1.9040 0.6560 1.9360 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.9080 1.9360 0.9400 ;
    LAYER V0 ;
      RECT 1.9040 1.4960 1.9360 1.5280 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.4040 2.0960 0.4360 ;
    LAYER V0 ;
      RECT 2.0640 0.5300 2.0960 0.5620 ;
    LAYER V0 ;
      RECT 2.0640 0.6560 2.0960 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V0 ;
      RECT 2.0640 1.4960 2.0960 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.4040 2.4160 0.4360 ;
    LAYER V0 ;
      RECT 2.3840 0.5300 2.4160 0.5620 ;
    LAYER V0 ;
      RECT 2.3840 0.6560 2.4160 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.9080 2.4160 0.9400 ;
    LAYER V0 ;
      RECT 2.3840 1.4960 2.4160 1.5280 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.5440 0.4040 2.5760 0.4360 ;
    LAYER V0 ;
      RECT 2.5440 0.5300 2.5760 0.5620 ;
    LAYER V0 ;
      RECT 2.5440 0.6560 2.5760 0.6880 ;
    LAYER V0 ;
      RECT 2.5440 0.9080 2.5760 0.9400 ;
    LAYER V0 ;
      RECT 2.5440 1.4960 2.5760 1.5280 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.7040 0.4040 2.7360 0.4360 ;
    LAYER V0 ;
      RECT 2.7040 0.5300 2.7360 0.5620 ;
    LAYER V0 ;
      RECT 2.7040 0.6560 2.7360 0.6880 ;
    LAYER V0 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V0 ;
      RECT 2.7040 1.4960 2.7360 1.5280 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
  END
END DP_NMOS_B_nfin96_n12_X8_Y1
MACRO Res_r400
  ORIGIN 0 0 ;
  FOREIGN Res_r400 0 0 ;
  SIZE 1.0400 BY 1.7640 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.3560 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6040 0.0680 0.9320 0.1000 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 1.7160 ;
    LAYER M1 ;
      RECT 0.3040 1.6640 0.4000 1.6960 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 1.7160 ;
    LAYER M1 ;
      RECT 0.3680 0.0680 0.4640 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 1.7160 ;
    LAYER M1 ;
      RECT 0.4320 1.6640 0.5280 1.6960 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 1.7160 ;
    LAYER M1 ;
      RECT 0.4960 0.0680 0.5920 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 1.7160 ;
    LAYER M1 ;
      RECT 0.5600 1.6640 0.6560 1.6960 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 1.7160 ;
    LAYER V1 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
  END
END Res_r400
MACRO Switch_NMOS_nfin288_n12_X6_Y4
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin288_n12_X6_Y4 0 0 ;
  SIZE 1.4400 BY 5.3760 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 5.0760 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 3.7320 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.8880 0.6600 4.4880 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.4000 0.3360 3.1440 ;
    LAYER M1 ;
      RECT 0.3040 3.2400 0.3360 3.4800 ;
    LAYER M1 ;
      RECT 0.3040 3.5760 0.3360 4.3200 ;
    LAYER M1 ;
      RECT 0.3040 4.4160 0.3360 4.6560 ;
    LAYER M1 ;
      RECT 0.3040 4.9200 0.3360 5.1600 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.2240 2.4000 0.2560 3.1440 ;
    LAYER M1 ;
      RECT 0.2240 3.5760 0.2560 4.3200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.4000 0.4160 3.1440 ;
    LAYER M1 ;
      RECT 0.3840 3.5760 0.4160 4.3200 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.4000 0.4960 3.1440 ;
    LAYER M1 ;
      RECT 0.4640 3.2400 0.4960 3.4800 ;
    LAYER M1 ;
      RECT 0.4640 3.5760 0.4960 4.3200 ;
    LAYER M1 ;
      RECT 0.4640 4.4160 0.4960 4.6560 ;
    LAYER M1 ;
      RECT 0.4640 4.9200 0.4960 5.1600 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 2.4000 0.5760 3.1440 ;
    LAYER M1 ;
      RECT 0.5440 3.5760 0.5760 4.3200 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.4000 0.6560 3.1440 ;
    LAYER M1 ;
      RECT 0.6240 3.2400 0.6560 3.4800 ;
    LAYER M1 ;
      RECT 0.6240 3.5760 0.6560 4.3200 ;
    LAYER M1 ;
      RECT 0.6240 4.4160 0.6560 4.6560 ;
    LAYER M1 ;
      RECT 0.6240 4.9200 0.6560 5.1600 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.4000 0.7360 3.1440 ;
    LAYER M1 ;
      RECT 0.7040 3.5760 0.7360 4.3200 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.4000 0.8160 3.1440 ;
    LAYER M1 ;
      RECT 0.7840 3.2400 0.8160 3.4800 ;
    LAYER M1 ;
      RECT 0.7840 3.5760 0.8160 4.3200 ;
    LAYER M1 ;
      RECT 0.7840 4.4160 0.8160 4.6560 ;
    LAYER M1 ;
      RECT 0.7840 4.9200 0.8160 5.1600 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.8640 2.4000 0.8960 3.1440 ;
    LAYER M1 ;
      RECT 0.8640 3.5760 0.8960 4.3200 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.2240 0.9760 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 2.0640 0.9760 2.3040 ;
    LAYER M1 ;
      RECT 0.9440 2.4000 0.9760 3.1440 ;
    LAYER M1 ;
      RECT 0.9440 3.2400 0.9760 3.4800 ;
    LAYER M1 ;
      RECT 0.9440 3.5760 0.9760 4.3200 ;
    LAYER M1 ;
      RECT 0.9440 4.4160 0.9760 4.6560 ;
    LAYER M1 ;
      RECT 0.9440 4.9200 0.9760 5.1600 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.4000 1.0560 3.1440 ;
    LAYER M1 ;
      RECT 1.0240 3.5760 1.0560 4.3200 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.2240 1.1360 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 2.0640 1.1360 2.3040 ;
    LAYER M1 ;
      RECT 1.1040 2.4000 1.1360 3.1440 ;
    LAYER M1 ;
      RECT 1.1040 3.2400 1.1360 3.4800 ;
    LAYER M1 ;
      RECT 1.1040 3.5760 1.1360 4.3200 ;
    LAYER M1 ;
      RECT 1.1040 4.4160 1.1360 4.6560 ;
    LAYER M1 ;
      RECT 1.1040 4.9200 1.1360 5.1600 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.1840 2.4000 1.2160 3.1440 ;
    LAYER M1 ;
      RECT 1.1840 3.5760 1.2160 4.3200 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 1.1560 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 1.1560 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.2360 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 1.1560 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 1.1560 2.1160 ;
    LAYER M2 ;
      RECT 0.2040 2.4200 1.2360 2.4520 ;
    LAYER M2 ;
      RECT 0.2840 2.5040 1.1560 2.5360 ;
    LAYER M2 ;
      RECT 0.2840 3.2600 1.1560 3.2920 ;
    LAYER M2 ;
      RECT 0.2040 3.5960 1.2360 3.6280 ;
    LAYER M2 ;
      RECT 0.2840 5.0240 1.1560 5.0560 ;
    LAYER M2 ;
      RECT 0.2840 3.6800 1.1560 3.7120 ;
    LAYER M2 ;
      RECT 0.2840 4.4360 1.1560 4.4680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 2.4200 0.2560 2.4520 ;
    LAYER V1 ;
      RECT 0.2240 3.5960 0.2560 3.6280 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 2.4200 0.4160 2.4520 ;
    LAYER V1 ;
      RECT 0.3840 3.5960 0.4160 3.6280 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 2.4200 0.5760 2.4520 ;
    LAYER V1 ;
      RECT 0.5440 3.5960 0.5760 3.6280 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 2.4200 0.7360 2.4520 ;
    LAYER V1 ;
      RECT 0.7040 3.5960 0.7360 3.6280 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 2.4200 0.8960 2.4520 ;
    LAYER V1 ;
      RECT 0.8640 3.5960 0.8960 3.6280 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V1 ;
      RECT 1.0240 2.4200 1.0560 2.4520 ;
    LAYER V1 ;
      RECT 1.0240 3.5960 1.0560 3.6280 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 2.4200 1.2160 2.4520 ;
    LAYER V1 ;
      RECT 1.1840 3.5960 1.2160 3.6280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER V1 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V1 ;
      RECT 0.3040 3.6800 0.3360 3.7120 ;
    LAYER V1 ;
      RECT 0.3040 4.4360 0.3360 4.4680 ;
    LAYER V1 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.5040 0.4960 2.5360 ;
    LAYER V1 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V1 ;
      RECT 0.4640 3.6800 0.4960 3.7120 ;
    LAYER V1 ;
      RECT 0.4640 4.4360 0.4960 4.4680 ;
    LAYER V1 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.5040 0.6560 2.5360 ;
    LAYER V1 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V1 ;
      RECT 0.6240 3.6800 0.6560 3.7120 ;
    LAYER V1 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V1 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.5040 0.8160 2.5360 ;
    LAYER V1 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V1 ;
      RECT 0.7840 3.6800 0.8160 3.7120 ;
    LAYER V1 ;
      RECT 0.7840 4.4360 0.8160 4.4680 ;
    LAYER V1 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.3280 0.9760 1.3600 ;
    LAYER V1 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V1 ;
      RECT 0.9440 2.5040 0.9760 2.5360 ;
    LAYER V1 ;
      RECT 0.9440 3.2600 0.9760 3.2920 ;
    LAYER V1 ;
      RECT 0.9440 3.6800 0.9760 3.7120 ;
    LAYER V1 ;
      RECT 0.9440 4.4360 0.9760 4.4680 ;
    LAYER V1 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V1 ;
      RECT 1.1040 0.1520 1.1360 0.1840 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.3280 1.1360 1.3600 ;
    LAYER V1 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V1 ;
      RECT 1.1040 2.5040 1.1360 2.5360 ;
    LAYER V1 ;
      RECT 1.1040 3.2600 1.1360 3.2920 ;
    LAYER V1 ;
      RECT 1.1040 3.6800 1.1360 3.7120 ;
    LAYER V1 ;
      RECT 1.1040 4.4360 1.1360 4.4680 ;
    LAYER V1 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.2440 0.4960 1.2760 ;
    LAYER V2 ;
      RECT 0.4640 2.4200 0.4960 2.4520 ;
    LAYER V2 ;
      RECT 0.4640 3.5960 0.4960 3.6280 ;
    LAYER V2 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V2 ;
      RECT 0.5440 0.1520 0.5760 0.1840 ;
    LAYER V2 ;
      RECT 0.5440 1.3280 0.5760 1.3600 ;
    LAYER V2 ;
      RECT 0.5440 2.5040 0.5760 2.5360 ;
    LAYER V2 ;
      RECT 0.5440 3.6800 0.5760 3.7120 ;
    LAYER V2 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V2 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V2 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V2 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.7560 0.3360 2.7880 ;
    LAYER V0 ;
      RECT 0.3040 2.8820 0.3360 2.9140 ;
    LAYER V0 ;
      RECT 0.3040 3.0080 0.3360 3.0400 ;
    LAYER V0 ;
      RECT 0.3040 3.2600 0.3360 3.2920 ;
    LAYER V0 ;
      RECT 0.3040 3.9320 0.3360 3.9640 ;
    LAYER V0 ;
      RECT 0.3040 4.0580 0.3360 4.0900 ;
    LAYER V0 ;
      RECT 0.3040 4.1840 0.3360 4.2160 ;
    LAYER V0 ;
      RECT 0.3040 4.4360 0.3360 4.4680 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.3040 5.0240 0.3360 5.0560 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.2240 2.7560 0.2560 2.7880 ;
    LAYER V0 ;
      RECT 0.2240 2.8820 0.2560 2.9140 ;
    LAYER V0 ;
      RECT 0.2240 3.0080 0.2560 3.0400 ;
    LAYER V0 ;
      RECT 0.2240 3.9320 0.2560 3.9640 ;
    LAYER V0 ;
      RECT 0.2240 4.0580 0.2560 4.0900 ;
    LAYER V0 ;
      RECT 0.2240 4.1840 0.2560 4.2160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.9320 0.4160 3.9640 ;
    LAYER V0 ;
      RECT 0.3840 3.9320 0.4160 3.9640 ;
    LAYER V0 ;
      RECT 0.3840 4.0580 0.4160 4.0900 ;
    LAYER V0 ;
      RECT 0.3840 4.0580 0.4160 4.0900 ;
    LAYER V0 ;
      RECT 0.3840 4.1840 0.4160 4.2160 ;
    LAYER V0 ;
      RECT 0.3840 4.1840 0.4160 4.2160 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.7560 0.4960 2.7880 ;
    LAYER V0 ;
      RECT 0.4640 2.8820 0.4960 2.9140 ;
    LAYER V0 ;
      RECT 0.4640 3.0080 0.4960 3.0400 ;
    LAYER V0 ;
      RECT 0.4640 3.2600 0.4960 3.2920 ;
    LAYER V0 ;
      RECT 0.4640 3.9320 0.4960 3.9640 ;
    LAYER V0 ;
      RECT 0.4640 4.0580 0.4960 4.0900 ;
    LAYER V0 ;
      RECT 0.4640 4.1840 0.4960 4.2160 ;
    LAYER V0 ;
      RECT 0.4640 4.4360 0.4960 4.4680 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.4640 5.0240 0.4960 5.0560 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.7560 0.6560 2.7880 ;
    LAYER V0 ;
      RECT 0.6240 2.8820 0.6560 2.9140 ;
    LAYER V0 ;
      RECT 0.6240 3.0080 0.6560 3.0400 ;
    LAYER V0 ;
      RECT 0.6240 3.2600 0.6560 3.2920 ;
    LAYER V0 ;
      RECT 0.6240 3.9320 0.6560 3.9640 ;
    LAYER V0 ;
      RECT 0.6240 4.0580 0.6560 4.0900 ;
    LAYER V0 ;
      RECT 0.6240 4.1840 0.6560 4.2160 ;
    LAYER V0 ;
      RECT 0.6240 4.4360 0.6560 4.4680 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.6240 5.0240 0.6560 5.0560 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.9320 0.7360 3.9640 ;
    LAYER V0 ;
      RECT 0.7040 3.9320 0.7360 3.9640 ;
    LAYER V0 ;
      RECT 0.7040 4.0580 0.7360 4.0900 ;
    LAYER V0 ;
      RECT 0.7040 4.0580 0.7360 4.0900 ;
    LAYER V0 ;
      RECT 0.7040 4.1840 0.7360 4.2160 ;
    LAYER V0 ;
      RECT 0.7040 4.1840 0.7360 4.2160 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.7560 0.8160 2.7880 ;
    LAYER V0 ;
      RECT 0.7840 2.8820 0.8160 2.9140 ;
    LAYER V0 ;
      RECT 0.7840 3.0080 0.8160 3.0400 ;
    LAYER V0 ;
      RECT 0.7840 3.2600 0.8160 3.2920 ;
    LAYER V0 ;
      RECT 0.7840 3.9320 0.8160 3.9640 ;
    LAYER V0 ;
      RECT 0.7840 4.0580 0.8160 4.0900 ;
    LAYER V0 ;
      RECT 0.7840 4.1840 0.8160 4.2160 ;
    LAYER V0 ;
      RECT 0.7840 4.4360 0.8160 4.4680 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.5800 0.9760 1.6120 ;
    LAYER V0 ;
      RECT 0.9440 1.7060 0.9760 1.7380 ;
    LAYER V0 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V0 ;
      RECT 0.9440 2.7560 0.9760 2.7880 ;
    LAYER V0 ;
      RECT 0.9440 2.8820 0.9760 2.9140 ;
    LAYER V0 ;
      RECT 0.9440 3.0080 0.9760 3.0400 ;
    LAYER V0 ;
      RECT 0.9440 3.2600 0.9760 3.2920 ;
    LAYER V0 ;
      RECT 0.9440 3.9320 0.9760 3.9640 ;
    LAYER V0 ;
      RECT 0.9440 4.0580 0.9760 4.0900 ;
    LAYER V0 ;
      RECT 0.9440 4.1840 0.9760 4.2160 ;
    LAYER V0 ;
      RECT 0.9440 4.4360 0.9760 4.4680 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 0.9440 5.0240 0.9760 5.0560 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.7560 1.0560 2.7880 ;
    LAYER V0 ;
      RECT 1.0240 2.7560 1.0560 2.7880 ;
    LAYER V0 ;
      RECT 1.0240 2.8820 1.0560 2.9140 ;
    LAYER V0 ;
      RECT 1.0240 2.8820 1.0560 2.9140 ;
    LAYER V0 ;
      RECT 1.0240 3.0080 1.0560 3.0400 ;
    LAYER V0 ;
      RECT 1.0240 3.0080 1.0560 3.0400 ;
    LAYER V0 ;
      RECT 1.0240 3.9320 1.0560 3.9640 ;
    LAYER V0 ;
      RECT 1.0240 3.9320 1.0560 3.9640 ;
    LAYER V0 ;
      RECT 1.0240 4.0580 1.0560 4.0900 ;
    LAYER V0 ;
      RECT 1.0240 4.0580 1.0560 4.0900 ;
    LAYER V0 ;
      RECT 1.0240 4.1840 1.0560 4.2160 ;
    LAYER V0 ;
      RECT 1.0240 4.1840 1.0560 4.2160 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.5800 1.1360 1.6120 ;
    LAYER V0 ;
      RECT 1.1040 1.7060 1.1360 1.7380 ;
    LAYER V0 ;
      RECT 1.1040 1.8320 1.1360 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V0 ;
      RECT 1.1040 2.7560 1.1360 2.7880 ;
    LAYER V0 ;
      RECT 1.1040 2.8820 1.1360 2.9140 ;
    LAYER V0 ;
      RECT 1.1040 3.0080 1.1360 3.0400 ;
    LAYER V0 ;
      RECT 1.1040 3.2600 1.1360 3.2920 ;
    LAYER V0 ;
      RECT 1.1040 3.9320 1.1360 3.9640 ;
    LAYER V0 ;
      RECT 1.1040 4.0580 1.1360 4.0900 ;
    LAYER V0 ;
      RECT 1.1040 4.1840 1.1360 4.2160 ;
    LAYER V0 ;
      RECT 1.1040 4.4360 1.1360 4.4680 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1040 5.0240 1.1360 5.0560 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 2.7560 1.2160 2.7880 ;
    LAYER V0 ;
      RECT 1.1840 2.8820 1.2160 2.9140 ;
    LAYER V0 ;
      RECT 1.1840 3.0080 1.2160 3.0400 ;
    LAYER V0 ;
      RECT 1.1840 3.9320 1.2160 3.9640 ;
    LAYER V0 ;
      RECT 1.1840 4.0580 1.2160 4.0900 ;
    LAYER V0 ;
      RECT 1.1840 4.1840 1.2160 4.2160 ;
  END
END Switch_NMOS_nfin288_n12_X6_Y4
MACRO Switch_NMOS_B_nfin72_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin72_n12_X3_Y2 0 0 ;
  SIZE 0.9600 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 1.2960 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.1320 0.3400 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.8880 0.4200 2.1360 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 0.6760 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.6760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.6760 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.7560 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 0.6760 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.6760 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V2 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V2 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V2 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V2 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
  END
END Switch_NMOS_B_nfin72_n12_X3_Y2
