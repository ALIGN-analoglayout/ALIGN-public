MACRO Switch_NMOS_nfin12_m1_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin12_m1_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_nfin12_m1_n12_X1_Y1
MACRO Switch_PMOS_nfin12_m1_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin12_m1_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_nfin12_m1_n12_X1_Y1
MACRO DP_NMOS_B_nfin12_m16_n12_X8_Y2
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin12_m16_n12_X8_Y2 0 0 ;
  SIZE 3.0400 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1800 0.0480 1.2200 1.2960 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2600 0.1320 1.3000 1.3800 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3400 0.2160 1.3800 1.4640 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4200 0.8880 1.4600 2.1360 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5000 0.9720 1.5400 2.2200 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 2.7560 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.5680 0.8160 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.2240 0.9760 1.9680 ;
    LAYER M1 ;
      RECT 0.9440 2.0640 0.9760 2.3040 ;
    LAYER M1 ;
      RECT 0.9440 2.5680 0.9760 2.8080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.2240 1.1360 1.9680 ;
    LAYER M1 ;
      RECT 1.1040 2.0640 1.1360 2.3040 ;
    LAYER M1 ;
      RECT 1.1040 2.5680 1.1360 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.8880 1.2960 1.1280 ;
    LAYER M1 ;
      RECT 1.2640 1.2240 1.2960 1.9680 ;
    LAYER M1 ;
      RECT 1.2640 2.0640 1.2960 2.3040 ;
    LAYER M1 ;
      RECT 1.2640 2.5680 1.2960 2.8080 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.4240 0.0480 1.4560 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.8880 1.4560 1.1280 ;
    LAYER M1 ;
      RECT 1.4240 1.2240 1.4560 1.9680 ;
    LAYER M1 ;
      RECT 1.4240 2.0640 1.4560 2.3040 ;
    LAYER M1 ;
      RECT 1.4240 2.5680 1.4560 2.8080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.2240 1.6160 1.9680 ;
    LAYER M1 ;
      RECT 1.5840 2.0640 1.6160 2.3040 ;
    LAYER M1 ;
      RECT 1.5840 2.5680 1.6160 2.8080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 1.2240 1.6960 1.9680 ;
    LAYER M1 ;
      RECT 1.7440 0.0480 1.7760 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.8880 1.7760 1.1280 ;
    LAYER M1 ;
      RECT 1.7440 1.2240 1.7760 1.9680 ;
    LAYER M1 ;
      RECT 1.7440 2.0640 1.7760 2.3040 ;
    LAYER M1 ;
      RECT 1.7440 2.5680 1.7760 2.8080 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.8240 1.2240 1.8560 1.9680 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.8880 1.9360 1.1280 ;
    LAYER M1 ;
      RECT 1.9040 1.2240 1.9360 1.9680 ;
    LAYER M1 ;
      RECT 1.9040 2.0640 1.9360 2.3040 ;
    LAYER M1 ;
      RECT 1.9040 2.5680 1.9360 2.8080 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 1.9840 1.2240 2.0160 1.9680 ;
    LAYER M1 ;
      RECT 2.0640 0.0480 2.0960 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.8880 2.0960 1.1280 ;
    LAYER M1 ;
      RECT 2.0640 1.2240 2.0960 1.9680 ;
    LAYER M1 ;
      RECT 2.0640 2.0640 2.0960 2.3040 ;
    LAYER M1 ;
      RECT 2.0640 2.5680 2.0960 2.8080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.1440 1.2240 2.1760 1.9680 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.2240 2.2560 1.9680 ;
    LAYER M1 ;
      RECT 2.2240 2.0640 2.2560 2.3040 ;
    LAYER M1 ;
      RECT 2.2240 2.5680 2.2560 2.8080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 1.2240 2.3360 1.9680 ;
    LAYER M1 ;
      RECT 2.3840 0.0480 2.4160 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.8880 2.4160 1.1280 ;
    LAYER M1 ;
      RECT 2.3840 1.2240 2.4160 1.9680 ;
    LAYER M1 ;
      RECT 2.3840 2.0640 2.4160 2.3040 ;
    LAYER M1 ;
      RECT 2.3840 2.5680 2.4160 2.8080 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER M1 ;
      RECT 2.4640 1.2240 2.4960 1.9680 ;
    LAYER M1 ;
      RECT 2.5440 0.0480 2.5760 0.7920 ;
    LAYER M1 ;
      RECT 2.5440 0.8880 2.5760 1.1280 ;
    LAYER M1 ;
      RECT 2.5440 1.2240 2.5760 1.9680 ;
    LAYER M1 ;
      RECT 2.5440 2.0640 2.5760 2.3040 ;
    LAYER M1 ;
      RECT 2.5440 2.5680 2.5760 2.8080 ;
    LAYER M1 ;
      RECT 2.6240 0.0480 2.6560 0.7920 ;
    LAYER M1 ;
      RECT 2.6240 1.2240 2.6560 1.9680 ;
    LAYER M1 ;
      RECT 2.7040 0.0480 2.7360 0.7920 ;
    LAYER M1 ;
      RECT 2.7040 0.8880 2.7360 1.1280 ;
    LAYER M1 ;
      RECT 2.7040 1.2240 2.7360 1.9680 ;
    LAYER M1 ;
      RECT 2.7040 2.0640 2.7360 2.3040 ;
    LAYER M1 ;
      RECT 2.7040 2.5680 2.7360 2.8080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER M1 ;
      RECT 2.7840 1.2240 2.8160 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 2.7560 0.1840 ;
    LAYER M2 ;
      RECT 0.4440 0.2360 2.5960 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 2.7560 0.9400 ;
    LAYER M2 ;
      RECT 0.4440 0.9920 2.5960 1.0240 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 2.8360 1.2760 ;
    LAYER M2 ;
      RECT 0.4440 1.3280 2.5960 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 1.4120 2.7560 1.4440 ;
    LAYER M2 ;
      RECT 0.4440 2.0840 2.5960 2.1160 ;
    LAYER M2 ;
      RECT 0.2840 2.1680 2.7560 2.2000 ;
    LAYER V1 ;
      RECT 2.6240 0.0680 2.6560 0.1000 ;
    LAYER V1 ;
      RECT 2.6240 1.2440 2.6560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 1.2440 2.8160 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.3440 0.0680 1.3760 0.1000 ;
    LAYER V1 ;
      RECT 1.3440 1.2440 1.3760 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 1.2440 1.6960 1.2760 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 1.2440 1.8560 1.2760 ;
    LAYER V1 ;
      RECT 1.9840 0.0680 2.0160 0.1000 ;
    LAYER V1 ;
      RECT 1.9840 1.2440 2.0160 1.2760 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 1.2440 2.1760 1.2760 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 1.2440 2.3360 1.2760 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 1.2440 2.4960 1.2760 ;
    LAYER V1 ;
      RECT 2.7040 0.1520 2.7360 0.1840 ;
    LAYER V1 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V1 ;
      RECT 2.7040 1.4120 2.7360 1.4440 ;
    LAYER V1 ;
      RECT 2.7040 2.1680 2.7360 2.2000 ;
    LAYER V1 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4120 0.3360 1.4440 ;
    LAYER V1 ;
      RECT 0.3040 2.1680 0.3360 2.2000 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4120 0.8160 1.4440 ;
    LAYER V1 ;
      RECT 0.7840 2.1680 0.8160 2.2000 ;
    LAYER V1 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4120 0.9760 1.4440 ;
    LAYER V1 ;
      RECT 0.9440 2.1680 0.9760 2.2000 ;
    LAYER V1 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V1 ;
      RECT 1.4240 0.1520 1.4560 0.1840 ;
    LAYER V1 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V1 ;
      RECT 1.4240 1.4120 1.4560 1.4440 ;
    LAYER V1 ;
      RECT 1.4240 2.1680 1.4560 2.2000 ;
    LAYER V1 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V1 ;
      RECT 1.5840 0.1520 1.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4120 1.6160 1.4440 ;
    LAYER V1 ;
      RECT 1.5840 2.1680 1.6160 2.2000 ;
    LAYER V1 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V1 ;
      RECT 2.0640 0.1520 2.0960 0.1840 ;
    LAYER V1 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V1 ;
      RECT 2.0640 1.4120 2.0960 1.4440 ;
    LAYER V1 ;
      RECT 2.0640 2.1680 2.0960 2.2000 ;
    LAYER V1 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.2240 1.4120 2.2560 1.4440 ;
    LAYER V1 ;
      RECT 2.2240 2.1680 2.2560 2.2000 ;
    LAYER V1 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V1 ;
      RECT 2.5440 0.2360 2.5760 0.2680 ;
    LAYER V1 ;
      RECT 2.5440 0.9920 2.5760 1.0240 ;
    LAYER V1 ;
      RECT 2.5440 1.3280 2.5760 1.3600 ;
    LAYER V1 ;
      RECT 2.5440 2.0840 2.5760 2.1160 ;
    LAYER V1 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9920 0.6560 1.0240 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.3280 1.1360 1.3600 ;
    LAYER V1 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V1 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V1 ;
      RECT 1.2640 0.2360 1.2960 0.2680 ;
    LAYER V1 ;
      RECT 1.2640 0.9920 1.2960 1.0240 ;
    LAYER V1 ;
      RECT 1.2640 1.3280 1.2960 1.3600 ;
    LAYER V1 ;
      RECT 1.2640 2.0840 1.2960 2.1160 ;
    LAYER V1 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V1 ;
      RECT 1.7440 0.2360 1.7760 0.2680 ;
    LAYER V1 ;
      RECT 1.7440 0.9920 1.7760 1.0240 ;
    LAYER V1 ;
      RECT 1.7440 1.3280 1.7760 1.3600 ;
    LAYER V1 ;
      RECT 1.7440 2.0840 1.7760 2.1160 ;
    LAYER V1 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V1 ;
      RECT 1.9040 0.2360 1.9360 0.2680 ;
    LAYER V1 ;
      RECT 1.9040 0.9920 1.9360 1.0240 ;
    LAYER V1 ;
      RECT 1.9040 1.3280 1.9360 1.3600 ;
    LAYER V1 ;
      RECT 1.9040 2.0840 1.9360 2.1160 ;
    LAYER V1 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V1 ;
      RECT 2.3840 0.2360 2.4160 0.2680 ;
    LAYER V1 ;
      RECT 2.3840 0.9920 2.4160 1.0240 ;
    LAYER V1 ;
      RECT 2.3840 1.3280 2.4160 1.3600 ;
    LAYER V1 ;
      RECT 2.3840 2.0840 2.4160 2.1160 ;
    LAYER V1 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V2 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V2 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V2 ;
      RECT 1.2640 0.1520 1.2960 0.1840 ;
    LAYER V2 ;
      RECT 1.2640 1.3280 1.2960 1.3600 ;
    LAYER V2 ;
      RECT 1.3440 0.2360 1.3760 0.2680 ;
    LAYER V2 ;
      RECT 1.3440 1.4120 1.3760 1.4440 ;
    LAYER V2 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V2 ;
      RECT 1.4240 2.0840 1.4560 2.1160 ;
    LAYER V2 ;
      RECT 1.5040 0.9920 1.5360 1.0240 ;
    LAYER V2 ;
      RECT 1.5040 2.1680 1.5360 2.2000 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.5800 0.9760 1.6120 ;
    LAYER V0 ;
      RECT 0.9440 1.7060 0.9760 1.7380 ;
    LAYER V0 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V0 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 0.9440 2.6720 0.9760 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.5800 1.1360 1.6120 ;
    LAYER V0 ;
      RECT 1.1040 1.7060 1.1360 1.7380 ;
    LAYER V0 ;
      RECT 1.1040 1.8320 1.1360 1.8640 ;
    LAYER V0 ;
      RECT 1.1040 2.0840 1.1360 2.1160 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1040 2.6720 1.1360 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.2640 0.4040 1.2960 0.4360 ;
    LAYER V0 ;
      RECT 1.2640 0.5300 1.2960 0.5620 ;
    LAYER V0 ;
      RECT 1.2640 0.6560 1.2960 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V0 ;
      RECT 1.2640 1.5800 1.2960 1.6120 ;
    LAYER V0 ;
      RECT 1.2640 1.7060 1.2960 1.7380 ;
    LAYER V0 ;
      RECT 1.2640 1.8320 1.2960 1.8640 ;
    LAYER V0 ;
      RECT 1.2640 2.0840 1.2960 2.1160 ;
    LAYER V0 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V0 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.4240 0.4040 1.4560 0.4360 ;
    LAYER V0 ;
      RECT 1.4240 0.5300 1.4560 0.5620 ;
    LAYER V0 ;
      RECT 1.4240 0.6560 1.4560 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V0 ;
      RECT 1.4240 1.5800 1.4560 1.6120 ;
    LAYER V0 ;
      RECT 1.4240 1.7060 1.4560 1.7380 ;
    LAYER V0 ;
      RECT 1.4240 1.8320 1.4560 1.8640 ;
    LAYER V0 ;
      RECT 1.4240 2.0840 1.4560 2.1160 ;
    LAYER V0 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V0 ;
      RECT 1.4240 2.6720 1.4560 2.7040 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.5800 1.6160 1.6120 ;
    LAYER V0 ;
      RECT 1.5840 1.7060 1.6160 1.7380 ;
    LAYER V0 ;
      RECT 1.5840 1.8320 1.6160 1.8640 ;
    LAYER V0 ;
      RECT 1.5840 2.0840 1.6160 2.1160 ;
    LAYER V0 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V0 ;
      RECT 1.5840 2.6720 1.6160 2.7040 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.7440 0.4040 1.7760 0.4360 ;
    LAYER V0 ;
      RECT 1.7440 0.5300 1.7760 0.5620 ;
    LAYER V0 ;
      RECT 1.7440 0.6560 1.7760 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.9080 1.7760 0.9400 ;
    LAYER V0 ;
      RECT 1.7440 1.5800 1.7760 1.6120 ;
    LAYER V0 ;
      RECT 1.7440 1.7060 1.7760 1.7380 ;
    LAYER V0 ;
      RECT 1.7440 1.8320 1.7760 1.8640 ;
    LAYER V0 ;
      RECT 1.7440 2.0840 1.7760 2.1160 ;
    LAYER V0 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V0 ;
      RECT 1.7440 2.6720 1.7760 2.7040 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.9040 0.4040 1.9360 0.4360 ;
    LAYER V0 ;
      RECT 1.9040 0.5300 1.9360 0.5620 ;
    LAYER V0 ;
      RECT 1.9040 0.6560 1.9360 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.9080 1.9360 0.9400 ;
    LAYER V0 ;
      RECT 1.9040 1.5800 1.9360 1.6120 ;
    LAYER V0 ;
      RECT 1.9040 1.7060 1.9360 1.7380 ;
    LAYER V0 ;
      RECT 1.9040 1.8320 1.9360 1.8640 ;
    LAYER V0 ;
      RECT 1.9040 2.0840 1.9360 2.1160 ;
    LAYER V0 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V0 ;
      RECT 1.9040 2.6720 1.9360 2.7040 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 1.5800 2.0160 1.6120 ;
    LAYER V0 ;
      RECT 1.9840 1.5800 2.0160 1.6120 ;
    LAYER V0 ;
      RECT 1.9840 1.7060 2.0160 1.7380 ;
    LAYER V0 ;
      RECT 1.9840 1.7060 2.0160 1.7380 ;
    LAYER V0 ;
      RECT 1.9840 1.8320 2.0160 1.8640 ;
    LAYER V0 ;
      RECT 1.9840 1.8320 2.0160 1.8640 ;
    LAYER V0 ;
      RECT 2.0640 0.4040 2.0960 0.4360 ;
    LAYER V0 ;
      RECT 2.0640 0.5300 2.0960 0.5620 ;
    LAYER V0 ;
      RECT 2.0640 0.6560 2.0960 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V0 ;
      RECT 2.0640 1.5800 2.0960 1.6120 ;
    LAYER V0 ;
      RECT 2.0640 1.7060 2.0960 1.7380 ;
    LAYER V0 ;
      RECT 2.0640 1.8320 2.0960 1.8640 ;
    LAYER V0 ;
      RECT 2.0640 2.0840 2.0960 2.1160 ;
    LAYER V0 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V0 ;
      RECT 2.0640 2.6720 2.0960 2.7040 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.5800 2.2560 1.6120 ;
    LAYER V0 ;
      RECT 2.2240 1.7060 2.2560 1.7380 ;
    LAYER V0 ;
      RECT 2.2240 1.8320 2.2560 1.8640 ;
    LAYER V0 ;
      RECT 2.2240 2.0840 2.2560 2.1160 ;
    LAYER V0 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V0 ;
      RECT 2.2240 2.6720 2.2560 2.7040 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 1.5800 2.3360 1.6120 ;
    LAYER V0 ;
      RECT 2.3040 1.5800 2.3360 1.6120 ;
    LAYER V0 ;
      RECT 2.3040 1.7060 2.3360 1.7380 ;
    LAYER V0 ;
      RECT 2.3040 1.7060 2.3360 1.7380 ;
    LAYER V0 ;
      RECT 2.3040 1.8320 2.3360 1.8640 ;
    LAYER V0 ;
      RECT 2.3040 1.8320 2.3360 1.8640 ;
    LAYER V0 ;
      RECT 2.3840 0.4040 2.4160 0.4360 ;
    LAYER V0 ;
      RECT 2.3840 0.5300 2.4160 0.5620 ;
    LAYER V0 ;
      RECT 2.3840 0.6560 2.4160 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.9080 2.4160 0.9400 ;
    LAYER V0 ;
      RECT 2.3840 1.5800 2.4160 1.6120 ;
    LAYER V0 ;
      RECT 2.3840 1.7060 2.4160 1.7380 ;
    LAYER V0 ;
      RECT 2.3840 1.8320 2.4160 1.8640 ;
    LAYER V0 ;
      RECT 2.3840 2.0840 2.4160 2.1160 ;
    LAYER V0 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V0 ;
      RECT 2.3840 2.6720 2.4160 2.7040 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.5440 0.4040 2.5760 0.4360 ;
    LAYER V0 ;
      RECT 2.5440 0.5300 2.5760 0.5620 ;
    LAYER V0 ;
      RECT 2.5440 0.6560 2.5760 0.6880 ;
    LAYER V0 ;
      RECT 2.5440 0.9080 2.5760 0.9400 ;
    LAYER V0 ;
      RECT 2.5440 1.5800 2.5760 1.6120 ;
    LAYER V0 ;
      RECT 2.5440 1.7060 2.5760 1.7380 ;
    LAYER V0 ;
      RECT 2.5440 1.8320 2.5760 1.8640 ;
    LAYER V0 ;
      RECT 2.5440 2.0840 2.5760 2.1160 ;
    LAYER V0 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V0 ;
      RECT 2.5440 2.6720 2.5760 2.7040 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 1.5800 2.6560 1.6120 ;
    LAYER V0 ;
      RECT 2.6240 1.5800 2.6560 1.6120 ;
    LAYER V0 ;
      RECT 2.6240 1.7060 2.6560 1.7380 ;
    LAYER V0 ;
      RECT 2.6240 1.7060 2.6560 1.7380 ;
    LAYER V0 ;
      RECT 2.6240 1.8320 2.6560 1.8640 ;
    LAYER V0 ;
      RECT 2.6240 1.8320 2.6560 1.8640 ;
    LAYER V0 ;
      RECT 2.7040 0.4040 2.7360 0.4360 ;
    LAYER V0 ;
      RECT 2.7040 0.5300 2.7360 0.5620 ;
    LAYER V0 ;
      RECT 2.7040 0.6560 2.7360 0.6880 ;
    LAYER V0 ;
      RECT 2.7040 0.9080 2.7360 0.9400 ;
    LAYER V0 ;
      RECT 2.7040 1.5800 2.7360 1.6120 ;
    LAYER V0 ;
      RECT 2.7040 1.7060 2.7360 1.7380 ;
    LAYER V0 ;
      RECT 2.7040 1.8320 2.7360 1.8640 ;
    LAYER V0 ;
      RECT 2.7040 2.0840 2.7360 2.1160 ;
    LAYER V0 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V0 ;
      RECT 2.7040 2.6720 2.7360 2.7040 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.7840 1.5800 2.8160 1.6120 ;
    LAYER V0 ;
      RECT 2.7840 1.7060 2.8160 1.7380 ;
    LAYER V0 ;
      RECT 2.7840 1.8320 2.8160 1.8640 ;
  END
END DP_NMOS_B_nfin12_m16_n12_X8_Y2
MACRO CCP_PMOS_nfin12_m4_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_nfin12_m4_n12_X2_Y2 0 0 ;
  SIZE 1.1200 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 2.7240 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 2.1360 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.2160 0.5000 2.2200 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.5680 0.8160 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 0.6760 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9920 0.8360 1.0240 ;
    LAYER M2 ;
      RECT 0.4440 0.2360 0.6760 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 2.6720 0.8360 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.8360 2.1160 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 0.6760 1.3600 ;
    LAYER M2 ;
      RECT 0.4440 2.1680 0.6760 2.2000 ;
    LAYER M2 ;
      RECT 0.2840 1.4120 0.8360 1.4440 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.1680 0.6560 2.2000 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.1680 0.4960 2.2000 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9920 0.8160 1.0240 ;
    LAYER V1 ;
      RECT 0.7840 1.4120 0.8160 1.4440 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4120 0.3360 1.4440 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V2 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V2 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V2 ;
      RECT 0.4640 1.4120 0.4960 1.4440 ;
    LAYER V2 ;
      RECT 0.4640 2.1680 0.4960 2.2000 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
  END
END CCP_PMOS_nfin12_m4_n12_X2_Y2
MACRO Switch_NMOS_nfin12_m8_n12_X4_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin12_m8_n12_X4_Y2 0 0 ;
  SIZE 1.1200 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.8880 0.5000 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.2240 0.6560 1.9680 ;
    LAYER M1 ;
      RECT 0.6240 2.0640 0.6560 2.3040 ;
    LAYER M1 ;
      RECT 0.6240 2.5680 0.6560 2.8080 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.2240 0.8160 1.9680 ;
    LAYER M1 ;
      RECT 0.7840 2.0640 0.8160 2.3040 ;
    LAYER M1 ;
      RECT 0.7840 2.5680 0.8160 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.8360 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 2.6720 0.8360 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 0.8360 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.8360 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 1.2440 0.7360 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.3280 0.6560 1.3600 ;
    LAYER V1 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V1 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.3280 0.8160 1.3600 ;
    LAYER V1 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V1 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.5800 0.6560 1.6120 ;
    LAYER V0 ;
      RECT 0.6240 1.7060 0.6560 1.7380 ;
    LAYER V0 ;
      RECT 0.6240 1.8320 0.6560 1.8640 ;
    LAYER V0 ;
      RECT 0.6240 2.0840 0.6560 2.1160 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.5800 0.8160 1.6120 ;
    LAYER V0 ;
      RECT 0.7840 1.7060 0.8160 1.7380 ;
    LAYER V0 ;
      RECT 0.7840 1.8320 0.8160 1.8640 ;
    LAYER V0 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.7840 2.6720 0.8160 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
  END
END Switch_NMOS_nfin12_m8_n12_X4_Y2
MACRO CCP_S_NMOS_B_nfin12_m8_n12_X8_Y1
  ORIGIN 0 0 ;
  FOREIGN CCP_S_NMOS_B_nfin12_m8_n12_X8_Y1 0 0 ;
  SIZE 10.2400 BY 1.8480 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 10.0360 0.1000 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.1520 9.3960 0.1840 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5.1000 0.2160 5.1400 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5.1800 0.3000 5.2200 1.0440 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 9.9560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.3920 1.6160 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.3920 2.2560 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7920 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.1280 ;
    LAYER M1 ;
      RECT 2.8640 1.3920 2.8960 1.6320 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7920 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7920 ;
    LAYER M1 ;
      RECT 3.5040 0.8880 3.5360 1.1280 ;
    LAYER M1 ;
      RECT 3.5040 1.3920 3.5360 1.6320 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7920 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7920 ;
    LAYER M1 ;
      RECT 4.1440 0.0480 4.1760 0.7920 ;
    LAYER M1 ;
      RECT 4.1440 0.8880 4.1760 1.1280 ;
    LAYER M1 ;
      RECT 4.1440 1.3920 4.1760 1.6320 ;
    LAYER M1 ;
      RECT 4.0640 0.0480 4.0960 0.7920 ;
    LAYER M1 ;
      RECT 4.2240 0.0480 4.2560 0.7920 ;
    LAYER M1 ;
      RECT 4.7840 0.0480 4.8160 0.7920 ;
    LAYER M1 ;
      RECT 4.7840 0.8880 4.8160 1.1280 ;
    LAYER M1 ;
      RECT 4.7840 1.3920 4.8160 1.6320 ;
    LAYER M1 ;
      RECT 4.7040 0.0480 4.7360 0.7920 ;
    LAYER M1 ;
      RECT 4.8640 0.0480 4.8960 0.7920 ;
    LAYER M1 ;
      RECT 5.4240 0.0480 5.4560 0.7920 ;
    LAYER M1 ;
      RECT 5.4240 0.8880 5.4560 1.1280 ;
    LAYER M1 ;
      RECT 5.4240 1.3920 5.4560 1.6320 ;
    LAYER M1 ;
      RECT 5.3440 0.0480 5.3760 0.7920 ;
    LAYER M1 ;
      RECT 5.5040 0.0480 5.5360 0.7920 ;
    LAYER M1 ;
      RECT 6.0640 0.0480 6.0960 0.7920 ;
    LAYER M1 ;
      RECT 6.0640 0.8880 6.0960 1.1280 ;
    LAYER M1 ;
      RECT 6.0640 1.3920 6.0960 1.6320 ;
    LAYER M1 ;
      RECT 5.9840 0.0480 6.0160 0.7920 ;
    LAYER M1 ;
      RECT 6.1440 0.0480 6.1760 0.7920 ;
    LAYER M1 ;
      RECT 6.7040 0.0480 6.7360 0.7920 ;
    LAYER M1 ;
      RECT 6.7040 0.8880 6.7360 1.1280 ;
    LAYER M1 ;
      RECT 6.7040 1.3920 6.7360 1.6320 ;
    LAYER M1 ;
      RECT 6.6240 0.0480 6.6560 0.7920 ;
    LAYER M1 ;
      RECT 6.7840 0.0480 6.8160 0.7920 ;
    LAYER M1 ;
      RECT 7.3440 0.0480 7.3760 0.7920 ;
    LAYER M1 ;
      RECT 7.3440 0.8880 7.3760 1.1280 ;
    LAYER M1 ;
      RECT 7.3440 1.3920 7.3760 1.6320 ;
    LAYER M1 ;
      RECT 7.2640 0.0480 7.2960 0.7920 ;
    LAYER M1 ;
      RECT 7.4240 0.0480 7.4560 0.7920 ;
    LAYER M1 ;
      RECT 7.9840 0.0480 8.0160 0.7920 ;
    LAYER M1 ;
      RECT 7.9840 0.8880 8.0160 1.1280 ;
    LAYER M1 ;
      RECT 7.9840 1.3920 8.0160 1.6320 ;
    LAYER M1 ;
      RECT 7.9040 0.0480 7.9360 0.7920 ;
    LAYER M1 ;
      RECT 8.0640 0.0480 8.0960 0.7920 ;
    LAYER M1 ;
      RECT 8.6240 0.0480 8.6560 0.7920 ;
    LAYER M1 ;
      RECT 8.6240 0.8880 8.6560 1.1280 ;
    LAYER M1 ;
      RECT 8.6240 1.3920 8.6560 1.6320 ;
    LAYER M1 ;
      RECT 8.5440 0.0480 8.5760 0.7920 ;
    LAYER M1 ;
      RECT 8.7040 0.0480 8.7360 0.7920 ;
    LAYER M1 ;
      RECT 9.2640 0.0480 9.2960 0.7920 ;
    LAYER M1 ;
      RECT 9.2640 0.8880 9.2960 1.1280 ;
    LAYER M1 ;
      RECT 9.2640 1.3920 9.2960 1.6320 ;
    LAYER M1 ;
      RECT 9.1840 0.0480 9.2160 0.7920 ;
    LAYER M1 ;
      RECT 9.3440 0.0480 9.3760 0.7920 ;
    LAYER M1 ;
      RECT 9.9040 0.0480 9.9360 0.7920 ;
    LAYER M1 ;
      RECT 9.9040 0.8880 9.9360 1.1280 ;
    LAYER M1 ;
      RECT 9.9040 1.3920 9.9360 1.6320 ;
    LAYER M1 ;
      RECT 9.8240 0.0480 9.8560 0.7920 ;
    LAYER M1 ;
      RECT 9.9840 0.0480 10.0160 0.7920 ;
    LAYER M2 ;
      RECT 0.9240 0.9080 9.3160 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 9.9560 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.9920 9.9560 1.0240 ;
    LAYER M2 ;
      RECT 0.9240 0.3200 9.3160 0.3520 ;
    LAYER V1 ;
      RECT 5.3440 0.0680 5.3760 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 7.9040 0.0680 7.9360 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 8.0640 0.0680 8.0960 0.1000 ;
    LAYER V1 ;
      RECT 5.5040 0.0680 5.5360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 9.8240 0.0680 9.8560 0.1000 ;
    LAYER V1 ;
      RECT 2.9440 0.0680 2.9760 0.1000 ;
    LAYER V1 ;
      RECT 4.7040 0.0680 4.7360 0.1000 ;
    LAYER V1 ;
      RECT 4.8640 0.0680 4.8960 0.1000 ;
    LAYER V1 ;
      RECT 7.4240 0.0680 7.4560 0.1000 ;
    LAYER V1 ;
      RECT 9.9840 0.0680 10.0160 0.1000 ;
    LAYER V1 ;
      RECT 7.2640 0.0680 7.2960 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.1520 0.8960 0.1840 ;
    LAYER V1 ;
      RECT 8.5440 0.1520 8.5760 0.1840 ;
    LAYER V1 ;
      RECT 3.5840 0.1520 3.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 8.7040 0.1520 8.7360 0.1840 ;
    LAYER V1 ;
      RECT 3.4240 0.1520 3.4560 0.1840 ;
    LAYER V1 ;
      RECT 6.1440 0.1520 6.1760 0.1840 ;
    LAYER V1 ;
      RECT 5.9840 0.1520 6.0160 0.1840 ;
    LAYER V1 ;
      RECT 9.1840 0.1520 9.2160 0.1840 ;
    LAYER V1 ;
      RECT 1.5040 0.1520 1.5360 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 6.6240 0.1520 6.6560 0.1840 ;
    LAYER V1 ;
      RECT 6.7840 0.1520 6.8160 0.1840 ;
    LAYER V1 ;
      RECT 4.2240 0.1520 4.2560 0.1840 ;
    LAYER V1 ;
      RECT 9.3440 0.1520 9.3760 0.1840 ;
    LAYER V1 ;
      RECT 4.0640 0.1520 4.0960 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 6.0640 0.3200 6.0960 0.3520 ;
    LAYER V1 ;
      RECT 6.0640 0.9080 6.0960 0.9400 ;
    LAYER V1 ;
      RECT 6.0640 1.4960 6.0960 1.5280 ;
    LAYER V1 ;
      RECT 8.6240 0.3200 8.6560 0.3520 ;
    LAYER V1 ;
      RECT 8.6240 0.9080 8.6560 0.9400 ;
    LAYER V1 ;
      RECT 8.6240 1.4960 8.6560 1.5280 ;
    LAYER V1 ;
      RECT 3.5040 0.3200 3.5360 0.3520 ;
    LAYER V1 ;
      RECT 3.5040 0.9080 3.5360 0.9400 ;
    LAYER V1 ;
      RECT 3.5040 1.4960 3.5360 1.5280 ;
    LAYER V1 ;
      RECT 1.5840 0.3200 1.6160 0.3520 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V1 ;
      RECT 6.7040 0.3200 6.7360 0.3520 ;
    LAYER V1 ;
      RECT 6.7040 0.9080 6.7360 0.9400 ;
    LAYER V1 ;
      RECT 6.7040 1.4960 6.7360 1.5280 ;
    LAYER V1 ;
      RECT 4.1440 0.3200 4.1760 0.3520 ;
    LAYER V1 ;
      RECT 4.1440 0.9080 4.1760 0.9400 ;
    LAYER V1 ;
      RECT 4.1440 1.4960 4.1760 1.5280 ;
    LAYER V1 ;
      RECT 9.2640 0.3200 9.2960 0.3520 ;
    LAYER V1 ;
      RECT 9.2640 0.9080 9.2960 0.9400 ;
    LAYER V1 ;
      RECT 9.2640 1.4960 9.2960 1.5280 ;
    LAYER V1 ;
      RECT 7.9840 0.2360 8.0160 0.2680 ;
    LAYER V1 ;
      RECT 7.9840 0.9920 8.0160 1.0240 ;
    LAYER V1 ;
      RECT 7.9840 1.4960 8.0160 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 5.4240 0.2360 5.4560 0.2680 ;
    LAYER V1 ;
      RECT 5.4240 0.9920 5.4560 1.0240 ;
    LAYER V1 ;
      RECT 5.4240 1.4960 5.4560 1.5280 ;
    LAYER V1 ;
      RECT 2.8640 0.2360 2.8960 0.2680 ;
    LAYER V1 ;
      RECT 2.8640 0.9920 2.8960 1.0240 ;
    LAYER V1 ;
      RECT 2.8640 1.4960 2.8960 1.5280 ;
    LAYER V1 ;
      RECT 2.2240 0.2360 2.2560 0.2680 ;
    LAYER V1 ;
      RECT 2.2240 0.9920 2.2560 1.0240 ;
    LAYER V1 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V1 ;
      RECT 4.7840 0.2360 4.8160 0.2680 ;
    LAYER V1 ;
      RECT 4.7840 0.9920 4.8160 1.0240 ;
    LAYER V1 ;
      RECT 4.7840 1.4960 4.8160 1.5280 ;
    LAYER V1 ;
      RECT 9.9040 0.2360 9.9360 0.2680 ;
    LAYER V1 ;
      RECT 9.9040 0.9920 9.9360 1.0240 ;
    LAYER V1 ;
      RECT 9.9040 1.4960 9.9360 1.5280 ;
    LAYER V1 ;
      RECT 7.3440 0.2360 7.3760 0.2680 ;
    LAYER V1 ;
      RECT 7.3440 0.9920 7.3760 1.0240 ;
    LAYER V1 ;
      RECT 7.3440 1.4960 7.3760 1.5280 ;
    LAYER V2 ;
      RECT 5.1040 0.2360 5.1360 0.2680 ;
    LAYER V2 ;
      RECT 5.1040 0.9080 5.1360 0.9400 ;
    LAYER V2 ;
      RECT 5.1840 0.3200 5.2160 0.3520 ;
    LAYER V2 ;
      RECT 5.1840 0.9920 5.2160 1.0240 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.8640 0.4040 2.8960 0.4360 ;
    LAYER V0 ;
      RECT 2.8640 0.5300 2.8960 0.5620 ;
    LAYER V0 ;
      RECT 2.8640 0.6560 2.8960 0.6880 ;
    LAYER V0 ;
      RECT 2.8640 0.9080 2.8960 0.9400 ;
    LAYER V0 ;
      RECT 2.8640 1.4960 2.8960 1.5280 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.9440 0.4040 2.9760 0.4360 ;
    LAYER V0 ;
      RECT 2.9440 0.5300 2.9760 0.5620 ;
    LAYER V0 ;
      RECT 2.9440 0.6560 2.9760 0.6880 ;
    LAYER V0 ;
      RECT 3.5040 0.4040 3.5360 0.4360 ;
    LAYER V0 ;
      RECT 3.5040 0.5300 3.5360 0.5620 ;
    LAYER V0 ;
      RECT 3.5040 0.6560 3.5360 0.6880 ;
    LAYER V0 ;
      RECT 3.5040 0.9080 3.5360 0.9400 ;
    LAYER V0 ;
      RECT 3.5040 1.4960 3.5360 1.5280 ;
    LAYER V0 ;
      RECT 3.4240 0.4040 3.4560 0.4360 ;
    LAYER V0 ;
      RECT 3.4240 0.5300 3.4560 0.5620 ;
    LAYER V0 ;
      RECT 3.4240 0.6560 3.4560 0.6880 ;
    LAYER V0 ;
      RECT 3.5840 0.4040 3.6160 0.4360 ;
    LAYER V0 ;
      RECT 3.5840 0.5300 3.6160 0.5620 ;
    LAYER V0 ;
      RECT 3.5840 0.6560 3.6160 0.6880 ;
    LAYER V0 ;
      RECT 4.1440 0.4040 4.1760 0.4360 ;
    LAYER V0 ;
      RECT 4.1440 0.5300 4.1760 0.5620 ;
    LAYER V0 ;
      RECT 4.1440 0.6560 4.1760 0.6880 ;
    LAYER V0 ;
      RECT 4.1440 0.9080 4.1760 0.9400 ;
    LAYER V0 ;
      RECT 4.1440 1.4960 4.1760 1.5280 ;
    LAYER V0 ;
      RECT 4.0640 0.4040 4.0960 0.4360 ;
    LAYER V0 ;
      RECT 4.0640 0.5300 4.0960 0.5620 ;
    LAYER V0 ;
      RECT 4.0640 0.6560 4.0960 0.6880 ;
    LAYER V0 ;
      RECT 4.2240 0.4040 4.2560 0.4360 ;
    LAYER V0 ;
      RECT 4.2240 0.5300 4.2560 0.5620 ;
    LAYER V0 ;
      RECT 4.2240 0.6560 4.2560 0.6880 ;
    LAYER V0 ;
      RECT 4.7840 0.4040 4.8160 0.4360 ;
    LAYER V0 ;
      RECT 4.7840 0.5300 4.8160 0.5620 ;
    LAYER V0 ;
      RECT 4.7840 0.6560 4.8160 0.6880 ;
    LAYER V0 ;
      RECT 4.7840 0.9080 4.8160 0.9400 ;
    LAYER V0 ;
      RECT 4.7840 1.4960 4.8160 1.5280 ;
    LAYER V0 ;
      RECT 4.7040 0.4040 4.7360 0.4360 ;
    LAYER V0 ;
      RECT 4.7040 0.5300 4.7360 0.5620 ;
    LAYER V0 ;
      RECT 4.7040 0.6560 4.7360 0.6880 ;
    LAYER V0 ;
      RECT 4.8640 0.4040 4.8960 0.4360 ;
    LAYER V0 ;
      RECT 4.8640 0.5300 4.8960 0.5620 ;
    LAYER V0 ;
      RECT 4.8640 0.6560 4.8960 0.6880 ;
    LAYER V0 ;
      RECT 5.4240 0.4040 5.4560 0.4360 ;
    LAYER V0 ;
      RECT 5.4240 0.5300 5.4560 0.5620 ;
    LAYER V0 ;
      RECT 5.4240 0.6560 5.4560 0.6880 ;
    LAYER V0 ;
      RECT 5.4240 0.9080 5.4560 0.9400 ;
    LAYER V0 ;
      RECT 5.4240 1.4960 5.4560 1.5280 ;
    LAYER V0 ;
      RECT 5.3440 0.4040 5.3760 0.4360 ;
    LAYER V0 ;
      RECT 5.3440 0.5300 5.3760 0.5620 ;
    LAYER V0 ;
      RECT 5.3440 0.6560 5.3760 0.6880 ;
    LAYER V0 ;
      RECT 5.5040 0.4040 5.5360 0.4360 ;
    LAYER V0 ;
      RECT 5.5040 0.5300 5.5360 0.5620 ;
    LAYER V0 ;
      RECT 5.5040 0.6560 5.5360 0.6880 ;
    LAYER V0 ;
      RECT 6.0640 0.4040 6.0960 0.4360 ;
    LAYER V0 ;
      RECT 6.0640 0.5300 6.0960 0.5620 ;
    LAYER V0 ;
      RECT 6.0640 0.6560 6.0960 0.6880 ;
    LAYER V0 ;
      RECT 6.0640 0.9080 6.0960 0.9400 ;
    LAYER V0 ;
      RECT 6.0640 1.4960 6.0960 1.5280 ;
    LAYER V0 ;
      RECT 5.9840 0.4040 6.0160 0.4360 ;
    LAYER V0 ;
      RECT 5.9840 0.5300 6.0160 0.5620 ;
    LAYER V0 ;
      RECT 5.9840 0.6560 6.0160 0.6880 ;
    LAYER V0 ;
      RECT 6.1440 0.4040 6.1760 0.4360 ;
    LAYER V0 ;
      RECT 6.1440 0.5300 6.1760 0.5620 ;
    LAYER V0 ;
      RECT 6.1440 0.6560 6.1760 0.6880 ;
    LAYER V0 ;
      RECT 6.7040 0.4040 6.7360 0.4360 ;
    LAYER V0 ;
      RECT 6.7040 0.5300 6.7360 0.5620 ;
    LAYER V0 ;
      RECT 6.7040 0.6560 6.7360 0.6880 ;
    LAYER V0 ;
      RECT 6.7040 0.9080 6.7360 0.9400 ;
    LAYER V0 ;
      RECT 6.7040 1.4960 6.7360 1.5280 ;
    LAYER V0 ;
      RECT 6.6240 0.4040 6.6560 0.4360 ;
    LAYER V0 ;
      RECT 6.6240 0.5300 6.6560 0.5620 ;
    LAYER V0 ;
      RECT 6.6240 0.6560 6.6560 0.6880 ;
    LAYER V0 ;
      RECT 6.7840 0.4040 6.8160 0.4360 ;
    LAYER V0 ;
      RECT 6.7840 0.5300 6.8160 0.5620 ;
    LAYER V0 ;
      RECT 6.7840 0.6560 6.8160 0.6880 ;
    LAYER V0 ;
      RECT 7.3440 0.4040 7.3760 0.4360 ;
    LAYER V0 ;
      RECT 7.3440 0.5300 7.3760 0.5620 ;
    LAYER V0 ;
      RECT 7.3440 0.6560 7.3760 0.6880 ;
    LAYER V0 ;
      RECT 7.3440 0.9080 7.3760 0.9400 ;
    LAYER V0 ;
      RECT 7.3440 1.4960 7.3760 1.5280 ;
    LAYER V0 ;
      RECT 7.2640 0.4040 7.2960 0.4360 ;
    LAYER V0 ;
      RECT 7.2640 0.5300 7.2960 0.5620 ;
    LAYER V0 ;
      RECT 7.2640 0.6560 7.2960 0.6880 ;
    LAYER V0 ;
      RECT 7.4240 0.4040 7.4560 0.4360 ;
    LAYER V0 ;
      RECT 7.4240 0.5300 7.4560 0.5620 ;
    LAYER V0 ;
      RECT 7.4240 0.6560 7.4560 0.6880 ;
    LAYER V0 ;
      RECT 7.9840 0.4040 8.0160 0.4360 ;
    LAYER V0 ;
      RECT 7.9840 0.5300 8.0160 0.5620 ;
    LAYER V0 ;
      RECT 7.9840 0.6560 8.0160 0.6880 ;
    LAYER V0 ;
      RECT 7.9840 0.9080 8.0160 0.9400 ;
    LAYER V0 ;
      RECT 7.9840 1.4960 8.0160 1.5280 ;
    LAYER V0 ;
      RECT 7.9040 0.4040 7.9360 0.4360 ;
    LAYER V0 ;
      RECT 7.9040 0.5300 7.9360 0.5620 ;
    LAYER V0 ;
      RECT 7.9040 0.6560 7.9360 0.6880 ;
    LAYER V0 ;
      RECT 8.0640 0.4040 8.0960 0.4360 ;
    LAYER V0 ;
      RECT 8.0640 0.5300 8.0960 0.5620 ;
    LAYER V0 ;
      RECT 8.0640 0.6560 8.0960 0.6880 ;
    LAYER V0 ;
      RECT 8.6240 0.4040 8.6560 0.4360 ;
    LAYER V0 ;
      RECT 8.6240 0.5300 8.6560 0.5620 ;
    LAYER V0 ;
      RECT 8.6240 0.6560 8.6560 0.6880 ;
    LAYER V0 ;
      RECT 8.6240 0.9080 8.6560 0.9400 ;
    LAYER V0 ;
      RECT 8.6240 1.4960 8.6560 1.5280 ;
    LAYER V0 ;
      RECT 8.5440 0.4040 8.5760 0.4360 ;
    LAYER V0 ;
      RECT 8.5440 0.5300 8.5760 0.5620 ;
    LAYER V0 ;
      RECT 8.5440 0.6560 8.5760 0.6880 ;
    LAYER V0 ;
      RECT 8.7040 0.4040 8.7360 0.4360 ;
    LAYER V0 ;
      RECT 8.7040 0.5300 8.7360 0.5620 ;
    LAYER V0 ;
      RECT 8.7040 0.6560 8.7360 0.6880 ;
    LAYER V0 ;
      RECT 9.2640 0.4040 9.2960 0.4360 ;
    LAYER V0 ;
      RECT 9.2640 0.5300 9.2960 0.5620 ;
    LAYER V0 ;
      RECT 9.2640 0.6560 9.2960 0.6880 ;
    LAYER V0 ;
      RECT 9.2640 0.9080 9.2960 0.9400 ;
    LAYER V0 ;
      RECT 9.2640 1.4960 9.2960 1.5280 ;
    LAYER V0 ;
      RECT 9.1840 0.4040 9.2160 0.4360 ;
    LAYER V0 ;
      RECT 9.1840 0.5300 9.2160 0.5620 ;
    LAYER V0 ;
      RECT 9.1840 0.6560 9.2160 0.6880 ;
    LAYER V0 ;
      RECT 9.3440 0.4040 9.3760 0.4360 ;
    LAYER V0 ;
      RECT 9.3440 0.5300 9.3760 0.5620 ;
    LAYER V0 ;
      RECT 9.3440 0.6560 9.3760 0.6880 ;
    LAYER V0 ;
      RECT 9.9040 0.4040 9.9360 0.4360 ;
    LAYER V0 ;
      RECT 9.9040 0.5300 9.9360 0.5620 ;
    LAYER V0 ;
      RECT 9.9040 0.6560 9.9360 0.6880 ;
    LAYER V0 ;
      RECT 9.9040 0.9080 9.9360 0.9400 ;
    LAYER V0 ;
      RECT 9.9040 1.4960 9.9360 1.5280 ;
    LAYER V0 ;
      RECT 9.8240 0.4040 9.8560 0.4360 ;
    LAYER V0 ;
      RECT 9.8240 0.5300 9.8560 0.5620 ;
    LAYER V0 ;
      RECT 9.8240 0.6560 9.8560 0.6880 ;
    LAYER V0 ;
      RECT 9.9840 0.4040 10.0160 0.4360 ;
    LAYER V0 ;
      RECT 9.9840 0.5300 10.0160 0.5620 ;
    LAYER V0 ;
      RECT 9.9840 0.6560 10.0160 0.6880 ;
  END
END CCP_S_NMOS_B_nfin12_m8_n12_X8_Y1
