VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RES_w1u_l14u
  UNITS 
    DATABASE MICRONS UNITS 1 ;
  END UNITS 

  ORIGIN 0 0 ;
  FOREIGN RES_w1u_l14u 0 0 ;
  SIZE 14.3 BY 1.2 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1 0.15 0.42 1.15 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.14 0.15 14.46 1.15 ;
    END
  END MINUS
END RES_w1u_l14u

