MACRO Switch_NMOS_n12_X4_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X4_Y2 0 0 ;
  SIZE 2.3400 BY 4.0320 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9980 0.3420 1.0300 1.7700 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.0760 0.4380 1.1080 1.8660 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1540 1.3020 1.1860 2.7300 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 3.3440 1.6740 3.3760 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.1260 0.9520 3.4980 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 0.3420 1.1080 1.1940 ;
    LAYER M1 ;
      RECT 1.0760 1.3020 1.1080 1.5780 ;
    LAYER M1 ;
      RECT 1.0760 1.6860 1.1080 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 2.6460 1.1080 2.9220 ;
    LAYER M1 ;
      RECT 1.1540 0.3420 1.1860 1.1940 ;
    LAYER M1 ;
      RECT 1.1540 1.6860 1.1860 2.5380 ;
    LAYER M1 ;
      RECT 1.2320 0.3420 1.2640 1.1940 ;
    LAYER M1 ;
      RECT 1.2320 1.3020 1.2640 1.5780 ;
    LAYER M1 ;
      RECT 1.2320 1.6860 1.2640 2.5380 ;
    LAYER M1 ;
      RECT 1.2320 2.6460 1.2640 2.9220 ;
    LAYER M1 ;
      RECT 1.3100 0.3420 1.3420 1.1940 ;
    LAYER M1 ;
      RECT 1.3100 1.6860 1.3420 2.5380 ;
    LAYER M1 ;
      RECT 1.3880 0.3420 1.4200 1.1940 ;
    LAYER M1 ;
      RECT 1.3880 1.3020 1.4200 1.5780 ;
    LAYER M1 ;
      RECT 1.3880 1.6860 1.4200 2.5380 ;
    LAYER M1 ;
      RECT 1.3880 2.6460 1.4200 2.9220 ;
    LAYER M1 ;
      RECT 1.3880 3.1260 1.4200 3.4980 ;
    LAYER M1 ;
      RECT 1.4660 0.3420 1.4980 1.1940 ;
    LAYER M1 ;
      RECT 1.4660 1.6860 1.4980 2.5380 ;
    LAYER M2 ;
      RECT 0.7380 0.3680 1.5240 0.4000 ;
    LAYER M2 ;
      RECT 0.8160 0.4640 1.4460 0.4960 ;
    LAYER M2 ;
      RECT 0.8160 1.3280 1.4460 1.3600 ;
    LAYER M2 ;
      RECT 0.7380 1.7120 1.5240 1.7440 ;
    LAYER M2 ;
      RECT 0.8160 1.8080 1.4460 1.8400 ;
    LAYER M2 ;
      RECT 0.8160 2.6720 1.4460 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 1.8080 0.9520 1.8400 ;
    LAYER V1 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V1 ;
      RECT 1.3880 0.4640 1.4200 0.4960 ;
    LAYER V1 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V1 ;
      RECT 1.3880 1.8080 1.4200 1.8400 ;
    LAYER V1 ;
      RECT 1.3880 2.6720 1.4200 2.7040 ;
    LAYER V1 ;
      RECT 1.3880 3.3440 1.4200 3.3760 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.8420 1.7120 0.8740 1.7440 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V1 ;
      RECT 1.1540 0.3680 1.1860 0.4000 ;
    LAYER V1 ;
      RECT 1.1540 1.7120 1.1860 1.7440 ;
    LAYER V1 ;
      RECT 1.3100 0.3680 1.3420 0.4000 ;
    LAYER V1 ;
      RECT 1.3100 1.7120 1.3420 1.7440 ;
    LAYER V1 ;
      RECT 1.4660 0.3680 1.4980 0.4000 ;
    LAYER V1 ;
      RECT 1.4660 1.7120 1.4980 1.7440 ;
    LAYER V1 ;
      RECT 1.2320 0.4640 1.2640 0.4960 ;
    LAYER V1 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V1 ;
      RECT 1.2320 1.8080 1.2640 1.8400 ;
    LAYER V1 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V1 ;
      RECT 1.0760 0.4640 1.1080 0.4960 ;
    LAYER V1 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V1 ;
      RECT 1.0760 1.8080 1.1080 1.8400 ;
    LAYER V1 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V2 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V2 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V2 ;
      RECT 1.0760 0.4640 1.1080 0.4960 ;
    LAYER V2 ;
      RECT 1.0760 1.8080 1.1080 1.8400 ;
    LAYER V2 ;
      RECT 1.1540 1.3280 1.1860 1.3600 ;
    LAYER V2 ;
      RECT 1.1540 2.6720 1.1860 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 0.7520 1.1080 0.7840 ;
    LAYER V0 ;
      RECT 1.0760 1.0400 1.1080 1.0720 ;
    LAYER V0 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V0 ;
      RECT 1.0760 2.0960 1.1080 2.1280 ;
    LAYER V0 ;
      RECT 1.0760 2.3840 1.1080 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.2320 0.7520 1.2640 0.7840 ;
    LAYER V0 ;
      RECT 1.2320 0.8960 1.2640 0.9280 ;
    LAYER V0 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V0 ;
      RECT 1.2320 2.0960 1.2640 2.1280 ;
    LAYER V0 ;
      RECT 1.2320 2.2400 1.2640 2.2720 ;
    LAYER V0 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3880 0.8960 1.4200 0.9280 ;
    LAYER V0 ;
      RECT 1.3880 1.0400 1.4200 1.0720 ;
    LAYER V0 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V0 ;
      RECT 1.3880 2.2400 1.4200 2.2720 ;
    LAYER V0 ;
      RECT 1.3880 2.3840 1.4200 2.4160 ;
    LAYER V0 ;
      RECT 1.3880 2.6720 1.4200 2.7040 ;
    LAYER V0 ;
      RECT 1.3880 3.3440 1.4200 3.3760 ;
    LAYER V0 ;
      RECT 1.3880 3.3440 1.4200 3.3760 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
  END
END Switch_NMOS_n12_X4_Y2
MACRO CCP_PMOS_S_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_S_n12_X2_Y2 0 0 ;
  SIZE 3.7440 BY 4.0320 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9340 0.3420 1.9660 1.7700 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.0120 0.4380 2.0440 2.7300 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.0900 0.5340 2.1220 2.8260 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 3.3440 3.0780 3.3760 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.1260 0.9520 3.4980 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 1.5440 0.3420 1.5760 1.1940 ;
    LAYER M1 ;
      RECT 1.5440 1.3020 1.5760 1.5780 ;
    LAYER M1 ;
      RECT 1.5440 1.6860 1.5760 2.5380 ;
    LAYER M1 ;
      RECT 1.5440 2.6460 1.5760 2.9220 ;
    LAYER M1 ;
      RECT 1.5440 3.1260 1.5760 3.4980 ;
    LAYER M1 ;
      RECT 1.4660 0.3420 1.4980 1.1940 ;
    LAYER M1 ;
      RECT 1.4660 1.6860 1.4980 2.5380 ;
    LAYER M1 ;
      RECT 1.6220 0.3420 1.6540 1.1940 ;
    LAYER M1 ;
      RECT 1.6220 1.6860 1.6540 2.5380 ;
    LAYER M1 ;
      RECT 2.1680 0.3420 2.2000 1.1940 ;
    LAYER M1 ;
      RECT 2.1680 1.3020 2.2000 1.5780 ;
    LAYER M1 ;
      RECT 2.1680 1.6860 2.2000 2.5380 ;
    LAYER M1 ;
      RECT 2.1680 2.6460 2.2000 2.9220 ;
    LAYER M1 ;
      RECT 2.1680 3.1260 2.2000 3.4980 ;
    LAYER M1 ;
      RECT 2.0900 0.3420 2.1220 1.1940 ;
    LAYER M1 ;
      RECT 2.0900 1.6860 2.1220 2.5380 ;
    LAYER M1 ;
      RECT 2.2460 0.3420 2.2780 1.1940 ;
    LAYER M1 ;
      RECT 2.2460 1.6860 2.2780 2.5380 ;
    LAYER M1 ;
      RECT 2.7920 0.3420 2.8240 1.1940 ;
    LAYER M1 ;
      RECT 2.7920 1.3020 2.8240 1.5780 ;
    LAYER M1 ;
      RECT 2.7920 1.6860 2.8240 2.5380 ;
    LAYER M1 ;
      RECT 2.7920 2.6460 2.8240 2.9220 ;
    LAYER M1 ;
      RECT 2.7920 3.1260 2.8240 3.4980 ;
    LAYER M1 ;
      RECT 2.7140 0.3420 2.7460 1.1940 ;
    LAYER M1 ;
      RECT 2.7140 1.6860 2.7460 2.5380 ;
    LAYER M1 ;
      RECT 2.8700 0.3420 2.9020 1.1940 ;
    LAYER M1 ;
      RECT 2.8700 1.6860 2.9020 2.5380 ;
    LAYER M2 ;
      RECT 0.7380 0.3680 2.9280 0.4000 ;
    LAYER M2 ;
      RECT 1.4400 1.3280 2.2260 1.3600 ;
    LAYER M2 ;
      RECT 0.8160 0.4640 2.8500 0.4960 ;
    LAYER M2 ;
      RECT 1.4400 0.5600 2.2260 0.5920 ;
    LAYER M2 ;
      RECT 0.8160 1.4240 2.8500 1.4560 ;
    LAYER M2 ;
      RECT 0.7380 1.7120 2.9280 1.7440 ;
    LAYER M2 ;
      RECT 1.4400 1.8080 2.2260 1.8400 ;
    LAYER M2 ;
      RECT 0.8160 2.6720 2.8500 2.7040 ;
    LAYER M2 ;
      RECT 1.4400 2.7680 2.2260 2.8000 ;
    LAYER M2 ;
      RECT 0.8160 1.9040 2.8500 1.9360 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.4240 0.9520 1.4560 ;
    LAYER V1 ;
      RECT 0.9200 1.9040 0.9520 1.9360 ;
    LAYER V1 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V1 ;
      RECT 1.5440 0.5600 1.5760 0.5920 ;
    LAYER V1 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V1 ;
      RECT 1.5440 1.8080 1.5760 1.8400 ;
    LAYER V1 ;
      RECT 1.5440 2.7680 1.5760 2.8000 ;
    LAYER V1 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V1 ;
      RECT 2.1680 0.5600 2.2000 0.5920 ;
    LAYER V1 ;
      RECT 2.1680 1.3280 2.2000 1.3600 ;
    LAYER V1 ;
      RECT 2.1680 1.8080 2.2000 1.8400 ;
    LAYER V1 ;
      RECT 2.1680 2.7680 2.2000 2.8000 ;
    LAYER V1 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V1 ;
      RECT 2.7920 0.4640 2.8240 0.4960 ;
    LAYER V1 ;
      RECT 2.7920 1.4240 2.8240 1.4560 ;
    LAYER V1 ;
      RECT 2.7920 1.9040 2.8240 1.9360 ;
    LAYER V1 ;
      RECT 2.7920 2.6720 2.8240 2.7040 ;
    LAYER V1 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.8420 1.7120 0.8740 1.7440 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V1 ;
      RECT 1.4660 0.3680 1.4980 0.4000 ;
    LAYER V1 ;
      RECT 1.4660 1.7120 1.4980 1.7440 ;
    LAYER V1 ;
      RECT 1.6220 0.3680 1.6540 0.4000 ;
    LAYER V1 ;
      RECT 1.6220 1.7120 1.6540 1.7440 ;
    LAYER V1 ;
      RECT 2.0900 0.3680 2.1220 0.4000 ;
    LAYER V1 ;
      RECT 2.0900 1.7120 2.1220 1.7440 ;
    LAYER V1 ;
      RECT 2.2460 0.3680 2.2780 0.4000 ;
    LAYER V1 ;
      RECT 2.2460 1.7120 2.2780 1.7440 ;
    LAYER V1 ;
      RECT 2.7140 0.3680 2.7460 0.4000 ;
    LAYER V1 ;
      RECT 2.7140 1.7120 2.7460 1.7440 ;
    LAYER V1 ;
      RECT 2.8700 0.3680 2.9020 0.4000 ;
    LAYER V1 ;
      RECT 2.8700 1.7120 2.9020 1.7440 ;
    LAYER V2 ;
      RECT 1.9340 0.3680 1.9660 0.4000 ;
    LAYER V2 ;
      RECT 1.9340 1.7120 1.9660 1.7440 ;
    LAYER V2 ;
      RECT 2.0120 0.4640 2.0440 0.4960 ;
    LAYER V2 ;
      RECT 2.0120 1.3280 2.0440 1.3600 ;
    LAYER V2 ;
      RECT 2.0120 1.8080 2.0440 1.8400 ;
    LAYER V2 ;
      RECT 2.0120 2.6720 2.0440 2.7040 ;
    LAYER V2 ;
      RECT 2.0900 0.5600 2.1220 0.5920 ;
    LAYER V2 ;
      RECT 2.0900 1.4240 2.1220 1.4560 ;
    LAYER V2 ;
      RECT 2.0900 1.9040 2.1220 1.9360 ;
    LAYER V2 ;
      RECT 2.0900 2.7680 2.1220 2.8000 ;
    LAYER V0 ;
      RECT 0.9200 0.7520 0.9520 0.7840 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.0960 0.9520 2.1280 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 1.5440 0.7520 1.5760 0.7840 ;
    LAYER V0 ;
      RECT 1.5440 0.8960 1.5760 0.9280 ;
    LAYER V0 ;
      RECT 1.5440 1.0400 1.5760 1.0720 ;
    LAYER V0 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V0 ;
      RECT 1.5440 2.0960 1.5760 2.1280 ;
    LAYER V0 ;
      RECT 1.5440 2.2400 1.5760 2.2720 ;
    LAYER V0 ;
      RECT 1.5440 2.3840 1.5760 2.4160 ;
    LAYER V0 ;
      RECT 1.5440 2.6720 1.5760 2.7040 ;
    LAYER V0 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V0 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
    LAYER V0 ;
      RECT 1.6220 0.7520 1.6540 0.7840 ;
    LAYER V0 ;
      RECT 1.6220 0.8960 1.6540 0.9280 ;
    LAYER V0 ;
      RECT 1.6220 1.0400 1.6540 1.0720 ;
    LAYER V0 ;
      RECT 1.6220 2.0960 1.6540 2.1280 ;
    LAYER V0 ;
      RECT 1.6220 2.2400 1.6540 2.2720 ;
    LAYER V0 ;
      RECT 1.6220 2.3840 1.6540 2.4160 ;
    LAYER V0 ;
      RECT 2.1680 0.7520 2.2000 0.7840 ;
    LAYER V0 ;
      RECT 2.1680 0.8960 2.2000 0.9280 ;
    LAYER V0 ;
      RECT 2.1680 1.0400 2.2000 1.0720 ;
    LAYER V0 ;
      RECT 2.1680 1.3280 2.2000 1.3600 ;
    LAYER V0 ;
      RECT 2.1680 2.0960 2.2000 2.1280 ;
    LAYER V0 ;
      RECT 2.1680 2.2400 2.2000 2.2720 ;
    LAYER V0 ;
      RECT 2.1680 2.3840 2.2000 2.4160 ;
    LAYER V0 ;
      RECT 2.1680 2.6720 2.2000 2.7040 ;
    LAYER V0 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V0 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V0 ;
      RECT 2.0900 0.7520 2.1220 0.7840 ;
    LAYER V0 ;
      RECT 2.0900 0.8960 2.1220 0.9280 ;
    LAYER V0 ;
      RECT 2.0900 1.0400 2.1220 1.0720 ;
    LAYER V0 ;
      RECT 2.0900 2.0960 2.1220 2.1280 ;
    LAYER V0 ;
      RECT 2.0900 2.2400 2.1220 2.2720 ;
    LAYER V0 ;
      RECT 2.0900 2.3840 2.1220 2.4160 ;
    LAYER V0 ;
      RECT 2.2460 0.7520 2.2780 0.7840 ;
    LAYER V0 ;
      RECT 2.2460 0.8960 2.2780 0.9280 ;
    LAYER V0 ;
      RECT 2.2460 1.0400 2.2780 1.0720 ;
    LAYER V0 ;
      RECT 2.2460 2.0960 2.2780 2.1280 ;
    LAYER V0 ;
      RECT 2.2460 2.2400 2.2780 2.2720 ;
    LAYER V0 ;
      RECT 2.2460 2.3840 2.2780 2.4160 ;
    LAYER V0 ;
      RECT 2.7920 0.7520 2.8240 0.7840 ;
    LAYER V0 ;
      RECT 2.7920 0.8960 2.8240 0.9280 ;
    LAYER V0 ;
      RECT 2.7920 1.0400 2.8240 1.0720 ;
    LAYER V0 ;
      RECT 2.7920 1.3280 2.8240 1.3600 ;
    LAYER V0 ;
      RECT 2.7920 2.0960 2.8240 2.1280 ;
    LAYER V0 ;
      RECT 2.7920 2.2400 2.8240 2.2720 ;
    LAYER V0 ;
      RECT 2.7920 2.3840 2.8240 2.4160 ;
    LAYER V0 ;
      RECT 2.7920 2.6720 2.8240 2.7040 ;
    LAYER V0 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V0 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V0 ;
      RECT 2.7140 0.7520 2.7460 0.7840 ;
    LAYER V0 ;
      RECT 2.7140 0.8960 2.7460 0.9280 ;
    LAYER V0 ;
      RECT 2.7140 1.0400 2.7460 1.0720 ;
    LAYER V0 ;
      RECT 2.7140 2.0960 2.7460 2.1280 ;
    LAYER V0 ;
      RECT 2.7140 2.2400 2.7460 2.2720 ;
    LAYER V0 ;
      RECT 2.7140 2.3840 2.7460 2.4160 ;
    LAYER V0 ;
      RECT 2.8700 0.7520 2.9020 0.7840 ;
    LAYER V0 ;
      RECT 2.8700 0.8960 2.9020 0.9280 ;
    LAYER V0 ;
      RECT 2.8700 1.0400 2.9020 1.0720 ;
    LAYER V0 ;
      RECT 2.8700 2.0960 2.9020 2.1280 ;
    LAYER V0 ;
      RECT 2.8700 2.2400 2.9020 2.2720 ;
    LAYER V0 ;
      RECT 2.8700 2.3840 2.9020 2.4160 ;
  END
END CCP_PMOS_S_n12_X2_Y2
MACRO Switch_PMOS_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y2 0 0 ;
  SIZE 2.0280 BY 4.0320 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8420 0.3420 0.8740 1.7700 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9200 0.4380 0.9520 1.8660 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9980 1.3020 1.0300 2.7300 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 3.3440 1.3620 3.3760 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.1260 0.9520 3.4980 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 0.3420 1.1080 1.1940 ;
    LAYER M1 ;
      RECT 1.0760 1.3020 1.1080 1.5780 ;
    LAYER M1 ;
      RECT 1.0760 1.6860 1.1080 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 2.6460 1.1080 2.9220 ;
    LAYER M1 ;
      RECT 1.1540 0.3420 1.1860 1.1940 ;
    LAYER M1 ;
      RECT 1.1540 1.6860 1.1860 2.5380 ;
    LAYER M2 ;
      RECT 0.7380 0.3680 1.2120 0.4000 ;
    LAYER M2 ;
      RECT 0.8160 0.4640 1.1340 0.4960 ;
    LAYER M2 ;
      RECT 0.8160 1.3280 1.1340 1.3600 ;
    LAYER M2 ;
      RECT 0.7380 1.7120 1.2120 1.7440 ;
    LAYER M2 ;
      RECT 0.8160 1.8080 1.1340 1.8400 ;
    LAYER M2 ;
      RECT 0.8160 2.6720 1.1340 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 1.8080 0.9520 1.8400 ;
    LAYER V1 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.8420 1.7120 0.8740 1.7440 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V1 ;
      RECT 1.1540 0.3680 1.1860 0.4000 ;
    LAYER V1 ;
      RECT 1.1540 1.7120 1.1860 1.7440 ;
    LAYER V1 ;
      RECT 1.0760 0.4640 1.1080 0.4960 ;
    LAYER V1 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V1 ;
      RECT 1.0760 1.8080 1.1080 1.8400 ;
    LAYER V1 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V2 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V2 ;
      RECT 0.8420 1.7120 0.8740 1.7440 ;
    LAYER V2 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V2 ;
      RECT 0.9200 1.8080 0.9520 1.8400 ;
    LAYER V2 ;
      RECT 0.9980 1.3280 1.0300 1.3600 ;
    LAYER V2 ;
      RECT 0.9980 2.6720 1.0300 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 0.7520 1.1080 0.7840 ;
    LAYER V0 ;
      RECT 1.0760 1.0400 1.1080 1.0720 ;
    LAYER V0 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V0 ;
      RECT 1.0760 2.0960 1.1080 2.1280 ;
    LAYER V0 ;
      RECT 1.0760 2.3840 1.1080 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
  END
END Switch_PMOS_n12_X2_Y2
MACRO DP_NMOS_n12_X4_Y4
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X4_Y4 0 0 ;
  SIZE 2.9640 BY 6.7200 ;
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2320 1.3020 1.2640 5.4180 ;
    END
  END GA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3100 0.3420 1.3420 4.4580 ;
    END
  END DA
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3880 0.4380 1.4200 4.5540 ;
    END
  END S
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4660 0.5340 1.4980 4.6500 ;
    END
  END DB
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5440 1.3980 1.5760 5.5140 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 6.0320 2.2980 6.0640 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.0300 0.9520 3.8820 ;
    LAYER M1 ;
      RECT 0.9200 3.9900 0.9520 4.2660 ;
    LAYER M1 ;
      RECT 0.9200 4.3740 0.9520 5.2260 ;
    LAYER M1 ;
      RECT 0.9200 5.3340 0.9520 5.6100 ;
    LAYER M1 ;
      RECT 0.9200 5.8140 0.9520 6.1860 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.8420 3.0300 0.8740 3.8820 ;
    LAYER M1 ;
      RECT 0.8420 4.3740 0.8740 5.2260 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 3.0300 1.0300 3.8820 ;
    LAYER M1 ;
      RECT 0.9980 4.3740 1.0300 5.2260 ;
    LAYER M1 ;
      RECT 1.0760 0.3420 1.1080 1.1940 ;
    LAYER M1 ;
      RECT 1.0760 1.3020 1.1080 1.5780 ;
    LAYER M1 ;
      RECT 1.0760 1.6860 1.1080 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 2.6460 1.1080 2.9220 ;
    LAYER M1 ;
      RECT 1.0760 3.0300 1.1080 3.8820 ;
    LAYER M1 ;
      RECT 1.0760 3.9900 1.1080 4.2660 ;
    LAYER M1 ;
      RECT 1.0760 4.3740 1.1080 5.2260 ;
    LAYER M1 ;
      RECT 1.0760 5.3340 1.1080 5.6100 ;
    LAYER M1 ;
      RECT 1.1540 0.3420 1.1860 1.1940 ;
    LAYER M1 ;
      RECT 1.1540 1.6860 1.1860 2.5380 ;
    LAYER M1 ;
      RECT 1.1540 3.0300 1.1860 3.8820 ;
    LAYER M1 ;
      RECT 1.1540 4.3740 1.1860 5.2260 ;
    LAYER M1 ;
      RECT 1.2320 0.3420 1.2640 1.1940 ;
    LAYER M1 ;
      RECT 1.2320 1.3020 1.2640 1.5780 ;
    LAYER M1 ;
      RECT 1.2320 1.6860 1.2640 2.5380 ;
    LAYER M1 ;
      RECT 1.2320 2.6460 1.2640 2.9220 ;
    LAYER M1 ;
      RECT 1.2320 3.0300 1.2640 3.8820 ;
    LAYER M1 ;
      RECT 1.2320 3.9900 1.2640 4.2660 ;
    LAYER M1 ;
      RECT 1.2320 4.3740 1.2640 5.2260 ;
    LAYER M1 ;
      RECT 1.2320 5.3340 1.2640 5.6100 ;
    LAYER M1 ;
      RECT 1.3100 0.3420 1.3420 1.1940 ;
    LAYER M1 ;
      RECT 1.3100 1.6860 1.3420 2.5380 ;
    LAYER M1 ;
      RECT 1.3100 3.0300 1.3420 3.8820 ;
    LAYER M1 ;
      RECT 1.3100 4.3740 1.3420 5.2260 ;
    LAYER M1 ;
      RECT 1.3880 0.3420 1.4200 1.1940 ;
    LAYER M1 ;
      RECT 1.3880 1.3020 1.4200 1.5780 ;
    LAYER M1 ;
      RECT 1.3880 1.6860 1.4200 2.5380 ;
    LAYER M1 ;
      RECT 1.3880 2.6460 1.4200 2.9220 ;
    LAYER M1 ;
      RECT 1.3880 3.0300 1.4200 3.8820 ;
    LAYER M1 ;
      RECT 1.3880 3.9900 1.4200 4.2660 ;
    LAYER M1 ;
      RECT 1.3880 4.3740 1.4200 5.2260 ;
    LAYER M1 ;
      RECT 1.3880 5.3340 1.4200 5.6100 ;
    LAYER M1 ;
      RECT 1.3880 5.8140 1.4200 6.1860 ;
    LAYER M1 ;
      RECT 1.4660 0.3420 1.4980 1.1940 ;
    LAYER M1 ;
      RECT 1.4660 1.6860 1.4980 2.5380 ;
    LAYER M1 ;
      RECT 1.4660 3.0300 1.4980 3.8820 ;
    LAYER M1 ;
      RECT 1.4660 4.3740 1.4980 5.2260 ;
    LAYER M1 ;
      RECT 1.5440 0.3420 1.5760 1.1940 ;
    LAYER M1 ;
      RECT 1.5440 1.3020 1.5760 1.5780 ;
    LAYER M1 ;
      RECT 1.5440 1.6860 1.5760 2.5380 ;
    LAYER M1 ;
      RECT 1.5440 2.6460 1.5760 2.9220 ;
    LAYER M1 ;
      RECT 1.5440 3.0300 1.5760 3.8820 ;
    LAYER M1 ;
      RECT 1.5440 3.9900 1.5760 4.2660 ;
    LAYER M1 ;
      RECT 1.5440 4.3740 1.5760 5.2260 ;
    LAYER M1 ;
      RECT 1.5440 5.3340 1.5760 5.6100 ;
    LAYER M1 ;
      RECT 1.6220 0.3420 1.6540 1.1940 ;
    LAYER M1 ;
      RECT 1.6220 1.6860 1.6540 2.5380 ;
    LAYER M1 ;
      RECT 1.6220 3.0300 1.6540 3.8820 ;
    LAYER M1 ;
      RECT 1.6220 4.3740 1.6540 5.2260 ;
    LAYER M1 ;
      RECT 1.7000 0.3420 1.7320 1.1940 ;
    LAYER M1 ;
      RECT 1.7000 1.3020 1.7320 1.5780 ;
    LAYER M1 ;
      RECT 1.7000 1.6860 1.7320 2.5380 ;
    LAYER M1 ;
      RECT 1.7000 2.6460 1.7320 2.9220 ;
    LAYER M1 ;
      RECT 1.7000 3.0300 1.7320 3.8820 ;
    LAYER M1 ;
      RECT 1.7000 3.9900 1.7320 4.2660 ;
    LAYER M1 ;
      RECT 1.7000 4.3740 1.7320 5.2260 ;
    LAYER M1 ;
      RECT 1.7000 5.3340 1.7320 5.6100 ;
    LAYER M1 ;
      RECT 1.7780 0.3420 1.8100 1.1940 ;
    LAYER M1 ;
      RECT 1.7780 1.6860 1.8100 2.5380 ;
    LAYER M1 ;
      RECT 1.7780 3.0300 1.8100 3.8820 ;
    LAYER M1 ;
      RECT 1.7780 4.3740 1.8100 5.2260 ;
    LAYER M1 ;
      RECT 1.8560 0.3420 1.8880 1.1940 ;
    LAYER M1 ;
      RECT 1.8560 1.3020 1.8880 1.5780 ;
    LAYER M1 ;
      RECT 1.8560 1.6860 1.8880 2.5380 ;
    LAYER M1 ;
      RECT 1.8560 2.6460 1.8880 2.9220 ;
    LAYER M1 ;
      RECT 1.8560 3.0300 1.8880 3.8820 ;
    LAYER M1 ;
      RECT 1.8560 3.9900 1.8880 4.2660 ;
    LAYER M1 ;
      RECT 1.8560 4.3740 1.8880 5.2260 ;
    LAYER M1 ;
      RECT 1.8560 5.3340 1.8880 5.6100 ;
    LAYER M1 ;
      RECT 1.8560 5.8140 1.8880 6.1860 ;
    LAYER M1 ;
      RECT 1.9340 0.3420 1.9660 1.1940 ;
    LAYER M1 ;
      RECT 1.9340 1.6860 1.9660 2.5380 ;
    LAYER M1 ;
      RECT 1.9340 3.0300 1.9660 3.8820 ;
    LAYER M1 ;
      RECT 1.9340 4.3740 1.9660 5.2260 ;
    LAYER M1 ;
      RECT 2.0120 0.3420 2.0440 1.1940 ;
    LAYER M1 ;
      RECT 2.0120 1.3020 2.0440 1.5780 ;
    LAYER M1 ;
      RECT 2.0120 1.6860 2.0440 2.5380 ;
    LAYER M1 ;
      RECT 2.0120 2.6460 2.0440 2.9220 ;
    LAYER M1 ;
      RECT 2.0120 3.0300 2.0440 3.8820 ;
    LAYER M1 ;
      RECT 2.0120 3.9900 2.0440 4.2660 ;
    LAYER M1 ;
      RECT 2.0120 4.3740 2.0440 5.2260 ;
    LAYER M1 ;
      RECT 2.0120 5.3340 2.0440 5.6100 ;
    LAYER M1 ;
      RECT 2.0900 0.3420 2.1220 1.1940 ;
    LAYER M1 ;
      RECT 2.0900 1.6860 2.1220 2.5380 ;
    LAYER M1 ;
      RECT 2.0900 3.0300 2.1220 3.8820 ;
    LAYER M1 ;
      RECT 2.0900 4.3740 2.1220 5.2260 ;
    LAYER M2 ;
      RECT 0.8160 1.3280 2.0700 1.3600 ;
    LAYER M2 ;
      RECT 0.8160 0.3680 2.0700 0.4000 ;
    LAYER M2 ;
      RECT 0.7380 0.4640 2.1480 0.4960 ;
    LAYER M2 ;
      RECT 0.9720 0.5600 1.9140 0.5920 ;
    LAYER M2 ;
      RECT 0.9720 1.4240 1.9140 1.4560 ;
    LAYER M2 ;
      RECT 0.9720 2.6720 1.9140 2.7040 ;
    LAYER M2 ;
      RECT 0.9720 1.7120 1.9140 1.7440 ;
    LAYER M2 ;
      RECT 0.7380 1.8080 2.1480 1.8400 ;
    LAYER M2 ;
      RECT 0.8160 1.9040 2.0700 1.9360 ;
    LAYER M2 ;
      RECT 0.8160 2.7680 2.0700 2.8000 ;
    LAYER M2 ;
      RECT 0.8160 4.0160 2.0700 4.0480 ;
    LAYER M2 ;
      RECT 0.8160 3.0560 2.0700 3.0880 ;
    LAYER M2 ;
      RECT 0.7380 3.1520 2.1480 3.1840 ;
    LAYER M2 ;
      RECT 0.9720 3.2480 1.9140 3.2800 ;
    LAYER M2 ;
      RECT 0.9720 4.1120 1.9140 4.1440 ;
    LAYER M2 ;
      RECT 0.9720 5.3600 1.9140 5.3920 ;
    LAYER M2 ;
      RECT 0.9720 4.4000 1.9140 4.4320 ;
    LAYER M2 ;
      RECT 0.7380 4.4960 2.1480 4.5280 ;
    LAYER M2 ;
      RECT 0.8160 4.5920 2.0700 4.6240 ;
    LAYER M2 ;
      RECT 0.8160 5.4560 2.0700 5.4880 ;
    LAYER V1 ;
      RECT 0.9200 0.3680 0.9520 0.4000 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 1.9040 0.9520 1.9360 ;
    LAYER V1 ;
      RECT 0.9200 2.7680 0.9520 2.8000 ;
    LAYER V1 ;
      RECT 0.9200 3.0560 0.9520 3.0880 ;
    LAYER V1 ;
      RECT 0.9200 4.0160 0.9520 4.0480 ;
    LAYER V1 ;
      RECT 0.9200 4.5920 0.9520 4.6240 ;
    LAYER V1 ;
      RECT 0.9200 5.4560 0.9520 5.4880 ;
    LAYER V1 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V1 ;
      RECT 1.3880 0.3680 1.4200 0.4000 ;
    LAYER V1 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V1 ;
      RECT 1.3880 1.9040 1.4200 1.9360 ;
    LAYER V1 ;
      RECT 1.3880 2.7680 1.4200 2.8000 ;
    LAYER V1 ;
      RECT 1.3880 3.0560 1.4200 3.0880 ;
    LAYER V1 ;
      RECT 1.3880 4.0160 1.4200 4.0480 ;
    LAYER V1 ;
      RECT 1.3880 4.5920 1.4200 4.6240 ;
    LAYER V1 ;
      RECT 1.3880 5.4560 1.4200 5.4880 ;
    LAYER V1 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V1 ;
      RECT 1.8560 0.5600 1.8880 0.5920 ;
    LAYER V1 ;
      RECT 1.8560 1.4240 1.8880 1.4560 ;
    LAYER V1 ;
      RECT 1.8560 1.7120 1.8880 1.7440 ;
    LAYER V1 ;
      RECT 1.8560 2.6720 1.8880 2.7040 ;
    LAYER V1 ;
      RECT 1.8560 3.2480 1.8880 3.2800 ;
    LAYER V1 ;
      RECT 1.8560 4.1120 1.8880 4.1440 ;
    LAYER V1 ;
      RECT 1.8560 4.4000 1.8880 4.4320 ;
    LAYER V1 ;
      RECT 1.8560 5.3600 1.8880 5.3920 ;
    LAYER V1 ;
      RECT 1.8560 6.0320 1.8880 6.0640 ;
    LAYER V1 ;
      RECT 2.0120 0.3680 2.0440 0.4000 ;
    LAYER V1 ;
      RECT 2.0120 1.3280 2.0440 1.3600 ;
    LAYER V1 ;
      RECT 2.0120 1.9040 2.0440 1.9360 ;
    LAYER V1 ;
      RECT 2.0120 2.7680 2.0440 2.8000 ;
    LAYER V1 ;
      RECT 2.0120 3.0560 2.0440 3.0880 ;
    LAYER V1 ;
      RECT 2.0120 4.0160 2.0440 4.0480 ;
    LAYER V1 ;
      RECT 2.0120 4.5920 2.0440 4.6240 ;
    LAYER V1 ;
      RECT 2.0120 5.4560 2.0440 5.4880 ;
    LAYER V1 ;
      RECT 1.5440 0.3680 1.5760 0.4000 ;
    LAYER V1 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V1 ;
      RECT 1.5440 1.9040 1.5760 1.9360 ;
    LAYER V1 ;
      RECT 1.5440 2.7680 1.5760 2.8000 ;
    LAYER V1 ;
      RECT 1.5440 3.0560 1.5760 3.0880 ;
    LAYER V1 ;
      RECT 1.5440 4.0160 1.5760 4.0480 ;
    LAYER V1 ;
      RECT 1.5440 4.5920 1.5760 4.6240 ;
    LAYER V1 ;
      RECT 1.5440 5.4560 1.5760 5.4880 ;
    LAYER V1 ;
      RECT 0.8420 0.4640 0.8740 0.4960 ;
    LAYER V1 ;
      RECT 0.8420 1.8080 0.8740 1.8400 ;
    LAYER V1 ;
      RECT 0.8420 3.1520 0.8740 3.1840 ;
    LAYER V1 ;
      RECT 0.8420 4.4960 0.8740 4.5280 ;
    LAYER V1 ;
      RECT 0.9980 0.4640 1.0300 0.4960 ;
    LAYER V1 ;
      RECT 0.9980 1.8080 1.0300 1.8400 ;
    LAYER V1 ;
      RECT 0.9980 3.1520 1.0300 3.1840 ;
    LAYER V1 ;
      RECT 0.9980 4.4960 1.0300 4.5280 ;
    LAYER V1 ;
      RECT 1.1540 0.4640 1.1860 0.4960 ;
    LAYER V1 ;
      RECT 1.1540 1.8080 1.1860 1.8400 ;
    LAYER V1 ;
      RECT 1.1540 3.1520 1.1860 3.1840 ;
    LAYER V1 ;
      RECT 1.1540 4.4960 1.1860 4.5280 ;
    LAYER V1 ;
      RECT 1.3100 0.4640 1.3420 0.4960 ;
    LAYER V1 ;
      RECT 1.3100 1.8080 1.3420 1.8400 ;
    LAYER V1 ;
      RECT 1.3100 3.1520 1.3420 3.1840 ;
    LAYER V1 ;
      RECT 1.3100 4.4960 1.3420 4.5280 ;
    LAYER V1 ;
      RECT 1.4660 0.4640 1.4980 0.4960 ;
    LAYER V1 ;
      RECT 1.4660 1.8080 1.4980 1.8400 ;
    LAYER V1 ;
      RECT 1.4660 3.1520 1.4980 3.1840 ;
    LAYER V1 ;
      RECT 1.4660 4.4960 1.4980 4.5280 ;
    LAYER V1 ;
      RECT 1.6220 0.4640 1.6540 0.4960 ;
    LAYER V1 ;
      RECT 1.6220 1.8080 1.6540 1.8400 ;
    LAYER V1 ;
      RECT 1.6220 3.1520 1.6540 3.1840 ;
    LAYER V1 ;
      RECT 1.6220 4.4960 1.6540 4.5280 ;
    LAYER V1 ;
      RECT 1.7780 0.4640 1.8100 0.4960 ;
    LAYER V1 ;
      RECT 1.7780 1.8080 1.8100 1.8400 ;
    LAYER V1 ;
      RECT 1.7780 3.1520 1.8100 3.1840 ;
    LAYER V1 ;
      RECT 1.7780 4.4960 1.8100 4.5280 ;
    LAYER V1 ;
      RECT 1.9340 0.4640 1.9660 0.4960 ;
    LAYER V1 ;
      RECT 1.9340 1.8080 1.9660 1.8400 ;
    LAYER V1 ;
      RECT 1.9340 3.1520 1.9660 3.1840 ;
    LAYER V1 ;
      RECT 1.9340 4.4960 1.9660 4.5280 ;
    LAYER V1 ;
      RECT 2.0900 0.4640 2.1220 0.4960 ;
    LAYER V1 ;
      RECT 2.0900 1.8080 2.1220 1.8400 ;
    LAYER V1 ;
      RECT 2.0900 3.1520 2.1220 3.1840 ;
    LAYER V1 ;
      RECT 2.0900 4.4960 2.1220 4.5280 ;
    LAYER V1 ;
      RECT 1.2320 0.5600 1.2640 0.5920 ;
    LAYER V1 ;
      RECT 1.2320 1.4240 1.2640 1.4560 ;
    LAYER V1 ;
      RECT 1.2320 1.7120 1.2640 1.7440 ;
    LAYER V1 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V1 ;
      RECT 1.2320 3.2480 1.2640 3.2800 ;
    LAYER V1 ;
      RECT 1.2320 4.1120 1.2640 4.1440 ;
    LAYER V1 ;
      RECT 1.2320 4.4000 1.2640 4.4320 ;
    LAYER V1 ;
      RECT 1.2320 5.3600 1.2640 5.3920 ;
    LAYER V1 ;
      RECT 1.0760 0.5600 1.1080 0.5920 ;
    LAYER V1 ;
      RECT 1.0760 1.4240 1.1080 1.4560 ;
    LAYER V1 ;
      RECT 1.0760 1.7120 1.1080 1.7440 ;
    LAYER V1 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V1 ;
      RECT 1.0760 3.2480 1.1080 3.2800 ;
    LAYER V1 ;
      RECT 1.0760 4.1120 1.1080 4.1440 ;
    LAYER V1 ;
      RECT 1.0760 4.4000 1.1080 4.4320 ;
    LAYER V1 ;
      RECT 1.0760 5.3600 1.1080 5.3920 ;
    LAYER V1 ;
      RECT 1.7000 0.5600 1.7320 0.5920 ;
    LAYER V1 ;
      RECT 1.7000 1.4240 1.7320 1.4560 ;
    LAYER V1 ;
      RECT 1.7000 1.7120 1.7320 1.7440 ;
    LAYER V1 ;
      RECT 1.7000 2.6720 1.7320 2.7040 ;
    LAYER V1 ;
      RECT 1.7000 3.2480 1.7320 3.2800 ;
    LAYER V1 ;
      RECT 1.7000 4.1120 1.7320 4.1440 ;
    LAYER V1 ;
      RECT 1.7000 4.4000 1.7320 4.4320 ;
    LAYER V1 ;
      RECT 1.7000 5.3600 1.7320 5.3920 ;
    LAYER V2 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V2 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V2 ;
      RECT 1.2320 4.0160 1.2640 4.0480 ;
    LAYER V2 ;
      RECT 1.2320 5.3600 1.2640 5.3920 ;
    LAYER V2 ;
      RECT 1.3100 0.3680 1.3420 0.4000 ;
    LAYER V2 ;
      RECT 1.3100 1.7120 1.3420 1.7440 ;
    LAYER V2 ;
      RECT 1.3100 3.0560 1.3420 3.0880 ;
    LAYER V2 ;
      RECT 1.3100 4.4000 1.3420 4.4320 ;
    LAYER V2 ;
      RECT 1.3880 0.4640 1.4200 0.4960 ;
    LAYER V2 ;
      RECT 1.3880 1.8080 1.4200 1.8400 ;
    LAYER V2 ;
      RECT 1.3880 3.1520 1.4200 3.1840 ;
    LAYER V2 ;
      RECT 1.3880 4.4960 1.4200 4.5280 ;
    LAYER V2 ;
      RECT 1.4660 0.5600 1.4980 0.5920 ;
    LAYER V2 ;
      RECT 1.4660 1.9040 1.4980 1.9360 ;
    LAYER V2 ;
      RECT 1.4660 3.2480 1.4980 3.2800 ;
    LAYER V2 ;
      RECT 1.4660 4.5920 1.4980 4.6240 ;
    LAYER V2 ;
      RECT 1.5440 1.4240 1.5760 1.4560 ;
    LAYER V2 ;
      RECT 1.5440 2.7680 1.5760 2.8000 ;
    LAYER V2 ;
      RECT 1.5440 4.1120 1.5760 4.1440 ;
    LAYER V2 ;
      RECT 1.5440 5.4560 1.5760 5.4880 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.5840 0.9520 3.6160 ;
    LAYER V0 ;
      RECT 0.9200 3.7280 0.9520 3.7600 ;
    LAYER V0 ;
      RECT 0.9200 4.0160 0.9520 4.0480 ;
    LAYER V0 ;
      RECT 0.9200 4.9280 0.9520 4.9600 ;
    LAYER V0 ;
      RECT 0.9200 5.0720 0.9520 5.1040 ;
    LAYER V0 ;
      RECT 0.9200 5.3600 0.9520 5.3920 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.8420 3.4400 0.8740 3.4720 ;
    LAYER V0 ;
      RECT 0.8420 3.5840 0.8740 3.6160 ;
    LAYER V0 ;
      RECT 0.8420 3.7280 0.8740 3.7600 ;
    LAYER V0 ;
      RECT 0.8420 4.7840 0.8740 4.8160 ;
    LAYER V0 ;
      RECT 0.8420 4.9280 0.8740 4.9600 ;
    LAYER V0 ;
      RECT 0.8420 5.0720 0.8740 5.1040 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 3.4400 1.0300 3.4720 ;
    LAYER V0 ;
      RECT 0.9980 3.4400 1.0300 3.4720 ;
    LAYER V0 ;
      RECT 0.9980 3.5840 1.0300 3.6160 ;
    LAYER V0 ;
      RECT 0.9980 3.5840 1.0300 3.6160 ;
    LAYER V0 ;
      RECT 0.9980 3.7280 1.0300 3.7600 ;
    LAYER V0 ;
      RECT 0.9980 3.7280 1.0300 3.7600 ;
    LAYER V0 ;
      RECT 0.9980 4.7840 1.0300 4.8160 ;
    LAYER V0 ;
      RECT 0.9980 4.7840 1.0300 4.8160 ;
    LAYER V0 ;
      RECT 0.9980 4.9280 1.0300 4.9600 ;
    LAYER V0 ;
      RECT 0.9980 4.9280 1.0300 4.9600 ;
    LAYER V0 ;
      RECT 0.9980 5.0720 1.0300 5.1040 ;
    LAYER V0 ;
      RECT 0.9980 5.0720 1.0300 5.1040 ;
    LAYER V0 ;
      RECT 1.0760 0.7520 1.1080 0.7840 ;
    LAYER V0 ;
      RECT 1.0760 1.0400 1.1080 1.0720 ;
    LAYER V0 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V0 ;
      RECT 1.0760 2.0960 1.1080 2.1280 ;
    LAYER V0 ;
      RECT 1.0760 2.3840 1.1080 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V0 ;
      RECT 1.0760 3.4400 1.1080 3.4720 ;
    LAYER V0 ;
      RECT 1.0760 3.7280 1.1080 3.7600 ;
    LAYER V0 ;
      RECT 1.0760 4.0160 1.1080 4.0480 ;
    LAYER V0 ;
      RECT 1.0760 4.7840 1.1080 4.8160 ;
    LAYER V0 ;
      RECT 1.0760 5.0720 1.1080 5.1040 ;
    LAYER V0 ;
      RECT 1.0760 5.3600 1.1080 5.3920 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.1540 3.4400 1.1860 3.4720 ;
    LAYER V0 ;
      RECT 1.1540 3.4400 1.1860 3.4720 ;
    LAYER V0 ;
      RECT 1.1540 3.5840 1.1860 3.6160 ;
    LAYER V0 ;
      RECT 1.1540 3.5840 1.1860 3.6160 ;
    LAYER V0 ;
      RECT 1.1540 3.7280 1.1860 3.7600 ;
    LAYER V0 ;
      RECT 1.1540 3.7280 1.1860 3.7600 ;
    LAYER V0 ;
      RECT 1.1540 4.7840 1.1860 4.8160 ;
    LAYER V0 ;
      RECT 1.1540 4.7840 1.1860 4.8160 ;
    LAYER V0 ;
      RECT 1.1540 4.9280 1.1860 4.9600 ;
    LAYER V0 ;
      RECT 1.1540 4.9280 1.1860 4.9600 ;
    LAYER V0 ;
      RECT 1.1540 5.0720 1.1860 5.1040 ;
    LAYER V0 ;
      RECT 1.1540 5.0720 1.1860 5.1040 ;
    LAYER V0 ;
      RECT 1.2320 0.7520 1.2640 0.7840 ;
    LAYER V0 ;
      RECT 1.2320 0.8960 1.2640 0.9280 ;
    LAYER V0 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V0 ;
      RECT 1.2320 2.0960 1.2640 2.1280 ;
    LAYER V0 ;
      RECT 1.2320 2.2400 1.2640 2.2720 ;
    LAYER V0 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V0 ;
      RECT 1.2320 3.4400 1.2640 3.4720 ;
    LAYER V0 ;
      RECT 1.2320 3.5840 1.2640 3.6160 ;
    LAYER V0 ;
      RECT 1.2320 4.0160 1.2640 4.0480 ;
    LAYER V0 ;
      RECT 1.2320 4.7840 1.2640 4.8160 ;
    LAYER V0 ;
      RECT 1.2320 4.9280 1.2640 4.9600 ;
    LAYER V0 ;
      RECT 1.2320 5.3600 1.2640 5.3920 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3100 3.4400 1.3420 3.4720 ;
    LAYER V0 ;
      RECT 1.3100 3.4400 1.3420 3.4720 ;
    LAYER V0 ;
      RECT 1.3100 3.5840 1.3420 3.6160 ;
    LAYER V0 ;
      RECT 1.3100 3.5840 1.3420 3.6160 ;
    LAYER V0 ;
      RECT 1.3100 3.7280 1.3420 3.7600 ;
    LAYER V0 ;
      RECT 1.3100 3.7280 1.3420 3.7600 ;
    LAYER V0 ;
      RECT 1.3100 4.7840 1.3420 4.8160 ;
    LAYER V0 ;
      RECT 1.3100 4.7840 1.3420 4.8160 ;
    LAYER V0 ;
      RECT 1.3100 4.9280 1.3420 4.9600 ;
    LAYER V0 ;
      RECT 1.3100 4.9280 1.3420 4.9600 ;
    LAYER V0 ;
      RECT 1.3100 5.0720 1.3420 5.1040 ;
    LAYER V0 ;
      RECT 1.3100 5.0720 1.3420 5.1040 ;
    LAYER V0 ;
      RECT 1.3880 0.8960 1.4200 0.9280 ;
    LAYER V0 ;
      RECT 1.3880 1.0400 1.4200 1.0720 ;
    LAYER V0 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V0 ;
      RECT 1.3880 2.2400 1.4200 2.2720 ;
    LAYER V0 ;
      RECT 1.3880 2.3840 1.4200 2.4160 ;
    LAYER V0 ;
      RECT 1.3880 2.6720 1.4200 2.7040 ;
    LAYER V0 ;
      RECT 1.3880 3.5840 1.4200 3.6160 ;
    LAYER V0 ;
      RECT 1.3880 3.7280 1.4200 3.7600 ;
    LAYER V0 ;
      RECT 1.3880 4.0160 1.4200 4.0480 ;
    LAYER V0 ;
      RECT 1.3880 4.9280 1.4200 4.9600 ;
    LAYER V0 ;
      RECT 1.3880 5.0720 1.4200 5.1040 ;
    LAYER V0 ;
      RECT 1.3880 5.3600 1.4200 5.3920 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
    LAYER V0 ;
      RECT 1.4660 3.4400 1.4980 3.4720 ;
    LAYER V0 ;
      RECT 1.4660 3.4400 1.4980 3.4720 ;
    LAYER V0 ;
      RECT 1.4660 3.5840 1.4980 3.6160 ;
    LAYER V0 ;
      RECT 1.4660 3.5840 1.4980 3.6160 ;
    LAYER V0 ;
      RECT 1.4660 3.7280 1.4980 3.7600 ;
    LAYER V0 ;
      RECT 1.4660 3.7280 1.4980 3.7600 ;
    LAYER V0 ;
      RECT 1.4660 4.7840 1.4980 4.8160 ;
    LAYER V0 ;
      RECT 1.4660 4.7840 1.4980 4.8160 ;
    LAYER V0 ;
      RECT 1.4660 4.9280 1.4980 4.9600 ;
    LAYER V0 ;
      RECT 1.4660 4.9280 1.4980 4.9600 ;
    LAYER V0 ;
      RECT 1.4660 5.0720 1.4980 5.1040 ;
    LAYER V0 ;
      RECT 1.4660 5.0720 1.4980 5.1040 ;
    LAYER V0 ;
      RECT 1.5440 0.7520 1.5760 0.7840 ;
    LAYER V0 ;
      RECT 1.5440 1.0400 1.5760 1.0720 ;
    LAYER V0 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V0 ;
      RECT 1.5440 2.0960 1.5760 2.1280 ;
    LAYER V0 ;
      RECT 1.5440 2.3840 1.5760 2.4160 ;
    LAYER V0 ;
      RECT 1.5440 2.6720 1.5760 2.7040 ;
    LAYER V0 ;
      RECT 1.5440 3.4400 1.5760 3.4720 ;
    LAYER V0 ;
      RECT 1.5440 3.7280 1.5760 3.7600 ;
    LAYER V0 ;
      RECT 1.5440 4.0160 1.5760 4.0480 ;
    LAYER V0 ;
      RECT 1.5440 4.7840 1.5760 4.8160 ;
    LAYER V0 ;
      RECT 1.5440 5.0720 1.5760 5.1040 ;
    LAYER V0 ;
      RECT 1.5440 5.3600 1.5760 5.3920 ;
    LAYER V0 ;
      RECT 1.6220 0.7520 1.6540 0.7840 ;
    LAYER V0 ;
      RECT 1.6220 0.7520 1.6540 0.7840 ;
    LAYER V0 ;
      RECT 1.6220 0.8960 1.6540 0.9280 ;
    LAYER V0 ;
      RECT 1.6220 0.8960 1.6540 0.9280 ;
    LAYER V0 ;
      RECT 1.6220 1.0400 1.6540 1.0720 ;
    LAYER V0 ;
      RECT 1.6220 1.0400 1.6540 1.0720 ;
    LAYER V0 ;
      RECT 1.6220 2.0960 1.6540 2.1280 ;
    LAYER V0 ;
      RECT 1.6220 2.0960 1.6540 2.1280 ;
    LAYER V0 ;
      RECT 1.6220 2.2400 1.6540 2.2720 ;
    LAYER V0 ;
      RECT 1.6220 2.2400 1.6540 2.2720 ;
    LAYER V0 ;
      RECT 1.6220 2.3840 1.6540 2.4160 ;
    LAYER V0 ;
      RECT 1.6220 2.3840 1.6540 2.4160 ;
    LAYER V0 ;
      RECT 1.6220 3.4400 1.6540 3.4720 ;
    LAYER V0 ;
      RECT 1.6220 3.4400 1.6540 3.4720 ;
    LAYER V0 ;
      RECT 1.6220 3.5840 1.6540 3.6160 ;
    LAYER V0 ;
      RECT 1.6220 3.5840 1.6540 3.6160 ;
    LAYER V0 ;
      RECT 1.6220 3.7280 1.6540 3.7600 ;
    LAYER V0 ;
      RECT 1.6220 3.7280 1.6540 3.7600 ;
    LAYER V0 ;
      RECT 1.6220 4.7840 1.6540 4.8160 ;
    LAYER V0 ;
      RECT 1.6220 4.7840 1.6540 4.8160 ;
    LAYER V0 ;
      RECT 1.6220 4.9280 1.6540 4.9600 ;
    LAYER V0 ;
      RECT 1.6220 4.9280 1.6540 4.9600 ;
    LAYER V0 ;
      RECT 1.6220 5.0720 1.6540 5.1040 ;
    LAYER V0 ;
      RECT 1.6220 5.0720 1.6540 5.1040 ;
    LAYER V0 ;
      RECT 1.7000 0.7520 1.7320 0.7840 ;
    LAYER V0 ;
      RECT 1.7000 0.8960 1.7320 0.9280 ;
    LAYER V0 ;
      RECT 1.7000 1.3280 1.7320 1.3600 ;
    LAYER V0 ;
      RECT 1.7000 2.0960 1.7320 2.1280 ;
    LAYER V0 ;
      RECT 1.7000 2.2400 1.7320 2.2720 ;
    LAYER V0 ;
      RECT 1.7000 2.6720 1.7320 2.7040 ;
    LAYER V0 ;
      RECT 1.7000 3.4400 1.7320 3.4720 ;
    LAYER V0 ;
      RECT 1.7000 3.5840 1.7320 3.6160 ;
    LAYER V0 ;
      RECT 1.7000 4.0160 1.7320 4.0480 ;
    LAYER V0 ;
      RECT 1.7000 4.7840 1.7320 4.8160 ;
    LAYER V0 ;
      RECT 1.7000 4.9280 1.7320 4.9600 ;
    LAYER V0 ;
      RECT 1.7000 5.3600 1.7320 5.3920 ;
    LAYER V0 ;
      RECT 1.7780 0.7520 1.8100 0.7840 ;
    LAYER V0 ;
      RECT 1.7780 0.7520 1.8100 0.7840 ;
    LAYER V0 ;
      RECT 1.7780 0.8960 1.8100 0.9280 ;
    LAYER V0 ;
      RECT 1.7780 0.8960 1.8100 0.9280 ;
    LAYER V0 ;
      RECT 1.7780 1.0400 1.8100 1.0720 ;
    LAYER V0 ;
      RECT 1.7780 1.0400 1.8100 1.0720 ;
    LAYER V0 ;
      RECT 1.7780 2.0960 1.8100 2.1280 ;
    LAYER V0 ;
      RECT 1.7780 2.0960 1.8100 2.1280 ;
    LAYER V0 ;
      RECT 1.7780 2.2400 1.8100 2.2720 ;
    LAYER V0 ;
      RECT 1.7780 2.2400 1.8100 2.2720 ;
    LAYER V0 ;
      RECT 1.7780 2.3840 1.8100 2.4160 ;
    LAYER V0 ;
      RECT 1.7780 2.3840 1.8100 2.4160 ;
    LAYER V0 ;
      RECT 1.7780 3.4400 1.8100 3.4720 ;
    LAYER V0 ;
      RECT 1.7780 3.4400 1.8100 3.4720 ;
    LAYER V0 ;
      RECT 1.7780 3.5840 1.8100 3.6160 ;
    LAYER V0 ;
      RECT 1.7780 3.5840 1.8100 3.6160 ;
    LAYER V0 ;
      RECT 1.7780 3.7280 1.8100 3.7600 ;
    LAYER V0 ;
      RECT 1.7780 3.7280 1.8100 3.7600 ;
    LAYER V0 ;
      RECT 1.7780 4.7840 1.8100 4.8160 ;
    LAYER V0 ;
      RECT 1.7780 4.7840 1.8100 4.8160 ;
    LAYER V0 ;
      RECT 1.7780 4.9280 1.8100 4.9600 ;
    LAYER V0 ;
      RECT 1.7780 4.9280 1.8100 4.9600 ;
    LAYER V0 ;
      RECT 1.7780 5.0720 1.8100 5.1040 ;
    LAYER V0 ;
      RECT 1.7780 5.0720 1.8100 5.1040 ;
    LAYER V0 ;
      RECT 1.8560 0.8960 1.8880 0.9280 ;
    LAYER V0 ;
      RECT 1.8560 1.0400 1.8880 1.0720 ;
    LAYER V0 ;
      RECT 1.8560 1.3280 1.8880 1.3600 ;
    LAYER V0 ;
      RECT 1.8560 2.2400 1.8880 2.2720 ;
    LAYER V0 ;
      RECT 1.8560 2.3840 1.8880 2.4160 ;
    LAYER V0 ;
      RECT 1.8560 2.6720 1.8880 2.7040 ;
    LAYER V0 ;
      RECT 1.8560 3.5840 1.8880 3.6160 ;
    LAYER V0 ;
      RECT 1.8560 3.7280 1.8880 3.7600 ;
    LAYER V0 ;
      RECT 1.8560 4.0160 1.8880 4.0480 ;
    LAYER V0 ;
      RECT 1.8560 4.9280 1.8880 4.9600 ;
    LAYER V0 ;
      RECT 1.8560 5.0720 1.8880 5.1040 ;
    LAYER V0 ;
      RECT 1.8560 5.3600 1.8880 5.3920 ;
    LAYER V0 ;
      RECT 1.8560 6.0320 1.8880 6.0640 ;
    LAYER V0 ;
      RECT 1.8560 6.0320 1.8880 6.0640 ;
    LAYER V0 ;
      RECT 1.8560 6.0320 1.8880 6.0640 ;
    LAYER V0 ;
      RECT 1.8560 6.0320 1.8880 6.0640 ;
    LAYER V0 ;
      RECT 1.9340 0.7520 1.9660 0.7840 ;
    LAYER V0 ;
      RECT 1.9340 0.7520 1.9660 0.7840 ;
    LAYER V0 ;
      RECT 1.9340 0.8960 1.9660 0.9280 ;
    LAYER V0 ;
      RECT 1.9340 0.8960 1.9660 0.9280 ;
    LAYER V0 ;
      RECT 1.9340 1.0400 1.9660 1.0720 ;
    LAYER V0 ;
      RECT 1.9340 1.0400 1.9660 1.0720 ;
    LAYER V0 ;
      RECT 1.9340 2.0960 1.9660 2.1280 ;
    LAYER V0 ;
      RECT 1.9340 2.0960 1.9660 2.1280 ;
    LAYER V0 ;
      RECT 1.9340 2.2400 1.9660 2.2720 ;
    LAYER V0 ;
      RECT 1.9340 2.2400 1.9660 2.2720 ;
    LAYER V0 ;
      RECT 1.9340 2.3840 1.9660 2.4160 ;
    LAYER V0 ;
      RECT 1.9340 2.3840 1.9660 2.4160 ;
    LAYER V0 ;
      RECT 1.9340 3.4400 1.9660 3.4720 ;
    LAYER V0 ;
      RECT 1.9340 3.4400 1.9660 3.4720 ;
    LAYER V0 ;
      RECT 1.9340 3.5840 1.9660 3.6160 ;
    LAYER V0 ;
      RECT 1.9340 3.5840 1.9660 3.6160 ;
    LAYER V0 ;
      RECT 1.9340 3.7280 1.9660 3.7600 ;
    LAYER V0 ;
      RECT 1.9340 3.7280 1.9660 3.7600 ;
    LAYER V0 ;
      RECT 1.9340 4.7840 1.9660 4.8160 ;
    LAYER V0 ;
      RECT 1.9340 4.7840 1.9660 4.8160 ;
    LAYER V0 ;
      RECT 1.9340 4.9280 1.9660 4.9600 ;
    LAYER V0 ;
      RECT 1.9340 4.9280 1.9660 4.9600 ;
    LAYER V0 ;
      RECT 1.9340 5.0720 1.9660 5.1040 ;
    LAYER V0 ;
      RECT 1.9340 5.0720 1.9660 5.1040 ;
    LAYER V0 ;
      RECT 2.0120 0.7520 2.0440 0.7840 ;
    LAYER V0 ;
      RECT 2.0120 1.0400 2.0440 1.0720 ;
    LAYER V0 ;
      RECT 2.0120 1.3280 2.0440 1.3600 ;
    LAYER V0 ;
      RECT 2.0120 2.0960 2.0440 2.1280 ;
    LAYER V0 ;
      RECT 2.0120 2.3840 2.0440 2.4160 ;
    LAYER V0 ;
      RECT 2.0120 2.6720 2.0440 2.7040 ;
    LAYER V0 ;
      RECT 2.0120 3.4400 2.0440 3.4720 ;
    LAYER V0 ;
      RECT 2.0120 3.7280 2.0440 3.7600 ;
    LAYER V0 ;
      RECT 2.0120 4.0160 2.0440 4.0480 ;
    LAYER V0 ;
      RECT 2.0120 4.7840 2.0440 4.8160 ;
    LAYER V0 ;
      RECT 2.0120 5.0720 2.0440 5.1040 ;
    LAYER V0 ;
      RECT 2.0120 5.3600 2.0440 5.3920 ;
    LAYER V0 ;
      RECT 2.0900 0.7520 2.1220 0.7840 ;
    LAYER V0 ;
      RECT 2.0900 0.8960 2.1220 0.9280 ;
    LAYER V0 ;
      RECT 2.0900 1.0400 2.1220 1.0720 ;
    LAYER V0 ;
      RECT 2.0900 2.0960 2.1220 2.1280 ;
    LAYER V0 ;
      RECT 2.0900 2.2400 2.1220 2.2720 ;
    LAYER V0 ;
      RECT 2.0900 2.3840 2.1220 2.4160 ;
    LAYER V0 ;
      RECT 2.0900 3.4400 2.1220 3.4720 ;
    LAYER V0 ;
      RECT 2.0900 3.5840 2.1220 3.6160 ;
    LAYER V0 ;
      RECT 2.0900 3.7280 2.1220 3.7600 ;
    LAYER V0 ;
      RECT 2.0900 4.7840 2.1220 4.8160 ;
    LAYER V0 ;
      RECT 2.0900 4.9280 2.1220 4.9600 ;
    LAYER V0 ;
      RECT 2.0900 5.0720 2.1220 5.1040 ;
  END
END DP_NMOS_n12_X4_Y4
MACRO Switch_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X1_Y1 0 0 ;
  SIZE 1.8720 BY 2.6880 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 0.3680 1.0560 0.4000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 0.4640 0.9780 0.4960 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 1.3280 0.9780 1.3600 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 2.0000 1.2060 2.0320 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.7820 0.9520 2.1540 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 2.0000 0.9520 2.0320 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.0000 0.9520 2.0320 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
  END
END Switch_NMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 1.8720 BY 2.6880 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 0.3680 1.0560 0.4000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 0.4640 0.9780 0.4960 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7380 1.3280 0.9780 1.3600 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 2.0000 1.2060 2.0320 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.7820 0.9520 2.1540 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 2.0000 0.9520 2.0320 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.0000 0.9520 2.0320 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_NMOS_n12_X4_Y4
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X4_Y4 0 0 ;
  SIZE 2.3400 BY 6.7200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9980 0.3420 1.0300 4.4580 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.0760 0.4380 1.1080 4.5540 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1540 1.3020 1.1860 5.4180 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 6.0320 1.6740 6.0640 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.0300 0.9520 3.8820 ;
    LAYER M1 ;
      RECT 0.9200 3.9900 0.9520 4.2660 ;
    LAYER M1 ;
      RECT 0.9200 4.3740 0.9520 5.2260 ;
    LAYER M1 ;
      RECT 0.9200 5.3340 0.9520 5.6100 ;
    LAYER M1 ;
      RECT 0.9200 5.8140 0.9520 6.1860 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.8420 3.0300 0.8740 3.8820 ;
    LAYER M1 ;
      RECT 0.8420 4.3740 0.8740 5.2260 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 3.0300 1.0300 3.8820 ;
    LAYER M1 ;
      RECT 0.9980 4.3740 1.0300 5.2260 ;
    LAYER M1 ;
      RECT 1.0760 0.3420 1.1080 1.1940 ;
    LAYER M1 ;
      RECT 1.0760 1.3020 1.1080 1.5780 ;
    LAYER M1 ;
      RECT 1.0760 1.6860 1.1080 2.5380 ;
    LAYER M1 ;
      RECT 1.0760 2.6460 1.1080 2.9220 ;
    LAYER M1 ;
      RECT 1.0760 3.0300 1.1080 3.8820 ;
    LAYER M1 ;
      RECT 1.0760 3.9900 1.1080 4.2660 ;
    LAYER M1 ;
      RECT 1.0760 4.3740 1.1080 5.2260 ;
    LAYER M1 ;
      RECT 1.0760 5.3340 1.1080 5.6100 ;
    LAYER M1 ;
      RECT 1.1540 0.3420 1.1860 1.1940 ;
    LAYER M1 ;
      RECT 1.1540 1.6860 1.1860 2.5380 ;
    LAYER M1 ;
      RECT 1.1540 3.0300 1.1860 3.8820 ;
    LAYER M1 ;
      RECT 1.1540 4.3740 1.1860 5.2260 ;
    LAYER M1 ;
      RECT 1.2320 0.3420 1.2640 1.1940 ;
    LAYER M1 ;
      RECT 1.2320 1.3020 1.2640 1.5780 ;
    LAYER M1 ;
      RECT 1.2320 1.6860 1.2640 2.5380 ;
    LAYER M1 ;
      RECT 1.2320 2.6460 1.2640 2.9220 ;
    LAYER M1 ;
      RECT 1.2320 3.0300 1.2640 3.8820 ;
    LAYER M1 ;
      RECT 1.2320 3.9900 1.2640 4.2660 ;
    LAYER M1 ;
      RECT 1.2320 4.3740 1.2640 5.2260 ;
    LAYER M1 ;
      RECT 1.2320 5.3340 1.2640 5.6100 ;
    LAYER M1 ;
      RECT 1.3100 0.3420 1.3420 1.1940 ;
    LAYER M1 ;
      RECT 1.3100 1.6860 1.3420 2.5380 ;
    LAYER M1 ;
      RECT 1.3100 3.0300 1.3420 3.8820 ;
    LAYER M1 ;
      RECT 1.3100 4.3740 1.3420 5.2260 ;
    LAYER M1 ;
      RECT 1.3880 0.3420 1.4200 1.1940 ;
    LAYER M1 ;
      RECT 1.3880 1.3020 1.4200 1.5780 ;
    LAYER M1 ;
      RECT 1.3880 1.6860 1.4200 2.5380 ;
    LAYER M1 ;
      RECT 1.3880 2.6460 1.4200 2.9220 ;
    LAYER M1 ;
      RECT 1.3880 3.0300 1.4200 3.8820 ;
    LAYER M1 ;
      RECT 1.3880 3.9900 1.4200 4.2660 ;
    LAYER M1 ;
      RECT 1.3880 4.3740 1.4200 5.2260 ;
    LAYER M1 ;
      RECT 1.3880 5.3340 1.4200 5.6100 ;
    LAYER M1 ;
      RECT 1.3880 5.8140 1.4200 6.1860 ;
    LAYER M1 ;
      RECT 1.4660 0.3420 1.4980 1.1940 ;
    LAYER M1 ;
      RECT 1.4660 1.6860 1.4980 2.5380 ;
    LAYER M1 ;
      RECT 1.4660 3.0300 1.4980 3.8820 ;
    LAYER M1 ;
      RECT 1.4660 4.3740 1.4980 5.2260 ;
    LAYER M2 ;
      RECT 0.7380 0.3680 1.5240 0.4000 ;
    LAYER M2 ;
      RECT 0.8160 0.4640 1.4460 0.4960 ;
    LAYER M2 ;
      RECT 0.8160 1.3280 1.4460 1.3600 ;
    LAYER M2 ;
      RECT 0.7380 1.7120 1.5240 1.7440 ;
    LAYER M2 ;
      RECT 0.8160 1.8080 1.4460 1.8400 ;
    LAYER M2 ;
      RECT 0.8160 2.6720 1.4460 2.7040 ;
    LAYER M2 ;
      RECT 0.7380 3.0560 1.5240 3.0880 ;
    LAYER M2 ;
      RECT 0.8160 3.1520 1.4460 3.1840 ;
    LAYER M2 ;
      RECT 0.8160 4.0160 1.4460 4.0480 ;
    LAYER M2 ;
      RECT 0.7380 4.4000 1.5240 4.4320 ;
    LAYER M2 ;
      RECT 0.8160 4.4960 1.4460 4.5280 ;
    LAYER M2 ;
      RECT 0.8160 5.3600 1.4460 5.3920 ;
    LAYER V1 ;
      RECT 0.9200 0.4640 0.9520 0.4960 ;
    LAYER V1 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V1 ;
      RECT 0.9200 1.8080 0.9520 1.8400 ;
    LAYER V1 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 3.1520 0.9520 3.1840 ;
    LAYER V1 ;
      RECT 0.9200 4.0160 0.9520 4.0480 ;
    LAYER V1 ;
      RECT 0.9200 4.4960 0.9520 4.5280 ;
    LAYER V1 ;
      RECT 0.9200 5.3600 0.9520 5.3920 ;
    LAYER V1 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V1 ;
      RECT 1.3880 0.4640 1.4200 0.4960 ;
    LAYER V1 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V1 ;
      RECT 1.3880 1.8080 1.4200 1.8400 ;
    LAYER V1 ;
      RECT 1.3880 2.6720 1.4200 2.7040 ;
    LAYER V1 ;
      RECT 1.3880 3.1520 1.4200 3.1840 ;
    LAYER V1 ;
      RECT 1.3880 4.0160 1.4200 4.0480 ;
    LAYER V1 ;
      RECT 1.3880 4.4960 1.4200 4.5280 ;
    LAYER V1 ;
      RECT 1.3880 5.3600 1.4200 5.3920 ;
    LAYER V1 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.8420 1.7120 0.8740 1.7440 ;
    LAYER V1 ;
      RECT 0.8420 3.0560 0.8740 3.0880 ;
    LAYER V1 ;
      RECT 0.8420 4.4000 0.8740 4.4320 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V1 ;
      RECT 0.9980 3.0560 1.0300 3.0880 ;
    LAYER V1 ;
      RECT 0.9980 4.4000 1.0300 4.4320 ;
    LAYER V1 ;
      RECT 1.1540 0.3680 1.1860 0.4000 ;
    LAYER V1 ;
      RECT 1.1540 1.7120 1.1860 1.7440 ;
    LAYER V1 ;
      RECT 1.1540 3.0560 1.1860 3.0880 ;
    LAYER V1 ;
      RECT 1.1540 4.4000 1.1860 4.4320 ;
    LAYER V1 ;
      RECT 1.3100 0.3680 1.3420 0.4000 ;
    LAYER V1 ;
      RECT 1.3100 1.7120 1.3420 1.7440 ;
    LAYER V1 ;
      RECT 1.3100 3.0560 1.3420 3.0880 ;
    LAYER V1 ;
      RECT 1.3100 4.4000 1.3420 4.4320 ;
    LAYER V1 ;
      RECT 1.4660 0.3680 1.4980 0.4000 ;
    LAYER V1 ;
      RECT 1.4660 1.7120 1.4980 1.7440 ;
    LAYER V1 ;
      RECT 1.4660 3.0560 1.4980 3.0880 ;
    LAYER V1 ;
      RECT 1.4660 4.4000 1.4980 4.4320 ;
    LAYER V1 ;
      RECT 1.2320 0.4640 1.2640 0.4960 ;
    LAYER V1 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V1 ;
      RECT 1.2320 1.8080 1.2640 1.8400 ;
    LAYER V1 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V1 ;
      RECT 1.2320 3.1520 1.2640 3.1840 ;
    LAYER V1 ;
      RECT 1.2320 4.0160 1.2640 4.0480 ;
    LAYER V1 ;
      RECT 1.2320 4.4960 1.2640 4.5280 ;
    LAYER V1 ;
      RECT 1.2320 5.3600 1.2640 5.3920 ;
    LAYER V1 ;
      RECT 1.0760 0.4640 1.1080 0.4960 ;
    LAYER V1 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V1 ;
      RECT 1.0760 1.8080 1.1080 1.8400 ;
    LAYER V1 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V1 ;
      RECT 1.0760 3.1520 1.1080 3.1840 ;
    LAYER V1 ;
      RECT 1.0760 4.0160 1.1080 4.0480 ;
    LAYER V1 ;
      RECT 1.0760 4.4960 1.1080 4.5280 ;
    LAYER V1 ;
      RECT 1.0760 5.3600 1.1080 5.3920 ;
    LAYER V2 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V2 ;
      RECT 0.9980 1.7120 1.0300 1.7440 ;
    LAYER V2 ;
      RECT 0.9980 3.0560 1.0300 3.0880 ;
    LAYER V2 ;
      RECT 0.9980 4.4000 1.0300 4.4320 ;
    LAYER V2 ;
      RECT 1.0760 0.4640 1.1080 0.4960 ;
    LAYER V2 ;
      RECT 1.0760 1.8080 1.1080 1.8400 ;
    LAYER V2 ;
      RECT 1.0760 3.1520 1.1080 3.1840 ;
    LAYER V2 ;
      RECT 1.0760 4.4960 1.1080 4.5280 ;
    LAYER V2 ;
      RECT 1.1540 1.3280 1.1860 1.3600 ;
    LAYER V2 ;
      RECT 1.1540 2.6720 1.1860 2.7040 ;
    LAYER V2 ;
      RECT 1.1540 4.0160 1.1860 4.0480 ;
    LAYER V2 ;
      RECT 1.1540 5.3600 1.1860 5.3920 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.5840 0.9520 3.6160 ;
    LAYER V0 ;
      RECT 0.9200 3.7280 0.9520 3.7600 ;
    LAYER V0 ;
      RECT 0.9200 4.0160 0.9520 4.0480 ;
    LAYER V0 ;
      RECT 0.9200 4.9280 0.9520 4.9600 ;
    LAYER V0 ;
      RECT 0.9200 5.0720 0.9520 5.1040 ;
    LAYER V0 ;
      RECT 0.9200 5.3600 0.9520 5.3920 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.9200 6.0320 0.9520 6.0640 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.8420 3.4400 0.8740 3.4720 ;
    LAYER V0 ;
      RECT 0.8420 3.5840 0.8740 3.6160 ;
    LAYER V0 ;
      RECT 0.8420 3.7280 0.8740 3.7600 ;
    LAYER V0 ;
      RECT 0.8420 4.7840 0.8740 4.8160 ;
    LAYER V0 ;
      RECT 0.8420 4.9280 0.8740 4.9600 ;
    LAYER V0 ;
      RECT 0.8420 5.0720 0.8740 5.1040 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 3.4400 1.0300 3.4720 ;
    LAYER V0 ;
      RECT 0.9980 3.4400 1.0300 3.4720 ;
    LAYER V0 ;
      RECT 0.9980 3.5840 1.0300 3.6160 ;
    LAYER V0 ;
      RECT 0.9980 3.5840 1.0300 3.6160 ;
    LAYER V0 ;
      RECT 0.9980 3.7280 1.0300 3.7600 ;
    LAYER V0 ;
      RECT 0.9980 3.7280 1.0300 3.7600 ;
    LAYER V0 ;
      RECT 0.9980 4.7840 1.0300 4.8160 ;
    LAYER V0 ;
      RECT 0.9980 4.7840 1.0300 4.8160 ;
    LAYER V0 ;
      RECT 0.9980 4.9280 1.0300 4.9600 ;
    LAYER V0 ;
      RECT 0.9980 4.9280 1.0300 4.9600 ;
    LAYER V0 ;
      RECT 0.9980 5.0720 1.0300 5.1040 ;
    LAYER V0 ;
      RECT 0.9980 5.0720 1.0300 5.1040 ;
    LAYER V0 ;
      RECT 1.0760 0.7520 1.1080 0.7840 ;
    LAYER V0 ;
      RECT 1.0760 1.0400 1.1080 1.0720 ;
    LAYER V0 ;
      RECT 1.0760 1.3280 1.1080 1.3600 ;
    LAYER V0 ;
      RECT 1.0760 2.0960 1.1080 2.1280 ;
    LAYER V0 ;
      RECT 1.0760 2.3840 1.1080 2.4160 ;
    LAYER V0 ;
      RECT 1.0760 2.6720 1.1080 2.7040 ;
    LAYER V0 ;
      RECT 1.0760 3.4400 1.1080 3.4720 ;
    LAYER V0 ;
      RECT 1.0760 3.7280 1.1080 3.7600 ;
    LAYER V0 ;
      RECT 1.0760 4.0160 1.1080 4.0480 ;
    LAYER V0 ;
      RECT 1.0760 4.7840 1.1080 4.8160 ;
    LAYER V0 ;
      RECT 1.0760 5.0720 1.1080 5.1040 ;
    LAYER V0 ;
      RECT 1.0760 5.3600 1.1080 5.3920 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.7520 1.1860 0.7840 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 0.8960 1.1860 0.9280 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 1.0400 1.1860 1.0720 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.0960 1.1860 2.1280 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.2400 1.1860 2.2720 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.1540 2.3840 1.1860 2.4160 ;
    LAYER V0 ;
      RECT 1.1540 3.4400 1.1860 3.4720 ;
    LAYER V0 ;
      RECT 1.1540 3.4400 1.1860 3.4720 ;
    LAYER V0 ;
      RECT 1.1540 3.5840 1.1860 3.6160 ;
    LAYER V0 ;
      RECT 1.1540 3.5840 1.1860 3.6160 ;
    LAYER V0 ;
      RECT 1.1540 3.7280 1.1860 3.7600 ;
    LAYER V0 ;
      RECT 1.1540 3.7280 1.1860 3.7600 ;
    LAYER V0 ;
      RECT 1.1540 4.7840 1.1860 4.8160 ;
    LAYER V0 ;
      RECT 1.1540 4.7840 1.1860 4.8160 ;
    LAYER V0 ;
      RECT 1.1540 4.9280 1.1860 4.9600 ;
    LAYER V0 ;
      RECT 1.1540 4.9280 1.1860 4.9600 ;
    LAYER V0 ;
      RECT 1.1540 5.0720 1.1860 5.1040 ;
    LAYER V0 ;
      RECT 1.1540 5.0720 1.1860 5.1040 ;
    LAYER V0 ;
      RECT 1.2320 0.7520 1.2640 0.7840 ;
    LAYER V0 ;
      RECT 1.2320 0.8960 1.2640 0.9280 ;
    LAYER V0 ;
      RECT 1.2320 1.3280 1.2640 1.3600 ;
    LAYER V0 ;
      RECT 1.2320 2.0960 1.2640 2.1280 ;
    LAYER V0 ;
      RECT 1.2320 2.2400 1.2640 2.2720 ;
    LAYER V0 ;
      RECT 1.2320 2.6720 1.2640 2.7040 ;
    LAYER V0 ;
      RECT 1.2320 3.4400 1.2640 3.4720 ;
    LAYER V0 ;
      RECT 1.2320 3.5840 1.2640 3.6160 ;
    LAYER V0 ;
      RECT 1.2320 4.0160 1.2640 4.0480 ;
    LAYER V0 ;
      RECT 1.2320 4.7840 1.2640 4.8160 ;
    LAYER V0 ;
      RECT 1.2320 4.9280 1.2640 4.9600 ;
    LAYER V0 ;
      RECT 1.2320 5.3600 1.2640 5.3920 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.7520 1.3420 0.7840 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 0.8960 1.3420 0.9280 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 1.0400 1.3420 1.0720 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.0960 1.3420 2.1280 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.2400 1.3420 2.2720 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3100 2.3840 1.3420 2.4160 ;
    LAYER V0 ;
      RECT 1.3100 3.4400 1.3420 3.4720 ;
    LAYER V0 ;
      RECT 1.3100 3.4400 1.3420 3.4720 ;
    LAYER V0 ;
      RECT 1.3100 3.5840 1.3420 3.6160 ;
    LAYER V0 ;
      RECT 1.3100 3.5840 1.3420 3.6160 ;
    LAYER V0 ;
      RECT 1.3100 3.7280 1.3420 3.7600 ;
    LAYER V0 ;
      RECT 1.3100 3.7280 1.3420 3.7600 ;
    LAYER V0 ;
      RECT 1.3100 4.7840 1.3420 4.8160 ;
    LAYER V0 ;
      RECT 1.3100 4.7840 1.3420 4.8160 ;
    LAYER V0 ;
      RECT 1.3100 4.9280 1.3420 4.9600 ;
    LAYER V0 ;
      RECT 1.3100 4.9280 1.3420 4.9600 ;
    LAYER V0 ;
      RECT 1.3100 5.0720 1.3420 5.1040 ;
    LAYER V0 ;
      RECT 1.3100 5.0720 1.3420 5.1040 ;
    LAYER V0 ;
      RECT 1.3880 0.8960 1.4200 0.9280 ;
    LAYER V0 ;
      RECT 1.3880 1.0400 1.4200 1.0720 ;
    LAYER V0 ;
      RECT 1.3880 1.3280 1.4200 1.3600 ;
    LAYER V0 ;
      RECT 1.3880 2.2400 1.4200 2.2720 ;
    LAYER V0 ;
      RECT 1.3880 2.3840 1.4200 2.4160 ;
    LAYER V0 ;
      RECT 1.3880 2.6720 1.4200 2.7040 ;
    LAYER V0 ;
      RECT 1.3880 3.5840 1.4200 3.6160 ;
    LAYER V0 ;
      RECT 1.3880 3.7280 1.4200 3.7600 ;
    LAYER V0 ;
      RECT 1.3880 4.0160 1.4200 4.0480 ;
    LAYER V0 ;
      RECT 1.3880 4.9280 1.4200 4.9600 ;
    LAYER V0 ;
      RECT 1.3880 5.0720 1.4200 5.1040 ;
    LAYER V0 ;
      RECT 1.3880 5.3600 1.4200 5.3920 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.3880 6.0320 1.4200 6.0640 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
    LAYER V0 ;
      RECT 1.4660 3.4400 1.4980 3.4720 ;
    LAYER V0 ;
      RECT 1.4660 3.5840 1.4980 3.6160 ;
    LAYER V0 ;
      RECT 1.4660 3.7280 1.4980 3.7600 ;
    LAYER V0 ;
      RECT 1.4660 4.7840 1.4980 4.8160 ;
    LAYER V0 ;
      RECT 1.4660 4.9280 1.4980 4.9600 ;
    LAYER V0 ;
      RECT 1.4660 5.0720 1.4980 5.1040 ;
  END
END Switch_NMOS_n12_X4_Y4
MACRO CCP_NMOS_n12_X4_Y2
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_n12_X4_Y2 0 0 ;
  SIZE 6.2400 BY 4.0320 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3.1820 0.3420 3.2140 1.7700 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3.2600 0.4380 3.2920 1.8660 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3.3380 0.5340 3.3700 2.7300 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3.4160 0.6300 3.4480 2.8260 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6660 3.3440 5.5740 3.3760 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.9200 0.3420 0.9520 1.1940 ;
    LAYER M1 ;
      RECT 0.9200 1.3020 0.9520 1.5780 ;
    LAYER M1 ;
      RECT 0.9200 1.6860 0.9520 2.5380 ;
    LAYER M1 ;
      RECT 0.9200 2.6460 0.9520 2.9220 ;
    LAYER M1 ;
      RECT 0.9200 3.1260 0.9520 3.4980 ;
    LAYER M1 ;
      RECT 0.8420 0.3420 0.8740 1.1940 ;
    LAYER M1 ;
      RECT 0.8420 1.6860 0.8740 2.5380 ;
    LAYER M1 ;
      RECT 0.9980 0.3420 1.0300 1.1940 ;
    LAYER M1 ;
      RECT 0.9980 1.6860 1.0300 2.5380 ;
    LAYER M1 ;
      RECT 1.5440 0.3420 1.5760 1.1940 ;
    LAYER M1 ;
      RECT 1.5440 1.3020 1.5760 1.5780 ;
    LAYER M1 ;
      RECT 1.5440 1.6860 1.5760 2.5380 ;
    LAYER M1 ;
      RECT 1.5440 2.6460 1.5760 2.9220 ;
    LAYER M1 ;
      RECT 1.5440 3.1260 1.5760 3.4980 ;
    LAYER M1 ;
      RECT 1.4660 0.3420 1.4980 1.1940 ;
    LAYER M1 ;
      RECT 1.4660 1.6860 1.4980 2.5380 ;
    LAYER M1 ;
      RECT 1.6220 0.3420 1.6540 1.1940 ;
    LAYER M1 ;
      RECT 1.6220 1.6860 1.6540 2.5380 ;
    LAYER M1 ;
      RECT 2.1680 0.3420 2.2000 1.1940 ;
    LAYER M1 ;
      RECT 2.1680 1.3020 2.2000 1.5780 ;
    LAYER M1 ;
      RECT 2.1680 1.6860 2.2000 2.5380 ;
    LAYER M1 ;
      RECT 2.1680 2.6460 2.2000 2.9220 ;
    LAYER M1 ;
      RECT 2.1680 3.1260 2.2000 3.4980 ;
    LAYER M1 ;
      RECT 2.0900 0.3420 2.1220 1.1940 ;
    LAYER M1 ;
      RECT 2.0900 1.6860 2.1220 2.5380 ;
    LAYER M1 ;
      RECT 2.2460 0.3420 2.2780 1.1940 ;
    LAYER M1 ;
      RECT 2.2460 1.6860 2.2780 2.5380 ;
    LAYER M1 ;
      RECT 2.7920 0.3420 2.8240 1.1940 ;
    LAYER M1 ;
      RECT 2.7920 1.3020 2.8240 1.5780 ;
    LAYER M1 ;
      RECT 2.7920 1.6860 2.8240 2.5380 ;
    LAYER M1 ;
      RECT 2.7920 2.6460 2.8240 2.9220 ;
    LAYER M1 ;
      RECT 2.7920 3.1260 2.8240 3.4980 ;
    LAYER M1 ;
      RECT 2.7140 0.3420 2.7460 1.1940 ;
    LAYER M1 ;
      RECT 2.7140 1.6860 2.7460 2.5380 ;
    LAYER M1 ;
      RECT 2.8700 0.3420 2.9020 1.1940 ;
    LAYER M1 ;
      RECT 2.8700 1.6860 2.9020 2.5380 ;
    LAYER M1 ;
      RECT 3.4160 0.3420 3.4480 1.1940 ;
    LAYER M1 ;
      RECT 3.4160 1.3020 3.4480 1.5780 ;
    LAYER M1 ;
      RECT 3.4160 1.6860 3.4480 2.5380 ;
    LAYER M1 ;
      RECT 3.4160 2.6460 3.4480 2.9220 ;
    LAYER M1 ;
      RECT 3.4160 3.1260 3.4480 3.4980 ;
    LAYER M1 ;
      RECT 3.3380 0.3420 3.3700 1.1940 ;
    LAYER M1 ;
      RECT 3.3380 1.6860 3.3700 2.5380 ;
    LAYER M1 ;
      RECT 3.4940 0.3420 3.5260 1.1940 ;
    LAYER M1 ;
      RECT 3.4940 1.6860 3.5260 2.5380 ;
    LAYER M1 ;
      RECT 4.0400 0.3420 4.0720 1.1940 ;
    LAYER M1 ;
      RECT 4.0400 1.3020 4.0720 1.5780 ;
    LAYER M1 ;
      RECT 4.0400 1.6860 4.0720 2.5380 ;
    LAYER M1 ;
      RECT 4.0400 2.6460 4.0720 2.9220 ;
    LAYER M1 ;
      RECT 4.0400 3.1260 4.0720 3.4980 ;
    LAYER M1 ;
      RECT 3.9620 0.3420 3.9940 1.1940 ;
    LAYER M1 ;
      RECT 3.9620 1.6860 3.9940 2.5380 ;
    LAYER M1 ;
      RECT 4.1180 0.3420 4.1500 1.1940 ;
    LAYER M1 ;
      RECT 4.1180 1.6860 4.1500 2.5380 ;
    LAYER M1 ;
      RECT 4.6640 0.3420 4.6960 1.1940 ;
    LAYER M1 ;
      RECT 4.6640 1.3020 4.6960 1.5780 ;
    LAYER M1 ;
      RECT 4.6640 1.6860 4.6960 2.5380 ;
    LAYER M1 ;
      RECT 4.6640 2.6460 4.6960 2.9220 ;
    LAYER M1 ;
      RECT 4.6640 3.1260 4.6960 3.4980 ;
    LAYER M1 ;
      RECT 4.5860 0.3420 4.6180 1.1940 ;
    LAYER M1 ;
      RECT 4.5860 1.6860 4.6180 2.5380 ;
    LAYER M1 ;
      RECT 4.7420 0.3420 4.7740 1.1940 ;
    LAYER M1 ;
      RECT 4.7420 1.6860 4.7740 2.5380 ;
    LAYER M1 ;
      RECT 5.2880 0.3420 5.3200 1.1940 ;
    LAYER M1 ;
      RECT 5.2880 1.3020 5.3200 1.5780 ;
    LAYER M1 ;
      RECT 5.2880 1.6860 5.3200 2.5380 ;
    LAYER M1 ;
      RECT 5.2880 2.6460 5.3200 2.9220 ;
    LAYER M1 ;
      RECT 5.2880 3.1260 5.3200 3.4980 ;
    LAYER M1 ;
      RECT 5.2100 0.3420 5.2420 1.1940 ;
    LAYER M1 ;
      RECT 5.2100 1.6860 5.2420 2.5380 ;
    LAYER M1 ;
      RECT 5.3660 0.3420 5.3980 1.1940 ;
    LAYER M1 ;
      RECT 5.3660 1.6860 5.3980 2.5380 ;
    LAYER M2 ;
      RECT 0.7380 0.3680 5.4240 0.4000 ;
    LAYER M2 ;
      RECT 1.3620 0.4640 4.8000 0.4960 ;
    LAYER M2 ;
      RECT 0.8160 0.5600 5.3460 0.5920 ;
    LAYER M2 ;
      RECT 1.4400 1.3280 4.7220 1.3600 ;
    LAYER M2 ;
      RECT 1.4400 0.6560 4.7220 0.6880 ;
    LAYER M2 ;
      RECT 0.8160 1.4240 5.3460 1.4560 ;
    LAYER M2 ;
      RECT 1.3620 1.7120 4.8000 1.7440 ;
    LAYER M2 ;
      RECT 0.7380 1.8080 5.4240 1.8400 ;
    LAYER M2 ;
      RECT 1.4400 1.9040 4.7220 1.9360 ;
    LAYER M2 ;
      RECT 0.8160 2.6720 5.3460 2.7040 ;
    LAYER M2 ;
      RECT 0.8160 2.0000 5.3460 2.0320 ;
    LAYER M2 ;
      RECT 1.4400 2.7680 4.7220 2.8000 ;
    LAYER V1 ;
      RECT 0.9200 0.5600 0.9520 0.5920 ;
    LAYER V1 ;
      RECT 0.9200 1.4240 0.9520 1.4560 ;
    LAYER V1 ;
      RECT 0.9200 2.0000 0.9520 2.0320 ;
    LAYER V1 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V1 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V1 ;
      RECT 1.5440 0.6560 1.5760 0.6880 ;
    LAYER V1 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V1 ;
      RECT 1.5440 1.9040 1.5760 1.9360 ;
    LAYER V1 ;
      RECT 1.5440 2.7680 1.5760 2.8000 ;
    LAYER V1 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V1 ;
      RECT 2.1680 0.6560 2.2000 0.6880 ;
    LAYER V1 ;
      RECT 2.1680 1.3280 2.2000 1.3600 ;
    LAYER V1 ;
      RECT 2.1680 1.9040 2.2000 1.9360 ;
    LAYER V1 ;
      RECT 2.1680 2.7680 2.2000 2.8000 ;
    LAYER V1 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V1 ;
      RECT 2.7920 0.5600 2.8240 0.5920 ;
    LAYER V1 ;
      RECT 2.7920 1.4240 2.8240 1.4560 ;
    LAYER V1 ;
      RECT 2.7920 2.0000 2.8240 2.0320 ;
    LAYER V1 ;
      RECT 2.7920 2.6720 2.8240 2.7040 ;
    LAYER V1 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V1 ;
      RECT 3.4160 0.5600 3.4480 0.5920 ;
    LAYER V1 ;
      RECT 3.4160 1.4240 3.4480 1.4560 ;
    LAYER V1 ;
      RECT 3.4160 2.0000 3.4480 2.0320 ;
    LAYER V1 ;
      RECT 3.4160 2.6720 3.4480 2.7040 ;
    LAYER V1 ;
      RECT 3.4160 3.3440 3.4480 3.3760 ;
    LAYER V1 ;
      RECT 4.0400 0.6560 4.0720 0.6880 ;
    LAYER V1 ;
      RECT 4.0400 1.3280 4.0720 1.3600 ;
    LAYER V1 ;
      RECT 4.0400 1.9040 4.0720 1.9360 ;
    LAYER V1 ;
      RECT 4.0400 2.7680 4.0720 2.8000 ;
    LAYER V1 ;
      RECT 4.0400 3.3440 4.0720 3.3760 ;
    LAYER V1 ;
      RECT 4.6640 0.6560 4.6960 0.6880 ;
    LAYER V1 ;
      RECT 4.6640 1.3280 4.6960 1.3600 ;
    LAYER V1 ;
      RECT 4.6640 1.9040 4.6960 1.9360 ;
    LAYER V1 ;
      RECT 4.6640 2.7680 4.6960 2.8000 ;
    LAYER V1 ;
      RECT 4.6640 3.3440 4.6960 3.3760 ;
    LAYER V1 ;
      RECT 5.2880 0.5600 5.3200 0.5920 ;
    LAYER V1 ;
      RECT 5.2880 1.4240 5.3200 1.4560 ;
    LAYER V1 ;
      RECT 5.2880 2.0000 5.3200 2.0320 ;
    LAYER V1 ;
      RECT 5.2880 2.6720 5.3200 2.7040 ;
    LAYER V1 ;
      RECT 5.2880 3.3440 5.3200 3.3760 ;
    LAYER V1 ;
      RECT 3.3380 0.3680 3.3700 0.4000 ;
    LAYER V1 ;
      RECT 3.3380 1.8080 3.3700 1.8400 ;
    LAYER V1 ;
      RECT 0.8420 0.3680 0.8740 0.4000 ;
    LAYER V1 ;
      RECT 0.8420 1.8080 0.8740 1.8400 ;
    LAYER V1 ;
      RECT 3.4940 0.3680 3.5260 0.4000 ;
    LAYER V1 ;
      RECT 3.4940 1.8080 3.5260 1.8400 ;
    LAYER V1 ;
      RECT 0.9980 0.3680 1.0300 0.4000 ;
    LAYER V1 ;
      RECT 0.9980 1.8080 1.0300 1.8400 ;
    LAYER V1 ;
      RECT 2.7140 0.3680 2.7460 0.4000 ;
    LAYER V1 ;
      RECT 2.7140 1.8080 2.7460 1.8400 ;
    LAYER V1 ;
      RECT 2.8700 0.3680 2.9020 0.4000 ;
    LAYER V1 ;
      RECT 2.8700 1.8080 2.9020 1.8400 ;
    LAYER V1 ;
      RECT 5.2100 0.3680 5.2420 0.4000 ;
    LAYER V1 ;
      RECT 5.2100 1.8080 5.2420 1.8400 ;
    LAYER V1 ;
      RECT 5.3660 0.3680 5.3980 0.4000 ;
    LAYER V1 ;
      RECT 5.3660 1.8080 5.3980 1.8400 ;
    LAYER V1 ;
      RECT 1.4660 0.4640 1.4980 0.4960 ;
    LAYER V1 ;
      RECT 1.4660 1.7120 1.4980 1.7440 ;
    LAYER V1 ;
      RECT 3.9620 0.4640 3.9940 0.4960 ;
    LAYER V1 ;
      RECT 3.9620 1.7120 3.9940 1.7440 ;
    LAYER V1 ;
      RECT 1.6220 0.4640 1.6540 0.4960 ;
    LAYER V1 ;
      RECT 1.6220 1.7120 1.6540 1.7440 ;
    LAYER V1 ;
      RECT 4.1180 0.4640 4.1500 0.4960 ;
    LAYER V1 ;
      RECT 4.1180 1.7120 4.1500 1.7440 ;
    LAYER V1 ;
      RECT 4.5860 0.4640 4.6180 0.4960 ;
    LAYER V1 ;
      RECT 4.5860 1.7120 4.6180 1.7440 ;
    LAYER V1 ;
      RECT 2.0900 0.4640 2.1220 0.4960 ;
    LAYER V1 ;
      RECT 2.0900 1.7120 2.1220 1.7440 ;
    LAYER V1 ;
      RECT 4.7420 0.4640 4.7740 0.4960 ;
    LAYER V1 ;
      RECT 4.7420 1.7120 4.7740 1.7440 ;
    LAYER V1 ;
      RECT 2.2460 0.4640 2.2780 0.4960 ;
    LAYER V1 ;
      RECT 2.2460 1.7120 2.2780 1.7440 ;
    LAYER V2 ;
      RECT 3.1820 0.3680 3.2140 0.4000 ;
    LAYER V2 ;
      RECT 3.1820 1.7120 3.2140 1.7440 ;
    LAYER V2 ;
      RECT 3.2600 0.4640 3.2920 0.4960 ;
    LAYER V2 ;
      RECT 3.2600 1.8080 3.2920 1.8400 ;
    LAYER V2 ;
      RECT 3.3380 0.5600 3.3700 0.5920 ;
    LAYER V2 ;
      RECT 3.3380 1.3280 3.3700 1.3600 ;
    LAYER V2 ;
      RECT 3.3380 1.9040 3.3700 1.9360 ;
    LAYER V2 ;
      RECT 3.3380 2.6720 3.3700 2.7040 ;
    LAYER V2 ;
      RECT 3.4160 0.6560 3.4480 0.6880 ;
    LAYER V2 ;
      RECT 3.4160 1.4240 3.4480 1.4560 ;
    LAYER V2 ;
      RECT 3.4160 2.0000 3.4480 2.0320 ;
    LAYER V2 ;
      RECT 3.4160 2.7680 3.4480 2.8000 ;
    LAYER V0 ;
      RECT 0.9200 0.7520 0.9520 0.7840 ;
    LAYER V0 ;
      RECT 0.9200 0.8960 0.9520 0.9280 ;
    LAYER V0 ;
      RECT 0.9200 1.0400 0.9520 1.0720 ;
    LAYER V0 ;
      RECT 0.9200 1.3280 0.9520 1.3600 ;
    LAYER V0 ;
      RECT 0.9200 2.0960 0.9520 2.1280 ;
    LAYER V0 ;
      RECT 0.9200 2.2400 0.9520 2.2720 ;
    LAYER V0 ;
      RECT 0.9200 2.3840 0.9520 2.4160 ;
    LAYER V0 ;
      RECT 0.9200 2.6720 0.9520 2.7040 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.9200 3.3440 0.9520 3.3760 ;
    LAYER V0 ;
      RECT 0.8420 0.7520 0.8740 0.7840 ;
    LAYER V0 ;
      RECT 0.8420 0.8960 0.8740 0.9280 ;
    LAYER V0 ;
      RECT 0.8420 1.0400 0.8740 1.0720 ;
    LAYER V0 ;
      RECT 0.8420 2.0960 0.8740 2.1280 ;
    LAYER V0 ;
      RECT 0.8420 2.2400 0.8740 2.2720 ;
    LAYER V0 ;
      RECT 0.8420 2.3840 0.8740 2.4160 ;
    LAYER V0 ;
      RECT 0.9980 0.7520 1.0300 0.7840 ;
    LAYER V0 ;
      RECT 0.9980 0.8960 1.0300 0.9280 ;
    LAYER V0 ;
      RECT 0.9980 1.0400 1.0300 1.0720 ;
    LAYER V0 ;
      RECT 0.9980 2.0960 1.0300 2.1280 ;
    LAYER V0 ;
      RECT 0.9980 2.2400 1.0300 2.2720 ;
    LAYER V0 ;
      RECT 0.9980 2.3840 1.0300 2.4160 ;
    LAYER V0 ;
      RECT 1.5440 0.7520 1.5760 0.7840 ;
    LAYER V0 ;
      RECT 1.5440 0.8960 1.5760 0.9280 ;
    LAYER V0 ;
      RECT 1.5440 1.0400 1.5760 1.0720 ;
    LAYER V0 ;
      RECT 1.5440 1.3280 1.5760 1.3600 ;
    LAYER V0 ;
      RECT 1.5440 2.0960 1.5760 2.1280 ;
    LAYER V0 ;
      RECT 1.5440 2.2400 1.5760 2.2720 ;
    LAYER V0 ;
      RECT 1.5440 2.3840 1.5760 2.4160 ;
    LAYER V0 ;
      RECT 1.5440 2.6720 1.5760 2.7040 ;
    LAYER V0 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V0 ;
      RECT 1.5440 3.3440 1.5760 3.3760 ;
    LAYER V0 ;
      RECT 1.4660 0.7520 1.4980 0.7840 ;
    LAYER V0 ;
      RECT 1.4660 0.8960 1.4980 0.9280 ;
    LAYER V0 ;
      RECT 1.4660 1.0400 1.4980 1.0720 ;
    LAYER V0 ;
      RECT 1.4660 2.0960 1.4980 2.1280 ;
    LAYER V0 ;
      RECT 1.4660 2.2400 1.4980 2.2720 ;
    LAYER V0 ;
      RECT 1.4660 2.3840 1.4980 2.4160 ;
    LAYER V0 ;
      RECT 1.6220 0.7520 1.6540 0.7840 ;
    LAYER V0 ;
      RECT 1.6220 0.8960 1.6540 0.9280 ;
    LAYER V0 ;
      RECT 1.6220 1.0400 1.6540 1.0720 ;
    LAYER V0 ;
      RECT 1.6220 2.0960 1.6540 2.1280 ;
    LAYER V0 ;
      RECT 1.6220 2.2400 1.6540 2.2720 ;
    LAYER V0 ;
      RECT 1.6220 2.3840 1.6540 2.4160 ;
    LAYER V0 ;
      RECT 2.1680 0.7520 2.2000 0.7840 ;
    LAYER V0 ;
      RECT 2.1680 0.8960 2.2000 0.9280 ;
    LAYER V0 ;
      RECT 2.1680 1.0400 2.2000 1.0720 ;
    LAYER V0 ;
      RECT 2.1680 1.3280 2.2000 1.3600 ;
    LAYER V0 ;
      RECT 2.1680 2.0960 2.2000 2.1280 ;
    LAYER V0 ;
      RECT 2.1680 2.2400 2.2000 2.2720 ;
    LAYER V0 ;
      RECT 2.1680 2.3840 2.2000 2.4160 ;
    LAYER V0 ;
      RECT 2.1680 2.6720 2.2000 2.7040 ;
    LAYER V0 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V0 ;
      RECT 2.1680 3.3440 2.2000 3.3760 ;
    LAYER V0 ;
      RECT 2.0900 0.7520 2.1220 0.7840 ;
    LAYER V0 ;
      RECT 2.0900 0.8960 2.1220 0.9280 ;
    LAYER V0 ;
      RECT 2.0900 1.0400 2.1220 1.0720 ;
    LAYER V0 ;
      RECT 2.0900 2.0960 2.1220 2.1280 ;
    LAYER V0 ;
      RECT 2.0900 2.2400 2.1220 2.2720 ;
    LAYER V0 ;
      RECT 2.0900 2.3840 2.1220 2.4160 ;
    LAYER V0 ;
      RECT 2.2460 0.7520 2.2780 0.7840 ;
    LAYER V0 ;
      RECT 2.2460 0.8960 2.2780 0.9280 ;
    LAYER V0 ;
      RECT 2.2460 1.0400 2.2780 1.0720 ;
    LAYER V0 ;
      RECT 2.2460 2.0960 2.2780 2.1280 ;
    LAYER V0 ;
      RECT 2.2460 2.2400 2.2780 2.2720 ;
    LAYER V0 ;
      RECT 2.2460 2.3840 2.2780 2.4160 ;
    LAYER V0 ;
      RECT 2.7920 0.7520 2.8240 0.7840 ;
    LAYER V0 ;
      RECT 2.7920 0.8960 2.8240 0.9280 ;
    LAYER V0 ;
      RECT 2.7920 1.0400 2.8240 1.0720 ;
    LAYER V0 ;
      RECT 2.7920 1.3280 2.8240 1.3600 ;
    LAYER V0 ;
      RECT 2.7920 2.0960 2.8240 2.1280 ;
    LAYER V0 ;
      RECT 2.7920 2.2400 2.8240 2.2720 ;
    LAYER V0 ;
      RECT 2.7920 2.3840 2.8240 2.4160 ;
    LAYER V0 ;
      RECT 2.7920 2.6720 2.8240 2.7040 ;
    LAYER V0 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V0 ;
      RECT 2.7920 3.3440 2.8240 3.3760 ;
    LAYER V0 ;
      RECT 2.7140 0.7520 2.7460 0.7840 ;
    LAYER V0 ;
      RECT 2.7140 0.8960 2.7460 0.9280 ;
    LAYER V0 ;
      RECT 2.7140 1.0400 2.7460 1.0720 ;
    LAYER V0 ;
      RECT 2.7140 2.0960 2.7460 2.1280 ;
    LAYER V0 ;
      RECT 2.7140 2.2400 2.7460 2.2720 ;
    LAYER V0 ;
      RECT 2.7140 2.3840 2.7460 2.4160 ;
    LAYER V0 ;
      RECT 2.8700 0.7520 2.9020 0.7840 ;
    LAYER V0 ;
      RECT 2.8700 0.8960 2.9020 0.9280 ;
    LAYER V0 ;
      RECT 2.8700 1.0400 2.9020 1.0720 ;
    LAYER V0 ;
      RECT 2.8700 2.0960 2.9020 2.1280 ;
    LAYER V0 ;
      RECT 2.8700 2.2400 2.9020 2.2720 ;
    LAYER V0 ;
      RECT 2.8700 2.3840 2.9020 2.4160 ;
    LAYER V0 ;
      RECT 3.4160 0.7520 3.4480 0.7840 ;
    LAYER V0 ;
      RECT 3.4160 0.8960 3.4480 0.9280 ;
    LAYER V0 ;
      RECT 3.4160 1.0400 3.4480 1.0720 ;
    LAYER V0 ;
      RECT 3.4160 1.3280 3.4480 1.3600 ;
    LAYER V0 ;
      RECT 3.4160 2.0960 3.4480 2.1280 ;
    LAYER V0 ;
      RECT 3.4160 2.2400 3.4480 2.2720 ;
    LAYER V0 ;
      RECT 3.4160 2.3840 3.4480 2.4160 ;
    LAYER V0 ;
      RECT 3.4160 2.6720 3.4480 2.7040 ;
    LAYER V0 ;
      RECT 3.4160 3.3440 3.4480 3.3760 ;
    LAYER V0 ;
      RECT 3.4160 3.3440 3.4480 3.3760 ;
    LAYER V0 ;
      RECT 3.3380 0.7520 3.3700 0.7840 ;
    LAYER V0 ;
      RECT 3.3380 0.8960 3.3700 0.9280 ;
    LAYER V0 ;
      RECT 3.3380 1.0400 3.3700 1.0720 ;
    LAYER V0 ;
      RECT 3.3380 2.0960 3.3700 2.1280 ;
    LAYER V0 ;
      RECT 3.3380 2.2400 3.3700 2.2720 ;
    LAYER V0 ;
      RECT 3.3380 2.3840 3.3700 2.4160 ;
    LAYER V0 ;
      RECT 3.4940 0.7520 3.5260 0.7840 ;
    LAYER V0 ;
      RECT 3.4940 0.8960 3.5260 0.9280 ;
    LAYER V0 ;
      RECT 3.4940 1.0400 3.5260 1.0720 ;
    LAYER V0 ;
      RECT 3.4940 2.0960 3.5260 2.1280 ;
    LAYER V0 ;
      RECT 3.4940 2.2400 3.5260 2.2720 ;
    LAYER V0 ;
      RECT 3.4940 2.3840 3.5260 2.4160 ;
    LAYER V0 ;
      RECT 4.0400 0.7520 4.0720 0.7840 ;
    LAYER V0 ;
      RECT 4.0400 0.8960 4.0720 0.9280 ;
    LAYER V0 ;
      RECT 4.0400 1.0400 4.0720 1.0720 ;
    LAYER V0 ;
      RECT 4.0400 1.3280 4.0720 1.3600 ;
    LAYER V0 ;
      RECT 4.0400 2.0960 4.0720 2.1280 ;
    LAYER V0 ;
      RECT 4.0400 2.2400 4.0720 2.2720 ;
    LAYER V0 ;
      RECT 4.0400 2.3840 4.0720 2.4160 ;
    LAYER V0 ;
      RECT 4.0400 2.6720 4.0720 2.7040 ;
    LAYER V0 ;
      RECT 4.0400 3.3440 4.0720 3.3760 ;
    LAYER V0 ;
      RECT 4.0400 3.3440 4.0720 3.3760 ;
    LAYER V0 ;
      RECT 3.9620 0.7520 3.9940 0.7840 ;
    LAYER V0 ;
      RECT 3.9620 0.8960 3.9940 0.9280 ;
    LAYER V0 ;
      RECT 3.9620 1.0400 3.9940 1.0720 ;
    LAYER V0 ;
      RECT 3.9620 2.0960 3.9940 2.1280 ;
    LAYER V0 ;
      RECT 3.9620 2.2400 3.9940 2.2720 ;
    LAYER V0 ;
      RECT 3.9620 2.3840 3.9940 2.4160 ;
    LAYER V0 ;
      RECT 4.1180 0.7520 4.1500 0.7840 ;
    LAYER V0 ;
      RECT 4.1180 0.8960 4.1500 0.9280 ;
    LAYER V0 ;
      RECT 4.1180 1.0400 4.1500 1.0720 ;
    LAYER V0 ;
      RECT 4.1180 2.0960 4.1500 2.1280 ;
    LAYER V0 ;
      RECT 4.1180 2.2400 4.1500 2.2720 ;
    LAYER V0 ;
      RECT 4.1180 2.3840 4.1500 2.4160 ;
    LAYER V0 ;
      RECT 4.6640 0.7520 4.6960 0.7840 ;
    LAYER V0 ;
      RECT 4.6640 0.8960 4.6960 0.9280 ;
    LAYER V0 ;
      RECT 4.6640 1.0400 4.6960 1.0720 ;
    LAYER V0 ;
      RECT 4.6640 1.3280 4.6960 1.3600 ;
    LAYER V0 ;
      RECT 4.6640 2.0960 4.6960 2.1280 ;
    LAYER V0 ;
      RECT 4.6640 2.2400 4.6960 2.2720 ;
    LAYER V0 ;
      RECT 4.6640 2.3840 4.6960 2.4160 ;
    LAYER V0 ;
      RECT 4.6640 2.6720 4.6960 2.7040 ;
    LAYER V0 ;
      RECT 4.6640 3.3440 4.6960 3.3760 ;
    LAYER V0 ;
      RECT 4.6640 3.3440 4.6960 3.3760 ;
    LAYER V0 ;
      RECT 4.5860 0.7520 4.6180 0.7840 ;
    LAYER V0 ;
      RECT 4.5860 0.8960 4.6180 0.9280 ;
    LAYER V0 ;
      RECT 4.5860 1.0400 4.6180 1.0720 ;
    LAYER V0 ;
      RECT 4.5860 2.0960 4.6180 2.1280 ;
    LAYER V0 ;
      RECT 4.5860 2.2400 4.6180 2.2720 ;
    LAYER V0 ;
      RECT 4.5860 2.3840 4.6180 2.4160 ;
    LAYER V0 ;
      RECT 4.7420 0.7520 4.7740 0.7840 ;
    LAYER V0 ;
      RECT 4.7420 0.8960 4.7740 0.9280 ;
    LAYER V0 ;
      RECT 4.7420 1.0400 4.7740 1.0720 ;
    LAYER V0 ;
      RECT 4.7420 2.0960 4.7740 2.1280 ;
    LAYER V0 ;
      RECT 4.7420 2.2400 4.7740 2.2720 ;
    LAYER V0 ;
      RECT 4.7420 2.3840 4.7740 2.4160 ;
    LAYER V0 ;
      RECT 5.2880 0.7520 5.3200 0.7840 ;
    LAYER V0 ;
      RECT 5.2880 0.8960 5.3200 0.9280 ;
    LAYER V0 ;
      RECT 5.2880 1.0400 5.3200 1.0720 ;
    LAYER V0 ;
      RECT 5.2880 1.3280 5.3200 1.3600 ;
    LAYER V0 ;
      RECT 5.2880 2.0960 5.3200 2.1280 ;
    LAYER V0 ;
      RECT 5.2880 2.2400 5.3200 2.2720 ;
    LAYER V0 ;
      RECT 5.2880 2.3840 5.3200 2.4160 ;
    LAYER V0 ;
      RECT 5.2880 2.6720 5.3200 2.7040 ;
    LAYER V0 ;
      RECT 5.2880 3.3440 5.3200 3.3760 ;
    LAYER V0 ;
      RECT 5.2880 3.3440 5.3200 3.3760 ;
    LAYER V0 ;
      RECT 5.2100 0.7520 5.2420 0.7840 ;
    LAYER V0 ;
      RECT 5.2100 0.8960 5.2420 0.9280 ;
    LAYER V0 ;
      RECT 5.2100 1.0400 5.2420 1.0720 ;
    LAYER V0 ;
      RECT 5.2100 2.0960 5.2420 2.1280 ;
    LAYER V0 ;
      RECT 5.2100 2.2400 5.2420 2.2720 ;
    LAYER V0 ;
      RECT 5.2100 2.3840 5.2420 2.4160 ;
    LAYER V0 ;
      RECT 5.3660 0.7520 5.3980 0.7840 ;
    LAYER V0 ;
      RECT 5.3660 0.8960 5.3980 0.9280 ;
    LAYER V0 ;
      RECT 5.3660 1.0400 5.3980 1.0720 ;
    LAYER V0 ;
      RECT 5.3660 2.0960 5.3980 2.1280 ;
    LAYER V0 ;
      RECT 5.3660 2.2400 5.3980 2.2720 ;
    LAYER V0 ;
      RECT 5.3660 2.3840 5.3980 2.4160 ;
  END
END CCP_NMOS_n12_X4_Y2
