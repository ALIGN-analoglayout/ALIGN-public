MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 15.76 BY 23.1 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.844 22.644 2.876 22.716 ;
      LAYER M2 ;
        RECT 2.824 22.664 2.896 22.696 ;
      LAYER M1 ;
        RECT 12.732 22.644 12.764 22.716 ;
      LAYER M2 ;
        RECT 12.712 22.664 12.784 22.696 ;
      LAYER M2 ;
        RECT 2.86 22.664 12.748 22.696 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.98 0.384 6.012 0.456 ;
      LAYER M2 ;
        RECT 5.96 0.404 6.032 0.436 ;
      LAYER M1 ;
        RECT 9.276 0.384 9.308 0.456 ;
      LAYER M2 ;
        RECT 9.256 0.404 9.328 0.436 ;
      LAYER M2 ;
        RECT 5.996 0.404 9.292 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.3 22.812 6.332 22.884 ;
      LAYER M2 ;
        RECT 6.28 22.832 6.352 22.864 ;
      LAYER M1 ;
        RECT 9.596 22.812 9.628 22.884 ;
      LAYER M2 ;
        RECT 9.576 22.832 9.648 22.864 ;
      LAYER M2 ;
        RECT 6.316 22.832 9.612 22.864 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.684 0.216 2.716 0.288 ;
      LAYER M2 ;
        RECT 2.664 0.236 2.736 0.268 ;
      LAYER M1 ;
        RECT 12.572 0.216 12.604 0.288 ;
      LAYER M2 ;
        RECT 12.552 0.236 12.624 0.268 ;
      LAYER M2 ;
        RECT 2.7 0.236 12.588 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 9.052 7.188 9.084 7.26 ;
  LAYER M2 ;
        RECT 9.032 7.208 9.104 7.24 ;
  LAYER M2 ;
        RECT 5.996 7.208 9.068 7.24 ;
  LAYER M1 ;
        RECT 5.98 7.188 6.012 7.26 ;
  LAYER M2 ;
        RECT 5.96 7.208 6.032 7.24 ;
  LAYER M1 ;
        RECT 9.052 13.404 9.084 13.476 ;
  LAYER M2 ;
        RECT 9.032 13.424 9.104 13.456 ;
  LAYER M2 ;
        RECT 5.996 13.424 9.068 13.456 ;
  LAYER M1 ;
        RECT 5.98 13.404 6.012 13.476 ;
  LAYER M2 ;
        RECT 5.96 13.424 6.032 13.456 ;
  LAYER M1 ;
        RECT 5.756 10.296 5.788 10.368 ;
  LAYER M2 ;
        RECT 5.736 10.316 5.808 10.348 ;
  LAYER M1 ;
        RECT 5.756 10.164 5.788 10.332 ;
  LAYER M1 ;
        RECT 5.756 10.128 5.788 10.2 ;
  LAYER M2 ;
        RECT 5.736 10.148 5.808 10.18 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.996 10.18 ;
  LAYER M1 ;
        RECT 5.98 10.128 6.012 10.2 ;
  LAYER M2 ;
        RECT 5.96 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 5.756 7.188 5.788 7.26 ;
  LAYER M2 ;
        RECT 5.736 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 5.756 7.056 5.788 7.224 ;
  LAYER M1 ;
        RECT 5.756 7.02 5.788 7.092 ;
  LAYER M2 ;
        RECT 5.736 7.04 5.808 7.072 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.996 7.072 ;
  LAYER M1 ;
        RECT 5.98 7.02 6.012 7.092 ;
  LAYER M2 ;
        RECT 5.96 7.04 6.032 7.072 ;
  LAYER M1 ;
        RECT 5.98 0.384 6.012 0.456 ;
  LAYER M2 ;
        RECT 5.96 0.404 6.032 0.436 ;
  LAYER M1 ;
        RECT 5.98 0.42 6.012 0.672 ;
  LAYER M1 ;
        RECT 5.98 0.672 6.012 13.44 ;
  LAYER M1 ;
        RECT 12.348 10.296 12.38 10.368 ;
  LAYER M2 ;
        RECT 12.328 10.316 12.4 10.348 ;
  LAYER M2 ;
        RECT 9.292 10.316 12.364 10.348 ;
  LAYER M1 ;
        RECT 9.276 10.296 9.308 10.368 ;
  LAYER M2 ;
        RECT 9.256 10.316 9.328 10.348 ;
  LAYER M1 ;
        RECT 12.348 13.404 12.38 13.476 ;
  LAYER M2 ;
        RECT 12.328 13.424 12.4 13.456 ;
  LAYER M2 ;
        RECT 9.292 13.424 12.364 13.456 ;
  LAYER M1 ;
        RECT 9.276 13.404 9.308 13.476 ;
  LAYER M2 ;
        RECT 9.256 13.424 9.328 13.456 ;
  LAYER M1 ;
        RECT 9.276 0.384 9.308 0.456 ;
  LAYER M2 ;
        RECT 9.256 0.404 9.328 0.436 ;
  LAYER M1 ;
        RECT 9.276 0.42 9.308 0.672 ;
  LAYER M1 ;
        RECT 9.276 0.672 9.308 13.44 ;
  LAYER M2 ;
        RECT 5.996 0.404 9.292 0.436 ;
  LAYER M1 ;
        RECT 5.756 13.404 5.788 13.476 ;
  LAYER M2 ;
        RECT 5.736 13.424 5.808 13.456 ;
  LAYER M2 ;
        RECT 2.7 13.424 5.772 13.456 ;
  LAYER M1 ;
        RECT 2.684 13.404 2.716 13.476 ;
  LAYER M2 ;
        RECT 2.664 13.424 2.736 13.456 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 16.584 ;
  LAYER M2 ;
        RECT 5.736 16.532 5.808 16.564 ;
  LAYER M2 ;
        RECT 2.7 16.532 5.772 16.564 ;
  LAYER M1 ;
        RECT 2.684 16.512 2.716 16.584 ;
  LAYER M2 ;
        RECT 2.664 16.532 2.736 16.564 ;
  LAYER M1 ;
        RECT 2.684 0.216 2.716 0.288 ;
  LAYER M2 ;
        RECT 2.664 0.236 2.736 0.268 ;
  LAYER M1 ;
        RECT 2.684 0.252 2.716 0.672 ;
  LAYER M1 ;
        RECT 2.684 0.672 2.716 16.548 ;
  LAYER M1 ;
        RECT 12.348 7.188 12.38 7.26 ;
  LAYER M2 ;
        RECT 12.328 7.208 12.4 7.24 ;
  LAYER M1 ;
        RECT 12.348 7.056 12.38 7.224 ;
  LAYER M1 ;
        RECT 12.348 7.02 12.38 7.092 ;
  LAYER M2 ;
        RECT 12.328 7.04 12.4 7.072 ;
  LAYER M2 ;
        RECT 12.364 7.04 12.588 7.072 ;
  LAYER M1 ;
        RECT 12.572 7.02 12.604 7.092 ;
  LAYER M2 ;
        RECT 12.552 7.04 12.624 7.072 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 4.152 ;
  LAYER M2 ;
        RECT 12.328 4.1 12.4 4.132 ;
  LAYER M1 ;
        RECT 12.348 3.948 12.38 4.116 ;
  LAYER M1 ;
        RECT 12.348 3.912 12.38 3.984 ;
  LAYER M2 ;
        RECT 12.328 3.932 12.4 3.964 ;
  LAYER M2 ;
        RECT 12.364 3.932 12.588 3.964 ;
  LAYER M1 ;
        RECT 12.572 3.912 12.604 3.984 ;
  LAYER M2 ;
        RECT 12.552 3.932 12.624 3.964 ;
  LAYER M1 ;
        RECT 12.572 0.216 12.604 0.288 ;
  LAYER M2 ;
        RECT 12.552 0.236 12.624 0.268 ;
  LAYER M1 ;
        RECT 12.572 0.252 12.604 0.672 ;
  LAYER M1 ;
        RECT 12.572 0.672 12.604 7.056 ;
  LAYER M2 ;
        RECT 2.7 0.236 12.588 0.268 ;
  LAYER M1 ;
        RECT 9.052 16.512 9.084 16.584 ;
  LAYER M2 ;
        RECT 9.032 16.532 9.104 16.564 ;
  LAYER M2 ;
        RECT 5.772 16.532 9.068 16.564 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 16.584 ;
  LAYER M2 ;
        RECT 5.736 16.532 5.808 16.564 ;
  LAYER M1 ;
        RECT 9.052 4.08 9.084 4.152 ;
  LAYER M2 ;
        RECT 9.032 4.1 9.104 4.132 ;
  LAYER M2 ;
        RECT 9.068 4.1 12.364 4.132 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 4.152 ;
  LAYER M2 ;
        RECT 12.328 4.1 12.4 4.132 ;
  LAYER M1 ;
        RECT 5.756 0.972 5.788 1.044 ;
  LAYER M2 ;
        RECT 5.736 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 5.756 0.84 5.788 1.008 ;
  LAYER M1 ;
        RECT 5.756 0.804 5.788 0.876 ;
  LAYER M2 ;
        RECT 5.736 0.824 5.808 0.856 ;
  LAYER M2 ;
        RECT 5.772 0.824 6.156 0.856 ;
  LAYER M1 ;
        RECT 6.14 0.804 6.172 0.876 ;
  LAYER M2 ;
        RECT 6.12 0.824 6.192 0.856 ;
  LAYER M1 ;
        RECT 5.756 4.08 5.788 4.152 ;
  LAYER M2 ;
        RECT 5.736 4.1 5.808 4.132 ;
  LAYER M1 ;
        RECT 5.756 3.948 5.788 4.116 ;
  LAYER M1 ;
        RECT 5.756 3.912 5.788 3.984 ;
  LAYER M2 ;
        RECT 5.736 3.932 5.808 3.964 ;
  LAYER M2 ;
        RECT 5.772 3.932 6.156 3.964 ;
  LAYER M1 ;
        RECT 6.14 3.912 6.172 3.984 ;
  LAYER M2 ;
        RECT 6.12 3.932 6.192 3.964 ;
  LAYER M1 ;
        RECT 5.756 19.62 5.788 19.692 ;
  LAYER M2 ;
        RECT 5.736 19.64 5.808 19.672 ;
  LAYER M1 ;
        RECT 5.756 19.488 5.788 19.656 ;
  LAYER M1 ;
        RECT 5.756 19.452 5.788 19.524 ;
  LAYER M2 ;
        RECT 5.736 19.472 5.808 19.504 ;
  LAYER M2 ;
        RECT 5.772 19.472 6.156 19.504 ;
  LAYER M1 ;
        RECT 6.14 19.452 6.172 19.524 ;
  LAYER M2 ;
        RECT 6.12 19.472 6.192 19.504 ;
  LAYER M1 ;
        RECT 9.052 0.972 9.084 1.044 ;
  LAYER M2 ;
        RECT 9.032 0.992 9.104 1.024 ;
  LAYER M2 ;
        RECT 6.156 0.992 9.068 1.024 ;
  LAYER M1 ;
        RECT 6.14 0.972 6.172 1.044 ;
  LAYER M2 ;
        RECT 6.12 0.992 6.192 1.024 ;
  LAYER M1 ;
        RECT 9.052 10.296 9.084 10.368 ;
  LAYER M2 ;
        RECT 9.032 10.316 9.104 10.348 ;
  LAYER M2 ;
        RECT 6.156 10.316 9.068 10.348 ;
  LAYER M1 ;
        RECT 6.14 10.296 6.172 10.368 ;
  LAYER M2 ;
        RECT 6.12 10.316 6.192 10.348 ;
  LAYER M1 ;
        RECT 9.052 19.62 9.084 19.692 ;
  LAYER M2 ;
        RECT 9.032 19.64 9.104 19.672 ;
  LAYER M2 ;
        RECT 6.156 19.64 9.068 19.672 ;
  LAYER M1 ;
        RECT 6.14 19.62 6.172 19.692 ;
  LAYER M2 ;
        RECT 6.12 19.64 6.192 19.672 ;
  LAYER M1 ;
        RECT 6.14 0.048 6.172 0.12 ;
  LAYER M2 ;
        RECT 6.12 0.068 6.192 0.1 ;
  LAYER M1 ;
        RECT 6.14 0.084 6.172 0.672 ;
  LAYER M1 ;
        RECT 6.14 0.672 6.172 19.656 ;
  LAYER M1 ;
        RECT 12.348 0.972 12.38 1.044 ;
  LAYER M2 ;
        RECT 12.328 0.992 12.4 1.024 ;
  LAYER M2 ;
        RECT 9.452 0.992 12.364 1.024 ;
  LAYER M1 ;
        RECT 9.436 0.972 9.468 1.044 ;
  LAYER M2 ;
        RECT 9.416 0.992 9.488 1.024 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 16.584 ;
  LAYER M2 ;
        RECT 12.328 16.532 12.4 16.564 ;
  LAYER M2 ;
        RECT 9.452 16.532 12.364 16.564 ;
  LAYER M1 ;
        RECT 9.436 16.512 9.468 16.584 ;
  LAYER M2 ;
        RECT 9.416 16.532 9.488 16.564 ;
  LAYER M1 ;
        RECT 12.348 19.62 12.38 19.692 ;
  LAYER M2 ;
        RECT 12.328 19.64 12.4 19.672 ;
  LAYER M2 ;
        RECT 9.452 19.64 12.364 19.672 ;
  LAYER M1 ;
        RECT 9.436 19.62 9.468 19.692 ;
  LAYER M2 ;
        RECT 9.416 19.64 9.488 19.672 ;
  LAYER M1 ;
        RECT 9.436 0.048 9.468 0.12 ;
  LAYER M2 ;
        RECT 9.416 0.068 9.488 0.1 ;
  LAYER M1 ;
        RECT 9.436 0.084 9.468 0.672 ;
  LAYER M1 ;
        RECT 9.436 0.672 9.468 19.656 ;
  LAYER M2 ;
        RECT 6.156 0.068 9.452 0.1 ;
  LAYER M1 ;
        RECT 2.46 19.62 2.492 19.692 ;
  LAYER M2 ;
        RECT 2.44 19.64 2.512 19.672 ;
  LAYER M2 ;
        RECT 2.476 19.64 5.772 19.672 ;
  LAYER M1 ;
        RECT 5.756 19.62 5.788 19.692 ;
  LAYER M2 ;
        RECT 5.736 19.64 5.808 19.672 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 16.548 2.492 19.656 ;
  LAYER M1 ;
        RECT 2.46 19.62 2.492 19.692 ;
  LAYER M2 ;
        RECT 2.44 19.64 2.512 19.672 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 13.44 2.492 16.548 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 10.332 2.492 13.44 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 7.224 2.492 10.332 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 2.46 4.116 2.492 7.224 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 1.044 ;
  LAYER M2 ;
        RECT 2.44 0.992 2.512 1.024 ;
  LAYER M1 ;
        RECT 2.46 1.008 2.492 4.116 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 15.644 19.62 15.676 19.692 ;
  LAYER M2 ;
        RECT 15.624 19.64 15.696 19.672 ;
  LAYER M2 ;
        RECT 12.364 19.64 15.66 19.672 ;
  LAYER M1 ;
        RECT 12.348 19.62 12.38 19.692 ;
  LAYER M2 ;
        RECT 12.328 19.64 12.4 19.672 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 16.584 ;
  LAYER M2 ;
        RECT 15.624 16.532 15.696 16.564 ;
  LAYER M2 ;
        RECT 12.364 16.532 15.66 16.564 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 16.584 ;
  LAYER M2 ;
        RECT 12.328 16.532 12.4 16.564 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 13.476 ;
  LAYER M2 ;
        RECT 15.624 13.424 15.696 13.456 ;
  LAYER M1 ;
        RECT 15.644 13.44 15.676 16.548 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 16.584 ;
  LAYER M2 ;
        RECT 15.624 16.532 15.696 16.564 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 10.368 ;
  LAYER M2 ;
        RECT 15.624 10.316 15.696 10.348 ;
  LAYER M1 ;
        RECT 15.644 10.332 15.676 13.44 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 13.476 ;
  LAYER M2 ;
        RECT 15.624 13.424 15.696 13.456 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 7.26 ;
  LAYER M2 ;
        RECT 15.624 7.208 15.696 7.24 ;
  LAYER M1 ;
        RECT 15.644 7.224 15.676 10.332 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 10.368 ;
  LAYER M2 ;
        RECT 15.624 10.316 15.696 10.348 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 4.152 ;
  LAYER M2 ;
        RECT 15.624 4.1 15.696 4.132 ;
  LAYER M1 ;
        RECT 15.644 4.116 15.676 7.224 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 7.26 ;
  LAYER M2 ;
        RECT 15.624 7.208 15.696 7.24 ;
  LAYER M1 ;
        RECT 15.644 0.972 15.676 1.044 ;
  LAYER M2 ;
        RECT 15.624 0.992 15.696 1.024 ;
  LAYER M1 ;
        RECT 15.644 1.008 15.676 4.116 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 4.152 ;
  LAYER M2 ;
        RECT 15.624 4.1 15.696 4.132 ;
  LAYER M1 ;
        RECT 3.388 12.732 3.42 12.804 ;
  LAYER M2 ;
        RECT 3.368 12.752 3.44 12.784 ;
  LAYER M2 ;
        RECT 2.86 12.752 3.404 12.784 ;
  LAYER M1 ;
        RECT 2.844 12.732 2.876 12.804 ;
  LAYER M2 ;
        RECT 2.824 12.752 2.896 12.784 ;
  LAYER M1 ;
        RECT 3.388 9.624 3.42 9.696 ;
  LAYER M2 ;
        RECT 3.368 9.644 3.44 9.676 ;
  LAYER M2 ;
        RECT 2.86 9.644 3.404 9.676 ;
  LAYER M1 ;
        RECT 2.844 9.624 2.876 9.696 ;
  LAYER M2 ;
        RECT 2.824 9.644 2.896 9.676 ;
  LAYER M1 ;
        RECT 2.844 22.644 2.876 22.716 ;
  LAYER M2 ;
        RECT 2.824 22.664 2.896 22.696 ;
  LAYER M1 ;
        RECT 2.844 22.428 2.876 22.68 ;
  LAYER M1 ;
        RECT 2.844 9.66 2.876 22.428 ;
  LAYER M1 ;
        RECT 9.98 12.732 10.012 12.804 ;
  LAYER M2 ;
        RECT 9.96 12.752 10.032 12.784 ;
  LAYER M1 ;
        RECT 9.98 12.768 10.012 12.936 ;
  LAYER M1 ;
        RECT 9.98 12.9 10.012 12.972 ;
  LAYER M2 ;
        RECT 9.96 12.92 10.032 12.952 ;
  LAYER M2 ;
        RECT 9.996 12.92 12.748 12.952 ;
  LAYER M1 ;
        RECT 12.732 12.9 12.764 12.972 ;
  LAYER M2 ;
        RECT 12.712 12.92 12.784 12.952 ;
  LAYER M1 ;
        RECT 9.98 15.84 10.012 15.912 ;
  LAYER M2 ;
        RECT 9.96 15.86 10.032 15.892 ;
  LAYER M1 ;
        RECT 9.98 15.876 10.012 16.044 ;
  LAYER M1 ;
        RECT 9.98 16.008 10.012 16.08 ;
  LAYER M2 ;
        RECT 9.96 16.028 10.032 16.06 ;
  LAYER M2 ;
        RECT 9.996 16.028 12.748 16.06 ;
  LAYER M1 ;
        RECT 12.732 16.008 12.764 16.08 ;
  LAYER M2 ;
        RECT 12.712 16.028 12.784 16.06 ;
  LAYER M1 ;
        RECT 12.732 22.644 12.764 22.716 ;
  LAYER M2 ;
        RECT 12.712 22.664 12.784 22.696 ;
  LAYER M1 ;
        RECT 12.732 22.428 12.764 22.68 ;
  LAYER M1 ;
        RECT 12.732 12.936 12.764 22.428 ;
  LAYER M2 ;
        RECT 2.86 22.664 12.748 22.696 ;
  LAYER M1 ;
        RECT 6.684 9.624 6.716 9.696 ;
  LAYER M2 ;
        RECT 6.664 9.644 6.736 9.676 ;
  LAYER M2 ;
        RECT 3.404 9.644 6.7 9.676 ;
  LAYER M1 ;
        RECT 3.388 9.624 3.42 9.696 ;
  LAYER M2 ;
        RECT 3.368 9.644 3.44 9.676 ;
  LAYER M1 ;
        RECT 6.684 15.84 6.716 15.912 ;
  LAYER M2 ;
        RECT 6.664 15.86 6.736 15.892 ;
  LAYER M2 ;
        RECT 6.7 15.86 9.996 15.892 ;
  LAYER M1 ;
        RECT 9.98 15.84 10.012 15.912 ;
  LAYER M2 ;
        RECT 9.96 15.86 10.032 15.892 ;
  LAYER M1 ;
        RECT 3.388 15.84 3.42 15.912 ;
  LAYER M2 ;
        RECT 3.368 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 3.388 15.876 3.42 16.044 ;
  LAYER M1 ;
        RECT 3.388 16.008 3.42 16.08 ;
  LAYER M2 ;
        RECT 3.368 16.028 3.44 16.06 ;
  LAYER M2 ;
        RECT 3.404 16.028 6.316 16.06 ;
  LAYER M1 ;
        RECT 6.3 16.008 6.332 16.08 ;
  LAYER M2 ;
        RECT 6.28 16.028 6.352 16.06 ;
  LAYER M1 ;
        RECT 6.684 6.516 6.716 6.588 ;
  LAYER M2 ;
        RECT 6.664 6.536 6.736 6.568 ;
  LAYER M2 ;
        RECT 6.316 6.536 6.7 6.568 ;
  LAYER M1 ;
        RECT 6.3 6.516 6.332 6.588 ;
  LAYER M2 ;
        RECT 6.28 6.536 6.352 6.568 ;
  LAYER M1 ;
        RECT 6.684 18.948 6.716 19.02 ;
  LAYER M2 ;
        RECT 6.664 18.968 6.736 19 ;
  LAYER M2 ;
        RECT 6.316 18.968 6.7 19 ;
  LAYER M1 ;
        RECT 6.3 18.948 6.332 19.02 ;
  LAYER M2 ;
        RECT 6.28 18.968 6.352 19 ;
  LAYER M1 ;
        RECT 3.388 18.948 3.42 19.02 ;
  LAYER M2 ;
        RECT 3.368 18.968 3.44 19 ;
  LAYER M1 ;
        RECT 3.388 18.984 3.42 19.152 ;
  LAYER M1 ;
        RECT 3.388 19.116 3.42 19.188 ;
  LAYER M2 ;
        RECT 3.368 19.136 3.44 19.168 ;
  LAYER M2 ;
        RECT 3.404 19.136 6.316 19.168 ;
  LAYER M1 ;
        RECT 6.3 19.116 6.332 19.188 ;
  LAYER M2 ;
        RECT 6.28 19.136 6.352 19.168 ;
  LAYER M1 ;
        RECT 6.3 22.812 6.332 22.884 ;
  LAYER M2 ;
        RECT 6.28 22.832 6.352 22.864 ;
  LAYER M1 ;
        RECT 6.3 22.428 6.332 22.848 ;
  LAYER M1 ;
        RECT 6.3 6.552 6.332 22.428 ;
  LAYER M1 ;
        RECT 9.98 9.624 10.012 9.696 ;
  LAYER M2 ;
        RECT 9.96 9.644 10.032 9.676 ;
  LAYER M2 ;
        RECT 9.612 9.644 9.996 9.676 ;
  LAYER M1 ;
        RECT 9.596 9.624 9.628 9.696 ;
  LAYER M2 ;
        RECT 9.576 9.644 9.648 9.676 ;
  LAYER M1 ;
        RECT 9.98 6.516 10.012 6.588 ;
  LAYER M2 ;
        RECT 9.96 6.536 10.032 6.568 ;
  LAYER M2 ;
        RECT 9.612 6.536 9.996 6.568 ;
  LAYER M1 ;
        RECT 9.596 6.516 9.628 6.588 ;
  LAYER M2 ;
        RECT 9.576 6.536 9.648 6.568 ;
  LAYER M1 ;
        RECT 9.596 22.812 9.628 22.884 ;
  LAYER M2 ;
        RECT 9.576 22.832 9.648 22.864 ;
  LAYER M1 ;
        RECT 9.596 22.428 9.628 22.848 ;
  LAYER M1 ;
        RECT 9.596 6.552 9.628 22.428 ;
  LAYER M2 ;
        RECT 6.316 22.832 9.612 22.864 ;
  LAYER M1 ;
        RECT 3.388 3.408 3.42 3.48 ;
  LAYER M2 ;
        RECT 3.368 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 3.388 3.444 3.42 3.612 ;
  LAYER M1 ;
        RECT 3.388 3.576 3.42 3.648 ;
  LAYER M2 ;
        RECT 3.368 3.596 3.44 3.628 ;
  LAYER M2 ;
        RECT 3.404 3.596 6.476 3.628 ;
  LAYER M1 ;
        RECT 6.46 3.576 6.492 3.648 ;
  LAYER M2 ;
        RECT 6.44 3.596 6.512 3.628 ;
  LAYER M1 ;
        RECT 3.388 6.516 3.42 6.588 ;
  LAYER M2 ;
        RECT 3.368 6.536 3.44 6.568 ;
  LAYER M1 ;
        RECT 3.388 6.552 3.42 6.72 ;
  LAYER M1 ;
        RECT 3.388 6.684 3.42 6.756 ;
  LAYER M2 ;
        RECT 3.368 6.704 3.44 6.736 ;
  LAYER M2 ;
        RECT 3.404 6.704 6.476 6.736 ;
  LAYER M1 ;
        RECT 6.46 6.684 6.492 6.756 ;
  LAYER M2 ;
        RECT 6.44 6.704 6.512 6.736 ;
  LAYER M1 ;
        RECT 3.388 22.056 3.42 22.128 ;
  LAYER M2 ;
        RECT 3.368 22.076 3.44 22.108 ;
  LAYER M1 ;
        RECT 3.388 22.092 3.42 22.26 ;
  LAYER M1 ;
        RECT 3.388 22.224 3.42 22.296 ;
  LAYER M2 ;
        RECT 3.368 22.244 3.44 22.276 ;
  LAYER M2 ;
        RECT 3.404 22.244 6.476 22.276 ;
  LAYER M1 ;
        RECT 6.46 22.224 6.492 22.296 ;
  LAYER M2 ;
        RECT 6.44 22.244 6.512 22.276 ;
  LAYER M1 ;
        RECT 6.684 3.408 6.716 3.48 ;
  LAYER M2 ;
        RECT 6.664 3.428 6.736 3.46 ;
  LAYER M2 ;
        RECT 6.476 3.428 6.7 3.46 ;
  LAYER M1 ;
        RECT 6.46 3.408 6.492 3.48 ;
  LAYER M2 ;
        RECT 6.44 3.428 6.512 3.46 ;
  LAYER M1 ;
        RECT 6.684 12.732 6.716 12.804 ;
  LAYER M2 ;
        RECT 6.664 12.752 6.736 12.784 ;
  LAYER M2 ;
        RECT 6.476 12.752 6.7 12.784 ;
  LAYER M1 ;
        RECT 6.46 12.732 6.492 12.804 ;
  LAYER M2 ;
        RECT 6.44 12.752 6.512 12.784 ;
  LAYER M1 ;
        RECT 6.684 22.056 6.716 22.128 ;
  LAYER M2 ;
        RECT 6.664 22.076 6.736 22.108 ;
  LAYER M2 ;
        RECT 6.476 22.076 6.7 22.108 ;
  LAYER M1 ;
        RECT 6.46 22.056 6.492 22.128 ;
  LAYER M2 ;
        RECT 6.44 22.076 6.512 22.108 ;
  LAYER M1 ;
        RECT 6.46 22.98 6.492 23.052 ;
  LAYER M2 ;
        RECT 6.44 23 6.512 23.032 ;
  LAYER M1 ;
        RECT 6.46 22.428 6.492 23.016 ;
  LAYER M1 ;
        RECT 6.46 3.444 6.492 22.428 ;
  LAYER M1 ;
        RECT 9.98 3.408 10.012 3.48 ;
  LAYER M2 ;
        RECT 9.96 3.428 10.032 3.46 ;
  LAYER M2 ;
        RECT 9.772 3.428 9.996 3.46 ;
  LAYER M1 ;
        RECT 9.756 3.408 9.788 3.48 ;
  LAYER M2 ;
        RECT 9.736 3.428 9.808 3.46 ;
  LAYER M1 ;
        RECT 9.98 18.948 10.012 19.02 ;
  LAYER M2 ;
        RECT 9.96 18.968 10.032 19 ;
  LAYER M2 ;
        RECT 9.772 18.968 9.996 19 ;
  LAYER M1 ;
        RECT 9.756 18.948 9.788 19.02 ;
  LAYER M2 ;
        RECT 9.736 18.968 9.808 19 ;
  LAYER M1 ;
        RECT 9.98 22.056 10.012 22.128 ;
  LAYER M2 ;
        RECT 9.96 22.076 10.032 22.108 ;
  LAYER M2 ;
        RECT 9.772 22.076 9.996 22.108 ;
  LAYER M1 ;
        RECT 9.756 22.056 9.788 22.128 ;
  LAYER M2 ;
        RECT 9.736 22.076 9.808 22.108 ;
  LAYER M1 ;
        RECT 9.756 22.98 9.788 23.052 ;
  LAYER M2 ;
        RECT 9.736 23 9.808 23.032 ;
  LAYER M1 ;
        RECT 9.756 22.428 9.788 23.016 ;
  LAYER M1 ;
        RECT 9.756 3.444 9.788 22.428 ;
  LAYER M2 ;
        RECT 6.476 23 9.772 23.032 ;
  LAYER M1 ;
        RECT 0.092 22.056 0.124 22.128 ;
  LAYER M2 ;
        RECT 0.072 22.076 0.144 22.108 ;
  LAYER M2 ;
        RECT 0.108 22.076 3.404 22.108 ;
  LAYER M1 ;
        RECT 3.388 22.056 3.42 22.128 ;
  LAYER M2 ;
        RECT 3.368 22.076 3.44 22.108 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 18.984 0.124 22.092 ;
  LAYER M1 ;
        RECT 0.092 22.056 0.124 22.128 ;
  LAYER M2 ;
        RECT 0.072 22.076 0.144 22.108 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 15.876 0.124 18.984 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 12.768 0.124 15.876 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 9.66 0.124 12.768 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 0.092 6.552 0.124 9.66 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 3.408 0.124 3.48 ;
  LAYER M2 ;
        RECT 0.072 3.428 0.144 3.46 ;
  LAYER M1 ;
        RECT 0.092 3.444 0.124 6.552 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 13.276 22.056 13.308 22.128 ;
  LAYER M2 ;
        RECT 13.256 22.076 13.328 22.108 ;
  LAYER M2 ;
        RECT 9.996 22.076 13.292 22.108 ;
  LAYER M1 ;
        RECT 9.98 22.056 10.012 22.128 ;
  LAYER M2 ;
        RECT 9.96 22.076 10.032 22.108 ;
  LAYER M1 ;
        RECT 13.276 18.948 13.308 19.02 ;
  LAYER M2 ;
        RECT 13.256 18.968 13.328 19 ;
  LAYER M2 ;
        RECT 9.996 18.968 13.292 19 ;
  LAYER M1 ;
        RECT 9.98 18.948 10.012 19.02 ;
  LAYER M2 ;
        RECT 9.96 18.968 10.032 19 ;
  LAYER M1 ;
        RECT 13.276 15.84 13.308 15.912 ;
  LAYER M2 ;
        RECT 13.256 15.86 13.328 15.892 ;
  LAYER M1 ;
        RECT 13.276 15.876 13.308 18.984 ;
  LAYER M1 ;
        RECT 13.276 18.948 13.308 19.02 ;
  LAYER M2 ;
        RECT 13.256 18.968 13.328 19 ;
  LAYER M1 ;
        RECT 13.276 12.732 13.308 12.804 ;
  LAYER M2 ;
        RECT 13.256 12.752 13.328 12.784 ;
  LAYER M1 ;
        RECT 13.276 12.768 13.308 15.876 ;
  LAYER M1 ;
        RECT 13.276 15.84 13.308 15.912 ;
  LAYER M2 ;
        RECT 13.256 15.86 13.328 15.892 ;
  LAYER M1 ;
        RECT 13.276 9.624 13.308 9.696 ;
  LAYER M2 ;
        RECT 13.256 9.644 13.328 9.676 ;
  LAYER M1 ;
        RECT 13.276 9.66 13.308 12.768 ;
  LAYER M1 ;
        RECT 13.276 12.732 13.308 12.804 ;
  LAYER M2 ;
        RECT 13.256 12.752 13.328 12.784 ;
  LAYER M1 ;
        RECT 13.276 6.516 13.308 6.588 ;
  LAYER M2 ;
        RECT 13.256 6.536 13.328 6.568 ;
  LAYER M1 ;
        RECT 13.276 6.552 13.308 9.66 ;
  LAYER M1 ;
        RECT 13.276 9.624 13.308 9.696 ;
  LAYER M2 ;
        RECT 13.256 9.644 13.328 9.676 ;
  LAYER M1 ;
        RECT 13.276 3.408 13.308 3.48 ;
  LAYER M2 ;
        RECT 13.256 3.428 13.328 3.46 ;
  LAYER M1 ;
        RECT 13.276 3.444 13.308 6.552 ;
  LAYER M1 ;
        RECT 13.276 6.516 13.308 6.588 ;
  LAYER M2 ;
        RECT 13.256 6.536 13.328 6.568 ;
  LAYER M1 ;
        RECT 0.092 0.972 0.124 3.48 ;
  LAYER M3 ;
        RECT 0.092 3.428 0.124 3.46 ;
  LAYER M1 ;
        RECT 0.156 0.972 0.188 3.48 ;
  LAYER M3 ;
        RECT 0.156 0.992 0.188 1.024 ;
  LAYER M1 ;
        RECT 0.22 0.972 0.252 3.48 ;
  LAYER M3 ;
        RECT 0.22 3.428 0.252 3.46 ;
  LAYER M1 ;
        RECT 0.284 0.972 0.316 3.48 ;
  LAYER M3 ;
        RECT 0.284 0.992 0.316 1.024 ;
  LAYER M1 ;
        RECT 0.348 0.972 0.38 3.48 ;
  LAYER M3 ;
        RECT 0.348 3.428 0.38 3.46 ;
  LAYER M1 ;
        RECT 0.412 0.972 0.444 3.48 ;
  LAYER M3 ;
        RECT 0.412 0.992 0.444 1.024 ;
  LAYER M1 ;
        RECT 0.476 0.972 0.508 3.48 ;
  LAYER M3 ;
        RECT 0.476 3.428 0.508 3.46 ;
  LAYER M1 ;
        RECT 0.54 0.972 0.572 3.48 ;
  LAYER M3 ;
        RECT 0.54 0.992 0.572 1.024 ;
  LAYER M1 ;
        RECT 0.604 0.972 0.636 3.48 ;
  LAYER M3 ;
        RECT 0.604 3.428 0.636 3.46 ;
  LAYER M1 ;
        RECT 0.668 0.972 0.7 3.48 ;
  LAYER M3 ;
        RECT 0.668 0.992 0.7 1.024 ;
  LAYER M1 ;
        RECT 0.732 0.972 0.764 3.48 ;
  LAYER M3 ;
        RECT 0.732 3.428 0.764 3.46 ;
  LAYER M1 ;
        RECT 0.796 0.972 0.828 3.48 ;
  LAYER M3 ;
        RECT 0.796 0.992 0.828 1.024 ;
  LAYER M1 ;
        RECT 0.86 0.972 0.892 3.48 ;
  LAYER M3 ;
        RECT 0.86 3.428 0.892 3.46 ;
  LAYER M1 ;
        RECT 0.924 0.972 0.956 3.48 ;
  LAYER M3 ;
        RECT 0.924 0.992 0.956 1.024 ;
  LAYER M1 ;
        RECT 0.988 0.972 1.02 3.48 ;
  LAYER M3 ;
        RECT 0.988 3.428 1.02 3.46 ;
  LAYER M1 ;
        RECT 1.052 0.972 1.084 3.48 ;
  LAYER M3 ;
        RECT 1.052 0.992 1.084 1.024 ;
  LAYER M1 ;
        RECT 1.116 0.972 1.148 3.48 ;
  LAYER M3 ;
        RECT 1.116 3.428 1.148 3.46 ;
  LAYER M1 ;
        RECT 1.18 0.972 1.212 3.48 ;
  LAYER M3 ;
        RECT 1.18 0.992 1.212 1.024 ;
  LAYER M1 ;
        RECT 1.244 0.972 1.276 3.48 ;
  LAYER M3 ;
        RECT 1.244 3.428 1.276 3.46 ;
  LAYER M1 ;
        RECT 1.308 0.972 1.34 3.48 ;
  LAYER M3 ;
        RECT 1.308 0.992 1.34 1.024 ;
  LAYER M1 ;
        RECT 1.372 0.972 1.404 3.48 ;
  LAYER M3 ;
        RECT 1.372 3.428 1.404 3.46 ;
  LAYER M1 ;
        RECT 1.436 0.972 1.468 3.48 ;
  LAYER M3 ;
        RECT 1.436 0.992 1.468 1.024 ;
  LAYER M1 ;
        RECT 1.5 0.972 1.532 3.48 ;
  LAYER M3 ;
        RECT 1.5 3.428 1.532 3.46 ;
  LAYER M1 ;
        RECT 1.564 0.972 1.596 3.48 ;
  LAYER M3 ;
        RECT 1.564 0.992 1.596 1.024 ;
  LAYER M1 ;
        RECT 1.628 0.972 1.66 3.48 ;
  LAYER M3 ;
        RECT 1.628 3.428 1.66 3.46 ;
  LAYER M1 ;
        RECT 1.692 0.972 1.724 3.48 ;
  LAYER M3 ;
        RECT 1.692 0.992 1.724 1.024 ;
  LAYER M1 ;
        RECT 1.756 0.972 1.788 3.48 ;
  LAYER M3 ;
        RECT 1.756 3.428 1.788 3.46 ;
  LAYER M1 ;
        RECT 1.82 0.972 1.852 3.48 ;
  LAYER M3 ;
        RECT 1.82 0.992 1.852 1.024 ;
  LAYER M1 ;
        RECT 1.884 0.972 1.916 3.48 ;
  LAYER M3 ;
        RECT 1.884 3.428 1.916 3.46 ;
  LAYER M1 ;
        RECT 1.948 0.972 1.98 3.48 ;
  LAYER M3 ;
        RECT 1.948 0.992 1.98 1.024 ;
  LAYER M1 ;
        RECT 2.012 0.972 2.044 3.48 ;
  LAYER M3 ;
        RECT 2.012 3.428 2.044 3.46 ;
  LAYER M1 ;
        RECT 2.076 0.972 2.108 3.48 ;
  LAYER M3 ;
        RECT 2.076 0.992 2.108 1.024 ;
  LAYER M1 ;
        RECT 2.14 0.972 2.172 3.48 ;
  LAYER M3 ;
        RECT 2.14 3.428 2.172 3.46 ;
  LAYER M1 ;
        RECT 2.204 0.972 2.236 3.48 ;
  LAYER M3 ;
        RECT 2.204 0.992 2.236 1.024 ;
  LAYER M1 ;
        RECT 2.268 0.972 2.3 3.48 ;
  LAYER M3 ;
        RECT 2.268 3.428 2.3 3.46 ;
  LAYER M1 ;
        RECT 2.332 0.972 2.364 3.48 ;
  LAYER M3 ;
        RECT 2.332 0.992 2.364 1.024 ;
  LAYER M1 ;
        RECT 2.396 0.972 2.428 3.48 ;
  LAYER M3 ;
        RECT 2.396 3.428 2.428 3.46 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 3.48 ;
  LAYER M3 ;
        RECT 0.092 1.056 0.124 1.088 ;
  LAYER M2 ;
        RECT 2.46 1.12 2.492 1.152 ;
  LAYER M2 ;
        RECT 0.092 1.184 0.124 1.216 ;
  LAYER M2 ;
        RECT 2.46 1.248 2.492 1.28 ;
  LAYER M2 ;
        RECT 0.092 1.312 0.124 1.344 ;
  LAYER M2 ;
        RECT 2.46 1.376 2.492 1.408 ;
  LAYER M2 ;
        RECT 0.092 1.44 0.124 1.472 ;
  LAYER M2 ;
        RECT 2.46 1.504 2.492 1.536 ;
  LAYER M2 ;
        RECT 0.092 1.568 0.124 1.6 ;
  LAYER M2 ;
        RECT 2.46 1.632 2.492 1.664 ;
  LAYER M2 ;
        RECT 0.092 1.696 0.124 1.728 ;
  LAYER M2 ;
        RECT 2.46 1.76 2.492 1.792 ;
  LAYER M2 ;
        RECT 0.092 1.824 0.124 1.856 ;
  LAYER M2 ;
        RECT 2.46 1.888 2.492 1.92 ;
  LAYER M2 ;
        RECT 0.092 1.952 0.124 1.984 ;
  LAYER M2 ;
        RECT 2.46 2.016 2.492 2.048 ;
  LAYER M2 ;
        RECT 0.092 2.08 0.124 2.112 ;
  LAYER M2 ;
        RECT 2.46 2.144 2.492 2.176 ;
  LAYER M2 ;
        RECT 0.092 2.208 0.124 2.24 ;
  LAYER M2 ;
        RECT 2.46 2.272 2.492 2.304 ;
  LAYER M2 ;
        RECT 0.092 2.336 0.124 2.368 ;
  LAYER M2 ;
        RECT 2.46 2.4 2.492 2.432 ;
  LAYER M2 ;
        RECT 0.092 2.464 0.124 2.496 ;
  LAYER M2 ;
        RECT 2.46 2.528 2.492 2.56 ;
  LAYER M2 ;
        RECT 0.092 2.592 0.124 2.624 ;
  LAYER M2 ;
        RECT 2.46 2.656 2.492 2.688 ;
  LAYER M2 ;
        RECT 0.092 2.72 0.124 2.752 ;
  LAYER M2 ;
        RECT 2.46 2.784 2.492 2.816 ;
  LAYER M2 ;
        RECT 0.092 2.848 0.124 2.88 ;
  LAYER M2 ;
        RECT 2.46 2.912 2.492 2.944 ;
  LAYER M2 ;
        RECT 0.092 2.976 0.124 3.008 ;
  LAYER M2 ;
        RECT 2.46 3.04 2.492 3.072 ;
  LAYER M2 ;
        RECT 0.092 3.104 0.124 3.136 ;
  LAYER M2 ;
        RECT 2.46 3.168 2.492 3.2 ;
  LAYER M2 ;
        RECT 0.092 3.232 0.124 3.264 ;
  LAYER M2 ;
        RECT 2.46 3.296 2.492 3.328 ;
  LAYER M2 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M1 ;
        RECT 0.092 4.08 0.124 6.588 ;
  LAYER M3 ;
        RECT 0.092 6.536 0.124 6.568 ;
  LAYER M1 ;
        RECT 0.156 4.08 0.188 6.588 ;
  LAYER M3 ;
        RECT 0.156 4.1 0.188 4.132 ;
  LAYER M1 ;
        RECT 0.22 4.08 0.252 6.588 ;
  LAYER M3 ;
        RECT 0.22 6.536 0.252 6.568 ;
  LAYER M1 ;
        RECT 0.284 4.08 0.316 6.588 ;
  LAYER M3 ;
        RECT 0.284 4.1 0.316 4.132 ;
  LAYER M1 ;
        RECT 0.348 4.08 0.38 6.588 ;
  LAYER M3 ;
        RECT 0.348 6.536 0.38 6.568 ;
  LAYER M1 ;
        RECT 0.412 4.08 0.444 6.588 ;
  LAYER M3 ;
        RECT 0.412 4.1 0.444 4.132 ;
  LAYER M1 ;
        RECT 0.476 4.08 0.508 6.588 ;
  LAYER M3 ;
        RECT 0.476 6.536 0.508 6.568 ;
  LAYER M1 ;
        RECT 0.54 4.08 0.572 6.588 ;
  LAYER M3 ;
        RECT 0.54 4.1 0.572 4.132 ;
  LAYER M1 ;
        RECT 0.604 4.08 0.636 6.588 ;
  LAYER M3 ;
        RECT 0.604 6.536 0.636 6.568 ;
  LAYER M1 ;
        RECT 0.668 4.08 0.7 6.588 ;
  LAYER M3 ;
        RECT 0.668 4.1 0.7 4.132 ;
  LAYER M1 ;
        RECT 0.732 4.08 0.764 6.588 ;
  LAYER M3 ;
        RECT 0.732 6.536 0.764 6.568 ;
  LAYER M1 ;
        RECT 0.796 4.08 0.828 6.588 ;
  LAYER M3 ;
        RECT 0.796 4.1 0.828 4.132 ;
  LAYER M1 ;
        RECT 0.86 4.08 0.892 6.588 ;
  LAYER M3 ;
        RECT 0.86 6.536 0.892 6.568 ;
  LAYER M1 ;
        RECT 0.924 4.08 0.956 6.588 ;
  LAYER M3 ;
        RECT 0.924 4.1 0.956 4.132 ;
  LAYER M1 ;
        RECT 0.988 4.08 1.02 6.588 ;
  LAYER M3 ;
        RECT 0.988 6.536 1.02 6.568 ;
  LAYER M1 ;
        RECT 1.052 4.08 1.084 6.588 ;
  LAYER M3 ;
        RECT 1.052 4.1 1.084 4.132 ;
  LAYER M1 ;
        RECT 1.116 4.08 1.148 6.588 ;
  LAYER M3 ;
        RECT 1.116 6.536 1.148 6.568 ;
  LAYER M1 ;
        RECT 1.18 4.08 1.212 6.588 ;
  LAYER M3 ;
        RECT 1.18 4.1 1.212 4.132 ;
  LAYER M1 ;
        RECT 1.244 4.08 1.276 6.588 ;
  LAYER M3 ;
        RECT 1.244 6.536 1.276 6.568 ;
  LAYER M1 ;
        RECT 1.308 4.08 1.34 6.588 ;
  LAYER M3 ;
        RECT 1.308 4.1 1.34 4.132 ;
  LAYER M1 ;
        RECT 1.372 4.08 1.404 6.588 ;
  LAYER M3 ;
        RECT 1.372 6.536 1.404 6.568 ;
  LAYER M1 ;
        RECT 1.436 4.08 1.468 6.588 ;
  LAYER M3 ;
        RECT 1.436 4.1 1.468 4.132 ;
  LAYER M1 ;
        RECT 1.5 4.08 1.532 6.588 ;
  LAYER M3 ;
        RECT 1.5 6.536 1.532 6.568 ;
  LAYER M1 ;
        RECT 1.564 4.08 1.596 6.588 ;
  LAYER M3 ;
        RECT 1.564 4.1 1.596 4.132 ;
  LAYER M1 ;
        RECT 1.628 4.08 1.66 6.588 ;
  LAYER M3 ;
        RECT 1.628 6.536 1.66 6.568 ;
  LAYER M1 ;
        RECT 1.692 4.08 1.724 6.588 ;
  LAYER M3 ;
        RECT 1.692 4.1 1.724 4.132 ;
  LAYER M1 ;
        RECT 1.756 4.08 1.788 6.588 ;
  LAYER M3 ;
        RECT 1.756 6.536 1.788 6.568 ;
  LAYER M1 ;
        RECT 1.82 4.08 1.852 6.588 ;
  LAYER M3 ;
        RECT 1.82 4.1 1.852 4.132 ;
  LAYER M1 ;
        RECT 1.884 4.08 1.916 6.588 ;
  LAYER M3 ;
        RECT 1.884 6.536 1.916 6.568 ;
  LAYER M1 ;
        RECT 1.948 4.08 1.98 6.588 ;
  LAYER M3 ;
        RECT 1.948 4.1 1.98 4.132 ;
  LAYER M1 ;
        RECT 2.012 4.08 2.044 6.588 ;
  LAYER M3 ;
        RECT 2.012 6.536 2.044 6.568 ;
  LAYER M1 ;
        RECT 2.076 4.08 2.108 6.588 ;
  LAYER M3 ;
        RECT 2.076 4.1 2.108 4.132 ;
  LAYER M1 ;
        RECT 2.14 4.08 2.172 6.588 ;
  LAYER M3 ;
        RECT 2.14 6.536 2.172 6.568 ;
  LAYER M1 ;
        RECT 2.204 4.08 2.236 6.588 ;
  LAYER M3 ;
        RECT 2.204 4.1 2.236 4.132 ;
  LAYER M1 ;
        RECT 2.268 4.08 2.3 6.588 ;
  LAYER M3 ;
        RECT 2.268 6.536 2.3 6.568 ;
  LAYER M1 ;
        RECT 2.332 4.08 2.364 6.588 ;
  LAYER M3 ;
        RECT 2.332 4.1 2.364 4.132 ;
  LAYER M1 ;
        RECT 2.396 4.08 2.428 6.588 ;
  LAYER M3 ;
        RECT 2.396 6.536 2.428 6.568 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 6.588 ;
  LAYER M3 ;
        RECT 0.092 4.164 0.124 4.196 ;
  LAYER M2 ;
        RECT 2.46 4.228 2.492 4.26 ;
  LAYER M2 ;
        RECT 0.092 4.292 0.124 4.324 ;
  LAYER M2 ;
        RECT 2.46 4.356 2.492 4.388 ;
  LAYER M2 ;
        RECT 0.092 4.42 0.124 4.452 ;
  LAYER M2 ;
        RECT 2.46 4.484 2.492 4.516 ;
  LAYER M2 ;
        RECT 0.092 4.548 0.124 4.58 ;
  LAYER M2 ;
        RECT 2.46 4.612 2.492 4.644 ;
  LAYER M2 ;
        RECT 0.092 4.676 0.124 4.708 ;
  LAYER M2 ;
        RECT 2.46 4.74 2.492 4.772 ;
  LAYER M2 ;
        RECT 0.092 4.804 0.124 4.836 ;
  LAYER M2 ;
        RECT 2.46 4.868 2.492 4.9 ;
  LAYER M2 ;
        RECT 0.092 4.932 0.124 4.964 ;
  LAYER M2 ;
        RECT 2.46 4.996 2.492 5.028 ;
  LAYER M2 ;
        RECT 0.092 5.06 0.124 5.092 ;
  LAYER M2 ;
        RECT 2.46 5.124 2.492 5.156 ;
  LAYER M2 ;
        RECT 0.092 5.188 0.124 5.22 ;
  LAYER M2 ;
        RECT 2.46 5.252 2.492 5.284 ;
  LAYER M2 ;
        RECT 0.092 5.316 0.124 5.348 ;
  LAYER M2 ;
        RECT 2.46 5.38 2.492 5.412 ;
  LAYER M2 ;
        RECT 0.092 5.444 0.124 5.476 ;
  LAYER M2 ;
        RECT 2.46 5.508 2.492 5.54 ;
  LAYER M2 ;
        RECT 0.092 5.572 0.124 5.604 ;
  LAYER M2 ;
        RECT 2.46 5.636 2.492 5.668 ;
  LAYER M2 ;
        RECT 0.092 5.7 0.124 5.732 ;
  LAYER M2 ;
        RECT 2.46 5.764 2.492 5.796 ;
  LAYER M2 ;
        RECT 0.092 5.828 0.124 5.86 ;
  LAYER M2 ;
        RECT 2.46 5.892 2.492 5.924 ;
  LAYER M2 ;
        RECT 0.092 5.956 0.124 5.988 ;
  LAYER M2 ;
        RECT 2.46 6.02 2.492 6.052 ;
  LAYER M2 ;
        RECT 0.092 6.084 0.124 6.116 ;
  LAYER M2 ;
        RECT 2.46 6.148 2.492 6.18 ;
  LAYER M2 ;
        RECT 0.092 6.212 0.124 6.244 ;
  LAYER M2 ;
        RECT 2.46 6.276 2.492 6.308 ;
  LAYER M2 ;
        RECT 0.092 6.34 0.124 6.372 ;
  LAYER M2 ;
        RECT 2.46 6.404 2.492 6.436 ;
  LAYER M2 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M1 ;
        RECT 0.092 7.188 0.124 9.696 ;
  LAYER M3 ;
        RECT 0.092 9.644 0.124 9.676 ;
  LAYER M1 ;
        RECT 0.156 7.188 0.188 9.696 ;
  LAYER M3 ;
        RECT 0.156 7.208 0.188 7.24 ;
  LAYER M1 ;
        RECT 0.22 7.188 0.252 9.696 ;
  LAYER M3 ;
        RECT 0.22 9.644 0.252 9.676 ;
  LAYER M1 ;
        RECT 0.284 7.188 0.316 9.696 ;
  LAYER M3 ;
        RECT 0.284 7.208 0.316 7.24 ;
  LAYER M1 ;
        RECT 0.348 7.188 0.38 9.696 ;
  LAYER M3 ;
        RECT 0.348 9.644 0.38 9.676 ;
  LAYER M1 ;
        RECT 0.412 7.188 0.444 9.696 ;
  LAYER M3 ;
        RECT 0.412 7.208 0.444 7.24 ;
  LAYER M1 ;
        RECT 0.476 7.188 0.508 9.696 ;
  LAYER M3 ;
        RECT 0.476 9.644 0.508 9.676 ;
  LAYER M1 ;
        RECT 0.54 7.188 0.572 9.696 ;
  LAYER M3 ;
        RECT 0.54 7.208 0.572 7.24 ;
  LAYER M1 ;
        RECT 0.604 7.188 0.636 9.696 ;
  LAYER M3 ;
        RECT 0.604 9.644 0.636 9.676 ;
  LAYER M1 ;
        RECT 0.668 7.188 0.7 9.696 ;
  LAYER M3 ;
        RECT 0.668 7.208 0.7 7.24 ;
  LAYER M1 ;
        RECT 0.732 7.188 0.764 9.696 ;
  LAYER M3 ;
        RECT 0.732 9.644 0.764 9.676 ;
  LAYER M1 ;
        RECT 0.796 7.188 0.828 9.696 ;
  LAYER M3 ;
        RECT 0.796 7.208 0.828 7.24 ;
  LAYER M1 ;
        RECT 0.86 7.188 0.892 9.696 ;
  LAYER M3 ;
        RECT 0.86 9.644 0.892 9.676 ;
  LAYER M1 ;
        RECT 0.924 7.188 0.956 9.696 ;
  LAYER M3 ;
        RECT 0.924 7.208 0.956 7.24 ;
  LAYER M1 ;
        RECT 0.988 7.188 1.02 9.696 ;
  LAYER M3 ;
        RECT 0.988 9.644 1.02 9.676 ;
  LAYER M1 ;
        RECT 1.052 7.188 1.084 9.696 ;
  LAYER M3 ;
        RECT 1.052 7.208 1.084 7.24 ;
  LAYER M1 ;
        RECT 1.116 7.188 1.148 9.696 ;
  LAYER M3 ;
        RECT 1.116 9.644 1.148 9.676 ;
  LAYER M1 ;
        RECT 1.18 7.188 1.212 9.696 ;
  LAYER M3 ;
        RECT 1.18 7.208 1.212 7.24 ;
  LAYER M1 ;
        RECT 1.244 7.188 1.276 9.696 ;
  LAYER M3 ;
        RECT 1.244 9.644 1.276 9.676 ;
  LAYER M1 ;
        RECT 1.308 7.188 1.34 9.696 ;
  LAYER M3 ;
        RECT 1.308 7.208 1.34 7.24 ;
  LAYER M1 ;
        RECT 1.372 7.188 1.404 9.696 ;
  LAYER M3 ;
        RECT 1.372 9.644 1.404 9.676 ;
  LAYER M1 ;
        RECT 1.436 7.188 1.468 9.696 ;
  LAYER M3 ;
        RECT 1.436 7.208 1.468 7.24 ;
  LAYER M1 ;
        RECT 1.5 7.188 1.532 9.696 ;
  LAYER M3 ;
        RECT 1.5 9.644 1.532 9.676 ;
  LAYER M1 ;
        RECT 1.564 7.188 1.596 9.696 ;
  LAYER M3 ;
        RECT 1.564 7.208 1.596 7.24 ;
  LAYER M1 ;
        RECT 1.628 7.188 1.66 9.696 ;
  LAYER M3 ;
        RECT 1.628 9.644 1.66 9.676 ;
  LAYER M1 ;
        RECT 1.692 7.188 1.724 9.696 ;
  LAYER M3 ;
        RECT 1.692 7.208 1.724 7.24 ;
  LAYER M1 ;
        RECT 1.756 7.188 1.788 9.696 ;
  LAYER M3 ;
        RECT 1.756 9.644 1.788 9.676 ;
  LAYER M1 ;
        RECT 1.82 7.188 1.852 9.696 ;
  LAYER M3 ;
        RECT 1.82 7.208 1.852 7.24 ;
  LAYER M1 ;
        RECT 1.884 7.188 1.916 9.696 ;
  LAYER M3 ;
        RECT 1.884 9.644 1.916 9.676 ;
  LAYER M1 ;
        RECT 1.948 7.188 1.98 9.696 ;
  LAYER M3 ;
        RECT 1.948 7.208 1.98 7.24 ;
  LAYER M1 ;
        RECT 2.012 7.188 2.044 9.696 ;
  LAYER M3 ;
        RECT 2.012 9.644 2.044 9.676 ;
  LAYER M1 ;
        RECT 2.076 7.188 2.108 9.696 ;
  LAYER M3 ;
        RECT 2.076 7.208 2.108 7.24 ;
  LAYER M1 ;
        RECT 2.14 7.188 2.172 9.696 ;
  LAYER M3 ;
        RECT 2.14 9.644 2.172 9.676 ;
  LAYER M1 ;
        RECT 2.204 7.188 2.236 9.696 ;
  LAYER M3 ;
        RECT 2.204 7.208 2.236 7.24 ;
  LAYER M1 ;
        RECT 2.268 7.188 2.3 9.696 ;
  LAYER M3 ;
        RECT 2.268 9.644 2.3 9.676 ;
  LAYER M1 ;
        RECT 2.332 7.188 2.364 9.696 ;
  LAYER M3 ;
        RECT 2.332 7.208 2.364 7.24 ;
  LAYER M1 ;
        RECT 2.396 7.188 2.428 9.696 ;
  LAYER M3 ;
        RECT 2.396 9.644 2.428 9.676 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 9.696 ;
  LAYER M3 ;
        RECT 0.092 7.272 0.124 7.304 ;
  LAYER M2 ;
        RECT 2.46 7.336 2.492 7.368 ;
  LAYER M2 ;
        RECT 0.092 7.4 0.124 7.432 ;
  LAYER M2 ;
        RECT 2.46 7.464 2.492 7.496 ;
  LAYER M2 ;
        RECT 0.092 7.528 0.124 7.56 ;
  LAYER M2 ;
        RECT 2.46 7.592 2.492 7.624 ;
  LAYER M2 ;
        RECT 0.092 7.656 0.124 7.688 ;
  LAYER M2 ;
        RECT 2.46 7.72 2.492 7.752 ;
  LAYER M2 ;
        RECT 0.092 7.784 0.124 7.816 ;
  LAYER M2 ;
        RECT 2.46 7.848 2.492 7.88 ;
  LAYER M2 ;
        RECT 0.092 7.912 0.124 7.944 ;
  LAYER M2 ;
        RECT 2.46 7.976 2.492 8.008 ;
  LAYER M2 ;
        RECT 0.092 8.04 0.124 8.072 ;
  LAYER M2 ;
        RECT 2.46 8.104 2.492 8.136 ;
  LAYER M2 ;
        RECT 0.092 8.168 0.124 8.2 ;
  LAYER M2 ;
        RECT 2.46 8.232 2.492 8.264 ;
  LAYER M2 ;
        RECT 0.092 8.296 0.124 8.328 ;
  LAYER M2 ;
        RECT 2.46 8.36 2.492 8.392 ;
  LAYER M2 ;
        RECT 0.092 8.424 0.124 8.456 ;
  LAYER M2 ;
        RECT 2.46 8.488 2.492 8.52 ;
  LAYER M2 ;
        RECT 0.092 8.552 0.124 8.584 ;
  LAYER M2 ;
        RECT 2.46 8.616 2.492 8.648 ;
  LAYER M2 ;
        RECT 0.092 8.68 0.124 8.712 ;
  LAYER M2 ;
        RECT 2.46 8.744 2.492 8.776 ;
  LAYER M2 ;
        RECT 0.092 8.808 0.124 8.84 ;
  LAYER M2 ;
        RECT 2.46 8.872 2.492 8.904 ;
  LAYER M2 ;
        RECT 0.092 8.936 0.124 8.968 ;
  LAYER M2 ;
        RECT 2.46 9 2.492 9.032 ;
  LAYER M2 ;
        RECT 0.092 9.064 0.124 9.096 ;
  LAYER M2 ;
        RECT 2.46 9.128 2.492 9.16 ;
  LAYER M2 ;
        RECT 0.092 9.192 0.124 9.224 ;
  LAYER M2 ;
        RECT 2.46 9.256 2.492 9.288 ;
  LAYER M2 ;
        RECT 0.092 9.32 0.124 9.352 ;
  LAYER M2 ;
        RECT 2.46 9.384 2.492 9.416 ;
  LAYER M2 ;
        RECT 0.092 9.448 0.124 9.48 ;
  LAYER M2 ;
        RECT 2.46 9.512 2.492 9.544 ;
  LAYER M2 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M1 ;
        RECT 0.092 10.296 0.124 12.804 ;
  LAYER M3 ;
        RECT 0.092 12.752 0.124 12.784 ;
  LAYER M1 ;
        RECT 0.156 10.296 0.188 12.804 ;
  LAYER M3 ;
        RECT 0.156 10.316 0.188 10.348 ;
  LAYER M1 ;
        RECT 0.22 10.296 0.252 12.804 ;
  LAYER M3 ;
        RECT 0.22 12.752 0.252 12.784 ;
  LAYER M1 ;
        RECT 0.284 10.296 0.316 12.804 ;
  LAYER M3 ;
        RECT 0.284 10.316 0.316 10.348 ;
  LAYER M1 ;
        RECT 0.348 10.296 0.38 12.804 ;
  LAYER M3 ;
        RECT 0.348 12.752 0.38 12.784 ;
  LAYER M1 ;
        RECT 0.412 10.296 0.444 12.804 ;
  LAYER M3 ;
        RECT 0.412 10.316 0.444 10.348 ;
  LAYER M1 ;
        RECT 0.476 10.296 0.508 12.804 ;
  LAYER M3 ;
        RECT 0.476 12.752 0.508 12.784 ;
  LAYER M1 ;
        RECT 0.54 10.296 0.572 12.804 ;
  LAYER M3 ;
        RECT 0.54 10.316 0.572 10.348 ;
  LAYER M1 ;
        RECT 0.604 10.296 0.636 12.804 ;
  LAYER M3 ;
        RECT 0.604 12.752 0.636 12.784 ;
  LAYER M1 ;
        RECT 0.668 10.296 0.7 12.804 ;
  LAYER M3 ;
        RECT 0.668 10.316 0.7 10.348 ;
  LAYER M1 ;
        RECT 0.732 10.296 0.764 12.804 ;
  LAYER M3 ;
        RECT 0.732 12.752 0.764 12.784 ;
  LAYER M1 ;
        RECT 0.796 10.296 0.828 12.804 ;
  LAYER M3 ;
        RECT 0.796 10.316 0.828 10.348 ;
  LAYER M1 ;
        RECT 0.86 10.296 0.892 12.804 ;
  LAYER M3 ;
        RECT 0.86 12.752 0.892 12.784 ;
  LAYER M1 ;
        RECT 0.924 10.296 0.956 12.804 ;
  LAYER M3 ;
        RECT 0.924 10.316 0.956 10.348 ;
  LAYER M1 ;
        RECT 0.988 10.296 1.02 12.804 ;
  LAYER M3 ;
        RECT 0.988 12.752 1.02 12.784 ;
  LAYER M1 ;
        RECT 1.052 10.296 1.084 12.804 ;
  LAYER M3 ;
        RECT 1.052 10.316 1.084 10.348 ;
  LAYER M1 ;
        RECT 1.116 10.296 1.148 12.804 ;
  LAYER M3 ;
        RECT 1.116 12.752 1.148 12.784 ;
  LAYER M1 ;
        RECT 1.18 10.296 1.212 12.804 ;
  LAYER M3 ;
        RECT 1.18 10.316 1.212 10.348 ;
  LAYER M1 ;
        RECT 1.244 10.296 1.276 12.804 ;
  LAYER M3 ;
        RECT 1.244 12.752 1.276 12.784 ;
  LAYER M1 ;
        RECT 1.308 10.296 1.34 12.804 ;
  LAYER M3 ;
        RECT 1.308 10.316 1.34 10.348 ;
  LAYER M1 ;
        RECT 1.372 10.296 1.404 12.804 ;
  LAYER M3 ;
        RECT 1.372 12.752 1.404 12.784 ;
  LAYER M1 ;
        RECT 1.436 10.296 1.468 12.804 ;
  LAYER M3 ;
        RECT 1.436 10.316 1.468 10.348 ;
  LAYER M1 ;
        RECT 1.5 10.296 1.532 12.804 ;
  LAYER M3 ;
        RECT 1.5 12.752 1.532 12.784 ;
  LAYER M1 ;
        RECT 1.564 10.296 1.596 12.804 ;
  LAYER M3 ;
        RECT 1.564 10.316 1.596 10.348 ;
  LAYER M1 ;
        RECT 1.628 10.296 1.66 12.804 ;
  LAYER M3 ;
        RECT 1.628 12.752 1.66 12.784 ;
  LAYER M1 ;
        RECT 1.692 10.296 1.724 12.804 ;
  LAYER M3 ;
        RECT 1.692 10.316 1.724 10.348 ;
  LAYER M1 ;
        RECT 1.756 10.296 1.788 12.804 ;
  LAYER M3 ;
        RECT 1.756 12.752 1.788 12.784 ;
  LAYER M1 ;
        RECT 1.82 10.296 1.852 12.804 ;
  LAYER M3 ;
        RECT 1.82 10.316 1.852 10.348 ;
  LAYER M1 ;
        RECT 1.884 10.296 1.916 12.804 ;
  LAYER M3 ;
        RECT 1.884 12.752 1.916 12.784 ;
  LAYER M1 ;
        RECT 1.948 10.296 1.98 12.804 ;
  LAYER M3 ;
        RECT 1.948 10.316 1.98 10.348 ;
  LAYER M1 ;
        RECT 2.012 10.296 2.044 12.804 ;
  LAYER M3 ;
        RECT 2.012 12.752 2.044 12.784 ;
  LAYER M1 ;
        RECT 2.076 10.296 2.108 12.804 ;
  LAYER M3 ;
        RECT 2.076 10.316 2.108 10.348 ;
  LAYER M1 ;
        RECT 2.14 10.296 2.172 12.804 ;
  LAYER M3 ;
        RECT 2.14 12.752 2.172 12.784 ;
  LAYER M1 ;
        RECT 2.204 10.296 2.236 12.804 ;
  LAYER M3 ;
        RECT 2.204 10.316 2.236 10.348 ;
  LAYER M1 ;
        RECT 2.268 10.296 2.3 12.804 ;
  LAYER M3 ;
        RECT 2.268 12.752 2.3 12.784 ;
  LAYER M1 ;
        RECT 2.332 10.296 2.364 12.804 ;
  LAYER M3 ;
        RECT 2.332 10.316 2.364 10.348 ;
  LAYER M1 ;
        RECT 2.396 10.296 2.428 12.804 ;
  LAYER M3 ;
        RECT 2.396 12.752 2.428 12.784 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 12.804 ;
  LAYER M3 ;
        RECT 0.092 10.38 0.124 10.412 ;
  LAYER M2 ;
        RECT 2.46 10.444 2.492 10.476 ;
  LAYER M2 ;
        RECT 0.092 10.508 0.124 10.54 ;
  LAYER M2 ;
        RECT 2.46 10.572 2.492 10.604 ;
  LAYER M2 ;
        RECT 0.092 10.636 0.124 10.668 ;
  LAYER M2 ;
        RECT 2.46 10.7 2.492 10.732 ;
  LAYER M2 ;
        RECT 0.092 10.764 0.124 10.796 ;
  LAYER M2 ;
        RECT 2.46 10.828 2.492 10.86 ;
  LAYER M2 ;
        RECT 0.092 10.892 0.124 10.924 ;
  LAYER M2 ;
        RECT 2.46 10.956 2.492 10.988 ;
  LAYER M2 ;
        RECT 0.092 11.02 0.124 11.052 ;
  LAYER M2 ;
        RECT 2.46 11.084 2.492 11.116 ;
  LAYER M2 ;
        RECT 0.092 11.148 0.124 11.18 ;
  LAYER M2 ;
        RECT 2.46 11.212 2.492 11.244 ;
  LAYER M2 ;
        RECT 0.092 11.276 0.124 11.308 ;
  LAYER M2 ;
        RECT 2.46 11.34 2.492 11.372 ;
  LAYER M2 ;
        RECT 0.092 11.404 0.124 11.436 ;
  LAYER M2 ;
        RECT 2.46 11.468 2.492 11.5 ;
  LAYER M2 ;
        RECT 0.092 11.532 0.124 11.564 ;
  LAYER M2 ;
        RECT 2.46 11.596 2.492 11.628 ;
  LAYER M2 ;
        RECT 0.092 11.66 0.124 11.692 ;
  LAYER M2 ;
        RECT 2.46 11.724 2.492 11.756 ;
  LAYER M2 ;
        RECT 0.092 11.788 0.124 11.82 ;
  LAYER M2 ;
        RECT 2.46 11.852 2.492 11.884 ;
  LAYER M2 ;
        RECT 0.092 11.916 0.124 11.948 ;
  LAYER M2 ;
        RECT 2.46 11.98 2.492 12.012 ;
  LAYER M2 ;
        RECT 0.092 12.044 0.124 12.076 ;
  LAYER M2 ;
        RECT 2.46 12.108 2.492 12.14 ;
  LAYER M2 ;
        RECT 0.092 12.172 0.124 12.204 ;
  LAYER M2 ;
        RECT 2.46 12.236 2.492 12.268 ;
  LAYER M2 ;
        RECT 0.092 12.3 0.124 12.332 ;
  LAYER M2 ;
        RECT 2.46 12.364 2.492 12.396 ;
  LAYER M2 ;
        RECT 0.092 12.428 0.124 12.46 ;
  LAYER M2 ;
        RECT 2.46 12.492 2.492 12.524 ;
  LAYER M2 ;
        RECT 0.092 12.556 0.124 12.588 ;
  LAYER M2 ;
        RECT 2.46 12.62 2.492 12.652 ;
  LAYER M2 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M1 ;
        RECT 0.092 13.404 0.124 15.912 ;
  LAYER M3 ;
        RECT 0.092 15.86 0.124 15.892 ;
  LAYER M1 ;
        RECT 0.156 13.404 0.188 15.912 ;
  LAYER M3 ;
        RECT 0.156 13.424 0.188 13.456 ;
  LAYER M1 ;
        RECT 0.22 13.404 0.252 15.912 ;
  LAYER M3 ;
        RECT 0.22 15.86 0.252 15.892 ;
  LAYER M1 ;
        RECT 0.284 13.404 0.316 15.912 ;
  LAYER M3 ;
        RECT 0.284 13.424 0.316 13.456 ;
  LAYER M1 ;
        RECT 0.348 13.404 0.38 15.912 ;
  LAYER M3 ;
        RECT 0.348 15.86 0.38 15.892 ;
  LAYER M1 ;
        RECT 0.412 13.404 0.444 15.912 ;
  LAYER M3 ;
        RECT 0.412 13.424 0.444 13.456 ;
  LAYER M1 ;
        RECT 0.476 13.404 0.508 15.912 ;
  LAYER M3 ;
        RECT 0.476 15.86 0.508 15.892 ;
  LAYER M1 ;
        RECT 0.54 13.404 0.572 15.912 ;
  LAYER M3 ;
        RECT 0.54 13.424 0.572 13.456 ;
  LAYER M1 ;
        RECT 0.604 13.404 0.636 15.912 ;
  LAYER M3 ;
        RECT 0.604 15.86 0.636 15.892 ;
  LAYER M1 ;
        RECT 0.668 13.404 0.7 15.912 ;
  LAYER M3 ;
        RECT 0.668 13.424 0.7 13.456 ;
  LAYER M1 ;
        RECT 0.732 13.404 0.764 15.912 ;
  LAYER M3 ;
        RECT 0.732 15.86 0.764 15.892 ;
  LAYER M1 ;
        RECT 0.796 13.404 0.828 15.912 ;
  LAYER M3 ;
        RECT 0.796 13.424 0.828 13.456 ;
  LAYER M1 ;
        RECT 0.86 13.404 0.892 15.912 ;
  LAYER M3 ;
        RECT 0.86 15.86 0.892 15.892 ;
  LAYER M1 ;
        RECT 0.924 13.404 0.956 15.912 ;
  LAYER M3 ;
        RECT 0.924 13.424 0.956 13.456 ;
  LAYER M1 ;
        RECT 0.988 13.404 1.02 15.912 ;
  LAYER M3 ;
        RECT 0.988 15.86 1.02 15.892 ;
  LAYER M1 ;
        RECT 1.052 13.404 1.084 15.912 ;
  LAYER M3 ;
        RECT 1.052 13.424 1.084 13.456 ;
  LAYER M1 ;
        RECT 1.116 13.404 1.148 15.912 ;
  LAYER M3 ;
        RECT 1.116 15.86 1.148 15.892 ;
  LAYER M1 ;
        RECT 1.18 13.404 1.212 15.912 ;
  LAYER M3 ;
        RECT 1.18 13.424 1.212 13.456 ;
  LAYER M1 ;
        RECT 1.244 13.404 1.276 15.912 ;
  LAYER M3 ;
        RECT 1.244 15.86 1.276 15.892 ;
  LAYER M1 ;
        RECT 1.308 13.404 1.34 15.912 ;
  LAYER M3 ;
        RECT 1.308 13.424 1.34 13.456 ;
  LAYER M1 ;
        RECT 1.372 13.404 1.404 15.912 ;
  LAYER M3 ;
        RECT 1.372 15.86 1.404 15.892 ;
  LAYER M1 ;
        RECT 1.436 13.404 1.468 15.912 ;
  LAYER M3 ;
        RECT 1.436 13.424 1.468 13.456 ;
  LAYER M1 ;
        RECT 1.5 13.404 1.532 15.912 ;
  LAYER M3 ;
        RECT 1.5 15.86 1.532 15.892 ;
  LAYER M1 ;
        RECT 1.564 13.404 1.596 15.912 ;
  LAYER M3 ;
        RECT 1.564 13.424 1.596 13.456 ;
  LAYER M1 ;
        RECT 1.628 13.404 1.66 15.912 ;
  LAYER M3 ;
        RECT 1.628 15.86 1.66 15.892 ;
  LAYER M1 ;
        RECT 1.692 13.404 1.724 15.912 ;
  LAYER M3 ;
        RECT 1.692 13.424 1.724 13.456 ;
  LAYER M1 ;
        RECT 1.756 13.404 1.788 15.912 ;
  LAYER M3 ;
        RECT 1.756 15.86 1.788 15.892 ;
  LAYER M1 ;
        RECT 1.82 13.404 1.852 15.912 ;
  LAYER M3 ;
        RECT 1.82 13.424 1.852 13.456 ;
  LAYER M1 ;
        RECT 1.884 13.404 1.916 15.912 ;
  LAYER M3 ;
        RECT 1.884 15.86 1.916 15.892 ;
  LAYER M1 ;
        RECT 1.948 13.404 1.98 15.912 ;
  LAYER M3 ;
        RECT 1.948 13.424 1.98 13.456 ;
  LAYER M1 ;
        RECT 2.012 13.404 2.044 15.912 ;
  LAYER M3 ;
        RECT 2.012 15.86 2.044 15.892 ;
  LAYER M1 ;
        RECT 2.076 13.404 2.108 15.912 ;
  LAYER M3 ;
        RECT 2.076 13.424 2.108 13.456 ;
  LAYER M1 ;
        RECT 2.14 13.404 2.172 15.912 ;
  LAYER M3 ;
        RECT 2.14 15.86 2.172 15.892 ;
  LAYER M1 ;
        RECT 2.204 13.404 2.236 15.912 ;
  LAYER M3 ;
        RECT 2.204 13.424 2.236 13.456 ;
  LAYER M1 ;
        RECT 2.268 13.404 2.3 15.912 ;
  LAYER M3 ;
        RECT 2.268 15.86 2.3 15.892 ;
  LAYER M1 ;
        RECT 2.332 13.404 2.364 15.912 ;
  LAYER M3 ;
        RECT 2.332 13.424 2.364 13.456 ;
  LAYER M1 ;
        RECT 2.396 13.404 2.428 15.912 ;
  LAYER M3 ;
        RECT 2.396 15.86 2.428 15.892 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 15.912 ;
  LAYER M3 ;
        RECT 0.092 13.488 0.124 13.52 ;
  LAYER M2 ;
        RECT 2.46 13.552 2.492 13.584 ;
  LAYER M2 ;
        RECT 0.092 13.616 0.124 13.648 ;
  LAYER M2 ;
        RECT 2.46 13.68 2.492 13.712 ;
  LAYER M2 ;
        RECT 0.092 13.744 0.124 13.776 ;
  LAYER M2 ;
        RECT 2.46 13.808 2.492 13.84 ;
  LAYER M2 ;
        RECT 0.092 13.872 0.124 13.904 ;
  LAYER M2 ;
        RECT 2.46 13.936 2.492 13.968 ;
  LAYER M2 ;
        RECT 0.092 14 0.124 14.032 ;
  LAYER M2 ;
        RECT 2.46 14.064 2.492 14.096 ;
  LAYER M2 ;
        RECT 0.092 14.128 0.124 14.16 ;
  LAYER M2 ;
        RECT 2.46 14.192 2.492 14.224 ;
  LAYER M2 ;
        RECT 0.092 14.256 0.124 14.288 ;
  LAYER M2 ;
        RECT 2.46 14.32 2.492 14.352 ;
  LAYER M2 ;
        RECT 0.092 14.384 0.124 14.416 ;
  LAYER M2 ;
        RECT 2.46 14.448 2.492 14.48 ;
  LAYER M2 ;
        RECT 0.092 14.512 0.124 14.544 ;
  LAYER M2 ;
        RECT 2.46 14.576 2.492 14.608 ;
  LAYER M2 ;
        RECT 0.092 14.64 0.124 14.672 ;
  LAYER M2 ;
        RECT 2.46 14.704 2.492 14.736 ;
  LAYER M2 ;
        RECT 0.092 14.768 0.124 14.8 ;
  LAYER M2 ;
        RECT 2.46 14.832 2.492 14.864 ;
  LAYER M2 ;
        RECT 0.092 14.896 0.124 14.928 ;
  LAYER M2 ;
        RECT 2.46 14.96 2.492 14.992 ;
  LAYER M2 ;
        RECT 0.092 15.024 0.124 15.056 ;
  LAYER M2 ;
        RECT 2.46 15.088 2.492 15.12 ;
  LAYER M2 ;
        RECT 0.092 15.152 0.124 15.184 ;
  LAYER M2 ;
        RECT 2.46 15.216 2.492 15.248 ;
  LAYER M2 ;
        RECT 0.092 15.28 0.124 15.312 ;
  LAYER M2 ;
        RECT 2.46 15.344 2.492 15.376 ;
  LAYER M2 ;
        RECT 0.092 15.408 0.124 15.44 ;
  LAYER M2 ;
        RECT 2.46 15.472 2.492 15.504 ;
  LAYER M2 ;
        RECT 0.092 15.536 0.124 15.568 ;
  LAYER M2 ;
        RECT 2.46 15.6 2.492 15.632 ;
  LAYER M2 ;
        RECT 0.092 15.664 0.124 15.696 ;
  LAYER M2 ;
        RECT 2.46 15.728 2.492 15.76 ;
  LAYER M2 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M1 ;
        RECT 0.092 16.512 0.124 19.02 ;
  LAYER M3 ;
        RECT 0.092 18.968 0.124 19 ;
  LAYER M1 ;
        RECT 0.156 16.512 0.188 19.02 ;
  LAYER M3 ;
        RECT 0.156 16.532 0.188 16.564 ;
  LAYER M1 ;
        RECT 0.22 16.512 0.252 19.02 ;
  LAYER M3 ;
        RECT 0.22 18.968 0.252 19 ;
  LAYER M1 ;
        RECT 0.284 16.512 0.316 19.02 ;
  LAYER M3 ;
        RECT 0.284 16.532 0.316 16.564 ;
  LAYER M1 ;
        RECT 0.348 16.512 0.38 19.02 ;
  LAYER M3 ;
        RECT 0.348 18.968 0.38 19 ;
  LAYER M1 ;
        RECT 0.412 16.512 0.444 19.02 ;
  LAYER M3 ;
        RECT 0.412 16.532 0.444 16.564 ;
  LAYER M1 ;
        RECT 0.476 16.512 0.508 19.02 ;
  LAYER M3 ;
        RECT 0.476 18.968 0.508 19 ;
  LAYER M1 ;
        RECT 0.54 16.512 0.572 19.02 ;
  LAYER M3 ;
        RECT 0.54 16.532 0.572 16.564 ;
  LAYER M1 ;
        RECT 0.604 16.512 0.636 19.02 ;
  LAYER M3 ;
        RECT 0.604 18.968 0.636 19 ;
  LAYER M1 ;
        RECT 0.668 16.512 0.7 19.02 ;
  LAYER M3 ;
        RECT 0.668 16.532 0.7 16.564 ;
  LAYER M1 ;
        RECT 0.732 16.512 0.764 19.02 ;
  LAYER M3 ;
        RECT 0.732 18.968 0.764 19 ;
  LAYER M1 ;
        RECT 0.796 16.512 0.828 19.02 ;
  LAYER M3 ;
        RECT 0.796 16.532 0.828 16.564 ;
  LAYER M1 ;
        RECT 0.86 16.512 0.892 19.02 ;
  LAYER M3 ;
        RECT 0.86 18.968 0.892 19 ;
  LAYER M1 ;
        RECT 0.924 16.512 0.956 19.02 ;
  LAYER M3 ;
        RECT 0.924 16.532 0.956 16.564 ;
  LAYER M1 ;
        RECT 0.988 16.512 1.02 19.02 ;
  LAYER M3 ;
        RECT 0.988 18.968 1.02 19 ;
  LAYER M1 ;
        RECT 1.052 16.512 1.084 19.02 ;
  LAYER M3 ;
        RECT 1.052 16.532 1.084 16.564 ;
  LAYER M1 ;
        RECT 1.116 16.512 1.148 19.02 ;
  LAYER M3 ;
        RECT 1.116 18.968 1.148 19 ;
  LAYER M1 ;
        RECT 1.18 16.512 1.212 19.02 ;
  LAYER M3 ;
        RECT 1.18 16.532 1.212 16.564 ;
  LAYER M1 ;
        RECT 1.244 16.512 1.276 19.02 ;
  LAYER M3 ;
        RECT 1.244 18.968 1.276 19 ;
  LAYER M1 ;
        RECT 1.308 16.512 1.34 19.02 ;
  LAYER M3 ;
        RECT 1.308 16.532 1.34 16.564 ;
  LAYER M1 ;
        RECT 1.372 16.512 1.404 19.02 ;
  LAYER M3 ;
        RECT 1.372 18.968 1.404 19 ;
  LAYER M1 ;
        RECT 1.436 16.512 1.468 19.02 ;
  LAYER M3 ;
        RECT 1.436 16.532 1.468 16.564 ;
  LAYER M1 ;
        RECT 1.5 16.512 1.532 19.02 ;
  LAYER M3 ;
        RECT 1.5 18.968 1.532 19 ;
  LAYER M1 ;
        RECT 1.564 16.512 1.596 19.02 ;
  LAYER M3 ;
        RECT 1.564 16.532 1.596 16.564 ;
  LAYER M1 ;
        RECT 1.628 16.512 1.66 19.02 ;
  LAYER M3 ;
        RECT 1.628 18.968 1.66 19 ;
  LAYER M1 ;
        RECT 1.692 16.512 1.724 19.02 ;
  LAYER M3 ;
        RECT 1.692 16.532 1.724 16.564 ;
  LAYER M1 ;
        RECT 1.756 16.512 1.788 19.02 ;
  LAYER M3 ;
        RECT 1.756 18.968 1.788 19 ;
  LAYER M1 ;
        RECT 1.82 16.512 1.852 19.02 ;
  LAYER M3 ;
        RECT 1.82 16.532 1.852 16.564 ;
  LAYER M1 ;
        RECT 1.884 16.512 1.916 19.02 ;
  LAYER M3 ;
        RECT 1.884 18.968 1.916 19 ;
  LAYER M1 ;
        RECT 1.948 16.512 1.98 19.02 ;
  LAYER M3 ;
        RECT 1.948 16.532 1.98 16.564 ;
  LAYER M1 ;
        RECT 2.012 16.512 2.044 19.02 ;
  LAYER M3 ;
        RECT 2.012 18.968 2.044 19 ;
  LAYER M1 ;
        RECT 2.076 16.512 2.108 19.02 ;
  LAYER M3 ;
        RECT 2.076 16.532 2.108 16.564 ;
  LAYER M1 ;
        RECT 2.14 16.512 2.172 19.02 ;
  LAYER M3 ;
        RECT 2.14 18.968 2.172 19 ;
  LAYER M1 ;
        RECT 2.204 16.512 2.236 19.02 ;
  LAYER M3 ;
        RECT 2.204 16.532 2.236 16.564 ;
  LAYER M1 ;
        RECT 2.268 16.512 2.3 19.02 ;
  LAYER M3 ;
        RECT 2.268 18.968 2.3 19 ;
  LAYER M1 ;
        RECT 2.332 16.512 2.364 19.02 ;
  LAYER M3 ;
        RECT 2.332 16.532 2.364 16.564 ;
  LAYER M1 ;
        RECT 2.396 16.512 2.428 19.02 ;
  LAYER M3 ;
        RECT 2.396 18.968 2.428 19 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 19.02 ;
  LAYER M3 ;
        RECT 0.092 16.596 0.124 16.628 ;
  LAYER M2 ;
        RECT 2.46 16.66 2.492 16.692 ;
  LAYER M2 ;
        RECT 0.092 16.724 0.124 16.756 ;
  LAYER M2 ;
        RECT 2.46 16.788 2.492 16.82 ;
  LAYER M2 ;
        RECT 0.092 16.852 0.124 16.884 ;
  LAYER M2 ;
        RECT 2.46 16.916 2.492 16.948 ;
  LAYER M2 ;
        RECT 0.092 16.98 0.124 17.012 ;
  LAYER M2 ;
        RECT 2.46 17.044 2.492 17.076 ;
  LAYER M2 ;
        RECT 0.092 17.108 0.124 17.14 ;
  LAYER M2 ;
        RECT 2.46 17.172 2.492 17.204 ;
  LAYER M2 ;
        RECT 0.092 17.236 0.124 17.268 ;
  LAYER M2 ;
        RECT 2.46 17.3 2.492 17.332 ;
  LAYER M2 ;
        RECT 0.092 17.364 0.124 17.396 ;
  LAYER M2 ;
        RECT 2.46 17.428 2.492 17.46 ;
  LAYER M2 ;
        RECT 0.092 17.492 0.124 17.524 ;
  LAYER M2 ;
        RECT 2.46 17.556 2.492 17.588 ;
  LAYER M2 ;
        RECT 0.092 17.62 0.124 17.652 ;
  LAYER M2 ;
        RECT 2.46 17.684 2.492 17.716 ;
  LAYER M2 ;
        RECT 0.092 17.748 0.124 17.78 ;
  LAYER M2 ;
        RECT 2.46 17.812 2.492 17.844 ;
  LAYER M2 ;
        RECT 0.092 17.876 0.124 17.908 ;
  LAYER M2 ;
        RECT 2.46 17.94 2.492 17.972 ;
  LAYER M2 ;
        RECT 0.092 18.004 0.124 18.036 ;
  LAYER M2 ;
        RECT 2.46 18.068 2.492 18.1 ;
  LAYER M2 ;
        RECT 0.092 18.132 0.124 18.164 ;
  LAYER M2 ;
        RECT 2.46 18.196 2.492 18.228 ;
  LAYER M2 ;
        RECT 0.092 18.26 0.124 18.292 ;
  LAYER M2 ;
        RECT 2.46 18.324 2.492 18.356 ;
  LAYER M2 ;
        RECT 0.092 18.388 0.124 18.42 ;
  LAYER M2 ;
        RECT 2.46 18.452 2.492 18.484 ;
  LAYER M2 ;
        RECT 0.092 18.516 0.124 18.548 ;
  LAYER M2 ;
        RECT 2.46 18.58 2.492 18.612 ;
  LAYER M2 ;
        RECT 0.092 18.644 0.124 18.676 ;
  LAYER M2 ;
        RECT 2.46 18.708 2.492 18.74 ;
  LAYER M2 ;
        RECT 0.092 18.772 0.124 18.804 ;
  LAYER M2 ;
        RECT 2.46 18.836 2.492 18.868 ;
  LAYER M2 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M1 ;
        RECT 0.092 19.62 0.124 22.128 ;
  LAYER M3 ;
        RECT 0.092 22.076 0.124 22.108 ;
  LAYER M1 ;
        RECT 0.156 19.62 0.188 22.128 ;
  LAYER M3 ;
        RECT 0.156 19.64 0.188 19.672 ;
  LAYER M1 ;
        RECT 0.22 19.62 0.252 22.128 ;
  LAYER M3 ;
        RECT 0.22 22.076 0.252 22.108 ;
  LAYER M1 ;
        RECT 0.284 19.62 0.316 22.128 ;
  LAYER M3 ;
        RECT 0.284 19.64 0.316 19.672 ;
  LAYER M1 ;
        RECT 0.348 19.62 0.38 22.128 ;
  LAYER M3 ;
        RECT 0.348 22.076 0.38 22.108 ;
  LAYER M1 ;
        RECT 0.412 19.62 0.444 22.128 ;
  LAYER M3 ;
        RECT 0.412 19.64 0.444 19.672 ;
  LAYER M1 ;
        RECT 0.476 19.62 0.508 22.128 ;
  LAYER M3 ;
        RECT 0.476 22.076 0.508 22.108 ;
  LAYER M1 ;
        RECT 0.54 19.62 0.572 22.128 ;
  LAYER M3 ;
        RECT 0.54 19.64 0.572 19.672 ;
  LAYER M1 ;
        RECT 0.604 19.62 0.636 22.128 ;
  LAYER M3 ;
        RECT 0.604 22.076 0.636 22.108 ;
  LAYER M1 ;
        RECT 0.668 19.62 0.7 22.128 ;
  LAYER M3 ;
        RECT 0.668 19.64 0.7 19.672 ;
  LAYER M1 ;
        RECT 0.732 19.62 0.764 22.128 ;
  LAYER M3 ;
        RECT 0.732 22.076 0.764 22.108 ;
  LAYER M1 ;
        RECT 0.796 19.62 0.828 22.128 ;
  LAYER M3 ;
        RECT 0.796 19.64 0.828 19.672 ;
  LAYER M1 ;
        RECT 0.86 19.62 0.892 22.128 ;
  LAYER M3 ;
        RECT 0.86 22.076 0.892 22.108 ;
  LAYER M1 ;
        RECT 0.924 19.62 0.956 22.128 ;
  LAYER M3 ;
        RECT 0.924 19.64 0.956 19.672 ;
  LAYER M1 ;
        RECT 0.988 19.62 1.02 22.128 ;
  LAYER M3 ;
        RECT 0.988 22.076 1.02 22.108 ;
  LAYER M1 ;
        RECT 1.052 19.62 1.084 22.128 ;
  LAYER M3 ;
        RECT 1.052 19.64 1.084 19.672 ;
  LAYER M1 ;
        RECT 1.116 19.62 1.148 22.128 ;
  LAYER M3 ;
        RECT 1.116 22.076 1.148 22.108 ;
  LAYER M1 ;
        RECT 1.18 19.62 1.212 22.128 ;
  LAYER M3 ;
        RECT 1.18 19.64 1.212 19.672 ;
  LAYER M1 ;
        RECT 1.244 19.62 1.276 22.128 ;
  LAYER M3 ;
        RECT 1.244 22.076 1.276 22.108 ;
  LAYER M1 ;
        RECT 1.308 19.62 1.34 22.128 ;
  LAYER M3 ;
        RECT 1.308 19.64 1.34 19.672 ;
  LAYER M1 ;
        RECT 1.372 19.62 1.404 22.128 ;
  LAYER M3 ;
        RECT 1.372 22.076 1.404 22.108 ;
  LAYER M1 ;
        RECT 1.436 19.62 1.468 22.128 ;
  LAYER M3 ;
        RECT 1.436 19.64 1.468 19.672 ;
  LAYER M1 ;
        RECT 1.5 19.62 1.532 22.128 ;
  LAYER M3 ;
        RECT 1.5 22.076 1.532 22.108 ;
  LAYER M1 ;
        RECT 1.564 19.62 1.596 22.128 ;
  LAYER M3 ;
        RECT 1.564 19.64 1.596 19.672 ;
  LAYER M1 ;
        RECT 1.628 19.62 1.66 22.128 ;
  LAYER M3 ;
        RECT 1.628 22.076 1.66 22.108 ;
  LAYER M1 ;
        RECT 1.692 19.62 1.724 22.128 ;
  LAYER M3 ;
        RECT 1.692 19.64 1.724 19.672 ;
  LAYER M1 ;
        RECT 1.756 19.62 1.788 22.128 ;
  LAYER M3 ;
        RECT 1.756 22.076 1.788 22.108 ;
  LAYER M1 ;
        RECT 1.82 19.62 1.852 22.128 ;
  LAYER M3 ;
        RECT 1.82 19.64 1.852 19.672 ;
  LAYER M1 ;
        RECT 1.884 19.62 1.916 22.128 ;
  LAYER M3 ;
        RECT 1.884 22.076 1.916 22.108 ;
  LAYER M1 ;
        RECT 1.948 19.62 1.98 22.128 ;
  LAYER M3 ;
        RECT 1.948 19.64 1.98 19.672 ;
  LAYER M1 ;
        RECT 2.012 19.62 2.044 22.128 ;
  LAYER M3 ;
        RECT 2.012 22.076 2.044 22.108 ;
  LAYER M1 ;
        RECT 2.076 19.62 2.108 22.128 ;
  LAYER M3 ;
        RECT 2.076 19.64 2.108 19.672 ;
  LAYER M1 ;
        RECT 2.14 19.62 2.172 22.128 ;
  LAYER M3 ;
        RECT 2.14 22.076 2.172 22.108 ;
  LAYER M1 ;
        RECT 2.204 19.62 2.236 22.128 ;
  LAYER M3 ;
        RECT 2.204 19.64 2.236 19.672 ;
  LAYER M1 ;
        RECT 2.268 19.62 2.3 22.128 ;
  LAYER M3 ;
        RECT 2.268 22.076 2.3 22.108 ;
  LAYER M1 ;
        RECT 2.332 19.62 2.364 22.128 ;
  LAYER M3 ;
        RECT 2.332 19.64 2.364 19.672 ;
  LAYER M1 ;
        RECT 2.396 19.62 2.428 22.128 ;
  LAYER M3 ;
        RECT 2.396 22.076 2.428 22.108 ;
  LAYER M1 ;
        RECT 2.46 19.62 2.492 22.128 ;
  LAYER M3 ;
        RECT 0.092 19.704 0.124 19.736 ;
  LAYER M2 ;
        RECT 2.46 19.768 2.492 19.8 ;
  LAYER M2 ;
        RECT 0.092 19.832 0.124 19.864 ;
  LAYER M2 ;
        RECT 2.46 19.896 2.492 19.928 ;
  LAYER M2 ;
        RECT 0.092 19.96 0.124 19.992 ;
  LAYER M2 ;
        RECT 2.46 20.024 2.492 20.056 ;
  LAYER M2 ;
        RECT 0.092 20.088 0.124 20.12 ;
  LAYER M2 ;
        RECT 2.46 20.152 2.492 20.184 ;
  LAYER M2 ;
        RECT 0.092 20.216 0.124 20.248 ;
  LAYER M2 ;
        RECT 2.46 20.28 2.492 20.312 ;
  LAYER M2 ;
        RECT 0.092 20.344 0.124 20.376 ;
  LAYER M2 ;
        RECT 2.46 20.408 2.492 20.44 ;
  LAYER M2 ;
        RECT 0.092 20.472 0.124 20.504 ;
  LAYER M2 ;
        RECT 2.46 20.536 2.492 20.568 ;
  LAYER M2 ;
        RECT 0.092 20.6 0.124 20.632 ;
  LAYER M2 ;
        RECT 2.46 20.664 2.492 20.696 ;
  LAYER M2 ;
        RECT 0.092 20.728 0.124 20.76 ;
  LAYER M2 ;
        RECT 2.46 20.792 2.492 20.824 ;
  LAYER M2 ;
        RECT 0.092 20.856 0.124 20.888 ;
  LAYER M2 ;
        RECT 2.46 20.92 2.492 20.952 ;
  LAYER M2 ;
        RECT 0.092 20.984 0.124 21.016 ;
  LAYER M2 ;
        RECT 2.46 21.048 2.492 21.08 ;
  LAYER M2 ;
        RECT 0.092 21.112 0.124 21.144 ;
  LAYER M2 ;
        RECT 2.46 21.176 2.492 21.208 ;
  LAYER M2 ;
        RECT 0.092 21.24 0.124 21.272 ;
  LAYER M2 ;
        RECT 2.46 21.304 2.492 21.336 ;
  LAYER M2 ;
        RECT 0.092 21.368 0.124 21.4 ;
  LAYER M2 ;
        RECT 2.46 21.432 2.492 21.464 ;
  LAYER M2 ;
        RECT 0.092 21.496 0.124 21.528 ;
  LAYER M2 ;
        RECT 2.46 21.56 2.492 21.592 ;
  LAYER M2 ;
        RECT 0.092 21.624 0.124 21.656 ;
  LAYER M2 ;
        RECT 2.46 21.688 2.492 21.72 ;
  LAYER M2 ;
        RECT 0.092 21.752 0.124 21.784 ;
  LAYER M2 ;
        RECT 2.46 21.816 2.492 21.848 ;
  LAYER M2 ;
        RECT 0.092 21.88 0.124 21.912 ;
  LAYER M2 ;
        RECT 2.46 21.944 2.492 21.976 ;
  LAYER M2 ;
        RECT 0.044 19.572 2.54 22.176 ;
  LAYER M1 ;
        RECT 3.388 0.972 3.42 3.48 ;
  LAYER M3 ;
        RECT 3.388 3.428 3.42 3.46 ;
  LAYER M1 ;
        RECT 3.452 0.972 3.484 3.48 ;
  LAYER M3 ;
        RECT 3.452 0.992 3.484 1.024 ;
  LAYER M1 ;
        RECT 3.516 0.972 3.548 3.48 ;
  LAYER M3 ;
        RECT 3.516 3.428 3.548 3.46 ;
  LAYER M1 ;
        RECT 3.58 0.972 3.612 3.48 ;
  LAYER M3 ;
        RECT 3.58 0.992 3.612 1.024 ;
  LAYER M1 ;
        RECT 3.644 0.972 3.676 3.48 ;
  LAYER M3 ;
        RECT 3.644 3.428 3.676 3.46 ;
  LAYER M1 ;
        RECT 3.708 0.972 3.74 3.48 ;
  LAYER M3 ;
        RECT 3.708 0.992 3.74 1.024 ;
  LAYER M1 ;
        RECT 3.772 0.972 3.804 3.48 ;
  LAYER M3 ;
        RECT 3.772 3.428 3.804 3.46 ;
  LAYER M1 ;
        RECT 3.836 0.972 3.868 3.48 ;
  LAYER M3 ;
        RECT 3.836 0.992 3.868 1.024 ;
  LAYER M1 ;
        RECT 3.9 0.972 3.932 3.48 ;
  LAYER M3 ;
        RECT 3.9 3.428 3.932 3.46 ;
  LAYER M1 ;
        RECT 3.964 0.972 3.996 3.48 ;
  LAYER M3 ;
        RECT 3.964 0.992 3.996 1.024 ;
  LAYER M1 ;
        RECT 4.028 0.972 4.06 3.48 ;
  LAYER M3 ;
        RECT 4.028 3.428 4.06 3.46 ;
  LAYER M1 ;
        RECT 4.092 0.972 4.124 3.48 ;
  LAYER M3 ;
        RECT 4.092 0.992 4.124 1.024 ;
  LAYER M1 ;
        RECT 4.156 0.972 4.188 3.48 ;
  LAYER M3 ;
        RECT 4.156 3.428 4.188 3.46 ;
  LAYER M1 ;
        RECT 4.22 0.972 4.252 3.48 ;
  LAYER M3 ;
        RECT 4.22 0.992 4.252 1.024 ;
  LAYER M1 ;
        RECT 4.284 0.972 4.316 3.48 ;
  LAYER M3 ;
        RECT 4.284 3.428 4.316 3.46 ;
  LAYER M1 ;
        RECT 4.348 0.972 4.38 3.48 ;
  LAYER M3 ;
        RECT 4.348 0.992 4.38 1.024 ;
  LAYER M1 ;
        RECT 4.412 0.972 4.444 3.48 ;
  LAYER M3 ;
        RECT 4.412 3.428 4.444 3.46 ;
  LAYER M1 ;
        RECT 4.476 0.972 4.508 3.48 ;
  LAYER M3 ;
        RECT 4.476 0.992 4.508 1.024 ;
  LAYER M1 ;
        RECT 4.54 0.972 4.572 3.48 ;
  LAYER M3 ;
        RECT 4.54 3.428 4.572 3.46 ;
  LAYER M1 ;
        RECT 4.604 0.972 4.636 3.48 ;
  LAYER M3 ;
        RECT 4.604 0.992 4.636 1.024 ;
  LAYER M1 ;
        RECT 4.668 0.972 4.7 3.48 ;
  LAYER M3 ;
        RECT 4.668 3.428 4.7 3.46 ;
  LAYER M1 ;
        RECT 4.732 0.972 4.764 3.48 ;
  LAYER M3 ;
        RECT 4.732 0.992 4.764 1.024 ;
  LAYER M1 ;
        RECT 4.796 0.972 4.828 3.48 ;
  LAYER M3 ;
        RECT 4.796 3.428 4.828 3.46 ;
  LAYER M1 ;
        RECT 4.86 0.972 4.892 3.48 ;
  LAYER M3 ;
        RECT 4.86 0.992 4.892 1.024 ;
  LAYER M1 ;
        RECT 4.924 0.972 4.956 3.48 ;
  LAYER M3 ;
        RECT 4.924 3.428 4.956 3.46 ;
  LAYER M1 ;
        RECT 4.988 0.972 5.02 3.48 ;
  LAYER M3 ;
        RECT 4.988 0.992 5.02 1.024 ;
  LAYER M1 ;
        RECT 5.052 0.972 5.084 3.48 ;
  LAYER M3 ;
        RECT 5.052 3.428 5.084 3.46 ;
  LAYER M1 ;
        RECT 5.116 0.972 5.148 3.48 ;
  LAYER M3 ;
        RECT 5.116 0.992 5.148 1.024 ;
  LAYER M1 ;
        RECT 5.18 0.972 5.212 3.48 ;
  LAYER M3 ;
        RECT 5.18 3.428 5.212 3.46 ;
  LAYER M1 ;
        RECT 5.244 0.972 5.276 3.48 ;
  LAYER M3 ;
        RECT 5.244 0.992 5.276 1.024 ;
  LAYER M1 ;
        RECT 5.308 0.972 5.34 3.48 ;
  LAYER M3 ;
        RECT 5.308 3.428 5.34 3.46 ;
  LAYER M1 ;
        RECT 5.372 0.972 5.404 3.48 ;
  LAYER M3 ;
        RECT 5.372 0.992 5.404 1.024 ;
  LAYER M1 ;
        RECT 5.436 0.972 5.468 3.48 ;
  LAYER M3 ;
        RECT 5.436 3.428 5.468 3.46 ;
  LAYER M1 ;
        RECT 5.5 0.972 5.532 3.48 ;
  LAYER M3 ;
        RECT 5.5 0.992 5.532 1.024 ;
  LAYER M1 ;
        RECT 5.564 0.972 5.596 3.48 ;
  LAYER M3 ;
        RECT 5.564 3.428 5.596 3.46 ;
  LAYER M1 ;
        RECT 5.628 0.972 5.66 3.48 ;
  LAYER M3 ;
        RECT 5.628 0.992 5.66 1.024 ;
  LAYER M1 ;
        RECT 5.692 0.972 5.724 3.48 ;
  LAYER M3 ;
        RECT 5.692 3.428 5.724 3.46 ;
  LAYER M1 ;
        RECT 5.756 0.972 5.788 3.48 ;
  LAYER M3 ;
        RECT 3.388 1.056 3.42 1.088 ;
  LAYER M2 ;
        RECT 5.756 1.12 5.788 1.152 ;
  LAYER M2 ;
        RECT 3.388 1.184 3.42 1.216 ;
  LAYER M2 ;
        RECT 5.756 1.248 5.788 1.28 ;
  LAYER M2 ;
        RECT 3.388 1.312 3.42 1.344 ;
  LAYER M2 ;
        RECT 5.756 1.376 5.788 1.408 ;
  LAYER M2 ;
        RECT 3.388 1.44 3.42 1.472 ;
  LAYER M2 ;
        RECT 5.756 1.504 5.788 1.536 ;
  LAYER M2 ;
        RECT 3.388 1.568 3.42 1.6 ;
  LAYER M2 ;
        RECT 5.756 1.632 5.788 1.664 ;
  LAYER M2 ;
        RECT 3.388 1.696 3.42 1.728 ;
  LAYER M2 ;
        RECT 5.756 1.76 5.788 1.792 ;
  LAYER M2 ;
        RECT 3.388 1.824 3.42 1.856 ;
  LAYER M2 ;
        RECT 5.756 1.888 5.788 1.92 ;
  LAYER M2 ;
        RECT 3.388 1.952 3.42 1.984 ;
  LAYER M2 ;
        RECT 5.756 2.016 5.788 2.048 ;
  LAYER M2 ;
        RECT 3.388 2.08 3.42 2.112 ;
  LAYER M2 ;
        RECT 5.756 2.144 5.788 2.176 ;
  LAYER M2 ;
        RECT 3.388 2.208 3.42 2.24 ;
  LAYER M2 ;
        RECT 5.756 2.272 5.788 2.304 ;
  LAYER M2 ;
        RECT 3.388 2.336 3.42 2.368 ;
  LAYER M2 ;
        RECT 5.756 2.4 5.788 2.432 ;
  LAYER M2 ;
        RECT 3.388 2.464 3.42 2.496 ;
  LAYER M2 ;
        RECT 5.756 2.528 5.788 2.56 ;
  LAYER M2 ;
        RECT 3.388 2.592 3.42 2.624 ;
  LAYER M2 ;
        RECT 5.756 2.656 5.788 2.688 ;
  LAYER M2 ;
        RECT 3.388 2.72 3.42 2.752 ;
  LAYER M2 ;
        RECT 5.756 2.784 5.788 2.816 ;
  LAYER M2 ;
        RECT 3.388 2.848 3.42 2.88 ;
  LAYER M2 ;
        RECT 5.756 2.912 5.788 2.944 ;
  LAYER M2 ;
        RECT 3.388 2.976 3.42 3.008 ;
  LAYER M2 ;
        RECT 5.756 3.04 5.788 3.072 ;
  LAYER M2 ;
        RECT 3.388 3.104 3.42 3.136 ;
  LAYER M2 ;
        RECT 5.756 3.168 5.788 3.2 ;
  LAYER M2 ;
        RECT 3.388 3.232 3.42 3.264 ;
  LAYER M2 ;
        RECT 5.756 3.296 5.788 3.328 ;
  LAYER M2 ;
        RECT 3.34 0.924 5.836 3.528 ;
  LAYER M1 ;
        RECT 3.388 4.08 3.42 6.588 ;
  LAYER M3 ;
        RECT 3.388 6.536 3.42 6.568 ;
  LAYER M1 ;
        RECT 3.452 4.08 3.484 6.588 ;
  LAYER M3 ;
        RECT 3.452 4.1 3.484 4.132 ;
  LAYER M1 ;
        RECT 3.516 4.08 3.548 6.588 ;
  LAYER M3 ;
        RECT 3.516 6.536 3.548 6.568 ;
  LAYER M1 ;
        RECT 3.58 4.08 3.612 6.588 ;
  LAYER M3 ;
        RECT 3.58 4.1 3.612 4.132 ;
  LAYER M1 ;
        RECT 3.644 4.08 3.676 6.588 ;
  LAYER M3 ;
        RECT 3.644 6.536 3.676 6.568 ;
  LAYER M1 ;
        RECT 3.708 4.08 3.74 6.588 ;
  LAYER M3 ;
        RECT 3.708 4.1 3.74 4.132 ;
  LAYER M1 ;
        RECT 3.772 4.08 3.804 6.588 ;
  LAYER M3 ;
        RECT 3.772 6.536 3.804 6.568 ;
  LAYER M1 ;
        RECT 3.836 4.08 3.868 6.588 ;
  LAYER M3 ;
        RECT 3.836 4.1 3.868 4.132 ;
  LAYER M1 ;
        RECT 3.9 4.08 3.932 6.588 ;
  LAYER M3 ;
        RECT 3.9 6.536 3.932 6.568 ;
  LAYER M1 ;
        RECT 3.964 4.08 3.996 6.588 ;
  LAYER M3 ;
        RECT 3.964 4.1 3.996 4.132 ;
  LAYER M1 ;
        RECT 4.028 4.08 4.06 6.588 ;
  LAYER M3 ;
        RECT 4.028 6.536 4.06 6.568 ;
  LAYER M1 ;
        RECT 4.092 4.08 4.124 6.588 ;
  LAYER M3 ;
        RECT 4.092 4.1 4.124 4.132 ;
  LAYER M1 ;
        RECT 4.156 4.08 4.188 6.588 ;
  LAYER M3 ;
        RECT 4.156 6.536 4.188 6.568 ;
  LAYER M1 ;
        RECT 4.22 4.08 4.252 6.588 ;
  LAYER M3 ;
        RECT 4.22 4.1 4.252 4.132 ;
  LAYER M1 ;
        RECT 4.284 4.08 4.316 6.588 ;
  LAYER M3 ;
        RECT 4.284 6.536 4.316 6.568 ;
  LAYER M1 ;
        RECT 4.348 4.08 4.38 6.588 ;
  LAYER M3 ;
        RECT 4.348 4.1 4.38 4.132 ;
  LAYER M1 ;
        RECT 4.412 4.08 4.444 6.588 ;
  LAYER M3 ;
        RECT 4.412 6.536 4.444 6.568 ;
  LAYER M1 ;
        RECT 4.476 4.08 4.508 6.588 ;
  LAYER M3 ;
        RECT 4.476 4.1 4.508 4.132 ;
  LAYER M1 ;
        RECT 4.54 4.08 4.572 6.588 ;
  LAYER M3 ;
        RECT 4.54 6.536 4.572 6.568 ;
  LAYER M1 ;
        RECT 4.604 4.08 4.636 6.588 ;
  LAYER M3 ;
        RECT 4.604 4.1 4.636 4.132 ;
  LAYER M1 ;
        RECT 4.668 4.08 4.7 6.588 ;
  LAYER M3 ;
        RECT 4.668 6.536 4.7 6.568 ;
  LAYER M1 ;
        RECT 4.732 4.08 4.764 6.588 ;
  LAYER M3 ;
        RECT 4.732 4.1 4.764 4.132 ;
  LAYER M1 ;
        RECT 4.796 4.08 4.828 6.588 ;
  LAYER M3 ;
        RECT 4.796 6.536 4.828 6.568 ;
  LAYER M1 ;
        RECT 4.86 4.08 4.892 6.588 ;
  LAYER M3 ;
        RECT 4.86 4.1 4.892 4.132 ;
  LAYER M1 ;
        RECT 4.924 4.08 4.956 6.588 ;
  LAYER M3 ;
        RECT 4.924 6.536 4.956 6.568 ;
  LAYER M1 ;
        RECT 4.988 4.08 5.02 6.588 ;
  LAYER M3 ;
        RECT 4.988 4.1 5.02 4.132 ;
  LAYER M1 ;
        RECT 5.052 4.08 5.084 6.588 ;
  LAYER M3 ;
        RECT 5.052 6.536 5.084 6.568 ;
  LAYER M1 ;
        RECT 5.116 4.08 5.148 6.588 ;
  LAYER M3 ;
        RECT 5.116 4.1 5.148 4.132 ;
  LAYER M1 ;
        RECT 5.18 4.08 5.212 6.588 ;
  LAYER M3 ;
        RECT 5.18 6.536 5.212 6.568 ;
  LAYER M1 ;
        RECT 5.244 4.08 5.276 6.588 ;
  LAYER M3 ;
        RECT 5.244 4.1 5.276 4.132 ;
  LAYER M1 ;
        RECT 5.308 4.08 5.34 6.588 ;
  LAYER M3 ;
        RECT 5.308 6.536 5.34 6.568 ;
  LAYER M1 ;
        RECT 5.372 4.08 5.404 6.588 ;
  LAYER M3 ;
        RECT 5.372 4.1 5.404 4.132 ;
  LAYER M1 ;
        RECT 5.436 4.08 5.468 6.588 ;
  LAYER M3 ;
        RECT 5.436 6.536 5.468 6.568 ;
  LAYER M1 ;
        RECT 5.5 4.08 5.532 6.588 ;
  LAYER M3 ;
        RECT 5.5 4.1 5.532 4.132 ;
  LAYER M1 ;
        RECT 5.564 4.08 5.596 6.588 ;
  LAYER M3 ;
        RECT 5.564 6.536 5.596 6.568 ;
  LAYER M1 ;
        RECT 5.628 4.08 5.66 6.588 ;
  LAYER M3 ;
        RECT 5.628 4.1 5.66 4.132 ;
  LAYER M1 ;
        RECT 5.692 4.08 5.724 6.588 ;
  LAYER M3 ;
        RECT 5.692 6.536 5.724 6.568 ;
  LAYER M1 ;
        RECT 5.756 4.08 5.788 6.588 ;
  LAYER M3 ;
        RECT 3.388 4.164 3.42 4.196 ;
  LAYER M2 ;
        RECT 5.756 4.228 5.788 4.26 ;
  LAYER M2 ;
        RECT 3.388 4.292 3.42 4.324 ;
  LAYER M2 ;
        RECT 5.756 4.356 5.788 4.388 ;
  LAYER M2 ;
        RECT 3.388 4.42 3.42 4.452 ;
  LAYER M2 ;
        RECT 5.756 4.484 5.788 4.516 ;
  LAYER M2 ;
        RECT 3.388 4.548 3.42 4.58 ;
  LAYER M2 ;
        RECT 5.756 4.612 5.788 4.644 ;
  LAYER M2 ;
        RECT 3.388 4.676 3.42 4.708 ;
  LAYER M2 ;
        RECT 5.756 4.74 5.788 4.772 ;
  LAYER M2 ;
        RECT 3.388 4.804 3.42 4.836 ;
  LAYER M2 ;
        RECT 5.756 4.868 5.788 4.9 ;
  LAYER M2 ;
        RECT 3.388 4.932 3.42 4.964 ;
  LAYER M2 ;
        RECT 5.756 4.996 5.788 5.028 ;
  LAYER M2 ;
        RECT 3.388 5.06 3.42 5.092 ;
  LAYER M2 ;
        RECT 5.756 5.124 5.788 5.156 ;
  LAYER M2 ;
        RECT 3.388 5.188 3.42 5.22 ;
  LAYER M2 ;
        RECT 5.756 5.252 5.788 5.284 ;
  LAYER M2 ;
        RECT 3.388 5.316 3.42 5.348 ;
  LAYER M2 ;
        RECT 5.756 5.38 5.788 5.412 ;
  LAYER M2 ;
        RECT 3.388 5.444 3.42 5.476 ;
  LAYER M2 ;
        RECT 5.756 5.508 5.788 5.54 ;
  LAYER M2 ;
        RECT 3.388 5.572 3.42 5.604 ;
  LAYER M2 ;
        RECT 5.756 5.636 5.788 5.668 ;
  LAYER M2 ;
        RECT 3.388 5.7 3.42 5.732 ;
  LAYER M2 ;
        RECT 5.756 5.764 5.788 5.796 ;
  LAYER M2 ;
        RECT 3.388 5.828 3.42 5.86 ;
  LAYER M2 ;
        RECT 5.756 5.892 5.788 5.924 ;
  LAYER M2 ;
        RECT 3.388 5.956 3.42 5.988 ;
  LAYER M2 ;
        RECT 5.756 6.02 5.788 6.052 ;
  LAYER M2 ;
        RECT 3.388 6.084 3.42 6.116 ;
  LAYER M2 ;
        RECT 5.756 6.148 5.788 6.18 ;
  LAYER M2 ;
        RECT 3.388 6.212 3.42 6.244 ;
  LAYER M2 ;
        RECT 5.756 6.276 5.788 6.308 ;
  LAYER M2 ;
        RECT 3.388 6.34 3.42 6.372 ;
  LAYER M2 ;
        RECT 5.756 6.404 5.788 6.436 ;
  LAYER M2 ;
        RECT 3.34 4.032 5.836 6.636 ;
  LAYER M1 ;
        RECT 3.388 7.188 3.42 9.696 ;
  LAYER M3 ;
        RECT 3.388 9.644 3.42 9.676 ;
  LAYER M1 ;
        RECT 3.452 7.188 3.484 9.696 ;
  LAYER M3 ;
        RECT 3.452 7.208 3.484 7.24 ;
  LAYER M1 ;
        RECT 3.516 7.188 3.548 9.696 ;
  LAYER M3 ;
        RECT 3.516 9.644 3.548 9.676 ;
  LAYER M1 ;
        RECT 3.58 7.188 3.612 9.696 ;
  LAYER M3 ;
        RECT 3.58 7.208 3.612 7.24 ;
  LAYER M1 ;
        RECT 3.644 7.188 3.676 9.696 ;
  LAYER M3 ;
        RECT 3.644 9.644 3.676 9.676 ;
  LAYER M1 ;
        RECT 3.708 7.188 3.74 9.696 ;
  LAYER M3 ;
        RECT 3.708 7.208 3.74 7.24 ;
  LAYER M1 ;
        RECT 3.772 7.188 3.804 9.696 ;
  LAYER M3 ;
        RECT 3.772 9.644 3.804 9.676 ;
  LAYER M1 ;
        RECT 3.836 7.188 3.868 9.696 ;
  LAYER M3 ;
        RECT 3.836 7.208 3.868 7.24 ;
  LAYER M1 ;
        RECT 3.9 7.188 3.932 9.696 ;
  LAYER M3 ;
        RECT 3.9 9.644 3.932 9.676 ;
  LAYER M1 ;
        RECT 3.964 7.188 3.996 9.696 ;
  LAYER M3 ;
        RECT 3.964 7.208 3.996 7.24 ;
  LAYER M1 ;
        RECT 4.028 7.188 4.06 9.696 ;
  LAYER M3 ;
        RECT 4.028 9.644 4.06 9.676 ;
  LAYER M1 ;
        RECT 4.092 7.188 4.124 9.696 ;
  LAYER M3 ;
        RECT 4.092 7.208 4.124 7.24 ;
  LAYER M1 ;
        RECT 4.156 7.188 4.188 9.696 ;
  LAYER M3 ;
        RECT 4.156 9.644 4.188 9.676 ;
  LAYER M1 ;
        RECT 4.22 7.188 4.252 9.696 ;
  LAYER M3 ;
        RECT 4.22 7.208 4.252 7.24 ;
  LAYER M1 ;
        RECT 4.284 7.188 4.316 9.696 ;
  LAYER M3 ;
        RECT 4.284 9.644 4.316 9.676 ;
  LAYER M1 ;
        RECT 4.348 7.188 4.38 9.696 ;
  LAYER M3 ;
        RECT 4.348 7.208 4.38 7.24 ;
  LAYER M1 ;
        RECT 4.412 7.188 4.444 9.696 ;
  LAYER M3 ;
        RECT 4.412 9.644 4.444 9.676 ;
  LAYER M1 ;
        RECT 4.476 7.188 4.508 9.696 ;
  LAYER M3 ;
        RECT 4.476 7.208 4.508 7.24 ;
  LAYER M1 ;
        RECT 4.54 7.188 4.572 9.696 ;
  LAYER M3 ;
        RECT 4.54 9.644 4.572 9.676 ;
  LAYER M1 ;
        RECT 4.604 7.188 4.636 9.696 ;
  LAYER M3 ;
        RECT 4.604 7.208 4.636 7.24 ;
  LAYER M1 ;
        RECT 4.668 7.188 4.7 9.696 ;
  LAYER M3 ;
        RECT 4.668 9.644 4.7 9.676 ;
  LAYER M1 ;
        RECT 4.732 7.188 4.764 9.696 ;
  LAYER M3 ;
        RECT 4.732 7.208 4.764 7.24 ;
  LAYER M1 ;
        RECT 4.796 7.188 4.828 9.696 ;
  LAYER M3 ;
        RECT 4.796 9.644 4.828 9.676 ;
  LAYER M1 ;
        RECT 4.86 7.188 4.892 9.696 ;
  LAYER M3 ;
        RECT 4.86 7.208 4.892 7.24 ;
  LAYER M1 ;
        RECT 4.924 7.188 4.956 9.696 ;
  LAYER M3 ;
        RECT 4.924 9.644 4.956 9.676 ;
  LAYER M1 ;
        RECT 4.988 7.188 5.02 9.696 ;
  LAYER M3 ;
        RECT 4.988 7.208 5.02 7.24 ;
  LAYER M1 ;
        RECT 5.052 7.188 5.084 9.696 ;
  LAYER M3 ;
        RECT 5.052 9.644 5.084 9.676 ;
  LAYER M1 ;
        RECT 5.116 7.188 5.148 9.696 ;
  LAYER M3 ;
        RECT 5.116 7.208 5.148 7.24 ;
  LAYER M1 ;
        RECT 5.18 7.188 5.212 9.696 ;
  LAYER M3 ;
        RECT 5.18 9.644 5.212 9.676 ;
  LAYER M1 ;
        RECT 5.244 7.188 5.276 9.696 ;
  LAYER M3 ;
        RECT 5.244 7.208 5.276 7.24 ;
  LAYER M1 ;
        RECT 5.308 7.188 5.34 9.696 ;
  LAYER M3 ;
        RECT 5.308 9.644 5.34 9.676 ;
  LAYER M1 ;
        RECT 5.372 7.188 5.404 9.696 ;
  LAYER M3 ;
        RECT 5.372 7.208 5.404 7.24 ;
  LAYER M1 ;
        RECT 5.436 7.188 5.468 9.696 ;
  LAYER M3 ;
        RECT 5.436 9.644 5.468 9.676 ;
  LAYER M1 ;
        RECT 5.5 7.188 5.532 9.696 ;
  LAYER M3 ;
        RECT 5.5 7.208 5.532 7.24 ;
  LAYER M1 ;
        RECT 5.564 7.188 5.596 9.696 ;
  LAYER M3 ;
        RECT 5.564 9.644 5.596 9.676 ;
  LAYER M1 ;
        RECT 5.628 7.188 5.66 9.696 ;
  LAYER M3 ;
        RECT 5.628 7.208 5.66 7.24 ;
  LAYER M1 ;
        RECT 5.692 7.188 5.724 9.696 ;
  LAYER M3 ;
        RECT 5.692 9.644 5.724 9.676 ;
  LAYER M1 ;
        RECT 5.756 7.188 5.788 9.696 ;
  LAYER M3 ;
        RECT 3.388 7.272 3.42 7.304 ;
  LAYER M2 ;
        RECT 5.756 7.336 5.788 7.368 ;
  LAYER M2 ;
        RECT 3.388 7.4 3.42 7.432 ;
  LAYER M2 ;
        RECT 5.756 7.464 5.788 7.496 ;
  LAYER M2 ;
        RECT 3.388 7.528 3.42 7.56 ;
  LAYER M2 ;
        RECT 5.756 7.592 5.788 7.624 ;
  LAYER M2 ;
        RECT 3.388 7.656 3.42 7.688 ;
  LAYER M2 ;
        RECT 5.756 7.72 5.788 7.752 ;
  LAYER M2 ;
        RECT 3.388 7.784 3.42 7.816 ;
  LAYER M2 ;
        RECT 5.756 7.848 5.788 7.88 ;
  LAYER M2 ;
        RECT 3.388 7.912 3.42 7.944 ;
  LAYER M2 ;
        RECT 5.756 7.976 5.788 8.008 ;
  LAYER M2 ;
        RECT 3.388 8.04 3.42 8.072 ;
  LAYER M2 ;
        RECT 5.756 8.104 5.788 8.136 ;
  LAYER M2 ;
        RECT 3.388 8.168 3.42 8.2 ;
  LAYER M2 ;
        RECT 5.756 8.232 5.788 8.264 ;
  LAYER M2 ;
        RECT 3.388 8.296 3.42 8.328 ;
  LAYER M2 ;
        RECT 5.756 8.36 5.788 8.392 ;
  LAYER M2 ;
        RECT 3.388 8.424 3.42 8.456 ;
  LAYER M2 ;
        RECT 5.756 8.488 5.788 8.52 ;
  LAYER M2 ;
        RECT 3.388 8.552 3.42 8.584 ;
  LAYER M2 ;
        RECT 5.756 8.616 5.788 8.648 ;
  LAYER M2 ;
        RECT 3.388 8.68 3.42 8.712 ;
  LAYER M2 ;
        RECT 5.756 8.744 5.788 8.776 ;
  LAYER M2 ;
        RECT 3.388 8.808 3.42 8.84 ;
  LAYER M2 ;
        RECT 5.756 8.872 5.788 8.904 ;
  LAYER M2 ;
        RECT 3.388 8.936 3.42 8.968 ;
  LAYER M2 ;
        RECT 5.756 9 5.788 9.032 ;
  LAYER M2 ;
        RECT 3.388 9.064 3.42 9.096 ;
  LAYER M2 ;
        RECT 5.756 9.128 5.788 9.16 ;
  LAYER M2 ;
        RECT 3.388 9.192 3.42 9.224 ;
  LAYER M2 ;
        RECT 5.756 9.256 5.788 9.288 ;
  LAYER M2 ;
        RECT 3.388 9.32 3.42 9.352 ;
  LAYER M2 ;
        RECT 5.756 9.384 5.788 9.416 ;
  LAYER M2 ;
        RECT 3.388 9.448 3.42 9.48 ;
  LAYER M2 ;
        RECT 5.756 9.512 5.788 9.544 ;
  LAYER M2 ;
        RECT 3.34 7.14 5.836 9.744 ;
  LAYER M1 ;
        RECT 3.388 10.296 3.42 12.804 ;
  LAYER M3 ;
        RECT 3.388 12.752 3.42 12.784 ;
  LAYER M1 ;
        RECT 3.452 10.296 3.484 12.804 ;
  LAYER M3 ;
        RECT 3.452 10.316 3.484 10.348 ;
  LAYER M1 ;
        RECT 3.516 10.296 3.548 12.804 ;
  LAYER M3 ;
        RECT 3.516 12.752 3.548 12.784 ;
  LAYER M1 ;
        RECT 3.58 10.296 3.612 12.804 ;
  LAYER M3 ;
        RECT 3.58 10.316 3.612 10.348 ;
  LAYER M1 ;
        RECT 3.644 10.296 3.676 12.804 ;
  LAYER M3 ;
        RECT 3.644 12.752 3.676 12.784 ;
  LAYER M1 ;
        RECT 3.708 10.296 3.74 12.804 ;
  LAYER M3 ;
        RECT 3.708 10.316 3.74 10.348 ;
  LAYER M1 ;
        RECT 3.772 10.296 3.804 12.804 ;
  LAYER M3 ;
        RECT 3.772 12.752 3.804 12.784 ;
  LAYER M1 ;
        RECT 3.836 10.296 3.868 12.804 ;
  LAYER M3 ;
        RECT 3.836 10.316 3.868 10.348 ;
  LAYER M1 ;
        RECT 3.9 10.296 3.932 12.804 ;
  LAYER M3 ;
        RECT 3.9 12.752 3.932 12.784 ;
  LAYER M1 ;
        RECT 3.964 10.296 3.996 12.804 ;
  LAYER M3 ;
        RECT 3.964 10.316 3.996 10.348 ;
  LAYER M1 ;
        RECT 4.028 10.296 4.06 12.804 ;
  LAYER M3 ;
        RECT 4.028 12.752 4.06 12.784 ;
  LAYER M1 ;
        RECT 4.092 10.296 4.124 12.804 ;
  LAYER M3 ;
        RECT 4.092 10.316 4.124 10.348 ;
  LAYER M1 ;
        RECT 4.156 10.296 4.188 12.804 ;
  LAYER M3 ;
        RECT 4.156 12.752 4.188 12.784 ;
  LAYER M1 ;
        RECT 4.22 10.296 4.252 12.804 ;
  LAYER M3 ;
        RECT 4.22 10.316 4.252 10.348 ;
  LAYER M1 ;
        RECT 4.284 10.296 4.316 12.804 ;
  LAYER M3 ;
        RECT 4.284 12.752 4.316 12.784 ;
  LAYER M1 ;
        RECT 4.348 10.296 4.38 12.804 ;
  LAYER M3 ;
        RECT 4.348 10.316 4.38 10.348 ;
  LAYER M1 ;
        RECT 4.412 10.296 4.444 12.804 ;
  LAYER M3 ;
        RECT 4.412 12.752 4.444 12.784 ;
  LAYER M1 ;
        RECT 4.476 10.296 4.508 12.804 ;
  LAYER M3 ;
        RECT 4.476 10.316 4.508 10.348 ;
  LAYER M1 ;
        RECT 4.54 10.296 4.572 12.804 ;
  LAYER M3 ;
        RECT 4.54 12.752 4.572 12.784 ;
  LAYER M1 ;
        RECT 4.604 10.296 4.636 12.804 ;
  LAYER M3 ;
        RECT 4.604 10.316 4.636 10.348 ;
  LAYER M1 ;
        RECT 4.668 10.296 4.7 12.804 ;
  LAYER M3 ;
        RECT 4.668 12.752 4.7 12.784 ;
  LAYER M1 ;
        RECT 4.732 10.296 4.764 12.804 ;
  LAYER M3 ;
        RECT 4.732 10.316 4.764 10.348 ;
  LAYER M1 ;
        RECT 4.796 10.296 4.828 12.804 ;
  LAYER M3 ;
        RECT 4.796 12.752 4.828 12.784 ;
  LAYER M1 ;
        RECT 4.86 10.296 4.892 12.804 ;
  LAYER M3 ;
        RECT 4.86 10.316 4.892 10.348 ;
  LAYER M1 ;
        RECT 4.924 10.296 4.956 12.804 ;
  LAYER M3 ;
        RECT 4.924 12.752 4.956 12.784 ;
  LAYER M1 ;
        RECT 4.988 10.296 5.02 12.804 ;
  LAYER M3 ;
        RECT 4.988 10.316 5.02 10.348 ;
  LAYER M1 ;
        RECT 5.052 10.296 5.084 12.804 ;
  LAYER M3 ;
        RECT 5.052 12.752 5.084 12.784 ;
  LAYER M1 ;
        RECT 5.116 10.296 5.148 12.804 ;
  LAYER M3 ;
        RECT 5.116 10.316 5.148 10.348 ;
  LAYER M1 ;
        RECT 5.18 10.296 5.212 12.804 ;
  LAYER M3 ;
        RECT 5.18 12.752 5.212 12.784 ;
  LAYER M1 ;
        RECT 5.244 10.296 5.276 12.804 ;
  LAYER M3 ;
        RECT 5.244 10.316 5.276 10.348 ;
  LAYER M1 ;
        RECT 5.308 10.296 5.34 12.804 ;
  LAYER M3 ;
        RECT 5.308 12.752 5.34 12.784 ;
  LAYER M1 ;
        RECT 5.372 10.296 5.404 12.804 ;
  LAYER M3 ;
        RECT 5.372 10.316 5.404 10.348 ;
  LAYER M1 ;
        RECT 5.436 10.296 5.468 12.804 ;
  LAYER M3 ;
        RECT 5.436 12.752 5.468 12.784 ;
  LAYER M1 ;
        RECT 5.5 10.296 5.532 12.804 ;
  LAYER M3 ;
        RECT 5.5 10.316 5.532 10.348 ;
  LAYER M1 ;
        RECT 5.564 10.296 5.596 12.804 ;
  LAYER M3 ;
        RECT 5.564 12.752 5.596 12.784 ;
  LAYER M1 ;
        RECT 5.628 10.296 5.66 12.804 ;
  LAYER M3 ;
        RECT 5.628 10.316 5.66 10.348 ;
  LAYER M1 ;
        RECT 5.692 10.296 5.724 12.804 ;
  LAYER M3 ;
        RECT 5.692 12.752 5.724 12.784 ;
  LAYER M1 ;
        RECT 5.756 10.296 5.788 12.804 ;
  LAYER M3 ;
        RECT 3.388 10.38 3.42 10.412 ;
  LAYER M2 ;
        RECT 5.756 10.444 5.788 10.476 ;
  LAYER M2 ;
        RECT 3.388 10.508 3.42 10.54 ;
  LAYER M2 ;
        RECT 5.756 10.572 5.788 10.604 ;
  LAYER M2 ;
        RECT 3.388 10.636 3.42 10.668 ;
  LAYER M2 ;
        RECT 5.756 10.7 5.788 10.732 ;
  LAYER M2 ;
        RECT 3.388 10.764 3.42 10.796 ;
  LAYER M2 ;
        RECT 5.756 10.828 5.788 10.86 ;
  LAYER M2 ;
        RECT 3.388 10.892 3.42 10.924 ;
  LAYER M2 ;
        RECT 5.756 10.956 5.788 10.988 ;
  LAYER M2 ;
        RECT 3.388 11.02 3.42 11.052 ;
  LAYER M2 ;
        RECT 5.756 11.084 5.788 11.116 ;
  LAYER M2 ;
        RECT 3.388 11.148 3.42 11.18 ;
  LAYER M2 ;
        RECT 5.756 11.212 5.788 11.244 ;
  LAYER M2 ;
        RECT 3.388 11.276 3.42 11.308 ;
  LAYER M2 ;
        RECT 5.756 11.34 5.788 11.372 ;
  LAYER M2 ;
        RECT 3.388 11.404 3.42 11.436 ;
  LAYER M2 ;
        RECT 5.756 11.468 5.788 11.5 ;
  LAYER M2 ;
        RECT 3.388 11.532 3.42 11.564 ;
  LAYER M2 ;
        RECT 5.756 11.596 5.788 11.628 ;
  LAYER M2 ;
        RECT 3.388 11.66 3.42 11.692 ;
  LAYER M2 ;
        RECT 5.756 11.724 5.788 11.756 ;
  LAYER M2 ;
        RECT 3.388 11.788 3.42 11.82 ;
  LAYER M2 ;
        RECT 5.756 11.852 5.788 11.884 ;
  LAYER M2 ;
        RECT 3.388 11.916 3.42 11.948 ;
  LAYER M2 ;
        RECT 5.756 11.98 5.788 12.012 ;
  LAYER M2 ;
        RECT 3.388 12.044 3.42 12.076 ;
  LAYER M2 ;
        RECT 5.756 12.108 5.788 12.14 ;
  LAYER M2 ;
        RECT 3.388 12.172 3.42 12.204 ;
  LAYER M2 ;
        RECT 5.756 12.236 5.788 12.268 ;
  LAYER M2 ;
        RECT 3.388 12.3 3.42 12.332 ;
  LAYER M2 ;
        RECT 5.756 12.364 5.788 12.396 ;
  LAYER M2 ;
        RECT 3.388 12.428 3.42 12.46 ;
  LAYER M2 ;
        RECT 5.756 12.492 5.788 12.524 ;
  LAYER M2 ;
        RECT 3.388 12.556 3.42 12.588 ;
  LAYER M2 ;
        RECT 5.756 12.62 5.788 12.652 ;
  LAYER M2 ;
        RECT 3.34 10.248 5.836 12.852 ;
  LAYER M1 ;
        RECT 3.388 13.404 3.42 15.912 ;
  LAYER M3 ;
        RECT 3.388 15.86 3.42 15.892 ;
  LAYER M1 ;
        RECT 3.452 13.404 3.484 15.912 ;
  LAYER M3 ;
        RECT 3.452 13.424 3.484 13.456 ;
  LAYER M1 ;
        RECT 3.516 13.404 3.548 15.912 ;
  LAYER M3 ;
        RECT 3.516 15.86 3.548 15.892 ;
  LAYER M1 ;
        RECT 3.58 13.404 3.612 15.912 ;
  LAYER M3 ;
        RECT 3.58 13.424 3.612 13.456 ;
  LAYER M1 ;
        RECT 3.644 13.404 3.676 15.912 ;
  LAYER M3 ;
        RECT 3.644 15.86 3.676 15.892 ;
  LAYER M1 ;
        RECT 3.708 13.404 3.74 15.912 ;
  LAYER M3 ;
        RECT 3.708 13.424 3.74 13.456 ;
  LAYER M1 ;
        RECT 3.772 13.404 3.804 15.912 ;
  LAYER M3 ;
        RECT 3.772 15.86 3.804 15.892 ;
  LAYER M1 ;
        RECT 3.836 13.404 3.868 15.912 ;
  LAYER M3 ;
        RECT 3.836 13.424 3.868 13.456 ;
  LAYER M1 ;
        RECT 3.9 13.404 3.932 15.912 ;
  LAYER M3 ;
        RECT 3.9 15.86 3.932 15.892 ;
  LAYER M1 ;
        RECT 3.964 13.404 3.996 15.912 ;
  LAYER M3 ;
        RECT 3.964 13.424 3.996 13.456 ;
  LAYER M1 ;
        RECT 4.028 13.404 4.06 15.912 ;
  LAYER M3 ;
        RECT 4.028 15.86 4.06 15.892 ;
  LAYER M1 ;
        RECT 4.092 13.404 4.124 15.912 ;
  LAYER M3 ;
        RECT 4.092 13.424 4.124 13.456 ;
  LAYER M1 ;
        RECT 4.156 13.404 4.188 15.912 ;
  LAYER M3 ;
        RECT 4.156 15.86 4.188 15.892 ;
  LAYER M1 ;
        RECT 4.22 13.404 4.252 15.912 ;
  LAYER M3 ;
        RECT 4.22 13.424 4.252 13.456 ;
  LAYER M1 ;
        RECT 4.284 13.404 4.316 15.912 ;
  LAYER M3 ;
        RECT 4.284 15.86 4.316 15.892 ;
  LAYER M1 ;
        RECT 4.348 13.404 4.38 15.912 ;
  LAYER M3 ;
        RECT 4.348 13.424 4.38 13.456 ;
  LAYER M1 ;
        RECT 4.412 13.404 4.444 15.912 ;
  LAYER M3 ;
        RECT 4.412 15.86 4.444 15.892 ;
  LAYER M1 ;
        RECT 4.476 13.404 4.508 15.912 ;
  LAYER M3 ;
        RECT 4.476 13.424 4.508 13.456 ;
  LAYER M1 ;
        RECT 4.54 13.404 4.572 15.912 ;
  LAYER M3 ;
        RECT 4.54 15.86 4.572 15.892 ;
  LAYER M1 ;
        RECT 4.604 13.404 4.636 15.912 ;
  LAYER M3 ;
        RECT 4.604 13.424 4.636 13.456 ;
  LAYER M1 ;
        RECT 4.668 13.404 4.7 15.912 ;
  LAYER M3 ;
        RECT 4.668 15.86 4.7 15.892 ;
  LAYER M1 ;
        RECT 4.732 13.404 4.764 15.912 ;
  LAYER M3 ;
        RECT 4.732 13.424 4.764 13.456 ;
  LAYER M1 ;
        RECT 4.796 13.404 4.828 15.912 ;
  LAYER M3 ;
        RECT 4.796 15.86 4.828 15.892 ;
  LAYER M1 ;
        RECT 4.86 13.404 4.892 15.912 ;
  LAYER M3 ;
        RECT 4.86 13.424 4.892 13.456 ;
  LAYER M1 ;
        RECT 4.924 13.404 4.956 15.912 ;
  LAYER M3 ;
        RECT 4.924 15.86 4.956 15.892 ;
  LAYER M1 ;
        RECT 4.988 13.404 5.02 15.912 ;
  LAYER M3 ;
        RECT 4.988 13.424 5.02 13.456 ;
  LAYER M1 ;
        RECT 5.052 13.404 5.084 15.912 ;
  LAYER M3 ;
        RECT 5.052 15.86 5.084 15.892 ;
  LAYER M1 ;
        RECT 5.116 13.404 5.148 15.912 ;
  LAYER M3 ;
        RECT 5.116 13.424 5.148 13.456 ;
  LAYER M1 ;
        RECT 5.18 13.404 5.212 15.912 ;
  LAYER M3 ;
        RECT 5.18 15.86 5.212 15.892 ;
  LAYER M1 ;
        RECT 5.244 13.404 5.276 15.912 ;
  LAYER M3 ;
        RECT 5.244 13.424 5.276 13.456 ;
  LAYER M1 ;
        RECT 5.308 13.404 5.34 15.912 ;
  LAYER M3 ;
        RECT 5.308 15.86 5.34 15.892 ;
  LAYER M1 ;
        RECT 5.372 13.404 5.404 15.912 ;
  LAYER M3 ;
        RECT 5.372 13.424 5.404 13.456 ;
  LAYER M1 ;
        RECT 5.436 13.404 5.468 15.912 ;
  LAYER M3 ;
        RECT 5.436 15.86 5.468 15.892 ;
  LAYER M1 ;
        RECT 5.5 13.404 5.532 15.912 ;
  LAYER M3 ;
        RECT 5.5 13.424 5.532 13.456 ;
  LAYER M1 ;
        RECT 5.564 13.404 5.596 15.912 ;
  LAYER M3 ;
        RECT 5.564 15.86 5.596 15.892 ;
  LAYER M1 ;
        RECT 5.628 13.404 5.66 15.912 ;
  LAYER M3 ;
        RECT 5.628 13.424 5.66 13.456 ;
  LAYER M1 ;
        RECT 5.692 13.404 5.724 15.912 ;
  LAYER M3 ;
        RECT 5.692 15.86 5.724 15.892 ;
  LAYER M1 ;
        RECT 5.756 13.404 5.788 15.912 ;
  LAYER M3 ;
        RECT 3.388 13.488 3.42 13.52 ;
  LAYER M2 ;
        RECT 5.756 13.552 5.788 13.584 ;
  LAYER M2 ;
        RECT 3.388 13.616 3.42 13.648 ;
  LAYER M2 ;
        RECT 5.756 13.68 5.788 13.712 ;
  LAYER M2 ;
        RECT 3.388 13.744 3.42 13.776 ;
  LAYER M2 ;
        RECT 5.756 13.808 5.788 13.84 ;
  LAYER M2 ;
        RECT 3.388 13.872 3.42 13.904 ;
  LAYER M2 ;
        RECT 5.756 13.936 5.788 13.968 ;
  LAYER M2 ;
        RECT 3.388 14 3.42 14.032 ;
  LAYER M2 ;
        RECT 5.756 14.064 5.788 14.096 ;
  LAYER M2 ;
        RECT 3.388 14.128 3.42 14.16 ;
  LAYER M2 ;
        RECT 5.756 14.192 5.788 14.224 ;
  LAYER M2 ;
        RECT 3.388 14.256 3.42 14.288 ;
  LAYER M2 ;
        RECT 5.756 14.32 5.788 14.352 ;
  LAYER M2 ;
        RECT 3.388 14.384 3.42 14.416 ;
  LAYER M2 ;
        RECT 5.756 14.448 5.788 14.48 ;
  LAYER M2 ;
        RECT 3.388 14.512 3.42 14.544 ;
  LAYER M2 ;
        RECT 5.756 14.576 5.788 14.608 ;
  LAYER M2 ;
        RECT 3.388 14.64 3.42 14.672 ;
  LAYER M2 ;
        RECT 5.756 14.704 5.788 14.736 ;
  LAYER M2 ;
        RECT 3.388 14.768 3.42 14.8 ;
  LAYER M2 ;
        RECT 5.756 14.832 5.788 14.864 ;
  LAYER M2 ;
        RECT 3.388 14.896 3.42 14.928 ;
  LAYER M2 ;
        RECT 5.756 14.96 5.788 14.992 ;
  LAYER M2 ;
        RECT 3.388 15.024 3.42 15.056 ;
  LAYER M2 ;
        RECT 5.756 15.088 5.788 15.12 ;
  LAYER M2 ;
        RECT 3.388 15.152 3.42 15.184 ;
  LAYER M2 ;
        RECT 5.756 15.216 5.788 15.248 ;
  LAYER M2 ;
        RECT 3.388 15.28 3.42 15.312 ;
  LAYER M2 ;
        RECT 5.756 15.344 5.788 15.376 ;
  LAYER M2 ;
        RECT 3.388 15.408 3.42 15.44 ;
  LAYER M2 ;
        RECT 5.756 15.472 5.788 15.504 ;
  LAYER M2 ;
        RECT 3.388 15.536 3.42 15.568 ;
  LAYER M2 ;
        RECT 5.756 15.6 5.788 15.632 ;
  LAYER M2 ;
        RECT 3.388 15.664 3.42 15.696 ;
  LAYER M2 ;
        RECT 5.756 15.728 5.788 15.76 ;
  LAYER M2 ;
        RECT 3.34 13.356 5.836 15.96 ;
  LAYER M1 ;
        RECT 3.388 16.512 3.42 19.02 ;
  LAYER M3 ;
        RECT 3.388 18.968 3.42 19 ;
  LAYER M1 ;
        RECT 3.452 16.512 3.484 19.02 ;
  LAYER M3 ;
        RECT 3.452 16.532 3.484 16.564 ;
  LAYER M1 ;
        RECT 3.516 16.512 3.548 19.02 ;
  LAYER M3 ;
        RECT 3.516 18.968 3.548 19 ;
  LAYER M1 ;
        RECT 3.58 16.512 3.612 19.02 ;
  LAYER M3 ;
        RECT 3.58 16.532 3.612 16.564 ;
  LAYER M1 ;
        RECT 3.644 16.512 3.676 19.02 ;
  LAYER M3 ;
        RECT 3.644 18.968 3.676 19 ;
  LAYER M1 ;
        RECT 3.708 16.512 3.74 19.02 ;
  LAYER M3 ;
        RECT 3.708 16.532 3.74 16.564 ;
  LAYER M1 ;
        RECT 3.772 16.512 3.804 19.02 ;
  LAYER M3 ;
        RECT 3.772 18.968 3.804 19 ;
  LAYER M1 ;
        RECT 3.836 16.512 3.868 19.02 ;
  LAYER M3 ;
        RECT 3.836 16.532 3.868 16.564 ;
  LAYER M1 ;
        RECT 3.9 16.512 3.932 19.02 ;
  LAYER M3 ;
        RECT 3.9 18.968 3.932 19 ;
  LAYER M1 ;
        RECT 3.964 16.512 3.996 19.02 ;
  LAYER M3 ;
        RECT 3.964 16.532 3.996 16.564 ;
  LAYER M1 ;
        RECT 4.028 16.512 4.06 19.02 ;
  LAYER M3 ;
        RECT 4.028 18.968 4.06 19 ;
  LAYER M1 ;
        RECT 4.092 16.512 4.124 19.02 ;
  LAYER M3 ;
        RECT 4.092 16.532 4.124 16.564 ;
  LAYER M1 ;
        RECT 4.156 16.512 4.188 19.02 ;
  LAYER M3 ;
        RECT 4.156 18.968 4.188 19 ;
  LAYER M1 ;
        RECT 4.22 16.512 4.252 19.02 ;
  LAYER M3 ;
        RECT 4.22 16.532 4.252 16.564 ;
  LAYER M1 ;
        RECT 4.284 16.512 4.316 19.02 ;
  LAYER M3 ;
        RECT 4.284 18.968 4.316 19 ;
  LAYER M1 ;
        RECT 4.348 16.512 4.38 19.02 ;
  LAYER M3 ;
        RECT 4.348 16.532 4.38 16.564 ;
  LAYER M1 ;
        RECT 4.412 16.512 4.444 19.02 ;
  LAYER M3 ;
        RECT 4.412 18.968 4.444 19 ;
  LAYER M1 ;
        RECT 4.476 16.512 4.508 19.02 ;
  LAYER M3 ;
        RECT 4.476 16.532 4.508 16.564 ;
  LAYER M1 ;
        RECT 4.54 16.512 4.572 19.02 ;
  LAYER M3 ;
        RECT 4.54 18.968 4.572 19 ;
  LAYER M1 ;
        RECT 4.604 16.512 4.636 19.02 ;
  LAYER M3 ;
        RECT 4.604 16.532 4.636 16.564 ;
  LAYER M1 ;
        RECT 4.668 16.512 4.7 19.02 ;
  LAYER M3 ;
        RECT 4.668 18.968 4.7 19 ;
  LAYER M1 ;
        RECT 4.732 16.512 4.764 19.02 ;
  LAYER M3 ;
        RECT 4.732 16.532 4.764 16.564 ;
  LAYER M1 ;
        RECT 4.796 16.512 4.828 19.02 ;
  LAYER M3 ;
        RECT 4.796 18.968 4.828 19 ;
  LAYER M1 ;
        RECT 4.86 16.512 4.892 19.02 ;
  LAYER M3 ;
        RECT 4.86 16.532 4.892 16.564 ;
  LAYER M1 ;
        RECT 4.924 16.512 4.956 19.02 ;
  LAYER M3 ;
        RECT 4.924 18.968 4.956 19 ;
  LAYER M1 ;
        RECT 4.988 16.512 5.02 19.02 ;
  LAYER M3 ;
        RECT 4.988 16.532 5.02 16.564 ;
  LAYER M1 ;
        RECT 5.052 16.512 5.084 19.02 ;
  LAYER M3 ;
        RECT 5.052 18.968 5.084 19 ;
  LAYER M1 ;
        RECT 5.116 16.512 5.148 19.02 ;
  LAYER M3 ;
        RECT 5.116 16.532 5.148 16.564 ;
  LAYER M1 ;
        RECT 5.18 16.512 5.212 19.02 ;
  LAYER M3 ;
        RECT 5.18 18.968 5.212 19 ;
  LAYER M1 ;
        RECT 5.244 16.512 5.276 19.02 ;
  LAYER M3 ;
        RECT 5.244 16.532 5.276 16.564 ;
  LAYER M1 ;
        RECT 5.308 16.512 5.34 19.02 ;
  LAYER M3 ;
        RECT 5.308 18.968 5.34 19 ;
  LAYER M1 ;
        RECT 5.372 16.512 5.404 19.02 ;
  LAYER M3 ;
        RECT 5.372 16.532 5.404 16.564 ;
  LAYER M1 ;
        RECT 5.436 16.512 5.468 19.02 ;
  LAYER M3 ;
        RECT 5.436 18.968 5.468 19 ;
  LAYER M1 ;
        RECT 5.5 16.512 5.532 19.02 ;
  LAYER M3 ;
        RECT 5.5 16.532 5.532 16.564 ;
  LAYER M1 ;
        RECT 5.564 16.512 5.596 19.02 ;
  LAYER M3 ;
        RECT 5.564 18.968 5.596 19 ;
  LAYER M1 ;
        RECT 5.628 16.512 5.66 19.02 ;
  LAYER M3 ;
        RECT 5.628 16.532 5.66 16.564 ;
  LAYER M1 ;
        RECT 5.692 16.512 5.724 19.02 ;
  LAYER M3 ;
        RECT 5.692 18.968 5.724 19 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 19.02 ;
  LAYER M3 ;
        RECT 3.388 16.596 3.42 16.628 ;
  LAYER M2 ;
        RECT 5.756 16.66 5.788 16.692 ;
  LAYER M2 ;
        RECT 3.388 16.724 3.42 16.756 ;
  LAYER M2 ;
        RECT 5.756 16.788 5.788 16.82 ;
  LAYER M2 ;
        RECT 3.388 16.852 3.42 16.884 ;
  LAYER M2 ;
        RECT 5.756 16.916 5.788 16.948 ;
  LAYER M2 ;
        RECT 3.388 16.98 3.42 17.012 ;
  LAYER M2 ;
        RECT 5.756 17.044 5.788 17.076 ;
  LAYER M2 ;
        RECT 3.388 17.108 3.42 17.14 ;
  LAYER M2 ;
        RECT 5.756 17.172 5.788 17.204 ;
  LAYER M2 ;
        RECT 3.388 17.236 3.42 17.268 ;
  LAYER M2 ;
        RECT 5.756 17.3 5.788 17.332 ;
  LAYER M2 ;
        RECT 3.388 17.364 3.42 17.396 ;
  LAYER M2 ;
        RECT 5.756 17.428 5.788 17.46 ;
  LAYER M2 ;
        RECT 3.388 17.492 3.42 17.524 ;
  LAYER M2 ;
        RECT 5.756 17.556 5.788 17.588 ;
  LAYER M2 ;
        RECT 3.388 17.62 3.42 17.652 ;
  LAYER M2 ;
        RECT 5.756 17.684 5.788 17.716 ;
  LAYER M2 ;
        RECT 3.388 17.748 3.42 17.78 ;
  LAYER M2 ;
        RECT 5.756 17.812 5.788 17.844 ;
  LAYER M2 ;
        RECT 3.388 17.876 3.42 17.908 ;
  LAYER M2 ;
        RECT 5.756 17.94 5.788 17.972 ;
  LAYER M2 ;
        RECT 3.388 18.004 3.42 18.036 ;
  LAYER M2 ;
        RECT 5.756 18.068 5.788 18.1 ;
  LAYER M2 ;
        RECT 3.388 18.132 3.42 18.164 ;
  LAYER M2 ;
        RECT 5.756 18.196 5.788 18.228 ;
  LAYER M2 ;
        RECT 3.388 18.26 3.42 18.292 ;
  LAYER M2 ;
        RECT 5.756 18.324 5.788 18.356 ;
  LAYER M2 ;
        RECT 3.388 18.388 3.42 18.42 ;
  LAYER M2 ;
        RECT 5.756 18.452 5.788 18.484 ;
  LAYER M2 ;
        RECT 3.388 18.516 3.42 18.548 ;
  LAYER M2 ;
        RECT 5.756 18.58 5.788 18.612 ;
  LAYER M2 ;
        RECT 3.388 18.644 3.42 18.676 ;
  LAYER M2 ;
        RECT 5.756 18.708 5.788 18.74 ;
  LAYER M2 ;
        RECT 3.388 18.772 3.42 18.804 ;
  LAYER M2 ;
        RECT 5.756 18.836 5.788 18.868 ;
  LAYER M2 ;
        RECT 3.34 16.464 5.836 19.068 ;
  LAYER M1 ;
        RECT 3.388 19.62 3.42 22.128 ;
  LAYER M3 ;
        RECT 3.388 22.076 3.42 22.108 ;
  LAYER M1 ;
        RECT 3.452 19.62 3.484 22.128 ;
  LAYER M3 ;
        RECT 3.452 19.64 3.484 19.672 ;
  LAYER M1 ;
        RECT 3.516 19.62 3.548 22.128 ;
  LAYER M3 ;
        RECT 3.516 22.076 3.548 22.108 ;
  LAYER M1 ;
        RECT 3.58 19.62 3.612 22.128 ;
  LAYER M3 ;
        RECT 3.58 19.64 3.612 19.672 ;
  LAYER M1 ;
        RECT 3.644 19.62 3.676 22.128 ;
  LAYER M3 ;
        RECT 3.644 22.076 3.676 22.108 ;
  LAYER M1 ;
        RECT 3.708 19.62 3.74 22.128 ;
  LAYER M3 ;
        RECT 3.708 19.64 3.74 19.672 ;
  LAYER M1 ;
        RECT 3.772 19.62 3.804 22.128 ;
  LAYER M3 ;
        RECT 3.772 22.076 3.804 22.108 ;
  LAYER M1 ;
        RECT 3.836 19.62 3.868 22.128 ;
  LAYER M3 ;
        RECT 3.836 19.64 3.868 19.672 ;
  LAYER M1 ;
        RECT 3.9 19.62 3.932 22.128 ;
  LAYER M3 ;
        RECT 3.9 22.076 3.932 22.108 ;
  LAYER M1 ;
        RECT 3.964 19.62 3.996 22.128 ;
  LAYER M3 ;
        RECT 3.964 19.64 3.996 19.672 ;
  LAYER M1 ;
        RECT 4.028 19.62 4.06 22.128 ;
  LAYER M3 ;
        RECT 4.028 22.076 4.06 22.108 ;
  LAYER M1 ;
        RECT 4.092 19.62 4.124 22.128 ;
  LAYER M3 ;
        RECT 4.092 19.64 4.124 19.672 ;
  LAYER M1 ;
        RECT 4.156 19.62 4.188 22.128 ;
  LAYER M3 ;
        RECT 4.156 22.076 4.188 22.108 ;
  LAYER M1 ;
        RECT 4.22 19.62 4.252 22.128 ;
  LAYER M3 ;
        RECT 4.22 19.64 4.252 19.672 ;
  LAYER M1 ;
        RECT 4.284 19.62 4.316 22.128 ;
  LAYER M3 ;
        RECT 4.284 22.076 4.316 22.108 ;
  LAYER M1 ;
        RECT 4.348 19.62 4.38 22.128 ;
  LAYER M3 ;
        RECT 4.348 19.64 4.38 19.672 ;
  LAYER M1 ;
        RECT 4.412 19.62 4.444 22.128 ;
  LAYER M3 ;
        RECT 4.412 22.076 4.444 22.108 ;
  LAYER M1 ;
        RECT 4.476 19.62 4.508 22.128 ;
  LAYER M3 ;
        RECT 4.476 19.64 4.508 19.672 ;
  LAYER M1 ;
        RECT 4.54 19.62 4.572 22.128 ;
  LAYER M3 ;
        RECT 4.54 22.076 4.572 22.108 ;
  LAYER M1 ;
        RECT 4.604 19.62 4.636 22.128 ;
  LAYER M3 ;
        RECT 4.604 19.64 4.636 19.672 ;
  LAYER M1 ;
        RECT 4.668 19.62 4.7 22.128 ;
  LAYER M3 ;
        RECT 4.668 22.076 4.7 22.108 ;
  LAYER M1 ;
        RECT 4.732 19.62 4.764 22.128 ;
  LAYER M3 ;
        RECT 4.732 19.64 4.764 19.672 ;
  LAYER M1 ;
        RECT 4.796 19.62 4.828 22.128 ;
  LAYER M3 ;
        RECT 4.796 22.076 4.828 22.108 ;
  LAYER M1 ;
        RECT 4.86 19.62 4.892 22.128 ;
  LAYER M3 ;
        RECT 4.86 19.64 4.892 19.672 ;
  LAYER M1 ;
        RECT 4.924 19.62 4.956 22.128 ;
  LAYER M3 ;
        RECT 4.924 22.076 4.956 22.108 ;
  LAYER M1 ;
        RECT 4.988 19.62 5.02 22.128 ;
  LAYER M3 ;
        RECT 4.988 19.64 5.02 19.672 ;
  LAYER M1 ;
        RECT 5.052 19.62 5.084 22.128 ;
  LAYER M3 ;
        RECT 5.052 22.076 5.084 22.108 ;
  LAYER M1 ;
        RECT 5.116 19.62 5.148 22.128 ;
  LAYER M3 ;
        RECT 5.116 19.64 5.148 19.672 ;
  LAYER M1 ;
        RECT 5.18 19.62 5.212 22.128 ;
  LAYER M3 ;
        RECT 5.18 22.076 5.212 22.108 ;
  LAYER M1 ;
        RECT 5.244 19.62 5.276 22.128 ;
  LAYER M3 ;
        RECT 5.244 19.64 5.276 19.672 ;
  LAYER M1 ;
        RECT 5.308 19.62 5.34 22.128 ;
  LAYER M3 ;
        RECT 5.308 22.076 5.34 22.108 ;
  LAYER M1 ;
        RECT 5.372 19.62 5.404 22.128 ;
  LAYER M3 ;
        RECT 5.372 19.64 5.404 19.672 ;
  LAYER M1 ;
        RECT 5.436 19.62 5.468 22.128 ;
  LAYER M3 ;
        RECT 5.436 22.076 5.468 22.108 ;
  LAYER M1 ;
        RECT 5.5 19.62 5.532 22.128 ;
  LAYER M3 ;
        RECT 5.5 19.64 5.532 19.672 ;
  LAYER M1 ;
        RECT 5.564 19.62 5.596 22.128 ;
  LAYER M3 ;
        RECT 5.564 22.076 5.596 22.108 ;
  LAYER M1 ;
        RECT 5.628 19.62 5.66 22.128 ;
  LAYER M3 ;
        RECT 5.628 19.64 5.66 19.672 ;
  LAYER M1 ;
        RECT 5.692 19.62 5.724 22.128 ;
  LAYER M3 ;
        RECT 5.692 22.076 5.724 22.108 ;
  LAYER M1 ;
        RECT 5.756 19.62 5.788 22.128 ;
  LAYER M3 ;
        RECT 3.388 19.704 3.42 19.736 ;
  LAYER M2 ;
        RECT 5.756 19.768 5.788 19.8 ;
  LAYER M2 ;
        RECT 3.388 19.832 3.42 19.864 ;
  LAYER M2 ;
        RECT 5.756 19.896 5.788 19.928 ;
  LAYER M2 ;
        RECT 3.388 19.96 3.42 19.992 ;
  LAYER M2 ;
        RECT 5.756 20.024 5.788 20.056 ;
  LAYER M2 ;
        RECT 3.388 20.088 3.42 20.12 ;
  LAYER M2 ;
        RECT 5.756 20.152 5.788 20.184 ;
  LAYER M2 ;
        RECT 3.388 20.216 3.42 20.248 ;
  LAYER M2 ;
        RECT 5.756 20.28 5.788 20.312 ;
  LAYER M2 ;
        RECT 3.388 20.344 3.42 20.376 ;
  LAYER M2 ;
        RECT 5.756 20.408 5.788 20.44 ;
  LAYER M2 ;
        RECT 3.388 20.472 3.42 20.504 ;
  LAYER M2 ;
        RECT 5.756 20.536 5.788 20.568 ;
  LAYER M2 ;
        RECT 3.388 20.6 3.42 20.632 ;
  LAYER M2 ;
        RECT 5.756 20.664 5.788 20.696 ;
  LAYER M2 ;
        RECT 3.388 20.728 3.42 20.76 ;
  LAYER M2 ;
        RECT 5.756 20.792 5.788 20.824 ;
  LAYER M2 ;
        RECT 3.388 20.856 3.42 20.888 ;
  LAYER M2 ;
        RECT 5.756 20.92 5.788 20.952 ;
  LAYER M2 ;
        RECT 3.388 20.984 3.42 21.016 ;
  LAYER M2 ;
        RECT 5.756 21.048 5.788 21.08 ;
  LAYER M2 ;
        RECT 3.388 21.112 3.42 21.144 ;
  LAYER M2 ;
        RECT 5.756 21.176 5.788 21.208 ;
  LAYER M2 ;
        RECT 3.388 21.24 3.42 21.272 ;
  LAYER M2 ;
        RECT 5.756 21.304 5.788 21.336 ;
  LAYER M2 ;
        RECT 3.388 21.368 3.42 21.4 ;
  LAYER M2 ;
        RECT 5.756 21.432 5.788 21.464 ;
  LAYER M2 ;
        RECT 3.388 21.496 3.42 21.528 ;
  LAYER M2 ;
        RECT 5.756 21.56 5.788 21.592 ;
  LAYER M2 ;
        RECT 3.388 21.624 3.42 21.656 ;
  LAYER M2 ;
        RECT 5.756 21.688 5.788 21.72 ;
  LAYER M2 ;
        RECT 3.388 21.752 3.42 21.784 ;
  LAYER M2 ;
        RECT 5.756 21.816 5.788 21.848 ;
  LAYER M2 ;
        RECT 3.388 21.88 3.42 21.912 ;
  LAYER M2 ;
        RECT 5.756 21.944 5.788 21.976 ;
  LAYER M2 ;
        RECT 3.34 19.572 5.836 22.176 ;
  LAYER M1 ;
        RECT 6.684 0.972 6.716 3.48 ;
  LAYER M3 ;
        RECT 6.684 3.428 6.716 3.46 ;
  LAYER M1 ;
        RECT 6.748 0.972 6.78 3.48 ;
  LAYER M3 ;
        RECT 6.748 0.992 6.78 1.024 ;
  LAYER M1 ;
        RECT 6.812 0.972 6.844 3.48 ;
  LAYER M3 ;
        RECT 6.812 3.428 6.844 3.46 ;
  LAYER M1 ;
        RECT 6.876 0.972 6.908 3.48 ;
  LAYER M3 ;
        RECT 6.876 0.992 6.908 1.024 ;
  LAYER M1 ;
        RECT 6.94 0.972 6.972 3.48 ;
  LAYER M3 ;
        RECT 6.94 3.428 6.972 3.46 ;
  LAYER M1 ;
        RECT 7.004 0.972 7.036 3.48 ;
  LAYER M3 ;
        RECT 7.004 0.992 7.036 1.024 ;
  LAYER M1 ;
        RECT 7.068 0.972 7.1 3.48 ;
  LAYER M3 ;
        RECT 7.068 3.428 7.1 3.46 ;
  LAYER M1 ;
        RECT 7.132 0.972 7.164 3.48 ;
  LAYER M3 ;
        RECT 7.132 0.992 7.164 1.024 ;
  LAYER M1 ;
        RECT 7.196 0.972 7.228 3.48 ;
  LAYER M3 ;
        RECT 7.196 3.428 7.228 3.46 ;
  LAYER M1 ;
        RECT 7.26 0.972 7.292 3.48 ;
  LAYER M3 ;
        RECT 7.26 0.992 7.292 1.024 ;
  LAYER M1 ;
        RECT 7.324 0.972 7.356 3.48 ;
  LAYER M3 ;
        RECT 7.324 3.428 7.356 3.46 ;
  LAYER M1 ;
        RECT 7.388 0.972 7.42 3.48 ;
  LAYER M3 ;
        RECT 7.388 0.992 7.42 1.024 ;
  LAYER M1 ;
        RECT 7.452 0.972 7.484 3.48 ;
  LAYER M3 ;
        RECT 7.452 3.428 7.484 3.46 ;
  LAYER M1 ;
        RECT 7.516 0.972 7.548 3.48 ;
  LAYER M3 ;
        RECT 7.516 0.992 7.548 1.024 ;
  LAYER M1 ;
        RECT 7.58 0.972 7.612 3.48 ;
  LAYER M3 ;
        RECT 7.58 3.428 7.612 3.46 ;
  LAYER M1 ;
        RECT 7.644 0.972 7.676 3.48 ;
  LAYER M3 ;
        RECT 7.644 0.992 7.676 1.024 ;
  LAYER M1 ;
        RECT 7.708 0.972 7.74 3.48 ;
  LAYER M3 ;
        RECT 7.708 3.428 7.74 3.46 ;
  LAYER M1 ;
        RECT 7.772 0.972 7.804 3.48 ;
  LAYER M3 ;
        RECT 7.772 0.992 7.804 1.024 ;
  LAYER M1 ;
        RECT 7.836 0.972 7.868 3.48 ;
  LAYER M3 ;
        RECT 7.836 3.428 7.868 3.46 ;
  LAYER M1 ;
        RECT 7.9 0.972 7.932 3.48 ;
  LAYER M3 ;
        RECT 7.9 0.992 7.932 1.024 ;
  LAYER M1 ;
        RECT 7.964 0.972 7.996 3.48 ;
  LAYER M3 ;
        RECT 7.964 3.428 7.996 3.46 ;
  LAYER M1 ;
        RECT 8.028 0.972 8.06 3.48 ;
  LAYER M3 ;
        RECT 8.028 0.992 8.06 1.024 ;
  LAYER M1 ;
        RECT 8.092 0.972 8.124 3.48 ;
  LAYER M3 ;
        RECT 8.092 3.428 8.124 3.46 ;
  LAYER M1 ;
        RECT 8.156 0.972 8.188 3.48 ;
  LAYER M3 ;
        RECT 8.156 0.992 8.188 1.024 ;
  LAYER M1 ;
        RECT 8.22 0.972 8.252 3.48 ;
  LAYER M3 ;
        RECT 8.22 3.428 8.252 3.46 ;
  LAYER M1 ;
        RECT 8.284 0.972 8.316 3.48 ;
  LAYER M3 ;
        RECT 8.284 0.992 8.316 1.024 ;
  LAYER M1 ;
        RECT 8.348 0.972 8.38 3.48 ;
  LAYER M3 ;
        RECT 8.348 3.428 8.38 3.46 ;
  LAYER M1 ;
        RECT 8.412 0.972 8.444 3.48 ;
  LAYER M3 ;
        RECT 8.412 0.992 8.444 1.024 ;
  LAYER M1 ;
        RECT 8.476 0.972 8.508 3.48 ;
  LAYER M3 ;
        RECT 8.476 3.428 8.508 3.46 ;
  LAYER M1 ;
        RECT 8.54 0.972 8.572 3.48 ;
  LAYER M3 ;
        RECT 8.54 0.992 8.572 1.024 ;
  LAYER M1 ;
        RECT 8.604 0.972 8.636 3.48 ;
  LAYER M3 ;
        RECT 8.604 3.428 8.636 3.46 ;
  LAYER M1 ;
        RECT 8.668 0.972 8.7 3.48 ;
  LAYER M3 ;
        RECT 8.668 0.992 8.7 1.024 ;
  LAYER M1 ;
        RECT 8.732 0.972 8.764 3.48 ;
  LAYER M3 ;
        RECT 8.732 3.428 8.764 3.46 ;
  LAYER M1 ;
        RECT 8.796 0.972 8.828 3.48 ;
  LAYER M3 ;
        RECT 8.796 0.992 8.828 1.024 ;
  LAYER M1 ;
        RECT 8.86 0.972 8.892 3.48 ;
  LAYER M3 ;
        RECT 8.86 3.428 8.892 3.46 ;
  LAYER M1 ;
        RECT 8.924 0.972 8.956 3.48 ;
  LAYER M3 ;
        RECT 8.924 0.992 8.956 1.024 ;
  LAYER M1 ;
        RECT 8.988 0.972 9.02 3.48 ;
  LAYER M3 ;
        RECT 8.988 3.428 9.02 3.46 ;
  LAYER M1 ;
        RECT 9.052 0.972 9.084 3.48 ;
  LAYER M3 ;
        RECT 6.684 1.056 6.716 1.088 ;
  LAYER M2 ;
        RECT 9.052 1.12 9.084 1.152 ;
  LAYER M2 ;
        RECT 6.684 1.184 6.716 1.216 ;
  LAYER M2 ;
        RECT 9.052 1.248 9.084 1.28 ;
  LAYER M2 ;
        RECT 6.684 1.312 6.716 1.344 ;
  LAYER M2 ;
        RECT 9.052 1.376 9.084 1.408 ;
  LAYER M2 ;
        RECT 6.684 1.44 6.716 1.472 ;
  LAYER M2 ;
        RECT 9.052 1.504 9.084 1.536 ;
  LAYER M2 ;
        RECT 6.684 1.568 6.716 1.6 ;
  LAYER M2 ;
        RECT 9.052 1.632 9.084 1.664 ;
  LAYER M2 ;
        RECT 6.684 1.696 6.716 1.728 ;
  LAYER M2 ;
        RECT 9.052 1.76 9.084 1.792 ;
  LAYER M2 ;
        RECT 6.684 1.824 6.716 1.856 ;
  LAYER M2 ;
        RECT 9.052 1.888 9.084 1.92 ;
  LAYER M2 ;
        RECT 6.684 1.952 6.716 1.984 ;
  LAYER M2 ;
        RECT 9.052 2.016 9.084 2.048 ;
  LAYER M2 ;
        RECT 6.684 2.08 6.716 2.112 ;
  LAYER M2 ;
        RECT 9.052 2.144 9.084 2.176 ;
  LAYER M2 ;
        RECT 6.684 2.208 6.716 2.24 ;
  LAYER M2 ;
        RECT 9.052 2.272 9.084 2.304 ;
  LAYER M2 ;
        RECT 6.684 2.336 6.716 2.368 ;
  LAYER M2 ;
        RECT 9.052 2.4 9.084 2.432 ;
  LAYER M2 ;
        RECT 6.684 2.464 6.716 2.496 ;
  LAYER M2 ;
        RECT 9.052 2.528 9.084 2.56 ;
  LAYER M2 ;
        RECT 6.684 2.592 6.716 2.624 ;
  LAYER M2 ;
        RECT 9.052 2.656 9.084 2.688 ;
  LAYER M2 ;
        RECT 6.684 2.72 6.716 2.752 ;
  LAYER M2 ;
        RECT 9.052 2.784 9.084 2.816 ;
  LAYER M2 ;
        RECT 6.684 2.848 6.716 2.88 ;
  LAYER M2 ;
        RECT 9.052 2.912 9.084 2.944 ;
  LAYER M2 ;
        RECT 6.684 2.976 6.716 3.008 ;
  LAYER M2 ;
        RECT 9.052 3.04 9.084 3.072 ;
  LAYER M2 ;
        RECT 6.684 3.104 6.716 3.136 ;
  LAYER M2 ;
        RECT 9.052 3.168 9.084 3.2 ;
  LAYER M2 ;
        RECT 6.684 3.232 6.716 3.264 ;
  LAYER M2 ;
        RECT 9.052 3.296 9.084 3.328 ;
  LAYER M2 ;
        RECT 6.636 0.924 9.132 3.528 ;
  LAYER M1 ;
        RECT 6.684 4.08 6.716 6.588 ;
  LAYER M3 ;
        RECT 6.684 6.536 6.716 6.568 ;
  LAYER M1 ;
        RECT 6.748 4.08 6.78 6.588 ;
  LAYER M3 ;
        RECT 6.748 4.1 6.78 4.132 ;
  LAYER M1 ;
        RECT 6.812 4.08 6.844 6.588 ;
  LAYER M3 ;
        RECT 6.812 6.536 6.844 6.568 ;
  LAYER M1 ;
        RECT 6.876 4.08 6.908 6.588 ;
  LAYER M3 ;
        RECT 6.876 4.1 6.908 4.132 ;
  LAYER M1 ;
        RECT 6.94 4.08 6.972 6.588 ;
  LAYER M3 ;
        RECT 6.94 6.536 6.972 6.568 ;
  LAYER M1 ;
        RECT 7.004 4.08 7.036 6.588 ;
  LAYER M3 ;
        RECT 7.004 4.1 7.036 4.132 ;
  LAYER M1 ;
        RECT 7.068 4.08 7.1 6.588 ;
  LAYER M3 ;
        RECT 7.068 6.536 7.1 6.568 ;
  LAYER M1 ;
        RECT 7.132 4.08 7.164 6.588 ;
  LAYER M3 ;
        RECT 7.132 4.1 7.164 4.132 ;
  LAYER M1 ;
        RECT 7.196 4.08 7.228 6.588 ;
  LAYER M3 ;
        RECT 7.196 6.536 7.228 6.568 ;
  LAYER M1 ;
        RECT 7.26 4.08 7.292 6.588 ;
  LAYER M3 ;
        RECT 7.26 4.1 7.292 4.132 ;
  LAYER M1 ;
        RECT 7.324 4.08 7.356 6.588 ;
  LAYER M3 ;
        RECT 7.324 6.536 7.356 6.568 ;
  LAYER M1 ;
        RECT 7.388 4.08 7.42 6.588 ;
  LAYER M3 ;
        RECT 7.388 4.1 7.42 4.132 ;
  LAYER M1 ;
        RECT 7.452 4.08 7.484 6.588 ;
  LAYER M3 ;
        RECT 7.452 6.536 7.484 6.568 ;
  LAYER M1 ;
        RECT 7.516 4.08 7.548 6.588 ;
  LAYER M3 ;
        RECT 7.516 4.1 7.548 4.132 ;
  LAYER M1 ;
        RECT 7.58 4.08 7.612 6.588 ;
  LAYER M3 ;
        RECT 7.58 6.536 7.612 6.568 ;
  LAYER M1 ;
        RECT 7.644 4.08 7.676 6.588 ;
  LAYER M3 ;
        RECT 7.644 4.1 7.676 4.132 ;
  LAYER M1 ;
        RECT 7.708 4.08 7.74 6.588 ;
  LAYER M3 ;
        RECT 7.708 6.536 7.74 6.568 ;
  LAYER M1 ;
        RECT 7.772 4.08 7.804 6.588 ;
  LAYER M3 ;
        RECT 7.772 4.1 7.804 4.132 ;
  LAYER M1 ;
        RECT 7.836 4.08 7.868 6.588 ;
  LAYER M3 ;
        RECT 7.836 6.536 7.868 6.568 ;
  LAYER M1 ;
        RECT 7.9 4.08 7.932 6.588 ;
  LAYER M3 ;
        RECT 7.9 4.1 7.932 4.132 ;
  LAYER M1 ;
        RECT 7.964 4.08 7.996 6.588 ;
  LAYER M3 ;
        RECT 7.964 6.536 7.996 6.568 ;
  LAYER M1 ;
        RECT 8.028 4.08 8.06 6.588 ;
  LAYER M3 ;
        RECT 8.028 4.1 8.06 4.132 ;
  LAYER M1 ;
        RECT 8.092 4.08 8.124 6.588 ;
  LAYER M3 ;
        RECT 8.092 6.536 8.124 6.568 ;
  LAYER M1 ;
        RECT 8.156 4.08 8.188 6.588 ;
  LAYER M3 ;
        RECT 8.156 4.1 8.188 4.132 ;
  LAYER M1 ;
        RECT 8.22 4.08 8.252 6.588 ;
  LAYER M3 ;
        RECT 8.22 6.536 8.252 6.568 ;
  LAYER M1 ;
        RECT 8.284 4.08 8.316 6.588 ;
  LAYER M3 ;
        RECT 8.284 4.1 8.316 4.132 ;
  LAYER M1 ;
        RECT 8.348 4.08 8.38 6.588 ;
  LAYER M3 ;
        RECT 8.348 6.536 8.38 6.568 ;
  LAYER M1 ;
        RECT 8.412 4.08 8.444 6.588 ;
  LAYER M3 ;
        RECT 8.412 4.1 8.444 4.132 ;
  LAYER M1 ;
        RECT 8.476 4.08 8.508 6.588 ;
  LAYER M3 ;
        RECT 8.476 6.536 8.508 6.568 ;
  LAYER M1 ;
        RECT 8.54 4.08 8.572 6.588 ;
  LAYER M3 ;
        RECT 8.54 4.1 8.572 4.132 ;
  LAYER M1 ;
        RECT 8.604 4.08 8.636 6.588 ;
  LAYER M3 ;
        RECT 8.604 6.536 8.636 6.568 ;
  LAYER M1 ;
        RECT 8.668 4.08 8.7 6.588 ;
  LAYER M3 ;
        RECT 8.668 4.1 8.7 4.132 ;
  LAYER M1 ;
        RECT 8.732 4.08 8.764 6.588 ;
  LAYER M3 ;
        RECT 8.732 6.536 8.764 6.568 ;
  LAYER M1 ;
        RECT 8.796 4.08 8.828 6.588 ;
  LAYER M3 ;
        RECT 8.796 4.1 8.828 4.132 ;
  LAYER M1 ;
        RECT 8.86 4.08 8.892 6.588 ;
  LAYER M3 ;
        RECT 8.86 6.536 8.892 6.568 ;
  LAYER M1 ;
        RECT 8.924 4.08 8.956 6.588 ;
  LAYER M3 ;
        RECT 8.924 4.1 8.956 4.132 ;
  LAYER M1 ;
        RECT 8.988 4.08 9.02 6.588 ;
  LAYER M3 ;
        RECT 8.988 6.536 9.02 6.568 ;
  LAYER M1 ;
        RECT 9.052 4.08 9.084 6.588 ;
  LAYER M3 ;
        RECT 6.684 4.164 6.716 4.196 ;
  LAYER M2 ;
        RECT 9.052 4.228 9.084 4.26 ;
  LAYER M2 ;
        RECT 6.684 4.292 6.716 4.324 ;
  LAYER M2 ;
        RECT 9.052 4.356 9.084 4.388 ;
  LAYER M2 ;
        RECT 6.684 4.42 6.716 4.452 ;
  LAYER M2 ;
        RECT 9.052 4.484 9.084 4.516 ;
  LAYER M2 ;
        RECT 6.684 4.548 6.716 4.58 ;
  LAYER M2 ;
        RECT 9.052 4.612 9.084 4.644 ;
  LAYER M2 ;
        RECT 6.684 4.676 6.716 4.708 ;
  LAYER M2 ;
        RECT 9.052 4.74 9.084 4.772 ;
  LAYER M2 ;
        RECT 6.684 4.804 6.716 4.836 ;
  LAYER M2 ;
        RECT 9.052 4.868 9.084 4.9 ;
  LAYER M2 ;
        RECT 6.684 4.932 6.716 4.964 ;
  LAYER M2 ;
        RECT 9.052 4.996 9.084 5.028 ;
  LAYER M2 ;
        RECT 6.684 5.06 6.716 5.092 ;
  LAYER M2 ;
        RECT 9.052 5.124 9.084 5.156 ;
  LAYER M2 ;
        RECT 6.684 5.188 6.716 5.22 ;
  LAYER M2 ;
        RECT 9.052 5.252 9.084 5.284 ;
  LAYER M2 ;
        RECT 6.684 5.316 6.716 5.348 ;
  LAYER M2 ;
        RECT 9.052 5.38 9.084 5.412 ;
  LAYER M2 ;
        RECT 6.684 5.444 6.716 5.476 ;
  LAYER M2 ;
        RECT 9.052 5.508 9.084 5.54 ;
  LAYER M2 ;
        RECT 6.684 5.572 6.716 5.604 ;
  LAYER M2 ;
        RECT 9.052 5.636 9.084 5.668 ;
  LAYER M2 ;
        RECT 6.684 5.7 6.716 5.732 ;
  LAYER M2 ;
        RECT 9.052 5.764 9.084 5.796 ;
  LAYER M2 ;
        RECT 6.684 5.828 6.716 5.86 ;
  LAYER M2 ;
        RECT 9.052 5.892 9.084 5.924 ;
  LAYER M2 ;
        RECT 6.684 5.956 6.716 5.988 ;
  LAYER M2 ;
        RECT 9.052 6.02 9.084 6.052 ;
  LAYER M2 ;
        RECT 6.684 6.084 6.716 6.116 ;
  LAYER M2 ;
        RECT 9.052 6.148 9.084 6.18 ;
  LAYER M2 ;
        RECT 6.684 6.212 6.716 6.244 ;
  LAYER M2 ;
        RECT 9.052 6.276 9.084 6.308 ;
  LAYER M2 ;
        RECT 6.684 6.34 6.716 6.372 ;
  LAYER M2 ;
        RECT 9.052 6.404 9.084 6.436 ;
  LAYER M2 ;
        RECT 6.636 4.032 9.132 6.636 ;
  LAYER M1 ;
        RECT 6.684 7.188 6.716 9.696 ;
  LAYER M3 ;
        RECT 6.684 9.644 6.716 9.676 ;
  LAYER M1 ;
        RECT 6.748 7.188 6.78 9.696 ;
  LAYER M3 ;
        RECT 6.748 7.208 6.78 7.24 ;
  LAYER M1 ;
        RECT 6.812 7.188 6.844 9.696 ;
  LAYER M3 ;
        RECT 6.812 9.644 6.844 9.676 ;
  LAYER M1 ;
        RECT 6.876 7.188 6.908 9.696 ;
  LAYER M3 ;
        RECT 6.876 7.208 6.908 7.24 ;
  LAYER M1 ;
        RECT 6.94 7.188 6.972 9.696 ;
  LAYER M3 ;
        RECT 6.94 9.644 6.972 9.676 ;
  LAYER M1 ;
        RECT 7.004 7.188 7.036 9.696 ;
  LAYER M3 ;
        RECT 7.004 7.208 7.036 7.24 ;
  LAYER M1 ;
        RECT 7.068 7.188 7.1 9.696 ;
  LAYER M3 ;
        RECT 7.068 9.644 7.1 9.676 ;
  LAYER M1 ;
        RECT 7.132 7.188 7.164 9.696 ;
  LAYER M3 ;
        RECT 7.132 7.208 7.164 7.24 ;
  LAYER M1 ;
        RECT 7.196 7.188 7.228 9.696 ;
  LAYER M3 ;
        RECT 7.196 9.644 7.228 9.676 ;
  LAYER M1 ;
        RECT 7.26 7.188 7.292 9.696 ;
  LAYER M3 ;
        RECT 7.26 7.208 7.292 7.24 ;
  LAYER M1 ;
        RECT 7.324 7.188 7.356 9.696 ;
  LAYER M3 ;
        RECT 7.324 9.644 7.356 9.676 ;
  LAYER M1 ;
        RECT 7.388 7.188 7.42 9.696 ;
  LAYER M3 ;
        RECT 7.388 7.208 7.42 7.24 ;
  LAYER M1 ;
        RECT 7.452 7.188 7.484 9.696 ;
  LAYER M3 ;
        RECT 7.452 9.644 7.484 9.676 ;
  LAYER M1 ;
        RECT 7.516 7.188 7.548 9.696 ;
  LAYER M3 ;
        RECT 7.516 7.208 7.548 7.24 ;
  LAYER M1 ;
        RECT 7.58 7.188 7.612 9.696 ;
  LAYER M3 ;
        RECT 7.58 9.644 7.612 9.676 ;
  LAYER M1 ;
        RECT 7.644 7.188 7.676 9.696 ;
  LAYER M3 ;
        RECT 7.644 7.208 7.676 7.24 ;
  LAYER M1 ;
        RECT 7.708 7.188 7.74 9.696 ;
  LAYER M3 ;
        RECT 7.708 9.644 7.74 9.676 ;
  LAYER M1 ;
        RECT 7.772 7.188 7.804 9.696 ;
  LAYER M3 ;
        RECT 7.772 7.208 7.804 7.24 ;
  LAYER M1 ;
        RECT 7.836 7.188 7.868 9.696 ;
  LAYER M3 ;
        RECT 7.836 9.644 7.868 9.676 ;
  LAYER M1 ;
        RECT 7.9 7.188 7.932 9.696 ;
  LAYER M3 ;
        RECT 7.9 7.208 7.932 7.24 ;
  LAYER M1 ;
        RECT 7.964 7.188 7.996 9.696 ;
  LAYER M3 ;
        RECT 7.964 9.644 7.996 9.676 ;
  LAYER M1 ;
        RECT 8.028 7.188 8.06 9.696 ;
  LAYER M3 ;
        RECT 8.028 7.208 8.06 7.24 ;
  LAYER M1 ;
        RECT 8.092 7.188 8.124 9.696 ;
  LAYER M3 ;
        RECT 8.092 9.644 8.124 9.676 ;
  LAYER M1 ;
        RECT 8.156 7.188 8.188 9.696 ;
  LAYER M3 ;
        RECT 8.156 7.208 8.188 7.24 ;
  LAYER M1 ;
        RECT 8.22 7.188 8.252 9.696 ;
  LAYER M3 ;
        RECT 8.22 9.644 8.252 9.676 ;
  LAYER M1 ;
        RECT 8.284 7.188 8.316 9.696 ;
  LAYER M3 ;
        RECT 8.284 7.208 8.316 7.24 ;
  LAYER M1 ;
        RECT 8.348 7.188 8.38 9.696 ;
  LAYER M3 ;
        RECT 8.348 9.644 8.38 9.676 ;
  LAYER M1 ;
        RECT 8.412 7.188 8.444 9.696 ;
  LAYER M3 ;
        RECT 8.412 7.208 8.444 7.24 ;
  LAYER M1 ;
        RECT 8.476 7.188 8.508 9.696 ;
  LAYER M3 ;
        RECT 8.476 9.644 8.508 9.676 ;
  LAYER M1 ;
        RECT 8.54 7.188 8.572 9.696 ;
  LAYER M3 ;
        RECT 8.54 7.208 8.572 7.24 ;
  LAYER M1 ;
        RECT 8.604 7.188 8.636 9.696 ;
  LAYER M3 ;
        RECT 8.604 9.644 8.636 9.676 ;
  LAYER M1 ;
        RECT 8.668 7.188 8.7 9.696 ;
  LAYER M3 ;
        RECT 8.668 7.208 8.7 7.24 ;
  LAYER M1 ;
        RECT 8.732 7.188 8.764 9.696 ;
  LAYER M3 ;
        RECT 8.732 9.644 8.764 9.676 ;
  LAYER M1 ;
        RECT 8.796 7.188 8.828 9.696 ;
  LAYER M3 ;
        RECT 8.796 7.208 8.828 7.24 ;
  LAYER M1 ;
        RECT 8.86 7.188 8.892 9.696 ;
  LAYER M3 ;
        RECT 8.86 9.644 8.892 9.676 ;
  LAYER M1 ;
        RECT 8.924 7.188 8.956 9.696 ;
  LAYER M3 ;
        RECT 8.924 7.208 8.956 7.24 ;
  LAYER M1 ;
        RECT 8.988 7.188 9.02 9.696 ;
  LAYER M3 ;
        RECT 8.988 9.644 9.02 9.676 ;
  LAYER M1 ;
        RECT 9.052 7.188 9.084 9.696 ;
  LAYER M3 ;
        RECT 6.684 7.272 6.716 7.304 ;
  LAYER M2 ;
        RECT 9.052 7.336 9.084 7.368 ;
  LAYER M2 ;
        RECT 6.684 7.4 6.716 7.432 ;
  LAYER M2 ;
        RECT 9.052 7.464 9.084 7.496 ;
  LAYER M2 ;
        RECT 6.684 7.528 6.716 7.56 ;
  LAYER M2 ;
        RECT 9.052 7.592 9.084 7.624 ;
  LAYER M2 ;
        RECT 6.684 7.656 6.716 7.688 ;
  LAYER M2 ;
        RECT 9.052 7.72 9.084 7.752 ;
  LAYER M2 ;
        RECT 6.684 7.784 6.716 7.816 ;
  LAYER M2 ;
        RECT 9.052 7.848 9.084 7.88 ;
  LAYER M2 ;
        RECT 6.684 7.912 6.716 7.944 ;
  LAYER M2 ;
        RECT 9.052 7.976 9.084 8.008 ;
  LAYER M2 ;
        RECT 6.684 8.04 6.716 8.072 ;
  LAYER M2 ;
        RECT 9.052 8.104 9.084 8.136 ;
  LAYER M2 ;
        RECT 6.684 8.168 6.716 8.2 ;
  LAYER M2 ;
        RECT 9.052 8.232 9.084 8.264 ;
  LAYER M2 ;
        RECT 6.684 8.296 6.716 8.328 ;
  LAYER M2 ;
        RECT 9.052 8.36 9.084 8.392 ;
  LAYER M2 ;
        RECT 6.684 8.424 6.716 8.456 ;
  LAYER M2 ;
        RECT 9.052 8.488 9.084 8.52 ;
  LAYER M2 ;
        RECT 6.684 8.552 6.716 8.584 ;
  LAYER M2 ;
        RECT 9.052 8.616 9.084 8.648 ;
  LAYER M2 ;
        RECT 6.684 8.68 6.716 8.712 ;
  LAYER M2 ;
        RECT 9.052 8.744 9.084 8.776 ;
  LAYER M2 ;
        RECT 6.684 8.808 6.716 8.84 ;
  LAYER M2 ;
        RECT 9.052 8.872 9.084 8.904 ;
  LAYER M2 ;
        RECT 6.684 8.936 6.716 8.968 ;
  LAYER M2 ;
        RECT 9.052 9 9.084 9.032 ;
  LAYER M2 ;
        RECT 6.684 9.064 6.716 9.096 ;
  LAYER M2 ;
        RECT 9.052 9.128 9.084 9.16 ;
  LAYER M2 ;
        RECT 6.684 9.192 6.716 9.224 ;
  LAYER M2 ;
        RECT 9.052 9.256 9.084 9.288 ;
  LAYER M2 ;
        RECT 6.684 9.32 6.716 9.352 ;
  LAYER M2 ;
        RECT 9.052 9.384 9.084 9.416 ;
  LAYER M2 ;
        RECT 6.684 9.448 6.716 9.48 ;
  LAYER M2 ;
        RECT 9.052 9.512 9.084 9.544 ;
  LAYER M2 ;
        RECT 6.636 7.14 9.132 9.744 ;
  LAYER M1 ;
        RECT 6.684 10.296 6.716 12.804 ;
  LAYER M3 ;
        RECT 6.684 12.752 6.716 12.784 ;
  LAYER M1 ;
        RECT 6.748 10.296 6.78 12.804 ;
  LAYER M3 ;
        RECT 6.748 10.316 6.78 10.348 ;
  LAYER M1 ;
        RECT 6.812 10.296 6.844 12.804 ;
  LAYER M3 ;
        RECT 6.812 12.752 6.844 12.784 ;
  LAYER M1 ;
        RECT 6.876 10.296 6.908 12.804 ;
  LAYER M3 ;
        RECT 6.876 10.316 6.908 10.348 ;
  LAYER M1 ;
        RECT 6.94 10.296 6.972 12.804 ;
  LAYER M3 ;
        RECT 6.94 12.752 6.972 12.784 ;
  LAYER M1 ;
        RECT 7.004 10.296 7.036 12.804 ;
  LAYER M3 ;
        RECT 7.004 10.316 7.036 10.348 ;
  LAYER M1 ;
        RECT 7.068 10.296 7.1 12.804 ;
  LAYER M3 ;
        RECT 7.068 12.752 7.1 12.784 ;
  LAYER M1 ;
        RECT 7.132 10.296 7.164 12.804 ;
  LAYER M3 ;
        RECT 7.132 10.316 7.164 10.348 ;
  LAYER M1 ;
        RECT 7.196 10.296 7.228 12.804 ;
  LAYER M3 ;
        RECT 7.196 12.752 7.228 12.784 ;
  LAYER M1 ;
        RECT 7.26 10.296 7.292 12.804 ;
  LAYER M3 ;
        RECT 7.26 10.316 7.292 10.348 ;
  LAYER M1 ;
        RECT 7.324 10.296 7.356 12.804 ;
  LAYER M3 ;
        RECT 7.324 12.752 7.356 12.784 ;
  LAYER M1 ;
        RECT 7.388 10.296 7.42 12.804 ;
  LAYER M3 ;
        RECT 7.388 10.316 7.42 10.348 ;
  LAYER M1 ;
        RECT 7.452 10.296 7.484 12.804 ;
  LAYER M3 ;
        RECT 7.452 12.752 7.484 12.784 ;
  LAYER M1 ;
        RECT 7.516 10.296 7.548 12.804 ;
  LAYER M3 ;
        RECT 7.516 10.316 7.548 10.348 ;
  LAYER M1 ;
        RECT 7.58 10.296 7.612 12.804 ;
  LAYER M3 ;
        RECT 7.58 12.752 7.612 12.784 ;
  LAYER M1 ;
        RECT 7.644 10.296 7.676 12.804 ;
  LAYER M3 ;
        RECT 7.644 10.316 7.676 10.348 ;
  LAYER M1 ;
        RECT 7.708 10.296 7.74 12.804 ;
  LAYER M3 ;
        RECT 7.708 12.752 7.74 12.784 ;
  LAYER M1 ;
        RECT 7.772 10.296 7.804 12.804 ;
  LAYER M3 ;
        RECT 7.772 10.316 7.804 10.348 ;
  LAYER M1 ;
        RECT 7.836 10.296 7.868 12.804 ;
  LAYER M3 ;
        RECT 7.836 12.752 7.868 12.784 ;
  LAYER M1 ;
        RECT 7.9 10.296 7.932 12.804 ;
  LAYER M3 ;
        RECT 7.9 10.316 7.932 10.348 ;
  LAYER M1 ;
        RECT 7.964 10.296 7.996 12.804 ;
  LAYER M3 ;
        RECT 7.964 12.752 7.996 12.784 ;
  LAYER M1 ;
        RECT 8.028 10.296 8.06 12.804 ;
  LAYER M3 ;
        RECT 8.028 10.316 8.06 10.348 ;
  LAYER M1 ;
        RECT 8.092 10.296 8.124 12.804 ;
  LAYER M3 ;
        RECT 8.092 12.752 8.124 12.784 ;
  LAYER M1 ;
        RECT 8.156 10.296 8.188 12.804 ;
  LAYER M3 ;
        RECT 8.156 10.316 8.188 10.348 ;
  LAYER M1 ;
        RECT 8.22 10.296 8.252 12.804 ;
  LAYER M3 ;
        RECT 8.22 12.752 8.252 12.784 ;
  LAYER M1 ;
        RECT 8.284 10.296 8.316 12.804 ;
  LAYER M3 ;
        RECT 8.284 10.316 8.316 10.348 ;
  LAYER M1 ;
        RECT 8.348 10.296 8.38 12.804 ;
  LAYER M3 ;
        RECT 8.348 12.752 8.38 12.784 ;
  LAYER M1 ;
        RECT 8.412 10.296 8.444 12.804 ;
  LAYER M3 ;
        RECT 8.412 10.316 8.444 10.348 ;
  LAYER M1 ;
        RECT 8.476 10.296 8.508 12.804 ;
  LAYER M3 ;
        RECT 8.476 12.752 8.508 12.784 ;
  LAYER M1 ;
        RECT 8.54 10.296 8.572 12.804 ;
  LAYER M3 ;
        RECT 8.54 10.316 8.572 10.348 ;
  LAYER M1 ;
        RECT 8.604 10.296 8.636 12.804 ;
  LAYER M3 ;
        RECT 8.604 12.752 8.636 12.784 ;
  LAYER M1 ;
        RECT 8.668 10.296 8.7 12.804 ;
  LAYER M3 ;
        RECT 8.668 10.316 8.7 10.348 ;
  LAYER M1 ;
        RECT 8.732 10.296 8.764 12.804 ;
  LAYER M3 ;
        RECT 8.732 12.752 8.764 12.784 ;
  LAYER M1 ;
        RECT 8.796 10.296 8.828 12.804 ;
  LAYER M3 ;
        RECT 8.796 10.316 8.828 10.348 ;
  LAYER M1 ;
        RECT 8.86 10.296 8.892 12.804 ;
  LAYER M3 ;
        RECT 8.86 12.752 8.892 12.784 ;
  LAYER M1 ;
        RECT 8.924 10.296 8.956 12.804 ;
  LAYER M3 ;
        RECT 8.924 10.316 8.956 10.348 ;
  LAYER M1 ;
        RECT 8.988 10.296 9.02 12.804 ;
  LAYER M3 ;
        RECT 8.988 12.752 9.02 12.784 ;
  LAYER M1 ;
        RECT 9.052 10.296 9.084 12.804 ;
  LAYER M3 ;
        RECT 6.684 10.38 6.716 10.412 ;
  LAYER M2 ;
        RECT 9.052 10.444 9.084 10.476 ;
  LAYER M2 ;
        RECT 6.684 10.508 6.716 10.54 ;
  LAYER M2 ;
        RECT 9.052 10.572 9.084 10.604 ;
  LAYER M2 ;
        RECT 6.684 10.636 6.716 10.668 ;
  LAYER M2 ;
        RECT 9.052 10.7 9.084 10.732 ;
  LAYER M2 ;
        RECT 6.684 10.764 6.716 10.796 ;
  LAYER M2 ;
        RECT 9.052 10.828 9.084 10.86 ;
  LAYER M2 ;
        RECT 6.684 10.892 6.716 10.924 ;
  LAYER M2 ;
        RECT 9.052 10.956 9.084 10.988 ;
  LAYER M2 ;
        RECT 6.684 11.02 6.716 11.052 ;
  LAYER M2 ;
        RECT 9.052 11.084 9.084 11.116 ;
  LAYER M2 ;
        RECT 6.684 11.148 6.716 11.18 ;
  LAYER M2 ;
        RECT 9.052 11.212 9.084 11.244 ;
  LAYER M2 ;
        RECT 6.684 11.276 6.716 11.308 ;
  LAYER M2 ;
        RECT 9.052 11.34 9.084 11.372 ;
  LAYER M2 ;
        RECT 6.684 11.404 6.716 11.436 ;
  LAYER M2 ;
        RECT 9.052 11.468 9.084 11.5 ;
  LAYER M2 ;
        RECT 6.684 11.532 6.716 11.564 ;
  LAYER M2 ;
        RECT 9.052 11.596 9.084 11.628 ;
  LAYER M2 ;
        RECT 6.684 11.66 6.716 11.692 ;
  LAYER M2 ;
        RECT 9.052 11.724 9.084 11.756 ;
  LAYER M2 ;
        RECT 6.684 11.788 6.716 11.82 ;
  LAYER M2 ;
        RECT 9.052 11.852 9.084 11.884 ;
  LAYER M2 ;
        RECT 6.684 11.916 6.716 11.948 ;
  LAYER M2 ;
        RECT 9.052 11.98 9.084 12.012 ;
  LAYER M2 ;
        RECT 6.684 12.044 6.716 12.076 ;
  LAYER M2 ;
        RECT 9.052 12.108 9.084 12.14 ;
  LAYER M2 ;
        RECT 6.684 12.172 6.716 12.204 ;
  LAYER M2 ;
        RECT 9.052 12.236 9.084 12.268 ;
  LAYER M2 ;
        RECT 6.684 12.3 6.716 12.332 ;
  LAYER M2 ;
        RECT 9.052 12.364 9.084 12.396 ;
  LAYER M2 ;
        RECT 6.684 12.428 6.716 12.46 ;
  LAYER M2 ;
        RECT 9.052 12.492 9.084 12.524 ;
  LAYER M2 ;
        RECT 6.684 12.556 6.716 12.588 ;
  LAYER M2 ;
        RECT 9.052 12.62 9.084 12.652 ;
  LAYER M2 ;
        RECT 6.636 10.248 9.132 12.852 ;
  LAYER M1 ;
        RECT 6.684 13.404 6.716 15.912 ;
  LAYER M3 ;
        RECT 6.684 15.86 6.716 15.892 ;
  LAYER M1 ;
        RECT 6.748 13.404 6.78 15.912 ;
  LAYER M3 ;
        RECT 6.748 13.424 6.78 13.456 ;
  LAYER M1 ;
        RECT 6.812 13.404 6.844 15.912 ;
  LAYER M3 ;
        RECT 6.812 15.86 6.844 15.892 ;
  LAYER M1 ;
        RECT 6.876 13.404 6.908 15.912 ;
  LAYER M3 ;
        RECT 6.876 13.424 6.908 13.456 ;
  LAYER M1 ;
        RECT 6.94 13.404 6.972 15.912 ;
  LAYER M3 ;
        RECT 6.94 15.86 6.972 15.892 ;
  LAYER M1 ;
        RECT 7.004 13.404 7.036 15.912 ;
  LAYER M3 ;
        RECT 7.004 13.424 7.036 13.456 ;
  LAYER M1 ;
        RECT 7.068 13.404 7.1 15.912 ;
  LAYER M3 ;
        RECT 7.068 15.86 7.1 15.892 ;
  LAYER M1 ;
        RECT 7.132 13.404 7.164 15.912 ;
  LAYER M3 ;
        RECT 7.132 13.424 7.164 13.456 ;
  LAYER M1 ;
        RECT 7.196 13.404 7.228 15.912 ;
  LAYER M3 ;
        RECT 7.196 15.86 7.228 15.892 ;
  LAYER M1 ;
        RECT 7.26 13.404 7.292 15.912 ;
  LAYER M3 ;
        RECT 7.26 13.424 7.292 13.456 ;
  LAYER M1 ;
        RECT 7.324 13.404 7.356 15.912 ;
  LAYER M3 ;
        RECT 7.324 15.86 7.356 15.892 ;
  LAYER M1 ;
        RECT 7.388 13.404 7.42 15.912 ;
  LAYER M3 ;
        RECT 7.388 13.424 7.42 13.456 ;
  LAYER M1 ;
        RECT 7.452 13.404 7.484 15.912 ;
  LAYER M3 ;
        RECT 7.452 15.86 7.484 15.892 ;
  LAYER M1 ;
        RECT 7.516 13.404 7.548 15.912 ;
  LAYER M3 ;
        RECT 7.516 13.424 7.548 13.456 ;
  LAYER M1 ;
        RECT 7.58 13.404 7.612 15.912 ;
  LAYER M3 ;
        RECT 7.58 15.86 7.612 15.892 ;
  LAYER M1 ;
        RECT 7.644 13.404 7.676 15.912 ;
  LAYER M3 ;
        RECT 7.644 13.424 7.676 13.456 ;
  LAYER M1 ;
        RECT 7.708 13.404 7.74 15.912 ;
  LAYER M3 ;
        RECT 7.708 15.86 7.74 15.892 ;
  LAYER M1 ;
        RECT 7.772 13.404 7.804 15.912 ;
  LAYER M3 ;
        RECT 7.772 13.424 7.804 13.456 ;
  LAYER M1 ;
        RECT 7.836 13.404 7.868 15.912 ;
  LAYER M3 ;
        RECT 7.836 15.86 7.868 15.892 ;
  LAYER M1 ;
        RECT 7.9 13.404 7.932 15.912 ;
  LAYER M3 ;
        RECT 7.9 13.424 7.932 13.456 ;
  LAYER M1 ;
        RECT 7.964 13.404 7.996 15.912 ;
  LAYER M3 ;
        RECT 7.964 15.86 7.996 15.892 ;
  LAYER M1 ;
        RECT 8.028 13.404 8.06 15.912 ;
  LAYER M3 ;
        RECT 8.028 13.424 8.06 13.456 ;
  LAYER M1 ;
        RECT 8.092 13.404 8.124 15.912 ;
  LAYER M3 ;
        RECT 8.092 15.86 8.124 15.892 ;
  LAYER M1 ;
        RECT 8.156 13.404 8.188 15.912 ;
  LAYER M3 ;
        RECT 8.156 13.424 8.188 13.456 ;
  LAYER M1 ;
        RECT 8.22 13.404 8.252 15.912 ;
  LAYER M3 ;
        RECT 8.22 15.86 8.252 15.892 ;
  LAYER M1 ;
        RECT 8.284 13.404 8.316 15.912 ;
  LAYER M3 ;
        RECT 8.284 13.424 8.316 13.456 ;
  LAYER M1 ;
        RECT 8.348 13.404 8.38 15.912 ;
  LAYER M3 ;
        RECT 8.348 15.86 8.38 15.892 ;
  LAYER M1 ;
        RECT 8.412 13.404 8.444 15.912 ;
  LAYER M3 ;
        RECT 8.412 13.424 8.444 13.456 ;
  LAYER M1 ;
        RECT 8.476 13.404 8.508 15.912 ;
  LAYER M3 ;
        RECT 8.476 15.86 8.508 15.892 ;
  LAYER M1 ;
        RECT 8.54 13.404 8.572 15.912 ;
  LAYER M3 ;
        RECT 8.54 13.424 8.572 13.456 ;
  LAYER M1 ;
        RECT 8.604 13.404 8.636 15.912 ;
  LAYER M3 ;
        RECT 8.604 15.86 8.636 15.892 ;
  LAYER M1 ;
        RECT 8.668 13.404 8.7 15.912 ;
  LAYER M3 ;
        RECT 8.668 13.424 8.7 13.456 ;
  LAYER M1 ;
        RECT 8.732 13.404 8.764 15.912 ;
  LAYER M3 ;
        RECT 8.732 15.86 8.764 15.892 ;
  LAYER M1 ;
        RECT 8.796 13.404 8.828 15.912 ;
  LAYER M3 ;
        RECT 8.796 13.424 8.828 13.456 ;
  LAYER M1 ;
        RECT 8.86 13.404 8.892 15.912 ;
  LAYER M3 ;
        RECT 8.86 15.86 8.892 15.892 ;
  LAYER M1 ;
        RECT 8.924 13.404 8.956 15.912 ;
  LAYER M3 ;
        RECT 8.924 13.424 8.956 13.456 ;
  LAYER M1 ;
        RECT 8.988 13.404 9.02 15.912 ;
  LAYER M3 ;
        RECT 8.988 15.86 9.02 15.892 ;
  LAYER M1 ;
        RECT 9.052 13.404 9.084 15.912 ;
  LAYER M3 ;
        RECT 6.684 13.488 6.716 13.52 ;
  LAYER M2 ;
        RECT 9.052 13.552 9.084 13.584 ;
  LAYER M2 ;
        RECT 6.684 13.616 6.716 13.648 ;
  LAYER M2 ;
        RECT 9.052 13.68 9.084 13.712 ;
  LAYER M2 ;
        RECT 6.684 13.744 6.716 13.776 ;
  LAYER M2 ;
        RECT 9.052 13.808 9.084 13.84 ;
  LAYER M2 ;
        RECT 6.684 13.872 6.716 13.904 ;
  LAYER M2 ;
        RECT 9.052 13.936 9.084 13.968 ;
  LAYER M2 ;
        RECT 6.684 14 6.716 14.032 ;
  LAYER M2 ;
        RECT 9.052 14.064 9.084 14.096 ;
  LAYER M2 ;
        RECT 6.684 14.128 6.716 14.16 ;
  LAYER M2 ;
        RECT 9.052 14.192 9.084 14.224 ;
  LAYER M2 ;
        RECT 6.684 14.256 6.716 14.288 ;
  LAYER M2 ;
        RECT 9.052 14.32 9.084 14.352 ;
  LAYER M2 ;
        RECT 6.684 14.384 6.716 14.416 ;
  LAYER M2 ;
        RECT 9.052 14.448 9.084 14.48 ;
  LAYER M2 ;
        RECT 6.684 14.512 6.716 14.544 ;
  LAYER M2 ;
        RECT 9.052 14.576 9.084 14.608 ;
  LAYER M2 ;
        RECT 6.684 14.64 6.716 14.672 ;
  LAYER M2 ;
        RECT 9.052 14.704 9.084 14.736 ;
  LAYER M2 ;
        RECT 6.684 14.768 6.716 14.8 ;
  LAYER M2 ;
        RECT 9.052 14.832 9.084 14.864 ;
  LAYER M2 ;
        RECT 6.684 14.896 6.716 14.928 ;
  LAYER M2 ;
        RECT 9.052 14.96 9.084 14.992 ;
  LAYER M2 ;
        RECT 6.684 15.024 6.716 15.056 ;
  LAYER M2 ;
        RECT 9.052 15.088 9.084 15.12 ;
  LAYER M2 ;
        RECT 6.684 15.152 6.716 15.184 ;
  LAYER M2 ;
        RECT 9.052 15.216 9.084 15.248 ;
  LAYER M2 ;
        RECT 6.684 15.28 6.716 15.312 ;
  LAYER M2 ;
        RECT 9.052 15.344 9.084 15.376 ;
  LAYER M2 ;
        RECT 6.684 15.408 6.716 15.44 ;
  LAYER M2 ;
        RECT 9.052 15.472 9.084 15.504 ;
  LAYER M2 ;
        RECT 6.684 15.536 6.716 15.568 ;
  LAYER M2 ;
        RECT 9.052 15.6 9.084 15.632 ;
  LAYER M2 ;
        RECT 6.684 15.664 6.716 15.696 ;
  LAYER M2 ;
        RECT 9.052 15.728 9.084 15.76 ;
  LAYER M2 ;
        RECT 6.636 13.356 9.132 15.96 ;
  LAYER M1 ;
        RECT 6.684 16.512 6.716 19.02 ;
  LAYER M3 ;
        RECT 6.684 18.968 6.716 19 ;
  LAYER M1 ;
        RECT 6.748 16.512 6.78 19.02 ;
  LAYER M3 ;
        RECT 6.748 16.532 6.78 16.564 ;
  LAYER M1 ;
        RECT 6.812 16.512 6.844 19.02 ;
  LAYER M3 ;
        RECT 6.812 18.968 6.844 19 ;
  LAYER M1 ;
        RECT 6.876 16.512 6.908 19.02 ;
  LAYER M3 ;
        RECT 6.876 16.532 6.908 16.564 ;
  LAYER M1 ;
        RECT 6.94 16.512 6.972 19.02 ;
  LAYER M3 ;
        RECT 6.94 18.968 6.972 19 ;
  LAYER M1 ;
        RECT 7.004 16.512 7.036 19.02 ;
  LAYER M3 ;
        RECT 7.004 16.532 7.036 16.564 ;
  LAYER M1 ;
        RECT 7.068 16.512 7.1 19.02 ;
  LAYER M3 ;
        RECT 7.068 18.968 7.1 19 ;
  LAYER M1 ;
        RECT 7.132 16.512 7.164 19.02 ;
  LAYER M3 ;
        RECT 7.132 16.532 7.164 16.564 ;
  LAYER M1 ;
        RECT 7.196 16.512 7.228 19.02 ;
  LAYER M3 ;
        RECT 7.196 18.968 7.228 19 ;
  LAYER M1 ;
        RECT 7.26 16.512 7.292 19.02 ;
  LAYER M3 ;
        RECT 7.26 16.532 7.292 16.564 ;
  LAYER M1 ;
        RECT 7.324 16.512 7.356 19.02 ;
  LAYER M3 ;
        RECT 7.324 18.968 7.356 19 ;
  LAYER M1 ;
        RECT 7.388 16.512 7.42 19.02 ;
  LAYER M3 ;
        RECT 7.388 16.532 7.42 16.564 ;
  LAYER M1 ;
        RECT 7.452 16.512 7.484 19.02 ;
  LAYER M3 ;
        RECT 7.452 18.968 7.484 19 ;
  LAYER M1 ;
        RECT 7.516 16.512 7.548 19.02 ;
  LAYER M3 ;
        RECT 7.516 16.532 7.548 16.564 ;
  LAYER M1 ;
        RECT 7.58 16.512 7.612 19.02 ;
  LAYER M3 ;
        RECT 7.58 18.968 7.612 19 ;
  LAYER M1 ;
        RECT 7.644 16.512 7.676 19.02 ;
  LAYER M3 ;
        RECT 7.644 16.532 7.676 16.564 ;
  LAYER M1 ;
        RECT 7.708 16.512 7.74 19.02 ;
  LAYER M3 ;
        RECT 7.708 18.968 7.74 19 ;
  LAYER M1 ;
        RECT 7.772 16.512 7.804 19.02 ;
  LAYER M3 ;
        RECT 7.772 16.532 7.804 16.564 ;
  LAYER M1 ;
        RECT 7.836 16.512 7.868 19.02 ;
  LAYER M3 ;
        RECT 7.836 18.968 7.868 19 ;
  LAYER M1 ;
        RECT 7.9 16.512 7.932 19.02 ;
  LAYER M3 ;
        RECT 7.9 16.532 7.932 16.564 ;
  LAYER M1 ;
        RECT 7.964 16.512 7.996 19.02 ;
  LAYER M3 ;
        RECT 7.964 18.968 7.996 19 ;
  LAYER M1 ;
        RECT 8.028 16.512 8.06 19.02 ;
  LAYER M3 ;
        RECT 8.028 16.532 8.06 16.564 ;
  LAYER M1 ;
        RECT 8.092 16.512 8.124 19.02 ;
  LAYER M3 ;
        RECT 8.092 18.968 8.124 19 ;
  LAYER M1 ;
        RECT 8.156 16.512 8.188 19.02 ;
  LAYER M3 ;
        RECT 8.156 16.532 8.188 16.564 ;
  LAYER M1 ;
        RECT 8.22 16.512 8.252 19.02 ;
  LAYER M3 ;
        RECT 8.22 18.968 8.252 19 ;
  LAYER M1 ;
        RECT 8.284 16.512 8.316 19.02 ;
  LAYER M3 ;
        RECT 8.284 16.532 8.316 16.564 ;
  LAYER M1 ;
        RECT 8.348 16.512 8.38 19.02 ;
  LAYER M3 ;
        RECT 8.348 18.968 8.38 19 ;
  LAYER M1 ;
        RECT 8.412 16.512 8.444 19.02 ;
  LAYER M3 ;
        RECT 8.412 16.532 8.444 16.564 ;
  LAYER M1 ;
        RECT 8.476 16.512 8.508 19.02 ;
  LAYER M3 ;
        RECT 8.476 18.968 8.508 19 ;
  LAYER M1 ;
        RECT 8.54 16.512 8.572 19.02 ;
  LAYER M3 ;
        RECT 8.54 16.532 8.572 16.564 ;
  LAYER M1 ;
        RECT 8.604 16.512 8.636 19.02 ;
  LAYER M3 ;
        RECT 8.604 18.968 8.636 19 ;
  LAYER M1 ;
        RECT 8.668 16.512 8.7 19.02 ;
  LAYER M3 ;
        RECT 8.668 16.532 8.7 16.564 ;
  LAYER M1 ;
        RECT 8.732 16.512 8.764 19.02 ;
  LAYER M3 ;
        RECT 8.732 18.968 8.764 19 ;
  LAYER M1 ;
        RECT 8.796 16.512 8.828 19.02 ;
  LAYER M3 ;
        RECT 8.796 16.532 8.828 16.564 ;
  LAYER M1 ;
        RECT 8.86 16.512 8.892 19.02 ;
  LAYER M3 ;
        RECT 8.86 18.968 8.892 19 ;
  LAYER M1 ;
        RECT 8.924 16.512 8.956 19.02 ;
  LAYER M3 ;
        RECT 8.924 16.532 8.956 16.564 ;
  LAYER M1 ;
        RECT 8.988 16.512 9.02 19.02 ;
  LAYER M3 ;
        RECT 8.988 18.968 9.02 19 ;
  LAYER M1 ;
        RECT 9.052 16.512 9.084 19.02 ;
  LAYER M3 ;
        RECT 6.684 16.596 6.716 16.628 ;
  LAYER M2 ;
        RECT 9.052 16.66 9.084 16.692 ;
  LAYER M2 ;
        RECT 6.684 16.724 6.716 16.756 ;
  LAYER M2 ;
        RECT 9.052 16.788 9.084 16.82 ;
  LAYER M2 ;
        RECT 6.684 16.852 6.716 16.884 ;
  LAYER M2 ;
        RECT 9.052 16.916 9.084 16.948 ;
  LAYER M2 ;
        RECT 6.684 16.98 6.716 17.012 ;
  LAYER M2 ;
        RECT 9.052 17.044 9.084 17.076 ;
  LAYER M2 ;
        RECT 6.684 17.108 6.716 17.14 ;
  LAYER M2 ;
        RECT 9.052 17.172 9.084 17.204 ;
  LAYER M2 ;
        RECT 6.684 17.236 6.716 17.268 ;
  LAYER M2 ;
        RECT 9.052 17.3 9.084 17.332 ;
  LAYER M2 ;
        RECT 6.684 17.364 6.716 17.396 ;
  LAYER M2 ;
        RECT 9.052 17.428 9.084 17.46 ;
  LAYER M2 ;
        RECT 6.684 17.492 6.716 17.524 ;
  LAYER M2 ;
        RECT 9.052 17.556 9.084 17.588 ;
  LAYER M2 ;
        RECT 6.684 17.62 6.716 17.652 ;
  LAYER M2 ;
        RECT 9.052 17.684 9.084 17.716 ;
  LAYER M2 ;
        RECT 6.684 17.748 6.716 17.78 ;
  LAYER M2 ;
        RECT 9.052 17.812 9.084 17.844 ;
  LAYER M2 ;
        RECT 6.684 17.876 6.716 17.908 ;
  LAYER M2 ;
        RECT 9.052 17.94 9.084 17.972 ;
  LAYER M2 ;
        RECT 6.684 18.004 6.716 18.036 ;
  LAYER M2 ;
        RECT 9.052 18.068 9.084 18.1 ;
  LAYER M2 ;
        RECT 6.684 18.132 6.716 18.164 ;
  LAYER M2 ;
        RECT 9.052 18.196 9.084 18.228 ;
  LAYER M2 ;
        RECT 6.684 18.26 6.716 18.292 ;
  LAYER M2 ;
        RECT 9.052 18.324 9.084 18.356 ;
  LAYER M2 ;
        RECT 6.684 18.388 6.716 18.42 ;
  LAYER M2 ;
        RECT 9.052 18.452 9.084 18.484 ;
  LAYER M2 ;
        RECT 6.684 18.516 6.716 18.548 ;
  LAYER M2 ;
        RECT 9.052 18.58 9.084 18.612 ;
  LAYER M2 ;
        RECT 6.684 18.644 6.716 18.676 ;
  LAYER M2 ;
        RECT 9.052 18.708 9.084 18.74 ;
  LAYER M2 ;
        RECT 6.684 18.772 6.716 18.804 ;
  LAYER M2 ;
        RECT 9.052 18.836 9.084 18.868 ;
  LAYER M2 ;
        RECT 6.636 16.464 9.132 19.068 ;
  LAYER M1 ;
        RECT 6.684 19.62 6.716 22.128 ;
  LAYER M3 ;
        RECT 6.684 22.076 6.716 22.108 ;
  LAYER M1 ;
        RECT 6.748 19.62 6.78 22.128 ;
  LAYER M3 ;
        RECT 6.748 19.64 6.78 19.672 ;
  LAYER M1 ;
        RECT 6.812 19.62 6.844 22.128 ;
  LAYER M3 ;
        RECT 6.812 22.076 6.844 22.108 ;
  LAYER M1 ;
        RECT 6.876 19.62 6.908 22.128 ;
  LAYER M3 ;
        RECT 6.876 19.64 6.908 19.672 ;
  LAYER M1 ;
        RECT 6.94 19.62 6.972 22.128 ;
  LAYER M3 ;
        RECT 6.94 22.076 6.972 22.108 ;
  LAYER M1 ;
        RECT 7.004 19.62 7.036 22.128 ;
  LAYER M3 ;
        RECT 7.004 19.64 7.036 19.672 ;
  LAYER M1 ;
        RECT 7.068 19.62 7.1 22.128 ;
  LAYER M3 ;
        RECT 7.068 22.076 7.1 22.108 ;
  LAYER M1 ;
        RECT 7.132 19.62 7.164 22.128 ;
  LAYER M3 ;
        RECT 7.132 19.64 7.164 19.672 ;
  LAYER M1 ;
        RECT 7.196 19.62 7.228 22.128 ;
  LAYER M3 ;
        RECT 7.196 22.076 7.228 22.108 ;
  LAYER M1 ;
        RECT 7.26 19.62 7.292 22.128 ;
  LAYER M3 ;
        RECT 7.26 19.64 7.292 19.672 ;
  LAYER M1 ;
        RECT 7.324 19.62 7.356 22.128 ;
  LAYER M3 ;
        RECT 7.324 22.076 7.356 22.108 ;
  LAYER M1 ;
        RECT 7.388 19.62 7.42 22.128 ;
  LAYER M3 ;
        RECT 7.388 19.64 7.42 19.672 ;
  LAYER M1 ;
        RECT 7.452 19.62 7.484 22.128 ;
  LAYER M3 ;
        RECT 7.452 22.076 7.484 22.108 ;
  LAYER M1 ;
        RECT 7.516 19.62 7.548 22.128 ;
  LAYER M3 ;
        RECT 7.516 19.64 7.548 19.672 ;
  LAYER M1 ;
        RECT 7.58 19.62 7.612 22.128 ;
  LAYER M3 ;
        RECT 7.58 22.076 7.612 22.108 ;
  LAYER M1 ;
        RECT 7.644 19.62 7.676 22.128 ;
  LAYER M3 ;
        RECT 7.644 19.64 7.676 19.672 ;
  LAYER M1 ;
        RECT 7.708 19.62 7.74 22.128 ;
  LAYER M3 ;
        RECT 7.708 22.076 7.74 22.108 ;
  LAYER M1 ;
        RECT 7.772 19.62 7.804 22.128 ;
  LAYER M3 ;
        RECT 7.772 19.64 7.804 19.672 ;
  LAYER M1 ;
        RECT 7.836 19.62 7.868 22.128 ;
  LAYER M3 ;
        RECT 7.836 22.076 7.868 22.108 ;
  LAYER M1 ;
        RECT 7.9 19.62 7.932 22.128 ;
  LAYER M3 ;
        RECT 7.9 19.64 7.932 19.672 ;
  LAYER M1 ;
        RECT 7.964 19.62 7.996 22.128 ;
  LAYER M3 ;
        RECT 7.964 22.076 7.996 22.108 ;
  LAYER M1 ;
        RECT 8.028 19.62 8.06 22.128 ;
  LAYER M3 ;
        RECT 8.028 19.64 8.06 19.672 ;
  LAYER M1 ;
        RECT 8.092 19.62 8.124 22.128 ;
  LAYER M3 ;
        RECT 8.092 22.076 8.124 22.108 ;
  LAYER M1 ;
        RECT 8.156 19.62 8.188 22.128 ;
  LAYER M3 ;
        RECT 8.156 19.64 8.188 19.672 ;
  LAYER M1 ;
        RECT 8.22 19.62 8.252 22.128 ;
  LAYER M3 ;
        RECT 8.22 22.076 8.252 22.108 ;
  LAYER M1 ;
        RECT 8.284 19.62 8.316 22.128 ;
  LAYER M3 ;
        RECT 8.284 19.64 8.316 19.672 ;
  LAYER M1 ;
        RECT 8.348 19.62 8.38 22.128 ;
  LAYER M3 ;
        RECT 8.348 22.076 8.38 22.108 ;
  LAYER M1 ;
        RECT 8.412 19.62 8.444 22.128 ;
  LAYER M3 ;
        RECT 8.412 19.64 8.444 19.672 ;
  LAYER M1 ;
        RECT 8.476 19.62 8.508 22.128 ;
  LAYER M3 ;
        RECT 8.476 22.076 8.508 22.108 ;
  LAYER M1 ;
        RECT 8.54 19.62 8.572 22.128 ;
  LAYER M3 ;
        RECT 8.54 19.64 8.572 19.672 ;
  LAYER M1 ;
        RECT 8.604 19.62 8.636 22.128 ;
  LAYER M3 ;
        RECT 8.604 22.076 8.636 22.108 ;
  LAYER M1 ;
        RECT 8.668 19.62 8.7 22.128 ;
  LAYER M3 ;
        RECT 8.668 19.64 8.7 19.672 ;
  LAYER M1 ;
        RECT 8.732 19.62 8.764 22.128 ;
  LAYER M3 ;
        RECT 8.732 22.076 8.764 22.108 ;
  LAYER M1 ;
        RECT 8.796 19.62 8.828 22.128 ;
  LAYER M3 ;
        RECT 8.796 19.64 8.828 19.672 ;
  LAYER M1 ;
        RECT 8.86 19.62 8.892 22.128 ;
  LAYER M3 ;
        RECT 8.86 22.076 8.892 22.108 ;
  LAYER M1 ;
        RECT 8.924 19.62 8.956 22.128 ;
  LAYER M3 ;
        RECT 8.924 19.64 8.956 19.672 ;
  LAYER M1 ;
        RECT 8.988 19.62 9.02 22.128 ;
  LAYER M3 ;
        RECT 8.988 22.076 9.02 22.108 ;
  LAYER M1 ;
        RECT 9.052 19.62 9.084 22.128 ;
  LAYER M3 ;
        RECT 6.684 19.704 6.716 19.736 ;
  LAYER M2 ;
        RECT 9.052 19.768 9.084 19.8 ;
  LAYER M2 ;
        RECT 6.684 19.832 6.716 19.864 ;
  LAYER M2 ;
        RECT 9.052 19.896 9.084 19.928 ;
  LAYER M2 ;
        RECT 6.684 19.96 6.716 19.992 ;
  LAYER M2 ;
        RECT 9.052 20.024 9.084 20.056 ;
  LAYER M2 ;
        RECT 6.684 20.088 6.716 20.12 ;
  LAYER M2 ;
        RECT 9.052 20.152 9.084 20.184 ;
  LAYER M2 ;
        RECT 6.684 20.216 6.716 20.248 ;
  LAYER M2 ;
        RECT 9.052 20.28 9.084 20.312 ;
  LAYER M2 ;
        RECT 6.684 20.344 6.716 20.376 ;
  LAYER M2 ;
        RECT 9.052 20.408 9.084 20.44 ;
  LAYER M2 ;
        RECT 6.684 20.472 6.716 20.504 ;
  LAYER M2 ;
        RECT 9.052 20.536 9.084 20.568 ;
  LAYER M2 ;
        RECT 6.684 20.6 6.716 20.632 ;
  LAYER M2 ;
        RECT 9.052 20.664 9.084 20.696 ;
  LAYER M2 ;
        RECT 6.684 20.728 6.716 20.76 ;
  LAYER M2 ;
        RECT 9.052 20.792 9.084 20.824 ;
  LAYER M2 ;
        RECT 6.684 20.856 6.716 20.888 ;
  LAYER M2 ;
        RECT 9.052 20.92 9.084 20.952 ;
  LAYER M2 ;
        RECT 6.684 20.984 6.716 21.016 ;
  LAYER M2 ;
        RECT 9.052 21.048 9.084 21.08 ;
  LAYER M2 ;
        RECT 6.684 21.112 6.716 21.144 ;
  LAYER M2 ;
        RECT 9.052 21.176 9.084 21.208 ;
  LAYER M2 ;
        RECT 6.684 21.24 6.716 21.272 ;
  LAYER M2 ;
        RECT 9.052 21.304 9.084 21.336 ;
  LAYER M2 ;
        RECT 6.684 21.368 6.716 21.4 ;
  LAYER M2 ;
        RECT 9.052 21.432 9.084 21.464 ;
  LAYER M2 ;
        RECT 6.684 21.496 6.716 21.528 ;
  LAYER M2 ;
        RECT 9.052 21.56 9.084 21.592 ;
  LAYER M2 ;
        RECT 6.684 21.624 6.716 21.656 ;
  LAYER M2 ;
        RECT 9.052 21.688 9.084 21.72 ;
  LAYER M2 ;
        RECT 6.684 21.752 6.716 21.784 ;
  LAYER M2 ;
        RECT 9.052 21.816 9.084 21.848 ;
  LAYER M2 ;
        RECT 6.684 21.88 6.716 21.912 ;
  LAYER M2 ;
        RECT 9.052 21.944 9.084 21.976 ;
  LAYER M2 ;
        RECT 6.636 19.572 9.132 22.176 ;
  LAYER M1 ;
        RECT 9.98 0.972 10.012 3.48 ;
  LAYER M3 ;
        RECT 9.98 3.428 10.012 3.46 ;
  LAYER M1 ;
        RECT 10.044 0.972 10.076 3.48 ;
  LAYER M3 ;
        RECT 10.044 0.992 10.076 1.024 ;
  LAYER M1 ;
        RECT 10.108 0.972 10.14 3.48 ;
  LAYER M3 ;
        RECT 10.108 3.428 10.14 3.46 ;
  LAYER M1 ;
        RECT 10.172 0.972 10.204 3.48 ;
  LAYER M3 ;
        RECT 10.172 0.992 10.204 1.024 ;
  LAYER M1 ;
        RECT 10.236 0.972 10.268 3.48 ;
  LAYER M3 ;
        RECT 10.236 3.428 10.268 3.46 ;
  LAYER M1 ;
        RECT 10.3 0.972 10.332 3.48 ;
  LAYER M3 ;
        RECT 10.3 0.992 10.332 1.024 ;
  LAYER M1 ;
        RECT 10.364 0.972 10.396 3.48 ;
  LAYER M3 ;
        RECT 10.364 3.428 10.396 3.46 ;
  LAYER M1 ;
        RECT 10.428 0.972 10.46 3.48 ;
  LAYER M3 ;
        RECT 10.428 0.992 10.46 1.024 ;
  LAYER M1 ;
        RECT 10.492 0.972 10.524 3.48 ;
  LAYER M3 ;
        RECT 10.492 3.428 10.524 3.46 ;
  LAYER M1 ;
        RECT 10.556 0.972 10.588 3.48 ;
  LAYER M3 ;
        RECT 10.556 0.992 10.588 1.024 ;
  LAYER M1 ;
        RECT 10.62 0.972 10.652 3.48 ;
  LAYER M3 ;
        RECT 10.62 3.428 10.652 3.46 ;
  LAYER M1 ;
        RECT 10.684 0.972 10.716 3.48 ;
  LAYER M3 ;
        RECT 10.684 0.992 10.716 1.024 ;
  LAYER M1 ;
        RECT 10.748 0.972 10.78 3.48 ;
  LAYER M3 ;
        RECT 10.748 3.428 10.78 3.46 ;
  LAYER M1 ;
        RECT 10.812 0.972 10.844 3.48 ;
  LAYER M3 ;
        RECT 10.812 0.992 10.844 1.024 ;
  LAYER M1 ;
        RECT 10.876 0.972 10.908 3.48 ;
  LAYER M3 ;
        RECT 10.876 3.428 10.908 3.46 ;
  LAYER M1 ;
        RECT 10.94 0.972 10.972 3.48 ;
  LAYER M3 ;
        RECT 10.94 0.992 10.972 1.024 ;
  LAYER M1 ;
        RECT 11.004 0.972 11.036 3.48 ;
  LAYER M3 ;
        RECT 11.004 3.428 11.036 3.46 ;
  LAYER M1 ;
        RECT 11.068 0.972 11.1 3.48 ;
  LAYER M3 ;
        RECT 11.068 0.992 11.1 1.024 ;
  LAYER M1 ;
        RECT 11.132 0.972 11.164 3.48 ;
  LAYER M3 ;
        RECT 11.132 3.428 11.164 3.46 ;
  LAYER M1 ;
        RECT 11.196 0.972 11.228 3.48 ;
  LAYER M3 ;
        RECT 11.196 0.992 11.228 1.024 ;
  LAYER M1 ;
        RECT 11.26 0.972 11.292 3.48 ;
  LAYER M3 ;
        RECT 11.26 3.428 11.292 3.46 ;
  LAYER M1 ;
        RECT 11.324 0.972 11.356 3.48 ;
  LAYER M3 ;
        RECT 11.324 0.992 11.356 1.024 ;
  LAYER M1 ;
        RECT 11.388 0.972 11.42 3.48 ;
  LAYER M3 ;
        RECT 11.388 3.428 11.42 3.46 ;
  LAYER M1 ;
        RECT 11.452 0.972 11.484 3.48 ;
  LAYER M3 ;
        RECT 11.452 0.992 11.484 1.024 ;
  LAYER M1 ;
        RECT 11.516 0.972 11.548 3.48 ;
  LAYER M3 ;
        RECT 11.516 3.428 11.548 3.46 ;
  LAYER M1 ;
        RECT 11.58 0.972 11.612 3.48 ;
  LAYER M3 ;
        RECT 11.58 0.992 11.612 1.024 ;
  LAYER M1 ;
        RECT 11.644 0.972 11.676 3.48 ;
  LAYER M3 ;
        RECT 11.644 3.428 11.676 3.46 ;
  LAYER M1 ;
        RECT 11.708 0.972 11.74 3.48 ;
  LAYER M3 ;
        RECT 11.708 0.992 11.74 1.024 ;
  LAYER M1 ;
        RECT 11.772 0.972 11.804 3.48 ;
  LAYER M3 ;
        RECT 11.772 3.428 11.804 3.46 ;
  LAYER M1 ;
        RECT 11.836 0.972 11.868 3.48 ;
  LAYER M3 ;
        RECT 11.836 0.992 11.868 1.024 ;
  LAYER M1 ;
        RECT 11.9 0.972 11.932 3.48 ;
  LAYER M3 ;
        RECT 11.9 3.428 11.932 3.46 ;
  LAYER M1 ;
        RECT 11.964 0.972 11.996 3.48 ;
  LAYER M3 ;
        RECT 11.964 0.992 11.996 1.024 ;
  LAYER M1 ;
        RECT 12.028 0.972 12.06 3.48 ;
  LAYER M3 ;
        RECT 12.028 3.428 12.06 3.46 ;
  LAYER M1 ;
        RECT 12.092 0.972 12.124 3.48 ;
  LAYER M3 ;
        RECT 12.092 0.992 12.124 1.024 ;
  LAYER M1 ;
        RECT 12.156 0.972 12.188 3.48 ;
  LAYER M3 ;
        RECT 12.156 3.428 12.188 3.46 ;
  LAYER M1 ;
        RECT 12.22 0.972 12.252 3.48 ;
  LAYER M3 ;
        RECT 12.22 0.992 12.252 1.024 ;
  LAYER M1 ;
        RECT 12.284 0.972 12.316 3.48 ;
  LAYER M3 ;
        RECT 12.284 3.428 12.316 3.46 ;
  LAYER M1 ;
        RECT 12.348 0.972 12.38 3.48 ;
  LAYER M3 ;
        RECT 9.98 1.056 10.012 1.088 ;
  LAYER M2 ;
        RECT 12.348 1.12 12.38 1.152 ;
  LAYER M2 ;
        RECT 9.98 1.184 10.012 1.216 ;
  LAYER M2 ;
        RECT 12.348 1.248 12.38 1.28 ;
  LAYER M2 ;
        RECT 9.98 1.312 10.012 1.344 ;
  LAYER M2 ;
        RECT 12.348 1.376 12.38 1.408 ;
  LAYER M2 ;
        RECT 9.98 1.44 10.012 1.472 ;
  LAYER M2 ;
        RECT 12.348 1.504 12.38 1.536 ;
  LAYER M2 ;
        RECT 9.98 1.568 10.012 1.6 ;
  LAYER M2 ;
        RECT 12.348 1.632 12.38 1.664 ;
  LAYER M2 ;
        RECT 9.98 1.696 10.012 1.728 ;
  LAYER M2 ;
        RECT 12.348 1.76 12.38 1.792 ;
  LAYER M2 ;
        RECT 9.98 1.824 10.012 1.856 ;
  LAYER M2 ;
        RECT 12.348 1.888 12.38 1.92 ;
  LAYER M2 ;
        RECT 9.98 1.952 10.012 1.984 ;
  LAYER M2 ;
        RECT 12.348 2.016 12.38 2.048 ;
  LAYER M2 ;
        RECT 9.98 2.08 10.012 2.112 ;
  LAYER M2 ;
        RECT 12.348 2.144 12.38 2.176 ;
  LAYER M2 ;
        RECT 9.98 2.208 10.012 2.24 ;
  LAYER M2 ;
        RECT 12.348 2.272 12.38 2.304 ;
  LAYER M2 ;
        RECT 9.98 2.336 10.012 2.368 ;
  LAYER M2 ;
        RECT 12.348 2.4 12.38 2.432 ;
  LAYER M2 ;
        RECT 9.98 2.464 10.012 2.496 ;
  LAYER M2 ;
        RECT 12.348 2.528 12.38 2.56 ;
  LAYER M2 ;
        RECT 9.98 2.592 10.012 2.624 ;
  LAYER M2 ;
        RECT 12.348 2.656 12.38 2.688 ;
  LAYER M2 ;
        RECT 9.98 2.72 10.012 2.752 ;
  LAYER M2 ;
        RECT 12.348 2.784 12.38 2.816 ;
  LAYER M2 ;
        RECT 9.98 2.848 10.012 2.88 ;
  LAYER M2 ;
        RECT 12.348 2.912 12.38 2.944 ;
  LAYER M2 ;
        RECT 9.98 2.976 10.012 3.008 ;
  LAYER M2 ;
        RECT 12.348 3.04 12.38 3.072 ;
  LAYER M2 ;
        RECT 9.98 3.104 10.012 3.136 ;
  LAYER M2 ;
        RECT 12.348 3.168 12.38 3.2 ;
  LAYER M2 ;
        RECT 9.98 3.232 10.012 3.264 ;
  LAYER M2 ;
        RECT 12.348 3.296 12.38 3.328 ;
  LAYER M2 ;
        RECT 9.932 0.924 12.428 3.528 ;
  LAYER M1 ;
        RECT 9.98 4.08 10.012 6.588 ;
  LAYER M3 ;
        RECT 9.98 6.536 10.012 6.568 ;
  LAYER M1 ;
        RECT 10.044 4.08 10.076 6.588 ;
  LAYER M3 ;
        RECT 10.044 4.1 10.076 4.132 ;
  LAYER M1 ;
        RECT 10.108 4.08 10.14 6.588 ;
  LAYER M3 ;
        RECT 10.108 6.536 10.14 6.568 ;
  LAYER M1 ;
        RECT 10.172 4.08 10.204 6.588 ;
  LAYER M3 ;
        RECT 10.172 4.1 10.204 4.132 ;
  LAYER M1 ;
        RECT 10.236 4.08 10.268 6.588 ;
  LAYER M3 ;
        RECT 10.236 6.536 10.268 6.568 ;
  LAYER M1 ;
        RECT 10.3 4.08 10.332 6.588 ;
  LAYER M3 ;
        RECT 10.3 4.1 10.332 4.132 ;
  LAYER M1 ;
        RECT 10.364 4.08 10.396 6.588 ;
  LAYER M3 ;
        RECT 10.364 6.536 10.396 6.568 ;
  LAYER M1 ;
        RECT 10.428 4.08 10.46 6.588 ;
  LAYER M3 ;
        RECT 10.428 4.1 10.46 4.132 ;
  LAYER M1 ;
        RECT 10.492 4.08 10.524 6.588 ;
  LAYER M3 ;
        RECT 10.492 6.536 10.524 6.568 ;
  LAYER M1 ;
        RECT 10.556 4.08 10.588 6.588 ;
  LAYER M3 ;
        RECT 10.556 4.1 10.588 4.132 ;
  LAYER M1 ;
        RECT 10.62 4.08 10.652 6.588 ;
  LAYER M3 ;
        RECT 10.62 6.536 10.652 6.568 ;
  LAYER M1 ;
        RECT 10.684 4.08 10.716 6.588 ;
  LAYER M3 ;
        RECT 10.684 4.1 10.716 4.132 ;
  LAYER M1 ;
        RECT 10.748 4.08 10.78 6.588 ;
  LAYER M3 ;
        RECT 10.748 6.536 10.78 6.568 ;
  LAYER M1 ;
        RECT 10.812 4.08 10.844 6.588 ;
  LAYER M3 ;
        RECT 10.812 4.1 10.844 4.132 ;
  LAYER M1 ;
        RECT 10.876 4.08 10.908 6.588 ;
  LAYER M3 ;
        RECT 10.876 6.536 10.908 6.568 ;
  LAYER M1 ;
        RECT 10.94 4.08 10.972 6.588 ;
  LAYER M3 ;
        RECT 10.94 4.1 10.972 4.132 ;
  LAYER M1 ;
        RECT 11.004 4.08 11.036 6.588 ;
  LAYER M3 ;
        RECT 11.004 6.536 11.036 6.568 ;
  LAYER M1 ;
        RECT 11.068 4.08 11.1 6.588 ;
  LAYER M3 ;
        RECT 11.068 4.1 11.1 4.132 ;
  LAYER M1 ;
        RECT 11.132 4.08 11.164 6.588 ;
  LAYER M3 ;
        RECT 11.132 6.536 11.164 6.568 ;
  LAYER M1 ;
        RECT 11.196 4.08 11.228 6.588 ;
  LAYER M3 ;
        RECT 11.196 4.1 11.228 4.132 ;
  LAYER M1 ;
        RECT 11.26 4.08 11.292 6.588 ;
  LAYER M3 ;
        RECT 11.26 6.536 11.292 6.568 ;
  LAYER M1 ;
        RECT 11.324 4.08 11.356 6.588 ;
  LAYER M3 ;
        RECT 11.324 4.1 11.356 4.132 ;
  LAYER M1 ;
        RECT 11.388 4.08 11.42 6.588 ;
  LAYER M3 ;
        RECT 11.388 6.536 11.42 6.568 ;
  LAYER M1 ;
        RECT 11.452 4.08 11.484 6.588 ;
  LAYER M3 ;
        RECT 11.452 4.1 11.484 4.132 ;
  LAYER M1 ;
        RECT 11.516 4.08 11.548 6.588 ;
  LAYER M3 ;
        RECT 11.516 6.536 11.548 6.568 ;
  LAYER M1 ;
        RECT 11.58 4.08 11.612 6.588 ;
  LAYER M3 ;
        RECT 11.58 4.1 11.612 4.132 ;
  LAYER M1 ;
        RECT 11.644 4.08 11.676 6.588 ;
  LAYER M3 ;
        RECT 11.644 6.536 11.676 6.568 ;
  LAYER M1 ;
        RECT 11.708 4.08 11.74 6.588 ;
  LAYER M3 ;
        RECT 11.708 4.1 11.74 4.132 ;
  LAYER M1 ;
        RECT 11.772 4.08 11.804 6.588 ;
  LAYER M3 ;
        RECT 11.772 6.536 11.804 6.568 ;
  LAYER M1 ;
        RECT 11.836 4.08 11.868 6.588 ;
  LAYER M3 ;
        RECT 11.836 4.1 11.868 4.132 ;
  LAYER M1 ;
        RECT 11.9 4.08 11.932 6.588 ;
  LAYER M3 ;
        RECT 11.9 6.536 11.932 6.568 ;
  LAYER M1 ;
        RECT 11.964 4.08 11.996 6.588 ;
  LAYER M3 ;
        RECT 11.964 4.1 11.996 4.132 ;
  LAYER M1 ;
        RECT 12.028 4.08 12.06 6.588 ;
  LAYER M3 ;
        RECT 12.028 6.536 12.06 6.568 ;
  LAYER M1 ;
        RECT 12.092 4.08 12.124 6.588 ;
  LAYER M3 ;
        RECT 12.092 4.1 12.124 4.132 ;
  LAYER M1 ;
        RECT 12.156 4.08 12.188 6.588 ;
  LAYER M3 ;
        RECT 12.156 6.536 12.188 6.568 ;
  LAYER M1 ;
        RECT 12.22 4.08 12.252 6.588 ;
  LAYER M3 ;
        RECT 12.22 4.1 12.252 4.132 ;
  LAYER M1 ;
        RECT 12.284 4.08 12.316 6.588 ;
  LAYER M3 ;
        RECT 12.284 6.536 12.316 6.568 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 6.588 ;
  LAYER M3 ;
        RECT 9.98 4.164 10.012 4.196 ;
  LAYER M2 ;
        RECT 12.348 4.228 12.38 4.26 ;
  LAYER M2 ;
        RECT 9.98 4.292 10.012 4.324 ;
  LAYER M2 ;
        RECT 12.348 4.356 12.38 4.388 ;
  LAYER M2 ;
        RECT 9.98 4.42 10.012 4.452 ;
  LAYER M2 ;
        RECT 12.348 4.484 12.38 4.516 ;
  LAYER M2 ;
        RECT 9.98 4.548 10.012 4.58 ;
  LAYER M2 ;
        RECT 12.348 4.612 12.38 4.644 ;
  LAYER M2 ;
        RECT 9.98 4.676 10.012 4.708 ;
  LAYER M2 ;
        RECT 12.348 4.74 12.38 4.772 ;
  LAYER M2 ;
        RECT 9.98 4.804 10.012 4.836 ;
  LAYER M2 ;
        RECT 12.348 4.868 12.38 4.9 ;
  LAYER M2 ;
        RECT 9.98 4.932 10.012 4.964 ;
  LAYER M2 ;
        RECT 12.348 4.996 12.38 5.028 ;
  LAYER M2 ;
        RECT 9.98 5.06 10.012 5.092 ;
  LAYER M2 ;
        RECT 12.348 5.124 12.38 5.156 ;
  LAYER M2 ;
        RECT 9.98 5.188 10.012 5.22 ;
  LAYER M2 ;
        RECT 12.348 5.252 12.38 5.284 ;
  LAYER M2 ;
        RECT 9.98 5.316 10.012 5.348 ;
  LAYER M2 ;
        RECT 12.348 5.38 12.38 5.412 ;
  LAYER M2 ;
        RECT 9.98 5.444 10.012 5.476 ;
  LAYER M2 ;
        RECT 12.348 5.508 12.38 5.54 ;
  LAYER M2 ;
        RECT 9.98 5.572 10.012 5.604 ;
  LAYER M2 ;
        RECT 12.348 5.636 12.38 5.668 ;
  LAYER M2 ;
        RECT 9.98 5.7 10.012 5.732 ;
  LAYER M2 ;
        RECT 12.348 5.764 12.38 5.796 ;
  LAYER M2 ;
        RECT 9.98 5.828 10.012 5.86 ;
  LAYER M2 ;
        RECT 12.348 5.892 12.38 5.924 ;
  LAYER M2 ;
        RECT 9.98 5.956 10.012 5.988 ;
  LAYER M2 ;
        RECT 12.348 6.02 12.38 6.052 ;
  LAYER M2 ;
        RECT 9.98 6.084 10.012 6.116 ;
  LAYER M2 ;
        RECT 12.348 6.148 12.38 6.18 ;
  LAYER M2 ;
        RECT 9.98 6.212 10.012 6.244 ;
  LAYER M2 ;
        RECT 12.348 6.276 12.38 6.308 ;
  LAYER M2 ;
        RECT 9.98 6.34 10.012 6.372 ;
  LAYER M2 ;
        RECT 12.348 6.404 12.38 6.436 ;
  LAYER M2 ;
        RECT 9.932 4.032 12.428 6.636 ;
  LAYER M1 ;
        RECT 9.98 7.188 10.012 9.696 ;
  LAYER M3 ;
        RECT 9.98 9.644 10.012 9.676 ;
  LAYER M1 ;
        RECT 10.044 7.188 10.076 9.696 ;
  LAYER M3 ;
        RECT 10.044 7.208 10.076 7.24 ;
  LAYER M1 ;
        RECT 10.108 7.188 10.14 9.696 ;
  LAYER M3 ;
        RECT 10.108 9.644 10.14 9.676 ;
  LAYER M1 ;
        RECT 10.172 7.188 10.204 9.696 ;
  LAYER M3 ;
        RECT 10.172 7.208 10.204 7.24 ;
  LAYER M1 ;
        RECT 10.236 7.188 10.268 9.696 ;
  LAYER M3 ;
        RECT 10.236 9.644 10.268 9.676 ;
  LAYER M1 ;
        RECT 10.3 7.188 10.332 9.696 ;
  LAYER M3 ;
        RECT 10.3 7.208 10.332 7.24 ;
  LAYER M1 ;
        RECT 10.364 7.188 10.396 9.696 ;
  LAYER M3 ;
        RECT 10.364 9.644 10.396 9.676 ;
  LAYER M1 ;
        RECT 10.428 7.188 10.46 9.696 ;
  LAYER M3 ;
        RECT 10.428 7.208 10.46 7.24 ;
  LAYER M1 ;
        RECT 10.492 7.188 10.524 9.696 ;
  LAYER M3 ;
        RECT 10.492 9.644 10.524 9.676 ;
  LAYER M1 ;
        RECT 10.556 7.188 10.588 9.696 ;
  LAYER M3 ;
        RECT 10.556 7.208 10.588 7.24 ;
  LAYER M1 ;
        RECT 10.62 7.188 10.652 9.696 ;
  LAYER M3 ;
        RECT 10.62 9.644 10.652 9.676 ;
  LAYER M1 ;
        RECT 10.684 7.188 10.716 9.696 ;
  LAYER M3 ;
        RECT 10.684 7.208 10.716 7.24 ;
  LAYER M1 ;
        RECT 10.748 7.188 10.78 9.696 ;
  LAYER M3 ;
        RECT 10.748 9.644 10.78 9.676 ;
  LAYER M1 ;
        RECT 10.812 7.188 10.844 9.696 ;
  LAYER M3 ;
        RECT 10.812 7.208 10.844 7.24 ;
  LAYER M1 ;
        RECT 10.876 7.188 10.908 9.696 ;
  LAYER M3 ;
        RECT 10.876 9.644 10.908 9.676 ;
  LAYER M1 ;
        RECT 10.94 7.188 10.972 9.696 ;
  LAYER M3 ;
        RECT 10.94 7.208 10.972 7.24 ;
  LAYER M1 ;
        RECT 11.004 7.188 11.036 9.696 ;
  LAYER M3 ;
        RECT 11.004 9.644 11.036 9.676 ;
  LAYER M1 ;
        RECT 11.068 7.188 11.1 9.696 ;
  LAYER M3 ;
        RECT 11.068 7.208 11.1 7.24 ;
  LAYER M1 ;
        RECT 11.132 7.188 11.164 9.696 ;
  LAYER M3 ;
        RECT 11.132 9.644 11.164 9.676 ;
  LAYER M1 ;
        RECT 11.196 7.188 11.228 9.696 ;
  LAYER M3 ;
        RECT 11.196 7.208 11.228 7.24 ;
  LAYER M1 ;
        RECT 11.26 7.188 11.292 9.696 ;
  LAYER M3 ;
        RECT 11.26 9.644 11.292 9.676 ;
  LAYER M1 ;
        RECT 11.324 7.188 11.356 9.696 ;
  LAYER M3 ;
        RECT 11.324 7.208 11.356 7.24 ;
  LAYER M1 ;
        RECT 11.388 7.188 11.42 9.696 ;
  LAYER M3 ;
        RECT 11.388 9.644 11.42 9.676 ;
  LAYER M1 ;
        RECT 11.452 7.188 11.484 9.696 ;
  LAYER M3 ;
        RECT 11.452 7.208 11.484 7.24 ;
  LAYER M1 ;
        RECT 11.516 7.188 11.548 9.696 ;
  LAYER M3 ;
        RECT 11.516 9.644 11.548 9.676 ;
  LAYER M1 ;
        RECT 11.58 7.188 11.612 9.696 ;
  LAYER M3 ;
        RECT 11.58 7.208 11.612 7.24 ;
  LAYER M1 ;
        RECT 11.644 7.188 11.676 9.696 ;
  LAYER M3 ;
        RECT 11.644 9.644 11.676 9.676 ;
  LAYER M1 ;
        RECT 11.708 7.188 11.74 9.696 ;
  LAYER M3 ;
        RECT 11.708 7.208 11.74 7.24 ;
  LAYER M1 ;
        RECT 11.772 7.188 11.804 9.696 ;
  LAYER M3 ;
        RECT 11.772 9.644 11.804 9.676 ;
  LAYER M1 ;
        RECT 11.836 7.188 11.868 9.696 ;
  LAYER M3 ;
        RECT 11.836 7.208 11.868 7.24 ;
  LAYER M1 ;
        RECT 11.9 7.188 11.932 9.696 ;
  LAYER M3 ;
        RECT 11.9 9.644 11.932 9.676 ;
  LAYER M1 ;
        RECT 11.964 7.188 11.996 9.696 ;
  LAYER M3 ;
        RECT 11.964 7.208 11.996 7.24 ;
  LAYER M1 ;
        RECT 12.028 7.188 12.06 9.696 ;
  LAYER M3 ;
        RECT 12.028 9.644 12.06 9.676 ;
  LAYER M1 ;
        RECT 12.092 7.188 12.124 9.696 ;
  LAYER M3 ;
        RECT 12.092 7.208 12.124 7.24 ;
  LAYER M1 ;
        RECT 12.156 7.188 12.188 9.696 ;
  LAYER M3 ;
        RECT 12.156 9.644 12.188 9.676 ;
  LAYER M1 ;
        RECT 12.22 7.188 12.252 9.696 ;
  LAYER M3 ;
        RECT 12.22 7.208 12.252 7.24 ;
  LAYER M1 ;
        RECT 12.284 7.188 12.316 9.696 ;
  LAYER M3 ;
        RECT 12.284 9.644 12.316 9.676 ;
  LAYER M1 ;
        RECT 12.348 7.188 12.38 9.696 ;
  LAYER M3 ;
        RECT 9.98 7.272 10.012 7.304 ;
  LAYER M2 ;
        RECT 12.348 7.336 12.38 7.368 ;
  LAYER M2 ;
        RECT 9.98 7.4 10.012 7.432 ;
  LAYER M2 ;
        RECT 12.348 7.464 12.38 7.496 ;
  LAYER M2 ;
        RECT 9.98 7.528 10.012 7.56 ;
  LAYER M2 ;
        RECT 12.348 7.592 12.38 7.624 ;
  LAYER M2 ;
        RECT 9.98 7.656 10.012 7.688 ;
  LAYER M2 ;
        RECT 12.348 7.72 12.38 7.752 ;
  LAYER M2 ;
        RECT 9.98 7.784 10.012 7.816 ;
  LAYER M2 ;
        RECT 12.348 7.848 12.38 7.88 ;
  LAYER M2 ;
        RECT 9.98 7.912 10.012 7.944 ;
  LAYER M2 ;
        RECT 12.348 7.976 12.38 8.008 ;
  LAYER M2 ;
        RECT 9.98 8.04 10.012 8.072 ;
  LAYER M2 ;
        RECT 12.348 8.104 12.38 8.136 ;
  LAYER M2 ;
        RECT 9.98 8.168 10.012 8.2 ;
  LAYER M2 ;
        RECT 12.348 8.232 12.38 8.264 ;
  LAYER M2 ;
        RECT 9.98 8.296 10.012 8.328 ;
  LAYER M2 ;
        RECT 12.348 8.36 12.38 8.392 ;
  LAYER M2 ;
        RECT 9.98 8.424 10.012 8.456 ;
  LAYER M2 ;
        RECT 12.348 8.488 12.38 8.52 ;
  LAYER M2 ;
        RECT 9.98 8.552 10.012 8.584 ;
  LAYER M2 ;
        RECT 12.348 8.616 12.38 8.648 ;
  LAYER M2 ;
        RECT 9.98 8.68 10.012 8.712 ;
  LAYER M2 ;
        RECT 12.348 8.744 12.38 8.776 ;
  LAYER M2 ;
        RECT 9.98 8.808 10.012 8.84 ;
  LAYER M2 ;
        RECT 12.348 8.872 12.38 8.904 ;
  LAYER M2 ;
        RECT 9.98 8.936 10.012 8.968 ;
  LAYER M2 ;
        RECT 12.348 9 12.38 9.032 ;
  LAYER M2 ;
        RECT 9.98 9.064 10.012 9.096 ;
  LAYER M2 ;
        RECT 12.348 9.128 12.38 9.16 ;
  LAYER M2 ;
        RECT 9.98 9.192 10.012 9.224 ;
  LAYER M2 ;
        RECT 12.348 9.256 12.38 9.288 ;
  LAYER M2 ;
        RECT 9.98 9.32 10.012 9.352 ;
  LAYER M2 ;
        RECT 12.348 9.384 12.38 9.416 ;
  LAYER M2 ;
        RECT 9.98 9.448 10.012 9.48 ;
  LAYER M2 ;
        RECT 12.348 9.512 12.38 9.544 ;
  LAYER M2 ;
        RECT 9.932 7.14 12.428 9.744 ;
  LAYER M1 ;
        RECT 9.98 10.296 10.012 12.804 ;
  LAYER M3 ;
        RECT 9.98 12.752 10.012 12.784 ;
  LAYER M1 ;
        RECT 10.044 10.296 10.076 12.804 ;
  LAYER M3 ;
        RECT 10.044 10.316 10.076 10.348 ;
  LAYER M1 ;
        RECT 10.108 10.296 10.14 12.804 ;
  LAYER M3 ;
        RECT 10.108 12.752 10.14 12.784 ;
  LAYER M1 ;
        RECT 10.172 10.296 10.204 12.804 ;
  LAYER M3 ;
        RECT 10.172 10.316 10.204 10.348 ;
  LAYER M1 ;
        RECT 10.236 10.296 10.268 12.804 ;
  LAYER M3 ;
        RECT 10.236 12.752 10.268 12.784 ;
  LAYER M1 ;
        RECT 10.3 10.296 10.332 12.804 ;
  LAYER M3 ;
        RECT 10.3 10.316 10.332 10.348 ;
  LAYER M1 ;
        RECT 10.364 10.296 10.396 12.804 ;
  LAYER M3 ;
        RECT 10.364 12.752 10.396 12.784 ;
  LAYER M1 ;
        RECT 10.428 10.296 10.46 12.804 ;
  LAYER M3 ;
        RECT 10.428 10.316 10.46 10.348 ;
  LAYER M1 ;
        RECT 10.492 10.296 10.524 12.804 ;
  LAYER M3 ;
        RECT 10.492 12.752 10.524 12.784 ;
  LAYER M1 ;
        RECT 10.556 10.296 10.588 12.804 ;
  LAYER M3 ;
        RECT 10.556 10.316 10.588 10.348 ;
  LAYER M1 ;
        RECT 10.62 10.296 10.652 12.804 ;
  LAYER M3 ;
        RECT 10.62 12.752 10.652 12.784 ;
  LAYER M1 ;
        RECT 10.684 10.296 10.716 12.804 ;
  LAYER M3 ;
        RECT 10.684 10.316 10.716 10.348 ;
  LAYER M1 ;
        RECT 10.748 10.296 10.78 12.804 ;
  LAYER M3 ;
        RECT 10.748 12.752 10.78 12.784 ;
  LAYER M1 ;
        RECT 10.812 10.296 10.844 12.804 ;
  LAYER M3 ;
        RECT 10.812 10.316 10.844 10.348 ;
  LAYER M1 ;
        RECT 10.876 10.296 10.908 12.804 ;
  LAYER M3 ;
        RECT 10.876 12.752 10.908 12.784 ;
  LAYER M1 ;
        RECT 10.94 10.296 10.972 12.804 ;
  LAYER M3 ;
        RECT 10.94 10.316 10.972 10.348 ;
  LAYER M1 ;
        RECT 11.004 10.296 11.036 12.804 ;
  LAYER M3 ;
        RECT 11.004 12.752 11.036 12.784 ;
  LAYER M1 ;
        RECT 11.068 10.296 11.1 12.804 ;
  LAYER M3 ;
        RECT 11.068 10.316 11.1 10.348 ;
  LAYER M1 ;
        RECT 11.132 10.296 11.164 12.804 ;
  LAYER M3 ;
        RECT 11.132 12.752 11.164 12.784 ;
  LAYER M1 ;
        RECT 11.196 10.296 11.228 12.804 ;
  LAYER M3 ;
        RECT 11.196 10.316 11.228 10.348 ;
  LAYER M1 ;
        RECT 11.26 10.296 11.292 12.804 ;
  LAYER M3 ;
        RECT 11.26 12.752 11.292 12.784 ;
  LAYER M1 ;
        RECT 11.324 10.296 11.356 12.804 ;
  LAYER M3 ;
        RECT 11.324 10.316 11.356 10.348 ;
  LAYER M1 ;
        RECT 11.388 10.296 11.42 12.804 ;
  LAYER M3 ;
        RECT 11.388 12.752 11.42 12.784 ;
  LAYER M1 ;
        RECT 11.452 10.296 11.484 12.804 ;
  LAYER M3 ;
        RECT 11.452 10.316 11.484 10.348 ;
  LAYER M1 ;
        RECT 11.516 10.296 11.548 12.804 ;
  LAYER M3 ;
        RECT 11.516 12.752 11.548 12.784 ;
  LAYER M1 ;
        RECT 11.58 10.296 11.612 12.804 ;
  LAYER M3 ;
        RECT 11.58 10.316 11.612 10.348 ;
  LAYER M1 ;
        RECT 11.644 10.296 11.676 12.804 ;
  LAYER M3 ;
        RECT 11.644 12.752 11.676 12.784 ;
  LAYER M1 ;
        RECT 11.708 10.296 11.74 12.804 ;
  LAYER M3 ;
        RECT 11.708 10.316 11.74 10.348 ;
  LAYER M1 ;
        RECT 11.772 10.296 11.804 12.804 ;
  LAYER M3 ;
        RECT 11.772 12.752 11.804 12.784 ;
  LAYER M1 ;
        RECT 11.836 10.296 11.868 12.804 ;
  LAYER M3 ;
        RECT 11.836 10.316 11.868 10.348 ;
  LAYER M1 ;
        RECT 11.9 10.296 11.932 12.804 ;
  LAYER M3 ;
        RECT 11.9 12.752 11.932 12.784 ;
  LAYER M1 ;
        RECT 11.964 10.296 11.996 12.804 ;
  LAYER M3 ;
        RECT 11.964 10.316 11.996 10.348 ;
  LAYER M1 ;
        RECT 12.028 10.296 12.06 12.804 ;
  LAYER M3 ;
        RECT 12.028 12.752 12.06 12.784 ;
  LAYER M1 ;
        RECT 12.092 10.296 12.124 12.804 ;
  LAYER M3 ;
        RECT 12.092 10.316 12.124 10.348 ;
  LAYER M1 ;
        RECT 12.156 10.296 12.188 12.804 ;
  LAYER M3 ;
        RECT 12.156 12.752 12.188 12.784 ;
  LAYER M1 ;
        RECT 12.22 10.296 12.252 12.804 ;
  LAYER M3 ;
        RECT 12.22 10.316 12.252 10.348 ;
  LAYER M1 ;
        RECT 12.284 10.296 12.316 12.804 ;
  LAYER M3 ;
        RECT 12.284 12.752 12.316 12.784 ;
  LAYER M1 ;
        RECT 12.348 10.296 12.38 12.804 ;
  LAYER M3 ;
        RECT 9.98 10.38 10.012 10.412 ;
  LAYER M2 ;
        RECT 12.348 10.444 12.38 10.476 ;
  LAYER M2 ;
        RECT 9.98 10.508 10.012 10.54 ;
  LAYER M2 ;
        RECT 12.348 10.572 12.38 10.604 ;
  LAYER M2 ;
        RECT 9.98 10.636 10.012 10.668 ;
  LAYER M2 ;
        RECT 12.348 10.7 12.38 10.732 ;
  LAYER M2 ;
        RECT 9.98 10.764 10.012 10.796 ;
  LAYER M2 ;
        RECT 12.348 10.828 12.38 10.86 ;
  LAYER M2 ;
        RECT 9.98 10.892 10.012 10.924 ;
  LAYER M2 ;
        RECT 12.348 10.956 12.38 10.988 ;
  LAYER M2 ;
        RECT 9.98 11.02 10.012 11.052 ;
  LAYER M2 ;
        RECT 12.348 11.084 12.38 11.116 ;
  LAYER M2 ;
        RECT 9.98 11.148 10.012 11.18 ;
  LAYER M2 ;
        RECT 12.348 11.212 12.38 11.244 ;
  LAYER M2 ;
        RECT 9.98 11.276 10.012 11.308 ;
  LAYER M2 ;
        RECT 12.348 11.34 12.38 11.372 ;
  LAYER M2 ;
        RECT 9.98 11.404 10.012 11.436 ;
  LAYER M2 ;
        RECT 12.348 11.468 12.38 11.5 ;
  LAYER M2 ;
        RECT 9.98 11.532 10.012 11.564 ;
  LAYER M2 ;
        RECT 12.348 11.596 12.38 11.628 ;
  LAYER M2 ;
        RECT 9.98 11.66 10.012 11.692 ;
  LAYER M2 ;
        RECT 12.348 11.724 12.38 11.756 ;
  LAYER M2 ;
        RECT 9.98 11.788 10.012 11.82 ;
  LAYER M2 ;
        RECT 12.348 11.852 12.38 11.884 ;
  LAYER M2 ;
        RECT 9.98 11.916 10.012 11.948 ;
  LAYER M2 ;
        RECT 12.348 11.98 12.38 12.012 ;
  LAYER M2 ;
        RECT 9.98 12.044 10.012 12.076 ;
  LAYER M2 ;
        RECT 12.348 12.108 12.38 12.14 ;
  LAYER M2 ;
        RECT 9.98 12.172 10.012 12.204 ;
  LAYER M2 ;
        RECT 12.348 12.236 12.38 12.268 ;
  LAYER M2 ;
        RECT 9.98 12.3 10.012 12.332 ;
  LAYER M2 ;
        RECT 12.348 12.364 12.38 12.396 ;
  LAYER M2 ;
        RECT 9.98 12.428 10.012 12.46 ;
  LAYER M2 ;
        RECT 12.348 12.492 12.38 12.524 ;
  LAYER M2 ;
        RECT 9.98 12.556 10.012 12.588 ;
  LAYER M2 ;
        RECT 12.348 12.62 12.38 12.652 ;
  LAYER M2 ;
        RECT 9.932 10.248 12.428 12.852 ;
  LAYER M1 ;
        RECT 9.98 13.404 10.012 15.912 ;
  LAYER M3 ;
        RECT 9.98 15.86 10.012 15.892 ;
  LAYER M1 ;
        RECT 10.044 13.404 10.076 15.912 ;
  LAYER M3 ;
        RECT 10.044 13.424 10.076 13.456 ;
  LAYER M1 ;
        RECT 10.108 13.404 10.14 15.912 ;
  LAYER M3 ;
        RECT 10.108 15.86 10.14 15.892 ;
  LAYER M1 ;
        RECT 10.172 13.404 10.204 15.912 ;
  LAYER M3 ;
        RECT 10.172 13.424 10.204 13.456 ;
  LAYER M1 ;
        RECT 10.236 13.404 10.268 15.912 ;
  LAYER M3 ;
        RECT 10.236 15.86 10.268 15.892 ;
  LAYER M1 ;
        RECT 10.3 13.404 10.332 15.912 ;
  LAYER M3 ;
        RECT 10.3 13.424 10.332 13.456 ;
  LAYER M1 ;
        RECT 10.364 13.404 10.396 15.912 ;
  LAYER M3 ;
        RECT 10.364 15.86 10.396 15.892 ;
  LAYER M1 ;
        RECT 10.428 13.404 10.46 15.912 ;
  LAYER M3 ;
        RECT 10.428 13.424 10.46 13.456 ;
  LAYER M1 ;
        RECT 10.492 13.404 10.524 15.912 ;
  LAYER M3 ;
        RECT 10.492 15.86 10.524 15.892 ;
  LAYER M1 ;
        RECT 10.556 13.404 10.588 15.912 ;
  LAYER M3 ;
        RECT 10.556 13.424 10.588 13.456 ;
  LAYER M1 ;
        RECT 10.62 13.404 10.652 15.912 ;
  LAYER M3 ;
        RECT 10.62 15.86 10.652 15.892 ;
  LAYER M1 ;
        RECT 10.684 13.404 10.716 15.912 ;
  LAYER M3 ;
        RECT 10.684 13.424 10.716 13.456 ;
  LAYER M1 ;
        RECT 10.748 13.404 10.78 15.912 ;
  LAYER M3 ;
        RECT 10.748 15.86 10.78 15.892 ;
  LAYER M1 ;
        RECT 10.812 13.404 10.844 15.912 ;
  LAYER M3 ;
        RECT 10.812 13.424 10.844 13.456 ;
  LAYER M1 ;
        RECT 10.876 13.404 10.908 15.912 ;
  LAYER M3 ;
        RECT 10.876 15.86 10.908 15.892 ;
  LAYER M1 ;
        RECT 10.94 13.404 10.972 15.912 ;
  LAYER M3 ;
        RECT 10.94 13.424 10.972 13.456 ;
  LAYER M1 ;
        RECT 11.004 13.404 11.036 15.912 ;
  LAYER M3 ;
        RECT 11.004 15.86 11.036 15.892 ;
  LAYER M1 ;
        RECT 11.068 13.404 11.1 15.912 ;
  LAYER M3 ;
        RECT 11.068 13.424 11.1 13.456 ;
  LAYER M1 ;
        RECT 11.132 13.404 11.164 15.912 ;
  LAYER M3 ;
        RECT 11.132 15.86 11.164 15.892 ;
  LAYER M1 ;
        RECT 11.196 13.404 11.228 15.912 ;
  LAYER M3 ;
        RECT 11.196 13.424 11.228 13.456 ;
  LAYER M1 ;
        RECT 11.26 13.404 11.292 15.912 ;
  LAYER M3 ;
        RECT 11.26 15.86 11.292 15.892 ;
  LAYER M1 ;
        RECT 11.324 13.404 11.356 15.912 ;
  LAYER M3 ;
        RECT 11.324 13.424 11.356 13.456 ;
  LAYER M1 ;
        RECT 11.388 13.404 11.42 15.912 ;
  LAYER M3 ;
        RECT 11.388 15.86 11.42 15.892 ;
  LAYER M1 ;
        RECT 11.452 13.404 11.484 15.912 ;
  LAYER M3 ;
        RECT 11.452 13.424 11.484 13.456 ;
  LAYER M1 ;
        RECT 11.516 13.404 11.548 15.912 ;
  LAYER M3 ;
        RECT 11.516 15.86 11.548 15.892 ;
  LAYER M1 ;
        RECT 11.58 13.404 11.612 15.912 ;
  LAYER M3 ;
        RECT 11.58 13.424 11.612 13.456 ;
  LAYER M1 ;
        RECT 11.644 13.404 11.676 15.912 ;
  LAYER M3 ;
        RECT 11.644 15.86 11.676 15.892 ;
  LAYER M1 ;
        RECT 11.708 13.404 11.74 15.912 ;
  LAYER M3 ;
        RECT 11.708 13.424 11.74 13.456 ;
  LAYER M1 ;
        RECT 11.772 13.404 11.804 15.912 ;
  LAYER M3 ;
        RECT 11.772 15.86 11.804 15.892 ;
  LAYER M1 ;
        RECT 11.836 13.404 11.868 15.912 ;
  LAYER M3 ;
        RECT 11.836 13.424 11.868 13.456 ;
  LAYER M1 ;
        RECT 11.9 13.404 11.932 15.912 ;
  LAYER M3 ;
        RECT 11.9 15.86 11.932 15.892 ;
  LAYER M1 ;
        RECT 11.964 13.404 11.996 15.912 ;
  LAYER M3 ;
        RECT 11.964 13.424 11.996 13.456 ;
  LAYER M1 ;
        RECT 12.028 13.404 12.06 15.912 ;
  LAYER M3 ;
        RECT 12.028 15.86 12.06 15.892 ;
  LAYER M1 ;
        RECT 12.092 13.404 12.124 15.912 ;
  LAYER M3 ;
        RECT 12.092 13.424 12.124 13.456 ;
  LAYER M1 ;
        RECT 12.156 13.404 12.188 15.912 ;
  LAYER M3 ;
        RECT 12.156 15.86 12.188 15.892 ;
  LAYER M1 ;
        RECT 12.22 13.404 12.252 15.912 ;
  LAYER M3 ;
        RECT 12.22 13.424 12.252 13.456 ;
  LAYER M1 ;
        RECT 12.284 13.404 12.316 15.912 ;
  LAYER M3 ;
        RECT 12.284 15.86 12.316 15.892 ;
  LAYER M1 ;
        RECT 12.348 13.404 12.38 15.912 ;
  LAYER M3 ;
        RECT 9.98 13.488 10.012 13.52 ;
  LAYER M2 ;
        RECT 12.348 13.552 12.38 13.584 ;
  LAYER M2 ;
        RECT 9.98 13.616 10.012 13.648 ;
  LAYER M2 ;
        RECT 12.348 13.68 12.38 13.712 ;
  LAYER M2 ;
        RECT 9.98 13.744 10.012 13.776 ;
  LAYER M2 ;
        RECT 12.348 13.808 12.38 13.84 ;
  LAYER M2 ;
        RECT 9.98 13.872 10.012 13.904 ;
  LAYER M2 ;
        RECT 12.348 13.936 12.38 13.968 ;
  LAYER M2 ;
        RECT 9.98 14 10.012 14.032 ;
  LAYER M2 ;
        RECT 12.348 14.064 12.38 14.096 ;
  LAYER M2 ;
        RECT 9.98 14.128 10.012 14.16 ;
  LAYER M2 ;
        RECT 12.348 14.192 12.38 14.224 ;
  LAYER M2 ;
        RECT 9.98 14.256 10.012 14.288 ;
  LAYER M2 ;
        RECT 12.348 14.32 12.38 14.352 ;
  LAYER M2 ;
        RECT 9.98 14.384 10.012 14.416 ;
  LAYER M2 ;
        RECT 12.348 14.448 12.38 14.48 ;
  LAYER M2 ;
        RECT 9.98 14.512 10.012 14.544 ;
  LAYER M2 ;
        RECT 12.348 14.576 12.38 14.608 ;
  LAYER M2 ;
        RECT 9.98 14.64 10.012 14.672 ;
  LAYER M2 ;
        RECT 12.348 14.704 12.38 14.736 ;
  LAYER M2 ;
        RECT 9.98 14.768 10.012 14.8 ;
  LAYER M2 ;
        RECT 12.348 14.832 12.38 14.864 ;
  LAYER M2 ;
        RECT 9.98 14.896 10.012 14.928 ;
  LAYER M2 ;
        RECT 12.348 14.96 12.38 14.992 ;
  LAYER M2 ;
        RECT 9.98 15.024 10.012 15.056 ;
  LAYER M2 ;
        RECT 12.348 15.088 12.38 15.12 ;
  LAYER M2 ;
        RECT 9.98 15.152 10.012 15.184 ;
  LAYER M2 ;
        RECT 12.348 15.216 12.38 15.248 ;
  LAYER M2 ;
        RECT 9.98 15.28 10.012 15.312 ;
  LAYER M2 ;
        RECT 12.348 15.344 12.38 15.376 ;
  LAYER M2 ;
        RECT 9.98 15.408 10.012 15.44 ;
  LAYER M2 ;
        RECT 12.348 15.472 12.38 15.504 ;
  LAYER M2 ;
        RECT 9.98 15.536 10.012 15.568 ;
  LAYER M2 ;
        RECT 12.348 15.6 12.38 15.632 ;
  LAYER M2 ;
        RECT 9.98 15.664 10.012 15.696 ;
  LAYER M2 ;
        RECT 12.348 15.728 12.38 15.76 ;
  LAYER M2 ;
        RECT 9.932 13.356 12.428 15.96 ;
  LAYER M1 ;
        RECT 9.98 16.512 10.012 19.02 ;
  LAYER M3 ;
        RECT 9.98 18.968 10.012 19 ;
  LAYER M1 ;
        RECT 10.044 16.512 10.076 19.02 ;
  LAYER M3 ;
        RECT 10.044 16.532 10.076 16.564 ;
  LAYER M1 ;
        RECT 10.108 16.512 10.14 19.02 ;
  LAYER M3 ;
        RECT 10.108 18.968 10.14 19 ;
  LAYER M1 ;
        RECT 10.172 16.512 10.204 19.02 ;
  LAYER M3 ;
        RECT 10.172 16.532 10.204 16.564 ;
  LAYER M1 ;
        RECT 10.236 16.512 10.268 19.02 ;
  LAYER M3 ;
        RECT 10.236 18.968 10.268 19 ;
  LAYER M1 ;
        RECT 10.3 16.512 10.332 19.02 ;
  LAYER M3 ;
        RECT 10.3 16.532 10.332 16.564 ;
  LAYER M1 ;
        RECT 10.364 16.512 10.396 19.02 ;
  LAYER M3 ;
        RECT 10.364 18.968 10.396 19 ;
  LAYER M1 ;
        RECT 10.428 16.512 10.46 19.02 ;
  LAYER M3 ;
        RECT 10.428 16.532 10.46 16.564 ;
  LAYER M1 ;
        RECT 10.492 16.512 10.524 19.02 ;
  LAYER M3 ;
        RECT 10.492 18.968 10.524 19 ;
  LAYER M1 ;
        RECT 10.556 16.512 10.588 19.02 ;
  LAYER M3 ;
        RECT 10.556 16.532 10.588 16.564 ;
  LAYER M1 ;
        RECT 10.62 16.512 10.652 19.02 ;
  LAYER M3 ;
        RECT 10.62 18.968 10.652 19 ;
  LAYER M1 ;
        RECT 10.684 16.512 10.716 19.02 ;
  LAYER M3 ;
        RECT 10.684 16.532 10.716 16.564 ;
  LAYER M1 ;
        RECT 10.748 16.512 10.78 19.02 ;
  LAYER M3 ;
        RECT 10.748 18.968 10.78 19 ;
  LAYER M1 ;
        RECT 10.812 16.512 10.844 19.02 ;
  LAYER M3 ;
        RECT 10.812 16.532 10.844 16.564 ;
  LAYER M1 ;
        RECT 10.876 16.512 10.908 19.02 ;
  LAYER M3 ;
        RECT 10.876 18.968 10.908 19 ;
  LAYER M1 ;
        RECT 10.94 16.512 10.972 19.02 ;
  LAYER M3 ;
        RECT 10.94 16.532 10.972 16.564 ;
  LAYER M1 ;
        RECT 11.004 16.512 11.036 19.02 ;
  LAYER M3 ;
        RECT 11.004 18.968 11.036 19 ;
  LAYER M1 ;
        RECT 11.068 16.512 11.1 19.02 ;
  LAYER M3 ;
        RECT 11.068 16.532 11.1 16.564 ;
  LAYER M1 ;
        RECT 11.132 16.512 11.164 19.02 ;
  LAYER M3 ;
        RECT 11.132 18.968 11.164 19 ;
  LAYER M1 ;
        RECT 11.196 16.512 11.228 19.02 ;
  LAYER M3 ;
        RECT 11.196 16.532 11.228 16.564 ;
  LAYER M1 ;
        RECT 11.26 16.512 11.292 19.02 ;
  LAYER M3 ;
        RECT 11.26 18.968 11.292 19 ;
  LAYER M1 ;
        RECT 11.324 16.512 11.356 19.02 ;
  LAYER M3 ;
        RECT 11.324 16.532 11.356 16.564 ;
  LAYER M1 ;
        RECT 11.388 16.512 11.42 19.02 ;
  LAYER M3 ;
        RECT 11.388 18.968 11.42 19 ;
  LAYER M1 ;
        RECT 11.452 16.512 11.484 19.02 ;
  LAYER M3 ;
        RECT 11.452 16.532 11.484 16.564 ;
  LAYER M1 ;
        RECT 11.516 16.512 11.548 19.02 ;
  LAYER M3 ;
        RECT 11.516 18.968 11.548 19 ;
  LAYER M1 ;
        RECT 11.58 16.512 11.612 19.02 ;
  LAYER M3 ;
        RECT 11.58 16.532 11.612 16.564 ;
  LAYER M1 ;
        RECT 11.644 16.512 11.676 19.02 ;
  LAYER M3 ;
        RECT 11.644 18.968 11.676 19 ;
  LAYER M1 ;
        RECT 11.708 16.512 11.74 19.02 ;
  LAYER M3 ;
        RECT 11.708 16.532 11.74 16.564 ;
  LAYER M1 ;
        RECT 11.772 16.512 11.804 19.02 ;
  LAYER M3 ;
        RECT 11.772 18.968 11.804 19 ;
  LAYER M1 ;
        RECT 11.836 16.512 11.868 19.02 ;
  LAYER M3 ;
        RECT 11.836 16.532 11.868 16.564 ;
  LAYER M1 ;
        RECT 11.9 16.512 11.932 19.02 ;
  LAYER M3 ;
        RECT 11.9 18.968 11.932 19 ;
  LAYER M1 ;
        RECT 11.964 16.512 11.996 19.02 ;
  LAYER M3 ;
        RECT 11.964 16.532 11.996 16.564 ;
  LAYER M1 ;
        RECT 12.028 16.512 12.06 19.02 ;
  LAYER M3 ;
        RECT 12.028 18.968 12.06 19 ;
  LAYER M1 ;
        RECT 12.092 16.512 12.124 19.02 ;
  LAYER M3 ;
        RECT 12.092 16.532 12.124 16.564 ;
  LAYER M1 ;
        RECT 12.156 16.512 12.188 19.02 ;
  LAYER M3 ;
        RECT 12.156 18.968 12.188 19 ;
  LAYER M1 ;
        RECT 12.22 16.512 12.252 19.02 ;
  LAYER M3 ;
        RECT 12.22 16.532 12.252 16.564 ;
  LAYER M1 ;
        RECT 12.284 16.512 12.316 19.02 ;
  LAYER M3 ;
        RECT 12.284 18.968 12.316 19 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 19.02 ;
  LAYER M3 ;
        RECT 9.98 16.596 10.012 16.628 ;
  LAYER M2 ;
        RECT 12.348 16.66 12.38 16.692 ;
  LAYER M2 ;
        RECT 9.98 16.724 10.012 16.756 ;
  LAYER M2 ;
        RECT 12.348 16.788 12.38 16.82 ;
  LAYER M2 ;
        RECT 9.98 16.852 10.012 16.884 ;
  LAYER M2 ;
        RECT 12.348 16.916 12.38 16.948 ;
  LAYER M2 ;
        RECT 9.98 16.98 10.012 17.012 ;
  LAYER M2 ;
        RECT 12.348 17.044 12.38 17.076 ;
  LAYER M2 ;
        RECT 9.98 17.108 10.012 17.14 ;
  LAYER M2 ;
        RECT 12.348 17.172 12.38 17.204 ;
  LAYER M2 ;
        RECT 9.98 17.236 10.012 17.268 ;
  LAYER M2 ;
        RECT 12.348 17.3 12.38 17.332 ;
  LAYER M2 ;
        RECT 9.98 17.364 10.012 17.396 ;
  LAYER M2 ;
        RECT 12.348 17.428 12.38 17.46 ;
  LAYER M2 ;
        RECT 9.98 17.492 10.012 17.524 ;
  LAYER M2 ;
        RECT 12.348 17.556 12.38 17.588 ;
  LAYER M2 ;
        RECT 9.98 17.62 10.012 17.652 ;
  LAYER M2 ;
        RECT 12.348 17.684 12.38 17.716 ;
  LAYER M2 ;
        RECT 9.98 17.748 10.012 17.78 ;
  LAYER M2 ;
        RECT 12.348 17.812 12.38 17.844 ;
  LAYER M2 ;
        RECT 9.98 17.876 10.012 17.908 ;
  LAYER M2 ;
        RECT 12.348 17.94 12.38 17.972 ;
  LAYER M2 ;
        RECT 9.98 18.004 10.012 18.036 ;
  LAYER M2 ;
        RECT 12.348 18.068 12.38 18.1 ;
  LAYER M2 ;
        RECT 9.98 18.132 10.012 18.164 ;
  LAYER M2 ;
        RECT 12.348 18.196 12.38 18.228 ;
  LAYER M2 ;
        RECT 9.98 18.26 10.012 18.292 ;
  LAYER M2 ;
        RECT 12.348 18.324 12.38 18.356 ;
  LAYER M2 ;
        RECT 9.98 18.388 10.012 18.42 ;
  LAYER M2 ;
        RECT 12.348 18.452 12.38 18.484 ;
  LAYER M2 ;
        RECT 9.98 18.516 10.012 18.548 ;
  LAYER M2 ;
        RECT 12.348 18.58 12.38 18.612 ;
  LAYER M2 ;
        RECT 9.98 18.644 10.012 18.676 ;
  LAYER M2 ;
        RECT 12.348 18.708 12.38 18.74 ;
  LAYER M2 ;
        RECT 9.98 18.772 10.012 18.804 ;
  LAYER M2 ;
        RECT 12.348 18.836 12.38 18.868 ;
  LAYER M2 ;
        RECT 9.932 16.464 12.428 19.068 ;
  LAYER M1 ;
        RECT 9.98 19.62 10.012 22.128 ;
  LAYER M3 ;
        RECT 9.98 22.076 10.012 22.108 ;
  LAYER M1 ;
        RECT 10.044 19.62 10.076 22.128 ;
  LAYER M3 ;
        RECT 10.044 19.64 10.076 19.672 ;
  LAYER M1 ;
        RECT 10.108 19.62 10.14 22.128 ;
  LAYER M3 ;
        RECT 10.108 22.076 10.14 22.108 ;
  LAYER M1 ;
        RECT 10.172 19.62 10.204 22.128 ;
  LAYER M3 ;
        RECT 10.172 19.64 10.204 19.672 ;
  LAYER M1 ;
        RECT 10.236 19.62 10.268 22.128 ;
  LAYER M3 ;
        RECT 10.236 22.076 10.268 22.108 ;
  LAYER M1 ;
        RECT 10.3 19.62 10.332 22.128 ;
  LAYER M3 ;
        RECT 10.3 19.64 10.332 19.672 ;
  LAYER M1 ;
        RECT 10.364 19.62 10.396 22.128 ;
  LAYER M3 ;
        RECT 10.364 22.076 10.396 22.108 ;
  LAYER M1 ;
        RECT 10.428 19.62 10.46 22.128 ;
  LAYER M3 ;
        RECT 10.428 19.64 10.46 19.672 ;
  LAYER M1 ;
        RECT 10.492 19.62 10.524 22.128 ;
  LAYER M3 ;
        RECT 10.492 22.076 10.524 22.108 ;
  LAYER M1 ;
        RECT 10.556 19.62 10.588 22.128 ;
  LAYER M3 ;
        RECT 10.556 19.64 10.588 19.672 ;
  LAYER M1 ;
        RECT 10.62 19.62 10.652 22.128 ;
  LAYER M3 ;
        RECT 10.62 22.076 10.652 22.108 ;
  LAYER M1 ;
        RECT 10.684 19.62 10.716 22.128 ;
  LAYER M3 ;
        RECT 10.684 19.64 10.716 19.672 ;
  LAYER M1 ;
        RECT 10.748 19.62 10.78 22.128 ;
  LAYER M3 ;
        RECT 10.748 22.076 10.78 22.108 ;
  LAYER M1 ;
        RECT 10.812 19.62 10.844 22.128 ;
  LAYER M3 ;
        RECT 10.812 19.64 10.844 19.672 ;
  LAYER M1 ;
        RECT 10.876 19.62 10.908 22.128 ;
  LAYER M3 ;
        RECT 10.876 22.076 10.908 22.108 ;
  LAYER M1 ;
        RECT 10.94 19.62 10.972 22.128 ;
  LAYER M3 ;
        RECT 10.94 19.64 10.972 19.672 ;
  LAYER M1 ;
        RECT 11.004 19.62 11.036 22.128 ;
  LAYER M3 ;
        RECT 11.004 22.076 11.036 22.108 ;
  LAYER M1 ;
        RECT 11.068 19.62 11.1 22.128 ;
  LAYER M3 ;
        RECT 11.068 19.64 11.1 19.672 ;
  LAYER M1 ;
        RECT 11.132 19.62 11.164 22.128 ;
  LAYER M3 ;
        RECT 11.132 22.076 11.164 22.108 ;
  LAYER M1 ;
        RECT 11.196 19.62 11.228 22.128 ;
  LAYER M3 ;
        RECT 11.196 19.64 11.228 19.672 ;
  LAYER M1 ;
        RECT 11.26 19.62 11.292 22.128 ;
  LAYER M3 ;
        RECT 11.26 22.076 11.292 22.108 ;
  LAYER M1 ;
        RECT 11.324 19.62 11.356 22.128 ;
  LAYER M3 ;
        RECT 11.324 19.64 11.356 19.672 ;
  LAYER M1 ;
        RECT 11.388 19.62 11.42 22.128 ;
  LAYER M3 ;
        RECT 11.388 22.076 11.42 22.108 ;
  LAYER M1 ;
        RECT 11.452 19.62 11.484 22.128 ;
  LAYER M3 ;
        RECT 11.452 19.64 11.484 19.672 ;
  LAYER M1 ;
        RECT 11.516 19.62 11.548 22.128 ;
  LAYER M3 ;
        RECT 11.516 22.076 11.548 22.108 ;
  LAYER M1 ;
        RECT 11.58 19.62 11.612 22.128 ;
  LAYER M3 ;
        RECT 11.58 19.64 11.612 19.672 ;
  LAYER M1 ;
        RECT 11.644 19.62 11.676 22.128 ;
  LAYER M3 ;
        RECT 11.644 22.076 11.676 22.108 ;
  LAYER M1 ;
        RECT 11.708 19.62 11.74 22.128 ;
  LAYER M3 ;
        RECT 11.708 19.64 11.74 19.672 ;
  LAYER M1 ;
        RECT 11.772 19.62 11.804 22.128 ;
  LAYER M3 ;
        RECT 11.772 22.076 11.804 22.108 ;
  LAYER M1 ;
        RECT 11.836 19.62 11.868 22.128 ;
  LAYER M3 ;
        RECT 11.836 19.64 11.868 19.672 ;
  LAYER M1 ;
        RECT 11.9 19.62 11.932 22.128 ;
  LAYER M3 ;
        RECT 11.9 22.076 11.932 22.108 ;
  LAYER M1 ;
        RECT 11.964 19.62 11.996 22.128 ;
  LAYER M3 ;
        RECT 11.964 19.64 11.996 19.672 ;
  LAYER M1 ;
        RECT 12.028 19.62 12.06 22.128 ;
  LAYER M3 ;
        RECT 12.028 22.076 12.06 22.108 ;
  LAYER M1 ;
        RECT 12.092 19.62 12.124 22.128 ;
  LAYER M3 ;
        RECT 12.092 19.64 12.124 19.672 ;
  LAYER M1 ;
        RECT 12.156 19.62 12.188 22.128 ;
  LAYER M3 ;
        RECT 12.156 22.076 12.188 22.108 ;
  LAYER M1 ;
        RECT 12.22 19.62 12.252 22.128 ;
  LAYER M3 ;
        RECT 12.22 19.64 12.252 19.672 ;
  LAYER M1 ;
        RECT 12.284 19.62 12.316 22.128 ;
  LAYER M3 ;
        RECT 12.284 22.076 12.316 22.108 ;
  LAYER M1 ;
        RECT 12.348 19.62 12.38 22.128 ;
  LAYER M3 ;
        RECT 9.98 19.704 10.012 19.736 ;
  LAYER M2 ;
        RECT 12.348 19.768 12.38 19.8 ;
  LAYER M2 ;
        RECT 9.98 19.832 10.012 19.864 ;
  LAYER M2 ;
        RECT 12.348 19.896 12.38 19.928 ;
  LAYER M2 ;
        RECT 9.98 19.96 10.012 19.992 ;
  LAYER M2 ;
        RECT 12.348 20.024 12.38 20.056 ;
  LAYER M2 ;
        RECT 9.98 20.088 10.012 20.12 ;
  LAYER M2 ;
        RECT 12.348 20.152 12.38 20.184 ;
  LAYER M2 ;
        RECT 9.98 20.216 10.012 20.248 ;
  LAYER M2 ;
        RECT 12.348 20.28 12.38 20.312 ;
  LAYER M2 ;
        RECT 9.98 20.344 10.012 20.376 ;
  LAYER M2 ;
        RECT 12.348 20.408 12.38 20.44 ;
  LAYER M2 ;
        RECT 9.98 20.472 10.012 20.504 ;
  LAYER M2 ;
        RECT 12.348 20.536 12.38 20.568 ;
  LAYER M2 ;
        RECT 9.98 20.6 10.012 20.632 ;
  LAYER M2 ;
        RECT 12.348 20.664 12.38 20.696 ;
  LAYER M2 ;
        RECT 9.98 20.728 10.012 20.76 ;
  LAYER M2 ;
        RECT 12.348 20.792 12.38 20.824 ;
  LAYER M2 ;
        RECT 9.98 20.856 10.012 20.888 ;
  LAYER M2 ;
        RECT 12.348 20.92 12.38 20.952 ;
  LAYER M2 ;
        RECT 9.98 20.984 10.012 21.016 ;
  LAYER M2 ;
        RECT 12.348 21.048 12.38 21.08 ;
  LAYER M2 ;
        RECT 9.98 21.112 10.012 21.144 ;
  LAYER M2 ;
        RECT 12.348 21.176 12.38 21.208 ;
  LAYER M2 ;
        RECT 9.98 21.24 10.012 21.272 ;
  LAYER M2 ;
        RECT 12.348 21.304 12.38 21.336 ;
  LAYER M2 ;
        RECT 9.98 21.368 10.012 21.4 ;
  LAYER M2 ;
        RECT 12.348 21.432 12.38 21.464 ;
  LAYER M2 ;
        RECT 9.98 21.496 10.012 21.528 ;
  LAYER M2 ;
        RECT 12.348 21.56 12.38 21.592 ;
  LAYER M2 ;
        RECT 9.98 21.624 10.012 21.656 ;
  LAYER M2 ;
        RECT 12.348 21.688 12.38 21.72 ;
  LAYER M2 ;
        RECT 9.98 21.752 10.012 21.784 ;
  LAYER M2 ;
        RECT 12.348 21.816 12.38 21.848 ;
  LAYER M2 ;
        RECT 9.98 21.88 10.012 21.912 ;
  LAYER M2 ;
        RECT 12.348 21.944 12.38 21.976 ;
  LAYER M2 ;
        RECT 9.932 19.572 12.428 22.176 ;
  LAYER M1 ;
        RECT 13.276 0.972 13.308 3.48 ;
  LAYER M3 ;
        RECT 13.276 3.428 13.308 3.46 ;
  LAYER M1 ;
        RECT 13.34 0.972 13.372 3.48 ;
  LAYER M3 ;
        RECT 13.34 0.992 13.372 1.024 ;
  LAYER M1 ;
        RECT 13.404 0.972 13.436 3.48 ;
  LAYER M3 ;
        RECT 13.404 3.428 13.436 3.46 ;
  LAYER M1 ;
        RECT 13.468 0.972 13.5 3.48 ;
  LAYER M3 ;
        RECT 13.468 0.992 13.5 1.024 ;
  LAYER M1 ;
        RECT 13.532 0.972 13.564 3.48 ;
  LAYER M3 ;
        RECT 13.532 3.428 13.564 3.46 ;
  LAYER M1 ;
        RECT 13.596 0.972 13.628 3.48 ;
  LAYER M3 ;
        RECT 13.596 0.992 13.628 1.024 ;
  LAYER M1 ;
        RECT 13.66 0.972 13.692 3.48 ;
  LAYER M3 ;
        RECT 13.66 3.428 13.692 3.46 ;
  LAYER M1 ;
        RECT 13.724 0.972 13.756 3.48 ;
  LAYER M3 ;
        RECT 13.724 0.992 13.756 1.024 ;
  LAYER M1 ;
        RECT 13.788 0.972 13.82 3.48 ;
  LAYER M3 ;
        RECT 13.788 3.428 13.82 3.46 ;
  LAYER M1 ;
        RECT 13.852 0.972 13.884 3.48 ;
  LAYER M3 ;
        RECT 13.852 0.992 13.884 1.024 ;
  LAYER M1 ;
        RECT 13.916 0.972 13.948 3.48 ;
  LAYER M3 ;
        RECT 13.916 3.428 13.948 3.46 ;
  LAYER M1 ;
        RECT 13.98 0.972 14.012 3.48 ;
  LAYER M3 ;
        RECT 13.98 0.992 14.012 1.024 ;
  LAYER M1 ;
        RECT 14.044 0.972 14.076 3.48 ;
  LAYER M3 ;
        RECT 14.044 3.428 14.076 3.46 ;
  LAYER M1 ;
        RECT 14.108 0.972 14.14 3.48 ;
  LAYER M3 ;
        RECT 14.108 0.992 14.14 1.024 ;
  LAYER M1 ;
        RECT 14.172 0.972 14.204 3.48 ;
  LAYER M3 ;
        RECT 14.172 3.428 14.204 3.46 ;
  LAYER M1 ;
        RECT 14.236 0.972 14.268 3.48 ;
  LAYER M3 ;
        RECT 14.236 0.992 14.268 1.024 ;
  LAYER M1 ;
        RECT 14.3 0.972 14.332 3.48 ;
  LAYER M3 ;
        RECT 14.3 3.428 14.332 3.46 ;
  LAYER M1 ;
        RECT 14.364 0.972 14.396 3.48 ;
  LAYER M3 ;
        RECT 14.364 0.992 14.396 1.024 ;
  LAYER M1 ;
        RECT 14.428 0.972 14.46 3.48 ;
  LAYER M3 ;
        RECT 14.428 3.428 14.46 3.46 ;
  LAYER M1 ;
        RECT 14.492 0.972 14.524 3.48 ;
  LAYER M3 ;
        RECT 14.492 0.992 14.524 1.024 ;
  LAYER M1 ;
        RECT 14.556 0.972 14.588 3.48 ;
  LAYER M3 ;
        RECT 14.556 3.428 14.588 3.46 ;
  LAYER M1 ;
        RECT 14.62 0.972 14.652 3.48 ;
  LAYER M3 ;
        RECT 14.62 0.992 14.652 1.024 ;
  LAYER M1 ;
        RECT 14.684 0.972 14.716 3.48 ;
  LAYER M3 ;
        RECT 14.684 3.428 14.716 3.46 ;
  LAYER M1 ;
        RECT 14.748 0.972 14.78 3.48 ;
  LAYER M3 ;
        RECT 14.748 0.992 14.78 1.024 ;
  LAYER M1 ;
        RECT 14.812 0.972 14.844 3.48 ;
  LAYER M3 ;
        RECT 14.812 3.428 14.844 3.46 ;
  LAYER M1 ;
        RECT 14.876 0.972 14.908 3.48 ;
  LAYER M3 ;
        RECT 14.876 0.992 14.908 1.024 ;
  LAYER M1 ;
        RECT 14.94 0.972 14.972 3.48 ;
  LAYER M3 ;
        RECT 14.94 3.428 14.972 3.46 ;
  LAYER M1 ;
        RECT 15.004 0.972 15.036 3.48 ;
  LAYER M3 ;
        RECT 15.004 0.992 15.036 1.024 ;
  LAYER M1 ;
        RECT 15.068 0.972 15.1 3.48 ;
  LAYER M3 ;
        RECT 15.068 3.428 15.1 3.46 ;
  LAYER M1 ;
        RECT 15.132 0.972 15.164 3.48 ;
  LAYER M3 ;
        RECT 15.132 0.992 15.164 1.024 ;
  LAYER M1 ;
        RECT 15.196 0.972 15.228 3.48 ;
  LAYER M3 ;
        RECT 15.196 3.428 15.228 3.46 ;
  LAYER M1 ;
        RECT 15.26 0.972 15.292 3.48 ;
  LAYER M3 ;
        RECT 15.26 0.992 15.292 1.024 ;
  LAYER M1 ;
        RECT 15.324 0.972 15.356 3.48 ;
  LAYER M3 ;
        RECT 15.324 3.428 15.356 3.46 ;
  LAYER M1 ;
        RECT 15.388 0.972 15.42 3.48 ;
  LAYER M3 ;
        RECT 15.388 0.992 15.42 1.024 ;
  LAYER M1 ;
        RECT 15.452 0.972 15.484 3.48 ;
  LAYER M3 ;
        RECT 15.452 3.428 15.484 3.46 ;
  LAYER M1 ;
        RECT 15.516 0.972 15.548 3.48 ;
  LAYER M3 ;
        RECT 15.516 0.992 15.548 1.024 ;
  LAYER M1 ;
        RECT 15.58 0.972 15.612 3.48 ;
  LAYER M3 ;
        RECT 15.58 3.428 15.612 3.46 ;
  LAYER M1 ;
        RECT 15.644 0.972 15.676 3.48 ;
  LAYER M3 ;
        RECT 13.276 1.056 13.308 1.088 ;
  LAYER M2 ;
        RECT 15.644 1.12 15.676 1.152 ;
  LAYER M2 ;
        RECT 13.276 1.184 13.308 1.216 ;
  LAYER M2 ;
        RECT 15.644 1.248 15.676 1.28 ;
  LAYER M2 ;
        RECT 13.276 1.312 13.308 1.344 ;
  LAYER M2 ;
        RECT 15.644 1.376 15.676 1.408 ;
  LAYER M2 ;
        RECT 13.276 1.44 13.308 1.472 ;
  LAYER M2 ;
        RECT 15.644 1.504 15.676 1.536 ;
  LAYER M2 ;
        RECT 13.276 1.568 13.308 1.6 ;
  LAYER M2 ;
        RECT 15.644 1.632 15.676 1.664 ;
  LAYER M2 ;
        RECT 13.276 1.696 13.308 1.728 ;
  LAYER M2 ;
        RECT 15.644 1.76 15.676 1.792 ;
  LAYER M2 ;
        RECT 13.276 1.824 13.308 1.856 ;
  LAYER M2 ;
        RECT 15.644 1.888 15.676 1.92 ;
  LAYER M2 ;
        RECT 13.276 1.952 13.308 1.984 ;
  LAYER M2 ;
        RECT 15.644 2.016 15.676 2.048 ;
  LAYER M2 ;
        RECT 13.276 2.08 13.308 2.112 ;
  LAYER M2 ;
        RECT 15.644 2.144 15.676 2.176 ;
  LAYER M2 ;
        RECT 13.276 2.208 13.308 2.24 ;
  LAYER M2 ;
        RECT 15.644 2.272 15.676 2.304 ;
  LAYER M2 ;
        RECT 13.276 2.336 13.308 2.368 ;
  LAYER M2 ;
        RECT 15.644 2.4 15.676 2.432 ;
  LAYER M2 ;
        RECT 13.276 2.464 13.308 2.496 ;
  LAYER M2 ;
        RECT 15.644 2.528 15.676 2.56 ;
  LAYER M2 ;
        RECT 13.276 2.592 13.308 2.624 ;
  LAYER M2 ;
        RECT 15.644 2.656 15.676 2.688 ;
  LAYER M2 ;
        RECT 13.276 2.72 13.308 2.752 ;
  LAYER M2 ;
        RECT 15.644 2.784 15.676 2.816 ;
  LAYER M2 ;
        RECT 13.276 2.848 13.308 2.88 ;
  LAYER M2 ;
        RECT 15.644 2.912 15.676 2.944 ;
  LAYER M2 ;
        RECT 13.276 2.976 13.308 3.008 ;
  LAYER M2 ;
        RECT 15.644 3.04 15.676 3.072 ;
  LAYER M2 ;
        RECT 13.276 3.104 13.308 3.136 ;
  LAYER M2 ;
        RECT 15.644 3.168 15.676 3.2 ;
  LAYER M2 ;
        RECT 13.276 3.232 13.308 3.264 ;
  LAYER M2 ;
        RECT 15.644 3.296 15.676 3.328 ;
  LAYER M2 ;
        RECT 13.228 0.924 15.724 3.528 ;
  LAYER M1 ;
        RECT 13.276 4.08 13.308 6.588 ;
  LAYER M3 ;
        RECT 13.276 6.536 13.308 6.568 ;
  LAYER M1 ;
        RECT 13.34 4.08 13.372 6.588 ;
  LAYER M3 ;
        RECT 13.34 4.1 13.372 4.132 ;
  LAYER M1 ;
        RECT 13.404 4.08 13.436 6.588 ;
  LAYER M3 ;
        RECT 13.404 6.536 13.436 6.568 ;
  LAYER M1 ;
        RECT 13.468 4.08 13.5 6.588 ;
  LAYER M3 ;
        RECT 13.468 4.1 13.5 4.132 ;
  LAYER M1 ;
        RECT 13.532 4.08 13.564 6.588 ;
  LAYER M3 ;
        RECT 13.532 6.536 13.564 6.568 ;
  LAYER M1 ;
        RECT 13.596 4.08 13.628 6.588 ;
  LAYER M3 ;
        RECT 13.596 4.1 13.628 4.132 ;
  LAYER M1 ;
        RECT 13.66 4.08 13.692 6.588 ;
  LAYER M3 ;
        RECT 13.66 6.536 13.692 6.568 ;
  LAYER M1 ;
        RECT 13.724 4.08 13.756 6.588 ;
  LAYER M3 ;
        RECT 13.724 4.1 13.756 4.132 ;
  LAYER M1 ;
        RECT 13.788 4.08 13.82 6.588 ;
  LAYER M3 ;
        RECT 13.788 6.536 13.82 6.568 ;
  LAYER M1 ;
        RECT 13.852 4.08 13.884 6.588 ;
  LAYER M3 ;
        RECT 13.852 4.1 13.884 4.132 ;
  LAYER M1 ;
        RECT 13.916 4.08 13.948 6.588 ;
  LAYER M3 ;
        RECT 13.916 6.536 13.948 6.568 ;
  LAYER M1 ;
        RECT 13.98 4.08 14.012 6.588 ;
  LAYER M3 ;
        RECT 13.98 4.1 14.012 4.132 ;
  LAYER M1 ;
        RECT 14.044 4.08 14.076 6.588 ;
  LAYER M3 ;
        RECT 14.044 6.536 14.076 6.568 ;
  LAYER M1 ;
        RECT 14.108 4.08 14.14 6.588 ;
  LAYER M3 ;
        RECT 14.108 4.1 14.14 4.132 ;
  LAYER M1 ;
        RECT 14.172 4.08 14.204 6.588 ;
  LAYER M3 ;
        RECT 14.172 6.536 14.204 6.568 ;
  LAYER M1 ;
        RECT 14.236 4.08 14.268 6.588 ;
  LAYER M3 ;
        RECT 14.236 4.1 14.268 4.132 ;
  LAYER M1 ;
        RECT 14.3 4.08 14.332 6.588 ;
  LAYER M3 ;
        RECT 14.3 6.536 14.332 6.568 ;
  LAYER M1 ;
        RECT 14.364 4.08 14.396 6.588 ;
  LAYER M3 ;
        RECT 14.364 4.1 14.396 4.132 ;
  LAYER M1 ;
        RECT 14.428 4.08 14.46 6.588 ;
  LAYER M3 ;
        RECT 14.428 6.536 14.46 6.568 ;
  LAYER M1 ;
        RECT 14.492 4.08 14.524 6.588 ;
  LAYER M3 ;
        RECT 14.492 4.1 14.524 4.132 ;
  LAYER M1 ;
        RECT 14.556 4.08 14.588 6.588 ;
  LAYER M3 ;
        RECT 14.556 6.536 14.588 6.568 ;
  LAYER M1 ;
        RECT 14.62 4.08 14.652 6.588 ;
  LAYER M3 ;
        RECT 14.62 4.1 14.652 4.132 ;
  LAYER M1 ;
        RECT 14.684 4.08 14.716 6.588 ;
  LAYER M3 ;
        RECT 14.684 6.536 14.716 6.568 ;
  LAYER M1 ;
        RECT 14.748 4.08 14.78 6.588 ;
  LAYER M3 ;
        RECT 14.748 4.1 14.78 4.132 ;
  LAYER M1 ;
        RECT 14.812 4.08 14.844 6.588 ;
  LAYER M3 ;
        RECT 14.812 6.536 14.844 6.568 ;
  LAYER M1 ;
        RECT 14.876 4.08 14.908 6.588 ;
  LAYER M3 ;
        RECT 14.876 4.1 14.908 4.132 ;
  LAYER M1 ;
        RECT 14.94 4.08 14.972 6.588 ;
  LAYER M3 ;
        RECT 14.94 6.536 14.972 6.568 ;
  LAYER M1 ;
        RECT 15.004 4.08 15.036 6.588 ;
  LAYER M3 ;
        RECT 15.004 4.1 15.036 4.132 ;
  LAYER M1 ;
        RECT 15.068 4.08 15.1 6.588 ;
  LAYER M3 ;
        RECT 15.068 6.536 15.1 6.568 ;
  LAYER M1 ;
        RECT 15.132 4.08 15.164 6.588 ;
  LAYER M3 ;
        RECT 15.132 4.1 15.164 4.132 ;
  LAYER M1 ;
        RECT 15.196 4.08 15.228 6.588 ;
  LAYER M3 ;
        RECT 15.196 6.536 15.228 6.568 ;
  LAYER M1 ;
        RECT 15.26 4.08 15.292 6.588 ;
  LAYER M3 ;
        RECT 15.26 4.1 15.292 4.132 ;
  LAYER M1 ;
        RECT 15.324 4.08 15.356 6.588 ;
  LAYER M3 ;
        RECT 15.324 6.536 15.356 6.568 ;
  LAYER M1 ;
        RECT 15.388 4.08 15.42 6.588 ;
  LAYER M3 ;
        RECT 15.388 4.1 15.42 4.132 ;
  LAYER M1 ;
        RECT 15.452 4.08 15.484 6.588 ;
  LAYER M3 ;
        RECT 15.452 6.536 15.484 6.568 ;
  LAYER M1 ;
        RECT 15.516 4.08 15.548 6.588 ;
  LAYER M3 ;
        RECT 15.516 4.1 15.548 4.132 ;
  LAYER M1 ;
        RECT 15.58 4.08 15.612 6.588 ;
  LAYER M3 ;
        RECT 15.58 6.536 15.612 6.568 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 6.588 ;
  LAYER M3 ;
        RECT 13.276 4.164 13.308 4.196 ;
  LAYER M2 ;
        RECT 15.644 4.228 15.676 4.26 ;
  LAYER M2 ;
        RECT 13.276 4.292 13.308 4.324 ;
  LAYER M2 ;
        RECT 15.644 4.356 15.676 4.388 ;
  LAYER M2 ;
        RECT 13.276 4.42 13.308 4.452 ;
  LAYER M2 ;
        RECT 15.644 4.484 15.676 4.516 ;
  LAYER M2 ;
        RECT 13.276 4.548 13.308 4.58 ;
  LAYER M2 ;
        RECT 15.644 4.612 15.676 4.644 ;
  LAYER M2 ;
        RECT 13.276 4.676 13.308 4.708 ;
  LAYER M2 ;
        RECT 15.644 4.74 15.676 4.772 ;
  LAYER M2 ;
        RECT 13.276 4.804 13.308 4.836 ;
  LAYER M2 ;
        RECT 15.644 4.868 15.676 4.9 ;
  LAYER M2 ;
        RECT 13.276 4.932 13.308 4.964 ;
  LAYER M2 ;
        RECT 15.644 4.996 15.676 5.028 ;
  LAYER M2 ;
        RECT 13.276 5.06 13.308 5.092 ;
  LAYER M2 ;
        RECT 15.644 5.124 15.676 5.156 ;
  LAYER M2 ;
        RECT 13.276 5.188 13.308 5.22 ;
  LAYER M2 ;
        RECT 15.644 5.252 15.676 5.284 ;
  LAYER M2 ;
        RECT 13.276 5.316 13.308 5.348 ;
  LAYER M2 ;
        RECT 15.644 5.38 15.676 5.412 ;
  LAYER M2 ;
        RECT 13.276 5.444 13.308 5.476 ;
  LAYER M2 ;
        RECT 15.644 5.508 15.676 5.54 ;
  LAYER M2 ;
        RECT 13.276 5.572 13.308 5.604 ;
  LAYER M2 ;
        RECT 15.644 5.636 15.676 5.668 ;
  LAYER M2 ;
        RECT 13.276 5.7 13.308 5.732 ;
  LAYER M2 ;
        RECT 15.644 5.764 15.676 5.796 ;
  LAYER M2 ;
        RECT 13.276 5.828 13.308 5.86 ;
  LAYER M2 ;
        RECT 15.644 5.892 15.676 5.924 ;
  LAYER M2 ;
        RECT 13.276 5.956 13.308 5.988 ;
  LAYER M2 ;
        RECT 15.644 6.02 15.676 6.052 ;
  LAYER M2 ;
        RECT 13.276 6.084 13.308 6.116 ;
  LAYER M2 ;
        RECT 15.644 6.148 15.676 6.18 ;
  LAYER M2 ;
        RECT 13.276 6.212 13.308 6.244 ;
  LAYER M2 ;
        RECT 15.644 6.276 15.676 6.308 ;
  LAYER M2 ;
        RECT 13.276 6.34 13.308 6.372 ;
  LAYER M2 ;
        RECT 15.644 6.404 15.676 6.436 ;
  LAYER M2 ;
        RECT 13.228 4.032 15.724 6.636 ;
  LAYER M1 ;
        RECT 13.276 7.188 13.308 9.696 ;
  LAYER M3 ;
        RECT 13.276 9.644 13.308 9.676 ;
  LAYER M1 ;
        RECT 13.34 7.188 13.372 9.696 ;
  LAYER M3 ;
        RECT 13.34 7.208 13.372 7.24 ;
  LAYER M1 ;
        RECT 13.404 7.188 13.436 9.696 ;
  LAYER M3 ;
        RECT 13.404 9.644 13.436 9.676 ;
  LAYER M1 ;
        RECT 13.468 7.188 13.5 9.696 ;
  LAYER M3 ;
        RECT 13.468 7.208 13.5 7.24 ;
  LAYER M1 ;
        RECT 13.532 7.188 13.564 9.696 ;
  LAYER M3 ;
        RECT 13.532 9.644 13.564 9.676 ;
  LAYER M1 ;
        RECT 13.596 7.188 13.628 9.696 ;
  LAYER M3 ;
        RECT 13.596 7.208 13.628 7.24 ;
  LAYER M1 ;
        RECT 13.66 7.188 13.692 9.696 ;
  LAYER M3 ;
        RECT 13.66 9.644 13.692 9.676 ;
  LAYER M1 ;
        RECT 13.724 7.188 13.756 9.696 ;
  LAYER M3 ;
        RECT 13.724 7.208 13.756 7.24 ;
  LAYER M1 ;
        RECT 13.788 7.188 13.82 9.696 ;
  LAYER M3 ;
        RECT 13.788 9.644 13.82 9.676 ;
  LAYER M1 ;
        RECT 13.852 7.188 13.884 9.696 ;
  LAYER M3 ;
        RECT 13.852 7.208 13.884 7.24 ;
  LAYER M1 ;
        RECT 13.916 7.188 13.948 9.696 ;
  LAYER M3 ;
        RECT 13.916 9.644 13.948 9.676 ;
  LAYER M1 ;
        RECT 13.98 7.188 14.012 9.696 ;
  LAYER M3 ;
        RECT 13.98 7.208 14.012 7.24 ;
  LAYER M1 ;
        RECT 14.044 7.188 14.076 9.696 ;
  LAYER M3 ;
        RECT 14.044 9.644 14.076 9.676 ;
  LAYER M1 ;
        RECT 14.108 7.188 14.14 9.696 ;
  LAYER M3 ;
        RECT 14.108 7.208 14.14 7.24 ;
  LAYER M1 ;
        RECT 14.172 7.188 14.204 9.696 ;
  LAYER M3 ;
        RECT 14.172 9.644 14.204 9.676 ;
  LAYER M1 ;
        RECT 14.236 7.188 14.268 9.696 ;
  LAYER M3 ;
        RECT 14.236 7.208 14.268 7.24 ;
  LAYER M1 ;
        RECT 14.3 7.188 14.332 9.696 ;
  LAYER M3 ;
        RECT 14.3 9.644 14.332 9.676 ;
  LAYER M1 ;
        RECT 14.364 7.188 14.396 9.696 ;
  LAYER M3 ;
        RECT 14.364 7.208 14.396 7.24 ;
  LAYER M1 ;
        RECT 14.428 7.188 14.46 9.696 ;
  LAYER M3 ;
        RECT 14.428 9.644 14.46 9.676 ;
  LAYER M1 ;
        RECT 14.492 7.188 14.524 9.696 ;
  LAYER M3 ;
        RECT 14.492 7.208 14.524 7.24 ;
  LAYER M1 ;
        RECT 14.556 7.188 14.588 9.696 ;
  LAYER M3 ;
        RECT 14.556 9.644 14.588 9.676 ;
  LAYER M1 ;
        RECT 14.62 7.188 14.652 9.696 ;
  LAYER M3 ;
        RECT 14.62 7.208 14.652 7.24 ;
  LAYER M1 ;
        RECT 14.684 7.188 14.716 9.696 ;
  LAYER M3 ;
        RECT 14.684 9.644 14.716 9.676 ;
  LAYER M1 ;
        RECT 14.748 7.188 14.78 9.696 ;
  LAYER M3 ;
        RECT 14.748 7.208 14.78 7.24 ;
  LAYER M1 ;
        RECT 14.812 7.188 14.844 9.696 ;
  LAYER M3 ;
        RECT 14.812 9.644 14.844 9.676 ;
  LAYER M1 ;
        RECT 14.876 7.188 14.908 9.696 ;
  LAYER M3 ;
        RECT 14.876 7.208 14.908 7.24 ;
  LAYER M1 ;
        RECT 14.94 7.188 14.972 9.696 ;
  LAYER M3 ;
        RECT 14.94 9.644 14.972 9.676 ;
  LAYER M1 ;
        RECT 15.004 7.188 15.036 9.696 ;
  LAYER M3 ;
        RECT 15.004 7.208 15.036 7.24 ;
  LAYER M1 ;
        RECT 15.068 7.188 15.1 9.696 ;
  LAYER M3 ;
        RECT 15.068 9.644 15.1 9.676 ;
  LAYER M1 ;
        RECT 15.132 7.188 15.164 9.696 ;
  LAYER M3 ;
        RECT 15.132 7.208 15.164 7.24 ;
  LAYER M1 ;
        RECT 15.196 7.188 15.228 9.696 ;
  LAYER M3 ;
        RECT 15.196 9.644 15.228 9.676 ;
  LAYER M1 ;
        RECT 15.26 7.188 15.292 9.696 ;
  LAYER M3 ;
        RECT 15.26 7.208 15.292 7.24 ;
  LAYER M1 ;
        RECT 15.324 7.188 15.356 9.696 ;
  LAYER M3 ;
        RECT 15.324 9.644 15.356 9.676 ;
  LAYER M1 ;
        RECT 15.388 7.188 15.42 9.696 ;
  LAYER M3 ;
        RECT 15.388 7.208 15.42 7.24 ;
  LAYER M1 ;
        RECT 15.452 7.188 15.484 9.696 ;
  LAYER M3 ;
        RECT 15.452 9.644 15.484 9.676 ;
  LAYER M1 ;
        RECT 15.516 7.188 15.548 9.696 ;
  LAYER M3 ;
        RECT 15.516 7.208 15.548 7.24 ;
  LAYER M1 ;
        RECT 15.58 7.188 15.612 9.696 ;
  LAYER M3 ;
        RECT 15.58 9.644 15.612 9.676 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 9.696 ;
  LAYER M3 ;
        RECT 13.276 7.272 13.308 7.304 ;
  LAYER M2 ;
        RECT 15.644 7.336 15.676 7.368 ;
  LAYER M2 ;
        RECT 13.276 7.4 13.308 7.432 ;
  LAYER M2 ;
        RECT 15.644 7.464 15.676 7.496 ;
  LAYER M2 ;
        RECT 13.276 7.528 13.308 7.56 ;
  LAYER M2 ;
        RECT 15.644 7.592 15.676 7.624 ;
  LAYER M2 ;
        RECT 13.276 7.656 13.308 7.688 ;
  LAYER M2 ;
        RECT 15.644 7.72 15.676 7.752 ;
  LAYER M2 ;
        RECT 13.276 7.784 13.308 7.816 ;
  LAYER M2 ;
        RECT 15.644 7.848 15.676 7.88 ;
  LAYER M2 ;
        RECT 13.276 7.912 13.308 7.944 ;
  LAYER M2 ;
        RECT 15.644 7.976 15.676 8.008 ;
  LAYER M2 ;
        RECT 13.276 8.04 13.308 8.072 ;
  LAYER M2 ;
        RECT 15.644 8.104 15.676 8.136 ;
  LAYER M2 ;
        RECT 13.276 8.168 13.308 8.2 ;
  LAYER M2 ;
        RECT 15.644 8.232 15.676 8.264 ;
  LAYER M2 ;
        RECT 13.276 8.296 13.308 8.328 ;
  LAYER M2 ;
        RECT 15.644 8.36 15.676 8.392 ;
  LAYER M2 ;
        RECT 13.276 8.424 13.308 8.456 ;
  LAYER M2 ;
        RECT 15.644 8.488 15.676 8.52 ;
  LAYER M2 ;
        RECT 13.276 8.552 13.308 8.584 ;
  LAYER M2 ;
        RECT 15.644 8.616 15.676 8.648 ;
  LAYER M2 ;
        RECT 13.276 8.68 13.308 8.712 ;
  LAYER M2 ;
        RECT 15.644 8.744 15.676 8.776 ;
  LAYER M2 ;
        RECT 13.276 8.808 13.308 8.84 ;
  LAYER M2 ;
        RECT 15.644 8.872 15.676 8.904 ;
  LAYER M2 ;
        RECT 13.276 8.936 13.308 8.968 ;
  LAYER M2 ;
        RECT 15.644 9 15.676 9.032 ;
  LAYER M2 ;
        RECT 13.276 9.064 13.308 9.096 ;
  LAYER M2 ;
        RECT 15.644 9.128 15.676 9.16 ;
  LAYER M2 ;
        RECT 13.276 9.192 13.308 9.224 ;
  LAYER M2 ;
        RECT 15.644 9.256 15.676 9.288 ;
  LAYER M2 ;
        RECT 13.276 9.32 13.308 9.352 ;
  LAYER M2 ;
        RECT 15.644 9.384 15.676 9.416 ;
  LAYER M2 ;
        RECT 13.276 9.448 13.308 9.48 ;
  LAYER M2 ;
        RECT 15.644 9.512 15.676 9.544 ;
  LAYER M2 ;
        RECT 13.228 7.14 15.724 9.744 ;
  LAYER M1 ;
        RECT 13.276 10.296 13.308 12.804 ;
  LAYER M3 ;
        RECT 13.276 12.752 13.308 12.784 ;
  LAYER M1 ;
        RECT 13.34 10.296 13.372 12.804 ;
  LAYER M3 ;
        RECT 13.34 10.316 13.372 10.348 ;
  LAYER M1 ;
        RECT 13.404 10.296 13.436 12.804 ;
  LAYER M3 ;
        RECT 13.404 12.752 13.436 12.784 ;
  LAYER M1 ;
        RECT 13.468 10.296 13.5 12.804 ;
  LAYER M3 ;
        RECT 13.468 10.316 13.5 10.348 ;
  LAYER M1 ;
        RECT 13.532 10.296 13.564 12.804 ;
  LAYER M3 ;
        RECT 13.532 12.752 13.564 12.784 ;
  LAYER M1 ;
        RECT 13.596 10.296 13.628 12.804 ;
  LAYER M3 ;
        RECT 13.596 10.316 13.628 10.348 ;
  LAYER M1 ;
        RECT 13.66 10.296 13.692 12.804 ;
  LAYER M3 ;
        RECT 13.66 12.752 13.692 12.784 ;
  LAYER M1 ;
        RECT 13.724 10.296 13.756 12.804 ;
  LAYER M3 ;
        RECT 13.724 10.316 13.756 10.348 ;
  LAYER M1 ;
        RECT 13.788 10.296 13.82 12.804 ;
  LAYER M3 ;
        RECT 13.788 12.752 13.82 12.784 ;
  LAYER M1 ;
        RECT 13.852 10.296 13.884 12.804 ;
  LAYER M3 ;
        RECT 13.852 10.316 13.884 10.348 ;
  LAYER M1 ;
        RECT 13.916 10.296 13.948 12.804 ;
  LAYER M3 ;
        RECT 13.916 12.752 13.948 12.784 ;
  LAYER M1 ;
        RECT 13.98 10.296 14.012 12.804 ;
  LAYER M3 ;
        RECT 13.98 10.316 14.012 10.348 ;
  LAYER M1 ;
        RECT 14.044 10.296 14.076 12.804 ;
  LAYER M3 ;
        RECT 14.044 12.752 14.076 12.784 ;
  LAYER M1 ;
        RECT 14.108 10.296 14.14 12.804 ;
  LAYER M3 ;
        RECT 14.108 10.316 14.14 10.348 ;
  LAYER M1 ;
        RECT 14.172 10.296 14.204 12.804 ;
  LAYER M3 ;
        RECT 14.172 12.752 14.204 12.784 ;
  LAYER M1 ;
        RECT 14.236 10.296 14.268 12.804 ;
  LAYER M3 ;
        RECT 14.236 10.316 14.268 10.348 ;
  LAYER M1 ;
        RECT 14.3 10.296 14.332 12.804 ;
  LAYER M3 ;
        RECT 14.3 12.752 14.332 12.784 ;
  LAYER M1 ;
        RECT 14.364 10.296 14.396 12.804 ;
  LAYER M3 ;
        RECT 14.364 10.316 14.396 10.348 ;
  LAYER M1 ;
        RECT 14.428 10.296 14.46 12.804 ;
  LAYER M3 ;
        RECT 14.428 12.752 14.46 12.784 ;
  LAYER M1 ;
        RECT 14.492 10.296 14.524 12.804 ;
  LAYER M3 ;
        RECT 14.492 10.316 14.524 10.348 ;
  LAYER M1 ;
        RECT 14.556 10.296 14.588 12.804 ;
  LAYER M3 ;
        RECT 14.556 12.752 14.588 12.784 ;
  LAYER M1 ;
        RECT 14.62 10.296 14.652 12.804 ;
  LAYER M3 ;
        RECT 14.62 10.316 14.652 10.348 ;
  LAYER M1 ;
        RECT 14.684 10.296 14.716 12.804 ;
  LAYER M3 ;
        RECT 14.684 12.752 14.716 12.784 ;
  LAYER M1 ;
        RECT 14.748 10.296 14.78 12.804 ;
  LAYER M3 ;
        RECT 14.748 10.316 14.78 10.348 ;
  LAYER M1 ;
        RECT 14.812 10.296 14.844 12.804 ;
  LAYER M3 ;
        RECT 14.812 12.752 14.844 12.784 ;
  LAYER M1 ;
        RECT 14.876 10.296 14.908 12.804 ;
  LAYER M3 ;
        RECT 14.876 10.316 14.908 10.348 ;
  LAYER M1 ;
        RECT 14.94 10.296 14.972 12.804 ;
  LAYER M3 ;
        RECT 14.94 12.752 14.972 12.784 ;
  LAYER M1 ;
        RECT 15.004 10.296 15.036 12.804 ;
  LAYER M3 ;
        RECT 15.004 10.316 15.036 10.348 ;
  LAYER M1 ;
        RECT 15.068 10.296 15.1 12.804 ;
  LAYER M3 ;
        RECT 15.068 12.752 15.1 12.784 ;
  LAYER M1 ;
        RECT 15.132 10.296 15.164 12.804 ;
  LAYER M3 ;
        RECT 15.132 10.316 15.164 10.348 ;
  LAYER M1 ;
        RECT 15.196 10.296 15.228 12.804 ;
  LAYER M3 ;
        RECT 15.196 12.752 15.228 12.784 ;
  LAYER M1 ;
        RECT 15.26 10.296 15.292 12.804 ;
  LAYER M3 ;
        RECT 15.26 10.316 15.292 10.348 ;
  LAYER M1 ;
        RECT 15.324 10.296 15.356 12.804 ;
  LAYER M3 ;
        RECT 15.324 12.752 15.356 12.784 ;
  LAYER M1 ;
        RECT 15.388 10.296 15.42 12.804 ;
  LAYER M3 ;
        RECT 15.388 10.316 15.42 10.348 ;
  LAYER M1 ;
        RECT 15.452 10.296 15.484 12.804 ;
  LAYER M3 ;
        RECT 15.452 12.752 15.484 12.784 ;
  LAYER M1 ;
        RECT 15.516 10.296 15.548 12.804 ;
  LAYER M3 ;
        RECT 15.516 10.316 15.548 10.348 ;
  LAYER M1 ;
        RECT 15.58 10.296 15.612 12.804 ;
  LAYER M3 ;
        RECT 15.58 12.752 15.612 12.784 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 12.804 ;
  LAYER M3 ;
        RECT 13.276 10.38 13.308 10.412 ;
  LAYER M2 ;
        RECT 15.644 10.444 15.676 10.476 ;
  LAYER M2 ;
        RECT 13.276 10.508 13.308 10.54 ;
  LAYER M2 ;
        RECT 15.644 10.572 15.676 10.604 ;
  LAYER M2 ;
        RECT 13.276 10.636 13.308 10.668 ;
  LAYER M2 ;
        RECT 15.644 10.7 15.676 10.732 ;
  LAYER M2 ;
        RECT 13.276 10.764 13.308 10.796 ;
  LAYER M2 ;
        RECT 15.644 10.828 15.676 10.86 ;
  LAYER M2 ;
        RECT 13.276 10.892 13.308 10.924 ;
  LAYER M2 ;
        RECT 15.644 10.956 15.676 10.988 ;
  LAYER M2 ;
        RECT 13.276 11.02 13.308 11.052 ;
  LAYER M2 ;
        RECT 15.644 11.084 15.676 11.116 ;
  LAYER M2 ;
        RECT 13.276 11.148 13.308 11.18 ;
  LAYER M2 ;
        RECT 15.644 11.212 15.676 11.244 ;
  LAYER M2 ;
        RECT 13.276 11.276 13.308 11.308 ;
  LAYER M2 ;
        RECT 15.644 11.34 15.676 11.372 ;
  LAYER M2 ;
        RECT 13.276 11.404 13.308 11.436 ;
  LAYER M2 ;
        RECT 15.644 11.468 15.676 11.5 ;
  LAYER M2 ;
        RECT 13.276 11.532 13.308 11.564 ;
  LAYER M2 ;
        RECT 15.644 11.596 15.676 11.628 ;
  LAYER M2 ;
        RECT 13.276 11.66 13.308 11.692 ;
  LAYER M2 ;
        RECT 15.644 11.724 15.676 11.756 ;
  LAYER M2 ;
        RECT 13.276 11.788 13.308 11.82 ;
  LAYER M2 ;
        RECT 15.644 11.852 15.676 11.884 ;
  LAYER M2 ;
        RECT 13.276 11.916 13.308 11.948 ;
  LAYER M2 ;
        RECT 15.644 11.98 15.676 12.012 ;
  LAYER M2 ;
        RECT 13.276 12.044 13.308 12.076 ;
  LAYER M2 ;
        RECT 15.644 12.108 15.676 12.14 ;
  LAYER M2 ;
        RECT 13.276 12.172 13.308 12.204 ;
  LAYER M2 ;
        RECT 15.644 12.236 15.676 12.268 ;
  LAYER M2 ;
        RECT 13.276 12.3 13.308 12.332 ;
  LAYER M2 ;
        RECT 15.644 12.364 15.676 12.396 ;
  LAYER M2 ;
        RECT 13.276 12.428 13.308 12.46 ;
  LAYER M2 ;
        RECT 15.644 12.492 15.676 12.524 ;
  LAYER M2 ;
        RECT 13.276 12.556 13.308 12.588 ;
  LAYER M2 ;
        RECT 15.644 12.62 15.676 12.652 ;
  LAYER M2 ;
        RECT 13.228 10.248 15.724 12.852 ;
  LAYER M1 ;
        RECT 13.276 13.404 13.308 15.912 ;
  LAYER M3 ;
        RECT 13.276 15.86 13.308 15.892 ;
  LAYER M1 ;
        RECT 13.34 13.404 13.372 15.912 ;
  LAYER M3 ;
        RECT 13.34 13.424 13.372 13.456 ;
  LAYER M1 ;
        RECT 13.404 13.404 13.436 15.912 ;
  LAYER M3 ;
        RECT 13.404 15.86 13.436 15.892 ;
  LAYER M1 ;
        RECT 13.468 13.404 13.5 15.912 ;
  LAYER M3 ;
        RECT 13.468 13.424 13.5 13.456 ;
  LAYER M1 ;
        RECT 13.532 13.404 13.564 15.912 ;
  LAYER M3 ;
        RECT 13.532 15.86 13.564 15.892 ;
  LAYER M1 ;
        RECT 13.596 13.404 13.628 15.912 ;
  LAYER M3 ;
        RECT 13.596 13.424 13.628 13.456 ;
  LAYER M1 ;
        RECT 13.66 13.404 13.692 15.912 ;
  LAYER M3 ;
        RECT 13.66 15.86 13.692 15.892 ;
  LAYER M1 ;
        RECT 13.724 13.404 13.756 15.912 ;
  LAYER M3 ;
        RECT 13.724 13.424 13.756 13.456 ;
  LAYER M1 ;
        RECT 13.788 13.404 13.82 15.912 ;
  LAYER M3 ;
        RECT 13.788 15.86 13.82 15.892 ;
  LAYER M1 ;
        RECT 13.852 13.404 13.884 15.912 ;
  LAYER M3 ;
        RECT 13.852 13.424 13.884 13.456 ;
  LAYER M1 ;
        RECT 13.916 13.404 13.948 15.912 ;
  LAYER M3 ;
        RECT 13.916 15.86 13.948 15.892 ;
  LAYER M1 ;
        RECT 13.98 13.404 14.012 15.912 ;
  LAYER M3 ;
        RECT 13.98 13.424 14.012 13.456 ;
  LAYER M1 ;
        RECT 14.044 13.404 14.076 15.912 ;
  LAYER M3 ;
        RECT 14.044 15.86 14.076 15.892 ;
  LAYER M1 ;
        RECT 14.108 13.404 14.14 15.912 ;
  LAYER M3 ;
        RECT 14.108 13.424 14.14 13.456 ;
  LAYER M1 ;
        RECT 14.172 13.404 14.204 15.912 ;
  LAYER M3 ;
        RECT 14.172 15.86 14.204 15.892 ;
  LAYER M1 ;
        RECT 14.236 13.404 14.268 15.912 ;
  LAYER M3 ;
        RECT 14.236 13.424 14.268 13.456 ;
  LAYER M1 ;
        RECT 14.3 13.404 14.332 15.912 ;
  LAYER M3 ;
        RECT 14.3 15.86 14.332 15.892 ;
  LAYER M1 ;
        RECT 14.364 13.404 14.396 15.912 ;
  LAYER M3 ;
        RECT 14.364 13.424 14.396 13.456 ;
  LAYER M1 ;
        RECT 14.428 13.404 14.46 15.912 ;
  LAYER M3 ;
        RECT 14.428 15.86 14.46 15.892 ;
  LAYER M1 ;
        RECT 14.492 13.404 14.524 15.912 ;
  LAYER M3 ;
        RECT 14.492 13.424 14.524 13.456 ;
  LAYER M1 ;
        RECT 14.556 13.404 14.588 15.912 ;
  LAYER M3 ;
        RECT 14.556 15.86 14.588 15.892 ;
  LAYER M1 ;
        RECT 14.62 13.404 14.652 15.912 ;
  LAYER M3 ;
        RECT 14.62 13.424 14.652 13.456 ;
  LAYER M1 ;
        RECT 14.684 13.404 14.716 15.912 ;
  LAYER M3 ;
        RECT 14.684 15.86 14.716 15.892 ;
  LAYER M1 ;
        RECT 14.748 13.404 14.78 15.912 ;
  LAYER M3 ;
        RECT 14.748 13.424 14.78 13.456 ;
  LAYER M1 ;
        RECT 14.812 13.404 14.844 15.912 ;
  LAYER M3 ;
        RECT 14.812 15.86 14.844 15.892 ;
  LAYER M1 ;
        RECT 14.876 13.404 14.908 15.912 ;
  LAYER M3 ;
        RECT 14.876 13.424 14.908 13.456 ;
  LAYER M1 ;
        RECT 14.94 13.404 14.972 15.912 ;
  LAYER M3 ;
        RECT 14.94 15.86 14.972 15.892 ;
  LAYER M1 ;
        RECT 15.004 13.404 15.036 15.912 ;
  LAYER M3 ;
        RECT 15.004 13.424 15.036 13.456 ;
  LAYER M1 ;
        RECT 15.068 13.404 15.1 15.912 ;
  LAYER M3 ;
        RECT 15.068 15.86 15.1 15.892 ;
  LAYER M1 ;
        RECT 15.132 13.404 15.164 15.912 ;
  LAYER M3 ;
        RECT 15.132 13.424 15.164 13.456 ;
  LAYER M1 ;
        RECT 15.196 13.404 15.228 15.912 ;
  LAYER M3 ;
        RECT 15.196 15.86 15.228 15.892 ;
  LAYER M1 ;
        RECT 15.26 13.404 15.292 15.912 ;
  LAYER M3 ;
        RECT 15.26 13.424 15.292 13.456 ;
  LAYER M1 ;
        RECT 15.324 13.404 15.356 15.912 ;
  LAYER M3 ;
        RECT 15.324 15.86 15.356 15.892 ;
  LAYER M1 ;
        RECT 15.388 13.404 15.42 15.912 ;
  LAYER M3 ;
        RECT 15.388 13.424 15.42 13.456 ;
  LAYER M1 ;
        RECT 15.452 13.404 15.484 15.912 ;
  LAYER M3 ;
        RECT 15.452 15.86 15.484 15.892 ;
  LAYER M1 ;
        RECT 15.516 13.404 15.548 15.912 ;
  LAYER M3 ;
        RECT 15.516 13.424 15.548 13.456 ;
  LAYER M1 ;
        RECT 15.58 13.404 15.612 15.912 ;
  LAYER M3 ;
        RECT 15.58 15.86 15.612 15.892 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 15.912 ;
  LAYER M3 ;
        RECT 13.276 13.488 13.308 13.52 ;
  LAYER M2 ;
        RECT 15.644 13.552 15.676 13.584 ;
  LAYER M2 ;
        RECT 13.276 13.616 13.308 13.648 ;
  LAYER M2 ;
        RECT 15.644 13.68 15.676 13.712 ;
  LAYER M2 ;
        RECT 13.276 13.744 13.308 13.776 ;
  LAYER M2 ;
        RECT 15.644 13.808 15.676 13.84 ;
  LAYER M2 ;
        RECT 13.276 13.872 13.308 13.904 ;
  LAYER M2 ;
        RECT 15.644 13.936 15.676 13.968 ;
  LAYER M2 ;
        RECT 13.276 14 13.308 14.032 ;
  LAYER M2 ;
        RECT 15.644 14.064 15.676 14.096 ;
  LAYER M2 ;
        RECT 13.276 14.128 13.308 14.16 ;
  LAYER M2 ;
        RECT 15.644 14.192 15.676 14.224 ;
  LAYER M2 ;
        RECT 13.276 14.256 13.308 14.288 ;
  LAYER M2 ;
        RECT 15.644 14.32 15.676 14.352 ;
  LAYER M2 ;
        RECT 13.276 14.384 13.308 14.416 ;
  LAYER M2 ;
        RECT 15.644 14.448 15.676 14.48 ;
  LAYER M2 ;
        RECT 13.276 14.512 13.308 14.544 ;
  LAYER M2 ;
        RECT 15.644 14.576 15.676 14.608 ;
  LAYER M2 ;
        RECT 13.276 14.64 13.308 14.672 ;
  LAYER M2 ;
        RECT 15.644 14.704 15.676 14.736 ;
  LAYER M2 ;
        RECT 13.276 14.768 13.308 14.8 ;
  LAYER M2 ;
        RECT 15.644 14.832 15.676 14.864 ;
  LAYER M2 ;
        RECT 13.276 14.896 13.308 14.928 ;
  LAYER M2 ;
        RECT 15.644 14.96 15.676 14.992 ;
  LAYER M2 ;
        RECT 13.276 15.024 13.308 15.056 ;
  LAYER M2 ;
        RECT 15.644 15.088 15.676 15.12 ;
  LAYER M2 ;
        RECT 13.276 15.152 13.308 15.184 ;
  LAYER M2 ;
        RECT 15.644 15.216 15.676 15.248 ;
  LAYER M2 ;
        RECT 13.276 15.28 13.308 15.312 ;
  LAYER M2 ;
        RECT 15.644 15.344 15.676 15.376 ;
  LAYER M2 ;
        RECT 13.276 15.408 13.308 15.44 ;
  LAYER M2 ;
        RECT 15.644 15.472 15.676 15.504 ;
  LAYER M2 ;
        RECT 13.276 15.536 13.308 15.568 ;
  LAYER M2 ;
        RECT 15.644 15.6 15.676 15.632 ;
  LAYER M2 ;
        RECT 13.276 15.664 13.308 15.696 ;
  LAYER M2 ;
        RECT 15.644 15.728 15.676 15.76 ;
  LAYER M2 ;
        RECT 13.228 13.356 15.724 15.96 ;
  LAYER M1 ;
        RECT 13.276 16.512 13.308 19.02 ;
  LAYER M3 ;
        RECT 13.276 18.968 13.308 19 ;
  LAYER M1 ;
        RECT 13.34 16.512 13.372 19.02 ;
  LAYER M3 ;
        RECT 13.34 16.532 13.372 16.564 ;
  LAYER M1 ;
        RECT 13.404 16.512 13.436 19.02 ;
  LAYER M3 ;
        RECT 13.404 18.968 13.436 19 ;
  LAYER M1 ;
        RECT 13.468 16.512 13.5 19.02 ;
  LAYER M3 ;
        RECT 13.468 16.532 13.5 16.564 ;
  LAYER M1 ;
        RECT 13.532 16.512 13.564 19.02 ;
  LAYER M3 ;
        RECT 13.532 18.968 13.564 19 ;
  LAYER M1 ;
        RECT 13.596 16.512 13.628 19.02 ;
  LAYER M3 ;
        RECT 13.596 16.532 13.628 16.564 ;
  LAYER M1 ;
        RECT 13.66 16.512 13.692 19.02 ;
  LAYER M3 ;
        RECT 13.66 18.968 13.692 19 ;
  LAYER M1 ;
        RECT 13.724 16.512 13.756 19.02 ;
  LAYER M3 ;
        RECT 13.724 16.532 13.756 16.564 ;
  LAYER M1 ;
        RECT 13.788 16.512 13.82 19.02 ;
  LAYER M3 ;
        RECT 13.788 18.968 13.82 19 ;
  LAYER M1 ;
        RECT 13.852 16.512 13.884 19.02 ;
  LAYER M3 ;
        RECT 13.852 16.532 13.884 16.564 ;
  LAYER M1 ;
        RECT 13.916 16.512 13.948 19.02 ;
  LAYER M3 ;
        RECT 13.916 18.968 13.948 19 ;
  LAYER M1 ;
        RECT 13.98 16.512 14.012 19.02 ;
  LAYER M3 ;
        RECT 13.98 16.532 14.012 16.564 ;
  LAYER M1 ;
        RECT 14.044 16.512 14.076 19.02 ;
  LAYER M3 ;
        RECT 14.044 18.968 14.076 19 ;
  LAYER M1 ;
        RECT 14.108 16.512 14.14 19.02 ;
  LAYER M3 ;
        RECT 14.108 16.532 14.14 16.564 ;
  LAYER M1 ;
        RECT 14.172 16.512 14.204 19.02 ;
  LAYER M3 ;
        RECT 14.172 18.968 14.204 19 ;
  LAYER M1 ;
        RECT 14.236 16.512 14.268 19.02 ;
  LAYER M3 ;
        RECT 14.236 16.532 14.268 16.564 ;
  LAYER M1 ;
        RECT 14.3 16.512 14.332 19.02 ;
  LAYER M3 ;
        RECT 14.3 18.968 14.332 19 ;
  LAYER M1 ;
        RECT 14.364 16.512 14.396 19.02 ;
  LAYER M3 ;
        RECT 14.364 16.532 14.396 16.564 ;
  LAYER M1 ;
        RECT 14.428 16.512 14.46 19.02 ;
  LAYER M3 ;
        RECT 14.428 18.968 14.46 19 ;
  LAYER M1 ;
        RECT 14.492 16.512 14.524 19.02 ;
  LAYER M3 ;
        RECT 14.492 16.532 14.524 16.564 ;
  LAYER M1 ;
        RECT 14.556 16.512 14.588 19.02 ;
  LAYER M3 ;
        RECT 14.556 18.968 14.588 19 ;
  LAYER M1 ;
        RECT 14.62 16.512 14.652 19.02 ;
  LAYER M3 ;
        RECT 14.62 16.532 14.652 16.564 ;
  LAYER M1 ;
        RECT 14.684 16.512 14.716 19.02 ;
  LAYER M3 ;
        RECT 14.684 18.968 14.716 19 ;
  LAYER M1 ;
        RECT 14.748 16.512 14.78 19.02 ;
  LAYER M3 ;
        RECT 14.748 16.532 14.78 16.564 ;
  LAYER M1 ;
        RECT 14.812 16.512 14.844 19.02 ;
  LAYER M3 ;
        RECT 14.812 18.968 14.844 19 ;
  LAYER M1 ;
        RECT 14.876 16.512 14.908 19.02 ;
  LAYER M3 ;
        RECT 14.876 16.532 14.908 16.564 ;
  LAYER M1 ;
        RECT 14.94 16.512 14.972 19.02 ;
  LAYER M3 ;
        RECT 14.94 18.968 14.972 19 ;
  LAYER M1 ;
        RECT 15.004 16.512 15.036 19.02 ;
  LAYER M3 ;
        RECT 15.004 16.532 15.036 16.564 ;
  LAYER M1 ;
        RECT 15.068 16.512 15.1 19.02 ;
  LAYER M3 ;
        RECT 15.068 18.968 15.1 19 ;
  LAYER M1 ;
        RECT 15.132 16.512 15.164 19.02 ;
  LAYER M3 ;
        RECT 15.132 16.532 15.164 16.564 ;
  LAYER M1 ;
        RECT 15.196 16.512 15.228 19.02 ;
  LAYER M3 ;
        RECT 15.196 18.968 15.228 19 ;
  LAYER M1 ;
        RECT 15.26 16.512 15.292 19.02 ;
  LAYER M3 ;
        RECT 15.26 16.532 15.292 16.564 ;
  LAYER M1 ;
        RECT 15.324 16.512 15.356 19.02 ;
  LAYER M3 ;
        RECT 15.324 18.968 15.356 19 ;
  LAYER M1 ;
        RECT 15.388 16.512 15.42 19.02 ;
  LAYER M3 ;
        RECT 15.388 16.532 15.42 16.564 ;
  LAYER M1 ;
        RECT 15.452 16.512 15.484 19.02 ;
  LAYER M3 ;
        RECT 15.452 18.968 15.484 19 ;
  LAYER M1 ;
        RECT 15.516 16.512 15.548 19.02 ;
  LAYER M3 ;
        RECT 15.516 16.532 15.548 16.564 ;
  LAYER M1 ;
        RECT 15.58 16.512 15.612 19.02 ;
  LAYER M3 ;
        RECT 15.58 18.968 15.612 19 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 19.02 ;
  LAYER M3 ;
        RECT 13.276 16.596 13.308 16.628 ;
  LAYER M2 ;
        RECT 15.644 16.66 15.676 16.692 ;
  LAYER M2 ;
        RECT 13.276 16.724 13.308 16.756 ;
  LAYER M2 ;
        RECT 15.644 16.788 15.676 16.82 ;
  LAYER M2 ;
        RECT 13.276 16.852 13.308 16.884 ;
  LAYER M2 ;
        RECT 15.644 16.916 15.676 16.948 ;
  LAYER M2 ;
        RECT 13.276 16.98 13.308 17.012 ;
  LAYER M2 ;
        RECT 15.644 17.044 15.676 17.076 ;
  LAYER M2 ;
        RECT 13.276 17.108 13.308 17.14 ;
  LAYER M2 ;
        RECT 15.644 17.172 15.676 17.204 ;
  LAYER M2 ;
        RECT 13.276 17.236 13.308 17.268 ;
  LAYER M2 ;
        RECT 15.644 17.3 15.676 17.332 ;
  LAYER M2 ;
        RECT 13.276 17.364 13.308 17.396 ;
  LAYER M2 ;
        RECT 15.644 17.428 15.676 17.46 ;
  LAYER M2 ;
        RECT 13.276 17.492 13.308 17.524 ;
  LAYER M2 ;
        RECT 15.644 17.556 15.676 17.588 ;
  LAYER M2 ;
        RECT 13.276 17.62 13.308 17.652 ;
  LAYER M2 ;
        RECT 15.644 17.684 15.676 17.716 ;
  LAYER M2 ;
        RECT 13.276 17.748 13.308 17.78 ;
  LAYER M2 ;
        RECT 15.644 17.812 15.676 17.844 ;
  LAYER M2 ;
        RECT 13.276 17.876 13.308 17.908 ;
  LAYER M2 ;
        RECT 15.644 17.94 15.676 17.972 ;
  LAYER M2 ;
        RECT 13.276 18.004 13.308 18.036 ;
  LAYER M2 ;
        RECT 15.644 18.068 15.676 18.1 ;
  LAYER M2 ;
        RECT 13.276 18.132 13.308 18.164 ;
  LAYER M2 ;
        RECT 15.644 18.196 15.676 18.228 ;
  LAYER M2 ;
        RECT 13.276 18.26 13.308 18.292 ;
  LAYER M2 ;
        RECT 15.644 18.324 15.676 18.356 ;
  LAYER M2 ;
        RECT 13.276 18.388 13.308 18.42 ;
  LAYER M2 ;
        RECT 15.644 18.452 15.676 18.484 ;
  LAYER M2 ;
        RECT 13.276 18.516 13.308 18.548 ;
  LAYER M2 ;
        RECT 15.644 18.58 15.676 18.612 ;
  LAYER M2 ;
        RECT 13.276 18.644 13.308 18.676 ;
  LAYER M2 ;
        RECT 15.644 18.708 15.676 18.74 ;
  LAYER M2 ;
        RECT 13.276 18.772 13.308 18.804 ;
  LAYER M2 ;
        RECT 15.644 18.836 15.676 18.868 ;
  LAYER M2 ;
        RECT 13.228 16.464 15.724 19.068 ;
  LAYER M1 ;
        RECT 13.276 19.62 13.308 22.128 ;
  LAYER M3 ;
        RECT 13.276 22.076 13.308 22.108 ;
  LAYER M1 ;
        RECT 13.34 19.62 13.372 22.128 ;
  LAYER M3 ;
        RECT 13.34 19.64 13.372 19.672 ;
  LAYER M1 ;
        RECT 13.404 19.62 13.436 22.128 ;
  LAYER M3 ;
        RECT 13.404 22.076 13.436 22.108 ;
  LAYER M1 ;
        RECT 13.468 19.62 13.5 22.128 ;
  LAYER M3 ;
        RECT 13.468 19.64 13.5 19.672 ;
  LAYER M1 ;
        RECT 13.532 19.62 13.564 22.128 ;
  LAYER M3 ;
        RECT 13.532 22.076 13.564 22.108 ;
  LAYER M1 ;
        RECT 13.596 19.62 13.628 22.128 ;
  LAYER M3 ;
        RECT 13.596 19.64 13.628 19.672 ;
  LAYER M1 ;
        RECT 13.66 19.62 13.692 22.128 ;
  LAYER M3 ;
        RECT 13.66 22.076 13.692 22.108 ;
  LAYER M1 ;
        RECT 13.724 19.62 13.756 22.128 ;
  LAYER M3 ;
        RECT 13.724 19.64 13.756 19.672 ;
  LAYER M1 ;
        RECT 13.788 19.62 13.82 22.128 ;
  LAYER M3 ;
        RECT 13.788 22.076 13.82 22.108 ;
  LAYER M1 ;
        RECT 13.852 19.62 13.884 22.128 ;
  LAYER M3 ;
        RECT 13.852 19.64 13.884 19.672 ;
  LAYER M1 ;
        RECT 13.916 19.62 13.948 22.128 ;
  LAYER M3 ;
        RECT 13.916 22.076 13.948 22.108 ;
  LAYER M1 ;
        RECT 13.98 19.62 14.012 22.128 ;
  LAYER M3 ;
        RECT 13.98 19.64 14.012 19.672 ;
  LAYER M1 ;
        RECT 14.044 19.62 14.076 22.128 ;
  LAYER M3 ;
        RECT 14.044 22.076 14.076 22.108 ;
  LAYER M1 ;
        RECT 14.108 19.62 14.14 22.128 ;
  LAYER M3 ;
        RECT 14.108 19.64 14.14 19.672 ;
  LAYER M1 ;
        RECT 14.172 19.62 14.204 22.128 ;
  LAYER M3 ;
        RECT 14.172 22.076 14.204 22.108 ;
  LAYER M1 ;
        RECT 14.236 19.62 14.268 22.128 ;
  LAYER M3 ;
        RECT 14.236 19.64 14.268 19.672 ;
  LAYER M1 ;
        RECT 14.3 19.62 14.332 22.128 ;
  LAYER M3 ;
        RECT 14.3 22.076 14.332 22.108 ;
  LAYER M1 ;
        RECT 14.364 19.62 14.396 22.128 ;
  LAYER M3 ;
        RECT 14.364 19.64 14.396 19.672 ;
  LAYER M1 ;
        RECT 14.428 19.62 14.46 22.128 ;
  LAYER M3 ;
        RECT 14.428 22.076 14.46 22.108 ;
  LAYER M1 ;
        RECT 14.492 19.62 14.524 22.128 ;
  LAYER M3 ;
        RECT 14.492 19.64 14.524 19.672 ;
  LAYER M1 ;
        RECT 14.556 19.62 14.588 22.128 ;
  LAYER M3 ;
        RECT 14.556 22.076 14.588 22.108 ;
  LAYER M1 ;
        RECT 14.62 19.62 14.652 22.128 ;
  LAYER M3 ;
        RECT 14.62 19.64 14.652 19.672 ;
  LAYER M1 ;
        RECT 14.684 19.62 14.716 22.128 ;
  LAYER M3 ;
        RECT 14.684 22.076 14.716 22.108 ;
  LAYER M1 ;
        RECT 14.748 19.62 14.78 22.128 ;
  LAYER M3 ;
        RECT 14.748 19.64 14.78 19.672 ;
  LAYER M1 ;
        RECT 14.812 19.62 14.844 22.128 ;
  LAYER M3 ;
        RECT 14.812 22.076 14.844 22.108 ;
  LAYER M1 ;
        RECT 14.876 19.62 14.908 22.128 ;
  LAYER M3 ;
        RECT 14.876 19.64 14.908 19.672 ;
  LAYER M1 ;
        RECT 14.94 19.62 14.972 22.128 ;
  LAYER M3 ;
        RECT 14.94 22.076 14.972 22.108 ;
  LAYER M1 ;
        RECT 15.004 19.62 15.036 22.128 ;
  LAYER M3 ;
        RECT 15.004 19.64 15.036 19.672 ;
  LAYER M1 ;
        RECT 15.068 19.62 15.1 22.128 ;
  LAYER M3 ;
        RECT 15.068 22.076 15.1 22.108 ;
  LAYER M1 ;
        RECT 15.132 19.62 15.164 22.128 ;
  LAYER M3 ;
        RECT 15.132 19.64 15.164 19.672 ;
  LAYER M1 ;
        RECT 15.196 19.62 15.228 22.128 ;
  LAYER M3 ;
        RECT 15.196 22.076 15.228 22.108 ;
  LAYER M1 ;
        RECT 15.26 19.62 15.292 22.128 ;
  LAYER M3 ;
        RECT 15.26 19.64 15.292 19.672 ;
  LAYER M1 ;
        RECT 15.324 19.62 15.356 22.128 ;
  LAYER M3 ;
        RECT 15.324 22.076 15.356 22.108 ;
  LAYER M1 ;
        RECT 15.388 19.62 15.42 22.128 ;
  LAYER M3 ;
        RECT 15.388 19.64 15.42 19.672 ;
  LAYER M1 ;
        RECT 15.452 19.62 15.484 22.128 ;
  LAYER M3 ;
        RECT 15.452 22.076 15.484 22.108 ;
  LAYER M1 ;
        RECT 15.516 19.62 15.548 22.128 ;
  LAYER M3 ;
        RECT 15.516 19.64 15.548 19.672 ;
  LAYER M1 ;
        RECT 15.58 19.62 15.612 22.128 ;
  LAYER M3 ;
        RECT 15.58 22.076 15.612 22.108 ;
  LAYER M1 ;
        RECT 15.644 19.62 15.676 22.128 ;
  LAYER M3 ;
        RECT 13.276 19.704 13.308 19.736 ;
  LAYER M2 ;
        RECT 15.644 19.768 15.676 19.8 ;
  LAYER M2 ;
        RECT 13.276 19.832 13.308 19.864 ;
  LAYER M2 ;
        RECT 15.644 19.896 15.676 19.928 ;
  LAYER M2 ;
        RECT 13.276 19.96 13.308 19.992 ;
  LAYER M2 ;
        RECT 15.644 20.024 15.676 20.056 ;
  LAYER M2 ;
        RECT 13.276 20.088 13.308 20.12 ;
  LAYER M2 ;
        RECT 15.644 20.152 15.676 20.184 ;
  LAYER M2 ;
        RECT 13.276 20.216 13.308 20.248 ;
  LAYER M2 ;
        RECT 15.644 20.28 15.676 20.312 ;
  LAYER M2 ;
        RECT 13.276 20.344 13.308 20.376 ;
  LAYER M2 ;
        RECT 15.644 20.408 15.676 20.44 ;
  LAYER M2 ;
        RECT 13.276 20.472 13.308 20.504 ;
  LAYER M2 ;
        RECT 15.644 20.536 15.676 20.568 ;
  LAYER M2 ;
        RECT 13.276 20.6 13.308 20.632 ;
  LAYER M2 ;
        RECT 15.644 20.664 15.676 20.696 ;
  LAYER M2 ;
        RECT 13.276 20.728 13.308 20.76 ;
  LAYER M2 ;
        RECT 15.644 20.792 15.676 20.824 ;
  LAYER M2 ;
        RECT 13.276 20.856 13.308 20.888 ;
  LAYER M2 ;
        RECT 15.644 20.92 15.676 20.952 ;
  LAYER M2 ;
        RECT 13.276 20.984 13.308 21.016 ;
  LAYER M2 ;
        RECT 15.644 21.048 15.676 21.08 ;
  LAYER M2 ;
        RECT 13.276 21.112 13.308 21.144 ;
  LAYER M2 ;
        RECT 15.644 21.176 15.676 21.208 ;
  LAYER M2 ;
        RECT 13.276 21.24 13.308 21.272 ;
  LAYER M2 ;
        RECT 15.644 21.304 15.676 21.336 ;
  LAYER M2 ;
        RECT 13.276 21.368 13.308 21.4 ;
  LAYER M2 ;
        RECT 15.644 21.432 15.676 21.464 ;
  LAYER M2 ;
        RECT 13.276 21.496 13.308 21.528 ;
  LAYER M2 ;
        RECT 15.644 21.56 15.676 21.592 ;
  LAYER M2 ;
        RECT 13.276 21.624 13.308 21.656 ;
  LAYER M2 ;
        RECT 15.644 21.688 15.676 21.72 ;
  LAYER M2 ;
        RECT 13.276 21.752 13.308 21.784 ;
  LAYER M2 ;
        RECT 15.644 21.816 15.676 21.848 ;
  LAYER M2 ;
        RECT 13.276 21.88 13.308 21.912 ;
  LAYER M2 ;
        RECT 15.644 21.944 15.676 21.976 ;
  LAYER M2 ;
        RECT 13.228 19.572 15.724 22.176 ;
  END 
END Cap_60fF_Cap_60fF
