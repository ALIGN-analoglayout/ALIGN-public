MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 16.64 BY 18.984 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.624 18.528 6.656 18.6 ;
      LAYER M2 ;
        RECT 6.604 18.548 6.676 18.58 ;
      LAYER M1 ;
        RECT 10.144 18.528 10.176 18.6 ;
      LAYER M2 ;
        RECT 10.124 18.548 10.196 18.58 ;
      LAYER M2 ;
        RECT 6.64 18.548 10.16 18.58 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.144 0.384 6.176 0.456 ;
      LAYER M2 ;
        RECT 6.124 0.404 6.196 0.436 ;
      LAYER M1 ;
        RECT 9.664 0.384 9.696 0.456 ;
      LAYER M2 ;
        RECT 9.644 0.404 9.716 0.436 ;
      LAYER M2 ;
        RECT 6.16 0.404 9.68 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.784 18.696 6.816 18.768 ;
      LAYER M2 ;
        RECT 6.764 18.716 6.836 18.748 ;
      LAYER M1 ;
        RECT 10.304 18.696 10.336 18.768 ;
      LAYER M2 ;
        RECT 10.284 18.716 10.356 18.748 ;
      LAYER M2 ;
        RECT 6.8 18.716 10.32 18.748 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.304 0.216 6.336 0.288 ;
      LAYER M2 ;
        RECT 6.284 0.236 6.356 0.268 ;
      LAYER M1 ;
        RECT 9.824 0.216 9.856 0.288 ;
      LAYER M2 ;
        RECT 9.804 0.236 9.876 0.268 ;
      LAYER M2 ;
        RECT 6.32 0.236 9.84 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 9.504 6.768 9.536 6.84 ;
  LAYER M2 ;
        RECT 9.484 6.788 9.556 6.82 ;
  LAYER M2 ;
        RECT 6.16 6.788 9.52 6.82 ;
  LAYER M1 ;
        RECT 6.144 6.768 6.176 6.84 ;
  LAYER M2 ;
        RECT 6.124 6.788 6.196 6.82 ;
  LAYER M1 ;
        RECT 5.984 12.648 6.016 12.72 ;
  LAYER M2 ;
        RECT 5.964 12.668 6.036 12.7 ;
  LAYER M1 ;
        RECT 5.984 12.516 6.016 12.684 ;
  LAYER M1 ;
        RECT 5.984 12.48 6.016 12.552 ;
  LAYER M2 ;
        RECT 5.964 12.5 6.036 12.532 ;
  LAYER M2 ;
        RECT 6 12.5 6.16 12.532 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 12.552 ;
  LAYER M2 ;
        RECT 6.124 12.5 6.196 12.532 ;
  LAYER M1 ;
        RECT 6.144 0.384 6.176 0.456 ;
  LAYER M2 ;
        RECT 6.124 0.404 6.196 0.436 ;
  LAYER M1 ;
        RECT 6.144 0.42 6.176 0.588 ;
  LAYER M1 ;
        RECT 6.144 0.588 6.176 12.516 ;
  LAYER M1 ;
        RECT 13.024 3.828 13.056 3.9 ;
  LAYER M2 ;
        RECT 13.004 3.848 13.076 3.88 ;
  LAYER M2 ;
        RECT 9.68 3.848 13.04 3.88 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 3.9 ;
  LAYER M2 ;
        RECT 9.644 3.848 9.716 3.88 ;
  LAYER M1 ;
        RECT 9.664 0.384 9.696 0.456 ;
  LAYER M2 ;
        RECT 9.644 0.404 9.716 0.436 ;
  LAYER M1 ;
        RECT 9.664 0.42 9.696 0.588 ;
  LAYER M1 ;
        RECT 9.664 0.588 9.696 3.864 ;
  LAYER M2 ;
        RECT 6.16 0.404 9.68 0.436 ;
  LAYER M1 ;
        RECT 5.984 6.768 6.016 6.84 ;
  LAYER M2 ;
        RECT 5.964 6.788 6.036 6.82 ;
  LAYER M1 ;
        RECT 5.984 6.636 6.016 6.804 ;
  LAYER M1 ;
        RECT 5.984 6.6 6.016 6.672 ;
  LAYER M2 ;
        RECT 5.964 6.62 6.036 6.652 ;
  LAYER M2 ;
        RECT 6 6.62 6.32 6.652 ;
  LAYER M1 ;
        RECT 6.304 6.6 6.336 6.672 ;
  LAYER M2 ;
        RECT 6.284 6.62 6.356 6.652 ;
  LAYER M1 ;
        RECT 5.984 9.708 6.016 9.78 ;
  LAYER M2 ;
        RECT 5.964 9.728 6.036 9.76 ;
  LAYER M1 ;
        RECT 5.984 9.576 6.016 9.744 ;
  LAYER M1 ;
        RECT 5.984 9.54 6.016 9.612 ;
  LAYER M2 ;
        RECT 5.964 9.56 6.036 9.592 ;
  LAYER M2 ;
        RECT 6 9.56 6.32 9.592 ;
  LAYER M1 ;
        RECT 6.304 9.54 6.336 9.612 ;
  LAYER M2 ;
        RECT 6.284 9.56 6.356 9.592 ;
  LAYER M1 ;
        RECT 9.504 3.828 9.536 3.9 ;
  LAYER M2 ;
        RECT 9.484 3.848 9.556 3.88 ;
  LAYER M2 ;
        RECT 6.32 3.848 9.52 3.88 ;
  LAYER M1 ;
        RECT 6.304 3.828 6.336 3.9 ;
  LAYER M2 ;
        RECT 6.284 3.848 6.356 3.88 ;
  LAYER M1 ;
        RECT 9.504 12.648 9.536 12.72 ;
  LAYER M2 ;
        RECT 9.484 12.668 9.556 12.7 ;
  LAYER M2 ;
        RECT 6.32 12.668 9.52 12.7 ;
  LAYER M1 ;
        RECT 6.304 12.648 6.336 12.72 ;
  LAYER M2 ;
        RECT 6.284 12.668 6.356 12.7 ;
  LAYER M1 ;
        RECT 6.304 0.216 6.336 0.288 ;
  LAYER M2 ;
        RECT 6.284 0.236 6.356 0.268 ;
  LAYER M1 ;
        RECT 6.304 0.252 6.336 0.588 ;
  LAYER M1 ;
        RECT 6.304 0.588 6.336 12.684 ;
  LAYER M1 ;
        RECT 13.024 9.708 13.056 9.78 ;
  LAYER M2 ;
        RECT 13.004 9.728 13.076 9.76 ;
  LAYER M2 ;
        RECT 9.84 9.728 13.04 9.76 ;
  LAYER M1 ;
        RECT 9.824 9.708 9.856 9.78 ;
  LAYER M2 ;
        RECT 9.804 9.728 9.876 9.76 ;
  LAYER M1 ;
        RECT 13.024 6.768 13.056 6.84 ;
  LAYER M2 ;
        RECT 13.004 6.788 13.076 6.82 ;
  LAYER M2 ;
        RECT 9.84 6.788 13.04 6.82 ;
  LAYER M1 ;
        RECT 9.824 6.768 9.856 6.84 ;
  LAYER M2 ;
        RECT 9.804 6.788 9.876 6.82 ;
  LAYER M1 ;
        RECT 9.824 0.216 9.856 0.288 ;
  LAYER M2 ;
        RECT 9.804 0.236 9.876 0.268 ;
  LAYER M1 ;
        RECT 9.824 0.252 9.856 0.588 ;
  LAYER M1 ;
        RECT 9.824 0.588 9.856 9.744 ;
  LAYER M2 ;
        RECT 6.32 0.236 9.84 0.268 ;
  LAYER M1 ;
        RECT 5.984 0.888 6.016 0.96 ;
  LAYER M2 ;
        RECT 5.964 0.908 6.036 0.94 ;
  LAYER M1 ;
        RECT 5.984 0.756 6.016 0.924 ;
  LAYER M1 ;
        RECT 5.984 0.72 6.016 0.792 ;
  LAYER M2 ;
        RECT 5.964 0.74 6.036 0.772 ;
  LAYER M2 ;
        RECT 6 0.74 6.48 0.772 ;
  LAYER M1 ;
        RECT 6.464 0.72 6.496 0.792 ;
  LAYER M2 ;
        RECT 6.444 0.74 6.516 0.772 ;
  LAYER M1 ;
        RECT 5.984 3.828 6.016 3.9 ;
  LAYER M2 ;
        RECT 5.964 3.848 6.036 3.88 ;
  LAYER M1 ;
        RECT 5.984 3.696 6.016 3.864 ;
  LAYER M1 ;
        RECT 5.984 3.66 6.016 3.732 ;
  LAYER M2 ;
        RECT 5.964 3.68 6.036 3.712 ;
  LAYER M2 ;
        RECT 6 3.68 6.48 3.712 ;
  LAYER M1 ;
        RECT 6.464 3.66 6.496 3.732 ;
  LAYER M2 ;
        RECT 6.444 3.68 6.516 3.712 ;
  LAYER M1 ;
        RECT 5.984 15.588 6.016 15.66 ;
  LAYER M2 ;
        RECT 5.964 15.608 6.036 15.64 ;
  LAYER M1 ;
        RECT 5.984 15.456 6.016 15.624 ;
  LAYER M1 ;
        RECT 5.984 15.42 6.016 15.492 ;
  LAYER M2 ;
        RECT 5.964 15.44 6.036 15.472 ;
  LAYER M2 ;
        RECT 6 15.44 6.48 15.472 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 15.492 ;
  LAYER M2 ;
        RECT 6.444 15.44 6.516 15.472 ;
  LAYER M1 ;
        RECT 9.504 0.888 9.536 0.96 ;
  LAYER M2 ;
        RECT 9.484 0.908 9.556 0.94 ;
  LAYER M2 ;
        RECT 6.48 0.908 9.52 0.94 ;
  LAYER M1 ;
        RECT 6.464 0.888 6.496 0.96 ;
  LAYER M2 ;
        RECT 6.444 0.908 6.516 0.94 ;
  LAYER M1 ;
        RECT 9.504 9.708 9.536 9.78 ;
  LAYER M2 ;
        RECT 9.484 9.728 9.556 9.76 ;
  LAYER M2 ;
        RECT 6.48 9.728 9.52 9.76 ;
  LAYER M1 ;
        RECT 6.464 9.708 6.496 9.78 ;
  LAYER M2 ;
        RECT 6.444 9.728 6.516 9.76 ;
  LAYER M1 ;
        RECT 9.504 15.588 9.536 15.66 ;
  LAYER M2 ;
        RECT 9.484 15.608 9.556 15.64 ;
  LAYER M2 ;
        RECT 6.48 15.608 9.52 15.64 ;
  LAYER M1 ;
        RECT 6.464 15.588 6.496 15.66 ;
  LAYER M2 ;
        RECT 6.444 15.608 6.516 15.64 ;
  LAYER M1 ;
        RECT 6.464 0.048 6.496 0.12 ;
  LAYER M2 ;
        RECT 6.444 0.068 6.516 0.1 ;
  LAYER M1 ;
        RECT 6.464 0.084 6.496 0.588 ;
  LAYER M1 ;
        RECT 6.464 0.588 6.496 15.624 ;
  LAYER M1 ;
        RECT 13.024 0.888 13.056 0.96 ;
  LAYER M2 ;
        RECT 13.004 0.908 13.076 0.94 ;
  LAYER M2 ;
        RECT 10 0.908 13.04 0.94 ;
  LAYER M1 ;
        RECT 9.984 0.888 10.016 0.96 ;
  LAYER M2 ;
        RECT 9.964 0.908 10.036 0.94 ;
  LAYER M1 ;
        RECT 13.024 12.648 13.056 12.72 ;
  LAYER M2 ;
        RECT 13.004 12.668 13.076 12.7 ;
  LAYER M2 ;
        RECT 10 12.668 13.04 12.7 ;
  LAYER M1 ;
        RECT 9.984 12.648 10.016 12.72 ;
  LAYER M2 ;
        RECT 9.964 12.668 10.036 12.7 ;
  LAYER M1 ;
        RECT 13.024 15.588 13.056 15.66 ;
  LAYER M2 ;
        RECT 13.004 15.608 13.076 15.64 ;
  LAYER M2 ;
        RECT 10 15.608 13.04 15.64 ;
  LAYER M1 ;
        RECT 9.984 15.588 10.016 15.66 ;
  LAYER M2 ;
        RECT 9.964 15.608 10.036 15.64 ;
  LAYER M1 ;
        RECT 9.984 0.048 10.016 0.12 ;
  LAYER M2 ;
        RECT 9.964 0.068 10.036 0.1 ;
  LAYER M1 ;
        RECT 9.984 0.084 10.016 0.588 ;
  LAYER M1 ;
        RECT 9.984 0.588 10.016 15.624 ;
  LAYER M2 ;
        RECT 6.48 0.068 10 0.1 ;
  LAYER M1 ;
        RECT 2.464 15.588 2.496 15.66 ;
  LAYER M2 ;
        RECT 2.444 15.608 2.516 15.64 ;
  LAYER M2 ;
        RECT 2.48 15.608 6 15.64 ;
  LAYER M1 ;
        RECT 5.984 15.588 6.016 15.66 ;
  LAYER M2 ;
        RECT 5.964 15.608 6.036 15.64 ;
  LAYER M1 ;
        RECT 2.464 12.648 2.496 12.72 ;
  LAYER M2 ;
        RECT 2.444 12.668 2.516 12.7 ;
  LAYER M1 ;
        RECT 2.464 12.684 2.496 15.624 ;
  LAYER M1 ;
        RECT 2.464 15.588 2.496 15.66 ;
  LAYER M2 ;
        RECT 2.444 15.608 2.516 15.64 ;
  LAYER M1 ;
        RECT 2.464 9.708 2.496 9.78 ;
  LAYER M2 ;
        RECT 2.444 9.728 2.516 9.76 ;
  LAYER M1 ;
        RECT 2.464 9.744 2.496 12.684 ;
  LAYER M1 ;
        RECT 2.464 12.648 2.496 12.72 ;
  LAYER M2 ;
        RECT 2.444 12.668 2.516 12.7 ;
  LAYER M1 ;
        RECT 2.464 6.768 2.496 6.84 ;
  LAYER M2 ;
        RECT 2.444 6.788 2.516 6.82 ;
  LAYER M1 ;
        RECT 2.464 6.804 2.496 9.744 ;
  LAYER M1 ;
        RECT 2.464 9.708 2.496 9.78 ;
  LAYER M2 ;
        RECT 2.444 9.728 2.516 9.76 ;
  LAYER M1 ;
        RECT 2.464 3.828 2.496 3.9 ;
  LAYER M2 ;
        RECT 2.444 3.848 2.516 3.88 ;
  LAYER M1 ;
        RECT 2.464 3.864 2.496 6.804 ;
  LAYER M1 ;
        RECT 2.464 6.768 2.496 6.84 ;
  LAYER M2 ;
        RECT 2.444 6.788 2.516 6.82 ;
  LAYER M1 ;
        RECT 2.464 0.888 2.496 0.96 ;
  LAYER M2 ;
        RECT 2.444 0.908 2.516 0.94 ;
  LAYER M1 ;
        RECT 2.464 0.924 2.496 3.864 ;
  LAYER M1 ;
        RECT 2.464 3.828 2.496 3.9 ;
  LAYER M2 ;
        RECT 2.444 3.848 2.516 3.88 ;
  LAYER M1 ;
        RECT 16.544 15.588 16.576 15.66 ;
  LAYER M2 ;
        RECT 16.524 15.608 16.596 15.64 ;
  LAYER M2 ;
        RECT 13.04 15.608 16.56 15.64 ;
  LAYER M1 ;
        RECT 13.024 15.588 13.056 15.66 ;
  LAYER M2 ;
        RECT 13.004 15.608 13.076 15.64 ;
  LAYER M1 ;
        RECT 16.544 12.648 16.576 12.72 ;
  LAYER M2 ;
        RECT 16.524 12.668 16.596 12.7 ;
  LAYER M2 ;
        RECT 13.04 12.668 16.56 12.7 ;
  LAYER M1 ;
        RECT 13.024 12.648 13.056 12.72 ;
  LAYER M2 ;
        RECT 13.004 12.668 13.076 12.7 ;
  LAYER M1 ;
        RECT 16.544 9.708 16.576 9.78 ;
  LAYER M2 ;
        RECT 16.524 9.728 16.596 9.76 ;
  LAYER M1 ;
        RECT 16.544 9.744 16.576 12.684 ;
  LAYER M1 ;
        RECT 16.544 12.648 16.576 12.72 ;
  LAYER M2 ;
        RECT 16.524 12.668 16.596 12.7 ;
  LAYER M1 ;
        RECT 16.544 6.768 16.576 6.84 ;
  LAYER M2 ;
        RECT 16.524 6.788 16.596 6.82 ;
  LAYER M1 ;
        RECT 16.544 6.804 16.576 9.744 ;
  LAYER M1 ;
        RECT 16.544 9.708 16.576 9.78 ;
  LAYER M2 ;
        RECT 16.524 9.728 16.596 9.76 ;
  LAYER M1 ;
        RECT 16.544 3.828 16.576 3.9 ;
  LAYER M2 ;
        RECT 16.524 3.848 16.596 3.88 ;
  LAYER M1 ;
        RECT 16.544 3.864 16.576 6.804 ;
  LAYER M1 ;
        RECT 16.544 6.768 16.576 6.84 ;
  LAYER M2 ;
        RECT 16.524 6.788 16.596 6.82 ;
  LAYER M1 ;
        RECT 16.544 0.888 16.576 0.96 ;
  LAYER M2 ;
        RECT 16.524 0.908 16.596 0.94 ;
  LAYER M1 ;
        RECT 16.544 0.924 16.576 3.864 ;
  LAYER M1 ;
        RECT 16.544 3.828 16.576 3.9 ;
  LAYER M2 ;
        RECT 16.524 3.848 16.596 3.88 ;
  LAYER M1 ;
        RECT 7.104 9.204 7.136 9.276 ;
  LAYER M2 ;
        RECT 7.084 9.224 7.156 9.256 ;
  LAYER M2 ;
        RECT 6.64 9.224 7.12 9.256 ;
  LAYER M1 ;
        RECT 6.624 9.204 6.656 9.276 ;
  LAYER M2 ;
        RECT 6.604 9.224 6.676 9.256 ;
  LAYER M1 ;
        RECT 3.584 15.084 3.616 15.156 ;
  LAYER M2 ;
        RECT 3.564 15.104 3.636 15.136 ;
  LAYER M1 ;
        RECT 3.584 15.12 3.616 15.288 ;
  LAYER M1 ;
        RECT 3.584 15.252 3.616 15.324 ;
  LAYER M2 ;
        RECT 3.564 15.272 3.636 15.304 ;
  LAYER M2 ;
        RECT 3.6 15.272 6.64 15.304 ;
  LAYER M1 ;
        RECT 6.624 15.252 6.656 15.324 ;
  LAYER M2 ;
        RECT 6.604 15.272 6.676 15.304 ;
  LAYER M1 ;
        RECT 6.624 18.528 6.656 18.6 ;
  LAYER M2 ;
        RECT 6.604 18.548 6.676 18.58 ;
  LAYER M1 ;
        RECT 6.624 18.396 6.656 18.564 ;
  LAYER M1 ;
        RECT 6.624 9.24 6.656 18.396 ;
  LAYER M1 ;
        RECT 10.624 6.264 10.656 6.336 ;
  LAYER M2 ;
        RECT 10.604 6.284 10.676 6.316 ;
  LAYER M2 ;
        RECT 10.16 6.284 10.64 6.316 ;
  LAYER M1 ;
        RECT 10.144 6.264 10.176 6.336 ;
  LAYER M2 ;
        RECT 10.124 6.284 10.196 6.316 ;
  LAYER M1 ;
        RECT 10.144 18.528 10.176 18.6 ;
  LAYER M2 ;
        RECT 10.124 18.548 10.196 18.58 ;
  LAYER M1 ;
        RECT 10.144 18.396 10.176 18.564 ;
  LAYER M1 ;
        RECT 10.144 6.3 10.176 18.396 ;
  LAYER M2 ;
        RECT 6.64 18.548 10.16 18.58 ;
  LAYER M1 ;
        RECT 3.584 9.204 3.616 9.276 ;
  LAYER M2 ;
        RECT 3.564 9.224 3.636 9.256 ;
  LAYER M1 ;
        RECT 3.584 9.24 3.616 9.408 ;
  LAYER M1 ;
        RECT 3.584 9.372 3.616 9.444 ;
  LAYER M2 ;
        RECT 3.564 9.392 3.636 9.424 ;
  LAYER M2 ;
        RECT 3.6 9.392 6.8 9.424 ;
  LAYER M1 ;
        RECT 6.784 9.372 6.816 9.444 ;
  LAYER M2 ;
        RECT 6.764 9.392 6.836 9.424 ;
  LAYER M1 ;
        RECT 3.584 12.144 3.616 12.216 ;
  LAYER M2 ;
        RECT 3.564 12.164 3.636 12.196 ;
  LAYER M1 ;
        RECT 3.584 12.18 3.616 12.348 ;
  LAYER M1 ;
        RECT 3.584 12.312 3.616 12.384 ;
  LAYER M2 ;
        RECT 3.564 12.332 3.636 12.364 ;
  LAYER M2 ;
        RECT 3.6 12.332 6.8 12.364 ;
  LAYER M1 ;
        RECT 6.784 12.312 6.816 12.384 ;
  LAYER M2 ;
        RECT 6.764 12.332 6.836 12.364 ;
  LAYER M1 ;
        RECT 7.104 6.264 7.136 6.336 ;
  LAYER M2 ;
        RECT 7.084 6.284 7.156 6.316 ;
  LAYER M2 ;
        RECT 6.8 6.284 7.12 6.316 ;
  LAYER M1 ;
        RECT 6.784 6.264 6.816 6.336 ;
  LAYER M2 ;
        RECT 6.764 6.284 6.836 6.316 ;
  LAYER M1 ;
        RECT 7.104 15.084 7.136 15.156 ;
  LAYER M2 ;
        RECT 7.084 15.104 7.156 15.136 ;
  LAYER M2 ;
        RECT 6.8 15.104 7.12 15.136 ;
  LAYER M1 ;
        RECT 6.784 15.084 6.816 15.156 ;
  LAYER M2 ;
        RECT 6.764 15.104 6.836 15.136 ;
  LAYER M1 ;
        RECT 6.784 18.696 6.816 18.768 ;
  LAYER M2 ;
        RECT 6.764 18.716 6.836 18.748 ;
  LAYER M1 ;
        RECT 6.784 18.396 6.816 18.732 ;
  LAYER M1 ;
        RECT 6.784 6.3 6.816 18.396 ;
  LAYER M1 ;
        RECT 10.624 12.144 10.656 12.216 ;
  LAYER M2 ;
        RECT 10.604 12.164 10.676 12.196 ;
  LAYER M2 ;
        RECT 10.32 12.164 10.64 12.196 ;
  LAYER M1 ;
        RECT 10.304 12.144 10.336 12.216 ;
  LAYER M2 ;
        RECT 10.284 12.164 10.356 12.196 ;
  LAYER M1 ;
        RECT 10.624 9.204 10.656 9.276 ;
  LAYER M2 ;
        RECT 10.604 9.224 10.676 9.256 ;
  LAYER M2 ;
        RECT 10.32 9.224 10.64 9.256 ;
  LAYER M1 ;
        RECT 10.304 9.204 10.336 9.276 ;
  LAYER M2 ;
        RECT 10.284 9.224 10.356 9.256 ;
  LAYER M1 ;
        RECT 10.304 18.696 10.336 18.768 ;
  LAYER M2 ;
        RECT 10.284 18.716 10.356 18.748 ;
  LAYER M1 ;
        RECT 10.304 18.396 10.336 18.732 ;
  LAYER M1 ;
        RECT 10.304 9.24 10.336 18.396 ;
  LAYER M2 ;
        RECT 6.8 18.716 10.32 18.748 ;
  LAYER M1 ;
        RECT 3.584 3.324 3.616 3.396 ;
  LAYER M2 ;
        RECT 3.564 3.344 3.636 3.376 ;
  LAYER M1 ;
        RECT 3.584 3.36 3.616 3.528 ;
  LAYER M1 ;
        RECT 3.584 3.492 3.616 3.564 ;
  LAYER M2 ;
        RECT 3.564 3.512 3.636 3.544 ;
  LAYER M2 ;
        RECT 3.6 3.512 6.96 3.544 ;
  LAYER M1 ;
        RECT 6.944 3.492 6.976 3.564 ;
  LAYER M2 ;
        RECT 6.924 3.512 6.996 3.544 ;
  LAYER M1 ;
        RECT 3.584 6.264 3.616 6.336 ;
  LAYER M2 ;
        RECT 3.564 6.284 3.636 6.316 ;
  LAYER M1 ;
        RECT 3.584 6.3 3.616 6.468 ;
  LAYER M1 ;
        RECT 3.584 6.432 3.616 6.504 ;
  LAYER M2 ;
        RECT 3.564 6.452 3.636 6.484 ;
  LAYER M2 ;
        RECT 3.6 6.452 6.96 6.484 ;
  LAYER M1 ;
        RECT 6.944 6.432 6.976 6.504 ;
  LAYER M2 ;
        RECT 6.924 6.452 6.996 6.484 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.06 3.616 18.228 ;
  LAYER M1 ;
        RECT 3.584 18.192 3.616 18.264 ;
  LAYER M2 ;
        RECT 3.564 18.212 3.636 18.244 ;
  LAYER M2 ;
        RECT 3.6 18.212 6.96 18.244 ;
  LAYER M1 ;
        RECT 6.944 18.192 6.976 18.264 ;
  LAYER M2 ;
        RECT 6.924 18.212 6.996 18.244 ;
  LAYER M1 ;
        RECT 7.104 3.324 7.136 3.396 ;
  LAYER M2 ;
        RECT 7.084 3.344 7.156 3.376 ;
  LAYER M2 ;
        RECT 6.96 3.344 7.12 3.376 ;
  LAYER M1 ;
        RECT 6.944 3.324 6.976 3.396 ;
  LAYER M2 ;
        RECT 6.924 3.344 6.996 3.376 ;
  LAYER M1 ;
        RECT 7.104 12.144 7.136 12.216 ;
  LAYER M2 ;
        RECT 7.084 12.164 7.156 12.196 ;
  LAYER M2 ;
        RECT 6.96 12.164 7.12 12.196 ;
  LAYER M1 ;
        RECT 6.944 12.144 6.976 12.216 ;
  LAYER M2 ;
        RECT 6.924 12.164 6.996 12.196 ;
  LAYER M1 ;
        RECT 7.104 18.024 7.136 18.096 ;
  LAYER M2 ;
        RECT 7.084 18.044 7.156 18.076 ;
  LAYER M2 ;
        RECT 6.96 18.044 7.12 18.076 ;
  LAYER M1 ;
        RECT 6.944 18.024 6.976 18.096 ;
  LAYER M2 ;
        RECT 6.924 18.044 6.996 18.076 ;
  LAYER M1 ;
        RECT 6.944 18.864 6.976 18.936 ;
  LAYER M2 ;
        RECT 6.924 18.884 6.996 18.916 ;
  LAYER M1 ;
        RECT 6.944 18.396 6.976 18.9 ;
  LAYER M1 ;
        RECT 6.944 3.36 6.976 18.396 ;
  LAYER M1 ;
        RECT 10.624 3.324 10.656 3.396 ;
  LAYER M2 ;
        RECT 10.604 3.344 10.676 3.376 ;
  LAYER M2 ;
        RECT 10.48 3.344 10.64 3.376 ;
  LAYER M1 ;
        RECT 10.464 3.324 10.496 3.396 ;
  LAYER M2 ;
        RECT 10.444 3.344 10.516 3.376 ;
  LAYER M1 ;
        RECT 10.624 15.084 10.656 15.156 ;
  LAYER M2 ;
        RECT 10.604 15.104 10.676 15.136 ;
  LAYER M2 ;
        RECT 10.48 15.104 10.64 15.136 ;
  LAYER M1 ;
        RECT 10.464 15.084 10.496 15.156 ;
  LAYER M2 ;
        RECT 10.444 15.104 10.516 15.136 ;
  LAYER M1 ;
        RECT 10.624 18.024 10.656 18.096 ;
  LAYER M2 ;
        RECT 10.604 18.044 10.676 18.076 ;
  LAYER M2 ;
        RECT 10.48 18.044 10.64 18.076 ;
  LAYER M1 ;
        RECT 10.464 18.024 10.496 18.096 ;
  LAYER M2 ;
        RECT 10.444 18.044 10.516 18.076 ;
  LAYER M1 ;
        RECT 10.464 18.864 10.496 18.936 ;
  LAYER M2 ;
        RECT 10.444 18.884 10.516 18.916 ;
  LAYER M1 ;
        RECT 10.464 18.396 10.496 18.9 ;
  LAYER M1 ;
        RECT 10.464 3.36 10.496 18.396 ;
  LAYER M2 ;
        RECT 6.96 18.884 10.48 18.916 ;
  LAYER M1 ;
        RECT 0.064 18.024 0.096 18.096 ;
  LAYER M2 ;
        RECT 0.044 18.044 0.116 18.076 ;
  LAYER M2 ;
        RECT 0.08 18.044 3.6 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M1 ;
        RECT 0.064 15.084 0.096 15.156 ;
  LAYER M2 ;
        RECT 0.044 15.104 0.116 15.136 ;
  LAYER M1 ;
        RECT 0.064 15.12 0.096 18.06 ;
  LAYER M1 ;
        RECT 0.064 18.024 0.096 18.096 ;
  LAYER M2 ;
        RECT 0.044 18.044 0.116 18.076 ;
  LAYER M1 ;
        RECT 0.064 12.144 0.096 12.216 ;
  LAYER M2 ;
        RECT 0.044 12.164 0.116 12.196 ;
  LAYER M1 ;
        RECT 0.064 12.18 0.096 15.12 ;
  LAYER M1 ;
        RECT 0.064 15.084 0.096 15.156 ;
  LAYER M2 ;
        RECT 0.044 15.104 0.116 15.136 ;
  LAYER M1 ;
        RECT 0.064 9.204 0.096 9.276 ;
  LAYER M2 ;
        RECT 0.044 9.224 0.116 9.256 ;
  LAYER M1 ;
        RECT 0.064 9.24 0.096 12.18 ;
  LAYER M1 ;
        RECT 0.064 12.144 0.096 12.216 ;
  LAYER M2 ;
        RECT 0.044 12.164 0.116 12.196 ;
  LAYER M1 ;
        RECT 0.064 6.264 0.096 6.336 ;
  LAYER M2 ;
        RECT 0.044 6.284 0.116 6.316 ;
  LAYER M1 ;
        RECT 0.064 6.3 0.096 9.24 ;
  LAYER M1 ;
        RECT 0.064 9.204 0.096 9.276 ;
  LAYER M2 ;
        RECT 0.044 9.224 0.116 9.256 ;
  LAYER M1 ;
        RECT 0.064 3.324 0.096 3.396 ;
  LAYER M2 ;
        RECT 0.044 3.344 0.116 3.376 ;
  LAYER M1 ;
        RECT 0.064 3.36 0.096 6.3 ;
  LAYER M1 ;
        RECT 0.064 6.264 0.096 6.336 ;
  LAYER M2 ;
        RECT 0.044 6.284 0.116 6.316 ;
  LAYER M1 ;
        RECT 14.144 18.024 14.176 18.096 ;
  LAYER M2 ;
        RECT 14.124 18.044 14.196 18.076 ;
  LAYER M2 ;
        RECT 10.64 18.044 14.16 18.076 ;
  LAYER M1 ;
        RECT 10.624 18.024 10.656 18.096 ;
  LAYER M2 ;
        RECT 10.604 18.044 10.676 18.076 ;
  LAYER M1 ;
        RECT 14.144 15.084 14.176 15.156 ;
  LAYER M2 ;
        RECT 14.124 15.104 14.196 15.136 ;
  LAYER M2 ;
        RECT 10.64 15.104 14.16 15.136 ;
  LAYER M1 ;
        RECT 10.624 15.084 10.656 15.156 ;
  LAYER M2 ;
        RECT 10.604 15.104 10.676 15.136 ;
  LAYER M1 ;
        RECT 14.144 12.144 14.176 12.216 ;
  LAYER M2 ;
        RECT 14.124 12.164 14.196 12.196 ;
  LAYER M1 ;
        RECT 14.144 12.18 14.176 15.12 ;
  LAYER M1 ;
        RECT 14.144 15.084 14.176 15.156 ;
  LAYER M2 ;
        RECT 14.124 15.104 14.196 15.136 ;
  LAYER M1 ;
        RECT 14.144 9.204 14.176 9.276 ;
  LAYER M2 ;
        RECT 14.124 9.224 14.196 9.256 ;
  LAYER M1 ;
        RECT 14.144 9.24 14.176 12.18 ;
  LAYER M1 ;
        RECT 14.144 12.144 14.176 12.216 ;
  LAYER M2 ;
        RECT 14.124 12.164 14.196 12.196 ;
  LAYER M1 ;
        RECT 14.144 6.264 14.176 6.336 ;
  LAYER M2 ;
        RECT 14.124 6.284 14.196 6.316 ;
  LAYER M1 ;
        RECT 14.144 6.3 14.176 9.24 ;
  LAYER M1 ;
        RECT 14.144 9.204 14.176 9.276 ;
  LAYER M2 ;
        RECT 14.124 9.224 14.196 9.256 ;
  LAYER M1 ;
        RECT 14.144 3.324 14.176 3.396 ;
  LAYER M2 ;
        RECT 14.124 3.344 14.196 3.376 ;
  LAYER M1 ;
        RECT 14.144 3.36 14.176 6.3 ;
  LAYER M1 ;
        RECT 14.144 6.264 14.176 6.336 ;
  LAYER M2 ;
        RECT 14.124 6.284 14.196 6.316 ;
  LAYER M1 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M2 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M3 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M1 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M2 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M3 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M1 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M2 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M3 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M1 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M2 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M3 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M1 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M2 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M3 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M1 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M2 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M3 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M1 ;
        RECT 3.6 0.924 6 3.36 ;
  LAYER M2 ;
        RECT 3.6 0.924 6 3.36 ;
  LAYER M3 ;
        RECT 3.6 0.924 6 3.36 ;
  LAYER M1 ;
        RECT 3.6 3.864 6 6.3 ;
  LAYER M2 ;
        RECT 3.6 3.864 6 6.3 ;
  LAYER M3 ;
        RECT 3.6 3.864 6 6.3 ;
  LAYER M1 ;
        RECT 3.6 6.804 6 9.24 ;
  LAYER M2 ;
        RECT 3.6 6.804 6 9.24 ;
  LAYER M3 ;
        RECT 3.6 6.804 6 9.24 ;
  LAYER M1 ;
        RECT 3.6 9.744 6 12.18 ;
  LAYER M2 ;
        RECT 3.6 9.744 6 12.18 ;
  LAYER M3 ;
        RECT 3.6 9.744 6 12.18 ;
  LAYER M1 ;
        RECT 3.6 12.684 6 15.12 ;
  LAYER M2 ;
        RECT 3.6 12.684 6 15.12 ;
  LAYER M3 ;
        RECT 3.6 12.684 6 15.12 ;
  LAYER M1 ;
        RECT 3.6 15.624 6 18.06 ;
  LAYER M2 ;
        RECT 3.6 15.624 6 18.06 ;
  LAYER M3 ;
        RECT 3.6 15.624 6 18.06 ;
  LAYER M1 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M2 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M3 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M1 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M2 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M3 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M1 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M2 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M3 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M1 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M2 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M3 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M1 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M2 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M3 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M1 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M2 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M3 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M1 ;
        RECT 10.64 0.924 13.04 3.36 ;
  LAYER M2 ;
        RECT 10.64 0.924 13.04 3.36 ;
  LAYER M3 ;
        RECT 10.64 0.924 13.04 3.36 ;
  LAYER M1 ;
        RECT 10.64 3.864 13.04 6.3 ;
  LAYER M2 ;
        RECT 10.64 3.864 13.04 6.3 ;
  LAYER M3 ;
        RECT 10.64 3.864 13.04 6.3 ;
  LAYER M1 ;
        RECT 10.64 6.804 13.04 9.24 ;
  LAYER M2 ;
        RECT 10.64 6.804 13.04 9.24 ;
  LAYER M3 ;
        RECT 10.64 6.804 13.04 9.24 ;
  LAYER M1 ;
        RECT 10.64 9.744 13.04 12.18 ;
  LAYER M2 ;
        RECT 10.64 9.744 13.04 12.18 ;
  LAYER M3 ;
        RECT 10.64 9.744 13.04 12.18 ;
  LAYER M1 ;
        RECT 10.64 12.684 13.04 15.12 ;
  LAYER M2 ;
        RECT 10.64 12.684 13.04 15.12 ;
  LAYER M3 ;
        RECT 10.64 12.684 13.04 15.12 ;
  LAYER M1 ;
        RECT 10.64 15.624 13.04 18.06 ;
  LAYER M2 ;
        RECT 10.64 15.624 13.04 18.06 ;
  LAYER M3 ;
        RECT 10.64 15.624 13.04 18.06 ;
  LAYER M1 ;
        RECT 14.16 0.924 16.56 3.36 ;
  LAYER M2 ;
        RECT 14.16 0.924 16.56 3.36 ;
  LAYER M3 ;
        RECT 14.16 0.924 16.56 3.36 ;
  LAYER M1 ;
        RECT 14.16 3.864 16.56 6.3 ;
  LAYER M2 ;
        RECT 14.16 3.864 16.56 6.3 ;
  LAYER M3 ;
        RECT 14.16 3.864 16.56 6.3 ;
  LAYER M1 ;
        RECT 14.16 6.804 16.56 9.24 ;
  LAYER M2 ;
        RECT 14.16 6.804 16.56 9.24 ;
  LAYER M3 ;
        RECT 14.16 6.804 16.56 9.24 ;
  LAYER M1 ;
        RECT 14.16 9.744 16.56 12.18 ;
  LAYER M2 ;
        RECT 14.16 9.744 16.56 12.18 ;
  LAYER M3 ;
        RECT 14.16 9.744 16.56 12.18 ;
  LAYER M1 ;
        RECT 14.16 12.684 16.56 15.12 ;
  LAYER M2 ;
        RECT 14.16 12.684 16.56 15.12 ;
  LAYER M3 ;
        RECT 14.16 12.684 16.56 15.12 ;
  LAYER M1 ;
        RECT 14.16 15.624 16.56 18.06 ;
  LAYER M2 ;
        RECT 14.16 15.624 16.56 18.06 ;
  LAYER M3 ;
        RECT 14.16 15.624 16.56 18.06 ;
  END 
END Cap_30fF_Cap_60fF
