MACRO switched_capacitor_filter
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_filter 0 0 ;
  SIZE 47.52 BY 39.48 ;
  PIN id
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.664 -0.016 23.696 0.016 ;
      LAYER M2 ;
        RECT 23.324 0.32 24.116 0.352 ;
      LAYER M2 ;
        RECT 23.744 0.32 23.776 0.352 ;
      LAYER M3 ;
        RECT 23.74 0.316 23.78 0.356 ;
      LAYER M4 ;
        RECT 23.74 0.316 23.78 0.356 ;
      LAYER M5 ;
        RECT 23.728 0 23.792 0.336 ;
      LAYER M4 ;
        RECT 23.76 -0.02 23.92 0.02 ;
      LAYER M3 ;
        RECT 23.9 -0.02 23.94 0.02 ;
      LAYER M2 ;
        RECT 23.68 -0.016 23.92 0.016 ;
    END
  END id
  PIN voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.824 39.464 15.856 39.496 ;
      LAYER M2 ;
        RECT 22.844 4.436 24.676 4.468 ;
      LAYER M2 ;
        RECT 22.684 3.008 25.316 3.04 ;
      LAYER M2 ;
        RECT 23.424 4.436 23.456 4.468 ;
      LAYER M3 ;
        RECT 23.42 3.192 23.46 4.452 ;
      LAYER M4 ;
        RECT 23.28 3.172 23.44 3.212 ;
      LAYER M5 ;
        RECT 23.248 3.024 23.312 3.192 ;
      LAYER M4 ;
        RECT 23.26 3.004 23.3 3.044 ;
      LAYER M3 ;
        RECT 23.26 3.004 23.3 3.044 ;
      LAYER M2 ;
        RECT 23.264 3.008 23.296 3.04 ;
      LAYER M2 ;
        RECT 7.964 0.824 8.036 0.856 ;
      LAYER M1 ;
        RECT 12.128 14.832 12.16 14.904 ;
      LAYER M2 ;
        RECT 12.108 14.852 12.18 14.884 ;
      LAYER M1 ;
        RECT 3.2 14.832 3.232 14.904 ;
      LAYER M2 ;
        RECT 3.18 14.852 3.252 14.884 ;
      LAYER M2 ;
        RECT 3.216 14.852 12.144 14.884 ;
      LAYER M2 ;
        RECT 7.984 0.824 8.016 0.856 ;
      LAYER M3 ;
        RECT 7.98 0.84 8.02 1.596 ;
      LAYER M4 ;
        RECT 7.84 1.576 8 1.616 ;
      LAYER M3 ;
        RECT 7.82 1.596 7.86 14.7 ;
      LAYER M4 ;
        RECT 7.84 14.68 8.16 14.72 ;
      LAYER M5 ;
        RECT 8.128 14.7 8.192 14.868 ;
      LAYER M4 ;
        RECT 8.14 14.848 8.18 14.888 ;
      LAYER M3 ;
        RECT 8.14 14.848 8.18 14.888 ;
      LAYER M2 ;
        RECT 8.144 14.852 8.176 14.884 ;
      LAYER M1 ;
        RECT 22.176 39.024 22.208 39.096 ;
      LAYER M2 ;
        RECT 22.156 39.044 22.228 39.076 ;
      LAYER M1 ;
        RECT 25.152 39.024 25.184 39.096 ;
      LAYER M2 ;
        RECT 25.132 39.044 25.204 39.076 ;
      LAYER M2 ;
        RECT 22.192 39.044 25.168 39.076 ;
      LAYER M2 ;
        RECT 15.28 3.008 22.72 3.04 ;
      LAYER M3 ;
        RECT 15.26 3.004 15.3 3.044 ;
      LAYER M4 ;
        RECT 7.84 3.004 15.28 3.044 ;
      LAYER M3 ;
        RECT 7.82 3.004 7.86 3.044 ;
      LAYER M2 ;
        RECT 12.16 14.852 12.4 14.884 ;
      LAYER M3 ;
        RECT 12.38 14.868 12.42 39.06 ;
      LAYER M2 ;
        RECT 12.4 39.044 22.24 39.076 ;
      LAYER M2 ;
        RECT 15.824 39.044 15.856 39.076 ;
      LAYER M3 ;
        RECT 15.82 39.06 15.86 39.312 ;
      LAYER M4 ;
        RECT 15.82 39.292 15.86 39.332 ;
      LAYER M5 ;
        RECT 15.808 39.312 15.872 39.48 ;
      LAYER M4 ;
        RECT 15.82 39.46 15.86 39.5 ;
      LAYER M3 ;
        RECT 15.82 39.46 15.86 39.5 ;
      LAYER M2 ;
        RECT 15.824 39.464 15.856 39.496 ;
    END
  END voutn
  PIN voutp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.664 39.464 31.696 39.496 ;
      LAYER M2 ;
        RECT 23.484 4.268 24.036 4.3 ;
      LAYER M2 ;
        RECT 22.044 3.176 24.676 3.208 ;
      LAYER M2 ;
        RECT 23.584 4.268 23.616 4.3 ;
      LAYER M3 ;
        RECT 23.58 4.032 23.62 4.284 ;
      LAYER M4 ;
        RECT 23.28 4.012 23.6 4.052 ;
      LAYER M5 ;
        RECT 23.248 3.696 23.312 4.032 ;
      LAYER M4 ;
        RECT 23.26 3.676 23.3 3.716 ;
      LAYER M3 ;
        RECT 23.26 3.192 23.3 3.696 ;
      LAYER M2 ;
        RECT 23.264 3.176 23.296 3.208 ;
      LAYER M2 ;
        RECT 39.484 0.824 39.556 0.856 ;
      LAYER M1 ;
        RECT 35.36 14.832 35.392 14.904 ;
      LAYER M2 ;
        RECT 35.34 14.852 35.412 14.884 ;
      LAYER M1 ;
        RECT 44.288 14.832 44.32 14.904 ;
      LAYER M2 ;
        RECT 44.268 14.852 44.34 14.884 ;
      LAYER M2 ;
        RECT 35.376 14.852 44.304 14.884 ;
      LAYER M2 ;
        RECT 39.504 0.824 39.536 0.856 ;
      LAYER M3 ;
        RECT 39.5 0.84 39.54 1.596 ;
      LAYER M4 ;
        RECT 39.52 1.576 39.68 1.616 ;
      LAYER M3 ;
        RECT 39.66 1.596 39.7 14.7 ;
      LAYER M4 ;
        RECT 39.36 14.68 39.68 14.72 ;
      LAYER M5 ;
        RECT 39.328 14.7 39.392 14.868 ;
      LAYER M4 ;
        RECT 39.34 14.848 39.38 14.888 ;
      LAYER M3 ;
        RECT 39.34 14.848 39.38 14.888 ;
      LAYER M2 ;
        RECT 39.344 14.852 39.376 14.884 ;
      LAYER M1 ;
        RECT 19.2 39.192 19.232 39.264 ;
      LAYER M2 ;
        RECT 19.18 39.212 19.252 39.244 ;
      LAYER M1 ;
        RECT 28.128 39.192 28.16 39.264 ;
      LAYER M2 ;
        RECT 28.108 39.212 28.18 39.244 ;
      LAYER M2 ;
        RECT 19.216 39.212 28.144 39.244 ;
      LAYER M2 ;
        RECT 24 4.268 31.68 4.3 ;
      LAYER M3 ;
        RECT 31.66 4.264 31.7 4.304 ;
      LAYER M4 ;
        RECT 31.68 4.264 39.68 4.304 ;
      LAYER M3 ;
        RECT 39.66 4.264 39.7 4.304 ;
      LAYER M2 ;
        RECT 31.28 14.852 35.36 14.884 ;
      LAYER M3 ;
        RECT 31.26 14.868 31.3 38.304 ;
      LAYER M4 ;
        RECT 28.8 38.284 31.28 38.324 ;
      LAYER M5 ;
        RECT 28.768 38.304 28.832 39.228 ;
      LAYER M4 ;
        RECT 28.78 39.208 28.82 39.248 ;
      LAYER M3 ;
        RECT 28.78 39.208 28.82 39.248 ;
      LAYER M2 ;
        RECT 28.08 39.212 28.8 39.244 ;
      LAYER M4 ;
        RECT 31.248 38.284 31.68 38.324 ;
      LAYER M5 ;
        RECT 31.648 38.304 31.712 39.48 ;
      LAYER M4 ;
        RECT 31.66 39.46 31.7 39.5 ;
      LAYER M3 ;
        RECT 31.66 39.46 31.7 39.5 ;
      LAYER M2 ;
        RECT 31.664 39.464 31.696 39.496 ;
    END
  END voutp
  PIN vss
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 24.064 -0.016 24.096 0.016 ;
      LAYER M2 ;
        RECT 21.564 0.236 26.116 0.268 ;
      LAYER M1 ;
        RECT 22.336 19.872 22.368 19.944 ;
      LAYER M2 ;
        RECT 22.316 19.892 22.388 19.924 ;
      LAYER M1 ;
        RECT 25.312 19.872 25.344 19.944 ;
      LAYER M2 ;
        RECT 25.292 19.892 25.364 19.924 ;
      LAYER M2 ;
        RECT 22.352 19.892 25.328 19.924 ;
      LAYER M1 ;
        RECT 19.36 19.704 19.392 19.776 ;
      LAYER M2 ;
        RECT 19.34 19.724 19.412 19.756 ;
      LAYER M1 ;
        RECT 28.288 19.704 28.32 19.776 ;
      LAYER M2 ;
        RECT 28.268 19.724 28.34 19.756 ;
      LAYER M2 ;
        RECT 19.376 19.724 28.304 19.756 ;
      LAYER M2 ;
        RECT 24.064 0.236 24.096 0.268 ;
      LAYER M3 ;
        RECT 24.06 0 24.1 0.252 ;
      LAYER M2 ;
        RECT 24.064 -0.016 24.096 0.016 ;
      LAYER M3 ;
        RECT 24.06 0.252 24.1 19.908 ;
      LAYER M2 ;
        RECT 24.064 19.892 24.096 19.924 ;
      LAYER M3 ;
        RECT 24.06 19.72 24.1 19.76 ;
      LAYER M2 ;
        RECT 24.064 19.724 24.096 19.756 ;
    END
  END vss
  PIN vinn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.744 -0.016 15.776 0.016 ;
      LAYER M2 ;
        RECT 15.724 0.236 15.796 0.268 ;
      LAYER M1 ;
        RECT 28.288 5.844 28.32 5.916 ;
      LAYER M2 ;
        RECT 28.268 5.864 28.34 5.896 ;
      LAYER M1 ;
        RECT 19.36 5.844 19.392 5.916 ;
      LAYER M2 ;
        RECT 19.34 5.864 19.412 5.896 ;
      LAYER M2 ;
        RECT 19.376 5.864 28.304 5.896 ;
      LAYER M2 ;
        RECT 15.744 0.236 15.776 0.268 ;
      LAYER M3 ;
        RECT 15.74 0 15.78 0.252 ;
      LAYER M2 ;
        RECT 15.744 -0.016 15.776 0.016 ;
      LAYER M3 ;
        RECT 15.74 0.084 15.78 1.596 ;
      LAYER M2 ;
        RECT 15.76 1.58 19.36 1.612 ;
      LAYER M3 ;
        RECT 19.34 1.596 19.38 5.88 ;
      LAYER M2 ;
        RECT 19.344 5.864 19.376 5.896 ;
    END
  END vinn
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.904 -0.016 15.936 0.016 ;
      LAYER M2 ;
        RECT 5.244 0.236 5.316 0.268 ;
      LAYER M2 ;
        RECT 5.964 0.74 6.036 0.772 ;
      LAYER M2 ;
        RECT 7.324 0.74 7.396 0.772 ;
      LAYER M2 ;
        RECT 5.28 0.236 6 0.268 ;
      LAYER M3 ;
        RECT 5.98 0.252 6.02 0.756 ;
      LAYER M2 ;
        RECT 5.984 0.74 6.016 0.772 ;
      LAYER M2 ;
        RECT 6 0.74 7.2 0.772 ;
      LAYER M3 ;
        RECT 7.18 0.736 7.22 0.776 ;
      LAYER M4 ;
        RECT 7.2 0.736 7.36 0.776 ;
      LAYER M3 ;
        RECT 7.34 0.736 7.38 0.776 ;
      LAYER M2 ;
        RECT 7.344 0.74 7.376 0.772 ;
      LAYER M2 ;
        RECT 42.204 0.236 42.276 0.268 ;
      LAYER M2 ;
        RECT 41.484 0.74 41.556 0.772 ;
      LAYER M2 ;
        RECT 40.124 0.74 40.196 0.772 ;
      LAYER M2 ;
        RECT 41.52 0.236 42.24 0.268 ;
      LAYER M3 ;
        RECT 41.5 0.252 41.54 0.756 ;
      LAYER M2 ;
        RECT 41.504 0.74 41.536 0.772 ;
      LAYER M2 ;
        RECT 40.32 0.74 41.52 0.772 ;
      LAYER M3 ;
        RECT 40.3 0.736 40.34 0.776 ;
      LAYER M4 ;
        RECT 40.16 0.736 40.32 0.776 ;
      LAYER M3 ;
        RECT 40.14 0.736 40.18 0.776 ;
      LAYER M2 ;
        RECT 40.144 0.74 40.176 0.772 ;
      LAYER M4 ;
        RECT 7.344 0.736 7.92 0.776 ;
      LAYER M5 ;
        RECT 7.888 0.756 7.952 3.36 ;
      LAYER M4 ;
        RECT 7.92 3.34 15.12 3.38 ;
      LAYER M5 ;
        RECT 15.088 0 15.152 3.36 ;
      LAYER M4 ;
        RECT 15.12 -0.02 15.92 0.02 ;
      LAYER M3 ;
        RECT 15.9 -0.02 15.94 0.02 ;
      LAYER M2 ;
        RECT 15.904 -0.016 15.936 0.016 ;
      LAYER M5 ;
        RECT 15.088 3.312 15.152 3.456 ;
      LAYER M6 ;
        RECT 15.12 3.424 17.28 3.488 ;
      LAYER M5 ;
        RECT 17.248 3.456 17.312 5.04 ;
      LAYER M4 ;
        RECT 17.28 5.02 41.616 5.06 ;
      LAYER M5 ;
        RECT 41.584 1.764 41.648 5.04 ;
      LAYER M4 ;
        RECT 41.616 1.744 41.76 1.784 ;
      LAYER M3 ;
        RECT 41.74 1.512 41.78 1.764 ;
      LAYER M2 ;
        RECT 41.52 1.496 41.76 1.528 ;
      LAYER M3 ;
        RECT 41.5 0.756 41.54 1.512 ;
    END
  END agnd
  PIN vinp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.744 -0.016 31.776 0.016 ;
      LAYER M2 ;
        RECT 31.724 0.236 31.796 0.268 ;
      LAYER M1 ;
        RECT 25.312 6.012 25.344 6.084 ;
      LAYER M2 ;
        RECT 25.292 6.032 25.364 6.064 ;
      LAYER M1 ;
        RECT 22.336 6.012 22.368 6.084 ;
      LAYER M2 ;
        RECT 22.316 6.032 22.388 6.064 ;
      LAYER M2 ;
        RECT 22.352 6.032 25.328 6.064 ;
      LAYER M2 ;
        RECT 30.56 0.236 31.76 0.268 ;
      LAYER M3 ;
        RECT 30.54 0.252 30.58 3.276 ;
      LAYER M2 ;
        RECT 25.76 3.26 30.56 3.292 ;
      LAYER M3 ;
        RECT 25.74 3.276 25.78 6.048 ;
      LAYER M2 ;
        RECT 25.28 6.032 25.76 6.064 ;
      LAYER M2 ;
        RECT 31.744 0.236 31.776 0.268 ;
      LAYER M3 ;
        RECT 31.74 0 31.78 0.252 ;
      LAYER M2 ;
        RECT 31.744 -0.016 31.776 0.016 ;
    END
  END vinp
  OBS 
  LAYER M2 ;
        RECT 22.124 3.26 25.396 3.292 ;
  LAYER M2 ;
        RECT 21.484 0.488 26.036 0.52 ;
  LAYER M2 ;
        RECT 23.404 5.024 24.116 5.056 ;
  LAYER M2 ;
        RECT 22.764 4.184 24.756 4.216 ;
  LAYER M2 ;
        RECT 23.484 4.772 24.196 4.804 ;
  LAYER M3 ;
        RECT 23.5 1.56 23.54 2.472 ;
  LAYER M2 ;
        RECT 40.844 0.824 40.916 0.856 ;
  LAYER M1 ;
        RECT 35.2 31.212 35.232 31.284 ;
  LAYER M2 ;
        RECT 35.18 31.232 35.252 31.264 ;
  LAYER M1 ;
        RECT 44.128 31.212 44.16 31.284 ;
  LAYER M2 ;
        RECT 44.108 31.232 44.18 31.264 ;
  LAYER M2 ;
        RECT 35.216 31.232 44.144 31.264 ;
  LAYER M2 ;
        RECT 40.88 0.824 41.12 0.856 ;
  LAYER M3 ;
        RECT 41.1 0.84 41.14 31.08 ;
  LAYER M4 ;
        RECT 40.8 31.06 41.12 31.1 ;
  LAYER M5 ;
        RECT 40.768 31.08 40.832 31.248 ;
  LAYER M4 ;
        RECT 40.78 31.228 40.82 31.268 ;
  LAYER M3 ;
        RECT 40.78 31.228 40.82 31.268 ;
  LAYER M2 ;
        RECT 40.784 31.232 40.816 31.264 ;
  LAYER M1 ;
        RECT 28.128 19.116 28.16 19.188 ;
  LAYER M2 ;
        RECT 28.108 19.136 28.18 19.168 ;
  LAYER M1 ;
        RECT 19.2 19.116 19.232 19.188 ;
  LAYER M2 ;
        RECT 19.18 19.136 19.252 19.168 ;
  LAYER M2 ;
        RECT 19.216 19.136 28.144 19.168 ;
  LAYER M3 ;
        RECT 23.5 2.416 23.54 2.456 ;
  LAYER M4 ;
        RECT 23.52 2.416 24 2.456 ;
  LAYER M3 ;
        RECT 23.98 2.436 24.02 3.444 ;
  LAYER M2 ;
        RECT 24 3.428 31.68 3.46 ;
  LAYER M3 ;
        RECT 31.66 3.424 31.7 3.464 ;
  LAYER M4 ;
        RECT 31.68 3.424 41.12 3.464 ;
  LAYER M3 ;
        RECT 41.1 3.424 41.14 3.464 ;
  LAYER M2 ;
        RECT 24.464 3.428 24.496 3.46 ;
  LAYER M3 ;
        RECT 24.46 3.444 24.5 6.216 ;
  LAYER M4 ;
        RECT 24.46 6.196 24.5 6.236 ;
  LAYER M5 ;
        RECT 24.448 6.216 24.512 19.152 ;
  LAYER M4 ;
        RECT 24.46 19.132 24.5 19.172 ;
  LAYER M3 ;
        RECT 24.46 19.132 24.5 19.172 ;
  LAYER M2 ;
        RECT 24.464 19.136 24.496 19.168 ;
  LAYER M3 ;
        RECT 23.82 1.476 23.86 2.388 ;
  LAYER M2 ;
        RECT 6.604 0.824 6.676 0.856 ;
  LAYER M1 ;
        RECT 12.288 31.212 12.32 31.284 ;
  LAYER M2 ;
        RECT 12.268 31.232 12.34 31.264 ;
  LAYER M1 ;
        RECT 3.36 31.212 3.392 31.284 ;
  LAYER M2 ;
        RECT 3.34 31.232 3.412 31.264 ;
  LAYER M2 ;
        RECT 3.376 31.232 12.304 31.264 ;
  LAYER M2 ;
        RECT 6.4 0.824 6.64 0.856 ;
  LAYER M3 ;
        RECT 6.38 0.84 6.42 31.08 ;
  LAYER M4 ;
        RECT 6.4 31.06 6.72 31.1 ;
  LAYER M5 ;
        RECT 6.688 31.08 6.752 31.248 ;
  LAYER M4 ;
        RECT 6.7 31.228 6.74 31.268 ;
  LAYER M3 ;
        RECT 6.7 31.228 6.74 31.268 ;
  LAYER M2 ;
        RECT 6.704 31.232 6.736 31.264 ;
  LAYER M1 ;
        RECT 25.152 18.948 25.184 19.02 ;
  LAYER M2 ;
        RECT 25.132 18.968 25.204 19 ;
  LAYER M1 ;
        RECT 22.176 18.948 22.208 19.02 ;
  LAYER M2 ;
        RECT 22.156 18.968 22.228 19 ;
  LAYER M2 ;
        RECT 22.192 18.968 25.168 19 ;
  LAYER M3 ;
        RECT 23.82 1.492 23.86 1.532 ;
  LAYER M4 ;
        RECT 23.2 1.492 23.84 1.532 ;
  LAYER M3 ;
        RECT 23.18 1.492 23.22 1.532 ;
  LAYER M2 ;
        RECT 6.4 1.496 23.2 1.528 ;
  LAYER M3 ;
        RECT 6.38 1.492 6.42 1.532 ;
  LAYER M3 ;
        RECT 6.38 18.46 6.42 18.5 ;
  LAYER M2 ;
        RECT 6.4 18.464 16.24 18.496 ;
  LAYER M3 ;
        RECT 16.22 18.48 16.26 18.984 ;
  LAYER M2 ;
        RECT 16.24 18.968 22.24 19 ;
  LAYER M2 ;
        RECT 15.644 0.404 15.716 0.436 ;
  LAYER M2 ;
        RECT 6.684 0.656 6.756 0.688 ;
  LAYER M2 ;
        RECT 8.044 0.656 8.116 0.688 ;
  LAYER M2 ;
        RECT 8.48 0.404 15.68 0.436 ;
  LAYER M3 ;
        RECT 8.46 0.42 8.5 0.672 ;
  LAYER M4 ;
        RECT 8.32 0.652 8.48 0.692 ;
  LAYER M3 ;
        RECT 8.3 0.652 8.34 0.692 ;
  LAYER M2 ;
        RECT 8.08 0.656 8.32 0.688 ;
  LAYER M2 ;
        RECT 6.72 0.656 8.16 0.688 ;
  LAYER M2 ;
        RECT 31.804 0.404 31.876 0.436 ;
  LAYER M2 ;
        RECT 40.764 0.656 40.836 0.688 ;
  LAYER M2 ;
        RECT 39.404 0.656 39.476 0.688 ;
  LAYER M2 ;
        RECT 31.84 0.404 39.04 0.436 ;
  LAYER M3 ;
        RECT 39.02 0.42 39.06 0.672 ;
  LAYER M4 ;
        RECT 39.04 0.652 39.2 0.692 ;
  LAYER M3 ;
        RECT 39.18 0.652 39.22 0.692 ;
  LAYER M2 ;
        RECT 39.2 0.656 39.44 0.688 ;
  LAYER M2 ;
        RECT 39.36 0.656 40.8 0.688 ;
  LAYER M2 ;
        RECT 14.384 0.404 14.416 0.436 ;
  LAYER M3 ;
        RECT 14.38 0.42 14.42 4.2 ;
  LAYER M4 ;
        RECT 14.4 4.18 15.984 4.22 ;
  LAYER M5 ;
        RECT 15.952 4.2 16.016 5.208 ;
  LAYER M4 ;
        RECT 15.984 5.188 17.28 5.228 ;
  LAYER M5 ;
        RECT 17.248 5.208 17.312 6.72 ;
  LAYER M4 ;
        RECT 17.28 6.7 31.68 6.74 ;
  LAYER M5 ;
        RECT 31.648 1.176 31.712 6.72 ;
  LAYER M4 ;
        RECT 31.68 1.156 31.84 1.196 ;
  LAYER M3 ;
        RECT 31.82 0.42 31.86 1.176 ;
  LAYER M2 ;
        RECT 31.824 0.404 31.856 0.436 ;
  LAYER M2 ;
        RECT 5.324 0.404 5.396 0.436 ;
  LAYER M2 ;
        RECT 6.044 0.572 6.116 0.604 ;
  LAYER M2 ;
        RECT 7.404 0.572 7.476 0.604 ;
  LAYER M2 ;
        RECT 5.36 0.404 5.84 0.436 ;
  LAYER M3 ;
        RECT 5.82 0.4 5.86 0.44 ;
  LAYER M4 ;
        RECT 5.84 0.4 6 0.44 ;
  LAYER M5 ;
        RECT 5.968 0.42 6.032 0.588 ;
  LAYER M4 ;
        RECT 5.84 0.568 6 0.608 ;
  LAYER M3 ;
        RECT 5.82 0.568 5.86 0.608 ;
  LAYER M2 ;
        RECT 5.84 0.572 6.08 0.604 ;
  LAYER M2 ;
        RECT 6 0.572 7.44 0.604 ;
  LAYER M2 ;
        RECT 42.124 0.404 42.196 0.436 ;
  LAYER M2 ;
        RECT 41.404 0.572 41.476 0.604 ;
  LAYER M2 ;
        RECT 40.044 0.572 40.116 0.604 ;
  LAYER M2 ;
        RECT 41.68 0.404 42.16 0.436 ;
  LAYER M3 ;
        RECT 41.66 0.4 41.7 0.44 ;
  LAYER M4 ;
        RECT 41.52 0.4 41.68 0.44 ;
  LAYER M5 ;
        RECT 41.488 0.42 41.552 0.588 ;
  LAYER M4 ;
        RECT 41.52 0.568 41.68 0.608 ;
  LAYER M3 ;
        RECT 41.66 0.568 41.7 0.608 ;
  LAYER M2 ;
        RECT 41.44 0.572 41.68 0.604 ;
  LAYER M2 ;
        RECT 40.08 0.572 41.52 0.604 ;
  LAYER M2 ;
        RECT 7.44 0.572 40.08 0.604 ;
  LAYER M2 ;
        RECT 23.964 4.856 24.036 4.888 ;
  LAYER M2 ;
        RECT 23.324 4.352 24.196 4.384 ;
  LAYER M2 ;
        RECT 23.984 4.856 24.016 4.888 ;
  LAYER M3 ;
        RECT 23.98 4.368 24.02 4.872 ;
  LAYER M2 ;
        RECT 23.984 4.352 24.016 4.384 ;
  LAYER M2 ;
        RECT 23.324 4.94 23.396 4.972 ;
  LAYER M2 ;
        RECT 22.684 4.52 24.836 4.552 ;
  LAYER M2 ;
        RECT 23.36 4.94 23.6 4.972 ;
  LAYER M3 ;
        RECT 23.58 4.704 23.62 4.956 ;
  LAYER M4 ;
        RECT 23.28 4.684 23.6 4.724 ;
  LAYER M5 ;
        RECT 23.248 4.536 23.312 4.704 ;
  LAYER M4 ;
        RECT 23.26 4.516 23.3 4.556 ;
  LAYER M3 ;
        RECT 23.26 4.516 23.3 4.556 ;
  LAYER M2 ;
        RECT 23.264 4.52 23.296 4.552 ;
  LAYER M3 ;
        RECT 23.58 1.728 23.62 2.64 ;
  LAYER M2 ;
        RECT 22.204 3.092 24.836 3.124 ;
  LAYER M3 ;
        RECT 23.58 2.604 23.62 3.108 ;
  LAYER M2 ;
        RECT 23.584 3.092 23.616 3.124 ;
  LAYER M3 ;
        RECT 23.66 1.812 23.7 2.724 ;
  LAYER M2 ;
        RECT 21.404 0.404 25.956 0.436 ;
  LAYER M3 ;
        RECT 23.66 0.42 23.7 1.932 ;
  LAYER M2 ;
        RECT 23.664 0.404 23.696 0.436 ;
  LAYER M3 ;
        RECT 23.74 1.644 23.78 2.556 ;
  LAYER M2 ;
        RECT 22.844 2.924 25.476 2.956 ;
  LAYER M3 ;
        RECT 23.74 2.436 23.78 2.94 ;
  LAYER M2 ;
        RECT 23.744 2.924 23.776 2.956 ;
  LAYER M1 ;
        RECT 24.064 4.752 24.096 5.412 ;
  LAYER M1 ;
        RECT 23.424 4.752 23.456 5.412 ;
  LAYER M1 ;
        RECT 24.144 4.752 24.176 5.412 ;
  LAYER M1 ;
        RECT 23.504 4.752 23.536 5.412 ;
  LAYER M1 ;
        RECT 23.984 4.752 24.016 5.412 ;
  LAYER M1 ;
        RECT 23.344 5.192 23.376 5.224 ;
  LAYER M1 ;
        RECT 22.144 2.064 22.176 2.724 ;
  LAYER M1 ;
        RECT 22.144 1.224 22.176 1.884 ;
  LAYER M1 ;
        RECT 23.424 2.064 23.456 2.724 ;
  LAYER M1 ;
        RECT 23.424 1.224 23.456 1.884 ;
  LAYER M1 ;
        RECT 24.704 2.064 24.736 2.724 ;
  LAYER M1 ;
        RECT 24.704 1.224 24.736 1.884 ;
  LAYER M1 ;
        RECT 22.784 2.064 22.816 2.724 ;
  LAYER M1 ;
        RECT 22.784 1.224 22.816 1.884 ;
  LAYER M1 ;
        RECT 24.064 2.064 24.096 2.724 ;
  LAYER M1 ;
        RECT 24.064 1.224 24.096 1.884 ;
  LAYER M1 ;
        RECT 25.344 2.064 25.376 2.724 ;
  LAYER M1 ;
        RECT 25.344 1.224 25.376 1.884 ;
  LAYER M1 ;
        RECT 22.064 2.064 22.096 2.724 ;
  LAYER M1 ;
        RECT 22.064 1.224 22.096 1.884 ;
  LAYER M1 ;
        RECT 23.344 2.064 23.376 2.724 ;
  LAYER M1 ;
        RECT 23.344 1.224 23.376 1.884 ;
  LAYER M1 ;
        RECT 24.624 2.064 24.656 2.724 ;
  LAYER M1 ;
        RECT 24.624 1.224 24.656 1.884 ;
  LAYER M1 ;
        RECT 22.704 2.064 22.736 2.724 ;
  LAYER M1 ;
        RECT 22.704 1.224 22.736 1.884 ;
  LAYER M1 ;
        RECT 23.984 2.064 24.016 2.724 ;
  LAYER M1 ;
        RECT 23.984 1.224 24.016 1.884 ;
  LAYER M1 ;
        RECT 25.264 2.064 25.296 2.724 ;
  LAYER M1 ;
        RECT 25.264 1.224 25.296 1.884 ;
  LAYER M1 ;
        RECT 22.224 2.064 22.256 2.724 ;
  LAYER M1 ;
        RECT 22.224 1.224 22.256 1.884 ;
  LAYER M1 ;
        RECT 23.504 2.064 23.536 2.724 ;
  LAYER M1 ;
        RECT 23.504 1.224 23.536 1.884 ;
  LAYER M1 ;
        RECT 24.784 2.064 24.816 2.724 ;
  LAYER M1 ;
        RECT 24.784 1.224 24.816 1.884 ;
  LAYER M1 ;
        RECT 22.864 2.064 22.896 2.724 ;
  LAYER M1 ;
        RECT 22.864 1.224 22.896 1.884 ;
  LAYER M1 ;
        RECT 24.144 2.064 24.176 2.724 ;
  LAYER M1 ;
        RECT 24.144 1.224 24.176 1.884 ;
  LAYER M1 ;
        RECT 25.424 2.064 25.456 2.724 ;
  LAYER M1 ;
        RECT 25.424 1.224 25.456 1.884 ;
  LAYER M2 ;
        RECT 22.044 2.672 25.316 2.704 ;
  LAYER M2 ;
        RECT 22.204 2.588 24.836 2.62 ;
  LAYER M2 ;
        RECT 22.844 2.504 25.476 2.536 ;
  LAYER M2 ;
        RECT 22.124 2.42 24.756 2.452 ;
  LAYER M2 ;
        RECT 22.764 2.336 25.396 2.368 ;
  LAYER M2 ;
        RECT 22.044 1.832 25.316 1.864 ;
  LAYER M2 ;
        RECT 22.844 1.748 25.476 1.78 ;
  LAYER M2 ;
        RECT 22.204 1.664 24.836 1.696 ;
  LAYER M2 ;
        RECT 22.764 1.58 25.396 1.612 ;
  LAYER M2 ;
        RECT 25.424 1.412 25.456 1.444 ;
  LAYER M1 ;
        RECT 24.064 0.216 24.096 0.876 ;
  LAYER M1 ;
        RECT 23.424 0.216 23.456 0.876 ;
  LAYER M1 ;
        RECT 25.984 0.216 26.016 0.876 ;
  LAYER M1 ;
        RECT 25.344 0.216 25.376 0.876 ;
  LAYER M1 ;
        RECT 24.704 0.216 24.736 0.876 ;
  LAYER M1 ;
        RECT 22.784 0.216 22.816 0.876 ;
  LAYER M1 ;
        RECT 22.144 0.216 22.176 0.876 ;
  LAYER M1 ;
        RECT 21.504 0.216 21.536 0.876 ;
  LAYER M1 ;
        RECT 24.144 0.216 24.176 0.876 ;
  LAYER M1 ;
        RECT 23.504 0.216 23.536 0.876 ;
  LAYER M1 ;
        RECT 26.064 0.216 26.096 0.876 ;
  LAYER M1 ;
        RECT 25.424 0.216 25.456 0.876 ;
  LAYER M1 ;
        RECT 24.784 0.216 24.816 0.876 ;
  LAYER M1 ;
        RECT 22.864 0.216 22.896 0.876 ;
  LAYER M1 ;
        RECT 22.224 0.216 22.256 0.876 ;
  LAYER M1 ;
        RECT 21.584 0.216 21.616 0.876 ;
  LAYER M1 ;
        RECT 23.984 0.216 24.016 0.876 ;
  LAYER M1 ;
        RECT 23.344 0.216 23.376 0.876 ;
  LAYER M1 ;
        RECT 25.904 0.216 25.936 0.876 ;
  LAYER M1 ;
        RECT 25.264 0.216 25.296 0.876 ;
  LAYER M1 ;
        RECT 24.624 0.216 24.656 0.876 ;
  LAYER M1 ;
        RECT 22.704 0.216 22.736 0.876 ;
  LAYER M1 ;
        RECT 22.064 0.216 22.096 0.876 ;
  LAYER M1 ;
        RECT 21.424 0.656 21.456 0.688 ;
  LAYER M1 ;
        RECT 22.784 3.912 22.816 4.572 ;
  LAYER M1 ;
        RECT 24.704 3.912 24.736 4.572 ;
  LAYER M1 ;
        RECT 23.424 3.912 23.456 4.572 ;
  LAYER M1 ;
        RECT 24.064 3.912 24.096 4.572 ;
  LAYER M1 ;
        RECT 22.704 3.912 22.736 4.572 ;
  LAYER M1 ;
        RECT 24.784 3.912 24.816 4.572 ;
  LAYER M1 ;
        RECT 23.344 3.912 23.376 4.572 ;
  LAYER M1 ;
        RECT 24.144 3.912 24.176 4.572 ;
  LAYER M1 ;
        RECT 22.864 3.912 22.896 4.572 ;
  LAYER M1 ;
        RECT 24.624 3.912 24.656 4.572 ;
  LAYER M1 ;
        RECT 23.504 3.912 23.536 4.572 ;
  LAYER M1 ;
        RECT 23.984 4.1 24.016 4.132 ;
  LAYER M1 ;
        RECT 25.344 2.904 25.376 3.564 ;
  LAYER M1 ;
        RECT 24.064 2.904 24.096 3.564 ;
  LAYER M1 ;
        RECT 22.784 2.904 22.816 3.564 ;
  LAYER M1 ;
        RECT 24.704 2.904 24.736 3.564 ;
  LAYER M1 ;
        RECT 23.424 2.904 23.456 3.564 ;
  LAYER M1 ;
        RECT 22.144 2.904 22.176 3.564 ;
  LAYER M1 ;
        RECT 25.424 2.904 25.456 3.564 ;
  LAYER M1 ;
        RECT 24.144 2.904 24.176 3.564 ;
  LAYER M1 ;
        RECT 22.864 2.904 22.896 3.564 ;
  LAYER M1 ;
        RECT 24.784 2.904 24.816 3.564 ;
  LAYER M1 ;
        RECT 23.504 2.904 23.536 3.564 ;
  LAYER M1 ;
        RECT 22.224 2.904 22.256 3.564 ;
  LAYER M1 ;
        RECT 25.264 2.904 25.296 3.564 ;
  LAYER M1 ;
        RECT 23.984 2.904 24.016 3.564 ;
  LAYER M1 ;
        RECT 22.704 2.904 22.736 3.564 ;
  LAYER M1 ;
        RECT 24.624 2.904 24.656 3.564 ;
  LAYER M1 ;
        RECT 23.344 2.904 23.376 3.564 ;
  LAYER M1 ;
        RECT 22.064 3.344 22.096 3.376 ;
  LAYER M1 ;
        RECT 6.416 14.244 6.448 14.316 ;
  LAYER M2 ;
        RECT 6.396 14.264 6.468 14.296 ;
  LAYER M1 ;
        RECT 9.392 14.244 9.424 14.316 ;
  LAYER M2 ;
        RECT 9.372 14.264 9.444 14.296 ;
  LAYER M2 ;
        RECT 6.432 14.264 9.408 14.296 ;
  LAYER M2 ;
        RECT 6.124 0.908 6.836 0.94 ;
  LAYER M1 ;
        RECT 9.312 31.044 9.344 31.116 ;
  LAYER M2 ;
        RECT 9.292 31.064 9.364 31.096 ;
  LAYER M1 ;
        RECT 6.336 31.044 6.368 31.116 ;
  LAYER M2 ;
        RECT 6.316 31.064 6.388 31.096 ;
  LAYER M2 ;
        RECT 6.352 31.064 9.328 31.096 ;
  LAYER M2 ;
        RECT 6.544 14.264 6.576 14.296 ;
  LAYER M3 ;
        RECT 6.54 0.924 6.58 14.28 ;
  LAYER M2 ;
        RECT 6.544 0.908 6.576 0.94 ;
  LAYER M2 ;
        RECT 8.864 14.264 8.896 14.296 ;
  LAYER M3 ;
        RECT 8.86 14.28 8.9 17.808 ;
  LAYER M4 ;
        RECT 8.86 17.788 8.9 17.828 ;
  LAYER M5 ;
        RECT 8.848 17.808 8.912 31.08 ;
  LAYER M4 ;
        RECT 8.86 31.06 8.9 31.1 ;
  LAYER M3 ;
        RECT 8.86 31.06 8.9 31.1 ;
  LAYER M2 ;
        RECT 8.864 31.064 8.896 31.096 ;
  LAYER M1 ;
        RECT 6.256 1.308 6.288 1.38 ;
  LAYER M2 ;
        RECT 6.236 1.328 6.308 1.36 ;
  LAYER M1 ;
        RECT 9.232 1.308 9.264 1.38 ;
  LAYER M2 ;
        RECT 9.212 1.328 9.284 1.36 ;
  LAYER M2 ;
        RECT 6.272 1.328 9.248 1.36 ;
  LAYER M2 ;
        RECT 5.404 0.32 5.476 0.352 ;
  LAYER M2 ;
        RECT 15.564 0.32 15.636 0.352 ;
  LAYER M2 ;
        RECT 5.76 1.328 6.24 1.36 ;
  LAYER M3 ;
        RECT 5.74 0.336 5.78 1.344 ;
  LAYER M4 ;
        RECT 5.44 0.316 5.76 0.356 ;
  LAYER M3 ;
        RECT 5.42 0.316 5.46 0.356 ;
  LAYER M2 ;
        RECT 5.424 0.32 5.456 0.352 ;
  LAYER M2 ;
        RECT 9.28 1.328 15.28 1.36 ;
  LAYER M3 ;
        RECT 15.26 0.336 15.3 1.344 ;
  LAYER M4 ;
        RECT 15.28 0.316 15.6 0.356 ;
  LAYER M3 ;
        RECT 15.58 0.316 15.62 0.356 ;
  LAYER M2 ;
        RECT 15.584 0.32 15.616 0.352 ;
  LAYER M2 ;
        RECT 7.484 0.908 8.196 0.94 ;
  LAYER M1 ;
        RECT 9.152 15 9.184 15.072 ;
  LAYER M2 ;
        RECT 9.132 15.02 9.204 15.052 ;
  LAYER M1 ;
        RECT 6.176 15 6.208 15.072 ;
  LAYER M2 ;
        RECT 6.156 15.02 6.228 15.052 ;
  LAYER M2 ;
        RECT 6.192 15.02 9.168 15.052 ;
  LAYER M2 ;
        RECT 7.504 0.908 7.536 0.94 ;
  LAYER M3 ;
        RECT 7.5 0.924 7.54 15.036 ;
  LAYER M2 ;
        RECT 7.504 15.02 7.536 15.052 ;
  LAYER M1 ;
        RECT 9.008 5.004 9.04 5.076 ;
  LAYER M2 ;
        RECT 8.988 5.024 9.06 5.056 ;
  LAYER M2 ;
        RECT 6.272 5.024 9.024 5.056 ;
  LAYER M1 ;
        RECT 6.256 5.004 6.288 5.076 ;
  LAYER M2 ;
        RECT 6.236 5.024 6.308 5.056 ;
  LAYER M1 ;
        RECT 9.008 8.112 9.04 8.184 ;
  LAYER M2 ;
        RECT 8.988 8.132 9.06 8.164 ;
  LAYER M2 ;
        RECT 6.272 8.132 9.024 8.164 ;
  LAYER M1 ;
        RECT 6.256 8.112 6.288 8.184 ;
  LAYER M2 ;
        RECT 6.236 8.132 6.308 8.164 ;
  LAYER M1 ;
        RECT 6.032 5.004 6.064 5.076 ;
  LAYER M2 ;
        RECT 6.012 5.024 6.084 5.056 ;
  LAYER M1 ;
        RECT 6.032 4.872 6.064 5.04 ;
  LAYER M1 ;
        RECT 6.032 4.836 6.064 4.908 ;
  LAYER M2 ;
        RECT 6.012 4.856 6.084 4.888 ;
  LAYER M2 ;
        RECT 6.048 4.856 6.272 4.888 ;
  LAYER M1 ;
        RECT 6.256 4.836 6.288 4.908 ;
  LAYER M2 ;
        RECT 6.236 4.856 6.308 4.888 ;
  LAYER M1 ;
        RECT 6.032 8.112 6.064 8.184 ;
  LAYER M2 ;
        RECT 6.012 8.132 6.084 8.164 ;
  LAYER M1 ;
        RECT 6.032 7.98 6.064 8.148 ;
  LAYER M1 ;
        RECT 6.032 7.944 6.064 8.016 ;
  LAYER M2 ;
        RECT 6.012 7.964 6.084 7.996 ;
  LAYER M2 ;
        RECT 6.048 7.964 6.272 7.996 ;
  LAYER M1 ;
        RECT 6.256 7.944 6.288 8.016 ;
  LAYER M2 ;
        RECT 6.236 7.964 6.308 7.996 ;
  LAYER M1 ;
        RECT 6.256 1.308 6.288 1.38 ;
  LAYER M2 ;
        RECT 6.236 1.328 6.308 1.36 ;
  LAYER M1 ;
        RECT 6.256 1.344 6.288 1.596 ;
  LAYER M1 ;
        RECT 6.256 1.596 6.288 8.148 ;
  LAYER M1 ;
        RECT 11.984 8.112 12.016 8.184 ;
  LAYER M2 ;
        RECT 11.964 8.132 12.036 8.164 ;
  LAYER M2 ;
        RECT 9.248 8.132 12 8.164 ;
  LAYER M1 ;
        RECT 9.232 8.112 9.264 8.184 ;
  LAYER M2 ;
        RECT 9.212 8.132 9.284 8.164 ;
  LAYER M1 ;
        RECT 11.984 5.004 12.016 5.076 ;
  LAYER M2 ;
        RECT 11.964 5.024 12.036 5.056 ;
  LAYER M2 ;
        RECT 9.248 5.024 12 5.056 ;
  LAYER M1 ;
        RECT 9.232 5.004 9.264 5.076 ;
  LAYER M2 ;
        RECT 9.212 5.024 9.284 5.056 ;
  LAYER M1 ;
        RECT 9.232 1.308 9.264 1.38 ;
  LAYER M2 ;
        RECT 9.212 1.328 9.284 1.36 ;
  LAYER M1 ;
        RECT 9.232 1.344 9.264 1.596 ;
  LAYER M1 ;
        RECT 9.232 1.596 9.264 8.148 ;
  LAYER M2 ;
        RECT 6.272 1.328 9.248 1.36 ;
  LAYER M1 ;
        RECT 3.056 1.896 3.088 1.968 ;
  LAYER M2 ;
        RECT 3.036 1.916 3.108 1.948 ;
  LAYER M1 ;
        RECT 3.056 1.764 3.088 1.932 ;
  LAYER M1 ;
        RECT 3.056 1.728 3.088 1.8 ;
  LAYER M2 ;
        RECT 3.036 1.748 3.108 1.78 ;
  LAYER M2 ;
        RECT 3.072 1.748 3.296 1.78 ;
  LAYER M1 ;
        RECT 3.28 1.728 3.312 1.8 ;
  LAYER M2 ;
        RECT 3.26 1.748 3.332 1.78 ;
  LAYER M1 ;
        RECT 3.056 5.004 3.088 5.076 ;
  LAYER M2 ;
        RECT 3.036 5.024 3.108 5.056 ;
  LAYER M1 ;
        RECT 3.056 4.872 3.088 5.04 ;
  LAYER M1 ;
        RECT 3.056 4.836 3.088 4.908 ;
  LAYER M2 ;
        RECT 3.036 4.856 3.108 4.888 ;
  LAYER M2 ;
        RECT 3.072 4.856 3.296 4.888 ;
  LAYER M1 ;
        RECT 3.28 4.836 3.312 4.908 ;
  LAYER M2 ;
        RECT 3.26 4.856 3.332 4.888 ;
  LAYER M1 ;
        RECT 3.056 8.112 3.088 8.184 ;
  LAYER M2 ;
        RECT 3.036 8.132 3.108 8.164 ;
  LAYER M1 ;
        RECT 3.056 7.98 3.088 8.148 ;
  LAYER M1 ;
        RECT 3.056 7.944 3.088 8.016 ;
  LAYER M2 ;
        RECT 3.036 7.964 3.108 7.996 ;
  LAYER M2 ;
        RECT 3.072 7.964 3.296 7.996 ;
  LAYER M1 ;
        RECT 3.28 7.944 3.312 8.016 ;
  LAYER M2 ;
        RECT 3.26 7.964 3.332 7.996 ;
  LAYER M1 ;
        RECT 3.056 11.22 3.088 11.292 ;
  LAYER M2 ;
        RECT 3.036 11.24 3.108 11.272 ;
  LAYER M1 ;
        RECT 3.056 11.088 3.088 11.256 ;
  LAYER M1 ;
        RECT 3.056 11.052 3.088 11.124 ;
  LAYER M2 ;
        RECT 3.036 11.072 3.108 11.104 ;
  LAYER M2 ;
        RECT 3.072 11.072 3.296 11.104 ;
  LAYER M1 ;
        RECT 3.28 11.052 3.312 11.124 ;
  LAYER M2 ;
        RECT 3.26 11.072 3.332 11.104 ;
  LAYER M1 ;
        RECT 6.032 1.896 6.064 1.968 ;
  LAYER M2 ;
        RECT 6.012 1.916 6.084 1.948 ;
  LAYER M2 ;
        RECT 3.296 1.916 6.048 1.948 ;
  LAYER M1 ;
        RECT 3.28 1.896 3.312 1.968 ;
  LAYER M2 ;
        RECT 3.26 1.916 3.332 1.948 ;
  LAYER M1 ;
        RECT 6.032 11.22 6.064 11.292 ;
  LAYER M2 ;
        RECT 6.012 11.24 6.084 11.272 ;
  LAYER M2 ;
        RECT 3.296 11.24 6.048 11.272 ;
  LAYER M1 ;
        RECT 3.28 11.22 3.312 11.292 ;
  LAYER M2 ;
        RECT 3.26 11.24 3.332 11.272 ;
  LAYER M1 ;
        RECT 3.28 1.14 3.312 1.212 ;
  LAYER M2 ;
        RECT 3.26 1.16 3.332 1.192 ;
  LAYER M1 ;
        RECT 3.28 1.176 3.312 1.596 ;
  LAYER M1 ;
        RECT 3.28 1.596 3.312 11.256 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 1.968 ;
  LAYER M2 ;
        RECT 11.964 1.916 12.036 1.948 ;
  LAYER M1 ;
        RECT 11.984 1.764 12.016 1.932 ;
  LAYER M1 ;
        RECT 11.984 1.728 12.016 1.8 ;
  LAYER M2 ;
        RECT 11.964 1.748 12.036 1.78 ;
  LAYER M2 ;
        RECT 12 1.748 12.224 1.78 ;
  LAYER M1 ;
        RECT 12.208 1.728 12.24 1.8 ;
  LAYER M2 ;
        RECT 12.188 1.748 12.26 1.78 ;
  LAYER M1 ;
        RECT 11.984 11.22 12.016 11.292 ;
  LAYER M2 ;
        RECT 11.964 11.24 12.036 11.272 ;
  LAYER M1 ;
        RECT 11.984 11.088 12.016 11.256 ;
  LAYER M1 ;
        RECT 11.984 11.052 12.016 11.124 ;
  LAYER M2 ;
        RECT 11.964 11.072 12.036 11.104 ;
  LAYER M2 ;
        RECT 12 11.072 12.224 11.104 ;
  LAYER M1 ;
        RECT 12.208 11.052 12.24 11.124 ;
  LAYER M2 ;
        RECT 12.188 11.072 12.26 11.104 ;
  LAYER M1 ;
        RECT 14.96 1.896 14.992 1.968 ;
  LAYER M2 ;
        RECT 14.94 1.916 15.012 1.948 ;
  LAYER M2 ;
        RECT 12.224 1.916 14.976 1.948 ;
  LAYER M1 ;
        RECT 12.208 1.896 12.24 1.968 ;
  LAYER M2 ;
        RECT 12.188 1.916 12.26 1.948 ;
  LAYER M1 ;
        RECT 14.96 5.004 14.992 5.076 ;
  LAYER M2 ;
        RECT 14.94 5.024 15.012 5.056 ;
  LAYER M2 ;
        RECT 12.224 5.024 14.976 5.056 ;
  LAYER M1 ;
        RECT 12.208 5.004 12.24 5.076 ;
  LAYER M2 ;
        RECT 12.188 5.024 12.26 5.056 ;
  LAYER M1 ;
        RECT 14.96 8.112 14.992 8.184 ;
  LAYER M2 ;
        RECT 14.94 8.132 15.012 8.164 ;
  LAYER M2 ;
        RECT 12.224 8.132 14.976 8.164 ;
  LAYER M1 ;
        RECT 12.208 8.112 12.24 8.184 ;
  LAYER M2 ;
        RECT 12.188 8.132 12.26 8.164 ;
  LAYER M1 ;
        RECT 14.96 11.22 14.992 11.292 ;
  LAYER M2 ;
        RECT 14.94 11.24 15.012 11.272 ;
  LAYER M2 ;
        RECT 12.224 11.24 14.976 11.272 ;
  LAYER M1 ;
        RECT 12.208 11.22 12.24 11.292 ;
  LAYER M2 ;
        RECT 12.188 11.24 12.26 11.272 ;
  LAYER M1 ;
        RECT 12.208 1.14 12.24 1.212 ;
  LAYER M2 ;
        RECT 12.188 1.16 12.26 1.192 ;
  LAYER M1 ;
        RECT 12.208 1.176 12.24 1.596 ;
  LAYER M1 ;
        RECT 12.208 1.596 12.24 11.256 ;
  LAYER M2 ;
        RECT 3.296 1.16 12.224 1.192 ;
  LAYER M1 ;
        RECT 9.008 11.22 9.04 11.292 ;
  LAYER M2 ;
        RECT 8.988 11.24 9.06 11.272 ;
  LAYER M2 ;
        RECT 6.048 11.24 9.024 11.272 ;
  LAYER M1 ;
        RECT 6.032 11.22 6.064 11.292 ;
  LAYER M2 ;
        RECT 6.012 11.24 6.084 11.272 ;
  LAYER M1 ;
        RECT 9.008 1.896 9.04 1.968 ;
  LAYER M2 ;
        RECT 8.988 1.916 9.06 1.948 ;
  LAYER M2 ;
        RECT 9.024 1.916 12 1.948 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 1.968 ;
  LAYER M2 ;
        RECT 11.964 1.916 12.036 1.948 ;
  LAYER M1 ;
        RECT 6.64 7.44 6.672 7.512 ;
  LAYER M2 ;
        RECT 6.62 7.46 6.692 7.492 ;
  LAYER M2 ;
        RECT 6.432 7.46 6.656 7.492 ;
  LAYER M1 ;
        RECT 6.416 7.44 6.448 7.512 ;
  LAYER M2 ;
        RECT 6.396 7.46 6.468 7.492 ;
  LAYER M1 ;
        RECT 6.64 10.548 6.672 10.62 ;
  LAYER M2 ;
        RECT 6.62 10.568 6.692 10.6 ;
  LAYER M2 ;
        RECT 6.432 10.568 6.656 10.6 ;
  LAYER M1 ;
        RECT 6.416 10.548 6.448 10.62 ;
  LAYER M2 ;
        RECT 6.396 10.568 6.468 10.6 ;
  LAYER M1 ;
        RECT 3.664 7.44 3.696 7.512 ;
  LAYER M2 ;
        RECT 3.644 7.46 3.716 7.492 ;
  LAYER M1 ;
        RECT 3.664 7.476 3.696 7.644 ;
  LAYER M1 ;
        RECT 3.664 7.608 3.696 7.68 ;
  LAYER M2 ;
        RECT 3.644 7.628 3.716 7.66 ;
  LAYER M2 ;
        RECT 3.68 7.628 6.432 7.66 ;
  LAYER M1 ;
        RECT 6.416 7.608 6.448 7.68 ;
  LAYER M2 ;
        RECT 6.396 7.628 6.468 7.66 ;
  LAYER M1 ;
        RECT 3.664 10.548 3.696 10.62 ;
  LAYER M2 ;
        RECT 3.644 10.568 3.716 10.6 ;
  LAYER M1 ;
        RECT 3.664 10.584 3.696 10.752 ;
  LAYER M1 ;
        RECT 3.664 10.716 3.696 10.788 ;
  LAYER M2 ;
        RECT 3.644 10.736 3.716 10.768 ;
  LAYER M2 ;
        RECT 3.68 10.736 6.432 10.768 ;
  LAYER M1 ;
        RECT 6.416 10.716 6.448 10.788 ;
  LAYER M2 ;
        RECT 6.396 10.736 6.468 10.768 ;
  LAYER M1 ;
        RECT 6.416 14.244 6.448 14.316 ;
  LAYER M2 ;
        RECT 6.396 14.264 6.468 14.296 ;
  LAYER M1 ;
        RECT 6.416 14.028 6.448 14.28 ;
  LAYER M1 ;
        RECT 6.416 7.476 6.448 14.028 ;
  LAYER M1 ;
        RECT 9.616 10.548 9.648 10.62 ;
  LAYER M2 ;
        RECT 9.596 10.568 9.668 10.6 ;
  LAYER M2 ;
        RECT 9.408 10.568 9.632 10.6 ;
  LAYER M1 ;
        RECT 9.392 10.548 9.424 10.62 ;
  LAYER M2 ;
        RECT 9.372 10.568 9.444 10.6 ;
  LAYER M1 ;
        RECT 9.616 7.44 9.648 7.512 ;
  LAYER M2 ;
        RECT 9.596 7.46 9.668 7.492 ;
  LAYER M2 ;
        RECT 9.408 7.46 9.632 7.492 ;
  LAYER M1 ;
        RECT 9.392 7.44 9.424 7.512 ;
  LAYER M2 ;
        RECT 9.372 7.46 9.444 7.492 ;
  LAYER M1 ;
        RECT 9.392 14.244 9.424 14.316 ;
  LAYER M2 ;
        RECT 9.372 14.264 9.444 14.296 ;
  LAYER M1 ;
        RECT 9.392 14.028 9.424 14.28 ;
  LAYER M1 ;
        RECT 9.392 7.476 9.424 14.028 ;
  LAYER M2 ;
        RECT 6.432 14.264 9.408 14.296 ;
  LAYER M1 ;
        RECT 0.688 4.332 0.72 4.404 ;
  LAYER M2 ;
        RECT 0.668 4.352 0.74 4.384 ;
  LAYER M2 ;
        RECT 0.32 4.352 0.704 4.384 ;
  LAYER M1 ;
        RECT 0.304 4.332 0.336 4.404 ;
  LAYER M2 ;
        RECT 0.284 4.352 0.356 4.384 ;
  LAYER M1 ;
        RECT 0.688 7.44 0.72 7.512 ;
  LAYER M2 ;
        RECT 0.668 7.46 0.74 7.492 ;
  LAYER M2 ;
        RECT 0.32 7.46 0.704 7.492 ;
  LAYER M1 ;
        RECT 0.304 7.44 0.336 7.512 ;
  LAYER M2 ;
        RECT 0.284 7.46 0.356 7.492 ;
  LAYER M1 ;
        RECT 0.688 10.548 0.72 10.62 ;
  LAYER M2 ;
        RECT 0.668 10.568 0.74 10.6 ;
  LAYER M2 ;
        RECT 0.32 10.568 0.704 10.6 ;
  LAYER M1 ;
        RECT 0.304 10.548 0.336 10.62 ;
  LAYER M2 ;
        RECT 0.284 10.568 0.356 10.6 ;
  LAYER M1 ;
        RECT 0.688 13.656 0.72 13.728 ;
  LAYER M2 ;
        RECT 0.668 13.676 0.74 13.708 ;
  LAYER M2 ;
        RECT 0.32 13.676 0.704 13.708 ;
  LAYER M1 ;
        RECT 0.304 13.656 0.336 13.728 ;
  LAYER M2 ;
        RECT 0.284 13.676 0.356 13.708 ;
  LAYER M1 ;
        RECT 0.304 14.412 0.336 14.484 ;
  LAYER M2 ;
        RECT 0.284 14.432 0.356 14.464 ;
  LAYER M1 ;
        RECT 0.304 14.028 0.336 14.448 ;
  LAYER M1 ;
        RECT 0.304 4.368 0.336 14.028 ;
  LAYER M1 ;
        RECT 12.592 4.332 12.624 4.404 ;
  LAYER M2 ;
        RECT 12.572 4.352 12.644 4.384 ;
  LAYER M1 ;
        RECT 12.592 4.368 12.624 4.536 ;
  LAYER M1 ;
        RECT 12.592 4.5 12.624 4.572 ;
  LAYER M2 ;
        RECT 12.572 4.52 12.644 4.552 ;
  LAYER M2 ;
        RECT 12.608 4.52 15.2 4.552 ;
  LAYER M1 ;
        RECT 15.184 4.5 15.216 4.572 ;
  LAYER M2 ;
        RECT 15.164 4.52 15.236 4.552 ;
  LAYER M1 ;
        RECT 12.592 7.44 12.624 7.512 ;
  LAYER M2 ;
        RECT 12.572 7.46 12.644 7.492 ;
  LAYER M1 ;
        RECT 12.592 7.476 12.624 7.644 ;
  LAYER M1 ;
        RECT 12.592 7.608 12.624 7.68 ;
  LAYER M2 ;
        RECT 12.572 7.628 12.644 7.66 ;
  LAYER M2 ;
        RECT 12.608 7.628 15.2 7.66 ;
  LAYER M1 ;
        RECT 15.184 7.608 15.216 7.68 ;
  LAYER M2 ;
        RECT 15.164 7.628 15.236 7.66 ;
  LAYER M1 ;
        RECT 12.592 10.548 12.624 10.62 ;
  LAYER M2 ;
        RECT 12.572 10.568 12.644 10.6 ;
  LAYER M1 ;
        RECT 12.592 10.584 12.624 10.752 ;
  LAYER M1 ;
        RECT 12.592 10.716 12.624 10.788 ;
  LAYER M2 ;
        RECT 12.572 10.736 12.644 10.768 ;
  LAYER M2 ;
        RECT 12.608 10.736 15.2 10.768 ;
  LAYER M1 ;
        RECT 15.184 10.716 15.216 10.788 ;
  LAYER M2 ;
        RECT 15.164 10.736 15.236 10.768 ;
  LAYER M1 ;
        RECT 12.592 13.656 12.624 13.728 ;
  LAYER M2 ;
        RECT 12.572 13.676 12.644 13.708 ;
  LAYER M1 ;
        RECT 12.592 13.692 12.624 13.86 ;
  LAYER M1 ;
        RECT 12.592 13.824 12.624 13.896 ;
  LAYER M2 ;
        RECT 12.572 13.844 12.644 13.876 ;
  LAYER M2 ;
        RECT 12.608 13.844 15.2 13.876 ;
  LAYER M1 ;
        RECT 15.184 13.824 15.216 13.896 ;
  LAYER M2 ;
        RECT 15.164 13.844 15.236 13.876 ;
  LAYER M1 ;
        RECT 15.184 14.412 15.216 14.484 ;
  LAYER M2 ;
        RECT 15.164 14.432 15.236 14.464 ;
  LAYER M1 ;
        RECT 15.184 14.028 15.216 14.448 ;
  LAYER M1 ;
        RECT 15.184 4.536 15.216 14.028 ;
  LAYER M2 ;
        RECT 0.32 14.432 15.2 14.464 ;
  LAYER M1 ;
        RECT 3.664 4.332 3.696 4.404 ;
  LAYER M2 ;
        RECT 3.644 4.352 3.716 4.384 ;
  LAYER M2 ;
        RECT 0.704 4.352 3.68 4.384 ;
  LAYER M1 ;
        RECT 0.688 4.332 0.72 4.404 ;
  LAYER M2 ;
        RECT 0.668 4.352 0.74 4.384 ;
  LAYER M1 ;
        RECT 3.664 13.656 3.696 13.728 ;
  LAYER M2 ;
        RECT 3.644 13.676 3.716 13.708 ;
  LAYER M2 ;
        RECT 0.704 13.676 3.68 13.708 ;
  LAYER M1 ;
        RECT 0.688 13.656 0.72 13.728 ;
  LAYER M2 ;
        RECT 0.668 13.676 0.74 13.708 ;
  LAYER M1 ;
        RECT 6.64 13.656 6.672 13.728 ;
  LAYER M2 ;
        RECT 6.62 13.676 6.692 13.708 ;
  LAYER M2 ;
        RECT 3.68 13.676 6.656 13.708 ;
  LAYER M1 ;
        RECT 3.664 13.656 3.696 13.728 ;
  LAYER M2 ;
        RECT 3.644 13.676 3.716 13.708 ;
  LAYER M1 ;
        RECT 9.616 13.656 9.648 13.728 ;
  LAYER M2 ;
        RECT 9.596 13.676 9.668 13.708 ;
  LAYER M2 ;
        RECT 6.656 13.676 9.632 13.708 ;
  LAYER M1 ;
        RECT 6.64 13.656 6.672 13.728 ;
  LAYER M2 ;
        RECT 6.62 13.676 6.692 13.708 ;
  LAYER M1 ;
        RECT 9.616 4.332 9.648 4.404 ;
  LAYER M2 ;
        RECT 9.596 4.352 9.668 4.384 ;
  LAYER M2 ;
        RECT 9.632 4.352 12.608 4.384 ;
  LAYER M1 ;
        RECT 12.592 4.332 12.624 4.404 ;
  LAYER M2 ;
        RECT 12.572 4.352 12.644 4.384 ;
  LAYER M1 ;
        RECT 6.64 4.332 6.672 4.404 ;
  LAYER M2 ;
        RECT 6.62 4.352 6.692 4.384 ;
  LAYER M2 ;
        RECT 6.656 4.352 9.632 4.384 ;
  LAYER M1 ;
        RECT 9.616 4.332 9.648 4.404 ;
  LAYER M2 ;
        RECT 9.596 4.352 9.668 4.384 ;
  LAYER M1 ;
        RECT 0.688 1.896 0.72 4.404 ;
  LAYER M3 ;
        RECT 0.688 4.352 0.72 4.384 ;
  LAYER M1 ;
        RECT 0.752 1.896 0.784 4.404 ;
  LAYER M3 ;
        RECT 0.752 1.916 0.784 1.948 ;
  LAYER M1 ;
        RECT 0.816 1.896 0.848 4.404 ;
  LAYER M3 ;
        RECT 0.816 4.352 0.848 4.384 ;
  LAYER M1 ;
        RECT 0.88 1.896 0.912 4.404 ;
  LAYER M3 ;
        RECT 0.88 1.916 0.912 1.948 ;
  LAYER M1 ;
        RECT 0.944 1.896 0.976 4.404 ;
  LAYER M3 ;
        RECT 0.944 4.352 0.976 4.384 ;
  LAYER M1 ;
        RECT 1.008 1.896 1.04 4.404 ;
  LAYER M3 ;
        RECT 1.008 1.916 1.04 1.948 ;
  LAYER M1 ;
        RECT 1.072 1.896 1.104 4.404 ;
  LAYER M3 ;
        RECT 1.072 4.352 1.104 4.384 ;
  LAYER M1 ;
        RECT 1.136 1.896 1.168 4.404 ;
  LAYER M3 ;
        RECT 1.136 1.916 1.168 1.948 ;
  LAYER M1 ;
        RECT 1.2 1.896 1.232 4.404 ;
  LAYER M3 ;
        RECT 1.2 4.352 1.232 4.384 ;
  LAYER M1 ;
        RECT 1.264 1.896 1.296 4.404 ;
  LAYER M3 ;
        RECT 1.264 1.916 1.296 1.948 ;
  LAYER M1 ;
        RECT 1.328 1.896 1.36 4.404 ;
  LAYER M3 ;
        RECT 1.328 4.352 1.36 4.384 ;
  LAYER M1 ;
        RECT 1.392 1.896 1.424 4.404 ;
  LAYER M3 ;
        RECT 1.392 1.916 1.424 1.948 ;
  LAYER M1 ;
        RECT 1.456 1.896 1.488 4.404 ;
  LAYER M3 ;
        RECT 1.456 4.352 1.488 4.384 ;
  LAYER M1 ;
        RECT 1.52 1.896 1.552 4.404 ;
  LAYER M3 ;
        RECT 1.52 1.916 1.552 1.948 ;
  LAYER M1 ;
        RECT 1.584 1.896 1.616 4.404 ;
  LAYER M3 ;
        RECT 1.584 4.352 1.616 4.384 ;
  LAYER M1 ;
        RECT 1.648 1.896 1.68 4.404 ;
  LAYER M3 ;
        RECT 1.648 1.916 1.68 1.948 ;
  LAYER M1 ;
        RECT 1.712 1.896 1.744 4.404 ;
  LAYER M3 ;
        RECT 1.712 4.352 1.744 4.384 ;
  LAYER M1 ;
        RECT 1.776 1.896 1.808 4.404 ;
  LAYER M3 ;
        RECT 1.776 1.916 1.808 1.948 ;
  LAYER M1 ;
        RECT 1.84 1.896 1.872 4.404 ;
  LAYER M3 ;
        RECT 1.84 4.352 1.872 4.384 ;
  LAYER M1 ;
        RECT 1.904 1.896 1.936 4.404 ;
  LAYER M3 ;
        RECT 1.904 1.916 1.936 1.948 ;
  LAYER M1 ;
        RECT 1.968 1.896 2 4.404 ;
  LAYER M3 ;
        RECT 1.968 4.352 2 4.384 ;
  LAYER M1 ;
        RECT 2.032 1.896 2.064 4.404 ;
  LAYER M3 ;
        RECT 2.032 1.916 2.064 1.948 ;
  LAYER M1 ;
        RECT 2.096 1.896 2.128 4.404 ;
  LAYER M3 ;
        RECT 2.096 4.352 2.128 4.384 ;
  LAYER M1 ;
        RECT 2.16 1.896 2.192 4.404 ;
  LAYER M3 ;
        RECT 2.16 1.916 2.192 1.948 ;
  LAYER M1 ;
        RECT 2.224 1.896 2.256 4.404 ;
  LAYER M3 ;
        RECT 2.224 4.352 2.256 4.384 ;
  LAYER M1 ;
        RECT 2.288 1.896 2.32 4.404 ;
  LAYER M3 ;
        RECT 2.288 1.916 2.32 1.948 ;
  LAYER M1 ;
        RECT 2.352 1.896 2.384 4.404 ;
  LAYER M3 ;
        RECT 2.352 4.352 2.384 4.384 ;
  LAYER M1 ;
        RECT 2.416 1.896 2.448 4.404 ;
  LAYER M3 ;
        RECT 2.416 1.916 2.448 1.948 ;
  LAYER M1 ;
        RECT 2.48 1.896 2.512 4.404 ;
  LAYER M3 ;
        RECT 2.48 4.352 2.512 4.384 ;
  LAYER M1 ;
        RECT 2.544 1.896 2.576 4.404 ;
  LAYER M3 ;
        RECT 2.544 1.916 2.576 1.948 ;
  LAYER M1 ;
        RECT 2.608 1.896 2.64 4.404 ;
  LAYER M3 ;
        RECT 2.608 4.352 2.64 4.384 ;
  LAYER M1 ;
        RECT 2.672 1.896 2.704 4.404 ;
  LAYER M3 ;
        RECT 2.672 1.916 2.704 1.948 ;
  LAYER M1 ;
        RECT 2.736 1.896 2.768 4.404 ;
  LAYER M3 ;
        RECT 2.736 4.352 2.768 4.384 ;
  LAYER M1 ;
        RECT 2.8 1.896 2.832 4.404 ;
  LAYER M3 ;
        RECT 2.8 1.916 2.832 1.948 ;
  LAYER M1 ;
        RECT 2.864 1.896 2.896 4.404 ;
  LAYER M3 ;
        RECT 2.864 4.352 2.896 4.384 ;
  LAYER M1 ;
        RECT 2.928 1.896 2.96 4.404 ;
  LAYER M3 ;
        RECT 2.928 1.916 2.96 1.948 ;
  LAYER M1 ;
        RECT 2.992 1.896 3.024 4.404 ;
  LAYER M3 ;
        RECT 2.992 4.352 3.024 4.384 ;
  LAYER M1 ;
        RECT 3.056 1.896 3.088 4.404 ;
  LAYER M3 ;
        RECT 0.688 1.98 0.72 2.012 ;
  LAYER M2 ;
        RECT 3.056 2.044 3.088 2.076 ;
  LAYER M2 ;
        RECT 0.688 2.108 0.72 2.14 ;
  LAYER M2 ;
        RECT 3.056 2.172 3.088 2.204 ;
  LAYER M2 ;
        RECT 0.688 2.236 0.72 2.268 ;
  LAYER M2 ;
        RECT 3.056 2.3 3.088 2.332 ;
  LAYER M2 ;
        RECT 0.688 2.364 0.72 2.396 ;
  LAYER M2 ;
        RECT 3.056 2.428 3.088 2.46 ;
  LAYER M2 ;
        RECT 0.688 2.492 0.72 2.524 ;
  LAYER M2 ;
        RECT 3.056 2.556 3.088 2.588 ;
  LAYER M2 ;
        RECT 0.688 2.62 0.72 2.652 ;
  LAYER M2 ;
        RECT 3.056 2.684 3.088 2.716 ;
  LAYER M2 ;
        RECT 0.688 2.748 0.72 2.78 ;
  LAYER M2 ;
        RECT 3.056 2.812 3.088 2.844 ;
  LAYER M2 ;
        RECT 0.688 2.876 0.72 2.908 ;
  LAYER M2 ;
        RECT 3.056 2.94 3.088 2.972 ;
  LAYER M2 ;
        RECT 0.688 3.004 0.72 3.036 ;
  LAYER M2 ;
        RECT 3.056 3.068 3.088 3.1 ;
  LAYER M2 ;
        RECT 0.688 3.132 0.72 3.164 ;
  LAYER M2 ;
        RECT 3.056 3.196 3.088 3.228 ;
  LAYER M2 ;
        RECT 0.688 3.26 0.72 3.292 ;
  LAYER M2 ;
        RECT 3.056 3.324 3.088 3.356 ;
  LAYER M2 ;
        RECT 0.688 3.388 0.72 3.42 ;
  LAYER M2 ;
        RECT 3.056 3.452 3.088 3.484 ;
  LAYER M2 ;
        RECT 0.688 3.516 0.72 3.548 ;
  LAYER M2 ;
        RECT 3.056 3.58 3.088 3.612 ;
  LAYER M2 ;
        RECT 0.688 3.644 0.72 3.676 ;
  LAYER M2 ;
        RECT 3.056 3.708 3.088 3.74 ;
  LAYER M2 ;
        RECT 0.688 3.772 0.72 3.804 ;
  LAYER M2 ;
        RECT 3.056 3.836 3.088 3.868 ;
  LAYER M2 ;
        RECT 0.688 3.9 0.72 3.932 ;
  LAYER M2 ;
        RECT 3.056 3.964 3.088 3.996 ;
  LAYER M2 ;
        RECT 0.688 4.028 0.72 4.06 ;
  LAYER M2 ;
        RECT 3.056 4.092 3.088 4.124 ;
  LAYER M2 ;
        RECT 0.688 4.156 0.72 4.188 ;
  LAYER M2 ;
        RECT 3.056 4.22 3.088 4.252 ;
  LAYER M2 ;
        RECT 0.64 1.848 3.136 4.452 ;
  LAYER M1 ;
        RECT 0.688 5.004 0.72 7.512 ;
  LAYER M3 ;
        RECT 0.688 7.46 0.72 7.492 ;
  LAYER M1 ;
        RECT 0.752 5.004 0.784 7.512 ;
  LAYER M3 ;
        RECT 0.752 5.024 0.784 5.056 ;
  LAYER M1 ;
        RECT 0.816 5.004 0.848 7.512 ;
  LAYER M3 ;
        RECT 0.816 7.46 0.848 7.492 ;
  LAYER M1 ;
        RECT 0.88 5.004 0.912 7.512 ;
  LAYER M3 ;
        RECT 0.88 5.024 0.912 5.056 ;
  LAYER M1 ;
        RECT 0.944 5.004 0.976 7.512 ;
  LAYER M3 ;
        RECT 0.944 7.46 0.976 7.492 ;
  LAYER M1 ;
        RECT 1.008 5.004 1.04 7.512 ;
  LAYER M3 ;
        RECT 1.008 5.024 1.04 5.056 ;
  LAYER M1 ;
        RECT 1.072 5.004 1.104 7.512 ;
  LAYER M3 ;
        RECT 1.072 7.46 1.104 7.492 ;
  LAYER M1 ;
        RECT 1.136 5.004 1.168 7.512 ;
  LAYER M3 ;
        RECT 1.136 5.024 1.168 5.056 ;
  LAYER M1 ;
        RECT 1.2 5.004 1.232 7.512 ;
  LAYER M3 ;
        RECT 1.2 7.46 1.232 7.492 ;
  LAYER M1 ;
        RECT 1.264 5.004 1.296 7.512 ;
  LAYER M3 ;
        RECT 1.264 5.024 1.296 5.056 ;
  LAYER M1 ;
        RECT 1.328 5.004 1.36 7.512 ;
  LAYER M3 ;
        RECT 1.328 7.46 1.36 7.492 ;
  LAYER M1 ;
        RECT 1.392 5.004 1.424 7.512 ;
  LAYER M3 ;
        RECT 1.392 5.024 1.424 5.056 ;
  LAYER M1 ;
        RECT 1.456 5.004 1.488 7.512 ;
  LAYER M3 ;
        RECT 1.456 7.46 1.488 7.492 ;
  LAYER M1 ;
        RECT 1.52 5.004 1.552 7.512 ;
  LAYER M3 ;
        RECT 1.52 5.024 1.552 5.056 ;
  LAYER M1 ;
        RECT 1.584 5.004 1.616 7.512 ;
  LAYER M3 ;
        RECT 1.584 7.46 1.616 7.492 ;
  LAYER M1 ;
        RECT 1.648 5.004 1.68 7.512 ;
  LAYER M3 ;
        RECT 1.648 5.024 1.68 5.056 ;
  LAYER M1 ;
        RECT 1.712 5.004 1.744 7.512 ;
  LAYER M3 ;
        RECT 1.712 7.46 1.744 7.492 ;
  LAYER M1 ;
        RECT 1.776 5.004 1.808 7.512 ;
  LAYER M3 ;
        RECT 1.776 5.024 1.808 5.056 ;
  LAYER M1 ;
        RECT 1.84 5.004 1.872 7.512 ;
  LAYER M3 ;
        RECT 1.84 7.46 1.872 7.492 ;
  LAYER M1 ;
        RECT 1.904 5.004 1.936 7.512 ;
  LAYER M3 ;
        RECT 1.904 5.024 1.936 5.056 ;
  LAYER M1 ;
        RECT 1.968 5.004 2 7.512 ;
  LAYER M3 ;
        RECT 1.968 7.46 2 7.492 ;
  LAYER M1 ;
        RECT 2.032 5.004 2.064 7.512 ;
  LAYER M3 ;
        RECT 2.032 5.024 2.064 5.056 ;
  LAYER M1 ;
        RECT 2.096 5.004 2.128 7.512 ;
  LAYER M3 ;
        RECT 2.096 7.46 2.128 7.492 ;
  LAYER M1 ;
        RECT 2.16 5.004 2.192 7.512 ;
  LAYER M3 ;
        RECT 2.16 5.024 2.192 5.056 ;
  LAYER M1 ;
        RECT 2.224 5.004 2.256 7.512 ;
  LAYER M3 ;
        RECT 2.224 7.46 2.256 7.492 ;
  LAYER M1 ;
        RECT 2.288 5.004 2.32 7.512 ;
  LAYER M3 ;
        RECT 2.288 5.024 2.32 5.056 ;
  LAYER M1 ;
        RECT 2.352 5.004 2.384 7.512 ;
  LAYER M3 ;
        RECT 2.352 7.46 2.384 7.492 ;
  LAYER M1 ;
        RECT 2.416 5.004 2.448 7.512 ;
  LAYER M3 ;
        RECT 2.416 5.024 2.448 5.056 ;
  LAYER M1 ;
        RECT 2.48 5.004 2.512 7.512 ;
  LAYER M3 ;
        RECT 2.48 7.46 2.512 7.492 ;
  LAYER M1 ;
        RECT 2.544 5.004 2.576 7.512 ;
  LAYER M3 ;
        RECT 2.544 5.024 2.576 5.056 ;
  LAYER M1 ;
        RECT 2.608 5.004 2.64 7.512 ;
  LAYER M3 ;
        RECT 2.608 7.46 2.64 7.492 ;
  LAYER M1 ;
        RECT 2.672 5.004 2.704 7.512 ;
  LAYER M3 ;
        RECT 2.672 5.024 2.704 5.056 ;
  LAYER M1 ;
        RECT 2.736 5.004 2.768 7.512 ;
  LAYER M3 ;
        RECT 2.736 7.46 2.768 7.492 ;
  LAYER M1 ;
        RECT 2.8 5.004 2.832 7.512 ;
  LAYER M3 ;
        RECT 2.8 5.024 2.832 5.056 ;
  LAYER M1 ;
        RECT 2.864 5.004 2.896 7.512 ;
  LAYER M3 ;
        RECT 2.864 7.46 2.896 7.492 ;
  LAYER M1 ;
        RECT 2.928 5.004 2.96 7.512 ;
  LAYER M3 ;
        RECT 2.928 5.024 2.96 5.056 ;
  LAYER M1 ;
        RECT 2.992 5.004 3.024 7.512 ;
  LAYER M3 ;
        RECT 2.992 7.46 3.024 7.492 ;
  LAYER M1 ;
        RECT 3.056 5.004 3.088 7.512 ;
  LAYER M3 ;
        RECT 0.688 5.088 0.72 5.12 ;
  LAYER M2 ;
        RECT 3.056 5.152 3.088 5.184 ;
  LAYER M2 ;
        RECT 0.688 5.216 0.72 5.248 ;
  LAYER M2 ;
        RECT 3.056 5.28 3.088 5.312 ;
  LAYER M2 ;
        RECT 0.688 5.344 0.72 5.376 ;
  LAYER M2 ;
        RECT 3.056 5.408 3.088 5.44 ;
  LAYER M2 ;
        RECT 0.688 5.472 0.72 5.504 ;
  LAYER M2 ;
        RECT 3.056 5.536 3.088 5.568 ;
  LAYER M2 ;
        RECT 0.688 5.6 0.72 5.632 ;
  LAYER M2 ;
        RECT 3.056 5.664 3.088 5.696 ;
  LAYER M2 ;
        RECT 0.688 5.728 0.72 5.76 ;
  LAYER M2 ;
        RECT 3.056 5.792 3.088 5.824 ;
  LAYER M2 ;
        RECT 0.688 5.856 0.72 5.888 ;
  LAYER M2 ;
        RECT 3.056 5.92 3.088 5.952 ;
  LAYER M2 ;
        RECT 0.688 5.984 0.72 6.016 ;
  LAYER M2 ;
        RECT 3.056 6.048 3.088 6.08 ;
  LAYER M2 ;
        RECT 0.688 6.112 0.72 6.144 ;
  LAYER M2 ;
        RECT 3.056 6.176 3.088 6.208 ;
  LAYER M2 ;
        RECT 0.688 6.24 0.72 6.272 ;
  LAYER M2 ;
        RECT 3.056 6.304 3.088 6.336 ;
  LAYER M2 ;
        RECT 0.688 6.368 0.72 6.4 ;
  LAYER M2 ;
        RECT 3.056 6.432 3.088 6.464 ;
  LAYER M2 ;
        RECT 0.688 6.496 0.72 6.528 ;
  LAYER M2 ;
        RECT 3.056 6.56 3.088 6.592 ;
  LAYER M2 ;
        RECT 0.688 6.624 0.72 6.656 ;
  LAYER M2 ;
        RECT 3.056 6.688 3.088 6.72 ;
  LAYER M2 ;
        RECT 0.688 6.752 0.72 6.784 ;
  LAYER M2 ;
        RECT 3.056 6.816 3.088 6.848 ;
  LAYER M2 ;
        RECT 0.688 6.88 0.72 6.912 ;
  LAYER M2 ;
        RECT 3.056 6.944 3.088 6.976 ;
  LAYER M2 ;
        RECT 0.688 7.008 0.72 7.04 ;
  LAYER M2 ;
        RECT 3.056 7.072 3.088 7.104 ;
  LAYER M2 ;
        RECT 0.688 7.136 0.72 7.168 ;
  LAYER M2 ;
        RECT 3.056 7.2 3.088 7.232 ;
  LAYER M2 ;
        RECT 0.688 7.264 0.72 7.296 ;
  LAYER M2 ;
        RECT 3.056 7.328 3.088 7.36 ;
  LAYER M2 ;
        RECT 0.64 4.956 3.136 7.56 ;
  LAYER M1 ;
        RECT 0.688 8.112 0.72 10.62 ;
  LAYER M3 ;
        RECT 0.688 10.568 0.72 10.6 ;
  LAYER M1 ;
        RECT 0.752 8.112 0.784 10.62 ;
  LAYER M3 ;
        RECT 0.752 8.132 0.784 8.164 ;
  LAYER M1 ;
        RECT 0.816 8.112 0.848 10.62 ;
  LAYER M3 ;
        RECT 0.816 10.568 0.848 10.6 ;
  LAYER M1 ;
        RECT 0.88 8.112 0.912 10.62 ;
  LAYER M3 ;
        RECT 0.88 8.132 0.912 8.164 ;
  LAYER M1 ;
        RECT 0.944 8.112 0.976 10.62 ;
  LAYER M3 ;
        RECT 0.944 10.568 0.976 10.6 ;
  LAYER M1 ;
        RECT 1.008 8.112 1.04 10.62 ;
  LAYER M3 ;
        RECT 1.008 8.132 1.04 8.164 ;
  LAYER M1 ;
        RECT 1.072 8.112 1.104 10.62 ;
  LAYER M3 ;
        RECT 1.072 10.568 1.104 10.6 ;
  LAYER M1 ;
        RECT 1.136 8.112 1.168 10.62 ;
  LAYER M3 ;
        RECT 1.136 8.132 1.168 8.164 ;
  LAYER M1 ;
        RECT 1.2 8.112 1.232 10.62 ;
  LAYER M3 ;
        RECT 1.2 10.568 1.232 10.6 ;
  LAYER M1 ;
        RECT 1.264 8.112 1.296 10.62 ;
  LAYER M3 ;
        RECT 1.264 8.132 1.296 8.164 ;
  LAYER M1 ;
        RECT 1.328 8.112 1.36 10.62 ;
  LAYER M3 ;
        RECT 1.328 10.568 1.36 10.6 ;
  LAYER M1 ;
        RECT 1.392 8.112 1.424 10.62 ;
  LAYER M3 ;
        RECT 1.392 8.132 1.424 8.164 ;
  LAYER M1 ;
        RECT 1.456 8.112 1.488 10.62 ;
  LAYER M3 ;
        RECT 1.456 10.568 1.488 10.6 ;
  LAYER M1 ;
        RECT 1.52 8.112 1.552 10.62 ;
  LAYER M3 ;
        RECT 1.52 8.132 1.552 8.164 ;
  LAYER M1 ;
        RECT 1.584 8.112 1.616 10.62 ;
  LAYER M3 ;
        RECT 1.584 10.568 1.616 10.6 ;
  LAYER M1 ;
        RECT 1.648 8.112 1.68 10.62 ;
  LAYER M3 ;
        RECT 1.648 8.132 1.68 8.164 ;
  LAYER M1 ;
        RECT 1.712 8.112 1.744 10.62 ;
  LAYER M3 ;
        RECT 1.712 10.568 1.744 10.6 ;
  LAYER M1 ;
        RECT 1.776 8.112 1.808 10.62 ;
  LAYER M3 ;
        RECT 1.776 8.132 1.808 8.164 ;
  LAYER M1 ;
        RECT 1.84 8.112 1.872 10.62 ;
  LAYER M3 ;
        RECT 1.84 10.568 1.872 10.6 ;
  LAYER M1 ;
        RECT 1.904 8.112 1.936 10.62 ;
  LAYER M3 ;
        RECT 1.904 8.132 1.936 8.164 ;
  LAYER M1 ;
        RECT 1.968 8.112 2 10.62 ;
  LAYER M3 ;
        RECT 1.968 10.568 2 10.6 ;
  LAYER M1 ;
        RECT 2.032 8.112 2.064 10.62 ;
  LAYER M3 ;
        RECT 2.032 8.132 2.064 8.164 ;
  LAYER M1 ;
        RECT 2.096 8.112 2.128 10.62 ;
  LAYER M3 ;
        RECT 2.096 10.568 2.128 10.6 ;
  LAYER M1 ;
        RECT 2.16 8.112 2.192 10.62 ;
  LAYER M3 ;
        RECT 2.16 8.132 2.192 8.164 ;
  LAYER M1 ;
        RECT 2.224 8.112 2.256 10.62 ;
  LAYER M3 ;
        RECT 2.224 10.568 2.256 10.6 ;
  LAYER M1 ;
        RECT 2.288 8.112 2.32 10.62 ;
  LAYER M3 ;
        RECT 2.288 8.132 2.32 8.164 ;
  LAYER M1 ;
        RECT 2.352 8.112 2.384 10.62 ;
  LAYER M3 ;
        RECT 2.352 10.568 2.384 10.6 ;
  LAYER M1 ;
        RECT 2.416 8.112 2.448 10.62 ;
  LAYER M3 ;
        RECT 2.416 8.132 2.448 8.164 ;
  LAYER M1 ;
        RECT 2.48 8.112 2.512 10.62 ;
  LAYER M3 ;
        RECT 2.48 10.568 2.512 10.6 ;
  LAYER M1 ;
        RECT 2.544 8.112 2.576 10.62 ;
  LAYER M3 ;
        RECT 2.544 8.132 2.576 8.164 ;
  LAYER M1 ;
        RECT 2.608 8.112 2.64 10.62 ;
  LAYER M3 ;
        RECT 2.608 10.568 2.64 10.6 ;
  LAYER M1 ;
        RECT 2.672 8.112 2.704 10.62 ;
  LAYER M3 ;
        RECT 2.672 8.132 2.704 8.164 ;
  LAYER M1 ;
        RECT 2.736 8.112 2.768 10.62 ;
  LAYER M3 ;
        RECT 2.736 10.568 2.768 10.6 ;
  LAYER M1 ;
        RECT 2.8 8.112 2.832 10.62 ;
  LAYER M3 ;
        RECT 2.8 8.132 2.832 8.164 ;
  LAYER M1 ;
        RECT 2.864 8.112 2.896 10.62 ;
  LAYER M3 ;
        RECT 2.864 10.568 2.896 10.6 ;
  LAYER M1 ;
        RECT 2.928 8.112 2.96 10.62 ;
  LAYER M3 ;
        RECT 2.928 8.132 2.96 8.164 ;
  LAYER M1 ;
        RECT 2.992 8.112 3.024 10.62 ;
  LAYER M3 ;
        RECT 2.992 10.568 3.024 10.6 ;
  LAYER M1 ;
        RECT 3.056 8.112 3.088 10.62 ;
  LAYER M3 ;
        RECT 0.688 8.196 0.72 8.228 ;
  LAYER M2 ;
        RECT 3.056 8.26 3.088 8.292 ;
  LAYER M2 ;
        RECT 0.688 8.324 0.72 8.356 ;
  LAYER M2 ;
        RECT 3.056 8.388 3.088 8.42 ;
  LAYER M2 ;
        RECT 0.688 8.452 0.72 8.484 ;
  LAYER M2 ;
        RECT 3.056 8.516 3.088 8.548 ;
  LAYER M2 ;
        RECT 0.688 8.58 0.72 8.612 ;
  LAYER M2 ;
        RECT 3.056 8.644 3.088 8.676 ;
  LAYER M2 ;
        RECT 0.688 8.708 0.72 8.74 ;
  LAYER M2 ;
        RECT 3.056 8.772 3.088 8.804 ;
  LAYER M2 ;
        RECT 0.688 8.836 0.72 8.868 ;
  LAYER M2 ;
        RECT 3.056 8.9 3.088 8.932 ;
  LAYER M2 ;
        RECT 0.688 8.964 0.72 8.996 ;
  LAYER M2 ;
        RECT 3.056 9.028 3.088 9.06 ;
  LAYER M2 ;
        RECT 0.688 9.092 0.72 9.124 ;
  LAYER M2 ;
        RECT 3.056 9.156 3.088 9.188 ;
  LAYER M2 ;
        RECT 0.688 9.22 0.72 9.252 ;
  LAYER M2 ;
        RECT 3.056 9.284 3.088 9.316 ;
  LAYER M2 ;
        RECT 0.688 9.348 0.72 9.38 ;
  LAYER M2 ;
        RECT 3.056 9.412 3.088 9.444 ;
  LAYER M2 ;
        RECT 0.688 9.476 0.72 9.508 ;
  LAYER M2 ;
        RECT 3.056 9.54 3.088 9.572 ;
  LAYER M2 ;
        RECT 0.688 9.604 0.72 9.636 ;
  LAYER M2 ;
        RECT 3.056 9.668 3.088 9.7 ;
  LAYER M2 ;
        RECT 0.688 9.732 0.72 9.764 ;
  LAYER M2 ;
        RECT 3.056 9.796 3.088 9.828 ;
  LAYER M2 ;
        RECT 0.688 9.86 0.72 9.892 ;
  LAYER M2 ;
        RECT 3.056 9.924 3.088 9.956 ;
  LAYER M2 ;
        RECT 0.688 9.988 0.72 10.02 ;
  LAYER M2 ;
        RECT 3.056 10.052 3.088 10.084 ;
  LAYER M2 ;
        RECT 0.688 10.116 0.72 10.148 ;
  LAYER M2 ;
        RECT 3.056 10.18 3.088 10.212 ;
  LAYER M2 ;
        RECT 0.688 10.244 0.72 10.276 ;
  LAYER M2 ;
        RECT 3.056 10.308 3.088 10.34 ;
  LAYER M2 ;
        RECT 0.688 10.372 0.72 10.404 ;
  LAYER M2 ;
        RECT 3.056 10.436 3.088 10.468 ;
  LAYER M2 ;
        RECT 0.64 8.064 3.136 10.668 ;
  LAYER M1 ;
        RECT 0.688 11.22 0.72 13.728 ;
  LAYER M3 ;
        RECT 0.688 13.676 0.72 13.708 ;
  LAYER M1 ;
        RECT 0.752 11.22 0.784 13.728 ;
  LAYER M3 ;
        RECT 0.752 11.24 0.784 11.272 ;
  LAYER M1 ;
        RECT 0.816 11.22 0.848 13.728 ;
  LAYER M3 ;
        RECT 0.816 13.676 0.848 13.708 ;
  LAYER M1 ;
        RECT 0.88 11.22 0.912 13.728 ;
  LAYER M3 ;
        RECT 0.88 11.24 0.912 11.272 ;
  LAYER M1 ;
        RECT 0.944 11.22 0.976 13.728 ;
  LAYER M3 ;
        RECT 0.944 13.676 0.976 13.708 ;
  LAYER M1 ;
        RECT 1.008 11.22 1.04 13.728 ;
  LAYER M3 ;
        RECT 1.008 11.24 1.04 11.272 ;
  LAYER M1 ;
        RECT 1.072 11.22 1.104 13.728 ;
  LAYER M3 ;
        RECT 1.072 13.676 1.104 13.708 ;
  LAYER M1 ;
        RECT 1.136 11.22 1.168 13.728 ;
  LAYER M3 ;
        RECT 1.136 11.24 1.168 11.272 ;
  LAYER M1 ;
        RECT 1.2 11.22 1.232 13.728 ;
  LAYER M3 ;
        RECT 1.2 13.676 1.232 13.708 ;
  LAYER M1 ;
        RECT 1.264 11.22 1.296 13.728 ;
  LAYER M3 ;
        RECT 1.264 11.24 1.296 11.272 ;
  LAYER M1 ;
        RECT 1.328 11.22 1.36 13.728 ;
  LAYER M3 ;
        RECT 1.328 13.676 1.36 13.708 ;
  LAYER M1 ;
        RECT 1.392 11.22 1.424 13.728 ;
  LAYER M3 ;
        RECT 1.392 11.24 1.424 11.272 ;
  LAYER M1 ;
        RECT 1.456 11.22 1.488 13.728 ;
  LAYER M3 ;
        RECT 1.456 13.676 1.488 13.708 ;
  LAYER M1 ;
        RECT 1.52 11.22 1.552 13.728 ;
  LAYER M3 ;
        RECT 1.52 11.24 1.552 11.272 ;
  LAYER M1 ;
        RECT 1.584 11.22 1.616 13.728 ;
  LAYER M3 ;
        RECT 1.584 13.676 1.616 13.708 ;
  LAYER M1 ;
        RECT 1.648 11.22 1.68 13.728 ;
  LAYER M3 ;
        RECT 1.648 11.24 1.68 11.272 ;
  LAYER M1 ;
        RECT 1.712 11.22 1.744 13.728 ;
  LAYER M3 ;
        RECT 1.712 13.676 1.744 13.708 ;
  LAYER M1 ;
        RECT 1.776 11.22 1.808 13.728 ;
  LAYER M3 ;
        RECT 1.776 11.24 1.808 11.272 ;
  LAYER M1 ;
        RECT 1.84 11.22 1.872 13.728 ;
  LAYER M3 ;
        RECT 1.84 13.676 1.872 13.708 ;
  LAYER M1 ;
        RECT 1.904 11.22 1.936 13.728 ;
  LAYER M3 ;
        RECT 1.904 11.24 1.936 11.272 ;
  LAYER M1 ;
        RECT 1.968 11.22 2 13.728 ;
  LAYER M3 ;
        RECT 1.968 13.676 2 13.708 ;
  LAYER M1 ;
        RECT 2.032 11.22 2.064 13.728 ;
  LAYER M3 ;
        RECT 2.032 11.24 2.064 11.272 ;
  LAYER M1 ;
        RECT 2.096 11.22 2.128 13.728 ;
  LAYER M3 ;
        RECT 2.096 13.676 2.128 13.708 ;
  LAYER M1 ;
        RECT 2.16 11.22 2.192 13.728 ;
  LAYER M3 ;
        RECT 2.16 11.24 2.192 11.272 ;
  LAYER M1 ;
        RECT 2.224 11.22 2.256 13.728 ;
  LAYER M3 ;
        RECT 2.224 13.676 2.256 13.708 ;
  LAYER M1 ;
        RECT 2.288 11.22 2.32 13.728 ;
  LAYER M3 ;
        RECT 2.288 11.24 2.32 11.272 ;
  LAYER M1 ;
        RECT 2.352 11.22 2.384 13.728 ;
  LAYER M3 ;
        RECT 2.352 13.676 2.384 13.708 ;
  LAYER M1 ;
        RECT 2.416 11.22 2.448 13.728 ;
  LAYER M3 ;
        RECT 2.416 11.24 2.448 11.272 ;
  LAYER M1 ;
        RECT 2.48 11.22 2.512 13.728 ;
  LAYER M3 ;
        RECT 2.48 13.676 2.512 13.708 ;
  LAYER M1 ;
        RECT 2.544 11.22 2.576 13.728 ;
  LAYER M3 ;
        RECT 2.544 11.24 2.576 11.272 ;
  LAYER M1 ;
        RECT 2.608 11.22 2.64 13.728 ;
  LAYER M3 ;
        RECT 2.608 13.676 2.64 13.708 ;
  LAYER M1 ;
        RECT 2.672 11.22 2.704 13.728 ;
  LAYER M3 ;
        RECT 2.672 11.24 2.704 11.272 ;
  LAYER M1 ;
        RECT 2.736 11.22 2.768 13.728 ;
  LAYER M3 ;
        RECT 2.736 13.676 2.768 13.708 ;
  LAYER M1 ;
        RECT 2.8 11.22 2.832 13.728 ;
  LAYER M3 ;
        RECT 2.8 11.24 2.832 11.272 ;
  LAYER M1 ;
        RECT 2.864 11.22 2.896 13.728 ;
  LAYER M3 ;
        RECT 2.864 13.676 2.896 13.708 ;
  LAYER M1 ;
        RECT 2.928 11.22 2.96 13.728 ;
  LAYER M3 ;
        RECT 2.928 11.24 2.96 11.272 ;
  LAYER M1 ;
        RECT 2.992 11.22 3.024 13.728 ;
  LAYER M3 ;
        RECT 2.992 13.676 3.024 13.708 ;
  LAYER M1 ;
        RECT 3.056 11.22 3.088 13.728 ;
  LAYER M3 ;
        RECT 0.688 11.304 0.72 11.336 ;
  LAYER M2 ;
        RECT 3.056 11.368 3.088 11.4 ;
  LAYER M2 ;
        RECT 0.688 11.432 0.72 11.464 ;
  LAYER M2 ;
        RECT 3.056 11.496 3.088 11.528 ;
  LAYER M2 ;
        RECT 0.688 11.56 0.72 11.592 ;
  LAYER M2 ;
        RECT 3.056 11.624 3.088 11.656 ;
  LAYER M2 ;
        RECT 0.688 11.688 0.72 11.72 ;
  LAYER M2 ;
        RECT 3.056 11.752 3.088 11.784 ;
  LAYER M2 ;
        RECT 0.688 11.816 0.72 11.848 ;
  LAYER M2 ;
        RECT 3.056 11.88 3.088 11.912 ;
  LAYER M2 ;
        RECT 0.688 11.944 0.72 11.976 ;
  LAYER M2 ;
        RECT 3.056 12.008 3.088 12.04 ;
  LAYER M2 ;
        RECT 0.688 12.072 0.72 12.104 ;
  LAYER M2 ;
        RECT 3.056 12.136 3.088 12.168 ;
  LAYER M2 ;
        RECT 0.688 12.2 0.72 12.232 ;
  LAYER M2 ;
        RECT 3.056 12.264 3.088 12.296 ;
  LAYER M2 ;
        RECT 0.688 12.328 0.72 12.36 ;
  LAYER M2 ;
        RECT 3.056 12.392 3.088 12.424 ;
  LAYER M2 ;
        RECT 0.688 12.456 0.72 12.488 ;
  LAYER M2 ;
        RECT 3.056 12.52 3.088 12.552 ;
  LAYER M2 ;
        RECT 0.688 12.584 0.72 12.616 ;
  LAYER M2 ;
        RECT 3.056 12.648 3.088 12.68 ;
  LAYER M2 ;
        RECT 0.688 12.712 0.72 12.744 ;
  LAYER M2 ;
        RECT 3.056 12.776 3.088 12.808 ;
  LAYER M2 ;
        RECT 0.688 12.84 0.72 12.872 ;
  LAYER M2 ;
        RECT 3.056 12.904 3.088 12.936 ;
  LAYER M2 ;
        RECT 0.688 12.968 0.72 13 ;
  LAYER M2 ;
        RECT 3.056 13.032 3.088 13.064 ;
  LAYER M2 ;
        RECT 0.688 13.096 0.72 13.128 ;
  LAYER M2 ;
        RECT 3.056 13.16 3.088 13.192 ;
  LAYER M2 ;
        RECT 0.688 13.224 0.72 13.256 ;
  LAYER M2 ;
        RECT 3.056 13.288 3.088 13.32 ;
  LAYER M2 ;
        RECT 0.688 13.352 0.72 13.384 ;
  LAYER M2 ;
        RECT 3.056 13.416 3.088 13.448 ;
  LAYER M2 ;
        RECT 0.688 13.48 0.72 13.512 ;
  LAYER M2 ;
        RECT 3.056 13.544 3.088 13.576 ;
  LAYER M2 ;
        RECT 0.64 11.172 3.136 13.776 ;
  LAYER M1 ;
        RECT 3.664 1.896 3.696 4.404 ;
  LAYER M3 ;
        RECT 3.664 4.352 3.696 4.384 ;
  LAYER M1 ;
        RECT 3.728 1.896 3.76 4.404 ;
  LAYER M3 ;
        RECT 3.728 1.916 3.76 1.948 ;
  LAYER M1 ;
        RECT 3.792 1.896 3.824 4.404 ;
  LAYER M3 ;
        RECT 3.792 4.352 3.824 4.384 ;
  LAYER M1 ;
        RECT 3.856 1.896 3.888 4.404 ;
  LAYER M3 ;
        RECT 3.856 1.916 3.888 1.948 ;
  LAYER M1 ;
        RECT 3.92 1.896 3.952 4.404 ;
  LAYER M3 ;
        RECT 3.92 4.352 3.952 4.384 ;
  LAYER M1 ;
        RECT 3.984 1.896 4.016 4.404 ;
  LAYER M3 ;
        RECT 3.984 1.916 4.016 1.948 ;
  LAYER M1 ;
        RECT 4.048 1.896 4.08 4.404 ;
  LAYER M3 ;
        RECT 4.048 4.352 4.08 4.384 ;
  LAYER M1 ;
        RECT 4.112 1.896 4.144 4.404 ;
  LAYER M3 ;
        RECT 4.112 1.916 4.144 1.948 ;
  LAYER M1 ;
        RECT 4.176 1.896 4.208 4.404 ;
  LAYER M3 ;
        RECT 4.176 4.352 4.208 4.384 ;
  LAYER M1 ;
        RECT 4.24 1.896 4.272 4.404 ;
  LAYER M3 ;
        RECT 4.24 1.916 4.272 1.948 ;
  LAYER M1 ;
        RECT 4.304 1.896 4.336 4.404 ;
  LAYER M3 ;
        RECT 4.304 4.352 4.336 4.384 ;
  LAYER M1 ;
        RECT 4.368 1.896 4.4 4.404 ;
  LAYER M3 ;
        RECT 4.368 1.916 4.4 1.948 ;
  LAYER M1 ;
        RECT 4.432 1.896 4.464 4.404 ;
  LAYER M3 ;
        RECT 4.432 4.352 4.464 4.384 ;
  LAYER M1 ;
        RECT 4.496 1.896 4.528 4.404 ;
  LAYER M3 ;
        RECT 4.496 1.916 4.528 1.948 ;
  LAYER M1 ;
        RECT 4.56 1.896 4.592 4.404 ;
  LAYER M3 ;
        RECT 4.56 4.352 4.592 4.384 ;
  LAYER M1 ;
        RECT 4.624 1.896 4.656 4.404 ;
  LAYER M3 ;
        RECT 4.624 1.916 4.656 1.948 ;
  LAYER M1 ;
        RECT 4.688 1.896 4.72 4.404 ;
  LAYER M3 ;
        RECT 4.688 4.352 4.72 4.384 ;
  LAYER M1 ;
        RECT 4.752 1.896 4.784 4.404 ;
  LAYER M3 ;
        RECT 4.752 1.916 4.784 1.948 ;
  LAYER M1 ;
        RECT 4.816 1.896 4.848 4.404 ;
  LAYER M3 ;
        RECT 4.816 4.352 4.848 4.384 ;
  LAYER M1 ;
        RECT 4.88 1.896 4.912 4.404 ;
  LAYER M3 ;
        RECT 4.88 1.916 4.912 1.948 ;
  LAYER M1 ;
        RECT 4.944 1.896 4.976 4.404 ;
  LAYER M3 ;
        RECT 4.944 4.352 4.976 4.384 ;
  LAYER M1 ;
        RECT 5.008 1.896 5.04 4.404 ;
  LAYER M3 ;
        RECT 5.008 1.916 5.04 1.948 ;
  LAYER M1 ;
        RECT 5.072 1.896 5.104 4.404 ;
  LAYER M3 ;
        RECT 5.072 4.352 5.104 4.384 ;
  LAYER M1 ;
        RECT 5.136 1.896 5.168 4.404 ;
  LAYER M3 ;
        RECT 5.136 1.916 5.168 1.948 ;
  LAYER M1 ;
        RECT 5.2 1.896 5.232 4.404 ;
  LAYER M3 ;
        RECT 5.2 4.352 5.232 4.384 ;
  LAYER M1 ;
        RECT 5.264 1.896 5.296 4.404 ;
  LAYER M3 ;
        RECT 5.264 1.916 5.296 1.948 ;
  LAYER M1 ;
        RECT 5.328 1.896 5.36 4.404 ;
  LAYER M3 ;
        RECT 5.328 4.352 5.36 4.384 ;
  LAYER M1 ;
        RECT 5.392 1.896 5.424 4.404 ;
  LAYER M3 ;
        RECT 5.392 1.916 5.424 1.948 ;
  LAYER M1 ;
        RECT 5.456 1.896 5.488 4.404 ;
  LAYER M3 ;
        RECT 5.456 4.352 5.488 4.384 ;
  LAYER M1 ;
        RECT 5.52 1.896 5.552 4.404 ;
  LAYER M3 ;
        RECT 5.52 1.916 5.552 1.948 ;
  LAYER M1 ;
        RECT 5.584 1.896 5.616 4.404 ;
  LAYER M3 ;
        RECT 5.584 4.352 5.616 4.384 ;
  LAYER M1 ;
        RECT 5.648 1.896 5.68 4.404 ;
  LAYER M3 ;
        RECT 5.648 1.916 5.68 1.948 ;
  LAYER M1 ;
        RECT 5.712 1.896 5.744 4.404 ;
  LAYER M3 ;
        RECT 5.712 4.352 5.744 4.384 ;
  LAYER M1 ;
        RECT 5.776 1.896 5.808 4.404 ;
  LAYER M3 ;
        RECT 5.776 1.916 5.808 1.948 ;
  LAYER M1 ;
        RECT 5.84 1.896 5.872 4.404 ;
  LAYER M3 ;
        RECT 5.84 4.352 5.872 4.384 ;
  LAYER M1 ;
        RECT 5.904 1.896 5.936 4.404 ;
  LAYER M3 ;
        RECT 5.904 1.916 5.936 1.948 ;
  LAYER M1 ;
        RECT 5.968 1.896 6 4.404 ;
  LAYER M3 ;
        RECT 5.968 4.352 6 4.384 ;
  LAYER M1 ;
        RECT 6.032 1.896 6.064 4.404 ;
  LAYER M3 ;
        RECT 3.664 1.98 3.696 2.012 ;
  LAYER M2 ;
        RECT 6.032 2.044 6.064 2.076 ;
  LAYER M2 ;
        RECT 3.664 2.108 3.696 2.14 ;
  LAYER M2 ;
        RECT 6.032 2.172 6.064 2.204 ;
  LAYER M2 ;
        RECT 3.664 2.236 3.696 2.268 ;
  LAYER M2 ;
        RECT 6.032 2.3 6.064 2.332 ;
  LAYER M2 ;
        RECT 3.664 2.364 3.696 2.396 ;
  LAYER M2 ;
        RECT 6.032 2.428 6.064 2.46 ;
  LAYER M2 ;
        RECT 3.664 2.492 3.696 2.524 ;
  LAYER M2 ;
        RECT 6.032 2.556 6.064 2.588 ;
  LAYER M2 ;
        RECT 3.664 2.62 3.696 2.652 ;
  LAYER M2 ;
        RECT 6.032 2.684 6.064 2.716 ;
  LAYER M2 ;
        RECT 3.664 2.748 3.696 2.78 ;
  LAYER M2 ;
        RECT 6.032 2.812 6.064 2.844 ;
  LAYER M2 ;
        RECT 3.664 2.876 3.696 2.908 ;
  LAYER M2 ;
        RECT 6.032 2.94 6.064 2.972 ;
  LAYER M2 ;
        RECT 3.664 3.004 3.696 3.036 ;
  LAYER M2 ;
        RECT 6.032 3.068 6.064 3.1 ;
  LAYER M2 ;
        RECT 3.664 3.132 3.696 3.164 ;
  LAYER M2 ;
        RECT 6.032 3.196 6.064 3.228 ;
  LAYER M2 ;
        RECT 3.664 3.26 3.696 3.292 ;
  LAYER M2 ;
        RECT 6.032 3.324 6.064 3.356 ;
  LAYER M2 ;
        RECT 3.664 3.388 3.696 3.42 ;
  LAYER M2 ;
        RECT 6.032 3.452 6.064 3.484 ;
  LAYER M2 ;
        RECT 3.664 3.516 3.696 3.548 ;
  LAYER M2 ;
        RECT 6.032 3.58 6.064 3.612 ;
  LAYER M2 ;
        RECT 3.664 3.644 3.696 3.676 ;
  LAYER M2 ;
        RECT 6.032 3.708 6.064 3.74 ;
  LAYER M2 ;
        RECT 3.664 3.772 3.696 3.804 ;
  LAYER M2 ;
        RECT 6.032 3.836 6.064 3.868 ;
  LAYER M2 ;
        RECT 3.664 3.9 3.696 3.932 ;
  LAYER M2 ;
        RECT 6.032 3.964 6.064 3.996 ;
  LAYER M2 ;
        RECT 3.664 4.028 3.696 4.06 ;
  LAYER M2 ;
        RECT 6.032 4.092 6.064 4.124 ;
  LAYER M2 ;
        RECT 3.664 4.156 3.696 4.188 ;
  LAYER M2 ;
        RECT 6.032 4.22 6.064 4.252 ;
  LAYER M2 ;
        RECT 3.616 1.848 6.112 4.452 ;
  LAYER M1 ;
        RECT 3.664 5.004 3.696 7.512 ;
  LAYER M3 ;
        RECT 3.664 7.46 3.696 7.492 ;
  LAYER M1 ;
        RECT 3.728 5.004 3.76 7.512 ;
  LAYER M3 ;
        RECT 3.728 5.024 3.76 5.056 ;
  LAYER M1 ;
        RECT 3.792 5.004 3.824 7.512 ;
  LAYER M3 ;
        RECT 3.792 7.46 3.824 7.492 ;
  LAYER M1 ;
        RECT 3.856 5.004 3.888 7.512 ;
  LAYER M3 ;
        RECT 3.856 5.024 3.888 5.056 ;
  LAYER M1 ;
        RECT 3.92 5.004 3.952 7.512 ;
  LAYER M3 ;
        RECT 3.92 7.46 3.952 7.492 ;
  LAYER M1 ;
        RECT 3.984 5.004 4.016 7.512 ;
  LAYER M3 ;
        RECT 3.984 5.024 4.016 5.056 ;
  LAYER M1 ;
        RECT 4.048 5.004 4.08 7.512 ;
  LAYER M3 ;
        RECT 4.048 7.46 4.08 7.492 ;
  LAYER M1 ;
        RECT 4.112 5.004 4.144 7.512 ;
  LAYER M3 ;
        RECT 4.112 5.024 4.144 5.056 ;
  LAYER M1 ;
        RECT 4.176 5.004 4.208 7.512 ;
  LAYER M3 ;
        RECT 4.176 7.46 4.208 7.492 ;
  LAYER M1 ;
        RECT 4.24 5.004 4.272 7.512 ;
  LAYER M3 ;
        RECT 4.24 5.024 4.272 5.056 ;
  LAYER M1 ;
        RECT 4.304 5.004 4.336 7.512 ;
  LAYER M3 ;
        RECT 4.304 7.46 4.336 7.492 ;
  LAYER M1 ;
        RECT 4.368 5.004 4.4 7.512 ;
  LAYER M3 ;
        RECT 4.368 5.024 4.4 5.056 ;
  LAYER M1 ;
        RECT 4.432 5.004 4.464 7.512 ;
  LAYER M3 ;
        RECT 4.432 7.46 4.464 7.492 ;
  LAYER M1 ;
        RECT 4.496 5.004 4.528 7.512 ;
  LAYER M3 ;
        RECT 4.496 5.024 4.528 5.056 ;
  LAYER M1 ;
        RECT 4.56 5.004 4.592 7.512 ;
  LAYER M3 ;
        RECT 4.56 7.46 4.592 7.492 ;
  LAYER M1 ;
        RECT 4.624 5.004 4.656 7.512 ;
  LAYER M3 ;
        RECT 4.624 5.024 4.656 5.056 ;
  LAYER M1 ;
        RECT 4.688 5.004 4.72 7.512 ;
  LAYER M3 ;
        RECT 4.688 7.46 4.72 7.492 ;
  LAYER M1 ;
        RECT 4.752 5.004 4.784 7.512 ;
  LAYER M3 ;
        RECT 4.752 5.024 4.784 5.056 ;
  LAYER M1 ;
        RECT 4.816 5.004 4.848 7.512 ;
  LAYER M3 ;
        RECT 4.816 7.46 4.848 7.492 ;
  LAYER M1 ;
        RECT 4.88 5.004 4.912 7.512 ;
  LAYER M3 ;
        RECT 4.88 5.024 4.912 5.056 ;
  LAYER M1 ;
        RECT 4.944 5.004 4.976 7.512 ;
  LAYER M3 ;
        RECT 4.944 7.46 4.976 7.492 ;
  LAYER M1 ;
        RECT 5.008 5.004 5.04 7.512 ;
  LAYER M3 ;
        RECT 5.008 5.024 5.04 5.056 ;
  LAYER M1 ;
        RECT 5.072 5.004 5.104 7.512 ;
  LAYER M3 ;
        RECT 5.072 7.46 5.104 7.492 ;
  LAYER M1 ;
        RECT 5.136 5.004 5.168 7.512 ;
  LAYER M3 ;
        RECT 5.136 5.024 5.168 5.056 ;
  LAYER M1 ;
        RECT 5.2 5.004 5.232 7.512 ;
  LAYER M3 ;
        RECT 5.2 7.46 5.232 7.492 ;
  LAYER M1 ;
        RECT 5.264 5.004 5.296 7.512 ;
  LAYER M3 ;
        RECT 5.264 5.024 5.296 5.056 ;
  LAYER M1 ;
        RECT 5.328 5.004 5.36 7.512 ;
  LAYER M3 ;
        RECT 5.328 7.46 5.36 7.492 ;
  LAYER M1 ;
        RECT 5.392 5.004 5.424 7.512 ;
  LAYER M3 ;
        RECT 5.392 5.024 5.424 5.056 ;
  LAYER M1 ;
        RECT 5.456 5.004 5.488 7.512 ;
  LAYER M3 ;
        RECT 5.456 7.46 5.488 7.492 ;
  LAYER M1 ;
        RECT 5.52 5.004 5.552 7.512 ;
  LAYER M3 ;
        RECT 5.52 5.024 5.552 5.056 ;
  LAYER M1 ;
        RECT 5.584 5.004 5.616 7.512 ;
  LAYER M3 ;
        RECT 5.584 7.46 5.616 7.492 ;
  LAYER M1 ;
        RECT 5.648 5.004 5.68 7.512 ;
  LAYER M3 ;
        RECT 5.648 5.024 5.68 5.056 ;
  LAYER M1 ;
        RECT 5.712 5.004 5.744 7.512 ;
  LAYER M3 ;
        RECT 5.712 7.46 5.744 7.492 ;
  LAYER M1 ;
        RECT 5.776 5.004 5.808 7.512 ;
  LAYER M3 ;
        RECT 5.776 5.024 5.808 5.056 ;
  LAYER M1 ;
        RECT 5.84 5.004 5.872 7.512 ;
  LAYER M3 ;
        RECT 5.84 7.46 5.872 7.492 ;
  LAYER M1 ;
        RECT 5.904 5.004 5.936 7.512 ;
  LAYER M3 ;
        RECT 5.904 5.024 5.936 5.056 ;
  LAYER M1 ;
        RECT 5.968 5.004 6 7.512 ;
  LAYER M3 ;
        RECT 5.968 7.46 6 7.492 ;
  LAYER M1 ;
        RECT 6.032 5.004 6.064 7.512 ;
  LAYER M3 ;
        RECT 3.664 5.088 3.696 5.12 ;
  LAYER M2 ;
        RECT 6.032 5.152 6.064 5.184 ;
  LAYER M2 ;
        RECT 3.664 5.216 3.696 5.248 ;
  LAYER M2 ;
        RECT 6.032 5.28 6.064 5.312 ;
  LAYER M2 ;
        RECT 3.664 5.344 3.696 5.376 ;
  LAYER M2 ;
        RECT 6.032 5.408 6.064 5.44 ;
  LAYER M2 ;
        RECT 3.664 5.472 3.696 5.504 ;
  LAYER M2 ;
        RECT 6.032 5.536 6.064 5.568 ;
  LAYER M2 ;
        RECT 3.664 5.6 3.696 5.632 ;
  LAYER M2 ;
        RECT 6.032 5.664 6.064 5.696 ;
  LAYER M2 ;
        RECT 3.664 5.728 3.696 5.76 ;
  LAYER M2 ;
        RECT 6.032 5.792 6.064 5.824 ;
  LAYER M2 ;
        RECT 3.664 5.856 3.696 5.888 ;
  LAYER M2 ;
        RECT 6.032 5.92 6.064 5.952 ;
  LAYER M2 ;
        RECT 3.664 5.984 3.696 6.016 ;
  LAYER M2 ;
        RECT 6.032 6.048 6.064 6.08 ;
  LAYER M2 ;
        RECT 3.664 6.112 3.696 6.144 ;
  LAYER M2 ;
        RECT 6.032 6.176 6.064 6.208 ;
  LAYER M2 ;
        RECT 3.664 6.24 3.696 6.272 ;
  LAYER M2 ;
        RECT 6.032 6.304 6.064 6.336 ;
  LAYER M2 ;
        RECT 3.664 6.368 3.696 6.4 ;
  LAYER M2 ;
        RECT 6.032 6.432 6.064 6.464 ;
  LAYER M2 ;
        RECT 3.664 6.496 3.696 6.528 ;
  LAYER M2 ;
        RECT 6.032 6.56 6.064 6.592 ;
  LAYER M2 ;
        RECT 3.664 6.624 3.696 6.656 ;
  LAYER M2 ;
        RECT 6.032 6.688 6.064 6.72 ;
  LAYER M2 ;
        RECT 3.664 6.752 3.696 6.784 ;
  LAYER M2 ;
        RECT 6.032 6.816 6.064 6.848 ;
  LAYER M2 ;
        RECT 3.664 6.88 3.696 6.912 ;
  LAYER M2 ;
        RECT 6.032 6.944 6.064 6.976 ;
  LAYER M2 ;
        RECT 3.664 7.008 3.696 7.04 ;
  LAYER M2 ;
        RECT 6.032 7.072 6.064 7.104 ;
  LAYER M2 ;
        RECT 3.664 7.136 3.696 7.168 ;
  LAYER M2 ;
        RECT 6.032 7.2 6.064 7.232 ;
  LAYER M2 ;
        RECT 3.664 7.264 3.696 7.296 ;
  LAYER M2 ;
        RECT 6.032 7.328 6.064 7.36 ;
  LAYER M2 ;
        RECT 3.616 4.956 6.112 7.56 ;
  LAYER M1 ;
        RECT 3.664 8.112 3.696 10.62 ;
  LAYER M3 ;
        RECT 3.664 10.568 3.696 10.6 ;
  LAYER M1 ;
        RECT 3.728 8.112 3.76 10.62 ;
  LAYER M3 ;
        RECT 3.728 8.132 3.76 8.164 ;
  LAYER M1 ;
        RECT 3.792 8.112 3.824 10.62 ;
  LAYER M3 ;
        RECT 3.792 10.568 3.824 10.6 ;
  LAYER M1 ;
        RECT 3.856 8.112 3.888 10.62 ;
  LAYER M3 ;
        RECT 3.856 8.132 3.888 8.164 ;
  LAYER M1 ;
        RECT 3.92 8.112 3.952 10.62 ;
  LAYER M3 ;
        RECT 3.92 10.568 3.952 10.6 ;
  LAYER M1 ;
        RECT 3.984 8.112 4.016 10.62 ;
  LAYER M3 ;
        RECT 3.984 8.132 4.016 8.164 ;
  LAYER M1 ;
        RECT 4.048 8.112 4.08 10.62 ;
  LAYER M3 ;
        RECT 4.048 10.568 4.08 10.6 ;
  LAYER M1 ;
        RECT 4.112 8.112 4.144 10.62 ;
  LAYER M3 ;
        RECT 4.112 8.132 4.144 8.164 ;
  LAYER M1 ;
        RECT 4.176 8.112 4.208 10.62 ;
  LAYER M3 ;
        RECT 4.176 10.568 4.208 10.6 ;
  LAYER M1 ;
        RECT 4.24 8.112 4.272 10.62 ;
  LAYER M3 ;
        RECT 4.24 8.132 4.272 8.164 ;
  LAYER M1 ;
        RECT 4.304 8.112 4.336 10.62 ;
  LAYER M3 ;
        RECT 4.304 10.568 4.336 10.6 ;
  LAYER M1 ;
        RECT 4.368 8.112 4.4 10.62 ;
  LAYER M3 ;
        RECT 4.368 8.132 4.4 8.164 ;
  LAYER M1 ;
        RECT 4.432 8.112 4.464 10.62 ;
  LAYER M3 ;
        RECT 4.432 10.568 4.464 10.6 ;
  LAYER M1 ;
        RECT 4.496 8.112 4.528 10.62 ;
  LAYER M3 ;
        RECT 4.496 8.132 4.528 8.164 ;
  LAYER M1 ;
        RECT 4.56 8.112 4.592 10.62 ;
  LAYER M3 ;
        RECT 4.56 10.568 4.592 10.6 ;
  LAYER M1 ;
        RECT 4.624 8.112 4.656 10.62 ;
  LAYER M3 ;
        RECT 4.624 8.132 4.656 8.164 ;
  LAYER M1 ;
        RECT 4.688 8.112 4.72 10.62 ;
  LAYER M3 ;
        RECT 4.688 10.568 4.72 10.6 ;
  LAYER M1 ;
        RECT 4.752 8.112 4.784 10.62 ;
  LAYER M3 ;
        RECT 4.752 8.132 4.784 8.164 ;
  LAYER M1 ;
        RECT 4.816 8.112 4.848 10.62 ;
  LAYER M3 ;
        RECT 4.816 10.568 4.848 10.6 ;
  LAYER M1 ;
        RECT 4.88 8.112 4.912 10.62 ;
  LAYER M3 ;
        RECT 4.88 8.132 4.912 8.164 ;
  LAYER M1 ;
        RECT 4.944 8.112 4.976 10.62 ;
  LAYER M3 ;
        RECT 4.944 10.568 4.976 10.6 ;
  LAYER M1 ;
        RECT 5.008 8.112 5.04 10.62 ;
  LAYER M3 ;
        RECT 5.008 8.132 5.04 8.164 ;
  LAYER M1 ;
        RECT 5.072 8.112 5.104 10.62 ;
  LAYER M3 ;
        RECT 5.072 10.568 5.104 10.6 ;
  LAYER M1 ;
        RECT 5.136 8.112 5.168 10.62 ;
  LAYER M3 ;
        RECT 5.136 8.132 5.168 8.164 ;
  LAYER M1 ;
        RECT 5.2 8.112 5.232 10.62 ;
  LAYER M3 ;
        RECT 5.2 10.568 5.232 10.6 ;
  LAYER M1 ;
        RECT 5.264 8.112 5.296 10.62 ;
  LAYER M3 ;
        RECT 5.264 8.132 5.296 8.164 ;
  LAYER M1 ;
        RECT 5.328 8.112 5.36 10.62 ;
  LAYER M3 ;
        RECT 5.328 10.568 5.36 10.6 ;
  LAYER M1 ;
        RECT 5.392 8.112 5.424 10.62 ;
  LAYER M3 ;
        RECT 5.392 8.132 5.424 8.164 ;
  LAYER M1 ;
        RECT 5.456 8.112 5.488 10.62 ;
  LAYER M3 ;
        RECT 5.456 10.568 5.488 10.6 ;
  LAYER M1 ;
        RECT 5.52 8.112 5.552 10.62 ;
  LAYER M3 ;
        RECT 5.52 8.132 5.552 8.164 ;
  LAYER M1 ;
        RECT 5.584 8.112 5.616 10.62 ;
  LAYER M3 ;
        RECT 5.584 10.568 5.616 10.6 ;
  LAYER M1 ;
        RECT 5.648 8.112 5.68 10.62 ;
  LAYER M3 ;
        RECT 5.648 8.132 5.68 8.164 ;
  LAYER M1 ;
        RECT 5.712 8.112 5.744 10.62 ;
  LAYER M3 ;
        RECT 5.712 10.568 5.744 10.6 ;
  LAYER M1 ;
        RECT 5.776 8.112 5.808 10.62 ;
  LAYER M3 ;
        RECT 5.776 8.132 5.808 8.164 ;
  LAYER M1 ;
        RECT 5.84 8.112 5.872 10.62 ;
  LAYER M3 ;
        RECT 5.84 10.568 5.872 10.6 ;
  LAYER M1 ;
        RECT 5.904 8.112 5.936 10.62 ;
  LAYER M3 ;
        RECT 5.904 8.132 5.936 8.164 ;
  LAYER M1 ;
        RECT 5.968 8.112 6 10.62 ;
  LAYER M3 ;
        RECT 5.968 10.568 6 10.6 ;
  LAYER M1 ;
        RECT 6.032 8.112 6.064 10.62 ;
  LAYER M3 ;
        RECT 3.664 8.196 3.696 8.228 ;
  LAYER M2 ;
        RECT 6.032 8.26 6.064 8.292 ;
  LAYER M2 ;
        RECT 3.664 8.324 3.696 8.356 ;
  LAYER M2 ;
        RECT 6.032 8.388 6.064 8.42 ;
  LAYER M2 ;
        RECT 3.664 8.452 3.696 8.484 ;
  LAYER M2 ;
        RECT 6.032 8.516 6.064 8.548 ;
  LAYER M2 ;
        RECT 3.664 8.58 3.696 8.612 ;
  LAYER M2 ;
        RECT 6.032 8.644 6.064 8.676 ;
  LAYER M2 ;
        RECT 3.664 8.708 3.696 8.74 ;
  LAYER M2 ;
        RECT 6.032 8.772 6.064 8.804 ;
  LAYER M2 ;
        RECT 3.664 8.836 3.696 8.868 ;
  LAYER M2 ;
        RECT 6.032 8.9 6.064 8.932 ;
  LAYER M2 ;
        RECT 3.664 8.964 3.696 8.996 ;
  LAYER M2 ;
        RECT 6.032 9.028 6.064 9.06 ;
  LAYER M2 ;
        RECT 3.664 9.092 3.696 9.124 ;
  LAYER M2 ;
        RECT 6.032 9.156 6.064 9.188 ;
  LAYER M2 ;
        RECT 3.664 9.22 3.696 9.252 ;
  LAYER M2 ;
        RECT 6.032 9.284 6.064 9.316 ;
  LAYER M2 ;
        RECT 3.664 9.348 3.696 9.38 ;
  LAYER M2 ;
        RECT 6.032 9.412 6.064 9.444 ;
  LAYER M2 ;
        RECT 3.664 9.476 3.696 9.508 ;
  LAYER M2 ;
        RECT 6.032 9.54 6.064 9.572 ;
  LAYER M2 ;
        RECT 3.664 9.604 3.696 9.636 ;
  LAYER M2 ;
        RECT 6.032 9.668 6.064 9.7 ;
  LAYER M2 ;
        RECT 3.664 9.732 3.696 9.764 ;
  LAYER M2 ;
        RECT 6.032 9.796 6.064 9.828 ;
  LAYER M2 ;
        RECT 3.664 9.86 3.696 9.892 ;
  LAYER M2 ;
        RECT 6.032 9.924 6.064 9.956 ;
  LAYER M2 ;
        RECT 3.664 9.988 3.696 10.02 ;
  LAYER M2 ;
        RECT 6.032 10.052 6.064 10.084 ;
  LAYER M2 ;
        RECT 3.664 10.116 3.696 10.148 ;
  LAYER M2 ;
        RECT 6.032 10.18 6.064 10.212 ;
  LAYER M2 ;
        RECT 3.664 10.244 3.696 10.276 ;
  LAYER M2 ;
        RECT 6.032 10.308 6.064 10.34 ;
  LAYER M2 ;
        RECT 3.664 10.372 3.696 10.404 ;
  LAYER M2 ;
        RECT 6.032 10.436 6.064 10.468 ;
  LAYER M2 ;
        RECT 3.616 8.064 6.112 10.668 ;
  LAYER M1 ;
        RECT 3.664 11.22 3.696 13.728 ;
  LAYER M3 ;
        RECT 3.664 13.676 3.696 13.708 ;
  LAYER M1 ;
        RECT 3.728 11.22 3.76 13.728 ;
  LAYER M3 ;
        RECT 3.728 11.24 3.76 11.272 ;
  LAYER M1 ;
        RECT 3.792 11.22 3.824 13.728 ;
  LAYER M3 ;
        RECT 3.792 13.676 3.824 13.708 ;
  LAYER M1 ;
        RECT 3.856 11.22 3.888 13.728 ;
  LAYER M3 ;
        RECT 3.856 11.24 3.888 11.272 ;
  LAYER M1 ;
        RECT 3.92 11.22 3.952 13.728 ;
  LAYER M3 ;
        RECT 3.92 13.676 3.952 13.708 ;
  LAYER M1 ;
        RECT 3.984 11.22 4.016 13.728 ;
  LAYER M3 ;
        RECT 3.984 11.24 4.016 11.272 ;
  LAYER M1 ;
        RECT 4.048 11.22 4.08 13.728 ;
  LAYER M3 ;
        RECT 4.048 13.676 4.08 13.708 ;
  LAYER M1 ;
        RECT 4.112 11.22 4.144 13.728 ;
  LAYER M3 ;
        RECT 4.112 11.24 4.144 11.272 ;
  LAYER M1 ;
        RECT 4.176 11.22 4.208 13.728 ;
  LAYER M3 ;
        RECT 4.176 13.676 4.208 13.708 ;
  LAYER M1 ;
        RECT 4.24 11.22 4.272 13.728 ;
  LAYER M3 ;
        RECT 4.24 11.24 4.272 11.272 ;
  LAYER M1 ;
        RECT 4.304 11.22 4.336 13.728 ;
  LAYER M3 ;
        RECT 4.304 13.676 4.336 13.708 ;
  LAYER M1 ;
        RECT 4.368 11.22 4.4 13.728 ;
  LAYER M3 ;
        RECT 4.368 11.24 4.4 11.272 ;
  LAYER M1 ;
        RECT 4.432 11.22 4.464 13.728 ;
  LAYER M3 ;
        RECT 4.432 13.676 4.464 13.708 ;
  LAYER M1 ;
        RECT 4.496 11.22 4.528 13.728 ;
  LAYER M3 ;
        RECT 4.496 11.24 4.528 11.272 ;
  LAYER M1 ;
        RECT 4.56 11.22 4.592 13.728 ;
  LAYER M3 ;
        RECT 4.56 13.676 4.592 13.708 ;
  LAYER M1 ;
        RECT 4.624 11.22 4.656 13.728 ;
  LAYER M3 ;
        RECT 4.624 11.24 4.656 11.272 ;
  LAYER M1 ;
        RECT 4.688 11.22 4.72 13.728 ;
  LAYER M3 ;
        RECT 4.688 13.676 4.72 13.708 ;
  LAYER M1 ;
        RECT 4.752 11.22 4.784 13.728 ;
  LAYER M3 ;
        RECT 4.752 11.24 4.784 11.272 ;
  LAYER M1 ;
        RECT 4.816 11.22 4.848 13.728 ;
  LAYER M3 ;
        RECT 4.816 13.676 4.848 13.708 ;
  LAYER M1 ;
        RECT 4.88 11.22 4.912 13.728 ;
  LAYER M3 ;
        RECT 4.88 11.24 4.912 11.272 ;
  LAYER M1 ;
        RECT 4.944 11.22 4.976 13.728 ;
  LAYER M3 ;
        RECT 4.944 13.676 4.976 13.708 ;
  LAYER M1 ;
        RECT 5.008 11.22 5.04 13.728 ;
  LAYER M3 ;
        RECT 5.008 11.24 5.04 11.272 ;
  LAYER M1 ;
        RECT 5.072 11.22 5.104 13.728 ;
  LAYER M3 ;
        RECT 5.072 13.676 5.104 13.708 ;
  LAYER M1 ;
        RECT 5.136 11.22 5.168 13.728 ;
  LAYER M3 ;
        RECT 5.136 11.24 5.168 11.272 ;
  LAYER M1 ;
        RECT 5.2 11.22 5.232 13.728 ;
  LAYER M3 ;
        RECT 5.2 13.676 5.232 13.708 ;
  LAYER M1 ;
        RECT 5.264 11.22 5.296 13.728 ;
  LAYER M3 ;
        RECT 5.264 11.24 5.296 11.272 ;
  LAYER M1 ;
        RECT 5.328 11.22 5.36 13.728 ;
  LAYER M3 ;
        RECT 5.328 13.676 5.36 13.708 ;
  LAYER M1 ;
        RECT 5.392 11.22 5.424 13.728 ;
  LAYER M3 ;
        RECT 5.392 11.24 5.424 11.272 ;
  LAYER M1 ;
        RECT 5.456 11.22 5.488 13.728 ;
  LAYER M3 ;
        RECT 5.456 13.676 5.488 13.708 ;
  LAYER M1 ;
        RECT 5.52 11.22 5.552 13.728 ;
  LAYER M3 ;
        RECT 5.52 11.24 5.552 11.272 ;
  LAYER M1 ;
        RECT 5.584 11.22 5.616 13.728 ;
  LAYER M3 ;
        RECT 5.584 13.676 5.616 13.708 ;
  LAYER M1 ;
        RECT 5.648 11.22 5.68 13.728 ;
  LAYER M3 ;
        RECT 5.648 11.24 5.68 11.272 ;
  LAYER M1 ;
        RECT 5.712 11.22 5.744 13.728 ;
  LAYER M3 ;
        RECT 5.712 13.676 5.744 13.708 ;
  LAYER M1 ;
        RECT 5.776 11.22 5.808 13.728 ;
  LAYER M3 ;
        RECT 5.776 11.24 5.808 11.272 ;
  LAYER M1 ;
        RECT 5.84 11.22 5.872 13.728 ;
  LAYER M3 ;
        RECT 5.84 13.676 5.872 13.708 ;
  LAYER M1 ;
        RECT 5.904 11.22 5.936 13.728 ;
  LAYER M3 ;
        RECT 5.904 11.24 5.936 11.272 ;
  LAYER M1 ;
        RECT 5.968 11.22 6 13.728 ;
  LAYER M3 ;
        RECT 5.968 13.676 6 13.708 ;
  LAYER M1 ;
        RECT 6.032 11.22 6.064 13.728 ;
  LAYER M3 ;
        RECT 3.664 11.304 3.696 11.336 ;
  LAYER M2 ;
        RECT 6.032 11.368 6.064 11.4 ;
  LAYER M2 ;
        RECT 3.664 11.432 3.696 11.464 ;
  LAYER M2 ;
        RECT 6.032 11.496 6.064 11.528 ;
  LAYER M2 ;
        RECT 3.664 11.56 3.696 11.592 ;
  LAYER M2 ;
        RECT 6.032 11.624 6.064 11.656 ;
  LAYER M2 ;
        RECT 3.664 11.688 3.696 11.72 ;
  LAYER M2 ;
        RECT 6.032 11.752 6.064 11.784 ;
  LAYER M2 ;
        RECT 3.664 11.816 3.696 11.848 ;
  LAYER M2 ;
        RECT 6.032 11.88 6.064 11.912 ;
  LAYER M2 ;
        RECT 3.664 11.944 3.696 11.976 ;
  LAYER M2 ;
        RECT 6.032 12.008 6.064 12.04 ;
  LAYER M2 ;
        RECT 3.664 12.072 3.696 12.104 ;
  LAYER M2 ;
        RECT 6.032 12.136 6.064 12.168 ;
  LAYER M2 ;
        RECT 3.664 12.2 3.696 12.232 ;
  LAYER M2 ;
        RECT 6.032 12.264 6.064 12.296 ;
  LAYER M2 ;
        RECT 3.664 12.328 3.696 12.36 ;
  LAYER M2 ;
        RECT 6.032 12.392 6.064 12.424 ;
  LAYER M2 ;
        RECT 3.664 12.456 3.696 12.488 ;
  LAYER M2 ;
        RECT 6.032 12.52 6.064 12.552 ;
  LAYER M2 ;
        RECT 3.664 12.584 3.696 12.616 ;
  LAYER M2 ;
        RECT 6.032 12.648 6.064 12.68 ;
  LAYER M2 ;
        RECT 3.664 12.712 3.696 12.744 ;
  LAYER M2 ;
        RECT 6.032 12.776 6.064 12.808 ;
  LAYER M2 ;
        RECT 3.664 12.84 3.696 12.872 ;
  LAYER M2 ;
        RECT 6.032 12.904 6.064 12.936 ;
  LAYER M2 ;
        RECT 3.664 12.968 3.696 13 ;
  LAYER M2 ;
        RECT 6.032 13.032 6.064 13.064 ;
  LAYER M2 ;
        RECT 3.664 13.096 3.696 13.128 ;
  LAYER M2 ;
        RECT 6.032 13.16 6.064 13.192 ;
  LAYER M2 ;
        RECT 3.664 13.224 3.696 13.256 ;
  LAYER M2 ;
        RECT 6.032 13.288 6.064 13.32 ;
  LAYER M2 ;
        RECT 3.664 13.352 3.696 13.384 ;
  LAYER M2 ;
        RECT 6.032 13.416 6.064 13.448 ;
  LAYER M2 ;
        RECT 3.664 13.48 3.696 13.512 ;
  LAYER M2 ;
        RECT 6.032 13.544 6.064 13.576 ;
  LAYER M2 ;
        RECT 3.616 11.172 6.112 13.776 ;
  LAYER M1 ;
        RECT 6.64 1.896 6.672 4.404 ;
  LAYER M3 ;
        RECT 6.64 4.352 6.672 4.384 ;
  LAYER M1 ;
        RECT 6.704 1.896 6.736 4.404 ;
  LAYER M3 ;
        RECT 6.704 1.916 6.736 1.948 ;
  LAYER M1 ;
        RECT 6.768 1.896 6.8 4.404 ;
  LAYER M3 ;
        RECT 6.768 4.352 6.8 4.384 ;
  LAYER M1 ;
        RECT 6.832 1.896 6.864 4.404 ;
  LAYER M3 ;
        RECT 6.832 1.916 6.864 1.948 ;
  LAYER M1 ;
        RECT 6.896 1.896 6.928 4.404 ;
  LAYER M3 ;
        RECT 6.896 4.352 6.928 4.384 ;
  LAYER M1 ;
        RECT 6.96 1.896 6.992 4.404 ;
  LAYER M3 ;
        RECT 6.96 1.916 6.992 1.948 ;
  LAYER M1 ;
        RECT 7.024 1.896 7.056 4.404 ;
  LAYER M3 ;
        RECT 7.024 4.352 7.056 4.384 ;
  LAYER M1 ;
        RECT 7.088 1.896 7.12 4.404 ;
  LAYER M3 ;
        RECT 7.088 1.916 7.12 1.948 ;
  LAYER M1 ;
        RECT 7.152 1.896 7.184 4.404 ;
  LAYER M3 ;
        RECT 7.152 4.352 7.184 4.384 ;
  LAYER M1 ;
        RECT 7.216 1.896 7.248 4.404 ;
  LAYER M3 ;
        RECT 7.216 1.916 7.248 1.948 ;
  LAYER M1 ;
        RECT 7.28 1.896 7.312 4.404 ;
  LAYER M3 ;
        RECT 7.28 4.352 7.312 4.384 ;
  LAYER M1 ;
        RECT 7.344 1.896 7.376 4.404 ;
  LAYER M3 ;
        RECT 7.344 1.916 7.376 1.948 ;
  LAYER M1 ;
        RECT 7.408 1.896 7.44 4.404 ;
  LAYER M3 ;
        RECT 7.408 4.352 7.44 4.384 ;
  LAYER M1 ;
        RECT 7.472 1.896 7.504 4.404 ;
  LAYER M3 ;
        RECT 7.472 1.916 7.504 1.948 ;
  LAYER M1 ;
        RECT 7.536 1.896 7.568 4.404 ;
  LAYER M3 ;
        RECT 7.536 4.352 7.568 4.384 ;
  LAYER M1 ;
        RECT 7.6 1.896 7.632 4.404 ;
  LAYER M3 ;
        RECT 7.6 1.916 7.632 1.948 ;
  LAYER M1 ;
        RECT 7.664 1.896 7.696 4.404 ;
  LAYER M3 ;
        RECT 7.664 4.352 7.696 4.384 ;
  LAYER M1 ;
        RECT 7.728 1.896 7.76 4.404 ;
  LAYER M3 ;
        RECT 7.728 1.916 7.76 1.948 ;
  LAYER M1 ;
        RECT 7.792 1.896 7.824 4.404 ;
  LAYER M3 ;
        RECT 7.792 4.352 7.824 4.384 ;
  LAYER M1 ;
        RECT 7.856 1.896 7.888 4.404 ;
  LAYER M3 ;
        RECT 7.856 1.916 7.888 1.948 ;
  LAYER M1 ;
        RECT 7.92 1.896 7.952 4.404 ;
  LAYER M3 ;
        RECT 7.92 4.352 7.952 4.384 ;
  LAYER M1 ;
        RECT 7.984 1.896 8.016 4.404 ;
  LAYER M3 ;
        RECT 7.984 1.916 8.016 1.948 ;
  LAYER M1 ;
        RECT 8.048 1.896 8.08 4.404 ;
  LAYER M3 ;
        RECT 8.048 4.352 8.08 4.384 ;
  LAYER M1 ;
        RECT 8.112 1.896 8.144 4.404 ;
  LAYER M3 ;
        RECT 8.112 1.916 8.144 1.948 ;
  LAYER M1 ;
        RECT 8.176 1.896 8.208 4.404 ;
  LAYER M3 ;
        RECT 8.176 4.352 8.208 4.384 ;
  LAYER M1 ;
        RECT 8.24 1.896 8.272 4.404 ;
  LAYER M3 ;
        RECT 8.24 1.916 8.272 1.948 ;
  LAYER M1 ;
        RECT 8.304 1.896 8.336 4.404 ;
  LAYER M3 ;
        RECT 8.304 4.352 8.336 4.384 ;
  LAYER M1 ;
        RECT 8.368 1.896 8.4 4.404 ;
  LAYER M3 ;
        RECT 8.368 1.916 8.4 1.948 ;
  LAYER M1 ;
        RECT 8.432 1.896 8.464 4.404 ;
  LAYER M3 ;
        RECT 8.432 4.352 8.464 4.384 ;
  LAYER M1 ;
        RECT 8.496 1.896 8.528 4.404 ;
  LAYER M3 ;
        RECT 8.496 1.916 8.528 1.948 ;
  LAYER M1 ;
        RECT 8.56 1.896 8.592 4.404 ;
  LAYER M3 ;
        RECT 8.56 4.352 8.592 4.384 ;
  LAYER M1 ;
        RECT 8.624 1.896 8.656 4.404 ;
  LAYER M3 ;
        RECT 8.624 1.916 8.656 1.948 ;
  LAYER M1 ;
        RECT 8.688 1.896 8.72 4.404 ;
  LAYER M3 ;
        RECT 8.688 4.352 8.72 4.384 ;
  LAYER M1 ;
        RECT 8.752 1.896 8.784 4.404 ;
  LAYER M3 ;
        RECT 8.752 1.916 8.784 1.948 ;
  LAYER M1 ;
        RECT 8.816 1.896 8.848 4.404 ;
  LAYER M3 ;
        RECT 8.816 4.352 8.848 4.384 ;
  LAYER M1 ;
        RECT 8.88 1.896 8.912 4.404 ;
  LAYER M3 ;
        RECT 8.88 1.916 8.912 1.948 ;
  LAYER M1 ;
        RECT 8.944 1.896 8.976 4.404 ;
  LAYER M3 ;
        RECT 8.944 4.352 8.976 4.384 ;
  LAYER M1 ;
        RECT 9.008 1.896 9.04 4.404 ;
  LAYER M3 ;
        RECT 6.64 1.98 6.672 2.012 ;
  LAYER M2 ;
        RECT 9.008 2.044 9.04 2.076 ;
  LAYER M2 ;
        RECT 6.64 2.108 6.672 2.14 ;
  LAYER M2 ;
        RECT 9.008 2.172 9.04 2.204 ;
  LAYER M2 ;
        RECT 6.64 2.236 6.672 2.268 ;
  LAYER M2 ;
        RECT 9.008 2.3 9.04 2.332 ;
  LAYER M2 ;
        RECT 6.64 2.364 6.672 2.396 ;
  LAYER M2 ;
        RECT 9.008 2.428 9.04 2.46 ;
  LAYER M2 ;
        RECT 6.64 2.492 6.672 2.524 ;
  LAYER M2 ;
        RECT 9.008 2.556 9.04 2.588 ;
  LAYER M2 ;
        RECT 6.64 2.62 6.672 2.652 ;
  LAYER M2 ;
        RECT 9.008 2.684 9.04 2.716 ;
  LAYER M2 ;
        RECT 6.64 2.748 6.672 2.78 ;
  LAYER M2 ;
        RECT 9.008 2.812 9.04 2.844 ;
  LAYER M2 ;
        RECT 6.64 2.876 6.672 2.908 ;
  LAYER M2 ;
        RECT 9.008 2.94 9.04 2.972 ;
  LAYER M2 ;
        RECT 6.64 3.004 6.672 3.036 ;
  LAYER M2 ;
        RECT 9.008 3.068 9.04 3.1 ;
  LAYER M2 ;
        RECT 6.64 3.132 6.672 3.164 ;
  LAYER M2 ;
        RECT 9.008 3.196 9.04 3.228 ;
  LAYER M2 ;
        RECT 6.64 3.26 6.672 3.292 ;
  LAYER M2 ;
        RECT 9.008 3.324 9.04 3.356 ;
  LAYER M2 ;
        RECT 6.64 3.388 6.672 3.42 ;
  LAYER M2 ;
        RECT 9.008 3.452 9.04 3.484 ;
  LAYER M2 ;
        RECT 6.64 3.516 6.672 3.548 ;
  LAYER M2 ;
        RECT 9.008 3.58 9.04 3.612 ;
  LAYER M2 ;
        RECT 6.64 3.644 6.672 3.676 ;
  LAYER M2 ;
        RECT 9.008 3.708 9.04 3.74 ;
  LAYER M2 ;
        RECT 6.64 3.772 6.672 3.804 ;
  LAYER M2 ;
        RECT 9.008 3.836 9.04 3.868 ;
  LAYER M2 ;
        RECT 6.64 3.9 6.672 3.932 ;
  LAYER M2 ;
        RECT 9.008 3.964 9.04 3.996 ;
  LAYER M2 ;
        RECT 6.64 4.028 6.672 4.06 ;
  LAYER M2 ;
        RECT 9.008 4.092 9.04 4.124 ;
  LAYER M2 ;
        RECT 6.64 4.156 6.672 4.188 ;
  LAYER M2 ;
        RECT 9.008 4.22 9.04 4.252 ;
  LAYER M2 ;
        RECT 6.592 1.848 9.088 4.452 ;
  LAYER M1 ;
        RECT 6.64 5.004 6.672 7.512 ;
  LAYER M3 ;
        RECT 6.64 7.46 6.672 7.492 ;
  LAYER M1 ;
        RECT 6.704 5.004 6.736 7.512 ;
  LAYER M3 ;
        RECT 6.704 5.024 6.736 5.056 ;
  LAYER M1 ;
        RECT 6.768 5.004 6.8 7.512 ;
  LAYER M3 ;
        RECT 6.768 7.46 6.8 7.492 ;
  LAYER M1 ;
        RECT 6.832 5.004 6.864 7.512 ;
  LAYER M3 ;
        RECT 6.832 5.024 6.864 5.056 ;
  LAYER M1 ;
        RECT 6.896 5.004 6.928 7.512 ;
  LAYER M3 ;
        RECT 6.896 7.46 6.928 7.492 ;
  LAYER M1 ;
        RECT 6.96 5.004 6.992 7.512 ;
  LAYER M3 ;
        RECT 6.96 5.024 6.992 5.056 ;
  LAYER M1 ;
        RECT 7.024 5.004 7.056 7.512 ;
  LAYER M3 ;
        RECT 7.024 7.46 7.056 7.492 ;
  LAYER M1 ;
        RECT 7.088 5.004 7.12 7.512 ;
  LAYER M3 ;
        RECT 7.088 5.024 7.12 5.056 ;
  LAYER M1 ;
        RECT 7.152 5.004 7.184 7.512 ;
  LAYER M3 ;
        RECT 7.152 7.46 7.184 7.492 ;
  LAYER M1 ;
        RECT 7.216 5.004 7.248 7.512 ;
  LAYER M3 ;
        RECT 7.216 5.024 7.248 5.056 ;
  LAYER M1 ;
        RECT 7.28 5.004 7.312 7.512 ;
  LAYER M3 ;
        RECT 7.28 7.46 7.312 7.492 ;
  LAYER M1 ;
        RECT 7.344 5.004 7.376 7.512 ;
  LAYER M3 ;
        RECT 7.344 5.024 7.376 5.056 ;
  LAYER M1 ;
        RECT 7.408 5.004 7.44 7.512 ;
  LAYER M3 ;
        RECT 7.408 7.46 7.44 7.492 ;
  LAYER M1 ;
        RECT 7.472 5.004 7.504 7.512 ;
  LAYER M3 ;
        RECT 7.472 5.024 7.504 5.056 ;
  LAYER M1 ;
        RECT 7.536 5.004 7.568 7.512 ;
  LAYER M3 ;
        RECT 7.536 7.46 7.568 7.492 ;
  LAYER M1 ;
        RECT 7.6 5.004 7.632 7.512 ;
  LAYER M3 ;
        RECT 7.6 5.024 7.632 5.056 ;
  LAYER M1 ;
        RECT 7.664 5.004 7.696 7.512 ;
  LAYER M3 ;
        RECT 7.664 7.46 7.696 7.492 ;
  LAYER M1 ;
        RECT 7.728 5.004 7.76 7.512 ;
  LAYER M3 ;
        RECT 7.728 5.024 7.76 5.056 ;
  LAYER M1 ;
        RECT 7.792 5.004 7.824 7.512 ;
  LAYER M3 ;
        RECT 7.792 7.46 7.824 7.492 ;
  LAYER M1 ;
        RECT 7.856 5.004 7.888 7.512 ;
  LAYER M3 ;
        RECT 7.856 5.024 7.888 5.056 ;
  LAYER M1 ;
        RECT 7.92 5.004 7.952 7.512 ;
  LAYER M3 ;
        RECT 7.92 7.46 7.952 7.492 ;
  LAYER M1 ;
        RECT 7.984 5.004 8.016 7.512 ;
  LAYER M3 ;
        RECT 7.984 5.024 8.016 5.056 ;
  LAYER M1 ;
        RECT 8.048 5.004 8.08 7.512 ;
  LAYER M3 ;
        RECT 8.048 7.46 8.08 7.492 ;
  LAYER M1 ;
        RECT 8.112 5.004 8.144 7.512 ;
  LAYER M3 ;
        RECT 8.112 5.024 8.144 5.056 ;
  LAYER M1 ;
        RECT 8.176 5.004 8.208 7.512 ;
  LAYER M3 ;
        RECT 8.176 7.46 8.208 7.492 ;
  LAYER M1 ;
        RECT 8.24 5.004 8.272 7.512 ;
  LAYER M3 ;
        RECT 8.24 5.024 8.272 5.056 ;
  LAYER M1 ;
        RECT 8.304 5.004 8.336 7.512 ;
  LAYER M3 ;
        RECT 8.304 7.46 8.336 7.492 ;
  LAYER M1 ;
        RECT 8.368 5.004 8.4 7.512 ;
  LAYER M3 ;
        RECT 8.368 5.024 8.4 5.056 ;
  LAYER M1 ;
        RECT 8.432 5.004 8.464 7.512 ;
  LAYER M3 ;
        RECT 8.432 7.46 8.464 7.492 ;
  LAYER M1 ;
        RECT 8.496 5.004 8.528 7.512 ;
  LAYER M3 ;
        RECT 8.496 5.024 8.528 5.056 ;
  LAYER M1 ;
        RECT 8.56 5.004 8.592 7.512 ;
  LAYER M3 ;
        RECT 8.56 7.46 8.592 7.492 ;
  LAYER M1 ;
        RECT 8.624 5.004 8.656 7.512 ;
  LAYER M3 ;
        RECT 8.624 5.024 8.656 5.056 ;
  LAYER M1 ;
        RECT 8.688 5.004 8.72 7.512 ;
  LAYER M3 ;
        RECT 8.688 7.46 8.72 7.492 ;
  LAYER M1 ;
        RECT 8.752 5.004 8.784 7.512 ;
  LAYER M3 ;
        RECT 8.752 5.024 8.784 5.056 ;
  LAYER M1 ;
        RECT 8.816 5.004 8.848 7.512 ;
  LAYER M3 ;
        RECT 8.816 7.46 8.848 7.492 ;
  LAYER M1 ;
        RECT 8.88 5.004 8.912 7.512 ;
  LAYER M3 ;
        RECT 8.88 5.024 8.912 5.056 ;
  LAYER M1 ;
        RECT 8.944 5.004 8.976 7.512 ;
  LAYER M3 ;
        RECT 8.944 7.46 8.976 7.492 ;
  LAYER M1 ;
        RECT 9.008 5.004 9.04 7.512 ;
  LAYER M3 ;
        RECT 6.64 5.088 6.672 5.12 ;
  LAYER M2 ;
        RECT 9.008 5.152 9.04 5.184 ;
  LAYER M2 ;
        RECT 6.64 5.216 6.672 5.248 ;
  LAYER M2 ;
        RECT 9.008 5.28 9.04 5.312 ;
  LAYER M2 ;
        RECT 6.64 5.344 6.672 5.376 ;
  LAYER M2 ;
        RECT 9.008 5.408 9.04 5.44 ;
  LAYER M2 ;
        RECT 6.64 5.472 6.672 5.504 ;
  LAYER M2 ;
        RECT 9.008 5.536 9.04 5.568 ;
  LAYER M2 ;
        RECT 6.64 5.6 6.672 5.632 ;
  LAYER M2 ;
        RECT 9.008 5.664 9.04 5.696 ;
  LAYER M2 ;
        RECT 6.64 5.728 6.672 5.76 ;
  LAYER M2 ;
        RECT 9.008 5.792 9.04 5.824 ;
  LAYER M2 ;
        RECT 6.64 5.856 6.672 5.888 ;
  LAYER M2 ;
        RECT 9.008 5.92 9.04 5.952 ;
  LAYER M2 ;
        RECT 6.64 5.984 6.672 6.016 ;
  LAYER M2 ;
        RECT 9.008 6.048 9.04 6.08 ;
  LAYER M2 ;
        RECT 6.64 6.112 6.672 6.144 ;
  LAYER M2 ;
        RECT 9.008 6.176 9.04 6.208 ;
  LAYER M2 ;
        RECT 6.64 6.24 6.672 6.272 ;
  LAYER M2 ;
        RECT 9.008 6.304 9.04 6.336 ;
  LAYER M2 ;
        RECT 6.64 6.368 6.672 6.4 ;
  LAYER M2 ;
        RECT 9.008 6.432 9.04 6.464 ;
  LAYER M2 ;
        RECT 6.64 6.496 6.672 6.528 ;
  LAYER M2 ;
        RECT 9.008 6.56 9.04 6.592 ;
  LAYER M2 ;
        RECT 6.64 6.624 6.672 6.656 ;
  LAYER M2 ;
        RECT 9.008 6.688 9.04 6.72 ;
  LAYER M2 ;
        RECT 6.64 6.752 6.672 6.784 ;
  LAYER M2 ;
        RECT 9.008 6.816 9.04 6.848 ;
  LAYER M2 ;
        RECT 6.64 6.88 6.672 6.912 ;
  LAYER M2 ;
        RECT 9.008 6.944 9.04 6.976 ;
  LAYER M2 ;
        RECT 6.64 7.008 6.672 7.04 ;
  LAYER M2 ;
        RECT 9.008 7.072 9.04 7.104 ;
  LAYER M2 ;
        RECT 6.64 7.136 6.672 7.168 ;
  LAYER M2 ;
        RECT 9.008 7.2 9.04 7.232 ;
  LAYER M2 ;
        RECT 6.64 7.264 6.672 7.296 ;
  LAYER M2 ;
        RECT 9.008 7.328 9.04 7.36 ;
  LAYER M2 ;
        RECT 6.592 4.956 9.088 7.56 ;
  LAYER M1 ;
        RECT 6.64 8.112 6.672 10.62 ;
  LAYER M3 ;
        RECT 6.64 10.568 6.672 10.6 ;
  LAYER M1 ;
        RECT 6.704 8.112 6.736 10.62 ;
  LAYER M3 ;
        RECT 6.704 8.132 6.736 8.164 ;
  LAYER M1 ;
        RECT 6.768 8.112 6.8 10.62 ;
  LAYER M3 ;
        RECT 6.768 10.568 6.8 10.6 ;
  LAYER M1 ;
        RECT 6.832 8.112 6.864 10.62 ;
  LAYER M3 ;
        RECT 6.832 8.132 6.864 8.164 ;
  LAYER M1 ;
        RECT 6.896 8.112 6.928 10.62 ;
  LAYER M3 ;
        RECT 6.896 10.568 6.928 10.6 ;
  LAYER M1 ;
        RECT 6.96 8.112 6.992 10.62 ;
  LAYER M3 ;
        RECT 6.96 8.132 6.992 8.164 ;
  LAYER M1 ;
        RECT 7.024 8.112 7.056 10.62 ;
  LAYER M3 ;
        RECT 7.024 10.568 7.056 10.6 ;
  LAYER M1 ;
        RECT 7.088 8.112 7.12 10.62 ;
  LAYER M3 ;
        RECT 7.088 8.132 7.12 8.164 ;
  LAYER M1 ;
        RECT 7.152 8.112 7.184 10.62 ;
  LAYER M3 ;
        RECT 7.152 10.568 7.184 10.6 ;
  LAYER M1 ;
        RECT 7.216 8.112 7.248 10.62 ;
  LAYER M3 ;
        RECT 7.216 8.132 7.248 8.164 ;
  LAYER M1 ;
        RECT 7.28 8.112 7.312 10.62 ;
  LAYER M3 ;
        RECT 7.28 10.568 7.312 10.6 ;
  LAYER M1 ;
        RECT 7.344 8.112 7.376 10.62 ;
  LAYER M3 ;
        RECT 7.344 8.132 7.376 8.164 ;
  LAYER M1 ;
        RECT 7.408 8.112 7.44 10.62 ;
  LAYER M3 ;
        RECT 7.408 10.568 7.44 10.6 ;
  LAYER M1 ;
        RECT 7.472 8.112 7.504 10.62 ;
  LAYER M3 ;
        RECT 7.472 8.132 7.504 8.164 ;
  LAYER M1 ;
        RECT 7.536 8.112 7.568 10.62 ;
  LAYER M3 ;
        RECT 7.536 10.568 7.568 10.6 ;
  LAYER M1 ;
        RECT 7.6 8.112 7.632 10.62 ;
  LAYER M3 ;
        RECT 7.6 8.132 7.632 8.164 ;
  LAYER M1 ;
        RECT 7.664 8.112 7.696 10.62 ;
  LAYER M3 ;
        RECT 7.664 10.568 7.696 10.6 ;
  LAYER M1 ;
        RECT 7.728 8.112 7.76 10.62 ;
  LAYER M3 ;
        RECT 7.728 8.132 7.76 8.164 ;
  LAYER M1 ;
        RECT 7.792 8.112 7.824 10.62 ;
  LAYER M3 ;
        RECT 7.792 10.568 7.824 10.6 ;
  LAYER M1 ;
        RECT 7.856 8.112 7.888 10.62 ;
  LAYER M3 ;
        RECT 7.856 8.132 7.888 8.164 ;
  LAYER M1 ;
        RECT 7.92 8.112 7.952 10.62 ;
  LAYER M3 ;
        RECT 7.92 10.568 7.952 10.6 ;
  LAYER M1 ;
        RECT 7.984 8.112 8.016 10.62 ;
  LAYER M3 ;
        RECT 7.984 8.132 8.016 8.164 ;
  LAYER M1 ;
        RECT 8.048 8.112 8.08 10.62 ;
  LAYER M3 ;
        RECT 8.048 10.568 8.08 10.6 ;
  LAYER M1 ;
        RECT 8.112 8.112 8.144 10.62 ;
  LAYER M3 ;
        RECT 8.112 8.132 8.144 8.164 ;
  LAYER M1 ;
        RECT 8.176 8.112 8.208 10.62 ;
  LAYER M3 ;
        RECT 8.176 10.568 8.208 10.6 ;
  LAYER M1 ;
        RECT 8.24 8.112 8.272 10.62 ;
  LAYER M3 ;
        RECT 8.24 8.132 8.272 8.164 ;
  LAYER M1 ;
        RECT 8.304 8.112 8.336 10.62 ;
  LAYER M3 ;
        RECT 8.304 10.568 8.336 10.6 ;
  LAYER M1 ;
        RECT 8.368 8.112 8.4 10.62 ;
  LAYER M3 ;
        RECT 8.368 8.132 8.4 8.164 ;
  LAYER M1 ;
        RECT 8.432 8.112 8.464 10.62 ;
  LAYER M3 ;
        RECT 8.432 10.568 8.464 10.6 ;
  LAYER M1 ;
        RECT 8.496 8.112 8.528 10.62 ;
  LAYER M3 ;
        RECT 8.496 8.132 8.528 8.164 ;
  LAYER M1 ;
        RECT 8.56 8.112 8.592 10.62 ;
  LAYER M3 ;
        RECT 8.56 10.568 8.592 10.6 ;
  LAYER M1 ;
        RECT 8.624 8.112 8.656 10.62 ;
  LAYER M3 ;
        RECT 8.624 8.132 8.656 8.164 ;
  LAYER M1 ;
        RECT 8.688 8.112 8.72 10.62 ;
  LAYER M3 ;
        RECT 8.688 10.568 8.72 10.6 ;
  LAYER M1 ;
        RECT 8.752 8.112 8.784 10.62 ;
  LAYER M3 ;
        RECT 8.752 8.132 8.784 8.164 ;
  LAYER M1 ;
        RECT 8.816 8.112 8.848 10.62 ;
  LAYER M3 ;
        RECT 8.816 10.568 8.848 10.6 ;
  LAYER M1 ;
        RECT 8.88 8.112 8.912 10.62 ;
  LAYER M3 ;
        RECT 8.88 8.132 8.912 8.164 ;
  LAYER M1 ;
        RECT 8.944 8.112 8.976 10.62 ;
  LAYER M3 ;
        RECT 8.944 10.568 8.976 10.6 ;
  LAYER M1 ;
        RECT 9.008 8.112 9.04 10.62 ;
  LAYER M3 ;
        RECT 6.64 8.196 6.672 8.228 ;
  LAYER M2 ;
        RECT 9.008 8.26 9.04 8.292 ;
  LAYER M2 ;
        RECT 6.64 8.324 6.672 8.356 ;
  LAYER M2 ;
        RECT 9.008 8.388 9.04 8.42 ;
  LAYER M2 ;
        RECT 6.64 8.452 6.672 8.484 ;
  LAYER M2 ;
        RECT 9.008 8.516 9.04 8.548 ;
  LAYER M2 ;
        RECT 6.64 8.58 6.672 8.612 ;
  LAYER M2 ;
        RECT 9.008 8.644 9.04 8.676 ;
  LAYER M2 ;
        RECT 6.64 8.708 6.672 8.74 ;
  LAYER M2 ;
        RECT 9.008 8.772 9.04 8.804 ;
  LAYER M2 ;
        RECT 6.64 8.836 6.672 8.868 ;
  LAYER M2 ;
        RECT 9.008 8.9 9.04 8.932 ;
  LAYER M2 ;
        RECT 6.64 8.964 6.672 8.996 ;
  LAYER M2 ;
        RECT 9.008 9.028 9.04 9.06 ;
  LAYER M2 ;
        RECT 6.64 9.092 6.672 9.124 ;
  LAYER M2 ;
        RECT 9.008 9.156 9.04 9.188 ;
  LAYER M2 ;
        RECT 6.64 9.22 6.672 9.252 ;
  LAYER M2 ;
        RECT 9.008 9.284 9.04 9.316 ;
  LAYER M2 ;
        RECT 6.64 9.348 6.672 9.38 ;
  LAYER M2 ;
        RECT 9.008 9.412 9.04 9.444 ;
  LAYER M2 ;
        RECT 6.64 9.476 6.672 9.508 ;
  LAYER M2 ;
        RECT 9.008 9.54 9.04 9.572 ;
  LAYER M2 ;
        RECT 6.64 9.604 6.672 9.636 ;
  LAYER M2 ;
        RECT 9.008 9.668 9.04 9.7 ;
  LAYER M2 ;
        RECT 6.64 9.732 6.672 9.764 ;
  LAYER M2 ;
        RECT 9.008 9.796 9.04 9.828 ;
  LAYER M2 ;
        RECT 6.64 9.86 6.672 9.892 ;
  LAYER M2 ;
        RECT 9.008 9.924 9.04 9.956 ;
  LAYER M2 ;
        RECT 6.64 9.988 6.672 10.02 ;
  LAYER M2 ;
        RECT 9.008 10.052 9.04 10.084 ;
  LAYER M2 ;
        RECT 6.64 10.116 6.672 10.148 ;
  LAYER M2 ;
        RECT 9.008 10.18 9.04 10.212 ;
  LAYER M2 ;
        RECT 6.64 10.244 6.672 10.276 ;
  LAYER M2 ;
        RECT 9.008 10.308 9.04 10.34 ;
  LAYER M2 ;
        RECT 6.64 10.372 6.672 10.404 ;
  LAYER M2 ;
        RECT 9.008 10.436 9.04 10.468 ;
  LAYER M2 ;
        RECT 6.592 8.064 9.088 10.668 ;
  LAYER M1 ;
        RECT 6.64 11.22 6.672 13.728 ;
  LAYER M3 ;
        RECT 6.64 13.676 6.672 13.708 ;
  LAYER M1 ;
        RECT 6.704 11.22 6.736 13.728 ;
  LAYER M3 ;
        RECT 6.704 11.24 6.736 11.272 ;
  LAYER M1 ;
        RECT 6.768 11.22 6.8 13.728 ;
  LAYER M3 ;
        RECT 6.768 13.676 6.8 13.708 ;
  LAYER M1 ;
        RECT 6.832 11.22 6.864 13.728 ;
  LAYER M3 ;
        RECT 6.832 11.24 6.864 11.272 ;
  LAYER M1 ;
        RECT 6.896 11.22 6.928 13.728 ;
  LAYER M3 ;
        RECT 6.896 13.676 6.928 13.708 ;
  LAYER M1 ;
        RECT 6.96 11.22 6.992 13.728 ;
  LAYER M3 ;
        RECT 6.96 11.24 6.992 11.272 ;
  LAYER M1 ;
        RECT 7.024 11.22 7.056 13.728 ;
  LAYER M3 ;
        RECT 7.024 13.676 7.056 13.708 ;
  LAYER M1 ;
        RECT 7.088 11.22 7.12 13.728 ;
  LAYER M3 ;
        RECT 7.088 11.24 7.12 11.272 ;
  LAYER M1 ;
        RECT 7.152 11.22 7.184 13.728 ;
  LAYER M3 ;
        RECT 7.152 13.676 7.184 13.708 ;
  LAYER M1 ;
        RECT 7.216 11.22 7.248 13.728 ;
  LAYER M3 ;
        RECT 7.216 11.24 7.248 11.272 ;
  LAYER M1 ;
        RECT 7.28 11.22 7.312 13.728 ;
  LAYER M3 ;
        RECT 7.28 13.676 7.312 13.708 ;
  LAYER M1 ;
        RECT 7.344 11.22 7.376 13.728 ;
  LAYER M3 ;
        RECT 7.344 11.24 7.376 11.272 ;
  LAYER M1 ;
        RECT 7.408 11.22 7.44 13.728 ;
  LAYER M3 ;
        RECT 7.408 13.676 7.44 13.708 ;
  LAYER M1 ;
        RECT 7.472 11.22 7.504 13.728 ;
  LAYER M3 ;
        RECT 7.472 11.24 7.504 11.272 ;
  LAYER M1 ;
        RECT 7.536 11.22 7.568 13.728 ;
  LAYER M3 ;
        RECT 7.536 13.676 7.568 13.708 ;
  LAYER M1 ;
        RECT 7.6 11.22 7.632 13.728 ;
  LAYER M3 ;
        RECT 7.6 11.24 7.632 11.272 ;
  LAYER M1 ;
        RECT 7.664 11.22 7.696 13.728 ;
  LAYER M3 ;
        RECT 7.664 13.676 7.696 13.708 ;
  LAYER M1 ;
        RECT 7.728 11.22 7.76 13.728 ;
  LAYER M3 ;
        RECT 7.728 11.24 7.76 11.272 ;
  LAYER M1 ;
        RECT 7.792 11.22 7.824 13.728 ;
  LAYER M3 ;
        RECT 7.792 13.676 7.824 13.708 ;
  LAYER M1 ;
        RECT 7.856 11.22 7.888 13.728 ;
  LAYER M3 ;
        RECT 7.856 11.24 7.888 11.272 ;
  LAYER M1 ;
        RECT 7.92 11.22 7.952 13.728 ;
  LAYER M3 ;
        RECT 7.92 13.676 7.952 13.708 ;
  LAYER M1 ;
        RECT 7.984 11.22 8.016 13.728 ;
  LAYER M3 ;
        RECT 7.984 11.24 8.016 11.272 ;
  LAYER M1 ;
        RECT 8.048 11.22 8.08 13.728 ;
  LAYER M3 ;
        RECT 8.048 13.676 8.08 13.708 ;
  LAYER M1 ;
        RECT 8.112 11.22 8.144 13.728 ;
  LAYER M3 ;
        RECT 8.112 11.24 8.144 11.272 ;
  LAYER M1 ;
        RECT 8.176 11.22 8.208 13.728 ;
  LAYER M3 ;
        RECT 8.176 13.676 8.208 13.708 ;
  LAYER M1 ;
        RECT 8.24 11.22 8.272 13.728 ;
  LAYER M3 ;
        RECT 8.24 11.24 8.272 11.272 ;
  LAYER M1 ;
        RECT 8.304 11.22 8.336 13.728 ;
  LAYER M3 ;
        RECT 8.304 13.676 8.336 13.708 ;
  LAYER M1 ;
        RECT 8.368 11.22 8.4 13.728 ;
  LAYER M3 ;
        RECT 8.368 11.24 8.4 11.272 ;
  LAYER M1 ;
        RECT 8.432 11.22 8.464 13.728 ;
  LAYER M3 ;
        RECT 8.432 13.676 8.464 13.708 ;
  LAYER M1 ;
        RECT 8.496 11.22 8.528 13.728 ;
  LAYER M3 ;
        RECT 8.496 11.24 8.528 11.272 ;
  LAYER M1 ;
        RECT 8.56 11.22 8.592 13.728 ;
  LAYER M3 ;
        RECT 8.56 13.676 8.592 13.708 ;
  LAYER M1 ;
        RECT 8.624 11.22 8.656 13.728 ;
  LAYER M3 ;
        RECT 8.624 11.24 8.656 11.272 ;
  LAYER M1 ;
        RECT 8.688 11.22 8.72 13.728 ;
  LAYER M3 ;
        RECT 8.688 13.676 8.72 13.708 ;
  LAYER M1 ;
        RECT 8.752 11.22 8.784 13.728 ;
  LAYER M3 ;
        RECT 8.752 11.24 8.784 11.272 ;
  LAYER M1 ;
        RECT 8.816 11.22 8.848 13.728 ;
  LAYER M3 ;
        RECT 8.816 13.676 8.848 13.708 ;
  LAYER M1 ;
        RECT 8.88 11.22 8.912 13.728 ;
  LAYER M3 ;
        RECT 8.88 11.24 8.912 11.272 ;
  LAYER M1 ;
        RECT 8.944 11.22 8.976 13.728 ;
  LAYER M3 ;
        RECT 8.944 13.676 8.976 13.708 ;
  LAYER M1 ;
        RECT 9.008 11.22 9.04 13.728 ;
  LAYER M3 ;
        RECT 6.64 11.304 6.672 11.336 ;
  LAYER M2 ;
        RECT 9.008 11.368 9.04 11.4 ;
  LAYER M2 ;
        RECT 6.64 11.432 6.672 11.464 ;
  LAYER M2 ;
        RECT 9.008 11.496 9.04 11.528 ;
  LAYER M2 ;
        RECT 6.64 11.56 6.672 11.592 ;
  LAYER M2 ;
        RECT 9.008 11.624 9.04 11.656 ;
  LAYER M2 ;
        RECT 6.64 11.688 6.672 11.72 ;
  LAYER M2 ;
        RECT 9.008 11.752 9.04 11.784 ;
  LAYER M2 ;
        RECT 6.64 11.816 6.672 11.848 ;
  LAYER M2 ;
        RECT 9.008 11.88 9.04 11.912 ;
  LAYER M2 ;
        RECT 6.64 11.944 6.672 11.976 ;
  LAYER M2 ;
        RECT 9.008 12.008 9.04 12.04 ;
  LAYER M2 ;
        RECT 6.64 12.072 6.672 12.104 ;
  LAYER M2 ;
        RECT 9.008 12.136 9.04 12.168 ;
  LAYER M2 ;
        RECT 6.64 12.2 6.672 12.232 ;
  LAYER M2 ;
        RECT 9.008 12.264 9.04 12.296 ;
  LAYER M2 ;
        RECT 6.64 12.328 6.672 12.36 ;
  LAYER M2 ;
        RECT 9.008 12.392 9.04 12.424 ;
  LAYER M2 ;
        RECT 6.64 12.456 6.672 12.488 ;
  LAYER M2 ;
        RECT 9.008 12.52 9.04 12.552 ;
  LAYER M2 ;
        RECT 6.64 12.584 6.672 12.616 ;
  LAYER M2 ;
        RECT 9.008 12.648 9.04 12.68 ;
  LAYER M2 ;
        RECT 6.64 12.712 6.672 12.744 ;
  LAYER M2 ;
        RECT 9.008 12.776 9.04 12.808 ;
  LAYER M2 ;
        RECT 6.64 12.84 6.672 12.872 ;
  LAYER M2 ;
        RECT 9.008 12.904 9.04 12.936 ;
  LAYER M2 ;
        RECT 6.64 12.968 6.672 13 ;
  LAYER M2 ;
        RECT 9.008 13.032 9.04 13.064 ;
  LAYER M2 ;
        RECT 6.64 13.096 6.672 13.128 ;
  LAYER M2 ;
        RECT 9.008 13.16 9.04 13.192 ;
  LAYER M2 ;
        RECT 6.64 13.224 6.672 13.256 ;
  LAYER M2 ;
        RECT 9.008 13.288 9.04 13.32 ;
  LAYER M2 ;
        RECT 6.64 13.352 6.672 13.384 ;
  LAYER M2 ;
        RECT 9.008 13.416 9.04 13.448 ;
  LAYER M2 ;
        RECT 6.64 13.48 6.672 13.512 ;
  LAYER M2 ;
        RECT 9.008 13.544 9.04 13.576 ;
  LAYER M2 ;
        RECT 6.592 11.172 9.088 13.776 ;
  LAYER M1 ;
        RECT 9.616 1.896 9.648 4.404 ;
  LAYER M3 ;
        RECT 9.616 4.352 9.648 4.384 ;
  LAYER M1 ;
        RECT 9.68 1.896 9.712 4.404 ;
  LAYER M3 ;
        RECT 9.68 1.916 9.712 1.948 ;
  LAYER M1 ;
        RECT 9.744 1.896 9.776 4.404 ;
  LAYER M3 ;
        RECT 9.744 4.352 9.776 4.384 ;
  LAYER M1 ;
        RECT 9.808 1.896 9.84 4.404 ;
  LAYER M3 ;
        RECT 9.808 1.916 9.84 1.948 ;
  LAYER M1 ;
        RECT 9.872 1.896 9.904 4.404 ;
  LAYER M3 ;
        RECT 9.872 4.352 9.904 4.384 ;
  LAYER M1 ;
        RECT 9.936 1.896 9.968 4.404 ;
  LAYER M3 ;
        RECT 9.936 1.916 9.968 1.948 ;
  LAYER M1 ;
        RECT 10 1.896 10.032 4.404 ;
  LAYER M3 ;
        RECT 10 4.352 10.032 4.384 ;
  LAYER M1 ;
        RECT 10.064 1.896 10.096 4.404 ;
  LAYER M3 ;
        RECT 10.064 1.916 10.096 1.948 ;
  LAYER M1 ;
        RECT 10.128 1.896 10.16 4.404 ;
  LAYER M3 ;
        RECT 10.128 4.352 10.16 4.384 ;
  LAYER M1 ;
        RECT 10.192 1.896 10.224 4.404 ;
  LAYER M3 ;
        RECT 10.192 1.916 10.224 1.948 ;
  LAYER M1 ;
        RECT 10.256 1.896 10.288 4.404 ;
  LAYER M3 ;
        RECT 10.256 4.352 10.288 4.384 ;
  LAYER M1 ;
        RECT 10.32 1.896 10.352 4.404 ;
  LAYER M3 ;
        RECT 10.32 1.916 10.352 1.948 ;
  LAYER M1 ;
        RECT 10.384 1.896 10.416 4.404 ;
  LAYER M3 ;
        RECT 10.384 4.352 10.416 4.384 ;
  LAYER M1 ;
        RECT 10.448 1.896 10.48 4.404 ;
  LAYER M3 ;
        RECT 10.448 1.916 10.48 1.948 ;
  LAYER M1 ;
        RECT 10.512 1.896 10.544 4.404 ;
  LAYER M3 ;
        RECT 10.512 4.352 10.544 4.384 ;
  LAYER M1 ;
        RECT 10.576 1.896 10.608 4.404 ;
  LAYER M3 ;
        RECT 10.576 1.916 10.608 1.948 ;
  LAYER M1 ;
        RECT 10.64 1.896 10.672 4.404 ;
  LAYER M3 ;
        RECT 10.64 4.352 10.672 4.384 ;
  LAYER M1 ;
        RECT 10.704 1.896 10.736 4.404 ;
  LAYER M3 ;
        RECT 10.704 1.916 10.736 1.948 ;
  LAYER M1 ;
        RECT 10.768 1.896 10.8 4.404 ;
  LAYER M3 ;
        RECT 10.768 4.352 10.8 4.384 ;
  LAYER M1 ;
        RECT 10.832 1.896 10.864 4.404 ;
  LAYER M3 ;
        RECT 10.832 1.916 10.864 1.948 ;
  LAYER M1 ;
        RECT 10.896 1.896 10.928 4.404 ;
  LAYER M3 ;
        RECT 10.896 4.352 10.928 4.384 ;
  LAYER M1 ;
        RECT 10.96 1.896 10.992 4.404 ;
  LAYER M3 ;
        RECT 10.96 1.916 10.992 1.948 ;
  LAYER M1 ;
        RECT 11.024 1.896 11.056 4.404 ;
  LAYER M3 ;
        RECT 11.024 4.352 11.056 4.384 ;
  LAYER M1 ;
        RECT 11.088 1.896 11.12 4.404 ;
  LAYER M3 ;
        RECT 11.088 1.916 11.12 1.948 ;
  LAYER M1 ;
        RECT 11.152 1.896 11.184 4.404 ;
  LAYER M3 ;
        RECT 11.152 4.352 11.184 4.384 ;
  LAYER M1 ;
        RECT 11.216 1.896 11.248 4.404 ;
  LAYER M3 ;
        RECT 11.216 1.916 11.248 1.948 ;
  LAYER M1 ;
        RECT 11.28 1.896 11.312 4.404 ;
  LAYER M3 ;
        RECT 11.28 4.352 11.312 4.384 ;
  LAYER M1 ;
        RECT 11.344 1.896 11.376 4.404 ;
  LAYER M3 ;
        RECT 11.344 1.916 11.376 1.948 ;
  LAYER M1 ;
        RECT 11.408 1.896 11.44 4.404 ;
  LAYER M3 ;
        RECT 11.408 4.352 11.44 4.384 ;
  LAYER M1 ;
        RECT 11.472 1.896 11.504 4.404 ;
  LAYER M3 ;
        RECT 11.472 1.916 11.504 1.948 ;
  LAYER M1 ;
        RECT 11.536 1.896 11.568 4.404 ;
  LAYER M3 ;
        RECT 11.536 4.352 11.568 4.384 ;
  LAYER M1 ;
        RECT 11.6 1.896 11.632 4.404 ;
  LAYER M3 ;
        RECT 11.6 1.916 11.632 1.948 ;
  LAYER M1 ;
        RECT 11.664 1.896 11.696 4.404 ;
  LAYER M3 ;
        RECT 11.664 4.352 11.696 4.384 ;
  LAYER M1 ;
        RECT 11.728 1.896 11.76 4.404 ;
  LAYER M3 ;
        RECT 11.728 1.916 11.76 1.948 ;
  LAYER M1 ;
        RECT 11.792 1.896 11.824 4.404 ;
  LAYER M3 ;
        RECT 11.792 4.352 11.824 4.384 ;
  LAYER M1 ;
        RECT 11.856 1.896 11.888 4.404 ;
  LAYER M3 ;
        RECT 11.856 1.916 11.888 1.948 ;
  LAYER M1 ;
        RECT 11.92 1.896 11.952 4.404 ;
  LAYER M3 ;
        RECT 11.92 4.352 11.952 4.384 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 4.404 ;
  LAYER M3 ;
        RECT 9.616 1.98 9.648 2.012 ;
  LAYER M2 ;
        RECT 11.984 2.044 12.016 2.076 ;
  LAYER M2 ;
        RECT 9.616 2.108 9.648 2.14 ;
  LAYER M2 ;
        RECT 11.984 2.172 12.016 2.204 ;
  LAYER M2 ;
        RECT 9.616 2.236 9.648 2.268 ;
  LAYER M2 ;
        RECT 11.984 2.3 12.016 2.332 ;
  LAYER M2 ;
        RECT 9.616 2.364 9.648 2.396 ;
  LAYER M2 ;
        RECT 11.984 2.428 12.016 2.46 ;
  LAYER M2 ;
        RECT 9.616 2.492 9.648 2.524 ;
  LAYER M2 ;
        RECT 11.984 2.556 12.016 2.588 ;
  LAYER M2 ;
        RECT 9.616 2.62 9.648 2.652 ;
  LAYER M2 ;
        RECT 11.984 2.684 12.016 2.716 ;
  LAYER M2 ;
        RECT 9.616 2.748 9.648 2.78 ;
  LAYER M2 ;
        RECT 11.984 2.812 12.016 2.844 ;
  LAYER M2 ;
        RECT 9.616 2.876 9.648 2.908 ;
  LAYER M2 ;
        RECT 11.984 2.94 12.016 2.972 ;
  LAYER M2 ;
        RECT 9.616 3.004 9.648 3.036 ;
  LAYER M2 ;
        RECT 11.984 3.068 12.016 3.1 ;
  LAYER M2 ;
        RECT 9.616 3.132 9.648 3.164 ;
  LAYER M2 ;
        RECT 11.984 3.196 12.016 3.228 ;
  LAYER M2 ;
        RECT 9.616 3.26 9.648 3.292 ;
  LAYER M2 ;
        RECT 11.984 3.324 12.016 3.356 ;
  LAYER M2 ;
        RECT 9.616 3.388 9.648 3.42 ;
  LAYER M2 ;
        RECT 11.984 3.452 12.016 3.484 ;
  LAYER M2 ;
        RECT 9.616 3.516 9.648 3.548 ;
  LAYER M2 ;
        RECT 11.984 3.58 12.016 3.612 ;
  LAYER M2 ;
        RECT 9.616 3.644 9.648 3.676 ;
  LAYER M2 ;
        RECT 11.984 3.708 12.016 3.74 ;
  LAYER M2 ;
        RECT 9.616 3.772 9.648 3.804 ;
  LAYER M2 ;
        RECT 11.984 3.836 12.016 3.868 ;
  LAYER M2 ;
        RECT 9.616 3.9 9.648 3.932 ;
  LAYER M2 ;
        RECT 11.984 3.964 12.016 3.996 ;
  LAYER M2 ;
        RECT 9.616 4.028 9.648 4.06 ;
  LAYER M2 ;
        RECT 11.984 4.092 12.016 4.124 ;
  LAYER M2 ;
        RECT 9.616 4.156 9.648 4.188 ;
  LAYER M2 ;
        RECT 11.984 4.22 12.016 4.252 ;
  LAYER M2 ;
        RECT 9.568 1.848 12.064 4.452 ;
  LAYER M1 ;
        RECT 9.616 5.004 9.648 7.512 ;
  LAYER M3 ;
        RECT 9.616 7.46 9.648 7.492 ;
  LAYER M1 ;
        RECT 9.68 5.004 9.712 7.512 ;
  LAYER M3 ;
        RECT 9.68 5.024 9.712 5.056 ;
  LAYER M1 ;
        RECT 9.744 5.004 9.776 7.512 ;
  LAYER M3 ;
        RECT 9.744 7.46 9.776 7.492 ;
  LAYER M1 ;
        RECT 9.808 5.004 9.84 7.512 ;
  LAYER M3 ;
        RECT 9.808 5.024 9.84 5.056 ;
  LAYER M1 ;
        RECT 9.872 5.004 9.904 7.512 ;
  LAYER M3 ;
        RECT 9.872 7.46 9.904 7.492 ;
  LAYER M1 ;
        RECT 9.936 5.004 9.968 7.512 ;
  LAYER M3 ;
        RECT 9.936 5.024 9.968 5.056 ;
  LAYER M1 ;
        RECT 10 5.004 10.032 7.512 ;
  LAYER M3 ;
        RECT 10 7.46 10.032 7.492 ;
  LAYER M1 ;
        RECT 10.064 5.004 10.096 7.512 ;
  LAYER M3 ;
        RECT 10.064 5.024 10.096 5.056 ;
  LAYER M1 ;
        RECT 10.128 5.004 10.16 7.512 ;
  LAYER M3 ;
        RECT 10.128 7.46 10.16 7.492 ;
  LAYER M1 ;
        RECT 10.192 5.004 10.224 7.512 ;
  LAYER M3 ;
        RECT 10.192 5.024 10.224 5.056 ;
  LAYER M1 ;
        RECT 10.256 5.004 10.288 7.512 ;
  LAYER M3 ;
        RECT 10.256 7.46 10.288 7.492 ;
  LAYER M1 ;
        RECT 10.32 5.004 10.352 7.512 ;
  LAYER M3 ;
        RECT 10.32 5.024 10.352 5.056 ;
  LAYER M1 ;
        RECT 10.384 5.004 10.416 7.512 ;
  LAYER M3 ;
        RECT 10.384 7.46 10.416 7.492 ;
  LAYER M1 ;
        RECT 10.448 5.004 10.48 7.512 ;
  LAYER M3 ;
        RECT 10.448 5.024 10.48 5.056 ;
  LAYER M1 ;
        RECT 10.512 5.004 10.544 7.512 ;
  LAYER M3 ;
        RECT 10.512 7.46 10.544 7.492 ;
  LAYER M1 ;
        RECT 10.576 5.004 10.608 7.512 ;
  LAYER M3 ;
        RECT 10.576 5.024 10.608 5.056 ;
  LAYER M1 ;
        RECT 10.64 5.004 10.672 7.512 ;
  LAYER M3 ;
        RECT 10.64 7.46 10.672 7.492 ;
  LAYER M1 ;
        RECT 10.704 5.004 10.736 7.512 ;
  LAYER M3 ;
        RECT 10.704 5.024 10.736 5.056 ;
  LAYER M1 ;
        RECT 10.768 5.004 10.8 7.512 ;
  LAYER M3 ;
        RECT 10.768 7.46 10.8 7.492 ;
  LAYER M1 ;
        RECT 10.832 5.004 10.864 7.512 ;
  LAYER M3 ;
        RECT 10.832 5.024 10.864 5.056 ;
  LAYER M1 ;
        RECT 10.896 5.004 10.928 7.512 ;
  LAYER M3 ;
        RECT 10.896 7.46 10.928 7.492 ;
  LAYER M1 ;
        RECT 10.96 5.004 10.992 7.512 ;
  LAYER M3 ;
        RECT 10.96 5.024 10.992 5.056 ;
  LAYER M1 ;
        RECT 11.024 5.004 11.056 7.512 ;
  LAYER M3 ;
        RECT 11.024 7.46 11.056 7.492 ;
  LAYER M1 ;
        RECT 11.088 5.004 11.12 7.512 ;
  LAYER M3 ;
        RECT 11.088 5.024 11.12 5.056 ;
  LAYER M1 ;
        RECT 11.152 5.004 11.184 7.512 ;
  LAYER M3 ;
        RECT 11.152 7.46 11.184 7.492 ;
  LAYER M1 ;
        RECT 11.216 5.004 11.248 7.512 ;
  LAYER M3 ;
        RECT 11.216 5.024 11.248 5.056 ;
  LAYER M1 ;
        RECT 11.28 5.004 11.312 7.512 ;
  LAYER M3 ;
        RECT 11.28 7.46 11.312 7.492 ;
  LAYER M1 ;
        RECT 11.344 5.004 11.376 7.512 ;
  LAYER M3 ;
        RECT 11.344 5.024 11.376 5.056 ;
  LAYER M1 ;
        RECT 11.408 5.004 11.44 7.512 ;
  LAYER M3 ;
        RECT 11.408 7.46 11.44 7.492 ;
  LAYER M1 ;
        RECT 11.472 5.004 11.504 7.512 ;
  LAYER M3 ;
        RECT 11.472 5.024 11.504 5.056 ;
  LAYER M1 ;
        RECT 11.536 5.004 11.568 7.512 ;
  LAYER M3 ;
        RECT 11.536 7.46 11.568 7.492 ;
  LAYER M1 ;
        RECT 11.6 5.004 11.632 7.512 ;
  LAYER M3 ;
        RECT 11.6 5.024 11.632 5.056 ;
  LAYER M1 ;
        RECT 11.664 5.004 11.696 7.512 ;
  LAYER M3 ;
        RECT 11.664 7.46 11.696 7.492 ;
  LAYER M1 ;
        RECT 11.728 5.004 11.76 7.512 ;
  LAYER M3 ;
        RECT 11.728 5.024 11.76 5.056 ;
  LAYER M1 ;
        RECT 11.792 5.004 11.824 7.512 ;
  LAYER M3 ;
        RECT 11.792 7.46 11.824 7.492 ;
  LAYER M1 ;
        RECT 11.856 5.004 11.888 7.512 ;
  LAYER M3 ;
        RECT 11.856 5.024 11.888 5.056 ;
  LAYER M1 ;
        RECT 11.92 5.004 11.952 7.512 ;
  LAYER M3 ;
        RECT 11.92 7.46 11.952 7.492 ;
  LAYER M1 ;
        RECT 11.984 5.004 12.016 7.512 ;
  LAYER M3 ;
        RECT 9.616 5.088 9.648 5.12 ;
  LAYER M2 ;
        RECT 11.984 5.152 12.016 5.184 ;
  LAYER M2 ;
        RECT 9.616 5.216 9.648 5.248 ;
  LAYER M2 ;
        RECT 11.984 5.28 12.016 5.312 ;
  LAYER M2 ;
        RECT 9.616 5.344 9.648 5.376 ;
  LAYER M2 ;
        RECT 11.984 5.408 12.016 5.44 ;
  LAYER M2 ;
        RECT 9.616 5.472 9.648 5.504 ;
  LAYER M2 ;
        RECT 11.984 5.536 12.016 5.568 ;
  LAYER M2 ;
        RECT 9.616 5.6 9.648 5.632 ;
  LAYER M2 ;
        RECT 11.984 5.664 12.016 5.696 ;
  LAYER M2 ;
        RECT 9.616 5.728 9.648 5.76 ;
  LAYER M2 ;
        RECT 11.984 5.792 12.016 5.824 ;
  LAYER M2 ;
        RECT 9.616 5.856 9.648 5.888 ;
  LAYER M2 ;
        RECT 11.984 5.92 12.016 5.952 ;
  LAYER M2 ;
        RECT 9.616 5.984 9.648 6.016 ;
  LAYER M2 ;
        RECT 11.984 6.048 12.016 6.08 ;
  LAYER M2 ;
        RECT 9.616 6.112 9.648 6.144 ;
  LAYER M2 ;
        RECT 11.984 6.176 12.016 6.208 ;
  LAYER M2 ;
        RECT 9.616 6.24 9.648 6.272 ;
  LAYER M2 ;
        RECT 11.984 6.304 12.016 6.336 ;
  LAYER M2 ;
        RECT 9.616 6.368 9.648 6.4 ;
  LAYER M2 ;
        RECT 11.984 6.432 12.016 6.464 ;
  LAYER M2 ;
        RECT 9.616 6.496 9.648 6.528 ;
  LAYER M2 ;
        RECT 11.984 6.56 12.016 6.592 ;
  LAYER M2 ;
        RECT 9.616 6.624 9.648 6.656 ;
  LAYER M2 ;
        RECT 11.984 6.688 12.016 6.72 ;
  LAYER M2 ;
        RECT 9.616 6.752 9.648 6.784 ;
  LAYER M2 ;
        RECT 11.984 6.816 12.016 6.848 ;
  LAYER M2 ;
        RECT 9.616 6.88 9.648 6.912 ;
  LAYER M2 ;
        RECT 11.984 6.944 12.016 6.976 ;
  LAYER M2 ;
        RECT 9.616 7.008 9.648 7.04 ;
  LAYER M2 ;
        RECT 11.984 7.072 12.016 7.104 ;
  LAYER M2 ;
        RECT 9.616 7.136 9.648 7.168 ;
  LAYER M2 ;
        RECT 11.984 7.2 12.016 7.232 ;
  LAYER M2 ;
        RECT 9.616 7.264 9.648 7.296 ;
  LAYER M2 ;
        RECT 11.984 7.328 12.016 7.36 ;
  LAYER M2 ;
        RECT 9.568 4.956 12.064 7.56 ;
  LAYER M1 ;
        RECT 9.616 8.112 9.648 10.62 ;
  LAYER M3 ;
        RECT 9.616 10.568 9.648 10.6 ;
  LAYER M1 ;
        RECT 9.68 8.112 9.712 10.62 ;
  LAYER M3 ;
        RECT 9.68 8.132 9.712 8.164 ;
  LAYER M1 ;
        RECT 9.744 8.112 9.776 10.62 ;
  LAYER M3 ;
        RECT 9.744 10.568 9.776 10.6 ;
  LAYER M1 ;
        RECT 9.808 8.112 9.84 10.62 ;
  LAYER M3 ;
        RECT 9.808 8.132 9.84 8.164 ;
  LAYER M1 ;
        RECT 9.872 8.112 9.904 10.62 ;
  LAYER M3 ;
        RECT 9.872 10.568 9.904 10.6 ;
  LAYER M1 ;
        RECT 9.936 8.112 9.968 10.62 ;
  LAYER M3 ;
        RECT 9.936 8.132 9.968 8.164 ;
  LAYER M1 ;
        RECT 10 8.112 10.032 10.62 ;
  LAYER M3 ;
        RECT 10 10.568 10.032 10.6 ;
  LAYER M1 ;
        RECT 10.064 8.112 10.096 10.62 ;
  LAYER M3 ;
        RECT 10.064 8.132 10.096 8.164 ;
  LAYER M1 ;
        RECT 10.128 8.112 10.16 10.62 ;
  LAYER M3 ;
        RECT 10.128 10.568 10.16 10.6 ;
  LAYER M1 ;
        RECT 10.192 8.112 10.224 10.62 ;
  LAYER M3 ;
        RECT 10.192 8.132 10.224 8.164 ;
  LAYER M1 ;
        RECT 10.256 8.112 10.288 10.62 ;
  LAYER M3 ;
        RECT 10.256 10.568 10.288 10.6 ;
  LAYER M1 ;
        RECT 10.32 8.112 10.352 10.62 ;
  LAYER M3 ;
        RECT 10.32 8.132 10.352 8.164 ;
  LAYER M1 ;
        RECT 10.384 8.112 10.416 10.62 ;
  LAYER M3 ;
        RECT 10.384 10.568 10.416 10.6 ;
  LAYER M1 ;
        RECT 10.448 8.112 10.48 10.62 ;
  LAYER M3 ;
        RECT 10.448 8.132 10.48 8.164 ;
  LAYER M1 ;
        RECT 10.512 8.112 10.544 10.62 ;
  LAYER M3 ;
        RECT 10.512 10.568 10.544 10.6 ;
  LAYER M1 ;
        RECT 10.576 8.112 10.608 10.62 ;
  LAYER M3 ;
        RECT 10.576 8.132 10.608 8.164 ;
  LAYER M1 ;
        RECT 10.64 8.112 10.672 10.62 ;
  LAYER M3 ;
        RECT 10.64 10.568 10.672 10.6 ;
  LAYER M1 ;
        RECT 10.704 8.112 10.736 10.62 ;
  LAYER M3 ;
        RECT 10.704 8.132 10.736 8.164 ;
  LAYER M1 ;
        RECT 10.768 8.112 10.8 10.62 ;
  LAYER M3 ;
        RECT 10.768 10.568 10.8 10.6 ;
  LAYER M1 ;
        RECT 10.832 8.112 10.864 10.62 ;
  LAYER M3 ;
        RECT 10.832 8.132 10.864 8.164 ;
  LAYER M1 ;
        RECT 10.896 8.112 10.928 10.62 ;
  LAYER M3 ;
        RECT 10.896 10.568 10.928 10.6 ;
  LAYER M1 ;
        RECT 10.96 8.112 10.992 10.62 ;
  LAYER M3 ;
        RECT 10.96 8.132 10.992 8.164 ;
  LAYER M1 ;
        RECT 11.024 8.112 11.056 10.62 ;
  LAYER M3 ;
        RECT 11.024 10.568 11.056 10.6 ;
  LAYER M1 ;
        RECT 11.088 8.112 11.12 10.62 ;
  LAYER M3 ;
        RECT 11.088 8.132 11.12 8.164 ;
  LAYER M1 ;
        RECT 11.152 8.112 11.184 10.62 ;
  LAYER M3 ;
        RECT 11.152 10.568 11.184 10.6 ;
  LAYER M1 ;
        RECT 11.216 8.112 11.248 10.62 ;
  LAYER M3 ;
        RECT 11.216 8.132 11.248 8.164 ;
  LAYER M1 ;
        RECT 11.28 8.112 11.312 10.62 ;
  LAYER M3 ;
        RECT 11.28 10.568 11.312 10.6 ;
  LAYER M1 ;
        RECT 11.344 8.112 11.376 10.62 ;
  LAYER M3 ;
        RECT 11.344 8.132 11.376 8.164 ;
  LAYER M1 ;
        RECT 11.408 8.112 11.44 10.62 ;
  LAYER M3 ;
        RECT 11.408 10.568 11.44 10.6 ;
  LAYER M1 ;
        RECT 11.472 8.112 11.504 10.62 ;
  LAYER M3 ;
        RECT 11.472 8.132 11.504 8.164 ;
  LAYER M1 ;
        RECT 11.536 8.112 11.568 10.62 ;
  LAYER M3 ;
        RECT 11.536 10.568 11.568 10.6 ;
  LAYER M1 ;
        RECT 11.6 8.112 11.632 10.62 ;
  LAYER M3 ;
        RECT 11.6 8.132 11.632 8.164 ;
  LAYER M1 ;
        RECT 11.664 8.112 11.696 10.62 ;
  LAYER M3 ;
        RECT 11.664 10.568 11.696 10.6 ;
  LAYER M1 ;
        RECT 11.728 8.112 11.76 10.62 ;
  LAYER M3 ;
        RECT 11.728 8.132 11.76 8.164 ;
  LAYER M1 ;
        RECT 11.792 8.112 11.824 10.62 ;
  LAYER M3 ;
        RECT 11.792 10.568 11.824 10.6 ;
  LAYER M1 ;
        RECT 11.856 8.112 11.888 10.62 ;
  LAYER M3 ;
        RECT 11.856 8.132 11.888 8.164 ;
  LAYER M1 ;
        RECT 11.92 8.112 11.952 10.62 ;
  LAYER M3 ;
        RECT 11.92 10.568 11.952 10.6 ;
  LAYER M1 ;
        RECT 11.984 8.112 12.016 10.62 ;
  LAYER M3 ;
        RECT 9.616 8.196 9.648 8.228 ;
  LAYER M2 ;
        RECT 11.984 8.26 12.016 8.292 ;
  LAYER M2 ;
        RECT 9.616 8.324 9.648 8.356 ;
  LAYER M2 ;
        RECT 11.984 8.388 12.016 8.42 ;
  LAYER M2 ;
        RECT 9.616 8.452 9.648 8.484 ;
  LAYER M2 ;
        RECT 11.984 8.516 12.016 8.548 ;
  LAYER M2 ;
        RECT 9.616 8.58 9.648 8.612 ;
  LAYER M2 ;
        RECT 11.984 8.644 12.016 8.676 ;
  LAYER M2 ;
        RECT 9.616 8.708 9.648 8.74 ;
  LAYER M2 ;
        RECT 11.984 8.772 12.016 8.804 ;
  LAYER M2 ;
        RECT 9.616 8.836 9.648 8.868 ;
  LAYER M2 ;
        RECT 11.984 8.9 12.016 8.932 ;
  LAYER M2 ;
        RECT 9.616 8.964 9.648 8.996 ;
  LAYER M2 ;
        RECT 11.984 9.028 12.016 9.06 ;
  LAYER M2 ;
        RECT 9.616 9.092 9.648 9.124 ;
  LAYER M2 ;
        RECT 11.984 9.156 12.016 9.188 ;
  LAYER M2 ;
        RECT 9.616 9.22 9.648 9.252 ;
  LAYER M2 ;
        RECT 11.984 9.284 12.016 9.316 ;
  LAYER M2 ;
        RECT 9.616 9.348 9.648 9.38 ;
  LAYER M2 ;
        RECT 11.984 9.412 12.016 9.444 ;
  LAYER M2 ;
        RECT 9.616 9.476 9.648 9.508 ;
  LAYER M2 ;
        RECT 11.984 9.54 12.016 9.572 ;
  LAYER M2 ;
        RECT 9.616 9.604 9.648 9.636 ;
  LAYER M2 ;
        RECT 11.984 9.668 12.016 9.7 ;
  LAYER M2 ;
        RECT 9.616 9.732 9.648 9.764 ;
  LAYER M2 ;
        RECT 11.984 9.796 12.016 9.828 ;
  LAYER M2 ;
        RECT 9.616 9.86 9.648 9.892 ;
  LAYER M2 ;
        RECT 11.984 9.924 12.016 9.956 ;
  LAYER M2 ;
        RECT 9.616 9.988 9.648 10.02 ;
  LAYER M2 ;
        RECT 11.984 10.052 12.016 10.084 ;
  LAYER M2 ;
        RECT 9.616 10.116 9.648 10.148 ;
  LAYER M2 ;
        RECT 11.984 10.18 12.016 10.212 ;
  LAYER M2 ;
        RECT 9.616 10.244 9.648 10.276 ;
  LAYER M2 ;
        RECT 11.984 10.308 12.016 10.34 ;
  LAYER M2 ;
        RECT 9.616 10.372 9.648 10.404 ;
  LAYER M2 ;
        RECT 11.984 10.436 12.016 10.468 ;
  LAYER M2 ;
        RECT 9.568 8.064 12.064 10.668 ;
  LAYER M1 ;
        RECT 9.616 11.22 9.648 13.728 ;
  LAYER M3 ;
        RECT 9.616 13.676 9.648 13.708 ;
  LAYER M1 ;
        RECT 9.68 11.22 9.712 13.728 ;
  LAYER M3 ;
        RECT 9.68 11.24 9.712 11.272 ;
  LAYER M1 ;
        RECT 9.744 11.22 9.776 13.728 ;
  LAYER M3 ;
        RECT 9.744 13.676 9.776 13.708 ;
  LAYER M1 ;
        RECT 9.808 11.22 9.84 13.728 ;
  LAYER M3 ;
        RECT 9.808 11.24 9.84 11.272 ;
  LAYER M1 ;
        RECT 9.872 11.22 9.904 13.728 ;
  LAYER M3 ;
        RECT 9.872 13.676 9.904 13.708 ;
  LAYER M1 ;
        RECT 9.936 11.22 9.968 13.728 ;
  LAYER M3 ;
        RECT 9.936 11.24 9.968 11.272 ;
  LAYER M1 ;
        RECT 10 11.22 10.032 13.728 ;
  LAYER M3 ;
        RECT 10 13.676 10.032 13.708 ;
  LAYER M1 ;
        RECT 10.064 11.22 10.096 13.728 ;
  LAYER M3 ;
        RECT 10.064 11.24 10.096 11.272 ;
  LAYER M1 ;
        RECT 10.128 11.22 10.16 13.728 ;
  LAYER M3 ;
        RECT 10.128 13.676 10.16 13.708 ;
  LAYER M1 ;
        RECT 10.192 11.22 10.224 13.728 ;
  LAYER M3 ;
        RECT 10.192 11.24 10.224 11.272 ;
  LAYER M1 ;
        RECT 10.256 11.22 10.288 13.728 ;
  LAYER M3 ;
        RECT 10.256 13.676 10.288 13.708 ;
  LAYER M1 ;
        RECT 10.32 11.22 10.352 13.728 ;
  LAYER M3 ;
        RECT 10.32 11.24 10.352 11.272 ;
  LAYER M1 ;
        RECT 10.384 11.22 10.416 13.728 ;
  LAYER M3 ;
        RECT 10.384 13.676 10.416 13.708 ;
  LAYER M1 ;
        RECT 10.448 11.22 10.48 13.728 ;
  LAYER M3 ;
        RECT 10.448 11.24 10.48 11.272 ;
  LAYER M1 ;
        RECT 10.512 11.22 10.544 13.728 ;
  LAYER M3 ;
        RECT 10.512 13.676 10.544 13.708 ;
  LAYER M1 ;
        RECT 10.576 11.22 10.608 13.728 ;
  LAYER M3 ;
        RECT 10.576 11.24 10.608 11.272 ;
  LAYER M1 ;
        RECT 10.64 11.22 10.672 13.728 ;
  LAYER M3 ;
        RECT 10.64 13.676 10.672 13.708 ;
  LAYER M1 ;
        RECT 10.704 11.22 10.736 13.728 ;
  LAYER M3 ;
        RECT 10.704 11.24 10.736 11.272 ;
  LAYER M1 ;
        RECT 10.768 11.22 10.8 13.728 ;
  LAYER M3 ;
        RECT 10.768 13.676 10.8 13.708 ;
  LAYER M1 ;
        RECT 10.832 11.22 10.864 13.728 ;
  LAYER M3 ;
        RECT 10.832 11.24 10.864 11.272 ;
  LAYER M1 ;
        RECT 10.896 11.22 10.928 13.728 ;
  LAYER M3 ;
        RECT 10.896 13.676 10.928 13.708 ;
  LAYER M1 ;
        RECT 10.96 11.22 10.992 13.728 ;
  LAYER M3 ;
        RECT 10.96 11.24 10.992 11.272 ;
  LAYER M1 ;
        RECT 11.024 11.22 11.056 13.728 ;
  LAYER M3 ;
        RECT 11.024 13.676 11.056 13.708 ;
  LAYER M1 ;
        RECT 11.088 11.22 11.12 13.728 ;
  LAYER M3 ;
        RECT 11.088 11.24 11.12 11.272 ;
  LAYER M1 ;
        RECT 11.152 11.22 11.184 13.728 ;
  LAYER M3 ;
        RECT 11.152 13.676 11.184 13.708 ;
  LAYER M1 ;
        RECT 11.216 11.22 11.248 13.728 ;
  LAYER M3 ;
        RECT 11.216 11.24 11.248 11.272 ;
  LAYER M1 ;
        RECT 11.28 11.22 11.312 13.728 ;
  LAYER M3 ;
        RECT 11.28 13.676 11.312 13.708 ;
  LAYER M1 ;
        RECT 11.344 11.22 11.376 13.728 ;
  LAYER M3 ;
        RECT 11.344 11.24 11.376 11.272 ;
  LAYER M1 ;
        RECT 11.408 11.22 11.44 13.728 ;
  LAYER M3 ;
        RECT 11.408 13.676 11.44 13.708 ;
  LAYER M1 ;
        RECT 11.472 11.22 11.504 13.728 ;
  LAYER M3 ;
        RECT 11.472 11.24 11.504 11.272 ;
  LAYER M1 ;
        RECT 11.536 11.22 11.568 13.728 ;
  LAYER M3 ;
        RECT 11.536 13.676 11.568 13.708 ;
  LAYER M1 ;
        RECT 11.6 11.22 11.632 13.728 ;
  LAYER M3 ;
        RECT 11.6 11.24 11.632 11.272 ;
  LAYER M1 ;
        RECT 11.664 11.22 11.696 13.728 ;
  LAYER M3 ;
        RECT 11.664 13.676 11.696 13.708 ;
  LAYER M1 ;
        RECT 11.728 11.22 11.76 13.728 ;
  LAYER M3 ;
        RECT 11.728 11.24 11.76 11.272 ;
  LAYER M1 ;
        RECT 11.792 11.22 11.824 13.728 ;
  LAYER M3 ;
        RECT 11.792 13.676 11.824 13.708 ;
  LAYER M1 ;
        RECT 11.856 11.22 11.888 13.728 ;
  LAYER M3 ;
        RECT 11.856 11.24 11.888 11.272 ;
  LAYER M1 ;
        RECT 11.92 11.22 11.952 13.728 ;
  LAYER M3 ;
        RECT 11.92 13.676 11.952 13.708 ;
  LAYER M1 ;
        RECT 11.984 11.22 12.016 13.728 ;
  LAYER M3 ;
        RECT 9.616 11.304 9.648 11.336 ;
  LAYER M2 ;
        RECT 11.984 11.368 12.016 11.4 ;
  LAYER M2 ;
        RECT 9.616 11.432 9.648 11.464 ;
  LAYER M2 ;
        RECT 11.984 11.496 12.016 11.528 ;
  LAYER M2 ;
        RECT 9.616 11.56 9.648 11.592 ;
  LAYER M2 ;
        RECT 11.984 11.624 12.016 11.656 ;
  LAYER M2 ;
        RECT 9.616 11.688 9.648 11.72 ;
  LAYER M2 ;
        RECT 11.984 11.752 12.016 11.784 ;
  LAYER M2 ;
        RECT 9.616 11.816 9.648 11.848 ;
  LAYER M2 ;
        RECT 11.984 11.88 12.016 11.912 ;
  LAYER M2 ;
        RECT 9.616 11.944 9.648 11.976 ;
  LAYER M2 ;
        RECT 11.984 12.008 12.016 12.04 ;
  LAYER M2 ;
        RECT 9.616 12.072 9.648 12.104 ;
  LAYER M2 ;
        RECT 11.984 12.136 12.016 12.168 ;
  LAYER M2 ;
        RECT 9.616 12.2 9.648 12.232 ;
  LAYER M2 ;
        RECT 11.984 12.264 12.016 12.296 ;
  LAYER M2 ;
        RECT 9.616 12.328 9.648 12.36 ;
  LAYER M2 ;
        RECT 11.984 12.392 12.016 12.424 ;
  LAYER M2 ;
        RECT 9.616 12.456 9.648 12.488 ;
  LAYER M2 ;
        RECT 11.984 12.52 12.016 12.552 ;
  LAYER M2 ;
        RECT 9.616 12.584 9.648 12.616 ;
  LAYER M2 ;
        RECT 11.984 12.648 12.016 12.68 ;
  LAYER M2 ;
        RECT 9.616 12.712 9.648 12.744 ;
  LAYER M2 ;
        RECT 11.984 12.776 12.016 12.808 ;
  LAYER M2 ;
        RECT 9.616 12.84 9.648 12.872 ;
  LAYER M2 ;
        RECT 11.984 12.904 12.016 12.936 ;
  LAYER M2 ;
        RECT 9.616 12.968 9.648 13 ;
  LAYER M2 ;
        RECT 11.984 13.032 12.016 13.064 ;
  LAYER M2 ;
        RECT 9.616 13.096 9.648 13.128 ;
  LAYER M2 ;
        RECT 11.984 13.16 12.016 13.192 ;
  LAYER M2 ;
        RECT 9.616 13.224 9.648 13.256 ;
  LAYER M2 ;
        RECT 11.984 13.288 12.016 13.32 ;
  LAYER M2 ;
        RECT 9.616 13.352 9.648 13.384 ;
  LAYER M2 ;
        RECT 11.984 13.416 12.016 13.448 ;
  LAYER M2 ;
        RECT 9.616 13.48 9.648 13.512 ;
  LAYER M2 ;
        RECT 11.984 13.544 12.016 13.576 ;
  LAYER M2 ;
        RECT 9.568 11.172 12.064 13.776 ;
  LAYER M1 ;
        RECT 12.592 1.896 12.624 4.404 ;
  LAYER M3 ;
        RECT 12.592 4.352 12.624 4.384 ;
  LAYER M1 ;
        RECT 12.656 1.896 12.688 4.404 ;
  LAYER M3 ;
        RECT 12.656 1.916 12.688 1.948 ;
  LAYER M1 ;
        RECT 12.72 1.896 12.752 4.404 ;
  LAYER M3 ;
        RECT 12.72 4.352 12.752 4.384 ;
  LAYER M1 ;
        RECT 12.784 1.896 12.816 4.404 ;
  LAYER M3 ;
        RECT 12.784 1.916 12.816 1.948 ;
  LAYER M1 ;
        RECT 12.848 1.896 12.88 4.404 ;
  LAYER M3 ;
        RECT 12.848 4.352 12.88 4.384 ;
  LAYER M1 ;
        RECT 12.912 1.896 12.944 4.404 ;
  LAYER M3 ;
        RECT 12.912 1.916 12.944 1.948 ;
  LAYER M1 ;
        RECT 12.976 1.896 13.008 4.404 ;
  LAYER M3 ;
        RECT 12.976 4.352 13.008 4.384 ;
  LAYER M1 ;
        RECT 13.04 1.896 13.072 4.404 ;
  LAYER M3 ;
        RECT 13.04 1.916 13.072 1.948 ;
  LAYER M1 ;
        RECT 13.104 1.896 13.136 4.404 ;
  LAYER M3 ;
        RECT 13.104 4.352 13.136 4.384 ;
  LAYER M1 ;
        RECT 13.168 1.896 13.2 4.404 ;
  LAYER M3 ;
        RECT 13.168 1.916 13.2 1.948 ;
  LAYER M1 ;
        RECT 13.232 1.896 13.264 4.404 ;
  LAYER M3 ;
        RECT 13.232 4.352 13.264 4.384 ;
  LAYER M1 ;
        RECT 13.296 1.896 13.328 4.404 ;
  LAYER M3 ;
        RECT 13.296 1.916 13.328 1.948 ;
  LAYER M1 ;
        RECT 13.36 1.896 13.392 4.404 ;
  LAYER M3 ;
        RECT 13.36 4.352 13.392 4.384 ;
  LAYER M1 ;
        RECT 13.424 1.896 13.456 4.404 ;
  LAYER M3 ;
        RECT 13.424 1.916 13.456 1.948 ;
  LAYER M1 ;
        RECT 13.488 1.896 13.52 4.404 ;
  LAYER M3 ;
        RECT 13.488 4.352 13.52 4.384 ;
  LAYER M1 ;
        RECT 13.552 1.896 13.584 4.404 ;
  LAYER M3 ;
        RECT 13.552 1.916 13.584 1.948 ;
  LAYER M1 ;
        RECT 13.616 1.896 13.648 4.404 ;
  LAYER M3 ;
        RECT 13.616 4.352 13.648 4.384 ;
  LAYER M1 ;
        RECT 13.68 1.896 13.712 4.404 ;
  LAYER M3 ;
        RECT 13.68 1.916 13.712 1.948 ;
  LAYER M1 ;
        RECT 13.744 1.896 13.776 4.404 ;
  LAYER M3 ;
        RECT 13.744 4.352 13.776 4.384 ;
  LAYER M1 ;
        RECT 13.808 1.896 13.84 4.404 ;
  LAYER M3 ;
        RECT 13.808 1.916 13.84 1.948 ;
  LAYER M1 ;
        RECT 13.872 1.896 13.904 4.404 ;
  LAYER M3 ;
        RECT 13.872 4.352 13.904 4.384 ;
  LAYER M1 ;
        RECT 13.936 1.896 13.968 4.404 ;
  LAYER M3 ;
        RECT 13.936 1.916 13.968 1.948 ;
  LAYER M1 ;
        RECT 14 1.896 14.032 4.404 ;
  LAYER M3 ;
        RECT 14 4.352 14.032 4.384 ;
  LAYER M1 ;
        RECT 14.064 1.896 14.096 4.404 ;
  LAYER M3 ;
        RECT 14.064 1.916 14.096 1.948 ;
  LAYER M1 ;
        RECT 14.128 1.896 14.16 4.404 ;
  LAYER M3 ;
        RECT 14.128 4.352 14.16 4.384 ;
  LAYER M1 ;
        RECT 14.192 1.896 14.224 4.404 ;
  LAYER M3 ;
        RECT 14.192 1.916 14.224 1.948 ;
  LAYER M1 ;
        RECT 14.256 1.896 14.288 4.404 ;
  LAYER M3 ;
        RECT 14.256 4.352 14.288 4.384 ;
  LAYER M1 ;
        RECT 14.32 1.896 14.352 4.404 ;
  LAYER M3 ;
        RECT 14.32 1.916 14.352 1.948 ;
  LAYER M1 ;
        RECT 14.384 1.896 14.416 4.404 ;
  LAYER M3 ;
        RECT 14.384 4.352 14.416 4.384 ;
  LAYER M1 ;
        RECT 14.448 1.896 14.48 4.404 ;
  LAYER M3 ;
        RECT 14.448 1.916 14.48 1.948 ;
  LAYER M1 ;
        RECT 14.512 1.896 14.544 4.404 ;
  LAYER M3 ;
        RECT 14.512 4.352 14.544 4.384 ;
  LAYER M1 ;
        RECT 14.576 1.896 14.608 4.404 ;
  LAYER M3 ;
        RECT 14.576 1.916 14.608 1.948 ;
  LAYER M1 ;
        RECT 14.64 1.896 14.672 4.404 ;
  LAYER M3 ;
        RECT 14.64 4.352 14.672 4.384 ;
  LAYER M1 ;
        RECT 14.704 1.896 14.736 4.404 ;
  LAYER M3 ;
        RECT 14.704 1.916 14.736 1.948 ;
  LAYER M1 ;
        RECT 14.768 1.896 14.8 4.404 ;
  LAYER M3 ;
        RECT 14.768 4.352 14.8 4.384 ;
  LAYER M1 ;
        RECT 14.832 1.896 14.864 4.404 ;
  LAYER M3 ;
        RECT 14.832 1.916 14.864 1.948 ;
  LAYER M1 ;
        RECT 14.896 1.896 14.928 4.404 ;
  LAYER M3 ;
        RECT 14.896 4.352 14.928 4.384 ;
  LAYER M1 ;
        RECT 14.96 1.896 14.992 4.404 ;
  LAYER M3 ;
        RECT 12.592 1.98 12.624 2.012 ;
  LAYER M2 ;
        RECT 14.96 2.044 14.992 2.076 ;
  LAYER M2 ;
        RECT 12.592 2.108 12.624 2.14 ;
  LAYER M2 ;
        RECT 14.96 2.172 14.992 2.204 ;
  LAYER M2 ;
        RECT 12.592 2.236 12.624 2.268 ;
  LAYER M2 ;
        RECT 14.96 2.3 14.992 2.332 ;
  LAYER M2 ;
        RECT 12.592 2.364 12.624 2.396 ;
  LAYER M2 ;
        RECT 14.96 2.428 14.992 2.46 ;
  LAYER M2 ;
        RECT 12.592 2.492 12.624 2.524 ;
  LAYER M2 ;
        RECT 14.96 2.556 14.992 2.588 ;
  LAYER M2 ;
        RECT 12.592 2.62 12.624 2.652 ;
  LAYER M2 ;
        RECT 14.96 2.684 14.992 2.716 ;
  LAYER M2 ;
        RECT 12.592 2.748 12.624 2.78 ;
  LAYER M2 ;
        RECT 14.96 2.812 14.992 2.844 ;
  LAYER M2 ;
        RECT 12.592 2.876 12.624 2.908 ;
  LAYER M2 ;
        RECT 14.96 2.94 14.992 2.972 ;
  LAYER M2 ;
        RECT 12.592 3.004 12.624 3.036 ;
  LAYER M2 ;
        RECT 14.96 3.068 14.992 3.1 ;
  LAYER M2 ;
        RECT 12.592 3.132 12.624 3.164 ;
  LAYER M2 ;
        RECT 14.96 3.196 14.992 3.228 ;
  LAYER M2 ;
        RECT 12.592 3.26 12.624 3.292 ;
  LAYER M2 ;
        RECT 14.96 3.324 14.992 3.356 ;
  LAYER M2 ;
        RECT 12.592 3.388 12.624 3.42 ;
  LAYER M2 ;
        RECT 14.96 3.452 14.992 3.484 ;
  LAYER M2 ;
        RECT 12.592 3.516 12.624 3.548 ;
  LAYER M2 ;
        RECT 14.96 3.58 14.992 3.612 ;
  LAYER M2 ;
        RECT 12.592 3.644 12.624 3.676 ;
  LAYER M2 ;
        RECT 14.96 3.708 14.992 3.74 ;
  LAYER M2 ;
        RECT 12.592 3.772 12.624 3.804 ;
  LAYER M2 ;
        RECT 14.96 3.836 14.992 3.868 ;
  LAYER M2 ;
        RECT 12.592 3.9 12.624 3.932 ;
  LAYER M2 ;
        RECT 14.96 3.964 14.992 3.996 ;
  LAYER M2 ;
        RECT 12.592 4.028 12.624 4.06 ;
  LAYER M2 ;
        RECT 14.96 4.092 14.992 4.124 ;
  LAYER M2 ;
        RECT 12.592 4.156 12.624 4.188 ;
  LAYER M2 ;
        RECT 14.96 4.22 14.992 4.252 ;
  LAYER M2 ;
        RECT 12.544 1.848 15.04 4.452 ;
  LAYER M1 ;
        RECT 12.592 5.004 12.624 7.512 ;
  LAYER M3 ;
        RECT 12.592 7.46 12.624 7.492 ;
  LAYER M1 ;
        RECT 12.656 5.004 12.688 7.512 ;
  LAYER M3 ;
        RECT 12.656 5.024 12.688 5.056 ;
  LAYER M1 ;
        RECT 12.72 5.004 12.752 7.512 ;
  LAYER M3 ;
        RECT 12.72 7.46 12.752 7.492 ;
  LAYER M1 ;
        RECT 12.784 5.004 12.816 7.512 ;
  LAYER M3 ;
        RECT 12.784 5.024 12.816 5.056 ;
  LAYER M1 ;
        RECT 12.848 5.004 12.88 7.512 ;
  LAYER M3 ;
        RECT 12.848 7.46 12.88 7.492 ;
  LAYER M1 ;
        RECT 12.912 5.004 12.944 7.512 ;
  LAYER M3 ;
        RECT 12.912 5.024 12.944 5.056 ;
  LAYER M1 ;
        RECT 12.976 5.004 13.008 7.512 ;
  LAYER M3 ;
        RECT 12.976 7.46 13.008 7.492 ;
  LAYER M1 ;
        RECT 13.04 5.004 13.072 7.512 ;
  LAYER M3 ;
        RECT 13.04 5.024 13.072 5.056 ;
  LAYER M1 ;
        RECT 13.104 5.004 13.136 7.512 ;
  LAYER M3 ;
        RECT 13.104 7.46 13.136 7.492 ;
  LAYER M1 ;
        RECT 13.168 5.004 13.2 7.512 ;
  LAYER M3 ;
        RECT 13.168 5.024 13.2 5.056 ;
  LAYER M1 ;
        RECT 13.232 5.004 13.264 7.512 ;
  LAYER M3 ;
        RECT 13.232 7.46 13.264 7.492 ;
  LAYER M1 ;
        RECT 13.296 5.004 13.328 7.512 ;
  LAYER M3 ;
        RECT 13.296 5.024 13.328 5.056 ;
  LAYER M1 ;
        RECT 13.36 5.004 13.392 7.512 ;
  LAYER M3 ;
        RECT 13.36 7.46 13.392 7.492 ;
  LAYER M1 ;
        RECT 13.424 5.004 13.456 7.512 ;
  LAYER M3 ;
        RECT 13.424 5.024 13.456 5.056 ;
  LAYER M1 ;
        RECT 13.488 5.004 13.52 7.512 ;
  LAYER M3 ;
        RECT 13.488 7.46 13.52 7.492 ;
  LAYER M1 ;
        RECT 13.552 5.004 13.584 7.512 ;
  LAYER M3 ;
        RECT 13.552 5.024 13.584 5.056 ;
  LAYER M1 ;
        RECT 13.616 5.004 13.648 7.512 ;
  LAYER M3 ;
        RECT 13.616 7.46 13.648 7.492 ;
  LAYER M1 ;
        RECT 13.68 5.004 13.712 7.512 ;
  LAYER M3 ;
        RECT 13.68 5.024 13.712 5.056 ;
  LAYER M1 ;
        RECT 13.744 5.004 13.776 7.512 ;
  LAYER M3 ;
        RECT 13.744 7.46 13.776 7.492 ;
  LAYER M1 ;
        RECT 13.808 5.004 13.84 7.512 ;
  LAYER M3 ;
        RECT 13.808 5.024 13.84 5.056 ;
  LAYER M1 ;
        RECT 13.872 5.004 13.904 7.512 ;
  LAYER M3 ;
        RECT 13.872 7.46 13.904 7.492 ;
  LAYER M1 ;
        RECT 13.936 5.004 13.968 7.512 ;
  LAYER M3 ;
        RECT 13.936 5.024 13.968 5.056 ;
  LAYER M1 ;
        RECT 14 5.004 14.032 7.512 ;
  LAYER M3 ;
        RECT 14 7.46 14.032 7.492 ;
  LAYER M1 ;
        RECT 14.064 5.004 14.096 7.512 ;
  LAYER M3 ;
        RECT 14.064 5.024 14.096 5.056 ;
  LAYER M1 ;
        RECT 14.128 5.004 14.16 7.512 ;
  LAYER M3 ;
        RECT 14.128 7.46 14.16 7.492 ;
  LAYER M1 ;
        RECT 14.192 5.004 14.224 7.512 ;
  LAYER M3 ;
        RECT 14.192 5.024 14.224 5.056 ;
  LAYER M1 ;
        RECT 14.256 5.004 14.288 7.512 ;
  LAYER M3 ;
        RECT 14.256 7.46 14.288 7.492 ;
  LAYER M1 ;
        RECT 14.32 5.004 14.352 7.512 ;
  LAYER M3 ;
        RECT 14.32 5.024 14.352 5.056 ;
  LAYER M1 ;
        RECT 14.384 5.004 14.416 7.512 ;
  LAYER M3 ;
        RECT 14.384 7.46 14.416 7.492 ;
  LAYER M1 ;
        RECT 14.448 5.004 14.48 7.512 ;
  LAYER M3 ;
        RECT 14.448 5.024 14.48 5.056 ;
  LAYER M1 ;
        RECT 14.512 5.004 14.544 7.512 ;
  LAYER M3 ;
        RECT 14.512 7.46 14.544 7.492 ;
  LAYER M1 ;
        RECT 14.576 5.004 14.608 7.512 ;
  LAYER M3 ;
        RECT 14.576 5.024 14.608 5.056 ;
  LAYER M1 ;
        RECT 14.64 5.004 14.672 7.512 ;
  LAYER M3 ;
        RECT 14.64 7.46 14.672 7.492 ;
  LAYER M1 ;
        RECT 14.704 5.004 14.736 7.512 ;
  LAYER M3 ;
        RECT 14.704 5.024 14.736 5.056 ;
  LAYER M1 ;
        RECT 14.768 5.004 14.8 7.512 ;
  LAYER M3 ;
        RECT 14.768 7.46 14.8 7.492 ;
  LAYER M1 ;
        RECT 14.832 5.004 14.864 7.512 ;
  LAYER M3 ;
        RECT 14.832 5.024 14.864 5.056 ;
  LAYER M1 ;
        RECT 14.896 5.004 14.928 7.512 ;
  LAYER M3 ;
        RECT 14.896 7.46 14.928 7.492 ;
  LAYER M1 ;
        RECT 14.96 5.004 14.992 7.512 ;
  LAYER M3 ;
        RECT 12.592 5.088 12.624 5.12 ;
  LAYER M2 ;
        RECT 14.96 5.152 14.992 5.184 ;
  LAYER M2 ;
        RECT 12.592 5.216 12.624 5.248 ;
  LAYER M2 ;
        RECT 14.96 5.28 14.992 5.312 ;
  LAYER M2 ;
        RECT 12.592 5.344 12.624 5.376 ;
  LAYER M2 ;
        RECT 14.96 5.408 14.992 5.44 ;
  LAYER M2 ;
        RECT 12.592 5.472 12.624 5.504 ;
  LAYER M2 ;
        RECT 14.96 5.536 14.992 5.568 ;
  LAYER M2 ;
        RECT 12.592 5.6 12.624 5.632 ;
  LAYER M2 ;
        RECT 14.96 5.664 14.992 5.696 ;
  LAYER M2 ;
        RECT 12.592 5.728 12.624 5.76 ;
  LAYER M2 ;
        RECT 14.96 5.792 14.992 5.824 ;
  LAYER M2 ;
        RECT 12.592 5.856 12.624 5.888 ;
  LAYER M2 ;
        RECT 14.96 5.92 14.992 5.952 ;
  LAYER M2 ;
        RECT 12.592 5.984 12.624 6.016 ;
  LAYER M2 ;
        RECT 14.96 6.048 14.992 6.08 ;
  LAYER M2 ;
        RECT 12.592 6.112 12.624 6.144 ;
  LAYER M2 ;
        RECT 14.96 6.176 14.992 6.208 ;
  LAYER M2 ;
        RECT 12.592 6.24 12.624 6.272 ;
  LAYER M2 ;
        RECT 14.96 6.304 14.992 6.336 ;
  LAYER M2 ;
        RECT 12.592 6.368 12.624 6.4 ;
  LAYER M2 ;
        RECT 14.96 6.432 14.992 6.464 ;
  LAYER M2 ;
        RECT 12.592 6.496 12.624 6.528 ;
  LAYER M2 ;
        RECT 14.96 6.56 14.992 6.592 ;
  LAYER M2 ;
        RECT 12.592 6.624 12.624 6.656 ;
  LAYER M2 ;
        RECT 14.96 6.688 14.992 6.72 ;
  LAYER M2 ;
        RECT 12.592 6.752 12.624 6.784 ;
  LAYER M2 ;
        RECT 14.96 6.816 14.992 6.848 ;
  LAYER M2 ;
        RECT 12.592 6.88 12.624 6.912 ;
  LAYER M2 ;
        RECT 14.96 6.944 14.992 6.976 ;
  LAYER M2 ;
        RECT 12.592 7.008 12.624 7.04 ;
  LAYER M2 ;
        RECT 14.96 7.072 14.992 7.104 ;
  LAYER M2 ;
        RECT 12.592 7.136 12.624 7.168 ;
  LAYER M2 ;
        RECT 14.96 7.2 14.992 7.232 ;
  LAYER M2 ;
        RECT 12.592 7.264 12.624 7.296 ;
  LAYER M2 ;
        RECT 14.96 7.328 14.992 7.36 ;
  LAYER M2 ;
        RECT 12.544 4.956 15.04 7.56 ;
  LAYER M1 ;
        RECT 12.592 8.112 12.624 10.62 ;
  LAYER M3 ;
        RECT 12.592 10.568 12.624 10.6 ;
  LAYER M1 ;
        RECT 12.656 8.112 12.688 10.62 ;
  LAYER M3 ;
        RECT 12.656 8.132 12.688 8.164 ;
  LAYER M1 ;
        RECT 12.72 8.112 12.752 10.62 ;
  LAYER M3 ;
        RECT 12.72 10.568 12.752 10.6 ;
  LAYER M1 ;
        RECT 12.784 8.112 12.816 10.62 ;
  LAYER M3 ;
        RECT 12.784 8.132 12.816 8.164 ;
  LAYER M1 ;
        RECT 12.848 8.112 12.88 10.62 ;
  LAYER M3 ;
        RECT 12.848 10.568 12.88 10.6 ;
  LAYER M1 ;
        RECT 12.912 8.112 12.944 10.62 ;
  LAYER M3 ;
        RECT 12.912 8.132 12.944 8.164 ;
  LAYER M1 ;
        RECT 12.976 8.112 13.008 10.62 ;
  LAYER M3 ;
        RECT 12.976 10.568 13.008 10.6 ;
  LAYER M1 ;
        RECT 13.04 8.112 13.072 10.62 ;
  LAYER M3 ;
        RECT 13.04 8.132 13.072 8.164 ;
  LAYER M1 ;
        RECT 13.104 8.112 13.136 10.62 ;
  LAYER M3 ;
        RECT 13.104 10.568 13.136 10.6 ;
  LAYER M1 ;
        RECT 13.168 8.112 13.2 10.62 ;
  LAYER M3 ;
        RECT 13.168 8.132 13.2 8.164 ;
  LAYER M1 ;
        RECT 13.232 8.112 13.264 10.62 ;
  LAYER M3 ;
        RECT 13.232 10.568 13.264 10.6 ;
  LAYER M1 ;
        RECT 13.296 8.112 13.328 10.62 ;
  LAYER M3 ;
        RECT 13.296 8.132 13.328 8.164 ;
  LAYER M1 ;
        RECT 13.36 8.112 13.392 10.62 ;
  LAYER M3 ;
        RECT 13.36 10.568 13.392 10.6 ;
  LAYER M1 ;
        RECT 13.424 8.112 13.456 10.62 ;
  LAYER M3 ;
        RECT 13.424 8.132 13.456 8.164 ;
  LAYER M1 ;
        RECT 13.488 8.112 13.52 10.62 ;
  LAYER M3 ;
        RECT 13.488 10.568 13.52 10.6 ;
  LAYER M1 ;
        RECT 13.552 8.112 13.584 10.62 ;
  LAYER M3 ;
        RECT 13.552 8.132 13.584 8.164 ;
  LAYER M1 ;
        RECT 13.616 8.112 13.648 10.62 ;
  LAYER M3 ;
        RECT 13.616 10.568 13.648 10.6 ;
  LAYER M1 ;
        RECT 13.68 8.112 13.712 10.62 ;
  LAYER M3 ;
        RECT 13.68 8.132 13.712 8.164 ;
  LAYER M1 ;
        RECT 13.744 8.112 13.776 10.62 ;
  LAYER M3 ;
        RECT 13.744 10.568 13.776 10.6 ;
  LAYER M1 ;
        RECT 13.808 8.112 13.84 10.62 ;
  LAYER M3 ;
        RECT 13.808 8.132 13.84 8.164 ;
  LAYER M1 ;
        RECT 13.872 8.112 13.904 10.62 ;
  LAYER M3 ;
        RECT 13.872 10.568 13.904 10.6 ;
  LAYER M1 ;
        RECT 13.936 8.112 13.968 10.62 ;
  LAYER M3 ;
        RECT 13.936 8.132 13.968 8.164 ;
  LAYER M1 ;
        RECT 14 8.112 14.032 10.62 ;
  LAYER M3 ;
        RECT 14 10.568 14.032 10.6 ;
  LAYER M1 ;
        RECT 14.064 8.112 14.096 10.62 ;
  LAYER M3 ;
        RECT 14.064 8.132 14.096 8.164 ;
  LAYER M1 ;
        RECT 14.128 8.112 14.16 10.62 ;
  LAYER M3 ;
        RECT 14.128 10.568 14.16 10.6 ;
  LAYER M1 ;
        RECT 14.192 8.112 14.224 10.62 ;
  LAYER M3 ;
        RECT 14.192 8.132 14.224 8.164 ;
  LAYER M1 ;
        RECT 14.256 8.112 14.288 10.62 ;
  LAYER M3 ;
        RECT 14.256 10.568 14.288 10.6 ;
  LAYER M1 ;
        RECT 14.32 8.112 14.352 10.62 ;
  LAYER M3 ;
        RECT 14.32 8.132 14.352 8.164 ;
  LAYER M1 ;
        RECT 14.384 8.112 14.416 10.62 ;
  LAYER M3 ;
        RECT 14.384 10.568 14.416 10.6 ;
  LAYER M1 ;
        RECT 14.448 8.112 14.48 10.62 ;
  LAYER M3 ;
        RECT 14.448 8.132 14.48 8.164 ;
  LAYER M1 ;
        RECT 14.512 8.112 14.544 10.62 ;
  LAYER M3 ;
        RECT 14.512 10.568 14.544 10.6 ;
  LAYER M1 ;
        RECT 14.576 8.112 14.608 10.62 ;
  LAYER M3 ;
        RECT 14.576 8.132 14.608 8.164 ;
  LAYER M1 ;
        RECT 14.64 8.112 14.672 10.62 ;
  LAYER M3 ;
        RECT 14.64 10.568 14.672 10.6 ;
  LAYER M1 ;
        RECT 14.704 8.112 14.736 10.62 ;
  LAYER M3 ;
        RECT 14.704 8.132 14.736 8.164 ;
  LAYER M1 ;
        RECT 14.768 8.112 14.8 10.62 ;
  LAYER M3 ;
        RECT 14.768 10.568 14.8 10.6 ;
  LAYER M1 ;
        RECT 14.832 8.112 14.864 10.62 ;
  LAYER M3 ;
        RECT 14.832 8.132 14.864 8.164 ;
  LAYER M1 ;
        RECT 14.896 8.112 14.928 10.62 ;
  LAYER M3 ;
        RECT 14.896 10.568 14.928 10.6 ;
  LAYER M1 ;
        RECT 14.96 8.112 14.992 10.62 ;
  LAYER M3 ;
        RECT 12.592 8.196 12.624 8.228 ;
  LAYER M2 ;
        RECT 14.96 8.26 14.992 8.292 ;
  LAYER M2 ;
        RECT 12.592 8.324 12.624 8.356 ;
  LAYER M2 ;
        RECT 14.96 8.388 14.992 8.42 ;
  LAYER M2 ;
        RECT 12.592 8.452 12.624 8.484 ;
  LAYER M2 ;
        RECT 14.96 8.516 14.992 8.548 ;
  LAYER M2 ;
        RECT 12.592 8.58 12.624 8.612 ;
  LAYER M2 ;
        RECT 14.96 8.644 14.992 8.676 ;
  LAYER M2 ;
        RECT 12.592 8.708 12.624 8.74 ;
  LAYER M2 ;
        RECT 14.96 8.772 14.992 8.804 ;
  LAYER M2 ;
        RECT 12.592 8.836 12.624 8.868 ;
  LAYER M2 ;
        RECT 14.96 8.9 14.992 8.932 ;
  LAYER M2 ;
        RECT 12.592 8.964 12.624 8.996 ;
  LAYER M2 ;
        RECT 14.96 9.028 14.992 9.06 ;
  LAYER M2 ;
        RECT 12.592 9.092 12.624 9.124 ;
  LAYER M2 ;
        RECT 14.96 9.156 14.992 9.188 ;
  LAYER M2 ;
        RECT 12.592 9.22 12.624 9.252 ;
  LAYER M2 ;
        RECT 14.96 9.284 14.992 9.316 ;
  LAYER M2 ;
        RECT 12.592 9.348 12.624 9.38 ;
  LAYER M2 ;
        RECT 14.96 9.412 14.992 9.444 ;
  LAYER M2 ;
        RECT 12.592 9.476 12.624 9.508 ;
  LAYER M2 ;
        RECT 14.96 9.54 14.992 9.572 ;
  LAYER M2 ;
        RECT 12.592 9.604 12.624 9.636 ;
  LAYER M2 ;
        RECT 14.96 9.668 14.992 9.7 ;
  LAYER M2 ;
        RECT 12.592 9.732 12.624 9.764 ;
  LAYER M2 ;
        RECT 14.96 9.796 14.992 9.828 ;
  LAYER M2 ;
        RECT 12.592 9.86 12.624 9.892 ;
  LAYER M2 ;
        RECT 14.96 9.924 14.992 9.956 ;
  LAYER M2 ;
        RECT 12.592 9.988 12.624 10.02 ;
  LAYER M2 ;
        RECT 14.96 10.052 14.992 10.084 ;
  LAYER M2 ;
        RECT 12.592 10.116 12.624 10.148 ;
  LAYER M2 ;
        RECT 14.96 10.18 14.992 10.212 ;
  LAYER M2 ;
        RECT 12.592 10.244 12.624 10.276 ;
  LAYER M2 ;
        RECT 14.96 10.308 14.992 10.34 ;
  LAYER M2 ;
        RECT 12.592 10.372 12.624 10.404 ;
  LAYER M2 ;
        RECT 14.96 10.436 14.992 10.468 ;
  LAYER M2 ;
        RECT 12.544 8.064 15.04 10.668 ;
  LAYER M1 ;
        RECT 12.592 11.22 12.624 13.728 ;
  LAYER M3 ;
        RECT 12.592 13.676 12.624 13.708 ;
  LAYER M1 ;
        RECT 12.656 11.22 12.688 13.728 ;
  LAYER M3 ;
        RECT 12.656 11.24 12.688 11.272 ;
  LAYER M1 ;
        RECT 12.72 11.22 12.752 13.728 ;
  LAYER M3 ;
        RECT 12.72 13.676 12.752 13.708 ;
  LAYER M1 ;
        RECT 12.784 11.22 12.816 13.728 ;
  LAYER M3 ;
        RECT 12.784 11.24 12.816 11.272 ;
  LAYER M1 ;
        RECT 12.848 11.22 12.88 13.728 ;
  LAYER M3 ;
        RECT 12.848 13.676 12.88 13.708 ;
  LAYER M1 ;
        RECT 12.912 11.22 12.944 13.728 ;
  LAYER M3 ;
        RECT 12.912 11.24 12.944 11.272 ;
  LAYER M1 ;
        RECT 12.976 11.22 13.008 13.728 ;
  LAYER M3 ;
        RECT 12.976 13.676 13.008 13.708 ;
  LAYER M1 ;
        RECT 13.04 11.22 13.072 13.728 ;
  LAYER M3 ;
        RECT 13.04 11.24 13.072 11.272 ;
  LAYER M1 ;
        RECT 13.104 11.22 13.136 13.728 ;
  LAYER M3 ;
        RECT 13.104 13.676 13.136 13.708 ;
  LAYER M1 ;
        RECT 13.168 11.22 13.2 13.728 ;
  LAYER M3 ;
        RECT 13.168 11.24 13.2 11.272 ;
  LAYER M1 ;
        RECT 13.232 11.22 13.264 13.728 ;
  LAYER M3 ;
        RECT 13.232 13.676 13.264 13.708 ;
  LAYER M1 ;
        RECT 13.296 11.22 13.328 13.728 ;
  LAYER M3 ;
        RECT 13.296 11.24 13.328 11.272 ;
  LAYER M1 ;
        RECT 13.36 11.22 13.392 13.728 ;
  LAYER M3 ;
        RECT 13.36 13.676 13.392 13.708 ;
  LAYER M1 ;
        RECT 13.424 11.22 13.456 13.728 ;
  LAYER M3 ;
        RECT 13.424 11.24 13.456 11.272 ;
  LAYER M1 ;
        RECT 13.488 11.22 13.52 13.728 ;
  LAYER M3 ;
        RECT 13.488 13.676 13.52 13.708 ;
  LAYER M1 ;
        RECT 13.552 11.22 13.584 13.728 ;
  LAYER M3 ;
        RECT 13.552 11.24 13.584 11.272 ;
  LAYER M1 ;
        RECT 13.616 11.22 13.648 13.728 ;
  LAYER M3 ;
        RECT 13.616 13.676 13.648 13.708 ;
  LAYER M1 ;
        RECT 13.68 11.22 13.712 13.728 ;
  LAYER M3 ;
        RECT 13.68 11.24 13.712 11.272 ;
  LAYER M1 ;
        RECT 13.744 11.22 13.776 13.728 ;
  LAYER M3 ;
        RECT 13.744 13.676 13.776 13.708 ;
  LAYER M1 ;
        RECT 13.808 11.22 13.84 13.728 ;
  LAYER M3 ;
        RECT 13.808 11.24 13.84 11.272 ;
  LAYER M1 ;
        RECT 13.872 11.22 13.904 13.728 ;
  LAYER M3 ;
        RECT 13.872 13.676 13.904 13.708 ;
  LAYER M1 ;
        RECT 13.936 11.22 13.968 13.728 ;
  LAYER M3 ;
        RECT 13.936 11.24 13.968 11.272 ;
  LAYER M1 ;
        RECT 14 11.22 14.032 13.728 ;
  LAYER M3 ;
        RECT 14 13.676 14.032 13.708 ;
  LAYER M1 ;
        RECT 14.064 11.22 14.096 13.728 ;
  LAYER M3 ;
        RECT 14.064 11.24 14.096 11.272 ;
  LAYER M1 ;
        RECT 14.128 11.22 14.16 13.728 ;
  LAYER M3 ;
        RECT 14.128 13.676 14.16 13.708 ;
  LAYER M1 ;
        RECT 14.192 11.22 14.224 13.728 ;
  LAYER M3 ;
        RECT 14.192 11.24 14.224 11.272 ;
  LAYER M1 ;
        RECT 14.256 11.22 14.288 13.728 ;
  LAYER M3 ;
        RECT 14.256 13.676 14.288 13.708 ;
  LAYER M1 ;
        RECT 14.32 11.22 14.352 13.728 ;
  LAYER M3 ;
        RECT 14.32 11.24 14.352 11.272 ;
  LAYER M1 ;
        RECT 14.384 11.22 14.416 13.728 ;
  LAYER M3 ;
        RECT 14.384 13.676 14.416 13.708 ;
  LAYER M1 ;
        RECT 14.448 11.22 14.48 13.728 ;
  LAYER M3 ;
        RECT 14.448 11.24 14.48 11.272 ;
  LAYER M1 ;
        RECT 14.512 11.22 14.544 13.728 ;
  LAYER M3 ;
        RECT 14.512 13.676 14.544 13.708 ;
  LAYER M1 ;
        RECT 14.576 11.22 14.608 13.728 ;
  LAYER M3 ;
        RECT 14.576 11.24 14.608 11.272 ;
  LAYER M1 ;
        RECT 14.64 11.22 14.672 13.728 ;
  LAYER M3 ;
        RECT 14.64 13.676 14.672 13.708 ;
  LAYER M1 ;
        RECT 14.704 11.22 14.736 13.728 ;
  LAYER M3 ;
        RECT 14.704 11.24 14.736 11.272 ;
  LAYER M1 ;
        RECT 14.768 11.22 14.8 13.728 ;
  LAYER M3 ;
        RECT 14.768 13.676 14.8 13.708 ;
  LAYER M1 ;
        RECT 14.832 11.22 14.864 13.728 ;
  LAYER M3 ;
        RECT 14.832 11.24 14.864 11.272 ;
  LAYER M1 ;
        RECT 14.896 11.22 14.928 13.728 ;
  LAYER M3 ;
        RECT 14.896 13.676 14.928 13.708 ;
  LAYER M1 ;
        RECT 14.96 11.22 14.992 13.728 ;
  LAYER M3 ;
        RECT 12.592 11.304 12.624 11.336 ;
  LAYER M2 ;
        RECT 14.96 11.368 14.992 11.4 ;
  LAYER M2 ;
        RECT 12.592 11.432 12.624 11.464 ;
  LAYER M2 ;
        RECT 14.96 11.496 14.992 11.528 ;
  LAYER M2 ;
        RECT 12.592 11.56 12.624 11.592 ;
  LAYER M2 ;
        RECT 14.96 11.624 14.992 11.656 ;
  LAYER M2 ;
        RECT 12.592 11.688 12.624 11.72 ;
  LAYER M2 ;
        RECT 14.96 11.752 14.992 11.784 ;
  LAYER M2 ;
        RECT 12.592 11.816 12.624 11.848 ;
  LAYER M2 ;
        RECT 14.96 11.88 14.992 11.912 ;
  LAYER M2 ;
        RECT 12.592 11.944 12.624 11.976 ;
  LAYER M2 ;
        RECT 14.96 12.008 14.992 12.04 ;
  LAYER M2 ;
        RECT 12.592 12.072 12.624 12.104 ;
  LAYER M2 ;
        RECT 14.96 12.136 14.992 12.168 ;
  LAYER M2 ;
        RECT 12.592 12.2 12.624 12.232 ;
  LAYER M2 ;
        RECT 14.96 12.264 14.992 12.296 ;
  LAYER M2 ;
        RECT 12.592 12.328 12.624 12.36 ;
  LAYER M2 ;
        RECT 14.96 12.392 14.992 12.424 ;
  LAYER M2 ;
        RECT 12.592 12.456 12.624 12.488 ;
  LAYER M2 ;
        RECT 14.96 12.52 14.992 12.552 ;
  LAYER M2 ;
        RECT 12.592 12.584 12.624 12.616 ;
  LAYER M2 ;
        RECT 14.96 12.648 14.992 12.68 ;
  LAYER M2 ;
        RECT 12.592 12.712 12.624 12.744 ;
  LAYER M2 ;
        RECT 14.96 12.776 14.992 12.808 ;
  LAYER M2 ;
        RECT 12.592 12.84 12.624 12.872 ;
  LAYER M2 ;
        RECT 14.96 12.904 14.992 12.936 ;
  LAYER M2 ;
        RECT 12.592 12.968 12.624 13 ;
  LAYER M2 ;
        RECT 14.96 13.032 14.992 13.064 ;
  LAYER M2 ;
        RECT 12.592 13.096 12.624 13.128 ;
  LAYER M2 ;
        RECT 14.96 13.16 14.992 13.192 ;
  LAYER M2 ;
        RECT 12.592 13.224 12.624 13.256 ;
  LAYER M2 ;
        RECT 14.96 13.288 14.992 13.32 ;
  LAYER M2 ;
        RECT 12.592 13.352 12.624 13.384 ;
  LAYER M2 ;
        RECT 14.96 13.416 14.992 13.448 ;
  LAYER M2 ;
        RECT 12.592 13.48 12.624 13.512 ;
  LAYER M2 ;
        RECT 14.96 13.544 14.992 13.576 ;
  LAYER M2 ;
        RECT 12.544 11.172 15.04 13.776 ;
  LAYER M1 ;
        RECT 5.344 0.216 5.376 0.876 ;
  LAYER M1 ;
        RECT 5.264 0.216 5.296 0.876 ;
  LAYER M1 ;
        RECT 5.424 0.656 5.456 0.688 ;
  LAYER M1 ;
        RECT 15.664 0.216 15.696 0.876 ;
  LAYER M1 ;
        RECT 15.744 0.216 15.776 0.876 ;
  LAYER M1 ;
        RECT 15.584 0.656 15.616 0.688 ;
  LAYER M1 ;
        RECT 6.704 0.3 6.736 0.96 ;
  LAYER M1 ;
        RECT 6.064 0.3 6.096 0.96 ;
  LAYER M1 ;
        RECT 6.784 0.3 6.816 0.96 ;
  LAYER M1 ;
        RECT 6.144 0.3 6.176 0.96 ;
  LAYER M1 ;
        RECT 6.624 0.3 6.656 0.96 ;
  LAYER M1 ;
        RECT 5.984 0.488 6.016 0.52 ;
  LAYER M1 ;
        RECT 8.064 0.3 8.096 0.96 ;
  LAYER M1 ;
        RECT 7.424 0.3 7.456 0.96 ;
  LAYER M1 ;
        RECT 8.144 0.3 8.176 0.96 ;
  LAYER M1 ;
        RECT 7.504 0.3 7.536 0.96 ;
  LAYER M1 ;
        RECT 7.984 0.3 8.016 0.96 ;
  LAYER M1 ;
        RECT 7.344 0.488 7.376 0.52 ;
  LAYER M1 ;
        RECT 6.56 24.24 6.592 24.312 ;
  LAYER M2 ;
        RECT 6.54 24.26 6.612 24.292 ;
  LAYER M2 ;
        RECT 6.576 24.26 9.328 24.292 ;
  LAYER M1 ;
        RECT 9.312 24.24 9.344 24.312 ;
  LAYER M2 ;
        RECT 9.292 24.26 9.364 24.292 ;
  LAYER M1 ;
        RECT 9.536 21.132 9.568 21.204 ;
  LAYER M2 ;
        RECT 9.516 21.152 9.588 21.184 ;
  LAYER M1 ;
        RECT 9.536 21.168 9.568 21.336 ;
  LAYER M1 ;
        RECT 9.536 21.3 9.568 21.372 ;
  LAYER M2 ;
        RECT 9.516 21.32 9.588 21.352 ;
  LAYER M2 ;
        RECT 9.328 21.32 9.552 21.352 ;
  LAYER M1 ;
        RECT 9.312 21.3 9.344 21.372 ;
  LAYER M2 ;
        RECT 9.292 21.32 9.364 21.352 ;
  LAYER M1 ;
        RECT 9.312 31.044 9.344 31.116 ;
  LAYER M2 ;
        RECT 9.292 31.064 9.364 31.096 ;
  LAYER M1 ;
        RECT 9.312 30.828 9.344 31.08 ;
  LAYER M1 ;
        RECT 9.312 21.336 9.344 30.828 ;
  LAYER M1 ;
        RECT 3.584 27.348 3.616 27.42 ;
  LAYER M2 ;
        RECT 3.564 27.368 3.636 27.4 ;
  LAYER M2 ;
        RECT 3.6 27.368 6.352 27.4 ;
  LAYER M1 ;
        RECT 6.336 27.348 6.368 27.42 ;
  LAYER M2 ;
        RECT 6.316 27.368 6.388 27.4 ;
  LAYER M1 ;
        RECT 6.336 31.044 6.368 31.116 ;
  LAYER M2 ;
        RECT 6.316 31.064 6.388 31.096 ;
  LAYER M1 ;
        RECT 6.336 30.828 6.368 31.08 ;
  LAYER M1 ;
        RECT 6.336 27.384 6.368 30.828 ;
  LAYER M2 ;
        RECT 6.352 31.064 9.328 31.096 ;
  LAYER M1 ;
        RECT 9.536 24.24 9.568 24.312 ;
  LAYER M2 ;
        RECT 9.516 24.26 9.588 24.292 ;
  LAYER M2 ;
        RECT 9.552 24.26 12.304 24.292 ;
  LAYER M1 ;
        RECT 12.288 24.24 12.32 24.312 ;
  LAYER M2 ;
        RECT 12.268 24.26 12.34 24.292 ;
  LAYER M1 ;
        RECT 9.536 27.348 9.568 27.42 ;
  LAYER M2 ;
        RECT 9.516 27.368 9.588 27.4 ;
  LAYER M2 ;
        RECT 9.552 27.368 12.304 27.4 ;
  LAYER M1 ;
        RECT 12.288 27.348 12.32 27.42 ;
  LAYER M2 ;
        RECT 12.268 27.368 12.34 27.4 ;
  LAYER M1 ;
        RECT 12.288 31.212 12.32 31.284 ;
  LAYER M2 ;
        RECT 12.268 31.232 12.34 31.264 ;
  LAYER M1 ;
        RECT 12.288 30.828 12.32 31.248 ;
  LAYER M1 ;
        RECT 12.288 24.276 12.32 30.828 ;
  LAYER M1 ;
        RECT 3.584 24.24 3.616 24.312 ;
  LAYER M2 ;
        RECT 3.564 24.26 3.636 24.292 ;
  LAYER M1 ;
        RECT 3.584 24.276 3.616 24.444 ;
  LAYER M1 ;
        RECT 3.584 24.408 3.616 24.48 ;
  LAYER M2 ;
        RECT 3.564 24.428 3.636 24.46 ;
  LAYER M2 ;
        RECT 3.376 24.428 3.6 24.46 ;
  LAYER M1 ;
        RECT 3.36 24.408 3.392 24.48 ;
  LAYER M2 ;
        RECT 3.34 24.428 3.412 24.46 ;
  LAYER M1 ;
        RECT 3.584 21.132 3.616 21.204 ;
  LAYER M2 ;
        RECT 3.564 21.152 3.636 21.184 ;
  LAYER M1 ;
        RECT 3.584 21.168 3.616 21.336 ;
  LAYER M1 ;
        RECT 3.584 21.3 3.616 21.372 ;
  LAYER M2 ;
        RECT 3.564 21.32 3.636 21.352 ;
  LAYER M2 ;
        RECT 3.376 21.32 3.6 21.352 ;
  LAYER M1 ;
        RECT 3.36 21.3 3.392 21.372 ;
  LAYER M2 ;
        RECT 3.34 21.32 3.412 21.352 ;
  LAYER M1 ;
        RECT 3.36 31.212 3.392 31.284 ;
  LAYER M2 ;
        RECT 3.34 31.232 3.412 31.264 ;
  LAYER M1 ;
        RECT 3.36 30.828 3.392 31.248 ;
  LAYER M1 ;
        RECT 3.36 21.336 3.392 30.828 ;
  LAYER M2 ;
        RECT 3.376 31.232 12.304 31.264 ;
  LAYER M1 ;
        RECT 6.56 27.348 6.592 27.42 ;
  LAYER M2 ;
        RECT 6.54 27.368 6.612 27.4 ;
  LAYER M2 ;
        RECT 6.576 27.368 9.552 27.4 ;
  LAYER M1 ;
        RECT 9.536 27.348 9.568 27.42 ;
  LAYER M2 ;
        RECT 9.516 27.368 9.588 27.4 ;
  LAYER M1 ;
        RECT 6.56 21.132 6.592 21.204 ;
  LAYER M2 ;
        RECT 6.54 21.152 6.612 21.184 ;
  LAYER M2 ;
        RECT 3.6 21.152 6.576 21.184 ;
  LAYER M1 ;
        RECT 3.584 21.132 3.616 21.204 ;
  LAYER M2 ;
        RECT 3.564 21.152 3.636 21.184 ;
  LAYER M1 ;
        RECT 12.512 30.456 12.544 30.528 ;
  LAYER M2 ;
        RECT 12.492 30.476 12.564 30.508 ;
  LAYER M2 ;
        RECT 12.528 30.476 15.28 30.508 ;
  LAYER M1 ;
        RECT 15.264 30.456 15.296 30.528 ;
  LAYER M2 ;
        RECT 15.244 30.476 15.316 30.508 ;
  LAYER M1 ;
        RECT 12.512 27.348 12.544 27.42 ;
  LAYER M2 ;
        RECT 12.492 27.368 12.564 27.4 ;
  LAYER M2 ;
        RECT 12.528 27.368 15.28 27.4 ;
  LAYER M1 ;
        RECT 15.264 27.348 15.296 27.42 ;
  LAYER M2 ;
        RECT 15.244 27.368 15.316 27.4 ;
  LAYER M1 ;
        RECT 12.512 24.24 12.544 24.312 ;
  LAYER M2 ;
        RECT 12.492 24.26 12.564 24.292 ;
  LAYER M2 ;
        RECT 12.528 24.26 15.28 24.292 ;
  LAYER M1 ;
        RECT 15.264 24.24 15.296 24.312 ;
  LAYER M2 ;
        RECT 15.244 24.26 15.316 24.292 ;
  LAYER M1 ;
        RECT 12.512 21.132 12.544 21.204 ;
  LAYER M2 ;
        RECT 12.492 21.152 12.564 21.184 ;
  LAYER M2 ;
        RECT 12.528 21.152 15.28 21.184 ;
  LAYER M1 ;
        RECT 15.264 21.132 15.296 21.204 ;
  LAYER M2 ;
        RECT 15.244 21.152 15.316 21.184 ;
  LAYER M1 ;
        RECT 12.512 18.024 12.544 18.096 ;
  LAYER M2 ;
        RECT 12.492 18.044 12.564 18.076 ;
  LAYER M2 ;
        RECT 12.528 18.044 15.28 18.076 ;
  LAYER M1 ;
        RECT 15.264 18.024 15.296 18.096 ;
  LAYER M2 ;
        RECT 15.244 18.044 15.316 18.076 ;
  LAYER M1 ;
        RECT 15.264 31.38 15.296 31.452 ;
  LAYER M2 ;
        RECT 15.244 31.4 15.316 31.432 ;
  LAYER M1 ;
        RECT 15.264 30.828 15.296 31.416 ;
  LAYER M1 ;
        RECT 15.264 18.06 15.296 30.828 ;
  LAYER M1 ;
        RECT 0.608 30.456 0.64 30.528 ;
  LAYER M2 ;
        RECT 0.588 30.476 0.66 30.508 ;
  LAYER M1 ;
        RECT 0.608 30.492 0.64 30.66 ;
  LAYER M1 ;
        RECT 0.608 30.624 0.64 30.696 ;
  LAYER M2 ;
        RECT 0.588 30.644 0.66 30.676 ;
  LAYER M2 ;
        RECT 0.4 30.644 0.624 30.676 ;
  LAYER M1 ;
        RECT 0.384 30.624 0.416 30.696 ;
  LAYER M2 ;
        RECT 0.364 30.644 0.436 30.676 ;
  LAYER M1 ;
        RECT 0.608 27.348 0.64 27.42 ;
  LAYER M2 ;
        RECT 0.588 27.368 0.66 27.4 ;
  LAYER M1 ;
        RECT 0.608 27.384 0.64 27.552 ;
  LAYER M1 ;
        RECT 0.608 27.516 0.64 27.588 ;
  LAYER M2 ;
        RECT 0.588 27.536 0.66 27.568 ;
  LAYER M2 ;
        RECT 0.4 27.536 0.624 27.568 ;
  LAYER M1 ;
        RECT 0.384 27.516 0.416 27.588 ;
  LAYER M2 ;
        RECT 0.364 27.536 0.436 27.568 ;
  LAYER M1 ;
        RECT 0.608 24.24 0.64 24.312 ;
  LAYER M2 ;
        RECT 0.588 24.26 0.66 24.292 ;
  LAYER M1 ;
        RECT 0.608 24.276 0.64 24.444 ;
  LAYER M1 ;
        RECT 0.608 24.408 0.64 24.48 ;
  LAYER M2 ;
        RECT 0.588 24.428 0.66 24.46 ;
  LAYER M2 ;
        RECT 0.4 24.428 0.624 24.46 ;
  LAYER M1 ;
        RECT 0.384 24.408 0.416 24.48 ;
  LAYER M2 ;
        RECT 0.364 24.428 0.436 24.46 ;
  LAYER M1 ;
        RECT 0.608 21.132 0.64 21.204 ;
  LAYER M2 ;
        RECT 0.588 21.152 0.66 21.184 ;
  LAYER M1 ;
        RECT 0.608 21.168 0.64 21.336 ;
  LAYER M1 ;
        RECT 0.608 21.3 0.64 21.372 ;
  LAYER M2 ;
        RECT 0.588 21.32 0.66 21.352 ;
  LAYER M2 ;
        RECT 0.4 21.32 0.624 21.352 ;
  LAYER M1 ;
        RECT 0.384 21.3 0.416 21.372 ;
  LAYER M2 ;
        RECT 0.364 21.32 0.436 21.352 ;
  LAYER M1 ;
        RECT 0.608 18.024 0.64 18.096 ;
  LAYER M2 ;
        RECT 0.588 18.044 0.66 18.076 ;
  LAYER M1 ;
        RECT 0.608 18.06 0.64 18.228 ;
  LAYER M1 ;
        RECT 0.608 18.192 0.64 18.264 ;
  LAYER M2 ;
        RECT 0.588 18.212 0.66 18.244 ;
  LAYER M2 ;
        RECT 0.4 18.212 0.624 18.244 ;
  LAYER M1 ;
        RECT 0.384 18.192 0.416 18.264 ;
  LAYER M2 ;
        RECT 0.364 18.212 0.436 18.244 ;
  LAYER M1 ;
        RECT 0.384 31.38 0.416 31.452 ;
  LAYER M2 ;
        RECT 0.364 31.4 0.436 31.432 ;
  LAYER M1 ;
        RECT 0.384 30.828 0.416 31.416 ;
  LAYER M1 ;
        RECT 0.384 18.228 0.416 30.828 ;
  LAYER M2 ;
        RECT 0.4 31.4 15.28 31.432 ;
  LAYER M1 ;
        RECT 9.536 30.456 9.568 30.528 ;
  LAYER M2 ;
        RECT 9.516 30.476 9.588 30.508 ;
  LAYER M2 ;
        RECT 9.552 30.476 12.528 30.508 ;
  LAYER M1 ;
        RECT 12.512 30.456 12.544 30.528 ;
  LAYER M2 ;
        RECT 12.492 30.476 12.564 30.508 ;
  LAYER M1 ;
        RECT 9.536 18.024 9.568 18.096 ;
  LAYER M2 ;
        RECT 9.516 18.044 9.588 18.076 ;
  LAYER M2 ;
        RECT 9.552 18.044 12.528 18.076 ;
  LAYER M1 ;
        RECT 12.512 18.024 12.544 18.096 ;
  LAYER M2 ;
        RECT 12.492 18.044 12.564 18.076 ;
  LAYER M1 ;
        RECT 6.56 18.024 6.592 18.096 ;
  LAYER M2 ;
        RECT 6.54 18.044 6.612 18.076 ;
  LAYER M2 ;
        RECT 6.576 18.044 9.552 18.076 ;
  LAYER M1 ;
        RECT 9.536 18.024 9.568 18.096 ;
  LAYER M2 ;
        RECT 9.516 18.044 9.588 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M2 ;
        RECT 3.6 18.044 6.576 18.076 ;
  LAYER M1 ;
        RECT 6.56 18.024 6.592 18.096 ;
  LAYER M2 ;
        RECT 6.54 18.044 6.612 18.076 ;
  LAYER M1 ;
        RECT 3.584 30.456 3.616 30.528 ;
  LAYER M2 ;
        RECT 3.564 30.476 3.636 30.508 ;
  LAYER M2 ;
        RECT 0.624 30.476 3.6 30.508 ;
  LAYER M1 ;
        RECT 0.608 30.456 0.64 30.528 ;
  LAYER M2 ;
        RECT 0.588 30.476 0.66 30.508 ;
  LAYER M1 ;
        RECT 6.56 30.456 6.592 30.528 ;
  LAYER M2 ;
        RECT 6.54 30.476 6.612 30.508 ;
  LAYER M2 ;
        RECT 3.6 30.476 6.576 30.508 ;
  LAYER M1 ;
        RECT 3.584 30.456 3.616 30.528 ;
  LAYER M2 ;
        RECT 3.564 30.476 3.636 30.508 ;
  LAYER M1 ;
        RECT 8.928 21.804 8.96 21.876 ;
  LAYER M2 ;
        RECT 8.908 21.824 8.98 21.856 ;
  LAYER M2 ;
        RECT 8.944 21.824 9.168 21.856 ;
  LAYER M1 ;
        RECT 9.152 21.804 9.184 21.876 ;
  LAYER M2 ;
        RECT 9.132 21.824 9.204 21.856 ;
  LAYER M1 ;
        RECT 11.904 18.696 11.936 18.768 ;
  LAYER M2 ;
        RECT 11.884 18.716 11.956 18.748 ;
  LAYER M1 ;
        RECT 11.904 18.564 11.936 18.732 ;
  LAYER M1 ;
        RECT 11.904 18.528 11.936 18.6 ;
  LAYER M2 ;
        RECT 11.884 18.548 11.956 18.58 ;
  LAYER M2 ;
        RECT 9.168 18.548 11.92 18.58 ;
  LAYER M1 ;
        RECT 9.152 18.528 9.184 18.6 ;
  LAYER M2 ;
        RECT 9.132 18.548 9.204 18.58 ;
  LAYER M1 ;
        RECT 9.152 15 9.184 15.072 ;
  LAYER M2 ;
        RECT 9.132 15.02 9.204 15.052 ;
  LAYER M1 ;
        RECT 9.152 15.036 9.184 15.288 ;
  LAYER M1 ;
        RECT 9.152 15.288 9.184 21.84 ;
  LAYER M1 ;
        RECT 5.952 24.912 5.984 24.984 ;
  LAYER M2 ;
        RECT 5.932 24.932 6.004 24.964 ;
  LAYER M2 ;
        RECT 5.968 24.932 6.192 24.964 ;
  LAYER M1 ;
        RECT 6.176 24.912 6.208 24.984 ;
  LAYER M2 ;
        RECT 6.156 24.932 6.228 24.964 ;
  LAYER M1 ;
        RECT 6.176 15 6.208 15.072 ;
  LAYER M2 ;
        RECT 6.156 15.02 6.228 15.052 ;
  LAYER M1 ;
        RECT 6.176 15.036 6.208 15.288 ;
  LAYER M1 ;
        RECT 6.176 15.288 6.208 24.948 ;
  LAYER M2 ;
        RECT 6.192 15.02 9.168 15.052 ;
  LAYER M1 ;
        RECT 11.904 21.804 11.936 21.876 ;
  LAYER M2 ;
        RECT 11.884 21.824 11.956 21.856 ;
  LAYER M2 ;
        RECT 11.92 21.824 12.144 21.856 ;
  LAYER M1 ;
        RECT 12.128 21.804 12.16 21.876 ;
  LAYER M2 ;
        RECT 12.108 21.824 12.18 21.856 ;
  LAYER M1 ;
        RECT 11.904 24.912 11.936 24.984 ;
  LAYER M2 ;
        RECT 11.884 24.932 11.956 24.964 ;
  LAYER M2 ;
        RECT 11.92 24.932 12.144 24.964 ;
  LAYER M1 ;
        RECT 12.128 24.912 12.16 24.984 ;
  LAYER M2 ;
        RECT 12.108 24.932 12.18 24.964 ;
  LAYER M1 ;
        RECT 12.128 14.832 12.16 14.904 ;
  LAYER M2 ;
        RECT 12.108 14.852 12.18 14.884 ;
  LAYER M1 ;
        RECT 12.128 14.868 12.16 15.288 ;
  LAYER M1 ;
        RECT 12.128 15.288 12.16 24.948 ;
  LAYER M1 ;
        RECT 5.952 21.804 5.984 21.876 ;
  LAYER M2 ;
        RECT 5.932 21.824 6.004 21.856 ;
  LAYER M1 ;
        RECT 5.952 21.672 5.984 21.84 ;
  LAYER M1 ;
        RECT 5.952 21.636 5.984 21.708 ;
  LAYER M2 ;
        RECT 5.932 21.656 6.004 21.688 ;
  LAYER M2 ;
        RECT 3.216 21.656 5.968 21.688 ;
  LAYER M1 ;
        RECT 3.2 21.636 3.232 21.708 ;
  LAYER M2 ;
        RECT 3.18 21.656 3.252 21.688 ;
  LAYER M1 ;
        RECT 5.952 18.696 5.984 18.768 ;
  LAYER M2 ;
        RECT 5.932 18.716 6.004 18.748 ;
  LAYER M1 ;
        RECT 5.952 18.564 5.984 18.732 ;
  LAYER M1 ;
        RECT 5.952 18.528 5.984 18.6 ;
  LAYER M2 ;
        RECT 5.932 18.548 6.004 18.58 ;
  LAYER M2 ;
        RECT 3.216 18.548 5.968 18.58 ;
  LAYER M1 ;
        RECT 3.2 18.528 3.232 18.6 ;
  LAYER M2 ;
        RECT 3.18 18.548 3.252 18.58 ;
  LAYER M1 ;
        RECT 3.2 14.832 3.232 14.904 ;
  LAYER M2 ;
        RECT 3.18 14.852 3.252 14.884 ;
  LAYER M1 ;
        RECT 3.2 14.868 3.232 15.288 ;
  LAYER M1 ;
        RECT 3.2 15.288 3.232 21.672 ;
  LAYER M2 ;
        RECT 3.216 14.852 12.144 14.884 ;
  LAYER M1 ;
        RECT 8.928 24.912 8.96 24.984 ;
  LAYER M2 ;
        RECT 8.908 24.932 8.98 24.964 ;
  LAYER M2 ;
        RECT 8.944 24.932 11.92 24.964 ;
  LAYER M1 ;
        RECT 11.904 24.912 11.936 24.984 ;
  LAYER M2 ;
        RECT 11.884 24.932 11.956 24.964 ;
  LAYER M1 ;
        RECT 8.928 18.696 8.96 18.768 ;
  LAYER M2 ;
        RECT 8.908 18.716 8.98 18.748 ;
  LAYER M2 ;
        RECT 5.968 18.716 8.944 18.748 ;
  LAYER M1 ;
        RECT 5.952 18.696 5.984 18.768 ;
  LAYER M2 ;
        RECT 5.932 18.716 6.004 18.748 ;
  LAYER M1 ;
        RECT 14.88 28.02 14.912 28.092 ;
  LAYER M2 ;
        RECT 14.86 28.04 14.932 28.072 ;
  LAYER M2 ;
        RECT 14.896 28.04 15.12 28.072 ;
  LAYER M1 ;
        RECT 15.104 28.02 15.136 28.092 ;
  LAYER M2 ;
        RECT 15.084 28.04 15.156 28.072 ;
  LAYER M1 ;
        RECT 14.88 24.912 14.912 24.984 ;
  LAYER M2 ;
        RECT 14.86 24.932 14.932 24.964 ;
  LAYER M2 ;
        RECT 14.896 24.932 15.12 24.964 ;
  LAYER M1 ;
        RECT 15.104 24.912 15.136 24.984 ;
  LAYER M2 ;
        RECT 15.084 24.932 15.156 24.964 ;
  LAYER M1 ;
        RECT 14.88 21.804 14.912 21.876 ;
  LAYER M2 ;
        RECT 14.86 21.824 14.932 21.856 ;
  LAYER M2 ;
        RECT 14.896 21.824 15.12 21.856 ;
  LAYER M1 ;
        RECT 15.104 21.804 15.136 21.876 ;
  LAYER M2 ;
        RECT 15.084 21.824 15.156 21.856 ;
  LAYER M1 ;
        RECT 14.88 18.696 14.912 18.768 ;
  LAYER M2 ;
        RECT 14.86 18.716 14.932 18.748 ;
  LAYER M2 ;
        RECT 14.896 18.716 15.12 18.748 ;
  LAYER M1 ;
        RECT 15.104 18.696 15.136 18.768 ;
  LAYER M2 ;
        RECT 15.084 18.716 15.156 18.748 ;
  LAYER M1 ;
        RECT 14.88 15.588 14.912 15.66 ;
  LAYER M2 ;
        RECT 14.86 15.608 14.932 15.64 ;
  LAYER M2 ;
        RECT 14.896 15.608 15.12 15.64 ;
  LAYER M1 ;
        RECT 15.104 15.588 15.136 15.66 ;
  LAYER M2 ;
        RECT 15.084 15.608 15.156 15.64 ;
  LAYER M1 ;
        RECT 15.104 14.664 15.136 14.736 ;
  LAYER M2 ;
        RECT 15.084 14.684 15.156 14.716 ;
  LAYER M1 ;
        RECT 15.104 14.7 15.136 15.288 ;
  LAYER M1 ;
        RECT 15.104 15.288 15.136 28.056 ;
  LAYER M1 ;
        RECT 2.976 28.02 3.008 28.092 ;
  LAYER M2 ;
        RECT 2.956 28.04 3.028 28.072 ;
  LAYER M1 ;
        RECT 2.976 27.888 3.008 28.056 ;
  LAYER M1 ;
        RECT 2.976 27.852 3.008 27.924 ;
  LAYER M2 ;
        RECT 2.956 27.872 3.028 27.904 ;
  LAYER M2 ;
        RECT 0.24 27.872 2.992 27.904 ;
  LAYER M1 ;
        RECT 0.224 27.852 0.256 27.924 ;
  LAYER M2 ;
        RECT 0.204 27.872 0.276 27.904 ;
  LAYER M1 ;
        RECT 2.976 24.912 3.008 24.984 ;
  LAYER M2 ;
        RECT 2.956 24.932 3.028 24.964 ;
  LAYER M1 ;
        RECT 2.976 24.78 3.008 24.948 ;
  LAYER M1 ;
        RECT 2.976 24.744 3.008 24.816 ;
  LAYER M2 ;
        RECT 2.956 24.764 3.028 24.796 ;
  LAYER M2 ;
        RECT 0.24 24.764 2.992 24.796 ;
  LAYER M1 ;
        RECT 0.224 24.744 0.256 24.816 ;
  LAYER M2 ;
        RECT 0.204 24.764 0.276 24.796 ;
  LAYER M1 ;
        RECT 2.976 21.804 3.008 21.876 ;
  LAYER M2 ;
        RECT 2.956 21.824 3.028 21.856 ;
  LAYER M1 ;
        RECT 2.976 21.672 3.008 21.84 ;
  LAYER M1 ;
        RECT 2.976 21.636 3.008 21.708 ;
  LAYER M2 ;
        RECT 2.956 21.656 3.028 21.688 ;
  LAYER M2 ;
        RECT 0.24 21.656 2.992 21.688 ;
  LAYER M1 ;
        RECT 0.224 21.636 0.256 21.708 ;
  LAYER M2 ;
        RECT 0.204 21.656 0.276 21.688 ;
  LAYER M1 ;
        RECT 2.976 18.696 3.008 18.768 ;
  LAYER M2 ;
        RECT 2.956 18.716 3.028 18.748 ;
  LAYER M1 ;
        RECT 2.976 18.564 3.008 18.732 ;
  LAYER M1 ;
        RECT 2.976 18.528 3.008 18.6 ;
  LAYER M2 ;
        RECT 2.956 18.548 3.028 18.58 ;
  LAYER M2 ;
        RECT 0.24 18.548 2.992 18.58 ;
  LAYER M1 ;
        RECT 0.224 18.528 0.256 18.6 ;
  LAYER M2 ;
        RECT 0.204 18.548 0.276 18.58 ;
  LAYER M1 ;
        RECT 2.976 15.588 3.008 15.66 ;
  LAYER M2 ;
        RECT 2.956 15.608 3.028 15.64 ;
  LAYER M1 ;
        RECT 2.976 15.456 3.008 15.624 ;
  LAYER M1 ;
        RECT 2.976 15.42 3.008 15.492 ;
  LAYER M2 ;
        RECT 2.956 15.44 3.028 15.472 ;
  LAYER M2 ;
        RECT 0.24 15.44 2.992 15.472 ;
  LAYER M1 ;
        RECT 0.224 15.42 0.256 15.492 ;
  LAYER M2 ;
        RECT 0.204 15.44 0.276 15.472 ;
  LAYER M1 ;
        RECT 0.224 14.664 0.256 14.736 ;
  LAYER M2 ;
        RECT 0.204 14.684 0.276 14.716 ;
  LAYER M1 ;
        RECT 0.224 14.7 0.256 15.288 ;
  LAYER M1 ;
        RECT 0.224 15.288 0.256 27.888 ;
  LAYER M2 ;
        RECT 0.24 14.684 15.12 14.716 ;
  LAYER M1 ;
        RECT 11.904 28.02 11.936 28.092 ;
  LAYER M2 ;
        RECT 11.884 28.04 11.956 28.072 ;
  LAYER M2 ;
        RECT 11.92 28.04 14.896 28.072 ;
  LAYER M1 ;
        RECT 14.88 28.02 14.912 28.092 ;
  LAYER M2 ;
        RECT 14.86 28.04 14.932 28.072 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 15.66 ;
  LAYER M2 ;
        RECT 11.884 15.608 11.956 15.64 ;
  LAYER M2 ;
        RECT 11.92 15.608 14.896 15.64 ;
  LAYER M1 ;
        RECT 14.88 15.588 14.912 15.66 ;
  LAYER M2 ;
        RECT 14.86 15.608 14.932 15.64 ;
  LAYER M1 ;
        RECT 8.928 15.588 8.96 15.66 ;
  LAYER M2 ;
        RECT 8.908 15.608 8.98 15.64 ;
  LAYER M2 ;
        RECT 8.944 15.608 11.92 15.64 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 15.66 ;
  LAYER M2 ;
        RECT 11.884 15.608 11.956 15.64 ;
  LAYER M1 ;
        RECT 5.952 15.588 5.984 15.66 ;
  LAYER M2 ;
        RECT 5.932 15.608 6.004 15.64 ;
  LAYER M2 ;
        RECT 5.968 15.608 8.944 15.64 ;
  LAYER M1 ;
        RECT 8.928 15.588 8.96 15.66 ;
  LAYER M2 ;
        RECT 8.908 15.608 8.98 15.64 ;
  LAYER M1 ;
        RECT 5.952 28.02 5.984 28.092 ;
  LAYER M2 ;
        RECT 5.932 28.04 6.004 28.072 ;
  LAYER M2 ;
        RECT 2.992 28.04 5.968 28.072 ;
  LAYER M1 ;
        RECT 2.976 28.02 3.008 28.092 ;
  LAYER M2 ;
        RECT 2.956 28.04 3.028 28.072 ;
  LAYER M1 ;
        RECT 8.928 28.02 8.96 28.092 ;
  LAYER M2 ;
        RECT 8.908 28.04 8.98 28.072 ;
  LAYER M2 ;
        RECT 5.968 28.04 8.944 28.072 ;
  LAYER M1 ;
        RECT 5.952 28.02 5.984 28.092 ;
  LAYER M2 ;
        RECT 5.932 28.04 6.004 28.072 ;
  LAYER M1 ;
        RECT 14.88 28.02 14.912 30.528 ;
  LAYER M3 ;
        RECT 14.88 28.04 14.912 28.072 ;
  LAYER M1 ;
        RECT 14.816 28.02 14.848 30.528 ;
  LAYER M3 ;
        RECT 14.816 30.476 14.848 30.508 ;
  LAYER M1 ;
        RECT 14.752 28.02 14.784 30.528 ;
  LAYER M3 ;
        RECT 14.752 28.04 14.784 28.072 ;
  LAYER M1 ;
        RECT 14.688 28.02 14.72 30.528 ;
  LAYER M3 ;
        RECT 14.688 30.476 14.72 30.508 ;
  LAYER M1 ;
        RECT 14.624 28.02 14.656 30.528 ;
  LAYER M3 ;
        RECT 14.624 28.04 14.656 28.072 ;
  LAYER M1 ;
        RECT 14.56 28.02 14.592 30.528 ;
  LAYER M3 ;
        RECT 14.56 30.476 14.592 30.508 ;
  LAYER M1 ;
        RECT 14.496 28.02 14.528 30.528 ;
  LAYER M3 ;
        RECT 14.496 28.04 14.528 28.072 ;
  LAYER M1 ;
        RECT 14.432 28.02 14.464 30.528 ;
  LAYER M3 ;
        RECT 14.432 30.476 14.464 30.508 ;
  LAYER M1 ;
        RECT 14.368 28.02 14.4 30.528 ;
  LAYER M3 ;
        RECT 14.368 28.04 14.4 28.072 ;
  LAYER M1 ;
        RECT 14.304 28.02 14.336 30.528 ;
  LAYER M3 ;
        RECT 14.304 30.476 14.336 30.508 ;
  LAYER M1 ;
        RECT 14.24 28.02 14.272 30.528 ;
  LAYER M3 ;
        RECT 14.24 28.04 14.272 28.072 ;
  LAYER M1 ;
        RECT 14.176 28.02 14.208 30.528 ;
  LAYER M3 ;
        RECT 14.176 30.476 14.208 30.508 ;
  LAYER M1 ;
        RECT 14.112 28.02 14.144 30.528 ;
  LAYER M3 ;
        RECT 14.112 28.04 14.144 28.072 ;
  LAYER M1 ;
        RECT 14.048 28.02 14.08 30.528 ;
  LAYER M3 ;
        RECT 14.048 30.476 14.08 30.508 ;
  LAYER M1 ;
        RECT 13.984 28.02 14.016 30.528 ;
  LAYER M3 ;
        RECT 13.984 28.04 14.016 28.072 ;
  LAYER M1 ;
        RECT 13.92 28.02 13.952 30.528 ;
  LAYER M3 ;
        RECT 13.92 30.476 13.952 30.508 ;
  LAYER M1 ;
        RECT 13.856 28.02 13.888 30.528 ;
  LAYER M3 ;
        RECT 13.856 28.04 13.888 28.072 ;
  LAYER M1 ;
        RECT 13.792 28.02 13.824 30.528 ;
  LAYER M3 ;
        RECT 13.792 30.476 13.824 30.508 ;
  LAYER M1 ;
        RECT 13.728 28.02 13.76 30.528 ;
  LAYER M3 ;
        RECT 13.728 28.04 13.76 28.072 ;
  LAYER M1 ;
        RECT 13.664 28.02 13.696 30.528 ;
  LAYER M3 ;
        RECT 13.664 30.476 13.696 30.508 ;
  LAYER M1 ;
        RECT 13.6 28.02 13.632 30.528 ;
  LAYER M3 ;
        RECT 13.6 28.04 13.632 28.072 ;
  LAYER M1 ;
        RECT 13.536 28.02 13.568 30.528 ;
  LAYER M3 ;
        RECT 13.536 30.476 13.568 30.508 ;
  LAYER M1 ;
        RECT 13.472 28.02 13.504 30.528 ;
  LAYER M3 ;
        RECT 13.472 28.04 13.504 28.072 ;
  LAYER M1 ;
        RECT 13.408 28.02 13.44 30.528 ;
  LAYER M3 ;
        RECT 13.408 30.476 13.44 30.508 ;
  LAYER M1 ;
        RECT 13.344 28.02 13.376 30.528 ;
  LAYER M3 ;
        RECT 13.344 28.04 13.376 28.072 ;
  LAYER M1 ;
        RECT 13.28 28.02 13.312 30.528 ;
  LAYER M3 ;
        RECT 13.28 30.476 13.312 30.508 ;
  LAYER M1 ;
        RECT 13.216 28.02 13.248 30.528 ;
  LAYER M3 ;
        RECT 13.216 28.04 13.248 28.072 ;
  LAYER M1 ;
        RECT 13.152 28.02 13.184 30.528 ;
  LAYER M3 ;
        RECT 13.152 30.476 13.184 30.508 ;
  LAYER M1 ;
        RECT 13.088 28.02 13.12 30.528 ;
  LAYER M3 ;
        RECT 13.088 28.04 13.12 28.072 ;
  LAYER M1 ;
        RECT 13.024 28.02 13.056 30.528 ;
  LAYER M3 ;
        RECT 13.024 30.476 13.056 30.508 ;
  LAYER M1 ;
        RECT 12.96 28.02 12.992 30.528 ;
  LAYER M3 ;
        RECT 12.96 28.04 12.992 28.072 ;
  LAYER M1 ;
        RECT 12.896 28.02 12.928 30.528 ;
  LAYER M3 ;
        RECT 12.896 30.476 12.928 30.508 ;
  LAYER M1 ;
        RECT 12.832 28.02 12.864 30.528 ;
  LAYER M3 ;
        RECT 12.832 28.04 12.864 28.072 ;
  LAYER M1 ;
        RECT 12.768 28.02 12.8 30.528 ;
  LAYER M3 ;
        RECT 12.768 30.476 12.8 30.508 ;
  LAYER M1 ;
        RECT 12.704 28.02 12.736 30.528 ;
  LAYER M3 ;
        RECT 12.704 28.04 12.736 28.072 ;
  LAYER M1 ;
        RECT 12.64 28.02 12.672 30.528 ;
  LAYER M3 ;
        RECT 12.64 30.476 12.672 30.508 ;
  LAYER M1 ;
        RECT 12.576 28.02 12.608 30.528 ;
  LAYER M3 ;
        RECT 12.576 28.04 12.608 28.072 ;
  LAYER M1 ;
        RECT 12.512 28.02 12.544 30.528 ;
  LAYER M3 ;
        RECT 14.88 30.412 14.912 30.444 ;
  LAYER M2 ;
        RECT 12.512 30.348 12.544 30.38 ;
  LAYER M2 ;
        RECT 14.88 30.284 14.912 30.316 ;
  LAYER M2 ;
        RECT 12.512 30.22 12.544 30.252 ;
  LAYER M2 ;
        RECT 14.88 30.156 14.912 30.188 ;
  LAYER M2 ;
        RECT 12.512 30.092 12.544 30.124 ;
  LAYER M2 ;
        RECT 14.88 30.028 14.912 30.06 ;
  LAYER M2 ;
        RECT 12.512 29.964 12.544 29.996 ;
  LAYER M2 ;
        RECT 14.88 29.9 14.912 29.932 ;
  LAYER M2 ;
        RECT 12.512 29.836 12.544 29.868 ;
  LAYER M2 ;
        RECT 14.88 29.772 14.912 29.804 ;
  LAYER M2 ;
        RECT 12.512 29.708 12.544 29.74 ;
  LAYER M2 ;
        RECT 14.88 29.644 14.912 29.676 ;
  LAYER M2 ;
        RECT 12.512 29.58 12.544 29.612 ;
  LAYER M2 ;
        RECT 14.88 29.516 14.912 29.548 ;
  LAYER M2 ;
        RECT 12.512 29.452 12.544 29.484 ;
  LAYER M2 ;
        RECT 14.88 29.388 14.912 29.42 ;
  LAYER M2 ;
        RECT 12.512 29.324 12.544 29.356 ;
  LAYER M2 ;
        RECT 14.88 29.26 14.912 29.292 ;
  LAYER M2 ;
        RECT 12.512 29.196 12.544 29.228 ;
  LAYER M2 ;
        RECT 14.88 29.132 14.912 29.164 ;
  LAYER M2 ;
        RECT 12.512 29.068 12.544 29.1 ;
  LAYER M2 ;
        RECT 14.88 29.004 14.912 29.036 ;
  LAYER M2 ;
        RECT 12.512 28.94 12.544 28.972 ;
  LAYER M2 ;
        RECT 14.88 28.876 14.912 28.908 ;
  LAYER M2 ;
        RECT 12.512 28.812 12.544 28.844 ;
  LAYER M2 ;
        RECT 14.88 28.748 14.912 28.78 ;
  LAYER M2 ;
        RECT 12.512 28.684 12.544 28.716 ;
  LAYER M2 ;
        RECT 14.88 28.62 14.912 28.652 ;
  LAYER M2 ;
        RECT 12.512 28.556 12.544 28.588 ;
  LAYER M2 ;
        RECT 14.88 28.492 14.912 28.524 ;
  LAYER M2 ;
        RECT 12.512 28.428 12.544 28.46 ;
  LAYER M2 ;
        RECT 14.88 28.364 14.912 28.396 ;
  LAYER M2 ;
        RECT 12.512 28.3 12.544 28.332 ;
  LAYER M2 ;
        RECT 14.88 28.236 14.912 28.268 ;
  LAYER M2 ;
        RECT 12.512 28.172 12.544 28.204 ;
  LAYER M2 ;
        RECT 12.464 27.972 14.96 30.576 ;
  LAYER M1 ;
        RECT 14.88 24.912 14.912 27.42 ;
  LAYER M3 ;
        RECT 14.88 24.932 14.912 24.964 ;
  LAYER M1 ;
        RECT 14.816 24.912 14.848 27.42 ;
  LAYER M3 ;
        RECT 14.816 27.368 14.848 27.4 ;
  LAYER M1 ;
        RECT 14.752 24.912 14.784 27.42 ;
  LAYER M3 ;
        RECT 14.752 24.932 14.784 24.964 ;
  LAYER M1 ;
        RECT 14.688 24.912 14.72 27.42 ;
  LAYER M3 ;
        RECT 14.688 27.368 14.72 27.4 ;
  LAYER M1 ;
        RECT 14.624 24.912 14.656 27.42 ;
  LAYER M3 ;
        RECT 14.624 24.932 14.656 24.964 ;
  LAYER M1 ;
        RECT 14.56 24.912 14.592 27.42 ;
  LAYER M3 ;
        RECT 14.56 27.368 14.592 27.4 ;
  LAYER M1 ;
        RECT 14.496 24.912 14.528 27.42 ;
  LAYER M3 ;
        RECT 14.496 24.932 14.528 24.964 ;
  LAYER M1 ;
        RECT 14.432 24.912 14.464 27.42 ;
  LAYER M3 ;
        RECT 14.432 27.368 14.464 27.4 ;
  LAYER M1 ;
        RECT 14.368 24.912 14.4 27.42 ;
  LAYER M3 ;
        RECT 14.368 24.932 14.4 24.964 ;
  LAYER M1 ;
        RECT 14.304 24.912 14.336 27.42 ;
  LAYER M3 ;
        RECT 14.304 27.368 14.336 27.4 ;
  LAYER M1 ;
        RECT 14.24 24.912 14.272 27.42 ;
  LAYER M3 ;
        RECT 14.24 24.932 14.272 24.964 ;
  LAYER M1 ;
        RECT 14.176 24.912 14.208 27.42 ;
  LAYER M3 ;
        RECT 14.176 27.368 14.208 27.4 ;
  LAYER M1 ;
        RECT 14.112 24.912 14.144 27.42 ;
  LAYER M3 ;
        RECT 14.112 24.932 14.144 24.964 ;
  LAYER M1 ;
        RECT 14.048 24.912 14.08 27.42 ;
  LAYER M3 ;
        RECT 14.048 27.368 14.08 27.4 ;
  LAYER M1 ;
        RECT 13.984 24.912 14.016 27.42 ;
  LAYER M3 ;
        RECT 13.984 24.932 14.016 24.964 ;
  LAYER M1 ;
        RECT 13.92 24.912 13.952 27.42 ;
  LAYER M3 ;
        RECT 13.92 27.368 13.952 27.4 ;
  LAYER M1 ;
        RECT 13.856 24.912 13.888 27.42 ;
  LAYER M3 ;
        RECT 13.856 24.932 13.888 24.964 ;
  LAYER M1 ;
        RECT 13.792 24.912 13.824 27.42 ;
  LAYER M3 ;
        RECT 13.792 27.368 13.824 27.4 ;
  LAYER M1 ;
        RECT 13.728 24.912 13.76 27.42 ;
  LAYER M3 ;
        RECT 13.728 24.932 13.76 24.964 ;
  LAYER M1 ;
        RECT 13.664 24.912 13.696 27.42 ;
  LAYER M3 ;
        RECT 13.664 27.368 13.696 27.4 ;
  LAYER M1 ;
        RECT 13.6 24.912 13.632 27.42 ;
  LAYER M3 ;
        RECT 13.6 24.932 13.632 24.964 ;
  LAYER M1 ;
        RECT 13.536 24.912 13.568 27.42 ;
  LAYER M3 ;
        RECT 13.536 27.368 13.568 27.4 ;
  LAYER M1 ;
        RECT 13.472 24.912 13.504 27.42 ;
  LAYER M3 ;
        RECT 13.472 24.932 13.504 24.964 ;
  LAYER M1 ;
        RECT 13.408 24.912 13.44 27.42 ;
  LAYER M3 ;
        RECT 13.408 27.368 13.44 27.4 ;
  LAYER M1 ;
        RECT 13.344 24.912 13.376 27.42 ;
  LAYER M3 ;
        RECT 13.344 24.932 13.376 24.964 ;
  LAYER M1 ;
        RECT 13.28 24.912 13.312 27.42 ;
  LAYER M3 ;
        RECT 13.28 27.368 13.312 27.4 ;
  LAYER M1 ;
        RECT 13.216 24.912 13.248 27.42 ;
  LAYER M3 ;
        RECT 13.216 24.932 13.248 24.964 ;
  LAYER M1 ;
        RECT 13.152 24.912 13.184 27.42 ;
  LAYER M3 ;
        RECT 13.152 27.368 13.184 27.4 ;
  LAYER M1 ;
        RECT 13.088 24.912 13.12 27.42 ;
  LAYER M3 ;
        RECT 13.088 24.932 13.12 24.964 ;
  LAYER M1 ;
        RECT 13.024 24.912 13.056 27.42 ;
  LAYER M3 ;
        RECT 13.024 27.368 13.056 27.4 ;
  LAYER M1 ;
        RECT 12.96 24.912 12.992 27.42 ;
  LAYER M3 ;
        RECT 12.96 24.932 12.992 24.964 ;
  LAYER M1 ;
        RECT 12.896 24.912 12.928 27.42 ;
  LAYER M3 ;
        RECT 12.896 27.368 12.928 27.4 ;
  LAYER M1 ;
        RECT 12.832 24.912 12.864 27.42 ;
  LAYER M3 ;
        RECT 12.832 24.932 12.864 24.964 ;
  LAYER M1 ;
        RECT 12.768 24.912 12.8 27.42 ;
  LAYER M3 ;
        RECT 12.768 27.368 12.8 27.4 ;
  LAYER M1 ;
        RECT 12.704 24.912 12.736 27.42 ;
  LAYER M3 ;
        RECT 12.704 24.932 12.736 24.964 ;
  LAYER M1 ;
        RECT 12.64 24.912 12.672 27.42 ;
  LAYER M3 ;
        RECT 12.64 27.368 12.672 27.4 ;
  LAYER M1 ;
        RECT 12.576 24.912 12.608 27.42 ;
  LAYER M3 ;
        RECT 12.576 24.932 12.608 24.964 ;
  LAYER M1 ;
        RECT 12.512 24.912 12.544 27.42 ;
  LAYER M3 ;
        RECT 14.88 27.304 14.912 27.336 ;
  LAYER M2 ;
        RECT 12.512 27.24 12.544 27.272 ;
  LAYER M2 ;
        RECT 14.88 27.176 14.912 27.208 ;
  LAYER M2 ;
        RECT 12.512 27.112 12.544 27.144 ;
  LAYER M2 ;
        RECT 14.88 27.048 14.912 27.08 ;
  LAYER M2 ;
        RECT 12.512 26.984 12.544 27.016 ;
  LAYER M2 ;
        RECT 14.88 26.92 14.912 26.952 ;
  LAYER M2 ;
        RECT 12.512 26.856 12.544 26.888 ;
  LAYER M2 ;
        RECT 14.88 26.792 14.912 26.824 ;
  LAYER M2 ;
        RECT 12.512 26.728 12.544 26.76 ;
  LAYER M2 ;
        RECT 14.88 26.664 14.912 26.696 ;
  LAYER M2 ;
        RECT 12.512 26.6 12.544 26.632 ;
  LAYER M2 ;
        RECT 14.88 26.536 14.912 26.568 ;
  LAYER M2 ;
        RECT 12.512 26.472 12.544 26.504 ;
  LAYER M2 ;
        RECT 14.88 26.408 14.912 26.44 ;
  LAYER M2 ;
        RECT 12.512 26.344 12.544 26.376 ;
  LAYER M2 ;
        RECT 14.88 26.28 14.912 26.312 ;
  LAYER M2 ;
        RECT 12.512 26.216 12.544 26.248 ;
  LAYER M2 ;
        RECT 14.88 26.152 14.912 26.184 ;
  LAYER M2 ;
        RECT 12.512 26.088 12.544 26.12 ;
  LAYER M2 ;
        RECT 14.88 26.024 14.912 26.056 ;
  LAYER M2 ;
        RECT 12.512 25.96 12.544 25.992 ;
  LAYER M2 ;
        RECT 14.88 25.896 14.912 25.928 ;
  LAYER M2 ;
        RECT 12.512 25.832 12.544 25.864 ;
  LAYER M2 ;
        RECT 14.88 25.768 14.912 25.8 ;
  LAYER M2 ;
        RECT 12.512 25.704 12.544 25.736 ;
  LAYER M2 ;
        RECT 14.88 25.64 14.912 25.672 ;
  LAYER M2 ;
        RECT 12.512 25.576 12.544 25.608 ;
  LAYER M2 ;
        RECT 14.88 25.512 14.912 25.544 ;
  LAYER M2 ;
        RECT 12.512 25.448 12.544 25.48 ;
  LAYER M2 ;
        RECT 14.88 25.384 14.912 25.416 ;
  LAYER M2 ;
        RECT 12.512 25.32 12.544 25.352 ;
  LAYER M2 ;
        RECT 14.88 25.256 14.912 25.288 ;
  LAYER M2 ;
        RECT 12.512 25.192 12.544 25.224 ;
  LAYER M2 ;
        RECT 14.88 25.128 14.912 25.16 ;
  LAYER M2 ;
        RECT 12.512 25.064 12.544 25.096 ;
  LAYER M2 ;
        RECT 12.464 24.864 14.96 27.468 ;
  LAYER M1 ;
        RECT 14.88 21.804 14.912 24.312 ;
  LAYER M3 ;
        RECT 14.88 21.824 14.912 21.856 ;
  LAYER M1 ;
        RECT 14.816 21.804 14.848 24.312 ;
  LAYER M3 ;
        RECT 14.816 24.26 14.848 24.292 ;
  LAYER M1 ;
        RECT 14.752 21.804 14.784 24.312 ;
  LAYER M3 ;
        RECT 14.752 21.824 14.784 21.856 ;
  LAYER M1 ;
        RECT 14.688 21.804 14.72 24.312 ;
  LAYER M3 ;
        RECT 14.688 24.26 14.72 24.292 ;
  LAYER M1 ;
        RECT 14.624 21.804 14.656 24.312 ;
  LAYER M3 ;
        RECT 14.624 21.824 14.656 21.856 ;
  LAYER M1 ;
        RECT 14.56 21.804 14.592 24.312 ;
  LAYER M3 ;
        RECT 14.56 24.26 14.592 24.292 ;
  LAYER M1 ;
        RECT 14.496 21.804 14.528 24.312 ;
  LAYER M3 ;
        RECT 14.496 21.824 14.528 21.856 ;
  LAYER M1 ;
        RECT 14.432 21.804 14.464 24.312 ;
  LAYER M3 ;
        RECT 14.432 24.26 14.464 24.292 ;
  LAYER M1 ;
        RECT 14.368 21.804 14.4 24.312 ;
  LAYER M3 ;
        RECT 14.368 21.824 14.4 21.856 ;
  LAYER M1 ;
        RECT 14.304 21.804 14.336 24.312 ;
  LAYER M3 ;
        RECT 14.304 24.26 14.336 24.292 ;
  LAYER M1 ;
        RECT 14.24 21.804 14.272 24.312 ;
  LAYER M3 ;
        RECT 14.24 21.824 14.272 21.856 ;
  LAYER M1 ;
        RECT 14.176 21.804 14.208 24.312 ;
  LAYER M3 ;
        RECT 14.176 24.26 14.208 24.292 ;
  LAYER M1 ;
        RECT 14.112 21.804 14.144 24.312 ;
  LAYER M3 ;
        RECT 14.112 21.824 14.144 21.856 ;
  LAYER M1 ;
        RECT 14.048 21.804 14.08 24.312 ;
  LAYER M3 ;
        RECT 14.048 24.26 14.08 24.292 ;
  LAYER M1 ;
        RECT 13.984 21.804 14.016 24.312 ;
  LAYER M3 ;
        RECT 13.984 21.824 14.016 21.856 ;
  LAYER M1 ;
        RECT 13.92 21.804 13.952 24.312 ;
  LAYER M3 ;
        RECT 13.92 24.26 13.952 24.292 ;
  LAYER M1 ;
        RECT 13.856 21.804 13.888 24.312 ;
  LAYER M3 ;
        RECT 13.856 21.824 13.888 21.856 ;
  LAYER M1 ;
        RECT 13.792 21.804 13.824 24.312 ;
  LAYER M3 ;
        RECT 13.792 24.26 13.824 24.292 ;
  LAYER M1 ;
        RECT 13.728 21.804 13.76 24.312 ;
  LAYER M3 ;
        RECT 13.728 21.824 13.76 21.856 ;
  LAYER M1 ;
        RECT 13.664 21.804 13.696 24.312 ;
  LAYER M3 ;
        RECT 13.664 24.26 13.696 24.292 ;
  LAYER M1 ;
        RECT 13.6 21.804 13.632 24.312 ;
  LAYER M3 ;
        RECT 13.6 21.824 13.632 21.856 ;
  LAYER M1 ;
        RECT 13.536 21.804 13.568 24.312 ;
  LAYER M3 ;
        RECT 13.536 24.26 13.568 24.292 ;
  LAYER M1 ;
        RECT 13.472 21.804 13.504 24.312 ;
  LAYER M3 ;
        RECT 13.472 21.824 13.504 21.856 ;
  LAYER M1 ;
        RECT 13.408 21.804 13.44 24.312 ;
  LAYER M3 ;
        RECT 13.408 24.26 13.44 24.292 ;
  LAYER M1 ;
        RECT 13.344 21.804 13.376 24.312 ;
  LAYER M3 ;
        RECT 13.344 21.824 13.376 21.856 ;
  LAYER M1 ;
        RECT 13.28 21.804 13.312 24.312 ;
  LAYER M3 ;
        RECT 13.28 24.26 13.312 24.292 ;
  LAYER M1 ;
        RECT 13.216 21.804 13.248 24.312 ;
  LAYER M3 ;
        RECT 13.216 21.824 13.248 21.856 ;
  LAYER M1 ;
        RECT 13.152 21.804 13.184 24.312 ;
  LAYER M3 ;
        RECT 13.152 24.26 13.184 24.292 ;
  LAYER M1 ;
        RECT 13.088 21.804 13.12 24.312 ;
  LAYER M3 ;
        RECT 13.088 21.824 13.12 21.856 ;
  LAYER M1 ;
        RECT 13.024 21.804 13.056 24.312 ;
  LAYER M3 ;
        RECT 13.024 24.26 13.056 24.292 ;
  LAYER M1 ;
        RECT 12.96 21.804 12.992 24.312 ;
  LAYER M3 ;
        RECT 12.96 21.824 12.992 21.856 ;
  LAYER M1 ;
        RECT 12.896 21.804 12.928 24.312 ;
  LAYER M3 ;
        RECT 12.896 24.26 12.928 24.292 ;
  LAYER M1 ;
        RECT 12.832 21.804 12.864 24.312 ;
  LAYER M3 ;
        RECT 12.832 21.824 12.864 21.856 ;
  LAYER M1 ;
        RECT 12.768 21.804 12.8 24.312 ;
  LAYER M3 ;
        RECT 12.768 24.26 12.8 24.292 ;
  LAYER M1 ;
        RECT 12.704 21.804 12.736 24.312 ;
  LAYER M3 ;
        RECT 12.704 21.824 12.736 21.856 ;
  LAYER M1 ;
        RECT 12.64 21.804 12.672 24.312 ;
  LAYER M3 ;
        RECT 12.64 24.26 12.672 24.292 ;
  LAYER M1 ;
        RECT 12.576 21.804 12.608 24.312 ;
  LAYER M3 ;
        RECT 12.576 21.824 12.608 21.856 ;
  LAYER M1 ;
        RECT 12.512 21.804 12.544 24.312 ;
  LAYER M3 ;
        RECT 14.88 24.196 14.912 24.228 ;
  LAYER M2 ;
        RECT 12.512 24.132 12.544 24.164 ;
  LAYER M2 ;
        RECT 14.88 24.068 14.912 24.1 ;
  LAYER M2 ;
        RECT 12.512 24.004 12.544 24.036 ;
  LAYER M2 ;
        RECT 14.88 23.94 14.912 23.972 ;
  LAYER M2 ;
        RECT 12.512 23.876 12.544 23.908 ;
  LAYER M2 ;
        RECT 14.88 23.812 14.912 23.844 ;
  LAYER M2 ;
        RECT 12.512 23.748 12.544 23.78 ;
  LAYER M2 ;
        RECT 14.88 23.684 14.912 23.716 ;
  LAYER M2 ;
        RECT 12.512 23.62 12.544 23.652 ;
  LAYER M2 ;
        RECT 14.88 23.556 14.912 23.588 ;
  LAYER M2 ;
        RECT 12.512 23.492 12.544 23.524 ;
  LAYER M2 ;
        RECT 14.88 23.428 14.912 23.46 ;
  LAYER M2 ;
        RECT 12.512 23.364 12.544 23.396 ;
  LAYER M2 ;
        RECT 14.88 23.3 14.912 23.332 ;
  LAYER M2 ;
        RECT 12.512 23.236 12.544 23.268 ;
  LAYER M2 ;
        RECT 14.88 23.172 14.912 23.204 ;
  LAYER M2 ;
        RECT 12.512 23.108 12.544 23.14 ;
  LAYER M2 ;
        RECT 14.88 23.044 14.912 23.076 ;
  LAYER M2 ;
        RECT 12.512 22.98 12.544 23.012 ;
  LAYER M2 ;
        RECT 14.88 22.916 14.912 22.948 ;
  LAYER M2 ;
        RECT 12.512 22.852 12.544 22.884 ;
  LAYER M2 ;
        RECT 14.88 22.788 14.912 22.82 ;
  LAYER M2 ;
        RECT 12.512 22.724 12.544 22.756 ;
  LAYER M2 ;
        RECT 14.88 22.66 14.912 22.692 ;
  LAYER M2 ;
        RECT 12.512 22.596 12.544 22.628 ;
  LAYER M2 ;
        RECT 14.88 22.532 14.912 22.564 ;
  LAYER M2 ;
        RECT 12.512 22.468 12.544 22.5 ;
  LAYER M2 ;
        RECT 14.88 22.404 14.912 22.436 ;
  LAYER M2 ;
        RECT 12.512 22.34 12.544 22.372 ;
  LAYER M2 ;
        RECT 14.88 22.276 14.912 22.308 ;
  LAYER M2 ;
        RECT 12.512 22.212 12.544 22.244 ;
  LAYER M2 ;
        RECT 14.88 22.148 14.912 22.18 ;
  LAYER M2 ;
        RECT 12.512 22.084 12.544 22.116 ;
  LAYER M2 ;
        RECT 14.88 22.02 14.912 22.052 ;
  LAYER M2 ;
        RECT 12.512 21.956 12.544 21.988 ;
  LAYER M2 ;
        RECT 12.464 21.756 14.96 24.36 ;
  LAYER M1 ;
        RECT 14.88 18.696 14.912 21.204 ;
  LAYER M3 ;
        RECT 14.88 18.716 14.912 18.748 ;
  LAYER M1 ;
        RECT 14.816 18.696 14.848 21.204 ;
  LAYER M3 ;
        RECT 14.816 21.152 14.848 21.184 ;
  LAYER M1 ;
        RECT 14.752 18.696 14.784 21.204 ;
  LAYER M3 ;
        RECT 14.752 18.716 14.784 18.748 ;
  LAYER M1 ;
        RECT 14.688 18.696 14.72 21.204 ;
  LAYER M3 ;
        RECT 14.688 21.152 14.72 21.184 ;
  LAYER M1 ;
        RECT 14.624 18.696 14.656 21.204 ;
  LAYER M3 ;
        RECT 14.624 18.716 14.656 18.748 ;
  LAYER M1 ;
        RECT 14.56 18.696 14.592 21.204 ;
  LAYER M3 ;
        RECT 14.56 21.152 14.592 21.184 ;
  LAYER M1 ;
        RECT 14.496 18.696 14.528 21.204 ;
  LAYER M3 ;
        RECT 14.496 18.716 14.528 18.748 ;
  LAYER M1 ;
        RECT 14.432 18.696 14.464 21.204 ;
  LAYER M3 ;
        RECT 14.432 21.152 14.464 21.184 ;
  LAYER M1 ;
        RECT 14.368 18.696 14.4 21.204 ;
  LAYER M3 ;
        RECT 14.368 18.716 14.4 18.748 ;
  LAYER M1 ;
        RECT 14.304 18.696 14.336 21.204 ;
  LAYER M3 ;
        RECT 14.304 21.152 14.336 21.184 ;
  LAYER M1 ;
        RECT 14.24 18.696 14.272 21.204 ;
  LAYER M3 ;
        RECT 14.24 18.716 14.272 18.748 ;
  LAYER M1 ;
        RECT 14.176 18.696 14.208 21.204 ;
  LAYER M3 ;
        RECT 14.176 21.152 14.208 21.184 ;
  LAYER M1 ;
        RECT 14.112 18.696 14.144 21.204 ;
  LAYER M3 ;
        RECT 14.112 18.716 14.144 18.748 ;
  LAYER M1 ;
        RECT 14.048 18.696 14.08 21.204 ;
  LAYER M3 ;
        RECT 14.048 21.152 14.08 21.184 ;
  LAYER M1 ;
        RECT 13.984 18.696 14.016 21.204 ;
  LAYER M3 ;
        RECT 13.984 18.716 14.016 18.748 ;
  LAYER M1 ;
        RECT 13.92 18.696 13.952 21.204 ;
  LAYER M3 ;
        RECT 13.92 21.152 13.952 21.184 ;
  LAYER M1 ;
        RECT 13.856 18.696 13.888 21.204 ;
  LAYER M3 ;
        RECT 13.856 18.716 13.888 18.748 ;
  LAYER M1 ;
        RECT 13.792 18.696 13.824 21.204 ;
  LAYER M3 ;
        RECT 13.792 21.152 13.824 21.184 ;
  LAYER M1 ;
        RECT 13.728 18.696 13.76 21.204 ;
  LAYER M3 ;
        RECT 13.728 18.716 13.76 18.748 ;
  LAYER M1 ;
        RECT 13.664 18.696 13.696 21.204 ;
  LAYER M3 ;
        RECT 13.664 21.152 13.696 21.184 ;
  LAYER M1 ;
        RECT 13.6 18.696 13.632 21.204 ;
  LAYER M3 ;
        RECT 13.6 18.716 13.632 18.748 ;
  LAYER M1 ;
        RECT 13.536 18.696 13.568 21.204 ;
  LAYER M3 ;
        RECT 13.536 21.152 13.568 21.184 ;
  LAYER M1 ;
        RECT 13.472 18.696 13.504 21.204 ;
  LAYER M3 ;
        RECT 13.472 18.716 13.504 18.748 ;
  LAYER M1 ;
        RECT 13.408 18.696 13.44 21.204 ;
  LAYER M3 ;
        RECT 13.408 21.152 13.44 21.184 ;
  LAYER M1 ;
        RECT 13.344 18.696 13.376 21.204 ;
  LAYER M3 ;
        RECT 13.344 18.716 13.376 18.748 ;
  LAYER M1 ;
        RECT 13.28 18.696 13.312 21.204 ;
  LAYER M3 ;
        RECT 13.28 21.152 13.312 21.184 ;
  LAYER M1 ;
        RECT 13.216 18.696 13.248 21.204 ;
  LAYER M3 ;
        RECT 13.216 18.716 13.248 18.748 ;
  LAYER M1 ;
        RECT 13.152 18.696 13.184 21.204 ;
  LAYER M3 ;
        RECT 13.152 21.152 13.184 21.184 ;
  LAYER M1 ;
        RECT 13.088 18.696 13.12 21.204 ;
  LAYER M3 ;
        RECT 13.088 18.716 13.12 18.748 ;
  LAYER M1 ;
        RECT 13.024 18.696 13.056 21.204 ;
  LAYER M3 ;
        RECT 13.024 21.152 13.056 21.184 ;
  LAYER M1 ;
        RECT 12.96 18.696 12.992 21.204 ;
  LAYER M3 ;
        RECT 12.96 18.716 12.992 18.748 ;
  LAYER M1 ;
        RECT 12.896 18.696 12.928 21.204 ;
  LAYER M3 ;
        RECT 12.896 21.152 12.928 21.184 ;
  LAYER M1 ;
        RECT 12.832 18.696 12.864 21.204 ;
  LAYER M3 ;
        RECT 12.832 18.716 12.864 18.748 ;
  LAYER M1 ;
        RECT 12.768 18.696 12.8 21.204 ;
  LAYER M3 ;
        RECT 12.768 21.152 12.8 21.184 ;
  LAYER M1 ;
        RECT 12.704 18.696 12.736 21.204 ;
  LAYER M3 ;
        RECT 12.704 18.716 12.736 18.748 ;
  LAYER M1 ;
        RECT 12.64 18.696 12.672 21.204 ;
  LAYER M3 ;
        RECT 12.64 21.152 12.672 21.184 ;
  LAYER M1 ;
        RECT 12.576 18.696 12.608 21.204 ;
  LAYER M3 ;
        RECT 12.576 18.716 12.608 18.748 ;
  LAYER M1 ;
        RECT 12.512 18.696 12.544 21.204 ;
  LAYER M3 ;
        RECT 14.88 21.088 14.912 21.12 ;
  LAYER M2 ;
        RECT 12.512 21.024 12.544 21.056 ;
  LAYER M2 ;
        RECT 14.88 20.96 14.912 20.992 ;
  LAYER M2 ;
        RECT 12.512 20.896 12.544 20.928 ;
  LAYER M2 ;
        RECT 14.88 20.832 14.912 20.864 ;
  LAYER M2 ;
        RECT 12.512 20.768 12.544 20.8 ;
  LAYER M2 ;
        RECT 14.88 20.704 14.912 20.736 ;
  LAYER M2 ;
        RECT 12.512 20.64 12.544 20.672 ;
  LAYER M2 ;
        RECT 14.88 20.576 14.912 20.608 ;
  LAYER M2 ;
        RECT 12.512 20.512 12.544 20.544 ;
  LAYER M2 ;
        RECT 14.88 20.448 14.912 20.48 ;
  LAYER M2 ;
        RECT 12.512 20.384 12.544 20.416 ;
  LAYER M2 ;
        RECT 14.88 20.32 14.912 20.352 ;
  LAYER M2 ;
        RECT 12.512 20.256 12.544 20.288 ;
  LAYER M2 ;
        RECT 14.88 20.192 14.912 20.224 ;
  LAYER M2 ;
        RECT 12.512 20.128 12.544 20.16 ;
  LAYER M2 ;
        RECT 14.88 20.064 14.912 20.096 ;
  LAYER M2 ;
        RECT 12.512 20 12.544 20.032 ;
  LAYER M2 ;
        RECT 14.88 19.936 14.912 19.968 ;
  LAYER M2 ;
        RECT 12.512 19.872 12.544 19.904 ;
  LAYER M2 ;
        RECT 14.88 19.808 14.912 19.84 ;
  LAYER M2 ;
        RECT 12.512 19.744 12.544 19.776 ;
  LAYER M2 ;
        RECT 14.88 19.68 14.912 19.712 ;
  LAYER M2 ;
        RECT 12.512 19.616 12.544 19.648 ;
  LAYER M2 ;
        RECT 14.88 19.552 14.912 19.584 ;
  LAYER M2 ;
        RECT 12.512 19.488 12.544 19.52 ;
  LAYER M2 ;
        RECT 14.88 19.424 14.912 19.456 ;
  LAYER M2 ;
        RECT 12.512 19.36 12.544 19.392 ;
  LAYER M2 ;
        RECT 14.88 19.296 14.912 19.328 ;
  LAYER M2 ;
        RECT 12.512 19.232 12.544 19.264 ;
  LAYER M2 ;
        RECT 14.88 19.168 14.912 19.2 ;
  LAYER M2 ;
        RECT 12.512 19.104 12.544 19.136 ;
  LAYER M2 ;
        RECT 14.88 19.04 14.912 19.072 ;
  LAYER M2 ;
        RECT 12.512 18.976 12.544 19.008 ;
  LAYER M2 ;
        RECT 14.88 18.912 14.912 18.944 ;
  LAYER M2 ;
        RECT 12.512 18.848 12.544 18.88 ;
  LAYER M2 ;
        RECT 12.464 18.648 14.96 21.252 ;
  LAYER M1 ;
        RECT 14.88 15.588 14.912 18.096 ;
  LAYER M3 ;
        RECT 14.88 15.608 14.912 15.64 ;
  LAYER M1 ;
        RECT 14.816 15.588 14.848 18.096 ;
  LAYER M3 ;
        RECT 14.816 18.044 14.848 18.076 ;
  LAYER M1 ;
        RECT 14.752 15.588 14.784 18.096 ;
  LAYER M3 ;
        RECT 14.752 15.608 14.784 15.64 ;
  LAYER M1 ;
        RECT 14.688 15.588 14.72 18.096 ;
  LAYER M3 ;
        RECT 14.688 18.044 14.72 18.076 ;
  LAYER M1 ;
        RECT 14.624 15.588 14.656 18.096 ;
  LAYER M3 ;
        RECT 14.624 15.608 14.656 15.64 ;
  LAYER M1 ;
        RECT 14.56 15.588 14.592 18.096 ;
  LAYER M3 ;
        RECT 14.56 18.044 14.592 18.076 ;
  LAYER M1 ;
        RECT 14.496 15.588 14.528 18.096 ;
  LAYER M3 ;
        RECT 14.496 15.608 14.528 15.64 ;
  LAYER M1 ;
        RECT 14.432 15.588 14.464 18.096 ;
  LAYER M3 ;
        RECT 14.432 18.044 14.464 18.076 ;
  LAYER M1 ;
        RECT 14.368 15.588 14.4 18.096 ;
  LAYER M3 ;
        RECT 14.368 15.608 14.4 15.64 ;
  LAYER M1 ;
        RECT 14.304 15.588 14.336 18.096 ;
  LAYER M3 ;
        RECT 14.304 18.044 14.336 18.076 ;
  LAYER M1 ;
        RECT 14.24 15.588 14.272 18.096 ;
  LAYER M3 ;
        RECT 14.24 15.608 14.272 15.64 ;
  LAYER M1 ;
        RECT 14.176 15.588 14.208 18.096 ;
  LAYER M3 ;
        RECT 14.176 18.044 14.208 18.076 ;
  LAYER M1 ;
        RECT 14.112 15.588 14.144 18.096 ;
  LAYER M3 ;
        RECT 14.112 15.608 14.144 15.64 ;
  LAYER M1 ;
        RECT 14.048 15.588 14.08 18.096 ;
  LAYER M3 ;
        RECT 14.048 18.044 14.08 18.076 ;
  LAYER M1 ;
        RECT 13.984 15.588 14.016 18.096 ;
  LAYER M3 ;
        RECT 13.984 15.608 14.016 15.64 ;
  LAYER M1 ;
        RECT 13.92 15.588 13.952 18.096 ;
  LAYER M3 ;
        RECT 13.92 18.044 13.952 18.076 ;
  LAYER M1 ;
        RECT 13.856 15.588 13.888 18.096 ;
  LAYER M3 ;
        RECT 13.856 15.608 13.888 15.64 ;
  LAYER M1 ;
        RECT 13.792 15.588 13.824 18.096 ;
  LAYER M3 ;
        RECT 13.792 18.044 13.824 18.076 ;
  LAYER M1 ;
        RECT 13.728 15.588 13.76 18.096 ;
  LAYER M3 ;
        RECT 13.728 15.608 13.76 15.64 ;
  LAYER M1 ;
        RECT 13.664 15.588 13.696 18.096 ;
  LAYER M3 ;
        RECT 13.664 18.044 13.696 18.076 ;
  LAYER M1 ;
        RECT 13.6 15.588 13.632 18.096 ;
  LAYER M3 ;
        RECT 13.6 15.608 13.632 15.64 ;
  LAYER M1 ;
        RECT 13.536 15.588 13.568 18.096 ;
  LAYER M3 ;
        RECT 13.536 18.044 13.568 18.076 ;
  LAYER M1 ;
        RECT 13.472 15.588 13.504 18.096 ;
  LAYER M3 ;
        RECT 13.472 15.608 13.504 15.64 ;
  LAYER M1 ;
        RECT 13.408 15.588 13.44 18.096 ;
  LAYER M3 ;
        RECT 13.408 18.044 13.44 18.076 ;
  LAYER M1 ;
        RECT 13.344 15.588 13.376 18.096 ;
  LAYER M3 ;
        RECT 13.344 15.608 13.376 15.64 ;
  LAYER M1 ;
        RECT 13.28 15.588 13.312 18.096 ;
  LAYER M3 ;
        RECT 13.28 18.044 13.312 18.076 ;
  LAYER M1 ;
        RECT 13.216 15.588 13.248 18.096 ;
  LAYER M3 ;
        RECT 13.216 15.608 13.248 15.64 ;
  LAYER M1 ;
        RECT 13.152 15.588 13.184 18.096 ;
  LAYER M3 ;
        RECT 13.152 18.044 13.184 18.076 ;
  LAYER M1 ;
        RECT 13.088 15.588 13.12 18.096 ;
  LAYER M3 ;
        RECT 13.088 15.608 13.12 15.64 ;
  LAYER M1 ;
        RECT 13.024 15.588 13.056 18.096 ;
  LAYER M3 ;
        RECT 13.024 18.044 13.056 18.076 ;
  LAYER M1 ;
        RECT 12.96 15.588 12.992 18.096 ;
  LAYER M3 ;
        RECT 12.96 15.608 12.992 15.64 ;
  LAYER M1 ;
        RECT 12.896 15.588 12.928 18.096 ;
  LAYER M3 ;
        RECT 12.896 18.044 12.928 18.076 ;
  LAYER M1 ;
        RECT 12.832 15.588 12.864 18.096 ;
  LAYER M3 ;
        RECT 12.832 15.608 12.864 15.64 ;
  LAYER M1 ;
        RECT 12.768 15.588 12.8 18.096 ;
  LAYER M3 ;
        RECT 12.768 18.044 12.8 18.076 ;
  LAYER M1 ;
        RECT 12.704 15.588 12.736 18.096 ;
  LAYER M3 ;
        RECT 12.704 15.608 12.736 15.64 ;
  LAYER M1 ;
        RECT 12.64 15.588 12.672 18.096 ;
  LAYER M3 ;
        RECT 12.64 18.044 12.672 18.076 ;
  LAYER M1 ;
        RECT 12.576 15.588 12.608 18.096 ;
  LAYER M3 ;
        RECT 12.576 15.608 12.608 15.64 ;
  LAYER M1 ;
        RECT 12.512 15.588 12.544 18.096 ;
  LAYER M3 ;
        RECT 14.88 17.98 14.912 18.012 ;
  LAYER M2 ;
        RECT 12.512 17.916 12.544 17.948 ;
  LAYER M2 ;
        RECT 14.88 17.852 14.912 17.884 ;
  LAYER M2 ;
        RECT 12.512 17.788 12.544 17.82 ;
  LAYER M2 ;
        RECT 14.88 17.724 14.912 17.756 ;
  LAYER M2 ;
        RECT 12.512 17.66 12.544 17.692 ;
  LAYER M2 ;
        RECT 14.88 17.596 14.912 17.628 ;
  LAYER M2 ;
        RECT 12.512 17.532 12.544 17.564 ;
  LAYER M2 ;
        RECT 14.88 17.468 14.912 17.5 ;
  LAYER M2 ;
        RECT 12.512 17.404 12.544 17.436 ;
  LAYER M2 ;
        RECT 14.88 17.34 14.912 17.372 ;
  LAYER M2 ;
        RECT 12.512 17.276 12.544 17.308 ;
  LAYER M2 ;
        RECT 14.88 17.212 14.912 17.244 ;
  LAYER M2 ;
        RECT 12.512 17.148 12.544 17.18 ;
  LAYER M2 ;
        RECT 14.88 17.084 14.912 17.116 ;
  LAYER M2 ;
        RECT 12.512 17.02 12.544 17.052 ;
  LAYER M2 ;
        RECT 14.88 16.956 14.912 16.988 ;
  LAYER M2 ;
        RECT 12.512 16.892 12.544 16.924 ;
  LAYER M2 ;
        RECT 14.88 16.828 14.912 16.86 ;
  LAYER M2 ;
        RECT 12.512 16.764 12.544 16.796 ;
  LAYER M2 ;
        RECT 14.88 16.7 14.912 16.732 ;
  LAYER M2 ;
        RECT 12.512 16.636 12.544 16.668 ;
  LAYER M2 ;
        RECT 14.88 16.572 14.912 16.604 ;
  LAYER M2 ;
        RECT 12.512 16.508 12.544 16.54 ;
  LAYER M2 ;
        RECT 14.88 16.444 14.912 16.476 ;
  LAYER M2 ;
        RECT 12.512 16.38 12.544 16.412 ;
  LAYER M2 ;
        RECT 14.88 16.316 14.912 16.348 ;
  LAYER M2 ;
        RECT 12.512 16.252 12.544 16.284 ;
  LAYER M2 ;
        RECT 14.88 16.188 14.912 16.22 ;
  LAYER M2 ;
        RECT 12.512 16.124 12.544 16.156 ;
  LAYER M2 ;
        RECT 14.88 16.06 14.912 16.092 ;
  LAYER M2 ;
        RECT 12.512 15.996 12.544 16.028 ;
  LAYER M2 ;
        RECT 14.88 15.932 14.912 15.964 ;
  LAYER M2 ;
        RECT 12.512 15.868 12.544 15.9 ;
  LAYER M2 ;
        RECT 14.88 15.804 14.912 15.836 ;
  LAYER M2 ;
        RECT 12.512 15.74 12.544 15.772 ;
  LAYER M2 ;
        RECT 12.464 15.54 14.96 18.144 ;
  LAYER M1 ;
        RECT 11.904 28.02 11.936 30.528 ;
  LAYER M3 ;
        RECT 11.904 28.04 11.936 28.072 ;
  LAYER M1 ;
        RECT 11.84 28.02 11.872 30.528 ;
  LAYER M3 ;
        RECT 11.84 30.476 11.872 30.508 ;
  LAYER M1 ;
        RECT 11.776 28.02 11.808 30.528 ;
  LAYER M3 ;
        RECT 11.776 28.04 11.808 28.072 ;
  LAYER M1 ;
        RECT 11.712 28.02 11.744 30.528 ;
  LAYER M3 ;
        RECT 11.712 30.476 11.744 30.508 ;
  LAYER M1 ;
        RECT 11.648 28.02 11.68 30.528 ;
  LAYER M3 ;
        RECT 11.648 28.04 11.68 28.072 ;
  LAYER M1 ;
        RECT 11.584 28.02 11.616 30.528 ;
  LAYER M3 ;
        RECT 11.584 30.476 11.616 30.508 ;
  LAYER M1 ;
        RECT 11.52 28.02 11.552 30.528 ;
  LAYER M3 ;
        RECT 11.52 28.04 11.552 28.072 ;
  LAYER M1 ;
        RECT 11.456 28.02 11.488 30.528 ;
  LAYER M3 ;
        RECT 11.456 30.476 11.488 30.508 ;
  LAYER M1 ;
        RECT 11.392 28.02 11.424 30.528 ;
  LAYER M3 ;
        RECT 11.392 28.04 11.424 28.072 ;
  LAYER M1 ;
        RECT 11.328 28.02 11.36 30.528 ;
  LAYER M3 ;
        RECT 11.328 30.476 11.36 30.508 ;
  LAYER M1 ;
        RECT 11.264 28.02 11.296 30.528 ;
  LAYER M3 ;
        RECT 11.264 28.04 11.296 28.072 ;
  LAYER M1 ;
        RECT 11.2 28.02 11.232 30.528 ;
  LAYER M3 ;
        RECT 11.2 30.476 11.232 30.508 ;
  LAYER M1 ;
        RECT 11.136 28.02 11.168 30.528 ;
  LAYER M3 ;
        RECT 11.136 28.04 11.168 28.072 ;
  LAYER M1 ;
        RECT 11.072 28.02 11.104 30.528 ;
  LAYER M3 ;
        RECT 11.072 30.476 11.104 30.508 ;
  LAYER M1 ;
        RECT 11.008 28.02 11.04 30.528 ;
  LAYER M3 ;
        RECT 11.008 28.04 11.04 28.072 ;
  LAYER M1 ;
        RECT 10.944 28.02 10.976 30.528 ;
  LAYER M3 ;
        RECT 10.944 30.476 10.976 30.508 ;
  LAYER M1 ;
        RECT 10.88 28.02 10.912 30.528 ;
  LAYER M3 ;
        RECT 10.88 28.04 10.912 28.072 ;
  LAYER M1 ;
        RECT 10.816 28.02 10.848 30.528 ;
  LAYER M3 ;
        RECT 10.816 30.476 10.848 30.508 ;
  LAYER M1 ;
        RECT 10.752 28.02 10.784 30.528 ;
  LAYER M3 ;
        RECT 10.752 28.04 10.784 28.072 ;
  LAYER M1 ;
        RECT 10.688 28.02 10.72 30.528 ;
  LAYER M3 ;
        RECT 10.688 30.476 10.72 30.508 ;
  LAYER M1 ;
        RECT 10.624 28.02 10.656 30.528 ;
  LAYER M3 ;
        RECT 10.624 28.04 10.656 28.072 ;
  LAYER M1 ;
        RECT 10.56 28.02 10.592 30.528 ;
  LAYER M3 ;
        RECT 10.56 30.476 10.592 30.508 ;
  LAYER M1 ;
        RECT 10.496 28.02 10.528 30.528 ;
  LAYER M3 ;
        RECT 10.496 28.04 10.528 28.072 ;
  LAYER M1 ;
        RECT 10.432 28.02 10.464 30.528 ;
  LAYER M3 ;
        RECT 10.432 30.476 10.464 30.508 ;
  LAYER M1 ;
        RECT 10.368 28.02 10.4 30.528 ;
  LAYER M3 ;
        RECT 10.368 28.04 10.4 28.072 ;
  LAYER M1 ;
        RECT 10.304 28.02 10.336 30.528 ;
  LAYER M3 ;
        RECT 10.304 30.476 10.336 30.508 ;
  LAYER M1 ;
        RECT 10.24 28.02 10.272 30.528 ;
  LAYER M3 ;
        RECT 10.24 28.04 10.272 28.072 ;
  LAYER M1 ;
        RECT 10.176 28.02 10.208 30.528 ;
  LAYER M3 ;
        RECT 10.176 30.476 10.208 30.508 ;
  LAYER M1 ;
        RECT 10.112 28.02 10.144 30.528 ;
  LAYER M3 ;
        RECT 10.112 28.04 10.144 28.072 ;
  LAYER M1 ;
        RECT 10.048 28.02 10.08 30.528 ;
  LAYER M3 ;
        RECT 10.048 30.476 10.08 30.508 ;
  LAYER M1 ;
        RECT 9.984 28.02 10.016 30.528 ;
  LAYER M3 ;
        RECT 9.984 28.04 10.016 28.072 ;
  LAYER M1 ;
        RECT 9.92 28.02 9.952 30.528 ;
  LAYER M3 ;
        RECT 9.92 30.476 9.952 30.508 ;
  LAYER M1 ;
        RECT 9.856 28.02 9.888 30.528 ;
  LAYER M3 ;
        RECT 9.856 28.04 9.888 28.072 ;
  LAYER M1 ;
        RECT 9.792 28.02 9.824 30.528 ;
  LAYER M3 ;
        RECT 9.792 30.476 9.824 30.508 ;
  LAYER M1 ;
        RECT 9.728 28.02 9.76 30.528 ;
  LAYER M3 ;
        RECT 9.728 28.04 9.76 28.072 ;
  LAYER M1 ;
        RECT 9.664 28.02 9.696 30.528 ;
  LAYER M3 ;
        RECT 9.664 30.476 9.696 30.508 ;
  LAYER M1 ;
        RECT 9.6 28.02 9.632 30.528 ;
  LAYER M3 ;
        RECT 9.6 28.04 9.632 28.072 ;
  LAYER M1 ;
        RECT 9.536 28.02 9.568 30.528 ;
  LAYER M3 ;
        RECT 11.904 30.412 11.936 30.444 ;
  LAYER M2 ;
        RECT 9.536 30.348 9.568 30.38 ;
  LAYER M2 ;
        RECT 11.904 30.284 11.936 30.316 ;
  LAYER M2 ;
        RECT 9.536 30.22 9.568 30.252 ;
  LAYER M2 ;
        RECT 11.904 30.156 11.936 30.188 ;
  LAYER M2 ;
        RECT 9.536 30.092 9.568 30.124 ;
  LAYER M2 ;
        RECT 11.904 30.028 11.936 30.06 ;
  LAYER M2 ;
        RECT 9.536 29.964 9.568 29.996 ;
  LAYER M2 ;
        RECT 11.904 29.9 11.936 29.932 ;
  LAYER M2 ;
        RECT 9.536 29.836 9.568 29.868 ;
  LAYER M2 ;
        RECT 11.904 29.772 11.936 29.804 ;
  LAYER M2 ;
        RECT 9.536 29.708 9.568 29.74 ;
  LAYER M2 ;
        RECT 11.904 29.644 11.936 29.676 ;
  LAYER M2 ;
        RECT 9.536 29.58 9.568 29.612 ;
  LAYER M2 ;
        RECT 11.904 29.516 11.936 29.548 ;
  LAYER M2 ;
        RECT 9.536 29.452 9.568 29.484 ;
  LAYER M2 ;
        RECT 11.904 29.388 11.936 29.42 ;
  LAYER M2 ;
        RECT 9.536 29.324 9.568 29.356 ;
  LAYER M2 ;
        RECT 11.904 29.26 11.936 29.292 ;
  LAYER M2 ;
        RECT 9.536 29.196 9.568 29.228 ;
  LAYER M2 ;
        RECT 11.904 29.132 11.936 29.164 ;
  LAYER M2 ;
        RECT 9.536 29.068 9.568 29.1 ;
  LAYER M2 ;
        RECT 11.904 29.004 11.936 29.036 ;
  LAYER M2 ;
        RECT 9.536 28.94 9.568 28.972 ;
  LAYER M2 ;
        RECT 11.904 28.876 11.936 28.908 ;
  LAYER M2 ;
        RECT 9.536 28.812 9.568 28.844 ;
  LAYER M2 ;
        RECT 11.904 28.748 11.936 28.78 ;
  LAYER M2 ;
        RECT 9.536 28.684 9.568 28.716 ;
  LAYER M2 ;
        RECT 11.904 28.62 11.936 28.652 ;
  LAYER M2 ;
        RECT 9.536 28.556 9.568 28.588 ;
  LAYER M2 ;
        RECT 11.904 28.492 11.936 28.524 ;
  LAYER M2 ;
        RECT 9.536 28.428 9.568 28.46 ;
  LAYER M2 ;
        RECT 11.904 28.364 11.936 28.396 ;
  LAYER M2 ;
        RECT 9.536 28.3 9.568 28.332 ;
  LAYER M2 ;
        RECT 11.904 28.236 11.936 28.268 ;
  LAYER M2 ;
        RECT 9.536 28.172 9.568 28.204 ;
  LAYER M2 ;
        RECT 9.488 27.972 11.984 30.576 ;
  LAYER M1 ;
        RECT 11.904 24.912 11.936 27.42 ;
  LAYER M3 ;
        RECT 11.904 24.932 11.936 24.964 ;
  LAYER M1 ;
        RECT 11.84 24.912 11.872 27.42 ;
  LAYER M3 ;
        RECT 11.84 27.368 11.872 27.4 ;
  LAYER M1 ;
        RECT 11.776 24.912 11.808 27.42 ;
  LAYER M3 ;
        RECT 11.776 24.932 11.808 24.964 ;
  LAYER M1 ;
        RECT 11.712 24.912 11.744 27.42 ;
  LAYER M3 ;
        RECT 11.712 27.368 11.744 27.4 ;
  LAYER M1 ;
        RECT 11.648 24.912 11.68 27.42 ;
  LAYER M3 ;
        RECT 11.648 24.932 11.68 24.964 ;
  LAYER M1 ;
        RECT 11.584 24.912 11.616 27.42 ;
  LAYER M3 ;
        RECT 11.584 27.368 11.616 27.4 ;
  LAYER M1 ;
        RECT 11.52 24.912 11.552 27.42 ;
  LAYER M3 ;
        RECT 11.52 24.932 11.552 24.964 ;
  LAYER M1 ;
        RECT 11.456 24.912 11.488 27.42 ;
  LAYER M3 ;
        RECT 11.456 27.368 11.488 27.4 ;
  LAYER M1 ;
        RECT 11.392 24.912 11.424 27.42 ;
  LAYER M3 ;
        RECT 11.392 24.932 11.424 24.964 ;
  LAYER M1 ;
        RECT 11.328 24.912 11.36 27.42 ;
  LAYER M3 ;
        RECT 11.328 27.368 11.36 27.4 ;
  LAYER M1 ;
        RECT 11.264 24.912 11.296 27.42 ;
  LAYER M3 ;
        RECT 11.264 24.932 11.296 24.964 ;
  LAYER M1 ;
        RECT 11.2 24.912 11.232 27.42 ;
  LAYER M3 ;
        RECT 11.2 27.368 11.232 27.4 ;
  LAYER M1 ;
        RECT 11.136 24.912 11.168 27.42 ;
  LAYER M3 ;
        RECT 11.136 24.932 11.168 24.964 ;
  LAYER M1 ;
        RECT 11.072 24.912 11.104 27.42 ;
  LAYER M3 ;
        RECT 11.072 27.368 11.104 27.4 ;
  LAYER M1 ;
        RECT 11.008 24.912 11.04 27.42 ;
  LAYER M3 ;
        RECT 11.008 24.932 11.04 24.964 ;
  LAYER M1 ;
        RECT 10.944 24.912 10.976 27.42 ;
  LAYER M3 ;
        RECT 10.944 27.368 10.976 27.4 ;
  LAYER M1 ;
        RECT 10.88 24.912 10.912 27.42 ;
  LAYER M3 ;
        RECT 10.88 24.932 10.912 24.964 ;
  LAYER M1 ;
        RECT 10.816 24.912 10.848 27.42 ;
  LAYER M3 ;
        RECT 10.816 27.368 10.848 27.4 ;
  LAYER M1 ;
        RECT 10.752 24.912 10.784 27.42 ;
  LAYER M3 ;
        RECT 10.752 24.932 10.784 24.964 ;
  LAYER M1 ;
        RECT 10.688 24.912 10.72 27.42 ;
  LAYER M3 ;
        RECT 10.688 27.368 10.72 27.4 ;
  LAYER M1 ;
        RECT 10.624 24.912 10.656 27.42 ;
  LAYER M3 ;
        RECT 10.624 24.932 10.656 24.964 ;
  LAYER M1 ;
        RECT 10.56 24.912 10.592 27.42 ;
  LAYER M3 ;
        RECT 10.56 27.368 10.592 27.4 ;
  LAYER M1 ;
        RECT 10.496 24.912 10.528 27.42 ;
  LAYER M3 ;
        RECT 10.496 24.932 10.528 24.964 ;
  LAYER M1 ;
        RECT 10.432 24.912 10.464 27.42 ;
  LAYER M3 ;
        RECT 10.432 27.368 10.464 27.4 ;
  LAYER M1 ;
        RECT 10.368 24.912 10.4 27.42 ;
  LAYER M3 ;
        RECT 10.368 24.932 10.4 24.964 ;
  LAYER M1 ;
        RECT 10.304 24.912 10.336 27.42 ;
  LAYER M3 ;
        RECT 10.304 27.368 10.336 27.4 ;
  LAYER M1 ;
        RECT 10.24 24.912 10.272 27.42 ;
  LAYER M3 ;
        RECT 10.24 24.932 10.272 24.964 ;
  LAYER M1 ;
        RECT 10.176 24.912 10.208 27.42 ;
  LAYER M3 ;
        RECT 10.176 27.368 10.208 27.4 ;
  LAYER M1 ;
        RECT 10.112 24.912 10.144 27.42 ;
  LAYER M3 ;
        RECT 10.112 24.932 10.144 24.964 ;
  LAYER M1 ;
        RECT 10.048 24.912 10.08 27.42 ;
  LAYER M3 ;
        RECT 10.048 27.368 10.08 27.4 ;
  LAYER M1 ;
        RECT 9.984 24.912 10.016 27.42 ;
  LAYER M3 ;
        RECT 9.984 24.932 10.016 24.964 ;
  LAYER M1 ;
        RECT 9.92 24.912 9.952 27.42 ;
  LAYER M3 ;
        RECT 9.92 27.368 9.952 27.4 ;
  LAYER M1 ;
        RECT 9.856 24.912 9.888 27.42 ;
  LAYER M3 ;
        RECT 9.856 24.932 9.888 24.964 ;
  LAYER M1 ;
        RECT 9.792 24.912 9.824 27.42 ;
  LAYER M3 ;
        RECT 9.792 27.368 9.824 27.4 ;
  LAYER M1 ;
        RECT 9.728 24.912 9.76 27.42 ;
  LAYER M3 ;
        RECT 9.728 24.932 9.76 24.964 ;
  LAYER M1 ;
        RECT 9.664 24.912 9.696 27.42 ;
  LAYER M3 ;
        RECT 9.664 27.368 9.696 27.4 ;
  LAYER M1 ;
        RECT 9.6 24.912 9.632 27.42 ;
  LAYER M3 ;
        RECT 9.6 24.932 9.632 24.964 ;
  LAYER M1 ;
        RECT 9.536 24.912 9.568 27.42 ;
  LAYER M3 ;
        RECT 11.904 27.304 11.936 27.336 ;
  LAYER M2 ;
        RECT 9.536 27.24 9.568 27.272 ;
  LAYER M2 ;
        RECT 11.904 27.176 11.936 27.208 ;
  LAYER M2 ;
        RECT 9.536 27.112 9.568 27.144 ;
  LAYER M2 ;
        RECT 11.904 27.048 11.936 27.08 ;
  LAYER M2 ;
        RECT 9.536 26.984 9.568 27.016 ;
  LAYER M2 ;
        RECT 11.904 26.92 11.936 26.952 ;
  LAYER M2 ;
        RECT 9.536 26.856 9.568 26.888 ;
  LAYER M2 ;
        RECT 11.904 26.792 11.936 26.824 ;
  LAYER M2 ;
        RECT 9.536 26.728 9.568 26.76 ;
  LAYER M2 ;
        RECT 11.904 26.664 11.936 26.696 ;
  LAYER M2 ;
        RECT 9.536 26.6 9.568 26.632 ;
  LAYER M2 ;
        RECT 11.904 26.536 11.936 26.568 ;
  LAYER M2 ;
        RECT 9.536 26.472 9.568 26.504 ;
  LAYER M2 ;
        RECT 11.904 26.408 11.936 26.44 ;
  LAYER M2 ;
        RECT 9.536 26.344 9.568 26.376 ;
  LAYER M2 ;
        RECT 11.904 26.28 11.936 26.312 ;
  LAYER M2 ;
        RECT 9.536 26.216 9.568 26.248 ;
  LAYER M2 ;
        RECT 11.904 26.152 11.936 26.184 ;
  LAYER M2 ;
        RECT 9.536 26.088 9.568 26.12 ;
  LAYER M2 ;
        RECT 11.904 26.024 11.936 26.056 ;
  LAYER M2 ;
        RECT 9.536 25.96 9.568 25.992 ;
  LAYER M2 ;
        RECT 11.904 25.896 11.936 25.928 ;
  LAYER M2 ;
        RECT 9.536 25.832 9.568 25.864 ;
  LAYER M2 ;
        RECT 11.904 25.768 11.936 25.8 ;
  LAYER M2 ;
        RECT 9.536 25.704 9.568 25.736 ;
  LAYER M2 ;
        RECT 11.904 25.64 11.936 25.672 ;
  LAYER M2 ;
        RECT 9.536 25.576 9.568 25.608 ;
  LAYER M2 ;
        RECT 11.904 25.512 11.936 25.544 ;
  LAYER M2 ;
        RECT 9.536 25.448 9.568 25.48 ;
  LAYER M2 ;
        RECT 11.904 25.384 11.936 25.416 ;
  LAYER M2 ;
        RECT 9.536 25.32 9.568 25.352 ;
  LAYER M2 ;
        RECT 11.904 25.256 11.936 25.288 ;
  LAYER M2 ;
        RECT 9.536 25.192 9.568 25.224 ;
  LAYER M2 ;
        RECT 11.904 25.128 11.936 25.16 ;
  LAYER M2 ;
        RECT 9.536 25.064 9.568 25.096 ;
  LAYER M2 ;
        RECT 9.488 24.864 11.984 27.468 ;
  LAYER M1 ;
        RECT 11.904 21.804 11.936 24.312 ;
  LAYER M3 ;
        RECT 11.904 21.824 11.936 21.856 ;
  LAYER M1 ;
        RECT 11.84 21.804 11.872 24.312 ;
  LAYER M3 ;
        RECT 11.84 24.26 11.872 24.292 ;
  LAYER M1 ;
        RECT 11.776 21.804 11.808 24.312 ;
  LAYER M3 ;
        RECT 11.776 21.824 11.808 21.856 ;
  LAYER M1 ;
        RECT 11.712 21.804 11.744 24.312 ;
  LAYER M3 ;
        RECT 11.712 24.26 11.744 24.292 ;
  LAYER M1 ;
        RECT 11.648 21.804 11.68 24.312 ;
  LAYER M3 ;
        RECT 11.648 21.824 11.68 21.856 ;
  LAYER M1 ;
        RECT 11.584 21.804 11.616 24.312 ;
  LAYER M3 ;
        RECT 11.584 24.26 11.616 24.292 ;
  LAYER M1 ;
        RECT 11.52 21.804 11.552 24.312 ;
  LAYER M3 ;
        RECT 11.52 21.824 11.552 21.856 ;
  LAYER M1 ;
        RECT 11.456 21.804 11.488 24.312 ;
  LAYER M3 ;
        RECT 11.456 24.26 11.488 24.292 ;
  LAYER M1 ;
        RECT 11.392 21.804 11.424 24.312 ;
  LAYER M3 ;
        RECT 11.392 21.824 11.424 21.856 ;
  LAYER M1 ;
        RECT 11.328 21.804 11.36 24.312 ;
  LAYER M3 ;
        RECT 11.328 24.26 11.36 24.292 ;
  LAYER M1 ;
        RECT 11.264 21.804 11.296 24.312 ;
  LAYER M3 ;
        RECT 11.264 21.824 11.296 21.856 ;
  LAYER M1 ;
        RECT 11.2 21.804 11.232 24.312 ;
  LAYER M3 ;
        RECT 11.2 24.26 11.232 24.292 ;
  LAYER M1 ;
        RECT 11.136 21.804 11.168 24.312 ;
  LAYER M3 ;
        RECT 11.136 21.824 11.168 21.856 ;
  LAYER M1 ;
        RECT 11.072 21.804 11.104 24.312 ;
  LAYER M3 ;
        RECT 11.072 24.26 11.104 24.292 ;
  LAYER M1 ;
        RECT 11.008 21.804 11.04 24.312 ;
  LAYER M3 ;
        RECT 11.008 21.824 11.04 21.856 ;
  LAYER M1 ;
        RECT 10.944 21.804 10.976 24.312 ;
  LAYER M3 ;
        RECT 10.944 24.26 10.976 24.292 ;
  LAYER M1 ;
        RECT 10.88 21.804 10.912 24.312 ;
  LAYER M3 ;
        RECT 10.88 21.824 10.912 21.856 ;
  LAYER M1 ;
        RECT 10.816 21.804 10.848 24.312 ;
  LAYER M3 ;
        RECT 10.816 24.26 10.848 24.292 ;
  LAYER M1 ;
        RECT 10.752 21.804 10.784 24.312 ;
  LAYER M3 ;
        RECT 10.752 21.824 10.784 21.856 ;
  LAYER M1 ;
        RECT 10.688 21.804 10.72 24.312 ;
  LAYER M3 ;
        RECT 10.688 24.26 10.72 24.292 ;
  LAYER M1 ;
        RECT 10.624 21.804 10.656 24.312 ;
  LAYER M3 ;
        RECT 10.624 21.824 10.656 21.856 ;
  LAYER M1 ;
        RECT 10.56 21.804 10.592 24.312 ;
  LAYER M3 ;
        RECT 10.56 24.26 10.592 24.292 ;
  LAYER M1 ;
        RECT 10.496 21.804 10.528 24.312 ;
  LAYER M3 ;
        RECT 10.496 21.824 10.528 21.856 ;
  LAYER M1 ;
        RECT 10.432 21.804 10.464 24.312 ;
  LAYER M3 ;
        RECT 10.432 24.26 10.464 24.292 ;
  LAYER M1 ;
        RECT 10.368 21.804 10.4 24.312 ;
  LAYER M3 ;
        RECT 10.368 21.824 10.4 21.856 ;
  LAYER M1 ;
        RECT 10.304 21.804 10.336 24.312 ;
  LAYER M3 ;
        RECT 10.304 24.26 10.336 24.292 ;
  LAYER M1 ;
        RECT 10.24 21.804 10.272 24.312 ;
  LAYER M3 ;
        RECT 10.24 21.824 10.272 21.856 ;
  LAYER M1 ;
        RECT 10.176 21.804 10.208 24.312 ;
  LAYER M3 ;
        RECT 10.176 24.26 10.208 24.292 ;
  LAYER M1 ;
        RECT 10.112 21.804 10.144 24.312 ;
  LAYER M3 ;
        RECT 10.112 21.824 10.144 21.856 ;
  LAYER M1 ;
        RECT 10.048 21.804 10.08 24.312 ;
  LAYER M3 ;
        RECT 10.048 24.26 10.08 24.292 ;
  LAYER M1 ;
        RECT 9.984 21.804 10.016 24.312 ;
  LAYER M3 ;
        RECT 9.984 21.824 10.016 21.856 ;
  LAYER M1 ;
        RECT 9.92 21.804 9.952 24.312 ;
  LAYER M3 ;
        RECT 9.92 24.26 9.952 24.292 ;
  LAYER M1 ;
        RECT 9.856 21.804 9.888 24.312 ;
  LAYER M3 ;
        RECT 9.856 21.824 9.888 21.856 ;
  LAYER M1 ;
        RECT 9.792 21.804 9.824 24.312 ;
  LAYER M3 ;
        RECT 9.792 24.26 9.824 24.292 ;
  LAYER M1 ;
        RECT 9.728 21.804 9.76 24.312 ;
  LAYER M3 ;
        RECT 9.728 21.824 9.76 21.856 ;
  LAYER M1 ;
        RECT 9.664 21.804 9.696 24.312 ;
  LAYER M3 ;
        RECT 9.664 24.26 9.696 24.292 ;
  LAYER M1 ;
        RECT 9.6 21.804 9.632 24.312 ;
  LAYER M3 ;
        RECT 9.6 21.824 9.632 21.856 ;
  LAYER M1 ;
        RECT 9.536 21.804 9.568 24.312 ;
  LAYER M3 ;
        RECT 11.904 24.196 11.936 24.228 ;
  LAYER M2 ;
        RECT 9.536 24.132 9.568 24.164 ;
  LAYER M2 ;
        RECT 11.904 24.068 11.936 24.1 ;
  LAYER M2 ;
        RECT 9.536 24.004 9.568 24.036 ;
  LAYER M2 ;
        RECT 11.904 23.94 11.936 23.972 ;
  LAYER M2 ;
        RECT 9.536 23.876 9.568 23.908 ;
  LAYER M2 ;
        RECT 11.904 23.812 11.936 23.844 ;
  LAYER M2 ;
        RECT 9.536 23.748 9.568 23.78 ;
  LAYER M2 ;
        RECT 11.904 23.684 11.936 23.716 ;
  LAYER M2 ;
        RECT 9.536 23.62 9.568 23.652 ;
  LAYER M2 ;
        RECT 11.904 23.556 11.936 23.588 ;
  LAYER M2 ;
        RECT 9.536 23.492 9.568 23.524 ;
  LAYER M2 ;
        RECT 11.904 23.428 11.936 23.46 ;
  LAYER M2 ;
        RECT 9.536 23.364 9.568 23.396 ;
  LAYER M2 ;
        RECT 11.904 23.3 11.936 23.332 ;
  LAYER M2 ;
        RECT 9.536 23.236 9.568 23.268 ;
  LAYER M2 ;
        RECT 11.904 23.172 11.936 23.204 ;
  LAYER M2 ;
        RECT 9.536 23.108 9.568 23.14 ;
  LAYER M2 ;
        RECT 11.904 23.044 11.936 23.076 ;
  LAYER M2 ;
        RECT 9.536 22.98 9.568 23.012 ;
  LAYER M2 ;
        RECT 11.904 22.916 11.936 22.948 ;
  LAYER M2 ;
        RECT 9.536 22.852 9.568 22.884 ;
  LAYER M2 ;
        RECT 11.904 22.788 11.936 22.82 ;
  LAYER M2 ;
        RECT 9.536 22.724 9.568 22.756 ;
  LAYER M2 ;
        RECT 11.904 22.66 11.936 22.692 ;
  LAYER M2 ;
        RECT 9.536 22.596 9.568 22.628 ;
  LAYER M2 ;
        RECT 11.904 22.532 11.936 22.564 ;
  LAYER M2 ;
        RECT 9.536 22.468 9.568 22.5 ;
  LAYER M2 ;
        RECT 11.904 22.404 11.936 22.436 ;
  LAYER M2 ;
        RECT 9.536 22.34 9.568 22.372 ;
  LAYER M2 ;
        RECT 11.904 22.276 11.936 22.308 ;
  LAYER M2 ;
        RECT 9.536 22.212 9.568 22.244 ;
  LAYER M2 ;
        RECT 11.904 22.148 11.936 22.18 ;
  LAYER M2 ;
        RECT 9.536 22.084 9.568 22.116 ;
  LAYER M2 ;
        RECT 11.904 22.02 11.936 22.052 ;
  LAYER M2 ;
        RECT 9.536 21.956 9.568 21.988 ;
  LAYER M2 ;
        RECT 9.488 21.756 11.984 24.36 ;
  LAYER M1 ;
        RECT 11.904 18.696 11.936 21.204 ;
  LAYER M3 ;
        RECT 11.904 18.716 11.936 18.748 ;
  LAYER M1 ;
        RECT 11.84 18.696 11.872 21.204 ;
  LAYER M3 ;
        RECT 11.84 21.152 11.872 21.184 ;
  LAYER M1 ;
        RECT 11.776 18.696 11.808 21.204 ;
  LAYER M3 ;
        RECT 11.776 18.716 11.808 18.748 ;
  LAYER M1 ;
        RECT 11.712 18.696 11.744 21.204 ;
  LAYER M3 ;
        RECT 11.712 21.152 11.744 21.184 ;
  LAYER M1 ;
        RECT 11.648 18.696 11.68 21.204 ;
  LAYER M3 ;
        RECT 11.648 18.716 11.68 18.748 ;
  LAYER M1 ;
        RECT 11.584 18.696 11.616 21.204 ;
  LAYER M3 ;
        RECT 11.584 21.152 11.616 21.184 ;
  LAYER M1 ;
        RECT 11.52 18.696 11.552 21.204 ;
  LAYER M3 ;
        RECT 11.52 18.716 11.552 18.748 ;
  LAYER M1 ;
        RECT 11.456 18.696 11.488 21.204 ;
  LAYER M3 ;
        RECT 11.456 21.152 11.488 21.184 ;
  LAYER M1 ;
        RECT 11.392 18.696 11.424 21.204 ;
  LAYER M3 ;
        RECT 11.392 18.716 11.424 18.748 ;
  LAYER M1 ;
        RECT 11.328 18.696 11.36 21.204 ;
  LAYER M3 ;
        RECT 11.328 21.152 11.36 21.184 ;
  LAYER M1 ;
        RECT 11.264 18.696 11.296 21.204 ;
  LAYER M3 ;
        RECT 11.264 18.716 11.296 18.748 ;
  LAYER M1 ;
        RECT 11.2 18.696 11.232 21.204 ;
  LAYER M3 ;
        RECT 11.2 21.152 11.232 21.184 ;
  LAYER M1 ;
        RECT 11.136 18.696 11.168 21.204 ;
  LAYER M3 ;
        RECT 11.136 18.716 11.168 18.748 ;
  LAYER M1 ;
        RECT 11.072 18.696 11.104 21.204 ;
  LAYER M3 ;
        RECT 11.072 21.152 11.104 21.184 ;
  LAYER M1 ;
        RECT 11.008 18.696 11.04 21.204 ;
  LAYER M3 ;
        RECT 11.008 18.716 11.04 18.748 ;
  LAYER M1 ;
        RECT 10.944 18.696 10.976 21.204 ;
  LAYER M3 ;
        RECT 10.944 21.152 10.976 21.184 ;
  LAYER M1 ;
        RECT 10.88 18.696 10.912 21.204 ;
  LAYER M3 ;
        RECT 10.88 18.716 10.912 18.748 ;
  LAYER M1 ;
        RECT 10.816 18.696 10.848 21.204 ;
  LAYER M3 ;
        RECT 10.816 21.152 10.848 21.184 ;
  LAYER M1 ;
        RECT 10.752 18.696 10.784 21.204 ;
  LAYER M3 ;
        RECT 10.752 18.716 10.784 18.748 ;
  LAYER M1 ;
        RECT 10.688 18.696 10.72 21.204 ;
  LAYER M3 ;
        RECT 10.688 21.152 10.72 21.184 ;
  LAYER M1 ;
        RECT 10.624 18.696 10.656 21.204 ;
  LAYER M3 ;
        RECT 10.624 18.716 10.656 18.748 ;
  LAYER M1 ;
        RECT 10.56 18.696 10.592 21.204 ;
  LAYER M3 ;
        RECT 10.56 21.152 10.592 21.184 ;
  LAYER M1 ;
        RECT 10.496 18.696 10.528 21.204 ;
  LAYER M3 ;
        RECT 10.496 18.716 10.528 18.748 ;
  LAYER M1 ;
        RECT 10.432 18.696 10.464 21.204 ;
  LAYER M3 ;
        RECT 10.432 21.152 10.464 21.184 ;
  LAYER M1 ;
        RECT 10.368 18.696 10.4 21.204 ;
  LAYER M3 ;
        RECT 10.368 18.716 10.4 18.748 ;
  LAYER M1 ;
        RECT 10.304 18.696 10.336 21.204 ;
  LAYER M3 ;
        RECT 10.304 21.152 10.336 21.184 ;
  LAYER M1 ;
        RECT 10.24 18.696 10.272 21.204 ;
  LAYER M3 ;
        RECT 10.24 18.716 10.272 18.748 ;
  LAYER M1 ;
        RECT 10.176 18.696 10.208 21.204 ;
  LAYER M3 ;
        RECT 10.176 21.152 10.208 21.184 ;
  LAYER M1 ;
        RECT 10.112 18.696 10.144 21.204 ;
  LAYER M3 ;
        RECT 10.112 18.716 10.144 18.748 ;
  LAYER M1 ;
        RECT 10.048 18.696 10.08 21.204 ;
  LAYER M3 ;
        RECT 10.048 21.152 10.08 21.184 ;
  LAYER M1 ;
        RECT 9.984 18.696 10.016 21.204 ;
  LAYER M3 ;
        RECT 9.984 18.716 10.016 18.748 ;
  LAYER M1 ;
        RECT 9.92 18.696 9.952 21.204 ;
  LAYER M3 ;
        RECT 9.92 21.152 9.952 21.184 ;
  LAYER M1 ;
        RECT 9.856 18.696 9.888 21.204 ;
  LAYER M3 ;
        RECT 9.856 18.716 9.888 18.748 ;
  LAYER M1 ;
        RECT 9.792 18.696 9.824 21.204 ;
  LAYER M3 ;
        RECT 9.792 21.152 9.824 21.184 ;
  LAYER M1 ;
        RECT 9.728 18.696 9.76 21.204 ;
  LAYER M3 ;
        RECT 9.728 18.716 9.76 18.748 ;
  LAYER M1 ;
        RECT 9.664 18.696 9.696 21.204 ;
  LAYER M3 ;
        RECT 9.664 21.152 9.696 21.184 ;
  LAYER M1 ;
        RECT 9.6 18.696 9.632 21.204 ;
  LAYER M3 ;
        RECT 9.6 18.716 9.632 18.748 ;
  LAYER M1 ;
        RECT 9.536 18.696 9.568 21.204 ;
  LAYER M3 ;
        RECT 11.904 21.088 11.936 21.12 ;
  LAYER M2 ;
        RECT 9.536 21.024 9.568 21.056 ;
  LAYER M2 ;
        RECT 11.904 20.96 11.936 20.992 ;
  LAYER M2 ;
        RECT 9.536 20.896 9.568 20.928 ;
  LAYER M2 ;
        RECT 11.904 20.832 11.936 20.864 ;
  LAYER M2 ;
        RECT 9.536 20.768 9.568 20.8 ;
  LAYER M2 ;
        RECT 11.904 20.704 11.936 20.736 ;
  LAYER M2 ;
        RECT 9.536 20.64 9.568 20.672 ;
  LAYER M2 ;
        RECT 11.904 20.576 11.936 20.608 ;
  LAYER M2 ;
        RECT 9.536 20.512 9.568 20.544 ;
  LAYER M2 ;
        RECT 11.904 20.448 11.936 20.48 ;
  LAYER M2 ;
        RECT 9.536 20.384 9.568 20.416 ;
  LAYER M2 ;
        RECT 11.904 20.32 11.936 20.352 ;
  LAYER M2 ;
        RECT 9.536 20.256 9.568 20.288 ;
  LAYER M2 ;
        RECT 11.904 20.192 11.936 20.224 ;
  LAYER M2 ;
        RECT 9.536 20.128 9.568 20.16 ;
  LAYER M2 ;
        RECT 11.904 20.064 11.936 20.096 ;
  LAYER M2 ;
        RECT 9.536 20 9.568 20.032 ;
  LAYER M2 ;
        RECT 11.904 19.936 11.936 19.968 ;
  LAYER M2 ;
        RECT 9.536 19.872 9.568 19.904 ;
  LAYER M2 ;
        RECT 11.904 19.808 11.936 19.84 ;
  LAYER M2 ;
        RECT 9.536 19.744 9.568 19.776 ;
  LAYER M2 ;
        RECT 11.904 19.68 11.936 19.712 ;
  LAYER M2 ;
        RECT 9.536 19.616 9.568 19.648 ;
  LAYER M2 ;
        RECT 11.904 19.552 11.936 19.584 ;
  LAYER M2 ;
        RECT 9.536 19.488 9.568 19.52 ;
  LAYER M2 ;
        RECT 11.904 19.424 11.936 19.456 ;
  LAYER M2 ;
        RECT 9.536 19.36 9.568 19.392 ;
  LAYER M2 ;
        RECT 11.904 19.296 11.936 19.328 ;
  LAYER M2 ;
        RECT 9.536 19.232 9.568 19.264 ;
  LAYER M2 ;
        RECT 11.904 19.168 11.936 19.2 ;
  LAYER M2 ;
        RECT 9.536 19.104 9.568 19.136 ;
  LAYER M2 ;
        RECT 11.904 19.04 11.936 19.072 ;
  LAYER M2 ;
        RECT 9.536 18.976 9.568 19.008 ;
  LAYER M2 ;
        RECT 11.904 18.912 11.936 18.944 ;
  LAYER M2 ;
        RECT 9.536 18.848 9.568 18.88 ;
  LAYER M2 ;
        RECT 9.488 18.648 11.984 21.252 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M3 ;
        RECT 11.904 15.608 11.936 15.64 ;
  LAYER M1 ;
        RECT 11.84 15.588 11.872 18.096 ;
  LAYER M3 ;
        RECT 11.84 18.044 11.872 18.076 ;
  LAYER M1 ;
        RECT 11.776 15.588 11.808 18.096 ;
  LAYER M3 ;
        RECT 11.776 15.608 11.808 15.64 ;
  LAYER M1 ;
        RECT 11.712 15.588 11.744 18.096 ;
  LAYER M3 ;
        RECT 11.712 18.044 11.744 18.076 ;
  LAYER M1 ;
        RECT 11.648 15.588 11.68 18.096 ;
  LAYER M3 ;
        RECT 11.648 15.608 11.68 15.64 ;
  LAYER M1 ;
        RECT 11.584 15.588 11.616 18.096 ;
  LAYER M3 ;
        RECT 11.584 18.044 11.616 18.076 ;
  LAYER M1 ;
        RECT 11.52 15.588 11.552 18.096 ;
  LAYER M3 ;
        RECT 11.52 15.608 11.552 15.64 ;
  LAYER M1 ;
        RECT 11.456 15.588 11.488 18.096 ;
  LAYER M3 ;
        RECT 11.456 18.044 11.488 18.076 ;
  LAYER M1 ;
        RECT 11.392 15.588 11.424 18.096 ;
  LAYER M3 ;
        RECT 11.392 15.608 11.424 15.64 ;
  LAYER M1 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M3 ;
        RECT 11.328 18.044 11.36 18.076 ;
  LAYER M1 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M3 ;
        RECT 11.264 15.608 11.296 15.64 ;
  LAYER M1 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M3 ;
        RECT 11.2 18.044 11.232 18.076 ;
  LAYER M1 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M3 ;
        RECT 11.136 15.608 11.168 15.64 ;
  LAYER M1 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M3 ;
        RECT 11.072 18.044 11.104 18.076 ;
  LAYER M1 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M3 ;
        RECT 11.008 15.608 11.04 15.64 ;
  LAYER M1 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M3 ;
        RECT 10.944 18.044 10.976 18.076 ;
  LAYER M1 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M3 ;
        RECT 10.88 15.608 10.912 15.64 ;
  LAYER M1 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M3 ;
        RECT 10.816 18.044 10.848 18.076 ;
  LAYER M1 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M3 ;
        RECT 10.752 15.608 10.784 15.64 ;
  LAYER M1 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M3 ;
        RECT 10.688 18.044 10.72 18.076 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M3 ;
        RECT 10.624 15.608 10.656 15.64 ;
  LAYER M1 ;
        RECT 10.56 15.588 10.592 18.096 ;
  LAYER M3 ;
        RECT 10.56 18.044 10.592 18.076 ;
  LAYER M1 ;
        RECT 10.496 15.588 10.528 18.096 ;
  LAYER M3 ;
        RECT 10.496 15.608 10.528 15.64 ;
  LAYER M1 ;
        RECT 10.432 15.588 10.464 18.096 ;
  LAYER M3 ;
        RECT 10.432 18.044 10.464 18.076 ;
  LAYER M1 ;
        RECT 10.368 15.588 10.4 18.096 ;
  LAYER M3 ;
        RECT 10.368 15.608 10.4 15.64 ;
  LAYER M1 ;
        RECT 10.304 15.588 10.336 18.096 ;
  LAYER M3 ;
        RECT 10.304 18.044 10.336 18.076 ;
  LAYER M1 ;
        RECT 10.24 15.588 10.272 18.096 ;
  LAYER M3 ;
        RECT 10.24 15.608 10.272 15.64 ;
  LAYER M1 ;
        RECT 10.176 15.588 10.208 18.096 ;
  LAYER M3 ;
        RECT 10.176 18.044 10.208 18.076 ;
  LAYER M1 ;
        RECT 10.112 15.588 10.144 18.096 ;
  LAYER M3 ;
        RECT 10.112 15.608 10.144 15.64 ;
  LAYER M1 ;
        RECT 10.048 15.588 10.08 18.096 ;
  LAYER M3 ;
        RECT 10.048 18.044 10.08 18.076 ;
  LAYER M1 ;
        RECT 9.984 15.588 10.016 18.096 ;
  LAYER M3 ;
        RECT 9.984 15.608 10.016 15.64 ;
  LAYER M1 ;
        RECT 9.92 15.588 9.952 18.096 ;
  LAYER M3 ;
        RECT 9.92 18.044 9.952 18.076 ;
  LAYER M1 ;
        RECT 9.856 15.588 9.888 18.096 ;
  LAYER M3 ;
        RECT 9.856 15.608 9.888 15.64 ;
  LAYER M1 ;
        RECT 9.792 15.588 9.824 18.096 ;
  LAYER M3 ;
        RECT 9.792 18.044 9.824 18.076 ;
  LAYER M1 ;
        RECT 9.728 15.588 9.76 18.096 ;
  LAYER M3 ;
        RECT 9.728 15.608 9.76 15.64 ;
  LAYER M1 ;
        RECT 9.664 15.588 9.696 18.096 ;
  LAYER M3 ;
        RECT 9.664 18.044 9.696 18.076 ;
  LAYER M1 ;
        RECT 9.6 15.588 9.632 18.096 ;
  LAYER M3 ;
        RECT 9.6 15.608 9.632 15.64 ;
  LAYER M1 ;
        RECT 9.536 15.588 9.568 18.096 ;
  LAYER M3 ;
        RECT 11.904 17.98 11.936 18.012 ;
  LAYER M2 ;
        RECT 9.536 17.916 9.568 17.948 ;
  LAYER M2 ;
        RECT 11.904 17.852 11.936 17.884 ;
  LAYER M2 ;
        RECT 9.536 17.788 9.568 17.82 ;
  LAYER M2 ;
        RECT 11.904 17.724 11.936 17.756 ;
  LAYER M2 ;
        RECT 9.536 17.66 9.568 17.692 ;
  LAYER M2 ;
        RECT 11.904 17.596 11.936 17.628 ;
  LAYER M2 ;
        RECT 9.536 17.532 9.568 17.564 ;
  LAYER M2 ;
        RECT 11.904 17.468 11.936 17.5 ;
  LAYER M2 ;
        RECT 9.536 17.404 9.568 17.436 ;
  LAYER M2 ;
        RECT 11.904 17.34 11.936 17.372 ;
  LAYER M2 ;
        RECT 9.536 17.276 9.568 17.308 ;
  LAYER M2 ;
        RECT 11.904 17.212 11.936 17.244 ;
  LAYER M2 ;
        RECT 9.536 17.148 9.568 17.18 ;
  LAYER M2 ;
        RECT 11.904 17.084 11.936 17.116 ;
  LAYER M2 ;
        RECT 9.536 17.02 9.568 17.052 ;
  LAYER M2 ;
        RECT 11.904 16.956 11.936 16.988 ;
  LAYER M2 ;
        RECT 9.536 16.892 9.568 16.924 ;
  LAYER M2 ;
        RECT 11.904 16.828 11.936 16.86 ;
  LAYER M2 ;
        RECT 9.536 16.764 9.568 16.796 ;
  LAYER M2 ;
        RECT 11.904 16.7 11.936 16.732 ;
  LAYER M2 ;
        RECT 9.536 16.636 9.568 16.668 ;
  LAYER M2 ;
        RECT 11.904 16.572 11.936 16.604 ;
  LAYER M2 ;
        RECT 9.536 16.508 9.568 16.54 ;
  LAYER M2 ;
        RECT 11.904 16.444 11.936 16.476 ;
  LAYER M2 ;
        RECT 9.536 16.38 9.568 16.412 ;
  LAYER M2 ;
        RECT 11.904 16.316 11.936 16.348 ;
  LAYER M2 ;
        RECT 9.536 16.252 9.568 16.284 ;
  LAYER M2 ;
        RECT 11.904 16.188 11.936 16.22 ;
  LAYER M2 ;
        RECT 9.536 16.124 9.568 16.156 ;
  LAYER M2 ;
        RECT 11.904 16.06 11.936 16.092 ;
  LAYER M2 ;
        RECT 9.536 15.996 9.568 16.028 ;
  LAYER M2 ;
        RECT 11.904 15.932 11.936 15.964 ;
  LAYER M2 ;
        RECT 9.536 15.868 9.568 15.9 ;
  LAYER M2 ;
        RECT 11.904 15.804 11.936 15.836 ;
  LAYER M2 ;
        RECT 9.536 15.74 9.568 15.772 ;
  LAYER M2 ;
        RECT 9.488 15.54 11.984 18.144 ;
  LAYER M1 ;
        RECT 8.928 28.02 8.96 30.528 ;
  LAYER M3 ;
        RECT 8.928 28.04 8.96 28.072 ;
  LAYER M1 ;
        RECT 8.864 28.02 8.896 30.528 ;
  LAYER M3 ;
        RECT 8.864 30.476 8.896 30.508 ;
  LAYER M1 ;
        RECT 8.8 28.02 8.832 30.528 ;
  LAYER M3 ;
        RECT 8.8 28.04 8.832 28.072 ;
  LAYER M1 ;
        RECT 8.736 28.02 8.768 30.528 ;
  LAYER M3 ;
        RECT 8.736 30.476 8.768 30.508 ;
  LAYER M1 ;
        RECT 8.672 28.02 8.704 30.528 ;
  LAYER M3 ;
        RECT 8.672 28.04 8.704 28.072 ;
  LAYER M1 ;
        RECT 8.608 28.02 8.64 30.528 ;
  LAYER M3 ;
        RECT 8.608 30.476 8.64 30.508 ;
  LAYER M1 ;
        RECT 8.544 28.02 8.576 30.528 ;
  LAYER M3 ;
        RECT 8.544 28.04 8.576 28.072 ;
  LAYER M1 ;
        RECT 8.48 28.02 8.512 30.528 ;
  LAYER M3 ;
        RECT 8.48 30.476 8.512 30.508 ;
  LAYER M1 ;
        RECT 8.416 28.02 8.448 30.528 ;
  LAYER M3 ;
        RECT 8.416 28.04 8.448 28.072 ;
  LAYER M1 ;
        RECT 8.352 28.02 8.384 30.528 ;
  LAYER M3 ;
        RECT 8.352 30.476 8.384 30.508 ;
  LAYER M1 ;
        RECT 8.288 28.02 8.32 30.528 ;
  LAYER M3 ;
        RECT 8.288 28.04 8.32 28.072 ;
  LAYER M1 ;
        RECT 8.224 28.02 8.256 30.528 ;
  LAYER M3 ;
        RECT 8.224 30.476 8.256 30.508 ;
  LAYER M1 ;
        RECT 8.16 28.02 8.192 30.528 ;
  LAYER M3 ;
        RECT 8.16 28.04 8.192 28.072 ;
  LAYER M1 ;
        RECT 8.096 28.02 8.128 30.528 ;
  LAYER M3 ;
        RECT 8.096 30.476 8.128 30.508 ;
  LAYER M1 ;
        RECT 8.032 28.02 8.064 30.528 ;
  LAYER M3 ;
        RECT 8.032 28.04 8.064 28.072 ;
  LAYER M1 ;
        RECT 7.968 28.02 8 30.528 ;
  LAYER M3 ;
        RECT 7.968 30.476 8 30.508 ;
  LAYER M1 ;
        RECT 7.904 28.02 7.936 30.528 ;
  LAYER M3 ;
        RECT 7.904 28.04 7.936 28.072 ;
  LAYER M1 ;
        RECT 7.84 28.02 7.872 30.528 ;
  LAYER M3 ;
        RECT 7.84 30.476 7.872 30.508 ;
  LAYER M1 ;
        RECT 7.776 28.02 7.808 30.528 ;
  LAYER M3 ;
        RECT 7.776 28.04 7.808 28.072 ;
  LAYER M1 ;
        RECT 7.712 28.02 7.744 30.528 ;
  LAYER M3 ;
        RECT 7.712 30.476 7.744 30.508 ;
  LAYER M1 ;
        RECT 7.648 28.02 7.68 30.528 ;
  LAYER M3 ;
        RECT 7.648 28.04 7.68 28.072 ;
  LAYER M1 ;
        RECT 7.584 28.02 7.616 30.528 ;
  LAYER M3 ;
        RECT 7.584 30.476 7.616 30.508 ;
  LAYER M1 ;
        RECT 7.52 28.02 7.552 30.528 ;
  LAYER M3 ;
        RECT 7.52 28.04 7.552 28.072 ;
  LAYER M1 ;
        RECT 7.456 28.02 7.488 30.528 ;
  LAYER M3 ;
        RECT 7.456 30.476 7.488 30.508 ;
  LAYER M1 ;
        RECT 7.392 28.02 7.424 30.528 ;
  LAYER M3 ;
        RECT 7.392 28.04 7.424 28.072 ;
  LAYER M1 ;
        RECT 7.328 28.02 7.36 30.528 ;
  LAYER M3 ;
        RECT 7.328 30.476 7.36 30.508 ;
  LAYER M1 ;
        RECT 7.264 28.02 7.296 30.528 ;
  LAYER M3 ;
        RECT 7.264 28.04 7.296 28.072 ;
  LAYER M1 ;
        RECT 7.2 28.02 7.232 30.528 ;
  LAYER M3 ;
        RECT 7.2 30.476 7.232 30.508 ;
  LAYER M1 ;
        RECT 7.136 28.02 7.168 30.528 ;
  LAYER M3 ;
        RECT 7.136 28.04 7.168 28.072 ;
  LAYER M1 ;
        RECT 7.072 28.02 7.104 30.528 ;
  LAYER M3 ;
        RECT 7.072 30.476 7.104 30.508 ;
  LAYER M1 ;
        RECT 7.008 28.02 7.04 30.528 ;
  LAYER M3 ;
        RECT 7.008 28.04 7.04 28.072 ;
  LAYER M1 ;
        RECT 6.944 28.02 6.976 30.528 ;
  LAYER M3 ;
        RECT 6.944 30.476 6.976 30.508 ;
  LAYER M1 ;
        RECT 6.88 28.02 6.912 30.528 ;
  LAYER M3 ;
        RECT 6.88 28.04 6.912 28.072 ;
  LAYER M1 ;
        RECT 6.816 28.02 6.848 30.528 ;
  LAYER M3 ;
        RECT 6.816 30.476 6.848 30.508 ;
  LAYER M1 ;
        RECT 6.752 28.02 6.784 30.528 ;
  LAYER M3 ;
        RECT 6.752 28.04 6.784 28.072 ;
  LAYER M1 ;
        RECT 6.688 28.02 6.72 30.528 ;
  LAYER M3 ;
        RECT 6.688 30.476 6.72 30.508 ;
  LAYER M1 ;
        RECT 6.624 28.02 6.656 30.528 ;
  LAYER M3 ;
        RECT 6.624 28.04 6.656 28.072 ;
  LAYER M1 ;
        RECT 6.56 28.02 6.592 30.528 ;
  LAYER M3 ;
        RECT 8.928 30.412 8.96 30.444 ;
  LAYER M2 ;
        RECT 6.56 30.348 6.592 30.38 ;
  LAYER M2 ;
        RECT 8.928 30.284 8.96 30.316 ;
  LAYER M2 ;
        RECT 6.56 30.22 6.592 30.252 ;
  LAYER M2 ;
        RECT 8.928 30.156 8.96 30.188 ;
  LAYER M2 ;
        RECT 6.56 30.092 6.592 30.124 ;
  LAYER M2 ;
        RECT 8.928 30.028 8.96 30.06 ;
  LAYER M2 ;
        RECT 6.56 29.964 6.592 29.996 ;
  LAYER M2 ;
        RECT 8.928 29.9 8.96 29.932 ;
  LAYER M2 ;
        RECT 6.56 29.836 6.592 29.868 ;
  LAYER M2 ;
        RECT 8.928 29.772 8.96 29.804 ;
  LAYER M2 ;
        RECT 6.56 29.708 6.592 29.74 ;
  LAYER M2 ;
        RECT 8.928 29.644 8.96 29.676 ;
  LAYER M2 ;
        RECT 6.56 29.58 6.592 29.612 ;
  LAYER M2 ;
        RECT 8.928 29.516 8.96 29.548 ;
  LAYER M2 ;
        RECT 6.56 29.452 6.592 29.484 ;
  LAYER M2 ;
        RECT 8.928 29.388 8.96 29.42 ;
  LAYER M2 ;
        RECT 6.56 29.324 6.592 29.356 ;
  LAYER M2 ;
        RECT 8.928 29.26 8.96 29.292 ;
  LAYER M2 ;
        RECT 6.56 29.196 6.592 29.228 ;
  LAYER M2 ;
        RECT 8.928 29.132 8.96 29.164 ;
  LAYER M2 ;
        RECT 6.56 29.068 6.592 29.1 ;
  LAYER M2 ;
        RECT 8.928 29.004 8.96 29.036 ;
  LAYER M2 ;
        RECT 6.56 28.94 6.592 28.972 ;
  LAYER M2 ;
        RECT 8.928 28.876 8.96 28.908 ;
  LAYER M2 ;
        RECT 6.56 28.812 6.592 28.844 ;
  LAYER M2 ;
        RECT 8.928 28.748 8.96 28.78 ;
  LAYER M2 ;
        RECT 6.56 28.684 6.592 28.716 ;
  LAYER M2 ;
        RECT 8.928 28.62 8.96 28.652 ;
  LAYER M2 ;
        RECT 6.56 28.556 6.592 28.588 ;
  LAYER M2 ;
        RECT 8.928 28.492 8.96 28.524 ;
  LAYER M2 ;
        RECT 6.56 28.428 6.592 28.46 ;
  LAYER M2 ;
        RECT 8.928 28.364 8.96 28.396 ;
  LAYER M2 ;
        RECT 6.56 28.3 6.592 28.332 ;
  LAYER M2 ;
        RECT 8.928 28.236 8.96 28.268 ;
  LAYER M2 ;
        RECT 6.56 28.172 6.592 28.204 ;
  LAYER M2 ;
        RECT 6.512 27.972 9.008 30.576 ;
  LAYER M1 ;
        RECT 8.928 24.912 8.96 27.42 ;
  LAYER M3 ;
        RECT 8.928 24.932 8.96 24.964 ;
  LAYER M1 ;
        RECT 8.864 24.912 8.896 27.42 ;
  LAYER M3 ;
        RECT 8.864 27.368 8.896 27.4 ;
  LAYER M1 ;
        RECT 8.8 24.912 8.832 27.42 ;
  LAYER M3 ;
        RECT 8.8 24.932 8.832 24.964 ;
  LAYER M1 ;
        RECT 8.736 24.912 8.768 27.42 ;
  LAYER M3 ;
        RECT 8.736 27.368 8.768 27.4 ;
  LAYER M1 ;
        RECT 8.672 24.912 8.704 27.42 ;
  LAYER M3 ;
        RECT 8.672 24.932 8.704 24.964 ;
  LAYER M1 ;
        RECT 8.608 24.912 8.64 27.42 ;
  LAYER M3 ;
        RECT 8.608 27.368 8.64 27.4 ;
  LAYER M1 ;
        RECT 8.544 24.912 8.576 27.42 ;
  LAYER M3 ;
        RECT 8.544 24.932 8.576 24.964 ;
  LAYER M1 ;
        RECT 8.48 24.912 8.512 27.42 ;
  LAYER M3 ;
        RECT 8.48 27.368 8.512 27.4 ;
  LAYER M1 ;
        RECT 8.416 24.912 8.448 27.42 ;
  LAYER M3 ;
        RECT 8.416 24.932 8.448 24.964 ;
  LAYER M1 ;
        RECT 8.352 24.912 8.384 27.42 ;
  LAYER M3 ;
        RECT 8.352 27.368 8.384 27.4 ;
  LAYER M1 ;
        RECT 8.288 24.912 8.32 27.42 ;
  LAYER M3 ;
        RECT 8.288 24.932 8.32 24.964 ;
  LAYER M1 ;
        RECT 8.224 24.912 8.256 27.42 ;
  LAYER M3 ;
        RECT 8.224 27.368 8.256 27.4 ;
  LAYER M1 ;
        RECT 8.16 24.912 8.192 27.42 ;
  LAYER M3 ;
        RECT 8.16 24.932 8.192 24.964 ;
  LAYER M1 ;
        RECT 8.096 24.912 8.128 27.42 ;
  LAYER M3 ;
        RECT 8.096 27.368 8.128 27.4 ;
  LAYER M1 ;
        RECT 8.032 24.912 8.064 27.42 ;
  LAYER M3 ;
        RECT 8.032 24.932 8.064 24.964 ;
  LAYER M1 ;
        RECT 7.968 24.912 8 27.42 ;
  LAYER M3 ;
        RECT 7.968 27.368 8 27.4 ;
  LAYER M1 ;
        RECT 7.904 24.912 7.936 27.42 ;
  LAYER M3 ;
        RECT 7.904 24.932 7.936 24.964 ;
  LAYER M1 ;
        RECT 7.84 24.912 7.872 27.42 ;
  LAYER M3 ;
        RECT 7.84 27.368 7.872 27.4 ;
  LAYER M1 ;
        RECT 7.776 24.912 7.808 27.42 ;
  LAYER M3 ;
        RECT 7.776 24.932 7.808 24.964 ;
  LAYER M1 ;
        RECT 7.712 24.912 7.744 27.42 ;
  LAYER M3 ;
        RECT 7.712 27.368 7.744 27.4 ;
  LAYER M1 ;
        RECT 7.648 24.912 7.68 27.42 ;
  LAYER M3 ;
        RECT 7.648 24.932 7.68 24.964 ;
  LAYER M1 ;
        RECT 7.584 24.912 7.616 27.42 ;
  LAYER M3 ;
        RECT 7.584 27.368 7.616 27.4 ;
  LAYER M1 ;
        RECT 7.52 24.912 7.552 27.42 ;
  LAYER M3 ;
        RECT 7.52 24.932 7.552 24.964 ;
  LAYER M1 ;
        RECT 7.456 24.912 7.488 27.42 ;
  LAYER M3 ;
        RECT 7.456 27.368 7.488 27.4 ;
  LAYER M1 ;
        RECT 7.392 24.912 7.424 27.42 ;
  LAYER M3 ;
        RECT 7.392 24.932 7.424 24.964 ;
  LAYER M1 ;
        RECT 7.328 24.912 7.36 27.42 ;
  LAYER M3 ;
        RECT 7.328 27.368 7.36 27.4 ;
  LAYER M1 ;
        RECT 7.264 24.912 7.296 27.42 ;
  LAYER M3 ;
        RECT 7.264 24.932 7.296 24.964 ;
  LAYER M1 ;
        RECT 7.2 24.912 7.232 27.42 ;
  LAYER M3 ;
        RECT 7.2 27.368 7.232 27.4 ;
  LAYER M1 ;
        RECT 7.136 24.912 7.168 27.42 ;
  LAYER M3 ;
        RECT 7.136 24.932 7.168 24.964 ;
  LAYER M1 ;
        RECT 7.072 24.912 7.104 27.42 ;
  LAYER M3 ;
        RECT 7.072 27.368 7.104 27.4 ;
  LAYER M1 ;
        RECT 7.008 24.912 7.04 27.42 ;
  LAYER M3 ;
        RECT 7.008 24.932 7.04 24.964 ;
  LAYER M1 ;
        RECT 6.944 24.912 6.976 27.42 ;
  LAYER M3 ;
        RECT 6.944 27.368 6.976 27.4 ;
  LAYER M1 ;
        RECT 6.88 24.912 6.912 27.42 ;
  LAYER M3 ;
        RECT 6.88 24.932 6.912 24.964 ;
  LAYER M1 ;
        RECT 6.816 24.912 6.848 27.42 ;
  LAYER M3 ;
        RECT 6.816 27.368 6.848 27.4 ;
  LAYER M1 ;
        RECT 6.752 24.912 6.784 27.42 ;
  LAYER M3 ;
        RECT 6.752 24.932 6.784 24.964 ;
  LAYER M1 ;
        RECT 6.688 24.912 6.72 27.42 ;
  LAYER M3 ;
        RECT 6.688 27.368 6.72 27.4 ;
  LAYER M1 ;
        RECT 6.624 24.912 6.656 27.42 ;
  LAYER M3 ;
        RECT 6.624 24.932 6.656 24.964 ;
  LAYER M1 ;
        RECT 6.56 24.912 6.592 27.42 ;
  LAYER M3 ;
        RECT 8.928 27.304 8.96 27.336 ;
  LAYER M2 ;
        RECT 6.56 27.24 6.592 27.272 ;
  LAYER M2 ;
        RECT 8.928 27.176 8.96 27.208 ;
  LAYER M2 ;
        RECT 6.56 27.112 6.592 27.144 ;
  LAYER M2 ;
        RECT 8.928 27.048 8.96 27.08 ;
  LAYER M2 ;
        RECT 6.56 26.984 6.592 27.016 ;
  LAYER M2 ;
        RECT 8.928 26.92 8.96 26.952 ;
  LAYER M2 ;
        RECT 6.56 26.856 6.592 26.888 ;
  LAYER M2 ;
        RECT 8.928 26.792 8.96 26.824 ;
  LAYER M2 ;
        RECT 6.56 26.728 6.592 26.76 ;
  LAYER M2 ;
        RECT 8.928 26.664 8.96 26.696 ;
  LAYER M2 ;
        RECT 6.56 26.6 6.592 26.632 ;
  LAYER M2 ;
        RECT 8.928 26.536 8.96 26.568 ;
  LAYER M2 ;
        RECT 6.56 26.472 6.592 26.504 ;
  LAYER M2 ;
        RECT 8.928 26.408 8.96 26.44 ;
  LAYER M2 ;
        RECT 6.56 26.344 6.592 26.376 ;
  LAYER M2 ;
        RECT 8.928 26.28 8.96 26.312 ;
  LAYER M2 ;
        RECT 6.56 26.216 6.592 26.248 ;
  LAYER M2 ;
        RECT 8.928 26.152 8.96 26.184 ;
  LAYER M2 ;
        RECT 6.56 26.088 6.592 26.12 ;
  LAYER M2 ;
        RECT 8.928 26.024 8.96 26.056 ;
  LAYER M2 ;
        RECT 6.56 25.96 6.592 25.992 ;
  LAYER M2 ;
        RECT 8.928 25.896 8.96 25.928 ;
  LAYER M2 ;
        RECT 6.56 25.832 6.592 25.864 ;
  LAYER M2 ;
        RECT 8.928 25.768 8.96 25.8 ;
  LAYER M2 ;
        RECT 6.56 25.704 6.592 25.736 ;
  LAYER M2 ;
        RECT 8.928 25.64 8.96 25.672 ;
  LAYER M2 ;
        RECT 6.56 25.576 6.592 25.608 ;
  LAYER M2 ;
        RECT 8.928 25.512 8.96 25.544 ;
  LAYER M2 ;
        RECT 6.56 25.448 6.592 25.48 ;
  LAYER M2 ;
        RECT 8.928 25.384 8.96 25.416 ;
  LAYER M2 ;
        RECT 6.56 25.32 6.592 25.352 ;
  LAYER M2 ;
        RECT 8.928 25.256 8.96 25.288 ;
  LAYER M2 ;
        RECT 6.56 25.192 6.592 25.224 ;
  LAYER M2 ;
        RECT 8.928 25.128 8.96 25.16 ;
  LAYER M2 ;
        RECT 6.56 25.064 6.592 25.096 ;
  LAYER M2 ;
        RECT 6.512 24.864 9.008 27.468 ;
  LAYER M1 ;
        RECT 8.928 21.804 8.96 24.312 ;
  LAYER M3 ;
        RECT 8.928 21.824 8.96 21.856 ;
  LAYER M1 ;
        RECT 8.864 21.804 8.896 24.312 ;
  LAYER M3 ;
        RECT 8.864 24.26 8.896 24.292 ;
  LAYER M1 ;
        RECT 8.8 21.804 8.832 24.312 ;
  LAYER M3 ;
        RECT 8.8 21.824 8.832 21.856 ;
  LAYER M1 ;
        RECT 8.736 21.804 8.768 24.312 ;
  LAYER M3 ;
        RECT 8.736 24.26 8.768 24.292 ;
  LAYER M1 ;
        RECT 8.672 21.804 8.704 24.312 ;
  LAYER M3 ;
        RECT 8.672 21.824 8.704 21.856 ;
  LAYER M1 ;
        RECT 8.608 21.804 8.64 24.312 ;
  LAYER M3 ;
        RECT 8.608 24.26 8.64 24.292 ;
  LAYER M1 ;
        RECT 8.544 21.804 8.576 24.312 ;
  LAYER M3 ;
        RECT 8.544 21.824 8.576 21.856 ;
  LAYER M1 ;
        RECT 8.48 21.804 8.512 24.312 ;
  LAYER M3 ;
        RECT 8.48 24.26 8.512 24.292 ;
  LAYER M1 ;
        RECT 8.416 21.804 8.448 24.312 ;
  LAYER M3 ;
        RECT 8.416 21.824 8.448 21.856 ;
  LAYER M1 ;
        RECT 8.352 21.804 8.384 24.312 ;
  LAYER M3 ;
        RECT 8.352 24.26 8.384 24.292 ;
  LAYER M1 ;
        RECT 8.288 21.804 8.32 24.312 ;
  LAYER M3 ;
        RECT 8.288 21.824 8.32 21.856 ;
  LAYER M1 ;
        RECT 8.224 21.804 8.256 24.312 ;
  LAYER M3 ;
        RECT 8.224 24.26 8.256 24.292 ;
  LAYER M1 ;
        RECT 8.16 21.804 8.192 24.312 ;
  LAYER M3 ;
        RECT 8.16 21.824 8.192 21.856 ;
  LAYER M1 ;
        RECT 8.096 21.804 8.128 24.312 ;
  LAYER M3 ;
        RECT 8.096 24.26 8.128 24.292 ;
  LAYER M1 ;
        RECT 8.032 21.804 8.064 24.312 ;
  LAYER M3 ;
        RECT 8.032 21.824 8.064 21.856 ;
  LAYER M1 ;
        RECT 7.968 21.804 8 24.312 ;
  LAYER M3 ;
        RECT 7.968 24.26 8 24.292 ;
  LAYER M1 ;
        RECT 7.904 21.804 7.936 24.312 ;
  LAYER M3 ;
        RECT 7.904 21.824 7.936 21.856 ;
  LAYER M1 ;
        RECT 7.84 21.804 7.872 24.312 ;
  LAYER M3 ;
        RECT 7.84 24.26 7.872 24.292 ;
  LAYER M1 ;
        RECT 7.776 21.804 7.808 24.312 ;
  LAYER M3 ;
        RECT 7.776 21.824 7.808 21.856 ;
  LAYER M1 ;
        RECT 7.712 21.804 7.744 24.312 ;
  LAYER M3 ;
        RECT 7.712 24.26 7.744 24.292 ;
  LAYER M1 ;
        RECT 7.648 21.804 7.68 24.312 ;
  LAYER M3 ;
        RECT 7.648 21.824 7.68 21.856 ;
  LAYER M1 ;
        RECT 7.584 21.804 7.616 24.312 ;
  LAYER M3 ;
        RECT 7.584 24.26 7.616 24.292 ;
  LAYER M1 ;
        RECT 7.52 21.804 7.552 24.312 ;
  LAYER M3 ;
        RECT 7.52 21.824 7.552 21.856 ;
  LAYER M1 ;
        RECT 7.456 21.804 7.488 24.312 ;
  LAYER M3 ;
        RECT 7.456 24.26 7.488 24.292 ;
  LAYER M1 ;
        RECT 7.392 21.804 7.424 24.312 ;
  LAYER M3 ;
        RECT 7.392 21.824 7.424 21.856 ;
  LAYER M1 ;
        RECT 7.328 21.804 7.36 24.312 ;
  LAYER M3 ;
        RECT 7.328 24.26 7.36 24.292 ;
  LAYER M1 ;
        RECT 7.264 21.804 7.296 24.312 ;
  LAYER M3 ;
        RECT 7.264 21.824 7.296 21.856 ;
  LAYER M1 ;
        RECT 7.2 21.804 7.232 24.312 ;
  LAYER M3 ;
        RECT 7.2 24.26 7.232 24.292 ;
  LAYER M1 ;
        RECT 7.136 21.804 7.168 24.312 ;
  LAYER M3 ;
        RECT 7.136 21.824 7.168 21.856 ;
  LAYER M1 ;
        RECT 7.072 21.804 7.104 24.312 ;
  LAYER M3 ;
        RECT 7.072 24.26 7.104 24.292 ;
  LAYER M1 ;
        RECT 7.008 21.804 7.04 24.312 ;
  LAYER M3 ;
        RECT 7.008 21.824 7.04 21.856 ;
  LAYER M1 ;
        RECT 6.944 21.804 6.976 24.312 ;
  LAYER M3 ;
        RECT 6.944 24.26 6.976 24.292 ;
  LAYER M1 ;
        RECT 6.88 21.804 6.912 24.312 ;
  LAYER M3 ;
        RECT 6.88 21.824 6.912 21.856 ;
  LAYER M1 ;
        RECT 6.816 21.804 6.848 24.312 ;
  LAYER M3 ;
        RECT 6.816 24.26 6.848 24.292 ;
  LAYER M1 ;
        RECT 6.752 21.804 6.784 24.312 ;
  LAYER M3 ;
        RECT 6.752 21.824 6.784 21.856 ;
  LAYER M1 ;
        RECT 6.688 21.804 6.72 24.312 ;
  LAYER M3 ;
        RECT 6.688 24.26 6.72 24.292 ;
  LAYER M1 ;
        RECT 6.624 21.804 6.656 24.312 ;
  LAYER M3 ;
        RECT 6.624 21.824 6.656 21.856 ;
  LAYER M1 ;
        RECT 6.56 21.804 6.592 24.312 ;
  LAYER M3 ;
        RECT 8.928 24.196 8.96 24.228 ;
  LAYER M2 ;
        RECT 6.56 24.132 6.592 24.164 ;
  LAYER M2 ;
        RECT 8.928 24.068 8.96 24.1 ;
  LAYER M2 ;
        RECT 6.56 24.004 6.592 24.036 ;
  LAYER M2 ;
        RECT 8.928 23.94 8.96 23.972 ;
  LAYER M2 ;
        RECT 6.56 23.876 6.592 23.908 ;
  LAYER M2 ;
        RECT 8.928 23.812 8.96 23.844 ;
  LAYER M2 ;
        RECT 6.56 23.748 6.592 23.78 ;
  LAYER M2 ;
        RECT 8.928 23.684 8.96 23.716 ;
  LAYER M2 ;
        RECT 6.56 23.62 6.592 23.652 ;
  LAYER M2 ;
        RECT 8.928 23.556 8.96 23.588 ;
  LAYER M2 ;
        RECT 6.56 23.492 6.592 23.524 ;
  LAYER M2 ;
        RECT 8.928 23.428 8.96 23.46 ;
  LAYER M2 ;
        RECT 6.56 23.364 6.592 23.396 ;
  LAYER M2 ;
        RECT 8.928 23.3 8.96 23.332 ;
  LAYER M2 ;
        RECT 6.56 23.236 6.592 23.268 ;
  LAYER M2 ;
        RECT 8.928 23.172 8.96 23.204 ;
  LAYER M2 ;
        RECT 6.56 23.108 6.592 23.14 ;
  LAYER M2 ;
        RECT 8.928 23.044 8.96 23.076 ;
  LAYER M2 ;
        RECT 6.56 22.98 6.592 23.012 ;
  LAYER M2 ;
        RECT 8.928 22.916 8.96 22.948 ;
  LAYER M2 ;
        RECT 6.56 22.852 6.592 22.884 ;
  LAYER M2 ;
        RECT 8.928 22.788 8.96 22.82 ;
  LAYER M2 ;
        RECT 6.56 22.724 6.592 22.756 ;
  LAYER M2 ;
        RECT 8.928 22.66 8.96 22.692 ;
  LAYER M2 ;
        RECT 6.56 22.596 6.592 22.628 ;
  LAYER M2 ;
        RECT 8.928 22.532 8.96 22.564 ;
  LAYER M2 ;
        RECT 6.56 22.468 6.592 22.5 ;
  LAYER M2 ;
        RECT 8.928 22.404 8.96 22.436 ;
  LAYER M2 ;
        RECT 6.56 22.34 6.592 22.372 ;
  LAYER M2 ;
        RECT 8.928 22.276 8.96 22.308 ;
  LAYER M2 ;
        RECT 6.56 22.212 6.592 22.244 ;
  LAYER M2 ;
        RECT 8.928 22.148 8.96 22.18 ;
  LAYER M2 ;
        RECT 6.56 22.084 6.592 22.116 ;
  LAYER M2 ;
        RECT 8.928 22.02 8.96 22.052 ;
  LAYER M2 ;
        RECT 6.56 21.956 6.592 21.988 ;
  LAYER M2 ;
        RECT 6.512 21.756 9.008 24.36 ;
  LAYER M1 ;
        RECT 8.928 18.696 8.96 21.204 ;
  LAYER M3 ;
        RECT 8.928 18.716 8.96 18.748 ;
  LAYER M1 ;
        RECT 8.864 18.696 8.896 21.204 ;
  LAYER M3 ;
        RECT 8.864 21.152 8.896 21.184 ;
  LAYER M1 ;
        RECT 8.8 18.696 8.832 21.204 ;
  LAYER M3 ;
        RECT 8.8 18.716 8.832 18.748 ;
  LAYER M1 ;
        RECT 8.736 18.696 8.768 21.204 ;
  LAYER M3 ;
        RECT 8.736 21.152 8.768 21.184 ;
  LAYER M1 ;
        RECT 8.672 18.696 8.704 21.204 ;
  LAYER M3 ;
        RECT 8.672 18.716 8.704 18.748 ;
  LAYER M1 ;
        RECT 8.608 18.696 8.64 21.204 ;
  LAYER M3 ;
        RECT 8.608 21.152 8.64 21.184 ;
  LAYER M1 ;
        RECT 8.544 18.696 8.576 21.204 ;
  LAYER M3 ;
        RECT 8.544 18.716 8.576 18.748 ;
  LAYER M1 ;
        RECT 8.48 18.696 8.512 21.204 ;
  LAYER M3 ;
        RECT 8.48 21.152 8.512 21.184 ;
  LAYER M1 ;
        RECT 8.416 18.696 8.448 21.204 ;
  LAYER M3 ;
        RECT 8.416 18.716 8.448 18.748 ;
  LAYER M1 ;
        RECT 8.352 18.696 8.384 21.204 ;
  LAYER M3 ;
        RECT 8.352 21.152 8.384 21.184 ;
  LAYER M1 ;
        RECT 8.288 18.696 8.32 21.204 ;
  LAYER M3 ;
        RECT 8.288 18.716 8.32 18.748 ;
  LAYER M1 ;
        RECT 8.224 18.696 8.256 21.204 ;
  LAYER M3 ;
        RECT 8.224 21.152 8.256 21.184 ;
  LAYER M1 ;
        RECT 8.16 18.696 8.192 21.204 ;
  LAYER M3 ;
        RECT 8.16 18.716 8.192 18.748 ;
  LAYER M1 ;
        RECT 8.096 18.696 8.128 21.204 ;
  LAYER M3 ;
        RECT 8.096 21.152 8.128 21.184 ;
  LAYER M1 ;
        RECT 8.032 18.696 8.064 21.204 ;
  LAYER M3 ;
        RECT 8.032 18.716 8.064 18.748 ;
  LAYER M1 ;
        RECT 7.968 18.696 8 21.204 ;
  LAYER M3 ;
        RECT 7.968 21.152 8 21.184 ;
  LAYER M1 ;
        RECT 7.904 18.696 7.936 21.204 ;
  LAYER M3 ;
        RECT 7.904 18.716 7.936 18.748 ;
  LAYER M1 ;
        RECT 7.84 18.696 7.872 21.204 ;
  LAYER M3 ;
        RECT 7.84 21.152 7.872 21.184 ;
  LAYER M1 ;
        RECT 7.776 18.696 7.808 21.204 ;
  LAYER M3 ;
        RECT 7.776 18.716 7.808 18.748 ;
  LAYER M1 ;
        RECT 7.712 18.696 7.744 21.204 ;
  LAYER M3 ;
        RECT 7.712 21.152 7.744 21.184 ;
  LAYER M1 ;
        RECT 7.648 18.696 7.68 21.204 ;
  LAYER M3 ;
        RECT 7.648 18.716 7.68 18.748 ;
  LAYER M1 ;
        RECT 7.584 18.696 7.616 21.204 ;
  LAYER M3 ;
        RECT 7.584 21.152 7.616 21.184 ;
  LAYER M1 ;
        RECT 7.52 18.696 7.552 21.204 ;
  LAYER M3 ;
        RECT 7.52 18.716 7.552 18.748 ;
  LAYER M1 ;
        RECT 7.456 18.696 7.488 21.204 ;
  LAYER M3 ;
        RECT 7.456 21.152 7.488 21.184 ;
  LAYER M1 ;
        RECT 7.392 18.696 7.424 21.204 ;
  LAYER M3 ;
        RECT 7.392 18.716 7.424 18.748 ;
  LAYER M1 ;
        RECT 7.328 18.696 7.36 21.204 ;
  LAYER M3 ;
        RECT 7.328 21.152 7.36 21.184 ;
  LAYER M1 ;
        RECT 7.264 18.696 7.296 21.204 ;
  LAYER M3 ;
        RECT 7.264 18.716 7.296 18.748 ;
  LAYER M1 ;
        RECT 7.2 18.696 7.232 21.204 ;
  LAYER M3 ;
        RECT 7.2 21.152 7.232 21.184 ;
  LAYER M1 ;
        RECT 7.136 18.696 7.168 21.204 ;
  LAYER M3 ;
        RECT 7.136 18.716 7.168 18.748 ;
  LAYER M1 ;
        RECT 7.072 18.696 7.104 21.204 ;
  LAYER M3 ;
        RECT 7.072 21.152 7.104 21.184 ;
  LAYER M1 ;
        RECT 7.008 18.696 7.04 21.204 ;
  LAYER M3 ;
        RECT 7.008 18.716 7.04 18.748 ;
  LAYER M1 ;
        RECT 6.944 18.696 6.976 21.204 ;
  LAYER M3 ;
        RECT 6.944 21.152 6.976 21.184 ;
  LAYER M1 ;
        RECT 6.88 18.696 6.912 21.204 ;
  LAYER M3 ;
        RECT 6.88 18.716 6.912 18.748 ;
  LAYER M1 ;
        RECT 6.816 18.696 6.848 21.204 ;
  LAYER M3 ;
        RECT 6.816 21.152 6.848 21.184 ;
  LAYER M1 ;
        RECT 6.752 18.696 6.784 21.204 ;
  LAYER M3 ;
        RECT 6.752 18.716 6.784 18.748 ;
  LAYER M1 ;
        RECT 6.688 18.696 6.72 21.204 ;
  LAYER M3 ;
        RECT 6.688 21.152 6.72 21.184 ;
  LAYER M1 ;
        RECT 6.624 18.696 6.656 21.204 ;
  LAYER M3 ;
        RECT 6.624 18.716 6.656 18.748 ;
  LAYER M1 ;
        RECT 6.56 18.696 6.592 21.204 ;
  LAYER M3 ;
        RECT 8.928 21.088 8.96 21.12 ;
  LAYER M2 ;
        RECT 6.56 21.024 6.592 21.056 ;
  LAYER M2 ;
        RECT 8.928 20.96 8.96 20.992 ;
  LAYER M2 ;
        RECT 6.56 20.896 6.592 20.928 ;
  LAYER M2 ;
        RECT 8.928 20.832 8.96 20.864 ;
  LAYER M2 ;
        RECT 6.56 20.768 6.592 20.8 ;
  LAYER M2 ;
        RECT 8.928 20.704 8.96 20.736 ;
  LAYER M2 ;
        RECT 6.56 20.64 6.592 20.672 ;
  LAYER M2 ;
        RECT 8.928 20.576 8.96 20.608 ;
  LAYER M2 ;
        RECT 6.56 20.512 6.592 20.544 ;
  LAYER M2 ;
        RECT 8.928 20.448 8.96 20.48 ;
  LAYER M2 ;
        RECT 6.56 20.384 6.592 20.416 ;
  LAYER M2 ;
        RECT 8.928 20.32 8.96 20.352 ;
  LAYER M2 ;
        RECT 6.56 20.256 6.592 20.288 ;
  LAYER M2 ;
        RECT 8.928 20.192 8.96 20.224 ;
  LAYER M2 ;
        RECT 6.56 20.128 6.592 20.16 ;
  LAYER M2 ;
        RECT 8.928 20.064 8.96 20.096 ;
  LAYER M2 ;
        RECT 6.56 20 6.592 20.032 ;
  LAYER M2 ;
        RECT 8.928 19.936 8.96 19.968 ;
  LAYER M2 ;
        RECT 6.56 19.872 6.592 19.904 ;
  LAYER M2 ;
        RECT 8.928 19.808 8.96 19.84 ;
  LAYER M2 ;
        RECT 6.56 19.744 6.592 19.776 ;
  LAYER M2 ;
        RECT 8.928 19.68 8.96 19.712 ;
  LAYER M2 ;
        RECT 6.56 19.616 6.592 19.648 ;
  LAYER M2 ;
        RECT 8.928 19.552 8.96 19.584 ;
  LAYER M2 ;
        RECT 6.56 19.488 6.592 19.52 ;
  LAYER M2 ;
        RECT 8.928 19.424 8.96 19.456 ;
  LAYER M2 ;
        RECT 6.56 19.36 6.592 19.392 ;
  LAYER M2 ;
        RECT 8.928 19.296 8.96 19.328 ;
  LAYER M2 ;
        RECT 6.56 19.232 6.592 19.264 ;
  LAYER M2 ;
        RECT 8.928 19.168 8.96 19.2 ;
  LAYER M2 ;
        RECT 6.56 19.104 6.592 19.136 ;
  LAYER M2 ;
        RECT 8.928 19.04 8.96 19.072 ;
  LAYER M2 ;
        RECT 6.56 18.976 6.592 19.008 ;
  LAYER M2 ;
        RECT 8.928 18.912 8.96 18.944 ;
  LAYER M2 ;
        RECT 6.56 18.848 6.592 18.88 ;
  LAYER M2 ;
        RECT 6.512 18.648 9.008 21.252 ;
  LAYER M1 ;
        RECT 8.928 15.588 8.96 18.096 ;
  LAYER M3 ;
        RECT 8.928 15.608 8.96 15.64 ;
  LAYER M1 ;
        RECT 8.864 15.588 8.896 18.096 ;
  LAYER M3 ;
        RECT 8.864 18.044 8.896 18.076 ;
  LAYER M1 ;
        RECT 8.8 15.588 8.832 18.096 ;
  LAYER M3 ;
        RECT 8.8 15.608 8.832 15.64 ;
  LAYER M1 ;
        RECT 8.736 15.588 8.768 18.096 ;
  LAYER M3 ;
        RECT 8.736 18.044 8.768 18.076 ;
  LAYER M1 ;
        RECT 8.672 15.588 8.704 18.096 ;
  LAYER M3 ;
        RECT 8.672 15.608 8.704 15.64 ;
  LAYER M1 ;
        RECT 8.608 15.588 8.64 18.096 ;
  LAYER M3 ;
        RECT 8.608 18.044 8.64 18.076 ;
  LAYER M1 ;
        RECT 8.544 15.588 8.576 18.096 ;
  LAYER M3 ;
        RECT 8.544 15.608 8.576 15.64 ;
  LAYER M1 ;
        RECT 8.48 15.588 8.512 18.096 ;
  LAYER M3 ;
        RECT 8.48 18.044 8.512 18.076 ;
  LAYER M1 ;
        RECT 8.416 15.588 8.448 18.096 ;
  LAYER M3 ;
        RECT 8.416 15.608 8.448 15.64 ;
  LAYER M1 ;
        RECT 8.352 15.588 8.384 18.096 ;
  LAYER M3 ;
        RECT 8.352 18.044 8.384 18.076 ;
  LAYER M1 ;
        RECT 8.288 15.588 8.32 18.096 ;
  LAYER M3 ;
        RECT 8.288 15.608 8.32 15.64 ;
  LAYER M1 ;
        RECT 8.224 15.588 8.256 18.096 ;
  LAYER M3 ;
        RECT 8.224 18.044 8.256 18.076 ;
  LAYER M1 ;
        RECT 8.16 15.588 8.192 18.096 ;
  LAYER M3 ;
        RECT 8.16 15.608 8.192 15.64 ;
  LAYER M1 ;
        RECT 8.096 15.588 8.128 18.096 ;
  LAYER M3 ;
        RECT 8.096 18.044 8.128 18.076 ;
  LAYER M1 ;
        RECT 8.032 15.588 8.064 18.096 ;
  LAYER M3 ;
        RECT 8.032 15.608 8.064 15.64 ;
  LAYER M1 ;
        RECT 7.968 15.588 8 18.096 ;
  LAYER M3 ;
        RECT 7.968 18.044 8 18.076 ;
  LAYER M1 ;
        RECT 7.904 15.588 7.936 18.096 ;
  LAYER M3 ;
        RECT 7.904 15.608 7.936 15.64 ;
  LAYER M1 ;
        RECT 7.84 15.588 7.872 18.096 ;
  LAYER M3 ;
        RECT 7.84 18.044 7.872 18.076 ;
  LAYER M1 ;
        RECT 7.776 15.588 7.808 18.096 ;
  LAYER M3 ;
        RECT 7.776 15.608 7.808 15.64 ;
  LAYER M1 ;
        RECT 7.712 15.588 7.744 18.096 ;
  LAYER M3 ;
        RECT 7.712 18.044 7.744 18.076 ;
  LAYER M1 ;
        RECT 7.648 15.588 7.68 18.096 ;
  LAYER M3 ;
        RECT 7.648 15.608 7.68 15.64 ;
  LAYER M1 ;
        RECT 7.584 15.588 7.616 18.096 ;
  LAYER M3 ;
        RECT 7.584 18.044 7.616 18.076 ;
  LAYER M1 ;
        RECT 7.52 15.588 7.552 18.096 ;
  LAYER M3 ;
        RECT 7.52 15.608 7.552 15.64 ;
  LAYER M1 ;
        RECT 7.456 15.588 7.488 18.096 ;
  LAYER M3 ;
        RECT 7.456 18.044 7.488 18.076 ;
  LAYER M1 ;
        RECT 7.392 15.588 7.424 18.096 ;
  LAYER M3 ;
        RECT 7.392 15.608 7.424 15.64 ;
  LAYER M1 ;
        RECT 7.328 15.588 7.36 18.096 ;
  LAYER M3 ;
        RECT 7.328 18.044 7.36 18.076 ;
  LAYER M1 ;
        RECT 7.264 15.588 7.296 18.096 ;
  LAYER M3 ;
        RECT 7.264 15.608 7.296 15.64 ;
  LAYER M1 ;
        RECT 7.2 15.588 7.232 18.096 ;
  LAYER M3 ;
        RECT 7.2 18.044 7.232 18.076 ;
  LAYER M1 ;
        RECT 7.136 15.588 7.168 18.096 ;
  LAYER M3 ;
        RECT 7.136 15.608 7.168 15.64 ;
  LAYER M1 ;
        RECT 7.072 15.588 7.104 18.096 ;
  LAYER M3 ;
        RECT 7.072 18.044 7.104 18.076 ;
  LAYER M1 ;
        RECT 7.008 15.588 7.04 18.096 ;
  LAYER M3 ;
        RECT 7.008 15.608 7.04 15.64 ;
  LAYER M1 ;
        RECT 6.944 15.588 6.976 18.096 ;
  LAYER M3 ;
        RECT 6.944 18.044 6.976 18.076 ;
  LAYER M1 ;
        RECT 6.88 15.588 6.912 18.096 ;
  LAYER M3 ;
        RECT 6.88 15.608 6.912 15.64 ;
  LAYER M1 ;
        RECT 6.816 15.588 6.848 18.096 ;
  LAYER M3 ;
        RECT 6.816 18.044 6.848 18.076 ;
  LAYER M1 ;
        RECT 6.752 15.588 6.784 18.096 ;
  LAYER M3 ;
        RECT 6.752 15.608 6.784 15.64 ;
  LAYER M1 ;
        RECT 6.688 15.588 6.72 18.096 ;
  LAYER M3 ;
        RECT 6.688 18.044 6.72 18.076 ;
  LAYER M1 ;
        RECT 6.624 15.588 6.656 18.096 ;
  LAYER M3 ;
        RECT 6.624 15.608 6.656 15.64 ;
  LAYER M1 ;
        RECT 6.56 15.588 6.592 18.096 ;
  LAYER M3 ;
        RECT 8.928 17.98 8.96 18.012 ;
  LAYER M2 ;
        RECT 6.56 17.916 6.592 17.948 ;
  LAYER M2 ;
        RECT 8.928 17.852 8.96 17.884 ;
  LAYER M2 ;
        RECT 6.56 17.788 6.592 17.82 ;
  LAYER M2 ;
        RECT 8.928 17.724 8.96 17.756 ;
  LAYER M2 ;
        RECT 6.56 17.66 6.592 17.692 ;
  LAYER M2 ;
        RECT 8.928 17.596 8.96 17.628 ;
  LAYER M2 ;
        RECT 6.56 17.532 6.592 17.564 ;
  LAYER M2 ;
        RECT 8.928 17.468 8.96 17.5 ;
  LAYER M2 ;
        RECT 6.56 17.404 6.592 17.436 ;
  LAYER M2 ;
        RECT 8.928 17.34 8.96 17.372 ;
  LAYER M2 ;
        RECT 6.56 17.276 6.592 17.308 ;
  LAYER M2 ;
        RECT 8.928 17.212 8.96 17.244 ;
  LAYER M2 ;
        RECT 6.56 17.148 6.592 17.18 ;
  LAYER M2 ;
        RECT 8.928 17.084 8.96 17.116 ;
  LAYER M2 ;
        RECT 6.56 17.02 6.592 17.052 ;
  LAYER M2 ;
        RECT 8.928 16.956 8.96 16.988 ;
  LAYER M2 ;
        RECT 6.56 16.892 6.592 16.924 ;
  LAYER M2 ;
        RECT 8.928 16.828 8.96 16.86 ;
  LAYER M2 ;
        RECT 6.56 16.764 6.592 16.796 ;
  LAYER M2 ;
        RECT 8.928 16.7 8.96 16.732 ;
  LAYER M2 ;
        RECT 6.56 16.636 6.592 16.668 ;
  LAYER M2 ;
        RECT 8.928 16.572 8.96 16.604 ;
  LAYER M2 ;
        RECT 6.56 16.508 6.592 16.54 ;
  LAYER M2 ;
        RECT 8.928 16.444 8.96 16.476 ;
  LAYER M2 ;
        RECT 6.56 16.38 6.592 16.412 ;
  LAYER M2 ;
        RECT 8.928 16.316 8.96 16.348 ;
  LAYER M2 ;
        RECT 6.56 16.252 6.592 16.284 ;
  LAYER M2 ;
        RECT 8.928 16.188 8.96 16.22 ;
  LAYER M2 ;
        RECT 6.56 16.124 6.592 16.156 ;
  LAYER M2 ;
        RECT 8.928 16.06 8.96 16.092 ;
  LAYER M2 ;
        RECT 6.56 15.996 6.592 16.028 ;
  LAYER M2 ;
        RECT 8.928 15.932 8.96 15.964 ;
  LAYER M2 ;
        RECT 6.56 15.868 6.592 15.9 ;
  LAYER M2 ;
        RECT 8.928 15.804 8.96 15.836 ;
  LAYER M2 ;
        RECT 6.56 15.74 6.592 15.772 ;
  LAYER M2 ;
        RECT 6.512 15.54 9.008 18.144 ;
  LAYER M1 ;
        RECT 5.952 28.02 5.984 30.528 ;
  LAYER M3 ;
        RECT 5.952 28.04 5.984 28.072 ;
  LAYER M1 ;
        RECT 5.888 28.02 5.92 30.528 ;
  LAYER M3 ;
        RECT 5.888 30.476 5.92 30.508 ;
  LAYER M1 ;
        RECT 5.824 28.02 5.856 30.528 ;
  LAYER M3 ;
        RECT 5.824 28.04 5.856 28.072 ;
  LAYER M1 ;
        RECT 5.76 28.02 5.792 30.528 ;
  LAYER M3 ;
        RECT 5.76 30.476 5.792 30.508 ;
  LAYER M1 ;
        RECT 5.696 28.02 5.728 30.528 ;
  LAYER M3 ;
        RECT 5.696 28.04 5.728 28.072 ;
  LAYER M1 ;
        RECT 5.632 28.02 5.664 30.528 ;
  LAYER M3 ;
        RECT 5.632 30.476 5.664 30.508 ;
  LAYER M1 ;
        RECT 5.568 28.02 5.6 30.528 ;
  LAYER M3 ;
        RECT 5.568 28.04 5.6 28.072 ;
  LAYER M1 ;
        RECT 5.504 28.02 5.536 30.528 ;
  LAYER M3 ;
        RECT 5.504 30.476 5.536 30.508 ;
  LAYER M1 ;
        RECT 5.44 28.02 5.472 30.528 ;
  LAYER M3 ;
        RECT 5.44 28.04 5.472 28.072 ;
  LAYER M1 ;
        RECT 5.376 28.02 5.408 30.528 ;
  LAYER M3 ;
        RECT 5.376 30.476 5.408 30.508 ;
  LAYER M1 ;
        RECT 5.312 28.02 5.344 30.528 ;
  LAYER M3 ;
        RECT 5.312 28.04 5.344 28.072 ;
  LAYER M1 ;
        RECT 5.248 28.02 5.28 30.528 ;
  LAYER M3 ;
        RECT 5.248 30.476 5.28 30.508 ;
  LAYER M1 ;
        RECT 5.184 28.02 5.216 30.528 ;
  LAYER M3 ;
        RECT 5.184 28.04 5.216 28.072 ;
  LAYER M1 ;
        RECT 5.12 28.02 5.152 30.528 ;
  LAYER M3 ;
        RECT 5.12 30.476 5.152 30.508 ;
  LAYER M1 ;
        RECT 5.056 28.02 5.088 30.528 ;
  LAYER M3 ;
        RECT 5.056 28.04 5.088 28.072 ;
  LAYER M1 ;
        RECT 4.992 28.02 5.024 30.528 ;
  LAYER M3 ;
        RECT 4.992 30.476 5.024 30.508 ;
  LAYER M1 ;
        RECT 4.928 28.02 4.96 30.528 ;
  LAYER M3 ;
        RECT 4.928 28.04 4.96 28.072 ;
  LAYER M1 ;
        RECT 4.864 28.02 4.896 30.528 ;
  LAYER M3 ;
        RECT 4.864 30.476 4.896 30.508 ;
  LAYER M1 ;
        RECT 4.8 28.02 4.832 30.528 ;
  LAYER M3 ;
        RECT 4.8 28.04 4.832 28.072 ;
  LAYER M1 ;
        RECT 4.736 28.02 4.768 30.528 ;
  LAYER M3 ;
        RECT 4.736 30.476 4.768 30.508 ;
  LAYER M1 ;
        RECT 4.672 28.02 4.704 30.528 ;
  LAYER M3 ;
        RECT 4.672 28.04 4.704 28.072 ;
  LAYER M1 ;
        RECT 4.608 28.02 4.64 30.528 ;
  LAYER M3 ;
        RECT 4.608 30.476 4.64 30.508 ;
  LAYER M1 ;
        RECT 4.544 28.02 4.576 30.528 ;
  LAYER M3 ;
        RECT 4.544 28.04 4.576 28.072 ;
  LAYER M1 ;
        RECT 4.48 28.02 4.512 30.528 ;
  LAYER M3 ;
        RECT 4.48 30.476 4.512 30.508 ;
  LAYER M1 ;
        RECT 4.416 28.02 4.448 30.528 ;
  LAYER M3 ;
        RECT 4.416 28.04 4.448 28.072 ;
  LAYER M1 ;
        RECT 4.352 28.02 4.384 30.528 ;
  LAYER M3 ;
        RECT 4.352 30.476 4.384 30.508 ;
  LAYER M1 ;
        RECT 4.288 28.02 4.32 30.528 ;
  LAYER M3 ;
        RECT 4.288 28.04 4.32 28.072 ;
  LAYER M1 ;
        RECT 4.224 28.02 4.256 30.528 ;
  LAYER M3 ;
        RECT 4.224 30.476 4.256 30.508 ;
  LAYER M1 ;
        RECT 4.16 28.02 4.192 30.528 ;
  LAYER M3 ;
        RECT 4.16 28.04 4.192 28.072 ;
  LAYER M1 ;
        RECT 4.096 28.02 4.128 30.528 ;
  LAYER M3 ;
        RECT 4.096 30.476 4.128 30.508 ;
  LAYER M1 ;
        RECT 4.032 28.02 4.064 30.528 ;
  LAYER M3 ;
        RECT 4.032 28.04 4.064 28.072 ;
  LAYER M1 ;
        RECT 3.968 28.02 4 30.528 ;
  LAYER M3 ;
        RECT 3.968 30.476 4 30.508 ;
  LAYER M1 ;
        RECT 3.904 28.02 3.936 30.528 ;
  LAYER M3 ;
        RECT 3.904 28.04 3.936 28.072 ;
  LAYER M1 ;
        RECT 3.84 28.02 3.872 30.528 ;
  LAYER M3 ;
        RECT 3.84 30.476 3.872 30.508 ;
  LAYER M1 ;
        RECT 3.776 28.02 3.808 30.528 ;
  LAYER M3 ;
        RECT 3.776 28.04 3.808 28.072 ;
  LAYER M1 ;
        RECT 3.712 28.02 3.744 30.528 ;
  LAYER M3 ;
        RECT 3.712 30.476 3.744 30.508 ;
  LAYER M1 ;
        RECT 3.648 28.02 3.68 30.528 ;
  LAYER M3 ;
        RECT 3.648 28.04 3.68 28.072 ;
  LAYER M1 ;
        RECT 3.584 28.02 3.616 30.528 ;
  LAYER M3 ;
        RECT 5.952 30.412 5.984 30.444 ;
  LAYER M2 ;
        RECT 3.584 30.348 3.616 30.38 ;
  LAYER M2 ;
        RECT 5.952 30.284 5.984 30.316 ;
  LAYER M2 ;
        RECT 3.584 30.22 3.616 30.252 ;
  LAYER M2 ;
        RECT 5.952 30.156 5.984 30.188 ;
  LAYER M2 ;
        RECT 3.584 30.092 3.616 30.124 ;
  LAYER M2 ;
        RECT 5.952 30.028 5.984 30.06 ;
  LAYER M2 ;
        RECT 3.584 29.964 3.616 29.996 ;
  LAYER M2 ;
        RECT 5.952 29.9 5.984 29.932 ;
  LAYER M2 ;
        RECT 3.584 29.836 3.616 29.868 ;
  LAYER M2 ;
        RECT 5.952 29.772 5.984 29.804 ;
  LAYER M2 ;
        RECT 3.584 29.708 3.616 29.74 ;
  LAYER M2 ;
        RECT 5.952 29.644 5.984 29.676 ;
  LAYER M2 ;
        RECT 3.584 29.58 3.616 29.612 ;
  LAYER M2 ;
        RECT 5.952 29.516 5.984 29.548 ;
  LAYER M2 ;
        RECT 3.584 29.452 3.616 29.484 ;
  LAYER M2 ;
        RECT 5.952 29.388 5.984 29.42 ;
  LAYER M2 ;
        RECT 3.584 29.324 3.616 29.356 ;
  LAYER M2 ;
        RECT 5.952 29.26 5.984 29.292 ;
  LAYER M2 ;
        RECT 3.584 29.196 3.616 29.228 ;
  LAYER M2 ;
        RECT 5.952 29.132 5.984 29.164 ;
  LAYER M2 ;
        RECT 3.584 29.068 3.616 29.1 ;
  LAYER M2 ;
        RECT 5.952 29.004 5.984 29.036 ;
  LAYER M2 ;
        RECT 3.584 28.94 3.616 28.972 ;
  LAYER M2 ;
        RECT 5.952 28.876 5.984 28.908 ;
  LAYER M2 ;
        RECT 3.584 28.812 3.616 28.844 ;
  LAYER M2 ;
        RECT 5.952 28.748 5.984 28.78 ;
  LAYER M2 ;
        RECT 3.584 28.684 3.616 28.716 ;
  LAYER M2 ;
        RECT 5.952 28.62 5.984 28.652 ;
  LAYER M2 ;
        RECT 3.584 28.556 3.616 28.588 ;
  LAYER M2 ;
        RECT 5.952 28.492 5.984 28.524 ;
  LAYER M2 ;
        RECT 3.584 28.428 3.616 28.46 ;
  LAYER M2 ;
        RECT 5.952 28.364 5.984 28.396 ;
  LAYER M2 ;
        RECT 3.584 28.3 3.616 28.332 ;
  LAYER M2 ;
        RECT 5.952 28.236 5.984 28.268 ;
  LAYER M2 ;
        RECT 3.584 28.172 3.616 28.204 ;
  LAYER M2 ;
        RECT 3.536 27.972 6.032 30.576 ;
  LAYER M1 ;
        RECT 5.952 24.912 5.984 27.42 ;
  LAYER M3 ;
        RECT 5.952 24.932 5.984 24.964 ;
  LAYER M1 ;
        RECT 5.888 24.912 5.92 27.42 ;
  LAYER M3 ;
        RECT 5.888 27.368 5.92 27.4 ;
  LAYER M1 ;
        RECT 5.824 24.912 5.856 27.42 ;
  LAYER M3 ;
        RECT 5.824 24.932 5.856 24.964 ;
  LAYER M1 ;
        RECT 5.76 24.912 5.792 27.42 ;
  LAYER M3 ;
        RECT 5.76 27.368 5.792 27.4 ;
  LAYER M1 ;
        RECT 5.696 24.912 5.728 27.42 ;
  LAYER M3 ;
        RECT 5.696 24.932 5.728 24.964 ;
  LAYER M1 ;
        RECT 5.632 24.912 5.664 27.42 ;
  LAYER M3 ;
        RECT 5.632 27.368 5.664 27.4 ;
  LAYER M1 ;
        RECT 5.568 24.912 5.6 27.42 ;
  LAYER M3 ;
        RECT 5.568 24.932 5.6 24.964 ;
  LAYER M1 ;
        RECT 5.504 24.912 5.536 27.42 ;
  LAYER M3 ;
        RECT 5.504 27.368 5.536 27.4 ;
  LAYER M1 ;
        RECT 5.44 24.912 5.472 27.42 ;
  LAYER M3 ;
        RECT 5.44 24.932 5.472 24.964 ;
  LAYER M1 ;
        RECT 5.376 24.912 5.408 27.42 ;
  LAYER M3 ;
        RECT 5.376 27.368 5.408 27.4 ;
  LAYER M1 ;
        RECT 5.312 24.912 5.344 27.42 ;
  LAYER M3 ;
        RECT 5.312 24.932 5.344 24.964 ;
  LAYER M1 ;
        RECT 5.248 24.912 5.28 27.42 ;
  LAYER M3 ;
        RECT 5.248 27.368 5.28 27.4 ;
  LAYER M1 ;
        RECT 5.184 24.912 5.216 27.42 ;
  LAYER M3 ;
        RECT 5.184 24.932 5.216 24.964 ;
  LAYER M1 ;
        RECT 5.12 24.912 5.152 27.42 ;
  LAYER M3 ;
        RECT 5.12 27.368 5.152 27.4 ;
  LAYER M1 ;
        RECT 5.056 24.912 5.088 27.42 ;
  LAYER M3 ;
        RECT 5.056 24.932 5.088 24.964 ;
  LAYER M1 ;
        RECT 4.992 24.912 5.024 27.42 ;
  LAYER M3 ;
        RECT 4.992 27.368 5.024 27.4 ;
  LAYER M1 ;
        RECT 4.928 24.912 4.96 27.42 ;
  LAYER M3 ;
        RECT 4.928 24.932 4.96 24.964 ;
  LAYER M1 ;
        RECT 4.864 24.912 4.896 27.42 ;
  LAYER M3 ;
        RECT 4.864 27.368 4.896 27.4 ;
  LAYER M1 ;
        RECT 4.8 24.912 4.832 27.42 ;
  LAYER M3 ;
        RECT 4.8 24.932 4.832 24.964 ;
  LAYER M1 ;
        RECT 4.736 24.912 4.768 27.42 ;
  LAYER M3 ;
        RECT 4.736 27.368 4.768 27.4 ;
  LAYER M1 ;
        RECT 4.672 24.912 4.704 27.42 ;
  LAYER M3 ;
        RECT 4.672 24.932 4.704 24.964 ;
  LAYER M1 ;
        RECT 4.608 24.912 4.64 27.42 ;
  LAYER M3 ;
        RECT 4.608 27.368 4.64 27.4 ;
  LAYER M1 ;
        RECT 4.544 24.912 4.576 27.42 ;
  LAYER M3 ;
        RECT 4.544 24.932 4.576 24.964 ;
  LAYER M1 ;
        RECT 4.48 24.912 4.512 27.42 ;
  LAYER M3 ;
        RECT 4.48 27.368 4.512 27.4 ;
  LAYER M1 ;
        RECT 4.416 24.912 4.448 27.42 ;
  LAYER M3 ;
        RECT 4.416 24.932 4.448 24.964 ;
  LAYER M1 ;
        RECT 4.352 24.912 4.384 27.42 ;
  LAYER M3 ;
        RECT 4.352 27.368 4.384 27.4 ;
  LAYER M1 ;
        RECT 4.288 24.912 4.32 27.42 ;
  LAYER M3 ;
        RECT 4.288 24.932 4.32 24.964 ;
  LAYER M1 ;
        RECT 4.224 24.912 4.256 27.42 ;
  LAYER M3 ;
        RECT 4.224 27.368 4.256 27.4 ;
  LAYER M1 ;
        RECT 4.16 24.912 4.192 27.42 ;
  LAYER M3 ;
        RECT 4.16 24.932 4.192 24.964 ;
  LAYER M1 ;
        RECT 4.096 24.912 4.128 27.42 ;
  LAYER M3 ;
        RECT 4.096 27.368 4.128 27.4 ;
  LAYER M1 ;
        RECT 4.032 24.912 4.064 27.42 ;
  LAYER M3 ;
        RECT 4.032 24.932 4.064 24.964 ;
  LAYER M1 ;
        RECT 3.968 24.912 4 27.42 ;
  LAYER M3 ;
        RECT 3.968 27.368 4 27.4 ;
  LAYER M1 ;
        RECT 3.904 24.912 3.936 27.42 ;
  LAYER M3 ;
        RECT 3.904 24.932 3.936 24.964 ;
  LAYER M1 ;
        RECT 3.84 24.912 3.872 27.42 ;
  LAYER M3 ;
        RECT 3.84 27.368 3.872 27.4 ;
  LAYER M1 ;
        RECT 3.776 24.912 3.808 27.42 ;
  LAYER M3 ;
        RECT 3.776 24.932 3.808 24.964 ;
  LAYER M1 ;
        RECT 3.712 24.912 3.744 27.42 ;
  LAYER M3 ;
        RECT 3.712 27.368 3.744 27.4 ;
  LAYER M1 ;
        RECT 3.648 24.912 3.68 27.42 ;
  LAYER M3 ;
        RECT 3.648 24.932 3.68 24.964 ;
  LAYER M1 ;
        RECT 3.584 24.912 3.616 27.42 ;
  LAYER M3 ;
        RECT 5.952 27.304 5.984 27.336 ;
  LAYER M2 ;
        RECT 3.584 27.24 3.616 27.272 ;
  LAYER M2 ;
        RECT 5.952 27.176 5.984 27.208 ;
  LAYER M2 ;
        RECT 3.584 27.112 3.616 27.144 ;
  LAYER M2 ;
        RECT 5.952 27.048 5.984 27.08 ;
  LAYER M2 ;
        RECT 3.584 26.984 3.616 27.016 ;
  LAYER M2 ;
        RECT 5.952 26.92 5.984 26.952 ;
  LAYER M2 ;
        RECT 3.584 26.856 3.616 26.888 ;
  LAYER M2 ;
        RECT 5.952 26.792 5.984 26.824 ;
  LAYER M2 ;
        RECT 3.584 26.728 3.616 26.76 ;
  LAYER M2 ;
        RECT 5.952 26.664 5.984 26.696 ;
  LAYER M2 ;
        RECT 3.584 26.6 3.616 26.632 ;
  LAYER M2 ;
        RECT 5.952 26.536 5.984 26.568 ;
  LAYER M2 ;
        RECT 3.584 26.472 3.616 26.504 ;
  LAYER M2 ;
        RECT 5.952 26.408 5.984 26.44 ;
  LAYER M2 ;
        RECT 3.584 26.344 3.616 26.376 ;
  LAYER M2 ;
        RECT 5.952 26.28 5.984 26.312 ;
  LAYER M2 ;
        RECT 3.584 26.216 3.616 26.248 ;
  LAYER M2 ;
        RECT 5.952 26.152 5.984 26.184 ;
  LAYER M2 ;
        RECT 3.584 26.088 3.616 26.12 ;
  LAYER M2 ;
        RECT 5.952 26.024 5.984 26.056 ;
  LAYER M2 ;
        RECT 3.584 25.96 3.616 25.992 ;
  LAYER M2 ;
        RECT 5.952 25.896 5.984 25.928 ;
  LAYER M2 ;
        RECT 3.584 25.832 3.616 25.864 ;
  LAYER M2 ;
        RECT 5.952 25.768 5.984 25.8 ;
  LAYER M2 ;
        RECT 3.584 25.704 3.616 25.736 ;
  LAYER M2 ;
        RECT 5.952 25.64 5.984 25.672 ;
  LAYER M2 ;
        RECT 3.584 25.576 3.616 25.608 ;
  LAYER M2 ;
        RECT 5.952 25.512 5.984 25.544 ;
  LAYER M2 ;
        RECT 3.584 25.448 3.616 25.48 ;
  LAYER M2 ;
        RECT 5.952 25.384 5.984 25.416 ;
  LAYER M2 ;
        RECT 3.584 25.32 3.616 25.352 ;
  LAYER M2 ;
        RECT 5.952 25.256 5.984 25.288 ;
  LAYER M2 ;
        RECT 3.584 25.192 3.616 25.224 ;
  LAYER M2 ;
        RECT 5.952 25.128 5.984 25.16 ;
  LAYER M2 ;
        RECT 3.584 25.064 3.616 25.096 ;
  LAYER M2 ;
        RECT 3.536 24.864 6.032 27.468 ;
  LAYER M1 ;
        RECT 5.952 21.804 5.984 24.312 ;
  LAYER M3 ;
        RECT 5.952 21.824 5.984 21.856 ;
  LAYER M1 ;
        RECT 5.888 21.804 5.92 24.312 ;
  LAYER M3 ;
        RECT 5.888 24.26 5.92 24.292 ;
  LAYER M1 ;
        RECT 5.824 21.804 5.856 24.312 ;
  LAYER M3 ;
        RECT 5.824 21.824 5.856 21.856 ;
  LAYER M1 ;
        RECT 5.76 21.804 5.792 24.312 ;
  LAYER M3 ;
        RECT 5.76 24.26 5.792 24.292 ;
  LAYER M1 ;
        RECT 5.696 21.804 5.728 24.312 ;
  LAYER M3 ;
        RECT 5.696 21.824 5.728 21.856 ;
  LAYER M1 ;
        RECT 5.632 21.804 5.664 24.312 ;
  LAYER M3 ;
        RECT 5.632 24.26 5.664 24.292 ;
  LAYER M1 ;
        RECT 5.568 21.804 5.6 24.312 ;
  LAYER M3 ;
        RECT 5.568 21.824 5.6 21.856 ;
  LAYER M1 ;
        RECT 5.504 21.804 5.536 24.312 ;
  LAYER M3 ;
        RECT 5.504 24.26 5.536 24.292 ;
  LAYER M1 ;
        RECT 5.44 21.804 5.472 24.312 ;
  LAYER M3 ;
        RECT 5.44 21.824 5.472 21.856 ;
  LAYER M1 ;
        RECT 5.376 21.804 5.408 24.312 ;
  LAYER M3 ;
        RECT 5.376 24.26 5.408 24.292 ;
  LAYER M1 ;
        RECT 5.312 21.804 5.344 24.312 ;
  LAYER M3 ;
        RECT 5.312 21.824 5.344 21.856 ;
  LAYER M1 ;
        RECT 5.248 21.804 5.28 24.312 ;
  LAYER M3 ;
        RECT 5.248 24.26 5.28 24.292 ;
  LAYER M1 ;
        RECT 5.184 21.804 5.216 24.312 ;
  LAYER M3 ;
        RECT 5.184 21.824 5.216 21.856 ;
  LAYER M1 ;
        RECT 5.12 21.804 5.152 24.312 ;
  LAYER M3 ;
        RECT 5.12 24.26 5.152 24.292 ;
  LAYER M1 ;
        RECT 5.056 21.804 5.088 24.312 ;
  LAYER M3 ;
        RECT 5.056 21.824 5.088 21.856 ;
  LAYER M1 ;
        RECT 4.992 21.804 5.024 24.312 ;
  LAYER M3 ;
        RECT 4.992 24.26 5.024 24.292 ;
  LAYER M1 ;
        RECT 4.928 21.804 4.96 24.312 ;
  LAYER M3 ;
        RECT 4.928 21.824 4.96 21.856 ;
  LAYER M1 ;
        RECT 4.864 21.804 4.896 24.312 ;
  LAYER M3 ;
        RECT 4.864 24.26 4.896 24.292 ;
  LAYER M1 ;
        RECT 4.8 21.804 4.832 24.312 ;
  LAYER M3 ;
        RECT 4.8 21.824 4.832 21.856 ;
  LAYER M1 ;
        RECT 4.736 21.804 4.768 24.312 ;
  LAYER M3 ;
        RECT 4.736 24.26 4.768 24.292 ;
  LAYER M1 ;
        RECT 4.672 21.804 4.704 24.312 ;
  LAYER M3 ;
        RECT 4.672 21.824 4.704 21.856 ;
  LAYER M1 ;
        RECT 4.608 21.804 4.64 24.312 ;
  LAYER M3 ;
        RECT 4.608 24.26 4.64 24.292 ;
  LAYER M1 ;
        RECT 4.544 21.804 4.576 24.312 ;
  LAYER M3 ;
        RECT 4.544 21.824 4.576 21.856 ;
  LAYER M1 ;
        RECT 4.48 21.804 4.512 24.312 ;
  LAYER M3 ;
        RECT 4.48 24.26 4.512 24.292 ;
  LAYER M1 ;
        RECT 4.416 21.804 4.448 24.312 ;
  LAYER M3 ;
        RECT 4.416 21.824 4.448 21.856 ;
  LAYER M1 ;
        RECT 4.352 21.804 4.384 24.312 ;
  LAYER M3 ;
        RECT 4.352 24.26 4.384 24.292 ;
  LAYER M1 ;
        RECT 4.288 21.804 4.32 24.312 ;
  LAYER M3 ;
        RECT 4.288 21.824 4.32 21.856 ;
  LAYER M1 ;
        RECT 4.224 21.804 4.256 24.312 ;
  LAYER M3 ;
        RECT 4.224 24.26 4.256 24.292 ;
  LAYER M1 ;
        RECT 4.16 21.804 4.192 24.312 ;
  LAYER M3 ;
        RECT 4.16 21.824 4.192 21.856 ;
  LAYER M1 ;
        RECT 4.096 21.804 4.128 24.312 ;
  LAYER M3 ;
        RECT 4.096 24.26 4.128 24.292 ;
  LAYER M1 ;
        RECT 4.032 21.804 4.064 24.312 ;
  LAYER M3 ;
        RECT 4.032 21.824 4.064 21.856 ;
  LAYER M1 ;
        RECT 3.968 21.804 4 24.312 ;
  LAYER M3 ;
        RECT 3.968 24.26 4 24.292 ;
  LAYER M1 ;
        RECT 3.904 21.804 3.936 24.312 ;
  LAYER M3 ;
        RECT 3.904 21.824 3.936 21.856 ;
  LAYER M1 ;
        RECT 3.84 21.804 3.872 24.312 ;
  LAYER M3 ;
        RECT 3.84 24.26 3.872 24.292 ;
  LAYER M1 ;
        RECT 3.776 21.804 3.808 24.312 ;
  LAYER M3 ;
        RECT 3.776 21.824 3.808 21.856 ;
  LAYER M1 ;
        RECT 3.712 21.804 3.744 24.312 ;
  LAYER M3 ;
        RECT 3.712 24.26 3.744 24.292 ;
  LAYER M1 ;
        RECT 3.648 21.804 3.68 24.312 ;
  LAYER M3 ;
        RECT 3.648 21.824 3.68 21.856 ;
  LAYER M1 ;
        RECT 3.584 21.804 3.616 24.312 ;
  LAYER M3 ;
        RECT 5.952 24.196 5.984 24.228 ;
  LAYER M2 ;
        RECT 3.584 24.132 3.616 24.164 ;
  LAYER M2 ;
        RECT 5.952 24.068 5.984 24.1 ;
  LAYER M2 ;
        RECT 3.584 24.004 3.616 24.036 ;
  LAYER M2 ;
        RECT 5.952 23.94 5.984 23.972 ;
  LAYER M2 ;
        RECT 3.584 23.876 3.616 23.908 ;
  LAYER M2 ;
        RECT 5.952 23.812 5.984 23.844 ;
  LAYER M2 ;
        RECT 3.584 23.748 3.616 23.78 ;
  LAYER M2 ;
        RECT 5.952 23.684 5.984 23.716 ;
  LAYER M2 ;
        RECT 3.584 23.62 3.616 23.652 ;
  LAYER M2 ;
        RECT 5.952 23.556 5.984 23.588 ;
  LAYER M2 ;
        RECT 3.584 23.492 3.616 23.524 ;
  LAYER M2 ;
        RECT 5.952 23.428 5.984 23.46 ;
  LAYER M2 ;
        RECT 3.584 23.364 3.616 23.396 ;
  LAYER M2 ;
        RECT 5.952 23.3 5.984 23.332 ;
  LAYER M2 ;
        RECT 3.584 23.236 3.616 23.268 ;
  LAYER M2 ;
        RECT 5.952 23.172 5.984 23.204 ;
  LAYER M2 ;
        RECT 3.584 23.108 3.616 23.14 ;
  LAYER M2 ;
        RECT 5.952 23.044 5.984 23.076 ;
  LAYER M2 ;
        RECT 3.584 22.98 3.616 23.012 ;
  LAYER M2 ;
        RECT 5.952 22.916 5.984 22.948 ;
  LAYER M2 ;
        RECT 3.584 22.852 3.616 22.884 ;
  LAYER M2 ;
        RECT 5.952 22.788 5.984 22.82 ;
  LAYER M2 ;
        RECT 3.584 22.724 3.616 22.756 ;
  LAYER M2 ;
        RECT 5.952 22.66 5.984 22.692 ;
  LAYER M2 ;
        RECT 3.584 22.596 3.616 22.628 ;
  LAYER M2 ;
        RECT 5.952 22.532 5.984 22.564 ;
  LAYER M2 ;
        RECT 3.584 22.468 3.616 22.5 ;
  LAYER M2 ;
        RECT 5.952 22.404 5.984 22.436 ;
  LAYER M2 ;
        RECT 3.584 22.34 3.616 22.372 ;
  LAYER M2 ;
        RECT 5.952 22.276 5.984 22.308 ;
  LAYER M2 ;
        RECT 3.584 22.212 3.616 22.244 ;
  LAYER M2 ;
        RECT 5.952 22.148 5.984 22.18 ;
  LAYER M2 ;
        RECT 3.584 22.084 3.616 22.116 ;
  LAYER M2 ;
        RECT 5.952 22.02 5.984 22.052 ;
  LAYER M2 ;
        RECT 3.584 21.956 3.616 21.988 ;
  LAYER M2 ;
        RECT 3.536 21.756 6.032 24.36 ;
  LAYER M1 ;
        RECT 5.952 18.696 5.984 21.204 ;
  LAYER M3 ;
        RECT 5.952 18.716 5.984 18.748 ;
  LAYER M1 ;
        RECT 5.888 18.696 5.92 21.204 ;
  LAYER M3 ;
        RECT 5.888 21.152 5.92 21.184 ;
  LAYER M1 ;
        RECT 5.824 18.696 5.856 21.204 ;
  LAYER M3 ;
        RECT 5.824 18.716 5.856 18.748 ;
  LAYER M1 ;
        RECT 5.76 18.696 5.792 21.204 ;
  LAYER M3 ;
        RECT 5.76 21.152 5.792 21.184 ;
  LAYER M1 ;
        RECT 5.696 18.696 5.728 21.204 ;
  LAYER M3 ;
        RECT 5.696 18.716 5.728 18.748 ;
  LAYER M1 ;
        RECT 5.632 18.696 5.664 21.204 ;
  LAYER M3 ;
        RECT 5.632 21.152 5.664 21.184 ;
  LAYER M1 ;
        RECT 5.568 18.696 5.6 21.204 ;
  LAYER M3 ;
        RECT 5.568 18.716 5.6 18.748 ;
  LAYER M1 ;
        RECT 5.504 18.696 5.536 21.204 ;
  LAYER M3 ;
        RECT 5.504 21.152 5.536 21.184 ;
  LAYER M1 ;
        RECT 5.44 18.696 5.472 21.204 ;
  LAYER M3 ;
        RECT 5.44 18.716 5.472 18.748 ;
  LAYER M1 ;
        RECT 5.376 18.696 5.408 21.204 ;
  LAYER M3 ;
        RECT 5.376 21.152 5.408 21.184 ;
  LAYER M1 ;
        RECT 5.312 18.696 5.344 21.204 ;
  LAYER M3 ;
        RECT 5.312 18.716 5.344 18.748 ;
  LAYER M1 ;
        RECT 5.248 18.696 5.28 21.204 ;
  LAYER M3 ;
        RECT 5.248 21.152 5.28 21.184 ;
  LAYER M1 ;
        RECT 5.184 18.696 5.216 21.204 ;
  LAYER M3 ;
        RECT 5.184 18.716 5.216 18.748 ;
  LAYER M1 ;
        RECT 5.12 18.696 5.152 21.204 ;
  LAYER M3 ;
        RECT 5.12 21.152 5.152 21.184 ;
  LAYER M1 ;
        RECT 5.056 18.696 5.088 21.204 ;
  LAYER M3 ;
        RECT 5.056 18.716 5.088 18.748 ;
  LAYER M1 ;
        RECT 4.992 18.696 5.024 21.204 ;
  LAYER M3 ;
        RECT 4.992 21.152 5.024 21.184 ;
  LAYER M1 ;
        RECT 4.928 18.696 4.96 21.204 ;
  LAYER M3 ;
        RECT 4.928 18.716 4.96 18.748 ;
  LAYER M1 ;
        RECT 4.864 18.696 4.896 21.204 ;
  LAYER M3 ;
        RECT 4.864 21.152 4.896 21.184 ;
  LAYER M1 ;
        RECT 4.8 18.696 4.832 21.204 ;
  LAYER M3 ;
        RECT 4.8 18.716 4.832 18.748 ;
  LAYER M1 ;
        RECT 4.736 18.696 4.768 21.204 ;
  LAYER M3 ;
        RECT 4.736 21.152 4.768 21.184 ;
  LAYER M1 ;
        RECT 4.672 18.696 4.704 21.204 ;
  LAYER M3 ;
        RECT 4.672 18.716 4.704 18.748 ;
  LAYER M1 ;
        RECT 4.608 18.696 4.64 21.204 ;
  LAYER M3 ;
        RECT 4.608 21.152 4.64 21.184 ;
  LAYER M1 ;
        RECT 4.544 18.696 4.576 21.204 ;
  LAYER M3 ;
        RECT 4.544 18.716 4.576 18.748 ;
  LAYER M1 ;
        RECT 4.48 18.696 4.512 21.204 ;
  LAYER M3 ;
        RECT 4.48 21.152 4.512 21.184 ;
  LAYER M1 ;
        RECT 4.416 18.696 4.448 21.204 ;
  LAYER M3 ;
        RECT 4.416 18.716 4.448 18.748 ;
  LAYER M1 ;
        RECT 4.352 18.696 4.384 21.204 ;
  LAYER M3 ;
        RECT 4.352 21.152 4.384 21.184 ;
  LAYER M1 ;
        RECT 4.288 18.696 4.32 21.204 ;
  LAYER M3 ;
        RECT 4.288 18.716 4.32 18.748 ;
  LAYER M1 ;
        RECT 4.224 18.696 4.256 21.204 ;
  LAYER M3 ;
        RECT 4.224 21.152 4.256 21.184 ;
  LAYER M1 ;
        RECT 4.16 18.696 4.192 21.204 ;
  LAYER M3 ;
        RECT 4.16 18.716 4.192 18.748 ;
  LAYER M1 ;
        RECT 4.096 18.696 4.128 21.204 ;
  LAYER M3 ;
        RECT 4.096 21.152 4.128 21.184 ;
  LAYER M1 ;
        RECT 4.032 18.696 4.064 21.204 ;
  LAYER M3 ;
        RECT 4.032 18.716 4.064 18.748 ;
  LAYER M1 ;
        RECT 3.968 18.696 4 21.204 ;
  LAYER M3 ;
        RECT 3.968 21.152 4 21.184 ;
  LAYER M1 ;
        RECT 3.904 18.696 3.936 21.204 ;
  LAYER M3 ;
        RECT 3.904 18.716 3.936 18.748 ;
  LAYER M1 ;
        RECT 3.84 18.696 3.872 21.204 ;
  LAYER M3 ;
        RECT 3.84 21.152 3.872 21.184 ;
  LAYER M1 ;
        RECT 3.776 18.696 3.808 21.204 ;
  LAYER M3 ;
        RECT 3.776 18.716 3.808 18.748 ;
  LAYER M1 ;
        RECT 3.712 18.696 3.744 21.204 ;
  LAYER M3 ;
        RECT 3.712 21.152 3.744 21.184 ;
  LAYER M1 ;
        RECT 3.648 18.696 3.68 21.204 ;
  LAYER M3 ;
        RECT 3.648 18.716 3.68 18.748 ;
  LAYER M1 ;
        RECT 3.584 18.696 3.616 21.204 ;
  LAYER M3 ;
        RECT 5.952 21.088 5.984 21.12 ;
  LAYER M2 ;
        RECT 3.584 21.024 3.616 21.056 ;
  LAYER M2 ;
        RECT 5.952 20.96 5.984 20.992 ;
  LAYER M2 ;
        RECT 3.584 20.896 3.616 20.928 ;
  LAYER M2 ;
        RECT 5.952 20.832 5.984 20.864 ;
  LAYER M2 ;
        RECT 3.584 20.768 3.616 20.8 ;
  LAYER M2 ;
        RECT 5.952 20.704 5.984 20.736 ;
  LAYER M2 ;
        RECT 3.584 20.64 3.616 20.672 ;
  LAYER M2 ;
        RECT 5.952 20.576 5.984 20.608 ;
  LAYER M2 ;
        RECT 3.584 20.512 3.616 20.544 ;
  LAYER M2 ;
        RECT 5.952 20.448 5.984 20.48 ;
  LAYER M2 ;
        RECT 3.584 20.384 3.616 20.416 ;
  LAYER M2 ;
        RECT 5.952 20.32 5.984 20.352 ;
  LAYER M2 ;
        RECT 3.584 20.256 3.616 20.288 ;
  LAYER M2 ;
        RECT 5.952 20.192 5.984 20.224 ;
  LAYER M2 ;
        RECT 3.584 20.128 3.616 20.16 ;
  LAYER M2 ;
        RECT 5.952 20.064 5.984 20.096 ;
  LAYER M2 ;
        RECT 3.584 20 3.616 20.032 ;
  LAYER M2 ;
        RECT 5.952 19.936 5.984 19.968 ;
  LAYER M2 ;
        RECT 3.584 19.872 3.616 19.904 ;
  LAYER M2 ;
        RECT 5.952 19.808 5.984 19.84 ;
  LAYER M2 ;
        RECT 3.584 19.744 3.616 19.776 ;
  LAYER M2 ;
        RECT 5.952 19.68 5.984 19.712 ;
  LAYER M2 ;
        RECT 3.584 19.616 3.616 19.648 ;
  LAYER M2 ;
        RECT 5.952 19.552 5.984 19.584 ;
  LAYER M2 ;
        RECT 3.584 19.488 3.616 19.52 ;
  LAYER M2 ;
        RECT 5.952 19.424 5.984 19.456 ;
  LAYER M2 ;
        RECT 3.584 19.36 3.616 19.392 ;
  LAYER M2 ;
        RECT 5.952 19.296 5.984 19.328 ;
  LAYER M2 ;
        RECT 3.584 19.232 3.616 19.264 ;
  LAYER M2 ;
        RECT 5.952 19.168 5.984 19.2 ;
  LAYER M2 ;
        RECT 3.584 19.104 3.616 19.136 ;
  LAYER M2 ;
        RECT 5.952 19.04 5.984 19.072 ;
  LAYER M2 ;
        RECT 3.584 18.976 3.616 19.008 ;
  LAYER M2 ;
        RECT 5.952 18.912 5.984 18.944 ;
  LAYER M2 ;
        RECT 3.584 18.848 3.616 18.88 ;
  LAYER M2 ;
        RECT 3.536 18.648 6.032 21.252 ;
  LAYER M1 ;
        RECT 5.952 15.588 5.984 18.096 ;
  LAYER M3 ;
        RECT 5.952 15.608 5.984 15.64 ;
  LAYER M1 ;
        RECT 5.888 15.588 5.92 18.096 ;
  LAYER M3 ;
        RECT 5.888 18.044 5.92 18.076 ;
  LAYER M1 ;
        RECT 5.824 15.588 5.856 18.096 ;
  LAYER M3 ;
        RECT 5.824 15.608 5.856 15.64 ;
  LAYER M1 ;
        RECT 5.76 15.588 5.792 18.096 ;
  LAYER M3 ;
        RECT 5.76 18.044 5.792 18.076 ;
  LAYER M1 ;
        RECT 5.696 15.588 5.728 18.096 ;
  LAYER M3 ;
        RECT 5.696 15.608 5.728 15.64 ;
  LAYER M1 ;
        RECT 5.632 15.588 5.664 18.096 ;
  LAYER M3 ;
        RECT 5.632 18.044 5.664 18.076 ;
  LAYER M1 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M3 ;
        RECT 5.568 15.608 5.6 15.64 ;
  LAYER M1 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M3 ;
        RECT 5.504 18.044 5.536 18.076 ;
  LAYER M1 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M3 ;
        RECT 5.44 15.608 5.472 15.64 ;
  LAYER M1 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M3 ;
        RECT 5.376 18.044 5.408 18.076 ;
  LAYER M1 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M3 ;
        RECT 5.312 15.608 5.344 15.64 ;
  LAYER M1 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M3 ;
        RECT 5.248 18.044 5.28 18.076 ;
  LAYER M1 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M3 ;
        RECT 5.184 15.608 5.216 15.64 ;
  LAYER M1 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M3 ;
        RECT 5.12 18.044 5.152 18.076 ;
  LAYER M1 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M3 ;
        RECT 5.056 15.608 5.088 15.64 ;
  LAYER M1 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M3 ;
        RECT 4.992 18.044 5.024 18.076 ;
  LAYER M1 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M3 ;
        RECT 4.928 15.608 4.96 15.64 ;
  LAYER M1 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M3 ;
        RECT 4.864 18.044 4.896 18.076 ;
  LAYER M1 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M3 ;
        RECT 4.8 15.608 4.832 15.64 ;
  LAYER M1 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M3 ;
        RECT 4.736 18.044 4.768 18.076 ;
  LAYER M1 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M3 ;
        RECT 4.672 15.608 4.704 15.64 ;
  LAYER M1 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M3 ;
        RECT 4.608 18.044 4.64 18.076 ;
  LAYER M1 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M3 ;
        RECT 4.544 15.608 4.576 15.64 ;
  LAYER M1 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M3 ;
        RECT 4.48 18.044 4.512 18.076 ;
  LAYER M1 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M3 ;
        RECT 4.416 15.608 4.448 15.64 ;
  LAYER M1 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M3 ;
        RECT 4.352 18.044 4.384 18.076 ;
  LAYER M1 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M3 ;
        RECT 4.288 15.608 4.32 15.64 ;
  LAYER M1 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M3 ;
        RECT 4.224 18.044 4.256 18.076 ;
  LAYER M1 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M3 ;
        RECT 4.16 15.608 4.192 15.64 ;
  LAYER M1 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M3 ;
        RECT 4.096 18.044 4.128 18.076 ;
  LAYER M1 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M3 ;
        RECT 4.032 15.608 4.064 15.64 ;
  LAYER M1 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M3 ;
        RECT 3.968 18.044 4 18.076 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M3 ;
        RECT 3.904 15.608 3.936 15.64 ;
  LAYER M1 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M3 ;
        RECT 3.84 18.044 3.872 18.076 ;
  LAYER M1 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M3 ;
        RECT 3.776 15.608 3.808 15.64 ;
  LAYER M1 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M3 ;
        RECT 3.712 18.044 3.744 18.076 ;
  LAYER M1 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M3 ;
        RECT 3.648 15.608 3.68 15.64 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M3 ;
        RECT 5.952 17.98 5.984 18.012 ;
  LAYER M2 ;
        RECT 3.584 17.916 3.616 17.948 ;
  LAYER M2 ;
        RECT 5.952 17.852 5.984 17.884 ;
  LAYER M2 ;
        RECT 3.584 17.788 3.616 17.82 ;
  LAYER M2 ;
        RECT 5.952 17.724 5.984 17.756 ;
  LAYER M2 ;
        RECT 3.584 17.66 3.616 17.692 ;
  LAYER M2 ;
        RECT 5.952 17.596 5.984 17.628 ;
  LAYER M2 ;
        RECT 3.584 17.532 3.616 17.564 ;
  LAYER M2 ;
        RECT 5.952 17.468 5.984 17.5 ;
  LAYER M2 ;
        RECT 3.584 17.404 3.616 17.436 ;
  LAYER M2 ;
        RECT 5.952 17.34 5.984 17.372 ;
  LAYER M2 ;
        RECT 3.584 17.276 3.616 17.308 ;
  LAYER M2 ;
        RECT 5.952 17.212 5.984 17.244 ;
  LAYER M2 ;
        RECT 3.584 17.148 3.616 17.18 ;
  LAYER M2 ;
        RECT 5.952 17.084 5.984 17.116 ;
  LAYER M2 ;
        RECT 3.584 17.02 3.616 17.052 ;
  LAYER M2 ;
        RECT 5.952 16.956 5.984 16.988 ;
  LAYER M2 ;
        RECT 3.584 16.892 3.616 16.924 ;
  LAYER M2 ;
        RECT 5.952 16.828 5.984 16.86 ;
  LAYER M2 ;
        RECT 3.584 16.764 3.616 16.796 ;
  LAYER M2 ;
        RECT 5.952 16.7 5.984 16.732 ;
  LAYER M2 ;
        RECT 3.584 16.636 3.616 16.668 ;
  LAYER M2 ;
        RECT 5.952 16.572 5.984 16.604 ;
  LAYER M2 ;
        RECT 3.584 16.508 3.616 16.54 ;
  LAYER M2 ;
        RECT 5.952 16.444 5.984 16.476 ;
  LAYER M2 ;
        RECT 3.584 16.38 3.616 16.412 ;
  LAYER M2 ;
        RECT 5.952 16.316 5.984 16.348 ;
  LAYER M2 ;
        RECT 3.584 16.252 3.616 16.284 ;
  LAYER M2 ;
        RECT 5.952 16.188 5.984 16.22 ;
  LAYER M2 ;
        RECT 3.584 16.124 3.616 16.156 ;
  LAYER M2 ;
        RECT 5.952 16.06 5.984 16.092 ;
  LAYER M2 ;
        RECT 3.584 15.996 3.616 16.028 ;
  LAYER M2 ;
        RECT 5.952 15.932 5.984 15.964 ;
  LAYER M2 ;
        RECT 3.584 15.868 3.616 15.9 ;
  LAYER M2 ;
        RECT 5.952 15.804 5.984 15.836 ;
  LAYER M2 ;
        RECT 3.584 15.74 3.616 15.772 ;
  LAYER M2 ;
        RECT 3.536 15.54 6.032 18.144 ;
  LAYER M1 ;
        RECT 2.976 28.02 3.008 30.528 ;
  LAYER M3 ;
        RECT 2.976 28.04 3.008 28.072 ;
  LAYER M1 ;
        RECT 2.912 28.02 2.944 30.528 ;
  LAYER M3 ;
        RECT 2.912 30.476 2.944 30.508 ;
  LAYER M1 ;
        RECT 2.848 28.02 2.88 30.528 ;
  LAYER M3 ;
        RECT 2.848 28.04 2.88 28.072 ;
  LAYER M1 ;
        RECT 2.784 28.02 2.816 30.528 ;
  LAYER M3 ;
        RECT 2.784 30.476 2.816 30.508 ;
  LAYER M1 ;
        RECT 2.72 28.02 2.752 30.528 ;
  LAYER M3 ;
        RECT 2.72 28.04 2.752 28.072 ;
  LAYER M1 ;
        RECT 2.656 28.02 2.688 30.528 ;
  LAYER M3 ;
        RECT 2.656 30.476 2.688 30.508 ;
  LAYER M1 ;
        RECT 2.592 28.02 2.624 30.528 ;
  LAYER M3 ;
        RECT 2.592 28.04 2.624 28.072 ;
  LAYER M1 ;
        RECT 2.528 28.02 2.56 30.528 ;
  LAYER M3 ;
        RECT 2.528 30.476 2.56 30.508 ;
  LAYER M1 ;
        RECT 2.464 28.02 2.496 30.528 ;
  LAYER M3 ;
        RECT 2.464 28.04 2.496 28.072 ;
  LAYER M1 ;
        RECT 2.4 28.02 2.432 30.528 ;
  LAYER M3 ;
        RECT 2.4 30.476 2.432 30.508 ;
  LAYER M1 ;
        RECT 2.336 28.02 2.368 30.528 ;
  LAYER M3 ;
        RECT 2.336 28.04 2.368 28.072 ;
  LAYER M1 ;
        RECT 2.272 28.02 2.304 30.528 ;
  LAYER M3 ;
        RECT 2.272 30.476 2.304 30.508 ;
  LAYER M1 ;
        RECT 2.208 28.02 2.24 30.528 ;
  LAYER M3 ;
        RECT 2.208 28.04 2.24 28.072 ;
  LAYER M1 ;
        RECT 2.144 28.02 2.176 30.528 ;
  LAYER M3 ;
        RECT 2.144 30.476 2.176 30.508 ;
  LAYER M1 ;
        RECT 2.08 28.02 2.112 30.528 ;
  LAYER M3 ;
        RECT 2.08 28.04 2.112 28.072 ;
  LAYER M1 ;
        RECT 2.016 28.02 2.048 30.528 ;
  LAYER M3 ;
        RECT 2.016 30.476 2.048 30.508 ;
  LAYER M1 ;
        RECT 1.952 28.02 1.984 30.528 ;
  LAYER M3 ;
        RECT 1.952 28.04 1.984 28.072 ;
  LAYER M1 ;
        RECT 1.888 28.02 1.92 30.528 ;
  LAYER M3 ;
        RECT 1.888 30.476 1.92 30.508 ;
  LAYER M1 ;
        RECT 1.824 28.02 1.856 30.528 ;
  LAYER M3 ;
        RECT 1.824 28.04 1.856 28.072 ;
  LAYER M1 ;
        RECT 1.76 28.02 1.792 30.528 ;
  LAYER M3 ;
        RECT 1.76 30.476 1.792 30.508 ;
  LAYER M1 ;
        RECT 1.696 28.02 1.728 30.528 ;
  LAYER M3 ;
        RECT 1.696 28.04 1.728 28.072 ;
  LAYER M1 ;
        RECT 1.632 28.02 1.664 30.528 ;
  LAYER M3 ;
        RECT 1.632 30.476 1.664 30.508 ;
  LAYER M1 ;
        RECT 1.568 28.02 1.6 30.528 ;
  LAYER M3 ;
        RECT 1.568 28.04 1.6 28.072 ;
  LAYER M1 ;
        RECT 1.504 28.02 1.536 30.528 ;
  LAYER M3 ;
        RECT 1.504 30.476 1.536 30.508 ;
  LAYER M1 ;
        RECT 1.44 28.02 1.472 30.528 ;
  LAYER M3 ;
        RECT 1.44 28.04 1.472 28.072 ;
  LAYER M1 ;
        RECT 1.376 28.02 1.408 30.528 ;
  LAYER M3 ;
        RECT 1.376 30.476 1.408 30.508 ;
  LAYER M1 ;
        RECT 1.312 28.02 1.344 30.528 ;
  LAYER M3 ;
        RECT 1.312 28.04 1.344 28.072 ;
  LAYER M1 ;
        RECT 1.248 28.02 1.28 30.528 ;
  LAYER M3 ;
        RECT 1.248 30.476 1.28 30.508 ;
  LAYER M1 ;
        RECT 1.184 28.02 1.216 30.528 ;
  LAYER M3 ;
        RECT 1.184 28.04 1.216 28.072 ;
  LAYER M1 ;
        RECT 1.12 28.02 1.152 30.528 ;
  LAYER M3 ;
        RECT 1.12 30.476 1.152 30.508 ;
  LAYER M1 ;
        RECT 1.056 28.02 1.088 30.528 ;
  LAYER M3 ;
        RECT 1.056 28.04 1.088 28.072 ;
  LAYER M1 ;
        RECT 0.992 28.02 1.024 30.528 ;
  LAYER M3 ;
        RECT 0.992 30.476 1.024 30.508 ;
  LAYER M1 ;
        RECT 0.928 28.02 0.96 30.528 ;
  LAYER M3 ;
        RECT 0.928 28.04 0.96 28.072 ;
  LAYER M1 ;
        RECT 0.864 28.02 0.896 30.528 ;
  LAYER M3 ;
        RECT 0.864 30.476 0.896 30.508 ;
  LAYER M1 ;
        RECT 0.8 28.02 0.832 30.528 ;
  LAYER M3 ;
        RECT 0.8 28.04 0.832 28.072 ;
  LAYER M1 ;
        RECT 0.736 28.02 0.768 30.528 ;
  LAYER M3 ;
        RECT 0.736 30.476 0.768 30.508 ;
  LAYER M1 ;
        RECT 0.672 28.02 0.704 30.528 ;
  LAYER M3 ;
        RECT 0.672 28.04 0.704 28.072 ;
  LAYER M1 ;
        RECT 0.608 28.02 0.64 30.528 ;
  LAYER M3 ;
        RECT 2.976 30.412 3.008 30.444 ;
  LAYER M2 ;
        RECT 0.608 30.348 0.64 30.38 ;
  LAYER M2 ;
        RECT 2.976 30.284 3.008 30.316 ;
  LAYER M2 ;
        RECT 0.608 30.22 0.64 30.252 ;
  LAYER M2 ;
        RECT 2.976 30.156 3.008 30.188 ;
  LAYER M2 ;
        RECT 0.608 30.092 0.64 30.124 ;
  LAYER M2 ;
        RECT 2.976 30.028 3.008 30.06 ;
  LAYER M2 ;
        RECT 0.608 29.964 0.64 29.996 ;
  LAYER M2 ;
        RECT 2.976 29.9 3.008 29.932 ;
  LAYER M2 ;
        RECT 0.608 29.836 0.64 29.868 ;
  LAYER M2 ;
        RECT 2.976 29.772 3.008 29.804 ;
  LAYER M2 ;
        RECT 0.608 29.708 0.64 29.74 ;
  LAYER M2 ;
        RECT 2.976 29.644 3.008 29.676 ;
  LAYER M2 ;
        RECT 0.608 29.58 0.64 29.612 ;
  LAYER M2 ;
        RECT 2.976 29.516 3.008 29.548 ;
  LAYER M2 ;
        RECT 0.608 29.452 0.64 29.484 ;
  LAYER M2 ;
        RECT 2.976 29.388 3.008 29.42 ;
  LAYER M2 ;
        RECT 0.608 29.324 0.64 29.356 ;
  LAYER M2 ;
        RECT 2.976 29.26 3.008 29.292 ;
  LAYER M2 ;
        RECT 0.608 29.196 0.64 29.228 ;
  LAYER M2 ;
        RECT 2.976 29.132 3.008 29.164 ;
  LAYER M2 ;
        RECT 0.608 29.068 0.64 29.1 ;
  LAYER M2 ;
        RECT 2.976 29.004 3.008 29.036 ;
  LAYER M2 ;
        RECT 0.608 28.94 0.64 28.972 ;
  LAYER M2 ;
        RECT 2.976 28.876 3.008 28.908 ;
  LAYER M2 ;
        RECT 0.608 28.812 0.64 28.844 ;
  LAYER M2 ;
        RECT 2.976 28.748 3.008 28.78 ;
  LAYER M2 ;
        RECT 0.608 28.684 0.64 28.716 ;
  LAYER M2 ;
        RECT 2.976 28.62 3.008 28.652 ;
  LAYER M2 ;
        RECT 0.608 28.556 0.64 28.588 ;
  LAYER M2 ;
        RECT 2.976 28.492 3.008 28.524 ;
  LAYER M2 ;
        RECT 0.608 28.428 0.64 28.46 ;
  LAYER M2 ;
        RECT 2.976 28.364 3.008 28.396 ;
  LAYER M2 ;
        RECT 0.608 28.3 0.64 28.332 ;
  LAYER M2 ;
        RECT 2.976 28.236 3.008 28.268 ;
  LAYER M2 ;
        RECT 0.608 28.172 0.64 28.204 ;
  LAYER M2 ;
        RECT 0.56 27.972 3.056 30.576 ;
  LAYER M1 ;
        RECT 2.976 24.912 3.008 27.42 ;
  LAYER M3 ;
        RECT 2.976 24.932 3.008 24.964 ;
  LAYER M1 ;
        RECT 2.912 24.912 2.944 27.42 ;
  LAYER M3 ;
        RECT 2.912 27.368 2.944 27.4 ;
  LAYER M1 ;
        RECT 2.848 24.912 2.88 27.42 ;
  LAYER M3 ;
        RECT 2.848 24.932 2.88 24.964 ;
  LAYER M1 ;
        RECT 2.784 24.912 2.816 27.42 ;
  LAYER M3 ;
        RECT 2.784 27.368 2.816 27.4 ;
  LAYER M1 ;
        RECT 2.72 24.912 2.752 27.42 ;
  LAYER M3 ;
        RECT 2.72 24.932 2.752 24.964 ;
  LAYER M1 ;
        RECT 2.656 24.912 2.688 27.42 ;
  LAYER M3 ;
        RECT 2.656 27.368 2.688 27.4 ;
  LAYER M1 ;
        RECT 2.592 24.912 2.624 27.42 ;
  LAYER M3 ;
        RECT 2.592 24.932 2.624 24.964 ;
  LAYER M1 ;
        RECT 2.528 24.912 2.56 27.42 ;
  LAYER M3 ;
        RECT 2.528 27.368 2.56 27.4 ;
  LAYER M1 ;
        RECT 2.464 24.912 2.496 27.42 ;
  LAYER M3 ;
        RECT 2.464 24.932 2.496 24.964 ;
  LAYER M1 ;
        RECT 2.4 24.912 2.432 27.42 ;
  LAYER M3 ;
        RECT 2.4 27.368 2.432 27.4 ;
  LAYER M1 ;
        RECT 2.336 24.912 2.368 27.42 ;
  LAYER M3 ;
        RECT 2.336 24.932 2.368 24.964 ;
  LAYER M1 ;
        RECT 2.272 24.912 2.304 27.42 ;
  LAYER M3 ;
        RECT 2.272 27.368 2.304 27.4 ;
  LAYER M1 ;
        RECT 2.208 24.912 2.24 27.42 ;
  LAYER M3 ;
        RECT 2.208 24.932 2.24 24.964 ;
  LAYER M1 ;
        RECT 2.144 24.912 2.176 27.42 ;
  LAYER M3 ;
        RECT 2.144 27.368 2.176 27.4 ;
  LAYER M1 ;
        RECT 2.08 24.912 2.112 27.42 ;
  LAYER M3 ;
        RECT 2.08 24.932 2.112 24.964 ;
  LAYER M1 ;
        RECT 2.016 24.912 2.048 27.42 ;
  LAYER M3 ;
        RECT 2.016 27.368 2.048 27.4 ;
  LAYER M1 ;
        RECT 1.952 24.912 1.984 27.42 ;
  LAYER M3 ;
        RECT 1.952 24.932 1.984 24.964 ;
  LAYER M1 ;
        RECT 1.888 24.912 1.92 27.42 ;
  LAYER M3 ;
        RECT 1.888 27.368 1.92 27.4 ;
  LAYER M1 ;
        RECT 1.824 24.912 1.856 27.42 ;
  LAYER M3 ;
        RECT 1.824 24.932 1.856 24.964 ;
  LAYER M1 ;
        RECT 1.76 24.912 1.792 27.42 ;
  LAYER M3 ;
        RECT 1.76 27.368 1.792 27.4 ;
  LAYER M1 ;
        RECT 1.696 24.912 1.728 27.42 ;
  LAYER M3 ;
        RECT 1.696 24.932 1.728 24.964 ;
  LAYER M1 ;
        RECT 1.632 24.912 1.664 27.42 ;
  LAYER M3 ;
        RECT 1.632 27.368 1.664 27.4 ;
  LAYER M1 ;
        RECT 1.568 24.912 1.6 27.42 ;
  LAYER M3 ;
        RECT 1.568 24.932 1.6 24.964 ;
  LAYER M1 ;
        RECT 1.504 24.912 1.536 27.42 ;
  LAYER M3 ;
        RECT 1.504 27.368 1.536 27.4 ;
  LAYER M1 ;
        RECT 1.44 24.912 1.472 27.42 ;
  LAYER M3 ;
        RECT 1.44 24.932 1.472 24.964 ;
  LAYER M1 ;
        RECT 1.376 24.912 1.408 27.42 ;
  LAYER M3 ;
        RECT 1.376 27.368 1.408 27.4 ;
  LAYER M1 ;
        RECT 1.312 24.912 1.344 27.42 ;
  LAYER M3 ;
        RECT 1.312 24.932 1.344 24.964 ;
  LAYER M1 ;
        RECT 1.248 24.912 1.28 27.42 ;
  LAYER M3 ;
        RECT 1.248 27.368 1.28 27.4 ;
  LAYER M1 ;
        RECT 1.184 24.912 1.216 27.42 ;
  LAYER M3 ;
        RECT 1.184 24.932 1.216 24.964 ;
  LAYER M1 ;
        RECT 1.12 24.912 1.152 27.42 ;
  LAYER M3 ;
        RECT 1.12 27.368 1.152 27.4 ;
  LAYER M1 ;
        RECT 1.056 24.912 1.088 27.42 ;
  LAYER M3 ;
        RECT 1.056 24.932 1.088 24.964 ;
  LAYER M1 ;
        RECT 0.992 24.912 1.024 27.42 ;
  LAYER M3 ;
        RECT 0.992 27.368 1.024 27.4 ;
  LAYER M1 ;
        RECT 0.928 24.912 0.96 27.42 ;
  LAYER M3 ;
        RECT 0.928 24.932 0.96 24.964 ;
  LAYER M1 ;
        RECT 0.864 24.912 0.896 27.42 ;
  LAYER M3 ;
        RECT 0.864 27.368 0.896 27.4 ;
  LAYER M1 ;
        RECT 0.8 24.912 0.832 27.42 ;
  LAYER M3 ;
        RECT 0.8 24.932 0.832 24.964 ;
  LAYER M1 ;
        RECT 0.736 24.912 0.768 27.42 ;
  LAYER M3 ;
        RECT 0.736 27.368 0.768 27.4 ;
  LAYER M1 ;
        RECT 0.672 24.912 0.704 27.42 ;
  LAYER M3 ;
        RECT 0.672 24.932 0.704 24.964 ;
  LAYER M1 ;
        RECT 0.608 24.912 0.64 27.42 ;
  LAYER M3 ;
        RECT 2.976 27.304 3.008 27.336 ;
  LAYER M2 ;
        RECT 0.608 27.24 0.64 27.272 ;
  LAYER M2 ;
        RECT 2.976 27.176 3.008 27.208 ;
  LAYER M2 ;
        RECT 0.608 27.112 0.64 27.144 ;
  LAYER M2 ;
        RECT 2.976 27.048 3.008 27.08 ;
  LAYER M2 ;
        RECT 0.608 26.984 0.64 27.016 ;
  LAYER M2 ;
        RECT 2.976 26.92 3.008 26.952 ;
  LAYER M2 ;
        RECT 0.608 26.856 0.64 26.888 ;
  LAYER M2 ;
        RECT 2.976 26.792 3.008 26.824 ;
  LAYER M2 ;
        RECT 0.608 26.728 0.64 26.76 ;
  LAYER M2 ;
        RECT 2.976 26.664 3.008 26.696 ;
  LAYER M2 ;
        RECT 0.608 26.6 0.64 26.632 ;
  LAYER M2 ;
        RECT 2.976 26.536 3.008 26.568 ;
  LAYER M2 ;
        RECT 0.608 26.472 0.64 26.504 ;
  LAYER M2 ;
        RECT 2.976 26.408 3.008 26.44 ;
  LAYER M2 ;
        RECT 0.608 26.344 0.64 26.376 ;
  LAYER M2 ;
        RECT 2.976 26.28 3.008 26.312 ;
  LAYER M2 ;
        RECT 0.608 26.216 0.64 26.248 ;
  LAYER M2 ;
        RECT 2.976 26.152 3.008 26.184 ;
  LAYER M2 ;
        RECT 0.608 26.088 0.64 26.12 ;
  LAYER M2 ;
        RECT 2.976 26.024 3.008 26.056 ;
  LAYER M2 ;
        RECT 0.608 25.96 0.64 25.992 ;
  LAYER M2 ;
        RECT 2.976 25.896 3.008 25.928 ;
  LAYER M2 ;
        RECT 0.608 25.832 0.64 25.864 ;
  LAYER M2 ;
        RECT 2.976 25.768 3.008 25.8 ;
  LAYER M2 ;
        RECT 0.608 25.704 0.64 25.736 ;
  LAYER M2 ;
        RECT 2.976 25.64 3.008 25.672 ;
  LAYER M2 ;
        RECT 0.608 25.576 0.64 25.608 ;
  LAYER M2 ;
        RECT 2.976 25.512 3.008 25.544 ;
  LAYER M2 ;
        RECT 0.608 25.448 0.64 25.48 ;
  LAYER M2 ;
        RECT 2.976 25.384 3.008 25.416 ;
  LAYER M2 ;
        RECT 0.608 25.32 0.64 25.352 ;
  LAYER M2 ;
        RECT 2.976 25.256 3.008 25.288 ;
  LAYER M2 ;
        RECT 0.608 25.192 0.64 25.224 ;
  LAYER M2 ;
        RECT 2.976 25.128 3.008 25.16 ;
  LAYER M2 ;
        RECT 0.608 25.064 0.64 25.096 ;
  LAYER M2 ;
        RECT 0.56 24.864 3.056 27.468 ;
  LAYER M1 ;
        RECT 2.976 21.804 3.008 24.312 ;
  LAYER M3 ;
        RECT 2.976 21.824 3.008 21.856 ;
  LAYER M1 ;
        RECT 2.912 21.804 2.944 24.312 ;
  LAYER M3 ;
        RECT 2.912 24.26 2.944 24.292 ;
  LAYER M1 ;
        RECT 2.848 21.804 2.88 24.312 ;
  LAYER M3 ;
        RECT 2.848 21.824 2.88 21.856 ;
  LAYER M1 ;
        RECT 2.784 21.804 2.816 24.312 ;
  LAYER M3 ;
        RECT 2.784 24.26 2.816 24.292 ;
  LAYER M1 ;
        RECT 2.72 21.804 2.752 24.312 ;
  LAYER M3 ;
        RECT 2.72 21.824 2.752 21.856 ;
  LAYER M1 ;
        RECT 2.656 21.804 2.688 24.312 ;
  LAYER M3 ;
        RECT 2.656 24.26 2.688 24.292 ;
  LAYER M1 ;
        RECT 2.592 21.804 2.624 24.312 ;
  LAYER M3 ;
        RECT 2.592 21.824 2.624 21.856 ;
  LAYER M1 ;
        RECT 2.528 21.804 2.56 24.312 ;
  LAYER M3 ;
        RECT 2.528 24.26 2.56 24.292 ;
  LAYER M1 ;
        RECT 2.464 21.804 2.496 24.312 ;
  LAYER M3 ;
        RECT 2.464 21.824 2.496 21.856 ;
  LAYER M1 ;
        RECT 2.4 21.804 2.432 24.312 ;
  LAYER M3 ;
        RECT 2.4 24.26 2.432 24.292 ;
  LAYER M1 ;
        RECT 2.336 21.804 2.368 24.312 ;
  LAYER M3 ;
        RECT 2.336 21.824 2.368 21.856 ;
  LAYER M1 ;
        RECT 2.272 21.804 2.304 24.312 ;
  LAYER M3 ;
        RECT 2.272 24.26 2.304 24.292 ;
  LAYER M1 ;
        RECT 2.208 21.804 2.24 24.312 ;
  LAYER M3 ;
        RECT 2.208 21.824 2.24 21.856 ;
  LAYER M1 ;
        RECT 2.144 21.804 2.176 24.312 ;
  LAYER M3 ;
        RECT 2.144 24.26 2.176 24.292 ;
  LAYER M1 ;
        RECT 2.08 21.804 2.112 24.312 ;
  LAYER M3 ;
        RECT 2.08 21.824 2.112 21.856 ;
  LAYER M1 ;
        RECT 2.016 21.804 2.048 24.312 ;
  LAYER M3 ;
        RECT 2.016 24.26 2.048 24.292 ;
  LAYER M1 ;
        RECT 1.952 21.804 1.984 24.312 ;
  LAYER M3 ;
        RECT 1.952 21.824 1.984 21.856 ;
  LAYER M1 ;
        RECT 1.888 21.804 1.92 24.312 ;
  LAYER M3 ;
        RECT 1.888 24.26 1.92 24.292 ;
  LAYER M1 ;
        RECT 1.824 21.804 1.856 24.312 ;
  LAYER M3 ;
        RECT 1.824 21.824 1.856 21.856 ;
  LAYER M1 ;
        RECT 1.76 21.804 1.792 24.312 ;
  LAYER M3 ;
        RECT 1.76 24.26 1.792 24.292 ;
  LAYER M1 ;
        RECT 1.696 21.804 1.728 24.312 ;
  LAYER M3 ;
        RECT 1.696 21.824 1.728 21.856 ;
  LAYER M1 ;
        RECT 1.632 21.804 1.664 24.312 ;
  LAYER M3 ;
        RECT 1.632 24.26 1.664 24.292 ;
  LAYER M1 ;
        RECT 1.568 21.804 1.6 24.312 ;
  LAYER M3 ;
        RECT 1.568 21.824 1.6 21.856 ;
  LAYER M1 ;
        RECT 1.504 21.804 1.536 24.312 ;
  LAYER M3 ;
        RECT 1.504 24.26 1.536 24.292 ;
  LAYER M1 ;
        RECT 1.44 21.804 1.472 24.312 ;
  LAYER M3 ;
        RECT 1.44 21.824 1.472 21.856 ;
  LAYER M1 ;
        RECT 1.376 21.804 1.408 24.312 ;
  LAYER M3 ;
        RECT 1.376 24.26 1.408 24.292 ;
  LAYER M1 ;
        RECT 1.312 21.804 1.344 24.312 ;
  LAYER M3 ;
        RECT 1.312 21.824 1.344 21.856 ;
  LAYER M1 ;
        RECT 1.248 21.804 1.28 24.312 ;
  LAYER M3 ;
        RECT 1.248 24.26 1.28 24.292 ;
  LAYER M1 ;
        RECT 1.184 21.804 1.216 24.312 ;
  LAYER M3 ;
        RECT 1.184 21.824 1.216 21.856 ;
  LAYER M1 ;
        RECT 1.12 21.804 1.152 24.312 ;
  LAYER M3 ;
        RECT 1.12 24.26 1.152 24.292 ;
  LAYER M1 ;
        RECT 1.056 21.804 1.088 24.312 ;
  LAYER M3 ;
        RECT 1.056 21.824 1.088 21.856 ;
  LAYER M1 ;
        RECT 0.992 21.804 1.024 24.312 ;
  LAYER M3 ;
        RECT 0.992 24.26 1.024 24.292 ;
  LAYER M1 ;
        RECT 0.928 21.804 0.96 24.312 ;
  LAYER M3 ;
        RECT 0.928 21.824 0.96 21.856 ;
  LAYER M1 ;
        RECT 0.864 21.804 0.896 24.312 ;
  LAYER M3 ;
        RECT 0.864 24.26 0.896 24.292 ;
  LAYER M1 ;
        RECT 0.8 21.804 0.832 24.312 ;
  LAYER M3 ;
        RECT 0.8 21.824 0.832 21.856 ;
  LAYER M1 ;
        RECT 0.736 21.804 0.768 24.312 ;
  LAYER M3 ;
        RECT 0.736 24.26 0.768 24.292 ;
  LAYER M1 ;
        RECT 0.672 21.804 0.704 24.312 ;
  LAYER M3 ;
        RECT 0.672 21.824 0.704 21.856 ;
  LAYER M1 ;
        RECT 0.608 21.804 0.64 24.312 ;
  LAYER M3 ;
        RECT 2.976 24.196 3.008 24.228 ;
  LAYER M2 ;
        RECT 0.608 24.132 0.64 24.164 ;
  LAYER M2 ;
        RECT 2.976 24.068 3.008 24.1 ;
  LAYER M2 ;
        RECT 0.608 24.004 0.64 24.036 ;
  LAYER M2 ;
        RECT 2.976 23.94 3.008 23.972 ;
  LAYER M2 ;
        RECT 0.608 23.876 0.64 23.908 ;
  LAYER M2 ;
        RECT 2.976 23.812 3.008 23.844 ;
  LAYER M2 ;
        RECT 0.608 23.748 0.64 23.78 ;
  LAYER M2 ;
        RECT 2.976 23.684 3.008 23.716 ;
  LAYER M2 ;
        RECT 0.608 23.62 0.64 23.652 ;
  LAYER M2 ;
        RECT 2.976 23.556 3.008 23.588 ;
  LAYER M2 ;
        RECT 0.608 23.492 0.64 23.524 ;
  LAYER M2 ;
        RECT 2.976 23.428 3.008 23.46 ;
  LAYER M2 ;
        RECT 0.608 23.364 0.64 23.396 ;
  LAYER M2 ;
        RECT 2.976 23.3 3.008 23.332 ;
  LAYER M2 ;
        RECT 0.608 23.236 0.64 23.268 ;
  LAYER M2 ;
        RECT 2.976 23.172 3.008 23.204 ;
  LAYER M2 ;
        RECT 0.608 23.108 0.64 23.14 ;
  LAYER M2 ;
        RECT 2.976 23.044 3.008 23.076 ;
  LAYER M2 ;
        RECT 0.608 22.98 0.64 23.012 ;
  LAYER M2 ;
        RECT 2.976 22.916 3.008 22.948 ;
  LAYER M2 ;
        RECT 0.608 22.852 0.64 22.884 ;
  LAYER M2 ;
        RECT 2.976 22.788 3.008 22.82 ;
  LAYER M2 ;
        RECT 0.608 22.724 0.64 22.756 ;
  LAYER M2 ;
        RECT 2.976 22.66 3.008 22.692 ;
  LAYER M2 ;
        RECT 0.608 22.596 0.64 22.628 ;
  LAYER M2 ;
        RECT 2.976 22.532 3.008 22.564 ;
  LAYER M2 ;
        RECT 0.608 22.468 0.64 22.5 ;
  LAYER M2 ;
        RECT 2.976 22.404 3.008 22.436 ;
  LAYER M2 ;
        RECT 0.608 22.34 0.64 22.372 ;
  LAYER M2 ;
        RECT 2.976 22.276 3.008 22.308 ;
  LAYER M2 ;
        RECT 0.608 22.212 0.64 22.244 ;
  LAYER M2 ;
        RECT 2.976 22.148 3.008 22.18 ;
  LAYER M2 ;
        RECT 0.608 22.084 0.64 22.116 ;
  LAYER M2 ;
        RECT 2.976 22.02 3.008 22.052 ;
  LAYER M2 ;
        RECT 0.608 21.956 0.64 21.988 ;
  LAYER M2 ;
        RECT 0.56 21.756 3.056 24.36 ;
  LAYER M1 ;
        RECT 2.976 18.696 3.008 21.204 ;
  LAYER M3 ;
        RECT 2.976 18.716 3.008 18.748 ;
  LAYER M1 ;
        RECT 2.912 18.696 2.944 21.204 ;
  LAYER M3 ;
        RECT 2.912 21.152 2.944 21.184 ;
  LAYER M1 ;
        RECT 2.848 18.696 2.88 21.204 ;
  LAYER M3 ;
        RECT 2.848 18.716 2.88 18.748 ;
  LAYER M1 ;
        RECT 2.784 18.696 2.816 21.204 ;
  LAYER M3 ;
        RECT 2.784 21.152 2.816 21.184 ;
  LAYER M1 ;
        RECT 2.72 18.696 2.752 21.204 ;
  LAYER M3 ;
        RECT 2.72 18.716 2.752 18.748 ;
  LAYER M1 ;
        RECT 2.656 18.696 2.688 21.204 ;
  LAYER M3 ;
        RECT 2.656 21.152 2.688 21.184 ;
  LAYER M1 ;
        RECT 2.592 18.696 2.624 21.204 ;
  LAYER M3 ;
        RECT 2.592 18.716 2.624 18.748 ;
  LAYER M1 ;
        RECT 2.528 18.696 2.56 21.204 ;
  LAYER M3 ;
        RECT 2.528 21.152 2.56 21.184 ;
  LAYER M1 ;
        RECT 2.464 18.696 2.496 21.204 ;
  LAYER M3 ;
        RECT 2.464 18.716 2.496 18.748 ;
  LAYER M1 ;
        RECT 2.4 18.696 2.432 21.204 ;
  LAYER M3 ;
        RECT 2.4 21.152 2.432 21.184 ;
  LAYER M1 ;
        RECT 2.336 18.696 2.368 21.204 ;
  LAYER M3 ;
        RECT 2.336 18.716 2.368 18.748 ;
  LAYER M1 ;
        RECT 2.272 18.696 2.304 21.204 ;
  LAYER M3 ;
        RECT 2.272 21.152 2.304 21.184 ;
  LAYER M1 ;
        RECT 2.208 18.696 2.24 21.204 ;
  LAYER M3 ;
        RECT 2.208 18.716 2.24 18.748 ;
  LAYER M1 ;
        RECT 2.144 18.696 2.176 21.204 ;
  LAYER M3 ;
        RECT 2.144 21.152 2.176 21.184 ;
  LAYER M1 ;
        RECT 2.08 18.696 2.112 21.204 ;
  LAYER M3 ;
        RECT 2.08 18.716 2.112 18.748 ;
  LAYER M1 ;
        RECT 2.016 18.696 2.048 21.204 ;
  LAYER M3 ;
        RECT 2.016 21.152 2.048 21.184 ;
  LAYER M1 ;
        RECT 1.952 18.696 1.984 21.204 ;
  LAYER M3 ;
        RECT 1.952 18.716 1.984 18.748 ;
  LAYER M1 ;
        RECT 1.888 18.696 1.92 21.204 ;
  LAYER M3 ;
        RECT 1.888 21.152 1.92 21.184 ;
  LAYER M1 ;
        RECT 1.824 18.696 1.856 21.204 ;
  LAYER M3 ;
        RECT 1.824 18.716 1.856 18.748 ;
  LAYER M1 ;
        RECT 1.76 18.696 1.792 21.204 ;
  LAYER M3 ;
        RECT 1.76 21.152 1.792 21.184 ;
  LAYER M1 ;
        RECT 1.696 18.696 1.728 21.204 ;
  LAYER M3 ;
        RECT 1.696 18.716 1.728 18.748 ;
  LAYER M1 ;
        RECT 1.632 18.696 1.664 21.204 ;
  LAYER M3 ;
        RECT 1.632 21.152 1.664 21.184 ;
  LAYER M1 ;
        RECT 1.568 18.696 1.6 21.204 ;
  LAYER M3 ;
        RECT 1.568 18.716 1.6 18.748 ;
  LAYER M1 ;
        RECT 1.504 18.696 1.536 21.204 ;
  LAYER M3 ;
        RECT 1.504 21.152 1.536 21.184 ;
  LAYER M1 ;
        RECT 1.44 18.696 1.472 21.204 ;
  LAYER M3 ;
        RECT 1.44 18.716 1.472 18.748 ;
  LAYER M1 ;
        RECT 1.376 18.696 1.408 21.204 ;
  LAYER M3 ;
        RECT 1.376 21.152 1.408 21.184 ;
  LAYER M1 ;
        RECT 1.312 18.696 1.344 21.204 ;
  LAYER M3 ;
        RECT 1.312 18.716 1.344 18.748 ;
  LAYER M1 ;
        RECT 1.248 18.696 1.28 21.204 ;
  LAYER M3 ;
        RECT 1.248 21.152 1.28 21.184 ;
  LAYER M1 ;
        RECT 1.184 18.696 1.216 21.204 ;
  LAYER M3 ;
        RECT 1.184 18.716 1.216 18.748 ;
  LAYER M1 ;
        RECT 1.12 18.696 1.152 21.204 ;
  LAYER M3 ;
        RECT 1.12 21.152 1.152 21.184 ;
  LAYER M1 ;
        RECT 1.056 18.696 1.088 21.204 ;
  LAYER M3 ;
        RECT 1.056 18.716 1.088 18.748 ;
  LAYER M1 ;
        RECT 0.992 18.696 1.024 21.204 ;
  LAYER M3 ;
        RECT 0.992 21.152 1.024 21.184 ;
  LAYER M1 ;
        RECT 0.928 18.696 0.96 21.204 ;
  LAYER M3 ;
        RECT 0.928 18.716 0.96 18.748 ;
  LAYER M1 ;
        RECT 0.864 18.696 0.896 21.204 ;
  LAYER M3 ;
        RECT 0.864 21.152 0.896 21.184 ;
  LAYER M1 ;
        RECT 0.8 18.696 0.832 21.204 ;
  LAYER M3 ;
        RECT 0.8 18.716 0.832 18.748 ;
  LAYER M1 ;
        RECT 0.736 18.696 0.768 21.204 ;
  LAYER M3 ;
        RECT 0.736 21.152 0.768 21.184 ;
  LAYER M1 ;
        RECT 0.672 18.696 0.704 21.204 ;
  LAYER M3 ;
        RECT 0.672 18.716 0.704 18.748 ;
  LAYER M1 ;
        RECT 0.608 18.696 0.64 21.204 ;
  LAYER M3 ;
        RECT 2.976 21.088 3.008 21.12 ;
  LAYER M2 ;
        RECT 0.608 21.024 0.64 21.056 ;
  LAYER M2 ;
        RECT 2.976 20.96 3.008 20.992 ;
  LAYER M2 ;
        RECT 0.608 20.896 0.64 20.928 ;
  LAYER M2 ;
        RECT 2.976 20.832 3.008 20.864 ;
  LAYER M2 ;
        RECT 0.608 20.768 0.64 20.8 ;
  LAYER M2 ;
        RECT 2.976 20.704 3.008 20.736 ;
  LAYER M2 ;
        RECT 0.608 20.64 0.64 20.672 ;
  LAYER M2 ;
        RECT 2.976 20.576 3.008 20.608 ;
  LAYER M2 ;
        RECT 0.608 20.512 0.64 20.544 ;
  LAYER M2 ;
        RECT 2.976 20.448 3.008 20.48 ;
  LAYER M2 ;
        RECT 0.608 20.384 0.64 20.416 ;
  LAYER M2 ;
        RECT 2.976 20.32 3.008 20.352 ;
  LAYER M2 ;
        RECT 0.608 20.256 0.64 20.288 ;
  LAYER M2 ;
        RECT 2.976 20.192 3.008 20.224 ;
  LAYER M2 ;
        RECT 0.608 20.128 0.64 20.16 ;
  LAYER M2 ;
        RECT 2.976 20.064 3.008 20.096 ;
  LAYER M2 ;
        RECT 0.608 20 0.64 20.032 ;
  LAYER M2 ;
        RECT 2.976 19.936 3.008 19.968 ;
  LAYER M2 ;
        RECT 0.608 19.872 0.64 19.904 ;
  LAYER M2 ;
        RECT 2.976 19.808 3.008 19.84 ;
  LAYER M2 ;
        RECT 0.608 19.744 0.64 19.776 ;
  LAYER M2 ;
        RECT 2.976 19.68 3.008 19.712 ;
  LAYER M2 ;
        RECT 0.608 19.616 0.64 19.648 ;
  LAYER M2 ;
        RECT 2.976 19.552 3.008 19.584 ;
  LAYER M2 ;
        RECT 0.608 19.488 0.64 19.52 ;
  LAYER M2 ;
        RECT 2.976 19.424 3.008 19.456 ;
  LAYER M2 ;
        RECT 0.608 19.36 0.64 19.392 ;
  LAYER M2 ;
        RECT 2.976 19.296 3.008 19.328 ;
  LAYER M2 ;
        RECT 0.608 19.232 0.64 19.264 ;
  LAYER M2 ;
        RECT 2.976 19.168 3.008 19.2 ;
  LAYER M2 ;
        RECT 0.608 19.104 0.64 19.136 ;
  LAYER M2 ;
        RECT 2.976 19.04 3.008 19.072 ;
  LAYER M2 ;
        RECT 0.608 18.976 0.64 19.008 ;
  LAYER M2 ;
        RECT 2.976 18.912 3.008 18.944 ;
  LAYER M2 ;
        RECT 0.608 18.848 0.64 18.88 ;
  LAYER M2 ;
        RECT 0.56 18.648 3.056 21.252 ;
  LAYER M1 ;
        RECT 2.976 15.588 3.008 18.096 ;
  LAYER M3 ;
        RECT 2.976 15.608 3.008 15.64 ;
  LAYER M1 ;
        RECT 2.912 15.588 2.944 18.096 ;
  LAYER M3 ;
        RECT 2.912 18.044 2.944 18.076 ;
  LAYER M1 ;
        RECT 2.848 15.588 2.88 18.096 ;
  LAYER M3 ;
        RECT 2.848 15.608 2.88 15.64 ;
  LAYER M1 ;
        RECT 2.784 15.588 2.816 18.096 ;
  LAYER M3 ;
        RECT 2.784 18.044 2.816 18.076 ;
  LAYER M1 ;
        RECT 2.72 15.588 2.752 18.096 ;
  LAYER M3 ;
        RECT 2.72 15.608 2.752 15.64 ;
  LAYER M1 ;
        RECT 2.656 15.588 2.688 18.096 ;
  LAYER M3 ;
        RECT 2.656 18.044 2.688 18.076 ;
  LAYER M1 ;
        RECT 2.592 15.588 2.624 18.096 ;
  LAYER M3 ;
        RECT 2.592 15.608 2.624 15.64 ;
  LAYER M1 ;
        RECT 2.528 15.588 2.56 18.096 ;
  LAYER M3 ;
        RECT 2.528 18.044 2.56 18.076 ;
  LAYER M1 ;
        RECT 2.464 15.588 2.496 18.096 ;
  LAYER M3 ;
        RECT 2.464 15.608 2.496 15.64 ;
  LAYER M1 ;
        RECT 2.4 15.588 2.432 18.096 ;
  LAYER M3 ;
        RECT 2.4 18.044 2.432 18.076 ;
  LAYER M1 ;
        RECT 2.336 15.588 2.368 18.096 ;
  LAYER M3 ;
        RECT 2.336 15.608 2.368 15.64 ;
  LAYER M1 ;
        RECT 2.272 15.588 2.304 18.096 ;
  LAYER M3 ;
        RECT 2.272 18.044 2.304 18.076 ;
  LAYER M1 ;
        RECT 2.208 15.588 2.24 18.096 ;
  LAYER M3 ;
        RECT 2.208 15.608 2.24 15.64 ;
  LAYER M1 ;
        RECT 2.144 15.588 2.176 18.096 ;
  LAYER M3 ;
        RECT 2.144 18.044 2.176 18.076 ;
  LAYER M1 ;
        RECT 2.08 15.588 2.112 18.096 ;
  LAYER M3 ;
        RECT 2.08 15.608 2.112 15.64 ;
  LAYER M1 ;
        RECT 2.016 15.588 2.048 18.096 ;
  LAYER M3 ;
        RECT 2.016 18.044 2.048 18.076 ;
  LAYER M1 ;
        RECT 1.952 15.588 1.984 18.096 ;
  LAYER M3 ;
        RECT 1.952 15.608 1.984 15.64 ;
  LAYER M1 ;
        RECT 1.888 15.588 1.92 18.096 ;
  LAYER M3 ;
        RECT 1.888 18.044 1.92 18.076 ;
  LAYER M1 ;
        RECT 1.824 15.588 1.856 18.096 ;
  LAYER M3 ;
        RECT 1.824 15.608 1.856 15.64 ;
  LAYER M1 ;
        RECT 1.76 15.588 1.792 18.096 ;
  LAYER M3 ;
        RECT 1.76 18.044 1.792 18.076 ;
  LAYER M1 ;
        RECT 1.696 15.588 1.728 18.096 ;
  LAYER M3 ;
        RECT 1.696 15.608 1.728 15.64 ;
  LAYER M1 ;
        RECT 1.632 15.588 1.664 18.096 ;
  LAYER M3 ;
        RECT 1.632 18.044 1.664 18.076 ;
  LAYER M1 ;
        RECT 1.568 15.588 1.6 18.096 ;
  LAYER M3 ;
        RECT 1.568 15.608 1.6 15.64 ;
  LAYER M1 ;
        RECT 1.504 15.588 1.536 18.096 ;
  LAYER M3 ;
        RECT 1.504 18.044 1.536 18.076 ;
  LAYER M1 ;
        RECT 1.44 15.588 1.472 18.096 ;
  LAYER M3 ;
        RECT 1.44 15.608 1.472 15.64 ;
  LAYER M1 ;
        RECT 1.376 15.588 1.408 18.096 ;
  LAYER M3 ;
        RECT 1.376 18.044 1.408 18.076 ;
  LAYER M1 ;
        RECT 1.312 15.588 1.344 18.096 ;
  LAYER M3 ;
        RECT 1.312 15.608 1.344 15.64 ;
  LAYER M1 ;
        RECT 1.248 15.588 1.28 18.096 ;
  LAYER M3 ;
        RECT 1.248 18.044 1.28 18.076 ;
  LAYER M1 ;
        RECT 1.184 15.588 1.216 18.096 ;
  LAYER M3 ;
        RECT 1.184 15.608 1.216 15.64 ;
  LAYER M1 ;
        RECT 1.12 15.588 1.152 18.096 ;
  LAYER M3 ;
        RECT 1.12 18.044 1.152 18.076 ;
  LAYER M1 ;
        RECT 1.056 15.588 1.088 18.096 ;
  LAYER M3 ;
        RECT 1.056 15.608 1.088 15.64 ;
  LAYER M1 ;
        RECT 0.992 15.588 1.024 18.096 ;
  LAYER M3 ;
        RECT 0.992 18.044 1.024 18.076 ;
  LAYER M1 ;
        RECT 0.928 15.588 0.96 18.096 ;
  LAYER M3 ;
        RECT 0.928 15.608 0.96 15.64 ;
  LAYER M1 ;
        RECT 0.864 15.588 0.896 18.096 ;
  LAYER M3 ;
        RECT 0.864 18.044 0.896 18.076 ;
  LAYER M1 ;
        RECT 0.8 15.588 0.832 18.096 ;
  LAYER M3 ;
        RECT 0.8 15.608 0.832 15.64 ;
  LAYER M1 ;
        RECT 0.736 15.588 0.768 18.096 ;
  LAYER M3 ;
        RECT 0.736 18.044 0.768 18.076 ;
  LAYER M1 ;
        RECT 0.672 15.588 0.704 18.096 ;
  LAYER M3 ;
        RECT 0.672 15.608 0.704 15.64 ;
  LAYER M1 ;
        RECT 0.608 15.588 0.64 18.096 ;
  LAYER M3 ;
        RECT 2.976 17.98 3.008 18.012 ;
  LAYER M2 ;
        RECT 0.608 17.916 0.64 17.948 ;
  LAYER M2 ;
        RECT 2.976 17.852 3.008 17.884 ;
  LAYER M2 ;
        RECT 0.608 17.788 0.64 17.82 ;
  LAYER M2 ;
        RECT 2.976 17.724 3.008 17.756 ;
  LAYER M2 ;
        RECT 0.608 17.66 0.64 17.692 ;
  LAYER M2 ;
        RECT 2.976 17.596 3.008 17.628 ;
  LAYER M2 ;
        RECT 0.608 17.532 0.64 17.564 ;
  LAYER M2 ;
        RECT 2.976 17.468 3.008 17.5 ;
  LAYER M2 ;
        RECT 0.608 17.404 0.64 17.436 ;
  LAYER M2 ;
        RECT 2.976 17.34 3.008 17.372 ;
  LAYER M2 ;
        RECT 0.608 17.276 0.64 17.308 ;
  LAYER M2 ;
        RECT 2.976 17.212 3.008 17.244 ;
  LAYER M2 ;
        RECT 0.608 17.148 0.64 17.18 ;
  LAYER M2 ;
        RECT 2.976 17.084 3.008 17.116 ;
  LAYER M2 ;
        RECT 0.608 17.02 0.64 17.052 ;
  LAYER M2 ;
        RECT 2.976 16.956 3.008 16.988 ;
  LAYER M2 ;
        RECT 0.608 16.892 0.64 16.924 ;
  LAYER M2 ;
        RECT 2.976 16.828 3.008 16.86 ;
  LAYER M2 ;
        RECT 0.608 16.764 0.64 16.796 ;
  LAYER M2 ;
        RECT 2.976 16.7 3.008 16.732 ;
  LAYER M2 ;
        RECT 0.608 16.636 0.64 16.668 ;
  LAYER M2 ;
        RECT 2.976 16.572 3.008 16.604 ;
  LAYER M2 ;
        RECT 0.608 16.508 0.64 16.54 ;
  LAYER M2 ;
        RECT 2.976 16.444 3.008 16.476 ;
  LAYER M2 ;
        RECT 0.608 16.38 0.64 16.412 ;
  LAYER M2 ;
        RECT 2.976 16.316 3.008 16.348 ;
  LAYER M2 ;
        RECT 0.608 16.252 0.64 16.284 ;
  LAYER M2 ;
        RECT 2.976 16.188 3.008 16.22 ;
  LAYER M2 ;
        RECT 0.608 16.124 0.64 16.156 ;
  LAYER M2 ;
        RECT 2.976 16.06 3.008 16.092 ;
  LAYER M2 ;
        RECT 0.608 15.996 0.64 16.028 ;
  LAYER M2 ;
        RECT 2.976 15.932 3.008 15.964 ;
  LAYER M2 ;
        RECT 0.608 15.868 0.64 15.9 ;
  LAYER M2 ;
        RECT 2.976 15.804 3.008 15.836 ;
  LAYER M2 ;
        RECT 0.608 15.74 0.64 15.772 ;
  LAYER M2 ;
        RECT 0.56 15.54 3.056 18.144 ;
  LAYER M1 ;
        RECT 41.072 14.244 41.104 14.316 ;
  LAYER M2 ;
        RECT 41.052 14.264 41.124 14.296 ;
  LAYER M1 ;
        RECT 38.096 14.244 38.128 14.316 ;
  LAYER M2 ;
        RECT 38.076 14.264 38.148 14.296 ;
  LAYER M2 ;
        RECT 38.112 14.264 41.088 14.296 ;
  LAYER M2 ;
        RECT 40.684 0.908 41.396 0.94 ;
  LAYER M1 ;
        RECT 38.176 31.044 38.208 31.116 ;
  LAYER M2 ;
        RECT 38.156 31.064 38.228 31.096 ;
  LAYER M1 ;
        RECT 41.152 31.044 41.184 31.116 ;
  LAYER M2 ;
        RECT 41.132 31.064 41.204 31.096 ;
  LAYER M2 ;
        RECT 38.192 31.064 41.168 31.096 ;
  LAYER M2 ;
        RECT 40.944 14.264 40.976 14.296 ;
  LAYER M3 ;
        RECT 40.94 0.924 40.98 14.28 ;
  LAYER M2 ;
        RECT 40.944 0.908 40.976 0.94 ;
  LAYER M2 ;
        RECT 38.624 14.264 38.656 14.296 ;
  LAYER M3 ;
        RECT 38.62 14.28 38.66 17.808 ;
  LAYER M4 ;
        RECT 38.62 17.788 38.66 17.828 ;
  LAYER M5 ;
        RECT 38.608 17.808 38.672 31.08 ;
  LAYER M4 ;
        RECT 38.62 31.06 38.66 31.1 ;
  LAYER M3 ;
        RECT 38.62 31.06 38.66 31.1 ;
  LAYER M2 ;
        RECT 38.624 31.064 38.656 31.096 ;
  LAYER M1 ;
        RECT 41.232 1.308 41.264 1.38 ;
  LAYER M2 ;
        RECT 41.212 1.328 41.284 1.36 ;
  LAYER M1 ;
        RECT 38.256 1.308 38.288 1.38 ;
  LAYER M2 ;
        RECT 38.236 1.328 38.308 1.36 ;
  LAYER M2 ;
        RECT 38.272 1.328 41.248 1.36 ;
  LAYER M2 ;
        RECT 42.044 0.32 42.116 0.352 ;
  LAYER M2 ;
        RECT 31.884 0.32 31.956 0.352 ;
  LAYER M2 ;
        RECT 41.28 1.328 41.76 1.36 ;
  LAYER M3 ;
        RECT 41.74 0.336 41.78 1.344 ;
  LAYER M4 ;
        RECT 41.76 0.316 42.08 0.356 ;
  LAYER M3 ;
        RECT 42.06 0.316 42.1 0.356 ;
  LAYER M2 ;
        RECT 42.064 0.32 42.096 0.352 ;
  LAYER M2 ;
        RECT 32.24 1.328 38.24 1.36 ;
  LAYER M3 ;
        RECT 32.22 0.336 32.26 1.344 ;
  LAYER M4 ;
        RECT 31.92 0.316 32.24 0.356 ;
  LAYER M3 ;
        RECT 31.9 0.316 31.94 0.356 ;
  LAYER M2 ;
        RECT 31.904 0.32 31.936 0.352 ;
  LAYER M2 ;
        RECT 39.324 0.908 40.036 0.94 ;
  LAYER M1 ;
        RECT 38.336 15 38.368 15.072 ;
  LAYER M2 ;
        RECT 38.316 15.02 38.388 15.052 ;
  LAYER M1 ;
        RECT 41.312 15 41.344 15.072 ;
  LAYER M2 ;
        RECT 41.292 15.02 41.364 15.052 ;
  LAYER M2 ;
        RECT 38.352 15.02 41.328 15.052 ;
  LAYER M2 ;
        RECT 39.984 0.908 40.016 0.94 ;
  LAYER M3 ;
        RECT 39.98 0.924 40.02 15.036 ;
  LAYER M2 ;
        RECT 39.984 15.02 40.016 15.052 ;
  LAYER M1 ;
        RECT 38.48 5.004 38.512 5.076 ;
  LAYER M2 ;
        RECT 38.46 5.024 38.532 5.056 ;
  LAYER M2 ;
        RECT 38.496 5.024 41.248 5.056 ;
  LAYER M1 ;
        RECT 41.232 5.004 41.264 5.076 ;
  LAYER M2 ;
        RECT 41.212 5.024 41.284 5.056 ;
  LAYER M1 ;
        RECT 38.48 8.112 38.512 8.184 ;
  LAYER M2 ;
        RECT 38.46 8.132 38.532 8.164 ;
  LAYER M2 ;
        RECT 38.496 8.132 41.248 8.164 ;
  LAYER M1 ;
        RECT 41.232 8.112 41.264 8.184 ;
  LAYER M2 ;
        RECT 41.212 8.132 41.284 8.164 ;
  LAYER M1 ;
        RECT 41.456 5.004 41.488 5.076 ;
  LAYER M2 ;
        RECT 41.436 5.024 41.508 5.056 ;
  LAYER M1 ;
        RECT 41.456 4.872 41.488 5.04 ;
  LAYER M1 ;
        RECT 41.456 4.836 41.488 4.908 ;
  LAYER M2 ;
        RECT 41.436 4.856 41.508 4.888 ;
  LAYER M2 ;
        RECT 41.248 4.856 41.472 4.888 ;
  LAYER M1 ;
        RECT 41.232 4.836 41.264 4.908 ;
  LAYER M2 ;
        RECT 41.212 4.856 41.284 4.888 ;
  LAYER M1 ;
        RECT 41.456 8.112 41.488 8.184 ;
  LAYER M2 ;
        RECT 41.436 8.132 41.508 8.164 ;
  LAYER M1 ;
        RECT 41.456 7.98 41.488 8.148 ;
  LAYER M1 ;
        RECT 41.456 7.944 41.488 8.016 ;
  LAYER M2 ;
        RECT 41.436 7.964 41.508 7.996 ;
  LAYER M2 ;
        RECT 41.248 7.964 41.472 7.996 ;
  LAYER M1 ;
        RECT 41.232 7.944 41.264 8.016 ;
  LAYER M2 ;
        RECT 41.212 7.964 41.284 7.996 ;
  LAYER M1 ;
        RECT 41.232 1.308 41.264 1.38 ;
  LAYER M2 ;
        RECT 41.212 1.328 41.284 1.36 ;
  LAYER M1 ;
        RECT 41.232 1.344 41.264 1.596 ;
  LAYER M1 ;
        RECT 41.232 1.596 41.264 8.148 ;
  LAYER M1 ;
        RECT 35.504 8.112 35.536 8.184 ;
  LAYER M2 ;
        RECT 35.484 8.132 35.556 8.164 ;
  LAYER M2 ;
        RECT 35.52 8.132 38.272 8.164 ;
  LAYER M1 ;
        RECT 38.256 8.112 38.288 8.184 ;
  LAYER M2 ;
        RECT 38.236 8.132 38.308 8.164 ;
  LAYER M1 ;
        RECT 35.504 5.004 35.536 5.076 ;
  LAYER M2 ;
        RECT 35.484 5.024 35.556 5.056 ;
  LAYER M2 ;
        RECT 35.52 5.024 38.272 5.056 ;
  LAYER M1 ;
        RECT 38.256 5.004 38.288 5.076 ;
  LAYER M2 ;
        RECT 38.236 5.024 38.308 5.056 ;
  LAYER M1 ;
        RECT 38.256 1.308 38.288 1.38 ;
  LAYER M2 ;
        RECT 38.236 1.328 38.308 1.36 ;
  LAYER M1 ;
        RECT 38.256 1.344 38.288 1.596 ;
  LAYER M1 ;
        RECT 38.256 1.596 38.288 8.148 ;
  LAYER M2 ;
        RECT 38.272 1.328 41.248 1.36 ;
  LAYER M1 ;
        RECT 44.432 1.896 44.464 1.968 ;
  LAYER M2 ;
        RECT 44.412 1.916 44.484 1.948 ;
  LAYER M1 ;
        RECT 44.432 1.764 44.464 1.932 ;
  LAYER M1 ;
        RECT 44.432 1.728 44.464 1.8 ;
  LAYER M2 ;
        RECT 44.412 1.748 44.484 1.78 ;
  LAYER M2 ;
        RECT 44.224 1.748 44.448 1.78 ;
  LAYER M1 ;
        RECT 44.208 1.728 44.24 1.8 ;
  LAYER M2 ;
        RECT 44.188 1.748 44.26 1.78 ;
  LAYER M1 ;
        RECT 44.432 5.004 44.464 5.076 ;
  LAYER M2 ;
        RECT 44.412 5.024 44.484 5.056 ;
  LAYER M1 ;
        RECT 44.432 4.872 44.464 5.04 ;
  LAYER M1 ;
        RECT 44.432 4.836 44.464 4.908 ;
  LAYER M2 ;
        RECT 44.412 4.856 44.484 4.888 ;
  LAYER M2 ;
        RECT 44.224 4.856 44.448 4.888 ;
  LAYER M1 ;
        RECT 44.208 4.836 44.24 4.908 ;
  LAYER M2 ;
        RECT 44.188 4.856 44.26 4.888 ;
  LAYER M1 ;
        RECT 44.432 8.112 44.464 8.184 ;
  LAYER M2 ;
        RECT 44.412 8.132 44.484 8.164 ;
  LAYER M1 ;
        RECT 44.432 7.98 44.464 8.148 ;
  LAYER M1 ;
        RECT 44.432 7.944 44.464 8.016 ;
  LAYER M2 ;
        RECT 44.412 7.964 44.484 7.996 ;
  LAYER M2 ;
        RECT 44.224 7.964 44.448 7.996 ;
  LAYER M1 ;
        RECT 44.208 7.944 44.24 8.016 ;
  LAYER M2 ;
        RECT 44.188 7.964 44.26 7.996 ;
  LAYER M1 ;
        RECT 44.432 11.22 44.464 11.292 ;
  LAYER M2 ;
        RECT 44.412 11.24 44.484 11.272 ;
  LAYER M1 ;
        RECT 44.432 11.088 44.464 11.256 ;
  LAYER M1 ;
        RECT 44.432 11.052 44.464 11.124 ;
  LAYER M2 ;
        RECT 44.412 11.072 44.484 11.104 ;
  LAYER M2 ;
        RECT 44.224 11.072 44.448 11.104 ;
  LAYER M1 ;
        RECT 44.208 11.052 44.24 11.124 ;
  LAYER M2 ;
        RECT 44.188 11.072 44.26 11.104 ;
  LAYER M1 ;
        RECT 41.456 1.896 41.488 1.968 ;
  LAYER M2 ;
        RECT 41.436 1.916 41.508 1.948 ;
  LAYER M2 ;
        RECT 41.472 1.916 44.224 1.948 ;
  LAYER M1 ;
        RECT 44.208 1.896 44.24 1.968 ;
  LAYER M2 ;
        RECT 44.188 1.916 44.26 1.948 ;
  LAYER M1 ;
        RECT 41.456 11.22 41.488 11.292 ;
  LAYER M2 ;
        RECT 41.436 11.24 41.508 11.272 ;
  LAYER M2 ;
        RECT 41.472 11.24 44.224 11.272 ;
  LAYER M1 ;
        RECT 44.208 11.22 44.24 11.292 ;
  LAYER M2 ;
        RECT 44.188 11.24 44.26 11.272 ;
  LAYER M1 ;
        RECT 44.208 1.14 44.24 1.212 ;
  LAYER M2 ;
        RECT 44.188 1.16 44.26 1.192 ;
  LAYER M1 ;
        RECT 44.208 1.176 44.24 1.596 ;
  LAYER M1 ;
        RECT 44.208 1.596 44.24 11.256 ;
  LAYER M1 ;
        RECT 35.504 1.896 35.536 1.968 ;
  LAYER M2 ;
        RECT 35.484 1.916 35.556 1.948 ;
  LAYER M1 ;
        RECT 35.504 1.764 35.536 1.932 ;
  LAYER M1 ;
        RECT 35.504 1.728 35.536 1.8 ;
  LAYER M2 ;
        RECT 35.484 1.748 35.556 1.78 ;
  LAYER M2 ;
        RECT 35.296 1.748 35.52 1.78 ;
  LAYER M1 ;
        RECT 35.28 1.728 35.312 1.8 ;
  LAYER M2 ;
        RECT 35.26 1.748 35.332 1.78 ;
  LAYER M1 ;
        RECT 35.504 11.22 35.536 11.292 ;
  LAYER M2 ;
        RECT 35.484 11.24 35.556 11.272 ;
  LAYER M1 ;
        RECT 35.504 11.088 35.536 11.256 ;
  LAYER M1 ;
        RECT 35.504 11.052 35.536 11.124 ;
  LAYER M2 ;
        RECT 35.484 11.072 35.556 11.104 ;
  LAYER M2 ;
        RECT 35.296 11.072 35.52 11.104 ;
  LAYER M1 ;
        RECT 35.28 11.052 35.312 11.124 ;
  LAYER M2 ;
        RECT 35.26 11.072 35.332 11.104 ;
  LAYER M1 ;
        RECT 32.528 1.896 32.56 1.968 ;
  LAYER M2 ;
        RECT 32.508 1.916 32.58 1.948 ;
  LAYER M2 ;
        RECT 32.544 1.916 35.296 1.948 ;
  LAYER M1 ;
        RECT 35.28 1.896 35.312 1.968 ;
  LAYER M2 ;
        RECT 35.26 1.916 35.332 1.948 ;
  LAYER M1 ;
        RECT 32.528 5.004 32.56 5.076 ;
  LAYER M2 ;
        RECT 32.508 5.024 32.58 5.056 ;
  LAYER M2 ;
        RECT 32.544 5.024 35.296 5.056 ;
  LAYER M1 ;
        RECT 35.28 5.004 35.312 5.076 ;
  LAYER M2 ;
        RECT 35.26 5.024 35.332 5.056 ;
  LAYER M1 ;
        RECT 32.528 8.112 32.56 8.184 ;
  LAYER M2 ;
        RECT 32.508 8.132 32.58 8.164 ;
  LAYER M2 ;
        RECT 32.544 8.132 35.296 8.164 ;
  LAYER M1 ;
        RECT 35.28 8.112 35.312 8.184 ;
  LAYER M2 ;
        RECT 35.26 8.132 35.332 8.164 ;
  LAYER M1 ;
        RECT 32.528 11.22 32.56 11.292 ;
  LAYER M2 ;
        RECT 32.508 11.24 32.58 11.272 ;
  LAYER M2 ;
        RECT 32.544 11.24 35.296 11.272 ;
  LAYER M1 ;
        RECT 35.28 11.22 35.312 11.292 ;
  LAYER M2 ;
        RECT 35.26 11.24 35.332 11.272 ;
  LAYER M1 ;
        RECT 35.28 1.14 35.312 1.212 ;
  LAYER M2 ;
        RECT 35.26 1.16 35.332 1.192 ;
  LAYER M1 ;
        RECT 35.28 1.176 35.312 1.596 ;
  LAYER M1 ;
        RECT 35.28 1.596 35.312 11.256 ;
  LAYER M2 ;
        RECT 35.296 1.16 44.224 1.192 ;
  LAYER M1 ;
        RECT 38.48 11.22 38.512 11.292 ;
  LAYER M2 ;
        RECT 38.46 11.24 38.532 11.272 ;
  LAYER M2 ;
        RECT 38.496 11.24 41.472 11.272 ;
  LAYER M1 ;
        RECT 41.456 11.22 41.488 11.292 ;
  LAYER M2 ;
        RECT 41.436 11.24 41.508 11.272 ;
  LAYER M1 ;
        RECT 38.48 1.896 38.512 1.968 ;
  LAYER M2 ;
        RECT 38.46 1.916 38.532 1.948 ;
  LAYER M2 ;
        RECT 35.52 1.916 38.496 1.948 ;
  LAYER M1 ;
        RECT 35.504 1.896 35.536 1.968 ;
  LAYER M2 ;
        RECT 35.484 1.916 35.556 1.948 ;
  LAYER M1 ;
        RECT 40.848 7.44 40.88 7.512 ;
  LAYER M2 ;
        RECT 40.828 7.46 40.9 7.492 ;
  LAYER M2 ;
        RECT 40.864 7.46 41.088 7.492 ;
  LAYER M1 ;
        RECT 41.072 7.44 41.104 7.512 ;
  LAYER M2 ;
        RECT 41.052 7.46 41.124 7.492 ;
  LAYER M1 ;
        RECT 40.848 10.548 40.88 10.62 ;
  LAYER M2 ;
        RECT 40.828 10.568 40.9 10.6 ;
  LAYER M2 ;
        RECT 40.864 10.568 41.088 10.6 ;
  LAYER M1 ;
        RECT 41.072 10.548 41.104 10.62 ;
  LAYER M2 ;
        RECT 41.052 10.568 41.124 10.6 ;
  LAYER M1 ;
        RECT 43.824 7.44 43.856 7.512 ;
  LAYER M2 ;
        RECT 43.804 7.46 43.876 7.492 ;
  LAYER M1 ;
        RECT 43.824 7.476 43.856 7.644 ;
  LAYER M1 ;
        RECT 43.824 7.608 43.856 7.68 ;
  LAYER M2 ;
        RECT 43.804 7.628 43.876 7.66 ;
  LAYER M2 ;
        RECT 41.088 7.628 43.84 7.66 ;
  LAYER M1 ;
        RECT 41.072 7.608 41.104 7.68 ;
  LAYER M2 ;
        RECT 41.052 7.628 41.124 7.66 ;
  LAYER M1 ;
        RECT 43.824 10.548 43.856 10.62 ;
  LAYER M2 ;
        RECT 43.804 10.568 43.876 10.6 ;
  LAYER M1 ;
        RECT 43.824 10.584 43.856 10.752 ;
  LAYER M1 ;
        RECT 43.824 10.716 43.856 10.788 ;
  LAYER M2 ;
        RECT 43.804 10.736 43.876 10.768 ;
  LAYER M2 ;
        RECT 41.088 10.736 43.84 10.768 ;
  LAYER M1 ;
        RECT 41.072 10.716 41.104 10.788 ;
  LAYER M2 ;
        RECT 41.052 10.736 41.124 10.768 ;
  LAYER M1 ;
        RECT 41.072 14.244 41.104 14.316 ;
  LAYER M2 ;
        RECT 41.052 14.264 41.124 14.296 ;
  LAYER M1 ;
        RECT 41.072 14.028 41.104 14.28 ;
  LAYER M1 ;
        RECT 41.072 7.476 41.104 14.028 ;
  LAYER M1 ;
        RECT 37.872 10.548 37.904 10.62 ;
  LAYER M2 ;
        RECT 37.852 10.568 37.924 10.6 ;
  LAYER M2 ;
        RECT 37.888 10.568 38.112 10.6 ;
  LAYER M1 ;
        RECT 38.096 10.548 38.128 10.62 ;
  LAYER M2 ;
        RECT 38.076 10.568 38.148 10.6 ;
  LAYER M1 ;
        RECT 37.872 7.44 37.904 7.512 ;
  LAYER M2 ;
        RECT 37.852 7.46 37.924 7.492 ;
  LAYER M2 ;
        RECT 37.888 7.46 38.112 7.492 ;
  LAYER M1 ;
        RECT 38.096 7.44 38.128 7.512 ;
  LAYER M2 ;
        RECT 38.076 7.46 38.148 7.492 ;
  LAYER M1 ;
        RECT 38.096 14.244 38.128 14.316 ;
  LAYER M2 ;
        RECT 38.076 14.264 38.148 14.296 ;
  LAYER M1 ;
        RECT 38.096 14.028 38.128 14.28 ;
  LAYER M1 ;
        RECT 38.096 7.476 38.128 14.028 ;
  LAYER M2 ;
        RECT 38.112 14.264 41.088 14.296 ;
  LAYER M1 ;
        RECT 46.8 4.332 46.832 4.404 ;
  LAYER M2 ;
        RECT 46.78 4.352 46.852 4.384 ;
  LAYER M2 ;
        RECT 46.816 4.352 47.2 4.384 ;
  LAYER M1 ;
        RECT 47.184 4.332 47.216 4.404 ;
  LAYER M2 ;
        RECT 47.164 4.352 47.236 4.384 ;
  LAYER M1 ;
        RECT 46.8 7.44 46.832 7.512 ;
  LAYER M2 ;
        RECT 46.78 7.46 46.852 7.492 ;
  LAYER M2 ;
        RECT 46.816 7.46 47.2 7.492 ;
  LAYER M1 ;
        RECT 47.184 7.44 47.216 7.512 ;
  LAYER M2 ;
        RECT 47.164 7.46 47.236 7.492 ;
  LAYER M1 ;
        RECT 46.8 10.548 46.832 10.62 ;
  LAYER M2 ;
        RECT 46.78 10.568 46.852 10.6 ;
  LAYER M2 ;
        RECT 46.816 10.568 47.2 10.6 ;
  LAYER M1 ;
        RECT 47.184 10.548 47.216 10.62 ;
  LAYER M2 ;
        RECT 47.164 10.568 47.236 10.6 ;
  LAYER M1 ;
        RECT 46.8 13.656 46.832 13.728 ;
  LAYER M2 ;
        RECT 46.78 13.676 46.852 13.708 ;
  LAYER M2 ;
        RECT 46.816 13.676 47.2 13.708 ;
  LAYER M1 ;
        RECT 47.184 13.656 47.216 13.728 ;
  LAYER M2 ;
        RECT 47.164 13.676 47.236 13.708 ;
  LAYER M1 ;
        RECT 47.184 14.412 47.216 14.484 ;
  LAYER M2 ;
        RECT 47.164 14.432 47.236 14.464 ;
  LAYER M1 ;
        RECT 47.184 14.028 47.216 14.448 ;
  LAYER M1 ;
        RECT 47.184 4.368 47.216 14.028 ;
  LAYER M1 ;
        RECT 34.896 4.332 34.928 4.404 ;
  LAYER M2 ;
        RECT 34.876 4.352 34.948 4.384 ;
  LAYER M1 ;
        RECT 34.896 4.368 34.928 4.536 ;
  LAYER M1 ;
        RECT 34.896 4.5 34.928 4.572 ;
  LAYER M2 ;
        RECT 34.876 4.52 34.948 4.552 ;
  LAYER M2 ;
        RECT 32.32 4.52 34.912 4.552 ;
  LAYER M1 ;
        RECT 32.304 4.5 32.336 4.572 ;
  LAYER M2 ;
        RECT 32.284 4.52 32.356 4.552 ;
  LAYER M1 ;
        RECT 34.896 7.44 34.928 7.512 ;
  LAYER M2 ;
        RECT 34.876 7.46 34.948 7.492 ;
  LAYER M1 ;
        RECT 34.896 7.476 34.928 7.644 ;
  LAYER M1 ;
        RECT 34.896 7.608 34.928 7.68 ;
  LAYER M2 ;
        RECT 34.876 7.628 34.948 7.66 ;
  LAYER M2 ;
        RECT 32.32 7.628 34.912 7.66 ;
  LAYER M1 ;
        RECT 32.304 7.608 32.336 7.68 ;
  LAYER M2 ;
        RECT 32.284 7.628 32.356 7.66 ;
  LAYER M1 ;
        RECT 34.896 10.548 34.928 10.62 ;
  LAYER M2 ;
        RECT 34.876 10.568 34.948 10.6 ;
  LAYER M1 ;
        RECT 34.896 10.584 34.928 10.752 ;
  LAYER M1 ;
        RECT 34.896 10.716 34.928 10.788 ;
  LAYER M2 ;
        RECT 34.876 10.736 34.948 10.768 ;
  LAYER M2 ;
        RECT 32.32 10.736 34.912 10.768 ;
  LAYER M1 ;
        RECT 32.304 10.716 32.336 10.788 ;
  LAYER M2 ;
        RECT 32.284 10.736 32.356 10.768 ;
  LAYER M1 ;
        RECT 34.896 13.656 34.928 13.728 ;
  LAYER M2 ;
        RECT 34.876 13.676 34.948 13.708 ;
  LAYER M1 ;
        RECT 34.896 13.692 34.928 13.86 ;
  LAYER M1 ;
        RECT 34.896 13.824 34.928 13.896 ;
  LAYER M2 ;
        RECT 34.876 13.844 34.948 13.876 ;
  LAYER M2 ;
        RECT 32.32 13.844 34.912 13.876 ;
  LAYER M1 ;
        RECT 32.304 13.824 32.336 13.896 ;
  LAYER M2 ;
        RECT 32.284 13.844 32.356 13.876 ;
  LAYER M1 ;
        RECT 32.304 14.412 32.336 14.484 ;
  LAYER M2 ;
        RECT 32.284 14.432 32.356 14.464 ;
  LAYER M1 ;
        RECT 32.304 14.028 32.336 14.448 ;
  LAYER M1 ;
        RECT 32.304 4.536 32.336 14.028 ;
  LAYER M2 ;
        RECT 32.32 14.432 47.2 14.464 ;
  LAYER M1 ;
        RECT 43.824 4.332 43.856 4.404 ;
  LAYER M2 ;
        RECT 43.804 4.352 43.876 4.384 ;
  LAYER M2 ;
        RECT 43.84 4.352 46.816 4.384 ;
  LAYER M1 ;
        RECT 46.8 4.332 46.832 4.404 ;
  LAYER M2 ;
        RECT 46.78 4.352 46.852 4.384 ;
  LAYER M1 ;
        RECT 43.824 13.656 43.856 13.728 ;
  LAYER M2 ;
        RECT 43.804 13.676 43.876 13.708 ;
  LAYER M2 ;
        RECT 43.84 13.676 46.816 13.708 ;
  LAYER M1 ;
        RECT 46.8 13.656 46.832 13.728 ;
  LAYER M2 ;
        RECT 46.78 13.676 46.852 13.708 ;
  LAYER M1 ;
        RECT 40.848 13.656 40.88 13.728 ;
  LAYER M2 ;
        RECT 40.828 13.676 40.9 13.708 ;
  LAYER M2 ;
        RECT 40.864 13.676 43.84 13.708 ;
  LAYER M1 ;
        RECT 43.824 13.656 43.856 13.728 ;
  LAYER M2 ;
        RECT 43.804 13.676 43.876 13.708 ;
  LAYER M1 ;
        RECT 37.872 13.656 37.904 13.728 ;
  LAYER M2 ;
        RECT 37.852 13.676 37.924 13.708 ;
  LAYER M2 ;
        RECT 37.888 13.676 40.864 13.708 ;
  LAYER M1 ;
        RECT 40.848 13.656 40.88 13.728 ;
  LAYER M2 ;
        RECT 40.828 13.676 40.9 13.708 ;
  LAYER M1 ;
        RECT 37.872 4.332 37.904 4.404 ;
  LAYER M2 ;
        RECT 37.852 4.352 37.924 4.384 ;
  LAYER M2 ;
        RECT 34.912 4.352 37.888 4.384 ;
  LAYER M1 ;
        RECT 34.896 4.332 34.928 4.404 ;
  LAYER M2 ;
        RECT 34.876 4.352 34.948 4.384 ;
  LAYER M1 ;
        RECT 40.848 4.332 40.88 4.404 ;
  LAYER M2 ;
        RECT 40.828 4.352 40.9 4.384 ;
  LAYER M2 ;
        RECT 37.888 4.352 40.864 4.384 ;
  LAYER M1 ;
        RECT 37.872 4.332 37.904 4.404 ;
  LAYER M2 ;
        RECT 37.852 4.352 37.924 4.384 ;
  LAYER M1 ;
        RECT 46.8 1.896 46.832 4.404 ;
  LAYER M3 ;
        RECT 46.8 4.352 46.832 4.384 ;
  LAYER M1 ;
        RECT 46.736 1.896 46.768 4.404 ;
  LAYER M3 ;
        RECT 46.736 1.916 46.768 1.948 ;
  LAYER M1 ;
        RECT 46.672 1.896 46.704 4.404 ;
  LAYER M3 ;
        RECT 46.672 4.352 46.704 4.384 ;
  LAYER M1 ;
        RECT 46.608 1.896 46.64 4.404 ;
  LAYER M3 ;
        RECT 46.608 1.916 46.64 1.948 ;
  LAYER M1 ;
        RECT 46.544 1.896 46.576 4.404 ;
  LAYER M3 ;
        RECT 46.544 4.352 46.576 4.384 ;
  LAYER M1 ;
        RECT 46.48 1.896 46.512 4.404 ;
  LAYER M3 ;
        RECT 46.48 1.916 46.512 1.948 ;
  LAYER M1 ;
        RECT 46.416 1.896 46.448 4.404 ;
  LAYER M3 ;
        RECT 46.416 4.352 46.448 4.384 ;
  LAYER M1 ;
        RECT 46.352 1.896 46.384 4.404 ;
  LAYER M3 ;
        RECT 46.352 1.916 46.384 1.948 ;
  LAYER M1 ;
        RECT 46.288 1.896 46.32 4.404 ;
  LAYER M3 ;
        RECT 46.288 4.352 46.32 4.384 ;
  LAYER M1 ;
        RECT 46.224 1.896 46.256 4.404 ;
  LAYER M3 ;
        RECT 46.224 1.916 46.256 1.948 ;
  LAYER M1 ;
        RECT 46.16 1.896 46.192 4.404 ;
  LAYER M3 ;
        RECT 46.16 4.352 46.192 4.384 ;
  LAYER M1 ;
        RECT 46.096 1.896 46.128 4.404 ;
  LAYER M3 ;
        RECT 46.096 1.916 46.128 1.948 ;
  LAYER M1 ;
        RECT 46.032 1.896 46.064 4.404 ;
  LAYER M3 ;
        RECT 46.032 4.352 46.064 4.384 ;
  LAYER M1 ;
        RECT 45.968 1.896 46 4.404 ;
  LAYER M3 ;
        RECT 45.968 1.916 46 1.948 ;
  LAYER M1 ;
        RECT 45.904 1.896 45.936 4.404 ;
  LAYER M3 ;
        RECT 45.904 4.352 45.936 4.384 ;
  LAYER M1 ;
        RECT 45.84 1.896 45.872 4.404 ;
  LAYER M3 ;
        RECT 45.84 1.916 45.872 1.948 ;
  LAYER M1 ;
        RECT 45.776 1.896 45.808 4.404 ;
  LAYER M3 ;
        RECT 45.776 4.352 45.808 4.384 ;
  LAYER M1 ;
        RECT 45.712 1.896 45.744 4.404 ;
  LAYER M3 ;
        RECT 45.712 1.916 45.744 1.948 ;
  LAYER M1 ;
        RECT 45.648 1.896 45.68 4.404 ;
  LAYER M3 ;
        RECT 45.648 4.352 45.68 4.384 ;
  LAYER M1 ;
        RECT 45.584 1.896 45.616 4.404 ;
  LAYER M3 ;
        RECT 45.584 1.916 45.616 1.948 ;
  LAYER M1 ;
        RECT 45.52 1.896 45.552 4.404 ;
  LAYER M3 ;
        RECT 45.52 4.352 45.552 4.384 ;
  LAYER M1 ;
        RECT 45.456 1.896 45.488 4.404 ;
  LAYER M3 ;
        RECT 45.456 1.916 45.488 1.948 ;
  LAYER M1 ;
        RECT 45.392 1.896 45.424 4.404 ;
  LAYER M3 ;
        RECT 45.392 4.352 45.424 4.384 ;
  LAYER M1 ;
        RECT 45.328 1.896 45.36 4.404 ;
  LAYER M3 ;
        RECT 45.328 1.916 45.36 1.948 ;
  LAYER M1 ;
        RECT 45.264 1.896 45.296 4.404 ;
  LAYER M3 ;
        RECT 45.264 4.352 45.296 4.384 ;
  LAYER M1 ;
        RECT 45.2 1.896 45.232 4.404 ;
  LAYER M3 ;
        RECT 45.2 1.916 45.232 1.948 ;
  LAYER M1 ;
        RECT 45.136 1.896 45.168 4.404 ;
  LAYER M3 ;
        RECT 45.136 4.352 45.168 4.384 ;
  LAYER M1 ;
        RECT 45.072 1.896 45.104 4.404 ;
  LAYER M3 ;
        RECT 45.072 1.916 45.104 1.948 ;
  LAYER M1 ;
        RECT 45.008 1.896 45.04 4.404 ;
  LAYER M3 ;
        RECT 45.008 4.352 45.04 4.384 ;
  LAYER M1 ;
        RECT 44.944 1.896 44.976 4.404 ;
  LAYER M3 ;
        RECT 44.944 1.916 44.976 1.948 ;
  LAYER M1 ;
        RECT 44.88 1.896 44.912 4.404 ;
  LAYER M3 ;
        RECT 44.88 4.352 44.912 4.384 ;
  LAYER M1 ;
        RECT 44.816 1.896 44.848 4.404 ;
  LAYER M3 ;
        RECT 44.816 1.916 44.848 1.948 ;
  LAYER M1 ;
        RECT 44.752 1.896 44.784 4.404 ;
  LAYER M3 ;
        RECT 44.752 4.352 44.784 4.384 ;
  LAYER M1 ;
        RECT 44.688 1.896 44.72 4.404 ;
  LAYER M3 ;
        RECT 44.688 1.916 44.72 1.948 ;
  LAYER M1 ;
        RECT 44.624 1.896 44.656 4.404 ;
  LAYER M3 ;
        RECT 44.624 4.352 44.656 4.384 ;
  LAYER M1 ;
        RECT 44.56 1.896 44.592 4.404 ;
  LAYER M3 ;
        RECT 44.56 1.916 44.592 1.948 ;
  LAYER M1 ;
        RECT 44.496 1.896 44.528 4.404 ;
  LAYER M3 ;
        RECT 44.496 4.352 44.528 4.384 ;
  LAYER M1 ;
        RECT 44.432 1.896 44.464 4.404 ;
  LAYER M3 ;
        RECT 46.8 1.98 46.832 2.012 ;
  LAYER M2 ;
        RECT 44.432 2.044 44.464 2.076 ;
  LAYER M2 ;
        RECT 46.8 2.108 46.832 2.14 ;
  LAYER M2 ;
        RECT 44.432 2.172 44.464 2.204 ;
  LAYER M2 ;
        RECT 46.8 2.236 46.832 2.268 ;
  LAYER M2 ;
        RECT 44.432 2.3 44.464 2.332 ;
  LAYER M2 ;
        RECT 46.8 2.364 46.832 2.396 ;
  LAYER M2 ;
        RECT 44.432 2.428 44.464 2.46 ;
  LAYER M2 ;
        RECT 46.8 2.492 46.832 2.524 ;
  LAYER M2 ;
        RECT 44.432 2.556 44.464 2.588 ;
  LAYER M2 ;
        RECT 46.8 2.62 46.832 2.652 ;
  LAYER M2 ;
        RECT 44.432 2.684 44.464 2.716 ;
  LAYER M2 ;
        RECT 46.8 2.748 46.832 2.78 ;
  LAYER M2 ;
        RECT 44.432 2.812 44.464 2.844 ;
  LAYER M2 ;
        RECT 46.8 2.876 46.832 2.908 ;
  LAYER M2 ;
        RECT 44.432 2.94 44.464 2.972 ;
  LAYER M2 ;
        RECT 46.8 3.004 46.832 3.036 ;
  LAYER M2 ;
        RECT 44.432 3.068 44.464 3.1 ;
  LAYER M2 ;
        RECT 46.8 3.132 46.832 3.164 ;
  LAYER M2 ;
        RECT 44.432 3.196 44.464 3.228 ;
  LAYER M2 ;
        RECT 46.8 3.26 46.832 3.292 ;
  LAYER M2 ;
        RECT 44.432 3.324 44.464 3.356 ;
  LAYER M2 ;
        RECT 46.8 3.388 46.832 3.42 ;
  LAYER M2 ;
        RECT 44.432 3.452 44.464 3.484 ;
  LAYER M2 ;
        RECT 46.8 3.516 46.832 3.548 ;
  LAYER M2 ;
        RECT 44.432 3.58 44.464 3.612 ;
  LAYER M2 ;
        RECT 46.8 3.644 46.832 3.676 ;
  LAYER M2 ;
        RECT 44.432 3.708 44.464 3.74 ;
  LAYER M2 ;
        RECT 46.8 3.772 46.832 3.804 ;
  LAYER M2 ;
        RECT 44.432 3.836 44.464 3.868 ;
  LAYER M2 ;
        RECT 46.8 3.9 46.832 3.932 ;
  LAYER M2 ;
        RECT 44.432 3.964 44.464 3.996 ;
  LAYER M2 ;
        RECT 46.8 4.028 46.832 4.06 ;
  LAYER M2 ;
        RECT 44.432 4.092 44.464 4.124 ;
  LAYER M2 ;
        RECT 46.8 4.156 46.832 4.188 ;
  LAYER M2 ;
        RECT 44.432 4.22 44.464 4.252 ;
  LAYER M2 ;
        RECT 44.384 1.848 46.88 4.452 ;
  LAYER M1 ;
        RECT 46.8 5.004 46.832 7.512 ;
  LAYER M3 ;
        RECT 46.8 7.46 46.832 7.492 ;
  LAYER M1 ;
        RECT 46.736 5.004 46.768 7.512 ;
  LAYER M3 ;
        RECT 46.736 5.024 46.768 5.056 ;
  LAYER M1 ;
        RECT 46.672 5.004 46.704 7.512 ;
  LAYER M3 ;
        RECT 46.672 7.46 46.704 7.492 ;
  LAYER M1 ;
        RECT 46.608 5.004 46.64 7.512 ;
  LAYER M3 ;
        RECT 46.608 5.024 46.64 5.056 ;
  LAYER M1 ;
        RECT 46.544 5.004 46.576 7.512 ;
  LAYER M3 ;
        RECT 46.544 7.46 46.576 7.492 ;
  LAYER M1 ;
        RECT 46.48 5.004 46.512 7.512 ;
  LAYER M3 ;
        RECT 46.48 5.024 46.512 5.056 ;
  LAYER M1 ;
        RECT 46.416 5.004 46.448 7.512 ;
  LAYER M3 ;
        RECT 46.416 7.46 46.448 7.492 ;
  LAYER M1 ;
        RECT 46.352 5.004 46.384 7.512 ;
  LAYER M3 ;
        RECT 46.352 5.024 46.384 5.056 ;
  LAYER M1 ;
        RECT 46.288 5.004 46.32 7.512 ;
  LAYER M3 ;
        RECT 46.288 7.46 46.32 7.492 ;
  LAYER M1 ;
        RECT 46.224 5.004 46.256 7.512 ;
  LAYER M3 ;
        RECT 46.224 5.024 46.256 5.056 ;
  LAYER M1 ;
        RECT 46.16 5.004 46.192 7.512 ;
  LAYER M3 ;
        RECT 46.16 7.46 46.192 7.492 ;
  LAYER M1 ;
        RECT 46.096 5.004 46.128 7.512 ;
  LAYER M3 ;
        RECT 46.096 5.024 46.128 5.056 ;
  LAYER M1 ;
        RECT 46.032 5.004 46.064 7.512 ;
  LAYER M3 ;
        RECT 46.032 7.46 46.064 7.492 ;
  LAYER M1 ;
        RECT 45.968 5.004 46 7.512 ;
  LAYER M3 ;
        RECT 45.968 5.024 46 5.056 ;
  LAYER M1 ;
        RECT 45.904 5.004 45.936 7.512 ;
  LAYER M3 ;
        RECT 45.904 7.46 45.936 7.492 ;
  LAYER M1 ;
        RECT 45.84 5.004 45.872 7.512 ;
  LAYER M3 ;
        RECT 45.84 5.024 45.872 5.056 ;
  LAYER M1 ;
        RECT 45.776 5.004 45.808 7.512 ;
  LAYER M3 ;
        RECT 45.776 7.46 45.808 7.492 ;
  LAYER M1 ;
        RECT 45.712 5.004 45.744 7.512 ;
  LAYER M3 ;
        RECT 45.712 5.024 45.744 5.056 ;
  LAYER M1 ;
        RECT 45.648 5.004 45.68 7.512 ;
  LAYER M3 ;
        RECT 45.648 7.46 45.68 7.492 ;
  LAYER M1 ;
        RECT 45.584 5.004 45.616 7.512 ;
  LAYER M3 ;
        RECT 45.584 5.024 45.616 5.056 ;
  LAYER M1 ;
        RECT 45.52 5.004 45.552 7.512 ;
  LAYER M3 ;
        RECT 45.52 7.46 45.552 7.492 ;
  LAYER M1 ;
        RECT 45.456 5.004 45.488 7.512 ;
  LAYER M3 ;
        RECT 45.456 5.024 45.488 5.056 ;
  LAYER M1 ;
        RECT 45.392 5.004 45.424 7.512 ;
  LAYER M3 ;
        RECT 45.392 7.46 45.424 7.492 ;
  LAYER M1 ;
        RECT 45.328 5.004 45.36 7.512 ;
  LAYER M3 ;
        RECT 45.328 5.024 45.36 5.056 ;
  LAYER M1 ;
        RECT 45.264 5.004 45.296 7.512 ;
  LAYER M3 ;
        RECT 45.264 7.46 45.296 7.492 ;
  LAYER M1 ;
        RECT 45.2 5.004 45.232 7.512 ;
  LAYER M3 ;
        RECT 45.2 5.024 45.232 5.056 ;
  LAYER M1 ;
        RECT 45.136 5.004 45.168 7.512 ;
  LAYER M3 ;
        RECT 45.136 7.46 45.168 7.492 ;
  LAYER M1 ;
        RECT 45.072 5.004 45.104 7.512 ;
  LAYER M3 ;
        RECT 45.072 5.024 45.104 5.056 ;
  LAYER M1 ;
        RECT 45.008 5.004 45.04 7.512 ;
  LAYER M3 ;
        RECT 45.008 7.46 45.04 7.492 ;
  LAYER M1 ;
        RECT 44.944 5.004 44.976 7.512 ;
  LAYER M3 ;
        RECT 44.944 5.024 44.976 5.056 ;
  LAYER M1 ;
        RECT 44.88 5.004 44.912 7.512 ;
  LAYER M3 ;
        RECT 44.88 7.46 44.912 7.492 ;
  LAYER M1 ;
        RECT 44.816 5.004 44.848 7.512 ;
  LAYER M3 ;
        RECT 44.816 5.024 44.848 5.056 ;
  LAYER M1 ;
        RECT 44.752 5.004 44.784 7.512 ;
  LAYER M3 ;
        RECT 44.752 7.46 44.784 7.492 ;
  LAYER M1 ;
        RECT 44.688 5.004 44.72 7.512 ;
  LAYER M3 ;
        RECT 44.688 5.024 44.72 5.056 ;
  LAYER M1 ;
        RECT 44.624 5.004 44.656 7.512 ;
  LAYER M3 ;
        RECT 44.624 7.46 44.656 7.492 ;
  LAYER M1 ;
        RECT 44.56 5.004 44.592 7.512 ;
  LAYER M3 ;
        RECT 44.56 5.024 44.592 5.056 ;
  LAYER M1 ;
        RECT 44.496 5.004 44.528 7.512 ;
  LAYER M3 ;
        RECT 44.496 7.46 44.528 7.492 ;
  LAYER M1 ;
        RECT 44.432 5.004 44.464 7.512 ;
  LAYER M3 ;
        RECT 46.8 5.088 46.832 5.12 ;
  LAYER M2 ;
        RECT 44.432 5.152 44.464 5.184 ;
  LAYER M2 ;
        RECT 46.8 5.216 46.832 5.248 ;
  LAYER M2 ;
        RECT 44.432 5.28 44.464 5.312 ;
  LAYER M2 ;
        RECT 46.8 5.344 46.832 5.376 ;
  LAYER M2 ;
        RECT 44.432 5.408 44.464 5.44 ;
  LAYER M2 ;
        RECT 46.8 5.472 46.832 5.504 ;
  LAYER M2 ;
        RECT 44.432 5.536 44.464 5.568 ;
  LAYER M2 ;
        RECT 46.8 5.6 46.832 5.632 ;
  LAYER M2 ;
        RECT 44.432 5.664 44.464 5.696 ;
  LAYER M2 ;
        RECT 46.8 5.728 46.832 5.76 ;
  LAYER M2 ;
        RECT 44.432 5.792 44.464 5.824 ;
  LAYER M2 ;
        RECT 46.8 5.856 46.832 5.888 ;
  LAYER M2 ;
        RECT 44.432 5.92 44.464 5.952 ;
  LAYER M2 ;
        RECT 46.8 5.984 46.832 6.016 ;
  LAYER M2 ;
        RECT 44.432 6.048 44.464 6.08 ;
  LAYER M2 ;
        RECT 46.8 6.112 46.832 6.144 ;
  LAYER M2 ;
        RECT 44.432 6.176 44.464 6.208 ;
  LAYER M2 ;
        RECT 46.8 6.24 46.832 6.272 ;
  LAYER M2 ;
        RECT 44.432 6.304 44.464 6.336 ;
  LAYER M2 ;
        RECT 46.8 6.368 46.832 6.4 ;
  LAYER M2 ;
        RECT 44.432 6.432 44.464 6.464 ;
  LAYER M2 ;
        RECT 46.8 6.496 46.832 6.528 ;
  LAYER M2 ;
        RECT 44.432 6.56 44.464 6.592 ;
  LAYER M2 ;
        RECT 46.8 6.624 46.832 6.656 ;
  LAYER M2 ;
        RECT 44.432 6.688 44.464 6.72 ;
  LAYER M2 ;
        RECT 46.8 6.752 46.832 6.784 ;
  LAYER M2 ;
        RECT 44.432 6.816 44.464 6.848 ;
  LAYER M2 ;
        RECT 46.8 6.88 46.832 6.912 ;
  LAYER M2 ;
        RECT 44.432 6.944 44.464 6.976 ;
  LAYER M2 ;
        RECT 46.8 7.008 46.832 7.04 ;
  LAYER M2 ;
        RECT 44.432 7.072 44.464 7.104 ;
  LAYER M2 ;
        RECT 46.8 7.136 46.832 7.168 ;
  LAYER M2 ;
        RECT 44.432 7.2 44.464 7.232 ;
  LAYER M2 ;
        RECT 46.8 7.264 46.832 7.296 ;
  LAYER M2 ;
        RECT 44.432 7.328 44.464 7.36 ;
  LAYER M2 ;
        RECT 44.384 4.956 46.88 7.56 ;
  LAYER M1 ;
        RECT 46.8 8.112 46.832 10.62 ;
  LAYER M3 ;
        RECT 46.8 10.568 46.832 10.6 ;
  LAYER M1 ;
        RECT 46.736 8.112 46.768 10.62 ;
  LAYER M3 ;
        RECT 46.736 8.132 46.768 8.164 ;
  LAYER M1 ;
        RECT 46.672 8.112 46.704 10.62 ;
  LAYER M3 ;
        RECT 46.672 10.568 46.704 10.6 ;
  LAYER M1 ;
        RECT 46.608 8.112 46.64 10.62 ;
  LAYER M3 ;
        RECT 46.608 8.132 46.64 8.164 ;
  LAYER M1 ;
        RECT 46.544 8.112 46.576 10.62 ;
  LAYER M3 ;
        RECT 46.544 10.568 46.576 10.6 ;
  LAYER M1 ;
        RECT 46.48 8.112 46.512 10.62 ;
  LAYER M3 ;
        RECT 46.48 8.132 46.512 8.164 ;
  LAYER M1 ;
        RECT 46.416 8.112 46.448 10.62 ;
  LAYER M3 ;
        RECT 46.416 10.568 46.448 10.6 ;
  LAYER M1 ;
        RECT 46.352 8.112 46.384 10.62 ;
  LAYER M3 ;
        RECT 46.352 8.132 46.384 8.164 ;
  LAYER M1 ;
        RECT 46.288 8.112 46.32 10.62 ;
  LAYER M3 ;
        RECT 46.288 10.568 46.32 10.6 ;
  LAYER M1 ;
        RECT 46.224 8.112 46.256 10.62 ;
  LAYER M3 ;
        RECT 46.224 8.132 46.256 8.164 ;
  LAYER M1 ;
        RECT 46.16 8.112 46.192 10.62 ;
  LAYER M3 ;
        RECT 46.16 10.568 46.192 10.6 ;
  LAYER M1 ;
        RECT 46.096 8.112 46.128 10.62 ;
  LAYER M3 ;
        RECT 46.096 8.132 46.128 8.164 ;
  LAYER M1 ;
        RECT 46.032 8.112 46.064 10.62 ;
  LAYER M3 ;
        RECT 46.032 10.568 46.064 10.6 ;
  LAYER M1 ;
        RECT 45.968 8.112 46 10.62 ;
  LAYER M3 ;
        RECT 45.968 8.132 46 8.164 ;
  LAYER M1 ;
        RECT 45.904 8.112 45.936 10.62 ;
  LAYER M3 ;
        RECT 45.904 10.568 45.936 10.6 ;
  LAYER M1 ;
        RECT 45.84 8.112 45.872 10.62 ;
  LAYER M3 ;
        RECT 45.84 8.132 45.872 8.164 ;
  LAYER M1 ;
        RECT 45.776 8.112 45.808 10.62 ;
  LAYER M3 ;
        RECT 45.776 10.568 45.808 10.6 ;
  LAYER M1 ;
        RECT 45.712 8.112 45.744 10.62 ;
  LAYER M3 ;
        RECT 45.712 8.132 45.744 8.164 ;
  LAYER M1 ;
        RECT 45.648 8.112 45.68 10.62 ;
  LAYER M3 ;
        RECT 45.648 10.568 45.68 10.6 ;
  LAYER M1 ;
        RECT 45.584 8.112 45.616 10.62 ;
  LAYER M3 ;
        RECT 45.584 8.132 45.616 8.164 ;
  LAYER M1 ;
        RECT 45.52 8.112 45.552 10.62 ;
  LAYER M3 ;
        RECT 45.52 10.568 45.552 10.6 ;
  LAYER M1 ;
        RECT 45.456 8.112 45.488 10.62 ;
  LAYER M3 ;
        RECT 45.456 8.132 45.488 8.164 ;
  LAYER M1 ;
        RECT 45.392 8.112 45.424 10.62 ;
  LAYER M3 ;
        RECT 45.392 10.568 45.424 10.6 ;
  LAYER M1 ;
        RECT 45.328 8.112 45.36 10.62 ;
  LAYER M3 ;
        RECT 45.328 8.132 45.36 8.164 ;
  LAYER M1 ;
        RECT 45.264 8.112 45.296 10.62 ;
  LAYER M3 ;
        RECT 45.264 10.568 45.296 10.6 ;
  LAYER M1 ;
        RECT 45.2 8.112 45.232 10.62 ;
  LAYER M3 ;
        RECT 45.2 8.132 45.232 8.164 ;
  LAYER M1 ;
        RECT 45.136 8.112 45.168 10.62 ;
  LAYER M3 ;
        RECT 45.136 10.568 45.168 10.6 ;
  LAYER M1 ;
        RECT 45.072 8.112 45.104 10.62 ;
  LAYER M3 ;
        RECT 45.072 8.132 45.104 8.164 ;
  LAYER M1 ;
        RECT 45.008 8.112 45.04 10.62 ;
  LAYER M3 ;
        RECT 45.008 10.568 45.04 10.6 ;
  LAYER M1 ;
        RECT 44.944 8.112 44.976 10.62 ;
  LAYER M3 ;
        RECT 44.944 8.132 44.976 8.164 ;
  LAYER M1 ;
        RECT 44.88 8.112 44.912 10.62 ;
  LAYER M3 ;
        RECT 44.88 10.568 44.912 10.6 ;
  LAYER M1 ;
        RECT 44.816 8.112 44.848 10.62 ;
  LAYER M3 ;
        RECT 44.816 8.132 44.848 8.164 ;
  LAYER M1 ;
        RECT 44.752 8.112 44.784 10.62 ;
  LAYER M3 ;
        RECT 44.752 10.568 44.784 10.6 ;
  LAYER M1 ;
        RECT 44.688 8.112 44.72 10.62 ;
  LAYER M3 ;
        RECT 44.688 8.132 44.72 8.164 ;
  LAYER M1 ;
        RECT 44.624 8.112 44.656 10.62 ;
  LAYER M3 ;
        RECT 44.624 10.568 44.656 10.6 ;
  LAYER M1 ;
        RECT 44.56 8.112 44.592 10.62 ;
  LAYER M3 ;
        RECT 44.56 8.132 44.592 8.164 ;
  LAYER M1 ;
        RECT 44.496 8.112 44.528 10.62 ;
  LAYER M3 ;
        RECT 44.496 10.568 44.528 10.6 ;
  LAYER M1 ;
        RECT 44.432 8.112 44.464 10.62 ;
  LAYER M3 ;
        RECT 46.8 8.196 46.832 8.228 ;
  LAYER M2 ;
        RECT 44.432 8.26 44.464 8.292 ;
  LAYER M2 ;
        RECT 46.8 8.324 46.832 8.356 ;
  LAYER M2 ;
        RECT 44.432 8.388 44.464 8.42 ;
  LAYER M2 ;
        RECT 46.8 8.452 46.832 8.484 ;
  LAYER M2 ;
        RECT 44.432 8.516 44.464 8.548 ;
  LAYER M2 ;
        RECT 46.8 8.58 46.832 8.612 ;
  LAYER M2 ;
        RECT 44.432 8.644 44.464 8.676 ;
  LAYER M2 ;
        RECT 46.8 8.708 46.832 8.74 ;
  LAYER M2 ;
        RECT 44.432 8.772 44.464 8.804 ;
  LAYER M2 ;
        RECT 46.8 8.836 46.832 8.868 ;
  LAYER M2 ;
        RECT 44.432 8.9 44.464 8.932 ;
  LAYER M2 ;
        RECT 46.8 8.964 46.832 8.996 ;
  LAYER M2 ;
        RECT 44.432 9.028 44.464 9.06 ;
  LAYER M2 ;
        RECT 46.8 9.092 46.832 9.124 ;
  LAYER M2 ;
        RECT 44.432 9.156 44.464 9.188 ;
  LAYER M2 ;
        RECT 46.8 9.22 46.832 9.252 ;
  LAYER M2 ;
        RECT 44.432 9.284 44.464 9.316 ;
  LAYER M2 ;
        RECT 46.8 9.348 46.832 9.38 ;
  LAYER M2 ;
        RECT 44.432 9.412 44.464 9.444 ;
  LAYER M2 ;
        RECT 46.8 9.476 46.832 9.508 ;
  LAYER M2 ;
        RECT 44.432 9.54 44.464 9.572 ;
  LAYER M2 ;
        RECT 46.8 9.604 46.832 9.636 ;
  LAYER M2 ;
        RECT 44.432 9.668 44.464 9.7 ;
  LAYER M2 ;
        RECT 46.8 9.732 46.832 9.764 ;
  LAYER M2 ;
        RECT 44.432 9.796 44.464 9.828 ;
  LAYER M2 ;
        RECT 46.8 9.86 46.832 9.892 ;
  LAYER M2 ;
        RECT 44.432 9.924 44.464 9.956 ;
  LAYER M2 ;
        RECT 46.8 9.988 46.832 10.02 ;
  LAYER M2 ;
        RECT 44.432 10.052 44.464 10.084 ;
  LAYER M2 ;
        RECT 46.8 10.116 46.832 10.148 ;
  LAYER M2 ;
        RECT 44.432 10.18 44.464 10.212 ;
  LAYER M2 ;
        RECT 46.8 10.244 46.832 10.276 ;
  LAYER M2 ;
        RECT 44.432 10.308 44.464 10.34 ;
  LAYER M2 ;
        RECT 46.8 10.372 46.832 10.404 ;
  LAYER M2 ;
        RECT 44.432 10.436 44.464 10.468 ;
  LAYER M2 ;
        RECT 44.384 8.064 46.88 10.668 ;
  LAYER M1 ;
        RECT 46.8 11.22 46.832 13.728 ;
  LAYER M3 ;
        RECT 46.8 13.676 46.832 13.708 ;
  LAYER M1 ;
        RECT 46.736 11.22 46.768 13.728 ;
  LAYER M3 ;
        RECT 46.736 11.24 46.768 11.272 ;
  LAYER M1 ;
        RECT 46.672 11.22 46.704 13.728 ;
  LAYER M3 ;
        RECT 46.672 13.676 46.704 13.708 ;
  LAYER M1 ;
        RECT 46.608 11.22 46.64 13.728 ;
  LAYER M3 ;
        RECT 46.608 11.24 46.64 11.272 ;
  LAYER M1 ;
        RECT 46.544 11.22 46.576 13.728 ;
  LAYER M3 ;
        RECT 46.544 13.676 46.576 13.708 ;
  LAYER M1 ;
        RECT 46.48 11.22 46.512 13.728 ;
  LAYER M3 ;
        RECT 46.48 11.24 46.512 11.272 ;
  LAYER M1 ;
        RECT 46.416 11.22 46.448 13.728 ;
  LAYER M3 ;
        RECT 46.416 13.676 46.448 13.708 ;
  LAYER M1 ;
        RECT 46.352 11.22 46.384 13.728 ;
  LAYER M3 ;
        RECT 46.352 11.24 46.384 11.272 ;
  LAYER M1 ;
        RECT 46.288 11.22 46.32 13.728 ;
  LAYER M3 ;
        RECT 46.288 13.676 46.32 13.708 ;
  LAYER M1 ;
        RECT 46.224 11.22 46.256 13.728 ;
  LAYER M3 ;
        RECT 46.224 11.24 46.256 11.272 ;
  LAYER M1 ;
        RECT 46.16 11.22 46.192 13.728 ;
  LAYER M3 ;
        RECT 46.16 13.676 46.192 13.708 ;
  LAYER M1 ;
        RECT 46.096 11.22 46.128 13.728 ;
  LAYER M3 ;
        RECT 46.096 11.24 46.128 11.272 ;
  LAYER M1 ;
        RECT 46.032 11.22 46.064 13.728 ;
  LAYER M3 ;
        RECT 46.032 13.676 46.064 13.708 ;
  LAYER M1 ;
        RECT 45.968 11.22 46 13.728 ;
  LAYER M3 ;
        RECT 45.968 11.24 46 11.272 ;
  LAYER M1 ;
        RECT 45.904 11.22 45.936 13.728 ;
  LAYER M3 ;
        RECT 45.904 13.676 45.936 13.708 ;
  LAYER M1 ;
        RECT 45.84 11.22 45.872 13.728 ;
  LAYER M3 ;
        RECT 45.84 11.24 45.872 11.272 ;
  LAYER M1 ;
        RECT 45.776 11.22 45.808 13.728 ;
  LAYER M3 ;
        RECT 45.776 13.676 45.808 13.708 ;
  LAYER M1 ;
        RECT 45.712 11.22 45.744 13.728 ;
  LAYER M3 ;
        RECT 45.712 11.24 45.744 11.272 ;
  LAYER M1 ;
        RECT 45.648 11.22 45.68 13.728 ;
  LAYER M3 ;
        RECT 45.648 13.676 45.68 13.708 ;
  LAYER M1 ;
        RECT 45.584 11.22 45.616 13.728 ;
  LAYER M3 ;
        RECT 45.584 11.24 45.616 11.272 ;
  LAYER M1 ;
        RECT 45.52 11.22 45.552 13.728 ;
  LAYER M3 ;
        RECT 45.52 13.676 45.552 13.708 ;
  LAYER M1 ;
        RECT 45.456 11.22 45.488 13.728 ;
  LAYER M3 ;
        RECT 45.456 11.24 45.488 11.272 ;
  LAYER M1 ;
        RECT 45.392 11.22 45.424 13.728 ;
  LAYER M3 ;
        RECT 45.392 13.676 45.424 13.708 ;
  LAYER M1 ;
        RECT 45.328 11.22 45.36 13.728 ;
  LAYER M3 ;
        RECT 45.328 11.24 45.36 11.272 ;
  LAYER M1 ;
        RECT 45.264 11.22 45.296 13.728 ;
  LAYER M3 ;
        RECT 45.264 13.676 45.296 13.708 ;
  LAYER M1 ;
        RECT 45.2 11.22 45.232 13.728 ;
  LAYER M3 ;
        RECT 45.2 11.24 45.232 11.272 ;
  LAYER M1 ;
        RECT 45.136 11.22 45.168 13.728 ;
  LAYER M3 ;
        RECT 45.136 13.676 45.168 13.708 ;
  LAYER M1 ;
        RECT 45.072 11.22 45.104 13.728 ;
  LAYER M3 ;
        RECT 45.072 11.24 45.104 11.272 ;
  LAYER M1 ;
        RECT 45.008 11.22 45.04 13.728 ;
  LAYER M3 ;
        RECT 45.008 13.676 45.04 13.708 ;
  LAYER M1 ;
        RECT 44.944 11.22 44.976 13.728 ;
  LAYER M3 ;
        RECT 44.944 11.24 44.976 11.272 ;
  LAYER M1 ;
        RECT 44.88 11.22 44.912 13.728 ;
  LAYER M3 ;
        RECT 44.88 13.676 44.912 13.708 ;
  LAYER M1 ;
        RECT 44.816 11.22 44.848 13.728 ;
  LAYER M3 ;
        RECT 44.816 11.24 44.848 11.272 ;
  LAYER M1 ;
        RECT 44.752 11.22 44.784 13.728 ;
  LAYER M3 ;
        RECT 44.752 13.676 44.784 13.708 ;
  LAYER M1 ;
        RECT 44.688 11.22 44.72 13.728 ;
  LAYER M3 ;
        RECT 44.688 11.24 44.72 11.272 ;
  LAYER M1 ;
        RECT 44.624 11.22 44.656 13.728 ;
  LAYER M3 ;
        RECT 44.624 13.676 44.656 13.708 ;
  LAYER M1 ;
        RECT 44.56 11.22 44.592 13.728 ;
  LAYER M3 ;
        RECT 44.56 11.24 44.592 11.272 ;
  LAYER M1 ;
        RECT 44.496 11.22 44.528 13.728 ;
  LAYER M3 ;
        RECT 44.496 13.676 44.528 13.708 ;
  LAYER M1 ;
        RECT 44.432 11.22 44.464 13.728 ;
  LAYER M3 ;
        RECT 46.8 11.304 46.832 11.336 ;
  LAYER M2 ;
        RECT 44.432 11.368 44.464 11.4 ;
  LAYER M2 ;
        RECT 46.8 11.432 46.832 11.464 ;
  LAYER M2 ;
        RECT 44.432 11.496 44.464 11.528 ;
  LAYER M2 ;
        RECT 46.8 11.56 46.832 11.592 ;
  LAYER M2 ;
        RECT 44.432 11.624 44.464 11.656 ;
  LAYER M2 ;
        RECT 46.8 11.688 46.832 11.72 ;
  LAYER M2 ;
        RECT 44.432 11.752 44.464 11.784 ;
  LAYER M2 ;
        RECT 46.8 11.816 46.832 11.848 ;
  LAYER M2 ;
        RECT 44.432 11.88 44.464 11.912 ;
  LAYER M2 ;
        RECT 46.8 11.944 46.832 11.976 ;
  LAYER M2 ;
        RECT 44.432 12.008 44.464 12.04 ;
  LAYER M2 ;
        RECT 46.8 12.072 46.832 12.104 ;
  LAYER M2 ;
        RECT 44.432 12.136 44.464 12.168 ;
  LAYER M2 ;
        RECT 46.8 12.2 46.832 12.232 ;
  LAYER M2 ;
        RECT 44.432 12.264 44.464 12.296 ;
  LAYER M2 ;
        RECT 46.8 12.328 46.832 12.36 ;
  LAYER M2 ;
        RECT 44.432 12.392 44.464 12.424 ;
  LAYER M2 ;
        RECT 46.8 12.456 46.832 12.488 ;
  LAYER M2 ;
        RECT 44.432 12.52 44.464 12.552 ;
  LAYER M2 ;
        RECT 46.8 12.584 46.832 12.616 ;
  LAYER M2 ;
        RECT 44.432 12.648 44.464 12.68 ;
  LAYER M2 ;
        RECT 46.8 12.712 46.832 12.744 ;
  LAYER M2 ;
        RECT 44.432 12.776 44.464 12.808 ;
  LAYER M2 ;
        RECT 46.8 12.84 46.832 12.872 ;
  LAYER M2 ;
        RECT 44.432 12.904 44.464 12.936 ;
  LAYER M2 ;
        RECT 46.8 12.968 46.832 13 ;
  LAYER M2 ;
        RECT 44.432 13.032 44.464 13.064 ;
  LAYER M2 ;
        RECT 46.8 13.096 46.832 13.128 ;
  LAYER M2 ;
        RECT 44.432 13.16 44.464 13.192 ;
  LAYER M2 ;
        RECT 46.8 13.224 46.832 13.256 ;
  LAYER M2 ;
        RECT 44.432 13.288 44.464 13.32 ;
  LAYER M2 ;
        RECT 46.8 13.352 46.832 13.384 ;
  LAYER M2 ;
        RECT 44.432 13.416 44.464 13.448 ;
  LAYER M2 ;
        RECT 46.8 13.48 46.832 13.512 ;
  LAYER M2 ;
        RECT 44.432 13.544 44.464 13.576 ;
  LAYER M2 ;
        RECT 44.384 11.172 46.88 13.776 ;
  LAYER M1 ;
        RECT 43.824 1.896 43.856 4.404 ;
  LAYER M3 ;
        RECT 43.824 4.352 43.856 4.384 ;
  LAYER M1 ;
        RECT 43.76 1.896 43.792 4.404 ;
  LAYER M3 ;
        RECT 43.76 1.916 43.792 1.948 ;
  LAYER M1 ;
        RECT 43.696 1.896 43.728 4.404 ;
  LAYER M3 ;
        RECT 43.696 4.352 43.728 4.384 ;
  LAYER M1 ;
        RECT 43.632 1.896 43.664 4.404 ;
  LAYER M3 ;
        RECT 43.632 1.916 43.664 1.948 ;
  LAYER M1 ;
        RECT 43.568 1.896 43.6 4.404 ;
  LAYER M3 ;
        RECT 43.568 4.352 43.6 4.384 ;
  LAYER M1 ;
        RECT 43.504 1.896 43.536 4.404 ;
  LAYER M3 ;
        RECT 43.504 1.916 43.536 1.948 ;
  LAYER M1 ;
        RECT 43.44 1.896 43.472 4.404 ;
  LAYER M3 ;
        RECT 43.44 4.352 43.472 4.384 ;
  LAYER M1 ;
        RECT 43.376 1.896 43.408 4.404 ;
  LAYER M3 ;
        RECT 43.376 1.916 43.408 1.948 ;
  LAYER M1 ;
        RECT 43.312 1.896 43.344 4.404 ;
  LAYER M3 ;
        RECT 43.312 4.352 43.344 4.384 ;
  LAYER M1 ;
        RECT 43.248 1.896 43.28 4.404 ;
  LAYER M3 ;
        RECT 43.248 1.916 43.28 1.948 ;
  LAYER M1 ;
        RECT 43.184 1.896 43.216 4.404 ;
  LAYER M3 ;
        RECT 43.184 4.352 43.216 4.384 ;
  LAYER M1 ;
        RECT 43.12 1.896 43.152 4.404 ;
  LAYER M3 ;
        RECT 43.12 1.916 43.152 1.948 ;
  LAYER M1 ;
        RECT 43.056 1.896 43.088 4.404 ;
  LAYER M3 ;
        RECT 43.056 4.352 43.088 4.384 ;
  LAYER M1 ;
        RECT 42.992 1.896 43.024 4.404 ;
  LAYER M3 ;
        RECT 42.992 1.916 43.024 1.948 ;
  LAYER M1 ;
        RECT 42.928 1.896 42.96 4.404 ;
  LAYER M3 ;
        RECT 42.928 4.352 42.96 4.384 ;
  LAYER M1 ;
        RECT 42.864 1.896 42.896 4.404 ;
  LAYER M3 ;
        RECT 42.864 1.916 42.896 1.948 ;
  LAYER M1 ;
        RECT 42.8 1.896 42.832 4.404 ;
  LAYER M3 ;
        RECT 42.8 4.352 42.832 4.384 ;
  LAYER M1 ;
        RECT 42.736 1.896 42.768 4.404 ;
  LAYER M3 ;
        RECT 42.736 1.916 42.768 1.948 ;
  LAYER M1 ;
        RECT 42.672 1.896 42.704 4.404 ;
  LAYER M3 ;
        RECT 42.672 4.352 42.704 4.384 ;
  LAYER M1 ;
        RECT 42.608 1.896 42.64 4.404 ;
  LAYER M3 ;
        RECT 42.608 1.916 42.64 1.948 ;
  LAYER M1 ;
        RECT 42.544 1.896 42.576 4.404 ;
  LAYER M3 ;
        RECT 42.544 4.352 42.576 4.384 ;
  LAYER M1 ;
        RECT 42.48 1.896 42.512 4.404 ;
  LAYER M3 ;
        RECT 42.48 1.916 42.512 1.948 ;
  LAYER M1 ;
        RECT 42.416 1.896 42.448 4.404 ;
  LAYER M3 ;
        RECT 42.416 4.352 42.448 4.384 ;
  LAYER M1 ;
        RECT 42.352 1.896 42.384 4.404 ;
  LAYER M3 ;
        RECT 42.352 1.916 42.384 1.948 ;
  LAYER M1 ;
        RECT 42.288 1.896 42.32 4.404 ;
  LAYER M3 ;
        RECT 42.288 4.352 42.32 4.384 ;
  LAYER M1 ;
        RECT 42.224 1.896 42.256 4.404 ;
  LAYER M3 ;
        RECT 42.224 1.916 42.256 1.948 ;
  LAYER M1 ;
        RECT 42.16 1.896 42.192 4.404 ;
  LAYER M3 ;
        RECT 42.16 4.352 42.192 4.384 ;
  LAYER M1 ;
        RECT 42.096 1.896 42.128 4.404 ;
  LAYER M3 ;
        RECT 42.096 1.916 42.128 1.948 ;
  LAYER M1 ;
        RECT 42.032 1.896 42.064 4.404 ;
  LAYER M3 ;
        RECT 42.032 4.352 42.064 4.384 ;
  LAYER M1 ;
        RECT 41.968 1.896 42 4.404 ;
  LAYER M3 ;
        RECT 41.968 1.916 42 1.948 ;
  LAYER M1 ;
        RECT 41.904 1.896 41.936 4.404 ;
  LAYER M3 ;
        RECT 41.904 4.352 41.936 4.384 ;
  LAYER M1 ;
        RECT 41.84 1.896 41.872 4.404 ;
  LAYER M3 ;
        RECT 41.84 1.916 41.872 1.948 ;
  LAYER M1 ;
        RECT 41.776 1.896 41.808 4.404 ;
  LAYER M3 ;
        RECT 41.776 4.352 41.808 4.384 ;
  LAYER M1 ;
        RECT 41.712 1.896 41.744 4.404 ;
  LAYER M3 ;
        RECT 41.712 1.916 41.744 1.948 ;
  LAYER M1 ;
        RECT 41.648 1.896 41.68 4.404 ;
  LAYER M3 ;
        RECT 41.648 4.352 41.68 4.384 ;
  LAYER M1 ;
        RECT 41.584 1.896 41.616 4.404 ;
  LAYER M3 ;
        RECT 41.584 1.916 41.616 1.948 ;
  LAYER M1 ;
        RECT 41.52 1.896 41.552 4.404 ;
  LAYER M3 ;
        RECT 41.52 4.352 41.552 4.384 ;
  LAYER M1 ;
        RECT 41.456 1.896 41.488 4.404 ;
  LAYER M3 ;
        RECT 43.824 1.98 43.856 2.012 ;
  LAYER M2 ;
        RECT 41.456 2.044 41.488 2.076 ;
  LAYER M2 ;
        RECT 43.824 2.108 43.856 2.14 ;
  LAYER M2 ;
        RECT 41.456 2.172 41.488 2.204 ;
  LAYER M2 ;
        RECT 43.824 2.236 43.856 2.268 ;
  LAYER M2 ;
        RECT 41.456 2.3 41.488 2.332 ;
  LAYER M2 ;
        RECT 43.824 2.364 43.856 2.396 ;
  LAYER M2 ;
        RECT 41.456 2.428 41.488 2.46 ;
  LAYER M2 ;
        RECT 43.824 2.492 43.856 2.524 ;
  LAYER M2 ;
        RECT 41.456 2.556 41.488 2.588 ;
  LAYER M2 ;
        RECT 43.824 2.62 43.856 2.652 ;
  LAYER M2 ;
        RECT 41.456 2.684 41.488 2.716 ;
  LAYER M2 ;
        RECT 43.824 2.748 43.856 2.78 ;
  LAYER M2 ;
        RECT 41.456 2.812 41.488 2.844 ;
  LAYER M2 ;
        RECT 43.824 2.876 43.856 2.908 ;
  LAYER M2 ;
        RECT 41.456 2.94 41.488 2.972 ;
  LAYER M2 ;
        RECT 43.824 3.004 43.856 3.036 ;
  LAYER M2 ;
        RECT 41.456 3.068 41.488 3.1 ;
  LAYER M2 ;
        RECT 43.824 3.132 43.856 3.164 ;
  LAYER M2 ;
        RECT 41.456 3.196 41.488 3.228 ;
  LAYER M2 ;
        RECT 43.824 3.26 43.856 3.292 ;
  LAYER M2 ;
        RECT 41.456 3.324 41.488 3.356 ;
  LAYER M2 ;
        RECT 43.824 3.388 43.856 3.42 ;
  LAYER M2 ;
        RECT 41.456 3.452 41.488 3.484 ;
  LAYER M2 ;
        RECT 43.824 3.516 43.856 3.548 ;
  LAYER M2 ;
        RECT 41.456 3.58 41.488 3.612 ;
  LAYER M2 ;
        RECT 43.824 3.644 43.856 3.676 ;
  LAYER M2 ;
        RECT 41.456 3.708 41.488 3.74 ;
  LAYER M2 ;
        RECT 43.824 3.772 43.856 3.804 ;
  LAYER M2 ;
        RECT 41.456 3.836 41.488 3.868 ;
  LAYER M2 ;
        RECT 43.824 3.9 43.856 3.932 ;
  LAYER M2 ;
        RECT 41.456 3.964 41.488 3.996 ;
  LAYER M2 ;
        RECT 43.824 4.028 43.856 4.06 ;
  LAYER M2 ;
        RECT 41.456 4.092 41.488 4.124 ;
  LAYER M2 ;
        RECT 43.824 4.156 43.856 4.188 ;
  LAYER M2 ;
        RECT 41.456 4.22 41.488 4.252 ;
  LAYER M2 ;
        RECT 41.408 1.848 43.904 4.452 ;
  LAYER M1 ;
        RECT 43.824 5.004 43.856 7.512 ;
  LAYER M3 ;
        RECT 43.824 7.46 43.856 7.492 ;
  LAYER M1 ;
        RECT 43.76 5.004 43.792 7.512 ;
  LAYER M3 ;
        RECT 43.76 5.024 43.792 5.056 ;
  LAYER M1 ;
        RECT 43.696 5.004 43.728 7.512 ;
  LAYER M3 ;
        RECT 43.696 7.46 43.728 7.492 ;
  LAYER M1 ;
        RECT 43.632 5.004 43.664 7.512 ;
  LAYER M3 ;
        RECT 43.632 5.024 43.664 5.056 ;
  LAYER M1 ;
        RECT 43.568 5.004 43.6 7.512 ;
  LAYER M3 ;
        RECT 43.568 7.46 43.6 7.492 ;
  LAYER M1 ;
        RECT 43.504 5.004 43.536 7.512 ;
  LAYER M3 ;
        RECT 43.504 5.024 43.536 5.056 ;
  LAYER M1 ;
        RECT 43.44 5.004 43.472 7.512 ;
  LAYER M3 ;
        RECT 43.44 7.46 43.472 7.492 ;
  LAYER M1 ;
        RECT 43.376 5.004 43.408 7.512 ;
  LAYER M3 ;
        RECT 43.376 5.024 43.408 5.056 ;
  LAYER M1 ;
        RECT 43.312 5.004 43.344 7.512 ;
  LAYER M3 ;
        RECT 43.312 7.46 43.344 7.492 ;
  LAYER M1 ;
        RECT 43.248 5.004 43.28 7.512 ;
  LAYER M3 ;
        RECT 43.248 5.024 43.28 5.056 ;
  LAYER M1 ;
        RECT 43.184 5.004 43.216 7.512 ;
  LAYER M3 ;
        RECT 43.184 7.46 43.216 7.492 ;
  LAYER M1 ;
        RECT 43.12 5.004 43.152 7.512 ;
  LAYER M3 ;
        RECT 43.12 5.024 43.152 5.056 ;
  LAYER M1 ;
        RECT 43.056 5.004 43.088 7.512 ;
  LAYER M3 ;
        RECT 43.056 7.46 43.088 7.492 ;
  LAYER M1 ;
        RECT 42.992 5.004 43.024 7.512 ;
  LAYER M3 ;
        RECT 42.992 5.024 43.024 5.056 ;
  LAYER M1 ;
        RECT 42.928 5.004 42.96 7.512 ;
  LAYER M3 ;
        RECT 42.928 7.46 42.96 7.492 ;
  LAYER M1 ;
        RECT 42.864 5.004 42.896 7.512 ;
  LAYER M3 ;
        RECT 42.864 5.024 42.896 5.056 ;
  LAYER M1 ;
        RECT 42.8 5.004 42.832 7.512 ;
  LAYER M3 ;
        RECT 42.8 7.46 42.832 7.492 ;
  LAYER M1 ;
        RECT 42.736 5.004 42.768 7.512 ;
  LAYER M3 ;
        RECT 42.736 5.024 42.768 5.056 ;
  LAYER M1 ;
        RECT 42.672 5.004 42.704 7.512 ;
  LAYER M3 ;
        RECT 42.672 7.46 42.704 7.492 ;
  LAYER M1 ;
        RECT 42.608 5.004 42.64 7.512 ;
  LAYER M3 ;
        RECT 42.608 5.024 42.64 5.056 ;
  LAYER M1 ;
        RECT 42.544 5.004 42.576 7.512 ;
  LAYER M3 ;
        RECT 42.544 7.46 42.576 7.492 ;
  LAYER M1 ;
        RECT 42.48 5.004 42.512 7.512 ;
  LAYER M3 ;
        RECT 42.48 5.024 42.512 5.056 ;
  LAYER M1 ;
        RECT 42.416 5.004 42.448 7.512 ;
  LAYER M3 ;
        RECT 42.416 7.46 42.448 7.492 ;
  LAYER M1 ;
        RECT 42.352 5.004 42.384 7.512 ;
  LAYER M3 ;
        RECT 42.352 5.024 42.384 5.056 ;
  LAYER M1 ;
        RECT 42.288 5.004 42.32 7.512 ;
  LAYER M3 ;
        RECT 42.288 7.46 42.32 7.492 ;
  LAYER M1 ;
        RECT 42.224 5.004 42.256 7.512 ;
  LAYER M3 ;
        RECT 42.224 5.024 42.256 5.056 ;
  LAYER M1 ;
        RECT 42.16 5.004 42.192 7.512 ;
  LAYER M3 ;
        RECT 42.16 7.46 42.192 7.492 ;
  LAYER M1 ;
        RECT 42.096 5.004 42.128 7.512 ;
  LAYER M3 ;
        RECT 42.096 5.024 42.128 5.056 ;
  LAYER M1 ;
        RECT 42.032 5.004 42.064 7.512 ;
  LAYER M3 ;
        RECT 42.032 7.46 42.064 7.492 ;
  LAYER M1 ;
        RECT 41.968 5.004 42 7.512 ;
  LAYER M3 ;
        RECT 41.968 5.024 42 5.056 ;
  LAYER M1 ;
        RECT 41.904 5.004 41.936 7.512 ;
  LAYER M3 ;
        RECT 41.904 7.46 41.936 7.492 ;
  LAYER M1 ;
        RECT 41.84 5.004 41.872 7.512 ;
  LAYER M3 ;
        RECT 41.84 5.024 41.872 5.056 ;
  LAYER M1 ;
        RECT 41.776 5.004 41.808 7.512 ;
  LAYER M3 ;
        RECT 41.776 7.46 41.808 7.492 ;
  LAYER M1 ;
        RECT 41.712 5.004 41.744 7.512 ;
  LAYER M3 ;
        RECT 41.712 5.024 41.744 5.056 ;
  LAYER M1 ;
        RECT 41.648 5.004 41.68 7.512 ;
  LAYER M3 ;
        RECT 41.648 7.46 41.68 7.492 ;
  LAYER M1 ;
        RECT 41.584 5.004 41.616 7.512 ;
  LAYER M3 ;
        RECT 41.584 5.024 41.616 5.056 ;
  LAYER M1 ;
        RECT 41.52 5.004 41.552 7.512 ;
  LAYER M3 ;
        RECT 41.52 7.46 41.552 7.492 ;
  LAYER M1 ;
        RECT 41.456 5.004 41.488 7.512 ;
  LAYER M3 ;
        RECT 43.824 5.088 43.856 5.12 ;
  LAYER M2 ;
        RECT 41.456 5.152 41.488 5.184 ;
  LAYER M2 ;
        RECT 43.824 5.216 43.856 5.248 ;
  LAYER M2 ;
        RECT 41.456 5.28 41.488 5.312 ;
  LAYER M2 ;
        RECT 43.824 5.344 43.856 5.376 ;
  LAYER M2 ;
        RECT 41.456 5.408 41.488 5.44 ;
  LAYER M2 ;
        RECT 43.824 5.472 43.856 5.504 ;
  LAYER M2 ;
        RECT 41.456 5.536 41.488 5.568 ;
  LAYER M2 ;
        RECT 43.824 5.6 43.856 5.632 ;
  LAYER M2 ;
        RECT 41.456 5.664 41.488 5.696 ;
  LAYER M2 ;
        RECT 43.824 5.728 43.856 5.76 ;
  LAYER M2 ;
        RECT 41.456 5.792 41.488 5.824 ;
  LAYER M2 ;
        RECT 43.824 5.856 43.856 5.888 ;
  LAYER M2 ;
        RECT 41.456 5.92 41.488 5.952 ;
  LAYER M2 ;
        RECT 43.824 5.984 43.856 6.016 ;
  LAYER M2 ;
        RECT 41.456 6.048 41.488 6.08 ;
  LAYER M2 ;
        RECT 43.824 6.112 43.856 6.144 ;
  LAYER M2 ;
        RECT 41.456 6.176 41.488 6.208 ;
  LAYER M2 ;
        RECT 43.824 6.24 43.856 6.272 ;
  LAYER M2 ;
        RECT 41.456 6.304 41.488 6.336 ;
  LAYER M2 ;
        RECT 43.824 6.368 43.856 6.4 ;
  LAYER M2 ;
        RECT 41.456 6.432 41.488 6.464 ;
  LAYER M2 ;
        RECT 43.824 6.496 43.856 6.528 ;
  LAYER M2 ;
        RECT 41.456 6.56 41.488 6.592 ;
  LAYER M2 ;
        RECT 43.824 6.624 43.856 6.656 ;
  LAYER M2 ;
        RECT 41.456 6.688 41.488 6.72 ;
  LAYER M2 ;
        RECT 43.824 6.752 43.856 6.784 ;
  LAYER M2 ;
        RECT 41.456 6.816 41.488 6.848 ;
  LAYER M2 ;
        RECT 43.824 6.88 43.856 6.912 ;
  LAYER M2 ;
        RECT 41.456 6.944 41.488 6.976 ;
  LAYER M2 ;
        RECT 43.824 7.008 43.856 7.04 ;
  LAYER M2 ;
        RECT 41.456 7.072 41.488 7.104 ;
  LAYER M2 ;
        RECT 43.824 7.136 43.856 7.168 ;
  LAYER M2 ;
        RECT 41.456 7.2 41.488 7.232 ;
  LAYER M2 ;
        RECT 43.824 7.264 43.856 7.296 ;
  LAYER M2 ;
        RECT 41.456 7.328 41.488 7.36 ;
  LAYER M2 ;
        RECT 41.408 4.956 43.904 7.56 ;
  LAYER M1 ;
        RECT 43.824 8.112 43.856 10.62 ;
  LAYER M3 ;
        RECT 43.824 10.568 43.856 10.6 ;
  LAYER M1 ;
        RECT 43.76 8.112 43.792 10.62 ;
  LAYER M3 ;
        RECT 43.76 8.132 43.792 8.164 ;
  LAYER M1 ;
        RECT 43.696 8.112 43.728 10.62 ;
  LAYER M3 ;
        RECT 43.696 10.568 43.728 10.6 ;
  LAYER M1 ;
        RECT 43.632 8.112 43.664 10.62 ;
  LAYER M3 ;
        RECT 43.632 8.132 43.664 8.164 ;
  LAYER M1 ;
        RECT 43.568 8.112 43.6 10.62 ;
  LAYER M3 ;
        RECT 43.568 10.568 43.6 10.6 ;
  LAYER M1 ;
        RECT 43.504 8.112 43.536 10.62 ;
  LAYER M3 ;
        RECT 43.504 8.132 43.536 8.164 ;
  LAYER M1 ;
        RECT 43.44 8.112 43.472 10.62 ;
  LAYER M3 ;
        RECT 43.44 10.568 43.472 10.6 ;
  LAYER M1 ;
        RECT 43.376 8.112 43.408 10.62 ;
  LAYER M3 ;
        RECT 43.376 8.132 43.408 8.164 ;
  LAYER M1 ;
        RECT 43.312 8.112 43.344 10.62 ;
  LAYER M3 ;
        RECT 43.312 10.568 43.344 10.6 ;
  LAYER M1 ;
        RECT 43.248 8.112 43.28 10.62 ;
  LAYER M3 ;
        RECT 43.248 8.132 43.28 8.164 ;
  LAYER M1 ;
        RECT 43.184 8.112 43.216 10.62 ;
  LAYER M3 ;
        RECT 43.184 10.568 43.216 10.6 ;
  LAYER M1 ;
        RECT 43.12 8.112 43.152 10.62 ;
  LAYER M3 ;
        RECT 43.12 8.132 43.152 8.164 ;
  LAYER M1 ;
        RECT 43.056 8.112 43.088 10.62 ;
  LAYER M3 ;
        RECT 43.056 10.568 43.088 10.6 ;
  LAYER M1 ;
        RECT 42.992 8.112 43.024 10.62 ;
  LAYER M3 ;
        RECT 42.992 8.132 43.024 8.164 ;
  LAYER M1 ;
        RECT 42.928 8.112 42.96 10.62 ;
  LAYER M3 ;
        RECT 42.928 10.568 42.96 10.6 ;
  LAYER M1 ;
        RECT 42.864 8.112 42.896 10.62 ;
  LAYER M3 ;
        RECT 42.864 8.132 42.896 8.164 ;
  LAYER M1 ;
        RECT 42.8 8.112 42.832 10.62 ;
  LAYER M3 ;
        RECT 42.8 10.568 42.832 10.6 ;
  LAYER M1 ;
        RECT 42.736 8.112 42.768 10.62 ;
  LAYER M3 ;
        RECT 42.736 8.132 42.768 8.164 ;
  LAYER M1 ;
        RECT 42.672 8.112 42.704 10.62 ;
  LAYER M3 ;
        RECT 42.672 10.568 42.704 10.6 ;
  LAYER M1 ;
        RECT 42.608 8.112 42.64 10.62 ;
  LAYER M3 ;
        RECT 42.608 8.132 42.64 8.164 ;
  LAYER M1 ;
        RECT 42.544 8.112 42.576 10.62 ;
  LAYER M3 ;
        RECT 42.544 10.568 42.576 10.6 ;
  LAYER M1 ;
        RECT 42.48 8.112 42.512 10.62 ;
  LAYER M3 ;
        RECT 42.48 8.132 42.512 8.164 ;
  LAYER M1 ;
        RECT 42.416 8.112 42.448 10.62 ;
  LAYER M3 ;
        RECT 42.416 10.568 42.448 10.6 ;
  LAYER M1 ;
        RECT 42.352 8.112 42.384 10.62 ;
  LAYER M3 ;
        RECT 42.352 8.132 42.384 8.164 ;
  LAYER M1 ;
        RECT 42.288 8.112 42.32 10.62 ;
  LAYER M3 ;
        RECT 42.288 10.568 42.32 10.6 ;
  LAYER M1 ;
        RECT 42.224 8.112 42.256 10.62 ;
  LAYER M3 ;
        RECT 42.224 8.132 42.256 8.164 ;
  LAYER M1 ;
        RECT 42.16 8.112 42.192 10.62 ;
  LAYER M3 ;
        RECT 42.16 10.568 42.192 10.6 ;
  LAYER M1 ;
        RECT 42.096 8.112 42.128 10.62 ;
  LAYER M3 ;
        RECT 42.096 8.132 42.128 8.164 ;
  LAYER M1 ;
        RECT 42.032 8.112 42.064 10.62 ;
  LAYER M3 ;
        RECT 42.032 10.568 42.064 10.6 ;
  LAYER M1 ;
        RECT 41.968 8.112 42 10.62 ;
  LAYER M3 ;
        RECT 41.968 8.132 42 8.164 ;
  LAYER M1 ;
        RECT 41.904 8.112 41.936 10.62 ;
  LAYER M3 ;
        RECT 41.904 10.568 41.936 10.6 ;
  LAYER M1 ;
        RECT 41.84 8.112 41.872 10.62 ;
  LAYER M3 ;
        RECT 41.84 8.132 41.872 8.164 ;
  LAYER M1 ;
        RECT 41.776 8.112 41.808 10.62 ;
  LAYER M3 ;
        RECT 41.776 10.568 41.808 10.6 ;
  LAYER M1 ;
        RECT 41.712 8.112 41.744 10.62 ;
  LAYER M3 ;
        RECT 41.712 8.132 41.744 8.164 ;
  LAYER M1 ;
        RECT 41.648 8.112 41.68 10.62 ;
  LAYER M3 ;
        RECT 41.648 10.568 41.68 10.6 ;
  LAYER M1 ;
        RECT 41.584 8.112 41.616 10.62 ;
  LAYER M3 ;
        RECT 41.584 8.132 41.616 8.164 ;
  LAYER M1 ;
        RECT 41.52 8.112 41.552 10.62 ;
  LAYER M3 ;
        RECT 41.52 10.568 41.552 10.6 ;
  LAYER M1 ;
        RECT 41.456 8.112 41.488 10.62 ;
  LAYER M3 ;
        RECT 43.824 8.196 43.856 8.228 ;
  LAYER M2 ;
        RECT 41.456 8.26 41.488 8.292 ;
  LAYER M2 ;
        RECT 43.824 8.324 43.856 8.356 ;
  LAYER M2 ;
        RECT 41.456 8.388 41.488 8.42 ;
  LAYER M2 ;
        RECT 43.824 8.452 43.856 8.484 ;
  LAYER M2 ;
        RECT 41.456 8.516 41.488 8.548 ;
  LAYER M2 ;
        RECT 43.824 8.58 43.856 8.612 ;
  LAYER M2 ;
        RECT 41.456 8.644 41.488 8.676 ;
  LAYER M2 ;
        RECT 43.824 8.708 43.856 8.74 ;
  LAYER M2 ;
        RECT 41.456 8.772 41.488 8.804 ;
  LAYER M2 ;
        RECT 43.824 8.836 43.856 8.868 ;
  LAYER M2 ;
        RECT 41.456 8.9 41.488 8.932 ;
  LAYER M2 ;
        RECT 43.824 8.964 43.856 8.996 ;
  LAYER M2 ;
        RECT 41.456 9.028 41.488 9.06 ;
  LAYER M2 ;
        RECT 43.824 9.092 43.856 9.124 ;
  LAYER M2 ;
        RECT 41.456 9.156 41.488 9.188 ;
  LAYER M2 ;
        RECT 43.824 9.22 43.856 9.252 ;
  LAYER M2 ;
        RECT 41.456 9.284 41.488 9.316 ;
  LAYER M2 ;
        RECT 43.824 9.348 43.856 9.38 ;
  LAYER M2 ;
        RECT 41.456 9.412 41.488 9.444 ;
  LAYER M2 ;
        RECT 43.824 9.476 43.856 9.508 ;
  LAYER M2 ;
        RECT 41.456 9.54 41.488 9.572 ;
  LAYER M2 ;
        RECT 43.824 9.604 43.856 9.636 ;
  LAYER M2 ;
        RECT 41.456 9.668 41.488 9.7 ;
  LAYER M2 ;
        RECT 43.824 9.732 43.856 9.764 ;
  LAYER M2 ;
        RECT 41.456 9.796 41.488 9.828 ;
  LAYER M2 ;
        RECT 43.824 9.86 43.856 9.892 ;
  LAYER M2 ;
        RECT 41.456 9.924 41.488 9.956 ;
  LAYER M2 ;
        RECT 43.824 9.988 43.856 10.02 ;
  LAYER M2 ;
        RECT 41.456 10.052 41.488 10.084 ;
  LAYER M2 ;
        RECT 43.824 10.116 43.856 10.148 ;
  LAYER M2 ;
        RECT 41.456 10.18 41.488 10.212 ;
  LAYER M2 ;
        RECT 43.824 10.244 43.856 10.276 ;
  LAYER M2 ;
        RECT 41.456 10.308 41.488 10.34 ;
  LAYER M2 ;
        RECT 43.824 10.372 43.856 10.404 ;
  LAYER M2 ;
        RECT 41.456 10.436 41.488 10.468 ;
  LAYER M2 ;
        RECT 41.408 8.064 43.904 10.668 ;
  LAYER M1 ;
        RECT 43.824 11.22 43.856 13.728 ;
  LAYER M3 ;
        RECT 43.824 13.676 43.856 13.708 ;
  LAYER M1 ;
        RECT 43.76 11.22 43.792 13.728 ;
  LAYER M3 ;
        RECT 43.76 11.24 43.792 11.272 ;
  LAYER M1 ;
        RECT 43.696 11.22 43.728 13.728 ;
  LAYER M3 ;
        RECT 43.696 13.676 43.728 13.708 ;
  LAYER M1 ;
        RECT 43.632 11.22 43.664 13.728 ;
  LAYER M3 ;
        RECT 43.632 11.24 43.664 11.272 ;
  LAYER M1 ;
        RECT 43.568 11.22 43.6 13.728 ;
  LAYER M3 ;
        RECT 43.568 13.676 43.6 13.708 ;
  LAYER M1 ;
        RECT 43.504 11.22 43.536 13.728 ;
  LAYER M3 ;
        RECT 43.504 11.24 43.536 11.272 ;
  LAYER M1 ;
        RECT 43.44 11.22 43.472 13.728 ;
  LAYER M3 ;
        RECT 43.44 13.676 43.472 13.708 ;
  LAYER M1 ;
        RECT 43.376 11.22 43.408 13.728 ;
  LAYER M3 ;
        RECT 43.376 11.24 43.408 11.272 ;
  LAYER M1 ;
        RECT 43.312 11.22 43.344 13.728 ;
  LAYER M3 ;
        RECT 43.312 13.676 43.344 13.708 ;
  LAYER M1 ;
        RECT 43.248 11.22 43.28 13.728 ;
  LAYER M3 ;
        RECT 43.248 11.24 43.28 11.272 ;
  LAYER M1 ;
        RECT 43.184 11.22 43.216 13.728 ;
  LAYER M3 ;
        RECT 43.184 13.676 43.216 13.708 ;
  LAYER M1 ;
        RECT 43.12 11.22 43.152 13.728 ;
  LAYER M3 ;
        RECT 43.12 11.24 43.152 11.272 ;
  LAYER M1 ;
        RECT 43.056 11.22 43.088 13.728 ;
  LAYER M3 ;
        RECT 43.056 13.676 43.088 13.708 ;
  LAYER M1 ;
        RECT 42.992 11.22 43.024 13.728 ;
  LAYER M3 ;
        RECT 42.992 11.24 43.024 11.272 ;
  LAYER M1 ;
        RECT 42.928 11.22 42.96 13.728 ;
  LAYER M3 ;
        RECT 42.928 13.676 42.96 13.708 ;
  LAYER M1 ;
        RECT 42.864 11.22 42.896 13.728 ;
  LAYER M3 ;
        RECT 42.864 11.24 42.896 11.272 ;
  LAYER M1 ;
        RECT 42.8 11.22 42.832 13.728 ;
  LAYER M3 ;
        RECT 42.8 13.676 42.832 13.708 ;
  LAYER M1 ;
        RECT 42.736 11.22 42.768 13.728 ;
  LAYER M3 ;
        RECT 42.736 11.24 42.768 11.272 ;
  LAYER M1 ;
        RECT 42.672 11.22 42.704 13.728 ;
  LAYER M3 ;
        RECT 42.672 13.676 42.704 13.708 ;
  LAYER M1 ;
        RECT 42.608 11.22 42.64 13.728 ;
  LAYER M3 ;
        RECT 42.608 11.24 42.64 11.272 ;
  LAYER M1 ;
        RECT 42.544 11.22 42.576 13.728 ;
  LAYER M3 ;
        RECT 42.544 13.676 42.576 13.708 ;
  LAYER M1 ;
        RECT 42.48 11.22 42.512 13.728 ;
  LAYER M3 ;
        RECT 42.48 11.24 42.512 11.272 ;
  LAYER M1 ;
        RECT 42.416 11.22 42.448 13.728 ;
  LAYER M3 ;
        RECT 42.416 13.676 42.448 13.708 ;
  LAYER M1 ;
        RECT 42.352 11.22 42.384 13.728 ;
  LAYER M3 ;
        RECT 42.352 11.24 42.384 11.272 ;
  LAYER M1 ;
        RECT 42.288 11.22 42.32 13.728 ;
  LAYER M3 ;
        RECT 42.288 13.676 42.32 13.708 ;
  LAYER M1 ;
        RECT 42.224 11.22 42.256 13.728 ;
  LAYER M3 ;
        RECT 42.224 11.24 42.256 11.272 ;
  LAYER M1 ;
        RECT 42.16 11.22 42.192 13.728 ;
  LAYER M3 ;
        RECT 42.16 13.676 42.192 13.708 ;
  LAYER M1 ;
        RECT 42.096 11.22 42.128 13.728 ;
  LAYER M3 ;
        RECT 42.096 11.24 42.128 11.272 ;
  LAYER M1 ;
        RECT 42.032 11.22 42.064 13.728 ;
  LAYER M3 ;
        RECT 42.032 13.676 42.064 13.708 ;
  LAYER M1 ;
        RECT 41.968 11.22 42 13.728 ;
  LAYER M3 ;
        RECT 41.968 11.24 42 11.272 ;
  LAYER M1 ;
        RECT 41.904 11.22 41.936 13.728 ;
  LAYER M3 ;
        RECT 41.904 13.676 41.936 13.708 ;
  LAYER M1 ;
        RECT 41.84 11.22 41.872 13.728 ;
  LAYER M3 ;
        RECT 41.84 11.24 41.872 11.272 ;
  LAYER M1 ;
        RECT 41.776 11.22 41.808 13.728 ;
  LAYER M3 ;
        RECT 41.776 13.676 41.808 13.708 ;
  LAYER M1 ;
        RECT 41.712 11.22 41.744 13.728 ;
  LAYER M3 ;
        RECT 41.712 11.24 41.744 11.272 ;
  LAYER M1 ;
        RECT 41.648 11.22 41.68 13.728 ;
  LAYER M3 ;
        RECT 41.648 13.676 41.68 13.708 ;
  LAYER M1 ;
        RECT 41.584 11.22 41.616 13.728 ;
  LAYER M3 ;
        RECT 41.584 11.24 41.616 11.272 ;
  LAYER M1 ;
        RECT 41.52 11.22 41.552 13.728 ;
  LAYER M3 ;
        RECT 41.52 13.676 41.552 13.708 ;
  LAYER M1 ;
        RECT 41.456 11.22 41.488 13.728 ;
  LAYER M3 ;
        RECT 43.824 11.304 43.856 11.336 ;
  LAYER M2 ;
        RECT 41.456 11.368 41.488 11.4 ;
  LAYER M2 ;
        RECT 43.824 11.432 43.856 11.464 ;
  LAYER M2 ;
        RECT 41.456 11.496 41.488 11.528 ;
  LAYER M2 ;
        RECT 43.824 11.56 43.856 11.592 ;
  LAYER M2 ;
        RECT 41.456 11.624 41.488 11.656 ;
  LAYER M2 ;
        RECT 43.824 11.688 43.856 11.72 ;
  LAYER M2 ;
        RECT 41.456 11.752 41.488 11.784 ;
  LAYER M2 ;
        RECT 43.824 11.816 43.856 11.848 ;
  LAYER M2 ;
        RECT 41.456 11.88 41.488 11.912 ;
  LAYER M2 ;
        RECT 43.824 11.944 43.856 11.976 ;
  LAYER M2 ;
        RECT 41.456 12.008 41.488 12.04 ;
  LAYER M2 ;
        RECT 43.824 12.072 43.856 12.104 ;
  LAYER M2 ;
        RECT 41.456 12.136 41.488 12.168 ;
  LAYER M2 ;
        RECT 43.824 12.2 43.856 12.232 ;
  LAYER M2 ;
        RECT 41.456 12.264 41.488 12.296 ;
  LAYER M2 ;
        RECT 43.824 12.328 43.856 12.36 ;
  LAYER M2 ;
        RECT 41.456 12.392 41.488 12.424 ;
  LAYER M2 ;
        RECT 43.824 12.456 43.856 12.488 ;
  LAYER M2 ;
        RECT 41.456 12.52 41.488 12.552 ;
  LAYER M2 ;
        RECT 43.824 12.584 43.856 12.616 ;
  LAYER M2 ;
        RECT 41.456 12.648 41.488 12.68 ;
  LAYER M2 ;
        RECT 43.824 12.712 43.856 12.744 ;
  LAYER M2 ;
        RECT 41.456 12.776 41.488 12.808 ;
  LAYER M2 ;
        RECT 43.824 12.84 43.856 12.872 ;
  LAYER M2 ;
        RECT 41.456 12.904 41.488 12.936 ;
  LAYER M2 ;
        RECT 43.824 12.968 43.856 13 ;
  LAYER M2 ;
        RECT 41.456 13.032 41.488 13.064 ;
  LAYER M2 ;
        RECT 43.824 13.096 43.856 13.128 ;
  LAYER M2 ;
        RECT 41.456 13.16 41.488 13.192 ;
  LAYER M2 ;
        RECT 43.824 13.224 43.856 13.256 ;
  LAYER M2 ;
        RECT 41.456 13.288 41.488 13.32 ;
  LAYER M2 ;
        RECT 43.824 13.352 43.856 13.384 ;
  LAYER M2 ;
        RECT 41.456 13.416 41.488 13.448 ;
  LAYER M2 ;
        RECT 43.824 13.48 43.856 13.512 ;
  LAYER M2 ;
        RECT 41.456 13.544 41.488 13.576 ;
  LAYER M2 ;
        RECT 41.408 11.172 43.904 13.776 ;
  LAYER M1 ;
        RECT 40.848 1.896 40.88 4.404 ;
  LAYER M3 ;
        RECT 40.848 4.352 40.88 4.384 ;
  LAYER M1 ;
        RECT 40.784 1.896 40.816 4.404 ;
  LAYER M3 ;
        RECT 40.784 1.916 40.816 1.948 ;
  LAYER M1 ;
        RECT 40.72 1.896 40.752 4.404 ;
  LAYER M3 ;
        RECT 40.72 4.352 40.752 4.384 ;
  LAYER M1 ;
        RECT 40.656 1.896 40.688 4.404 ;
  LAYER M3 ;
        RECT 40.656 1.916 40.688 1.948 ;
  LAYER M1 ;
        RECT 40.592 1.896 40.624 4.404 ;
  LAYER M3 ;
        RECT 40.592 4.352 40.624 4.384 ;
  LAYER M1 ;
        RECT 40.528 1.896 40.56 4.404 ;
  LAYER M3 ;
        RECT 40.528 1.916 40.56 1.948 ;
  LAYER M1 ;
        RECT 40.464 1.896 40.496 4.404 ;
  LAYER M3 ;
        RECT 40.464 4.352 40.496 4.384 ;
  LAYER M1 ;
        RECT 40.4 1.896 40.432 4.404 ;
  LAYER M3 ;
        RECT 40.4 1.916 40.432 1.948 ;
  LAYER M1 ;
        RECT 40.336 1.896 40.368 4.404 ;
  LAYER M3 ;
        RECT 40.336 4.352 40.368 4.384 ;
  LAYER M1 ;
        RECT 40.272 1.896 40.304 4.404 ;
  LAYER M3 ;
        RECT 40.272 1.916 40.304 1.948 ;
  LAYER M1 ;
        RECT 40.208 1.896 40.24 4.404 ;
  LAYER M3 ;
        RECT 40.208 4.352 40.24 4.384 ;
  LAYER M1 ;
        RECT 40.144 1.896 40.176 4.404 ;
  LAYER M3 ;
        RECT 40.144 1.916 40.176 1.948 ;
  LAYER M1 ;
        RECT 40.08 1.896 40.112 4.404 ;
  LAYER M3 ;
        RECT 40.08 4.352 40.112 4.384 ;
  LAYER M1 ;
        RECT 40.016 1.896 40.048 4.404 ;
  LAYER M3 ;
        RECT 40.016 1.916 40.048 1.948 ;
  LAYER M1 ;
        RECT 39.952 1.896 39.984 4.404 ;
  LAYER M3 ;
        RECT 39.952 4.352 39.984 4.384 ;
  LAYER M1 ;
        RECT 39.888 1.896 39.92 4.404 ;
  LAYER M3 ;
        RECT 39.888 1.916 39.92 1.948 ;
  LAYER M1 ;
        RECT 39.824 1.896 39.856 4.404 ;
  LAYER M3 ;
        RECT 39.824 4.352 39.856 4.384 ;
  LAYER M1 ;
        RECT 39.76 1.896 39.792 4.404 ;
  LAYER M3 ;
        RECT 39.76 1.916 39.792 1.948 ;
  LAYER M1 ;
        RECT 39.696 1.896 39.728 4.404 ;
  LAYER M3 ;
        RECT 39.696 4.352 39.728 4.384 ;
  LAYER M1 ;
        RECT 39.632 1.896 39.664 4.404 ;
  LAYER M3 ;
        RECT 39.632 1.916 39.664 1.948 ;
  LAYER M1 ;
        RECT 39.568 1.896 39.6 4.404 ;
  LAYER M3 ;
        RECT 39.568 4.352 39.6 4.384 ;
  LAYER M1 ;
        RECT 39.504 1.896 39.536 4.404 ;
  LAYER M3 ;
        RECT 39.504 1.916 39.536 1.948 ;
  LAYER M1 ;
        RECT 39.44 1.896 39.472 4.404 ;
  LAYER M3 ;
        RECT 39.44 4.352 39.472 4.384 ;
  LAYER M1 ;
        RECT 39.376 1.896 39.408 4.404 ;
  LAYER M3 ;
        RECT 39.376 1.916 39.408 1.948 ;
  LAYER M1 ;
        RECT 39.312 1.896 39.344 4.404 ;
  LAYER M3 ;
        RECT 39.312 4.352 39.344 4.384 ;
  LAYER M1 ;
        RECT 39.248 1.896 39.28 4.404 ;
  LAYER M3 ;
        RECT 39.248 1.916 39.28 1.948 ;
  LAYER M1 ;
        RECT 39.184 1.896 39.216 4.404 ;
  LAYER M3 ;
        RECT 39.184 4.352 39.216 4.384 ;
  LAYER M1 ;
        RECT 39.12 1.896 39.152 4.404 ;
  LAYER M3 ;
        RECT 39.12 1.916 39.152 1.948 ;
  LAYER M1 ;
        RECT 39.056 1.896 39.088 4.404 ;
  LAYER M3 ;
        RECT 39.056 4.352 39.088 4.384 ;
  LAYER M1 ;
        RECT 38.992 1.896 39.024 4.404 ;
  LAYER M3 ;
        RECT 38.992 1.916 39.024 1.948 ;
  LAYER M1 ;
        RECT 38.928 1.896 38.96 4.404 ;
  LAYER M3 ;
        RECT 38.928 4.352 38.96 4.384 ;
  LAYER M1 ;
        RECT 38.864 1.896 38.896 4.404 ;
  LAYER M3 ;
        RECT 38.864 1.916 38.896 1.948 ;
  LAYER M1 ;
        RECT 38.8 1.896 38.832 4.404 ;
  LAYER M3 ;
        RECT 38.8 4.352 38.832 4.384 ;
  LAYER M1 ;
        RECT 38.736 1.896 38.768 4.404 ;
  LAYER M3 ;
        RECT 38.736 1.916 38.768 1.948 ;
  LAYER M1 ;
        RECT 38.672 1.896 38.704 4.404 ;
  LAYER M3 ;
        RECT 38.672 4.352 38.704 4.384 ;
  LAYER M1 ;
        RECT 38.608 1.896 38.64 4.404 ;
  LAYER M3 ;
        RECT 38.608 1.916 38.64 1.948 ;
  LAYER M1 ;
        RECT 38.544 1.896 38.576 4.404 ;
  LAYER M3 ;
        RECT 38.544 4.352 38.576 4.384 ;
  LAYER M1 ;
        RECT 38.48 1.896 38.512 4.404 ;
  LAYER M3 ;
        RECT 40.848 1.98 40.88 2.012 ;
  LAYER M2 ;
        RECT 38.48 2.044 38.512 2.076 ;
  LAYER M2 ;
        RECT 40.848 2.108 40.88 2.14 ;
  LAYER M2 ;
        RECT 38.48 2.172 38.512 2.204 ;
  LAYER M2 ;
        RECT 40.848 2.236 40.88 2.268 ;
  LAYER M2 ;
        RECT 38.48 2.3 38.512 2.332 ;
  LAYER M2 ;
        RECT 40.848 2.364 40.88 2.396 ;
  LAYER M2 ;
        RECT 38.48 2.428 38.512 2.46 ;
  LAYER M2 ;
        RECT 40.848 2.492 40.88 2.524 ;
  LAYER M2 ;
        RECT 38.48 2.556 38.512 2.588 ;
  LAYER M2 ;
        RECT 40.848 2.62 40.88 2.652 ;
  LAYER M2 ;
        RECT 38.48 2.684 38.512 2.716 ;
  LAYER M2 ;
        RECT 40.848 2.748 40.88 2.78 ;
  LAYER M2 ;
        RECT 38.48 2.812 38.512 2.844 ;
  LAYER M2 ;
        RECT 40.848 2.876 40.88 2.908 ;
  LAYER M2 ;
        RECT 38.48 2.94 38.512 2.972 ;
  LAYER M2 ;
        RECT 40.848 3.004 40.88 3.036 ;
  LAYER M2 ;
        RECT 38.48 3.068 38.512 3.1 ;
  LAYER M2 ;
        RECT 40.848 3.132 40.88 3.164 ;
  LAYER M2 ;
        RECT 38.48 3.196 38.512 3.228 ;
  LAYER M2 ;
        RECT 40.848 3.26 40.88 3.292 ;
  LAYER M2 ;
        RECT 38.48 3.324 38.512 3.356 ;
  LAYER M2 ;
        RECT 40.848 3.388 40.88 3.42 ;
  LAYER M2 ;
        RECT 38.48 3.452 38.512 3.484 ;
  LAYER M2 ;
        RECT 40.848 3.516 40.88 3.548 ;
  LAYER M2 ;
        RECT 38.48 3.58 38.512 3.612 ;
  LAYER M2 ;
        RECT 40.848 3.644 40.88 3.676 ;
  LAYER M2 ;
        RECT 38.48 3.708 38.512 3.74 ;
  LAYER M2 ;
        RECT 40.848 3.772 40.88 3.804 ;
  LAYER M2 ;
        RECT 38.48 3.836 38.512 3.868 ;
  LAYER M2 ;
        RECT 40.848 3.9 40.88 3.932 ;
  LAYER M2 ;
        RECT 38.48 3.964 38.512 3.996 ;
  LAYER M2 ;
        RECT 40.848 4.028 40.88 4.06 ;
  LAYER M2 ;
        RECT 38.48 4.092 38.512 4.124 ;
  LAYER M2 ;
        RECT 40.848 4.156 40.88 4.188 ;
  LAYER M2 ;
        RECT 38.48 4.22 38.512 4.252 ;
  LAYER M2 ;
        RECT 38.432 1.848 40.928 4.452 ;
  LAYER M1 ;
        RECT 40.848 5.004 40.88 7.512 ;
  LAYER M3 ;
        RECT 40.848 7.46 40.88 7.492 ;
  LAYER M1 ;
        RECT 40.784 5.004 40.816 7.512 ;
  LAYER M3 ;
        RECT 40.784 5.024 40.816 5.056 ;
  LAYER M1 ;
        RECT 40.72 5.004 40.752 7.512 ;
  LAYER M3 ;
        RECT 40.72 7.46 40.752 7.492 ;
  LAYER M1 ;
        RECT 40.656 5.004 40.688 7.512 ;
  LAYER M3 ;
        RECT 40.656 5.024 40.688 5.056 ;
  LAYER M1 ;
        RECT 40.592 5.004 40.624 7.512 ;
  LAYER M3 ;
        RECT 40.592 7.46 40.624 7.492 ;
  LAYER M1 ;
        RECT 40.528 5.004 40.56 7.512 ;
  LAYER M3 ;
        RECT 40.528 5.024 40.56 5.056 ;
  LAYER M1 ;
        RECT 40.464 5.004 40.496 7.512 ;
  LAYER M3 ;
        RECT 40.464 7.46 40.496 7.492 ;
  LAYER M1 ;
        RECT 40.4 5.004 40.432 7.512 ;
  LAYER M3 ;
        RECT 40.4 5.024 40.432 5.056 ;
  LAYER M1 ;
        RECT 40.336 5.004 40.368 7.512 ;
  LAYER M3 ;
        RECT 40.336 7.46 40.368 7.492 ;
  LAYER M1 ;
        RECT 40.272 5.004 40.304 7.512 ;
  LAYER M3 ;
        RECT 40.272 5.024 40.304 5.056 ;
  LAYER M1 ;
        RECT 40.208 5.004 40.24 7.512 ;
  LAYER M3 ;
        RECT 40.208 7.46 40.24 7.492 ;
  LAYER M1 ;
        RECT 40.144 5.004 40.176 7.512 ;
  LAYER M3 ;
        RECT 40.144 5.024 40.176 5.056 ;
  LAYER M1 ;
        RECT 40.08 5.004 40.112 7.512 ;
  LAYER M3 ;
        RECT 40.08 7.46 40.112 7.492 ;
  LAYER M1 ;
        RECT 40.016 5.004 40.048 7.512 ;
  LAYER M3 ;
        RECT 40.016 5.024 40.048 5.056 ;
  LAYER M1 ;
        RECT 39.952 5.004 39.984 7.512 ;
  LAYER M3 ;
        RECT 39.952 7.46 39.984 7.492 ;
  LAYER M1 ;
        RECT 39.888 5.004 39.92 7.512 ;
  LAYER M3 ;
        RECT 39.888 5.024 39.92 5.056 ;
  LAYER M1 ;
        RECT 39.824 5.004 39.856 7.512 ;
  LAYER M3 ;
        RECT 39.824 7.46 39.856 7.492 ;
  LAYER M1 ;
        RECT 39.76 5.004 39.792 7.512 ;
  LAYER M3 ;
        RECT 39.76 5.024 39.792 5.056 ;
  LAYER M1 ;
        RECT 39.696 5.004 39.728 7.512 ;
  LAYER M3 ;
        RECT 39.696 7.46 39.728 7.492 ;
  LAYER M1 ;
        RECT 39.632 5.004 39.664 7.512 ;
  LAYER M3 ;
        RECT 39.632 5.024 39.664 5.056 ;
  LAYER M1 ;
        RECT 39.568 5.004 39.6 7.512 ;
  LAYER M3 ;
        RECT 39.568 7.46 39.6 7.492 ;
  LAYER M1 ;
        RECT 39.504 5.004 39.536 7.512 ;
  LAYER M3 ;
        RECT 39.504 5.024 39.536 5.056 ;
  LAYER M1 ;
        RECT 39.44 5.004 39.472 7.512 ;
  LAYER M3 ;
        RECT 39.44 7.46 39.472 7.492 ;
  LAYER M1 ;
        RECT 39.376 5.004 39.408 7.512 ;
  LAYER M3 ;
        RECT 39.376 5.024 39.408 5.056 ;
  LAYER M1 ;
        RECT 39.312 5.004 39.344 7.512 ;
  LAYER M3 ;
        RECT 39.312 7.46 39.344 7.492 ;
  LAYER M1 ;
        RECT 39.248 5.004 39.28 7.512 ;
  LAYER M3 ;
        RECT 39.248 5.024 39.28 5.056 ;
  LAYER M1 ;
        RECT 39.184 5.004 39.216 7.512 ;
  LAYER M3 ;
        RECT 39.184 7.46 39.216 7.492 ;
  LAYER M1 ;
        RECT 39.12 5.004 39.152 7.512 ;
  LAYER M3 ;
        RECT 39.12 5.024 39.152 5.056 ;
  LAYER M1 ;
        RECT 39.056 5.004 39.088 7.512 ;
  LAYER M3 ;
        RECT 39.056 7.46 39.088 7.492 ;
  LAYER M1 ;
        RECT 38.992 5.004 39.024 7.512 ;
  LAYER M3 ;
        RECT 38.992 5.024 39.024 5.056 ;
  LAYER M1 ;
        RECT 38.928 5.004 38.96 7.512 ;
  LAYER M3 ;
        RECT 38.928 7.46 38.96 7.492 ;
  LAYER M1 ;
        RECT 38.864 5.004 38.896 7.512 ;
  LAYER M3 ;
        RECT 38.864 5.024 38.896 5.056 ;
  LAYER M1 ;
        RECT 38.8 5.004 38.832 7.512 ;
  LAYER M3 ;
        RECT 38.8 7.46 38.832 7.492 ;
  LAYER M1 ;
        RECT 38.736 5.004 38.768 7.512 ;
  LAYER M3 ;
        RECT 38.736 5.024 38.768 5.056 ;
  LAYER M1 ;
        RECT 38.672 5.004 38.704 7.512 ;
  LAYER M3 ;
        RECT 38.672 7.46 38.704 7.492 ;
  LAYER M1 ;
        RECT 38.608 5.004 38.64 7.512 ;
  LAYER M3 ;
        RECT 38.608 5.024 38.64 5.056 ;
  LAYER M1 ;
        RECT 38.544 5.004 38.576 7.512 ;
  LAYER M3 ;
        RECT 38.544 7.46 38.576 7.492 ;
  LAYER M1 ;
        RECT 38.48 5.004 38.512 7.512 ;
  LAYER M3 ;
        RECT 40.848 5.088 40.88 5.12 ;
  LAYER M2 ;
        RECT 38.48 5.152 38.512 5.184 ;
  LAYER M2 ;
        RECT 40.848 5.216 40.88 5.248 ;
  LAYER M2 ;
        RECT 38.48 5.28 38.512 5.312 ;
  LAYER M2 ;
        RECT 40.848 5.344 40.88 5.376 ;
  LAYER M2 ;
        RECT 38.48 5.408 38.512 5.44 ;
  LAYER M2 ;
        RECT 40.848 5.472 40.88 5.504 ;
  LAYER M2 ;
        RECT 38.48 5.536 38.512 5.568 ;
  LAYER M2 ;
        RECT 40.848 5.6 40.88 5.632 ;
  LAYER M2 ;
        RECT 38.48 5.664 38.512 5.696 ;
  LAYER M2 ;
        RECT 40.848 5.728 40.88 5.76 ;
  LAYER M2 ;
        RECT 38.48 5.792 38.512 5.824 ;
  LAYER M2 ;
        RECT 40.848 5.856 40.88 5.888 ;
  LAYER M2 ;
        RECT 38.48 5.92 38.512 5.952 ;
  LAYER M2 ;
        RECT 40.848 5.984 40.88 6.016 ;
  LAYER M2 ;
        RECT 38.48 6.048 38.512 6.08 ;
  LAYER M2 ;
        RECT 40.848 6.112 40.88 6.144 ;
  LAYER M2 ;
        RECT 38.48 6.176 38.512 6.208 ;
  LAYER M2 ;
        RECT 40.848 6.24 40.88 6.272 ;
  LAYER M2 ;
        RECT 38.48 6.304 38.512 6.336 ;
  LAYER M2 ;
        RECT 40.848 6.368 40.88 6.4 ;
  LAYER M2 ;
        RECT 38.48 6.432 38.512 6.464 ;
  LAYER M2 ;
        RECT 40.848 6.496 40.88 6.528 ;
  LAYER M2 ;
        RECT 38.48 6.56 38.512 6.592 ;
  LAYER M2 ;
        RECT 40.848 6.624 40.88 6.656 ;
  LAYER M2 ;
        RECT 38.48 6.688 38.512 6.72 ;
  LAYER M2 ;
        RECT 40.848 6.752 40.88 6.784 ;
  LAYER M2 ;
        RECT 38.48 6.816 38.512 6.848 ;
  LAYER M2 ;
        RECT 40.848 6.88 40.88 6.912 ;
  LAYER M2 ;
        RECT 38.48 6.944 38.512 6.976 ;
  LAYER M2 ;
        RECT 40.848 7.008 40.88 7.04 ;
  LAYER M2 ;
        RECT 38.48 7.072 38.512 7.104 ;
  LAYER M2 ;
        RECT 40.848 7.136 40.88 7.168 ;
  LAYER M2 ;
        RECT 38.48 7.2 38.512 7.232 ;
  LAYER M2 ;
        RECT 40.848 7.264 40.88 7.296 ;
  LAYER M2 ;
        RECT 38.48 7.328 38.512 7.36 ;
  LAYER M2 ;
        RECT 38.432 4.956 40.928 7.56 ;
  LAYER M1 ;
        RECT 40.848 8.112 40.88 10.62 ;
  LAYER M3 ;
        RECT 40.848 10.568 40.88 10.6 ;
  LAYER M1 ;
        RECT 40.784 8.112 40.816 10.62 ;
  LAYER M3 ;
        RECT 40.784 8.132 40.816 8.164 ;
  LAYER M1 ;
        RECT 40.72 8.112 40.752 10.62 ;
  LAYER M3 ;
        RECT 40.72 10.568 40.752 10.6 ;
  LAYER M1 ;
        RECT 40.656 8.112 40.688 10.62 ;
  LAYER M3 ;
        RECT 40.656 8.132 40.688 8.164 ;
  LAYER M1 ;
        RECT 40.592 8.112 40.624 10.62 ;
  LAYER M3 ;
        RECT 40.592 10.568 40.624 10.6 ;
  LAYER M1 ;
        RECT 40.528 8.112 40.56 10.62 ;
  LAYER M3 ;
        RECT 40.528 8.132 40.56 8.164 ;
  LAYER M1 ;
        RECT 40.464 8.112 40.496 10.62 ;
  LAYER M3 ;
        RECT 40.464 10.568 40.496 10.6 ;
  LAYER M1 ;
        RECT 40.4 8.112 40.432 10.62 ;
  LAYER M3 ;
        RECT 40.4 8.132 40.432 8.164 ;
  LAYER M1 ;
        RECT 40.336 8.112 40.368 10.62 ;
  LAYER M3 ;
        RECT 40.336 10.568 40.368 10.6 ;
  LAYER M1 ;
        RECT 40.272 8.112 40.304 10.62 ;
  LAYER M3 ;
        RECT 40.272 8.132 40.304 8.164 ;
  LAYER M1 ;
        RECT 40.208 8.112 40.24 10.62 ;
  LAYER M3 ;
        RECT 40.208 10.568 40.24 10.6 ;
  LAYER M1 ;
        RECT 40.144 8.112 40.176 10.62 ;
  LAYER M3 ;
        RECT 40.144 8.132 40.176 8.164 ;
  LAYER M1 ;
        RECT 40.08 8.112 40.112 10.62 ;
  LAYER M3 ;
        RECT 40.08 10.568 40.112 10.6 ;
  LAYER M1 ;
        RECT 40.016 8.112 40.048 10.62 ;
  LAYER M3 ;
        RECT 40.016 8.132 40.048 8.164 ;
  LAYER M1 ;
        RECT 39.952 8.112 39.984 10.62 ;
  LAYER M3 ;
        RECT 39.952 10.568 39.984 10.6 ;
  LAYER M1 ;
        RECT 39.888 8.112 39.92 10.62 ;
  LAYER M3 ;
        RECT 39.888 8.132 39.92 8.164 ;
  LAYER M1 ;
        RECT 39.824 8.112 39.856 10.62 ;
  LAYER M3 ;
        RECT 39.824 10.568 39.856 10.6 ;
  LAYER M1 ;
        RECT 39.76 8.112 39.792 10.62 ;
  LAYER M3 ;
        RECT 39.76 8.132 39.792 8.164 ;
  LAYER M1 ;
        RECT 39.696 8.112 39.728 10.62 ;
  LAYER M3 ;
        RECT 39.696 10.568 39.728 10.6 ;
  LAYER M1 ;
        RECT 39.632 8.112 39.664 10.62 ;
  LAYER M3 ;
        RECT 39.632 8.132 39.664 8.164 ;
  LAYER M1 ;
        RECT 39.568 8.112 39.6 10.62 ;
  LAYER M3 ;
        RECT 39.568 10.568 39.6 10.6 ;
  LAYER M1 ;
        RECT 39.504 8.112 39.536 10.62 ;
  LAYER M3 ;
        RECT 39.504 8.132 39.536 8.164 ;
  LAYER M1 ;
        RECT 39.44 8.112 39.472 10.62 ;
  LAYER M3 ;
        RECT 39.44 10.568 39.472 10.6 ;
  LAYER M1 ;
        RECT 39.376 8.112 39.408 10.62 ;
  LAYER M3 ;
        RECT 39.376 8.132 39.408 8.164 ;
  LAYER M1 ;
        RECT 39.312 8.112 39.344 10.62 ;
  LAYER M3 ;
        RECT 39.312 10.568 39.344 10.6 ;
  LAYER M1 ;
        RECT 39.248 8.112 39.28 10.62 ;
  LAYER M3 ;
        RECT 39.248 8.132 39.28 8.164 ;
  LAYER M1 ;
        RECT 39.184 8.112 39.216 10.62 ;
  LAYER M3 ;
        RECT 39.184 10.568 39.216 10.6 ;
  LAYER M1 ;
        RECT 39.12 8.112 39.152 10.62 ;
  LAYER M3 ;
        RECT 39.12 8.132 39.152 8.164 ;
  LAYER M1 ;
        RECT 39.056 8.112 39.088 10.62 ;
  LAYER M3 ;
        RECT 39.056 10.568 39.088 10.6 ;
  LAYER M1 ;
        RECT 38.992 8.112 39.024 10.62 ;
  LAYER M3 ;
        RECT 38.992 8.132 39.024 8.164 ;
  LAYER M1 ;
        RECT 38.928 8.112 38.96 10.62 ;
  LAYER M3 ;
        RECT 38.928 10.568 38.96 10.6 ;
  LAYER M1 ;
        RECT 38.864 8.112 38.896 10.62 ;
  LAYER M3 ;
        RECT 38.864 8.132 38.896 8.164 ;
  LAYER M1 ;
        RECT 38.8 8.112 38.832 10.62 ;
  LAYER M3 ;
        RECT 38.8 10.568 38.832 10.6 ;
  LAYER M1 ;
        RECT 38.736 8.112 38.768 10.62 ;
  LAYER M3 ;
        RECT 38.736 8.132 38.768 8.164 ;
  LAYER M1 ;
        RECT 38.672 8.112 38.704 10.62 ;
  LAYER M3 ;
        RECT 38.672 10.568 38.704 10.6 ;
  LAYER M1 ;
        RECT 38.608 8.112 38.64 10.62 ;
  LAYER M3 ;
        RECT 38.608 8.132 38.64 8.164 ;
  LAYER M1 ;
        RECT 38.544 8.112 38.576 10.62 ;
  LAYER M3 ;
        RECT 38.544 10.568 38.576 10.6 ;
  LAYER M1 ;
        RECT 38.48 8.112 38.512 10.62 ;
  LAYER M3 ;
        RECT 40.848 8.196 40.88 8.228 ;
  LAYER M2 ;
        RECT 38.48 8.26 38.512 8.292 ;
  LAYER M2 ;
        RECT 40.848 8.324 40.88 8.356 ;
  LAYER M2 ;
        RECT 38.48 8.388 38.512 8.42 ;
  LAYER M2 ;
        RECT 40.848 8.452 40.88 8.484 ;
  LAYER M2 ;
        RECT 38.48 8.516 38.512 8.548 ;
  LAYER M2 ;
        RECT 40.848 8.58 40.88 8.612 ;
  LAYER M2 ;
        RECT 38.48 8.644 38.512 8.676 ;
  LAYER M2 ;
        RECT 40.848 8.708 40.88 8.74 ;
  LAYER M2 ;
        RECT 38.48 8.772 38.512 8.804 ;
  LAYER M2 ;
        RECT 40.848 8.836 40.88 8.868 ;
  LAYER M2 ;
        RECT 38.48 8.9 38.512 8.932 ;
  LAYER M2 ;
        RECT 40.848 8.964 40.88 8.996 ;
  LAYER M2 ;
        RECT 38.48 9.028 38.512 9.06 ;
  LAYER M2 ;
        RECT 40.848 9.092 40.88 9.124 ;
  LAYER M2 ;
        RECT 38.48 9.156 38.512 9.188 ;
  LAYER M2 ;
        RECT 40.848 9.22 40.88 9.252 ;
  LAYER M2 ;
        RECT 38.48 9.284 38.512 9.316 ;
  LAYER M2 ;
        RECT 40.848 9.348 40.88 9.38 ;
  LAYER M2 ;
        RECT 38.48 9.412 38.512 9.444 ;
  LAYER M2 ;
        RECT 40.848 9.476 40.88 9.508 ;
  LAYER M2 ;
        RECT 38.48 9.54 38.512 9.572 ;
  LAYER M2 ;
        RECT 40.848 9.604 40.88 9.636 ;
  LAYER M2 ;
        RECT 38.48 9.668 38.512 9.7 ;
  LAYER M2 ;
        RECT 40.848 9.732 40.88 9.764 ;
  LAYER M2 ;
        RECT 38.48 9.796 38.512 9.828 ;
  LAYER M2 ;
        RECT 40.848 9.86 40.88 9.892 ;
  LAYER M2 ;
        RECT 38.48 9.924 38.512 9.956 ;
  LAYER M2 ;
        RECT 40.848 9.988 40.88 10.02 ;
  LAYER M2 ;
        RECT 38.48 10.052 38.512 10.084 ;
  LAYER M2 ;
        RECT 40.848 10.116 40.88 10.148 ;
  LAYER M2 ;
        RECT 38.48 10.18 38.512 10.212 ;
  LAYER M2 ;
        RECT 40.848 10.244 40.88 10.276 ;
  LAYER M2 ;
        RECT 38.48 10.308 38.512 10.34 ;
  LAYER M2 ;
        RECT 40.848 10.372 40.88 10.404 ;
  LAYER M2 ;
        RECT 38.48 10.436 38.512 10.468 ;
  LAYER M2 ;
        RECT 38.432 8.064 40.928 10.668 ;
  LAYER M1 ;
        RECT 40.848 11.22 40.88 13.728 ;
  LAYER M3 ;
        RECT 40.848 13.676 40.88 13.708 ;
  LAYER M1 ;
        RECT 40.784 11.22 40.816 13.728 ;
  LAYER M3 ;
        RECT 40.784 11.24 40.816 11.272 ;
  LAYER M1 ;
        RECT 40.72 11.22 40.752 13.728 ;
  LAYER M3 ;
        RECT 40.72 13.676 40.752 13.708 ;
  LAYER M1 ;
        RECT 40.656 11.22 40.688 13.728 ;
  LAYER M3 ;
        RECT 40.656 11.24 40.688 11.272 ;
  LAYER M1 ;
        RECT 40.592 11.22 40.624 13.728 ;
  LAYER M3 ;
        RECT 40.592 13.676 40.624 13.708 ;
  LAYER M1 ;
        RECT 40.528 11.22 40.56 13.728 ;
  LAYER M3 ;
        RECT 40.528 11.24 40.56 11.272 ;
  LAYER M1 ;
        RECT 40.464 11.22 40.496 13.728 ;
  LAYER M3 ;
        RECT 40.464 13.676 40.496 13.708 ;
  LAYER M1 ;
        RECT 40.4 11.22 40.432 13.728 ;
  LAYER M3 ;
        RECT 40.4 11.24 40.432 11.272 ;
  LAYER M1 ;
        RECT 40.336 11.22 40.368 13.728 ;
  LAYER M3 ;
        RECT 40.336 13.676 40.368 13.708 ;
  LAYER M1 ;
        RECT 40.272 11.22 40.304 13.728 ;
  LAYER M3 ;
        RECT 40.272 11.24 40.304 11.272 ;
  LAYER M1 ;
        RECT 40.208 11.22 40.24 13.728 ;
  LAYER M3 ;
        RECT 40.208 13.676 40.24 13.708 ;
  LAYER M1 ;
        RECT 40.144 11.22 40.176 13.728 ;
  LAYER M3 ;
        RECT 40.144 11.24 40.176 11.272 ;
  LAYER M1 ;
        RECT 40.08 11.22 40.112 13.728 ;
  LAYER M3 ;
        RECT 40.08 13.676 40.112 13.708 ;
  LAYER M1 ;
        RECT 40.016 11.22 40.048 13.728 ;
  LAYER M3 ;
        RECT 40.016 11.24 40.048 11.272 ;
  LAYER M1 ;
        RECT 39.952 11.22 39.984 13.728 ;
  LAYER M3 ;
        RECT 39.952 13.676 39.984 13.708 ;
  LAYER M1 ;
        RECT 39.888 11.22 39.92 13.728 ;
  LAYER M3 ;
        RECT 39.888 11.24 39.92 11.272 ;
  LAYER M1 ;
        RECT 39.824 11.22 39.856 13.728 ;
  LAYER M3 ;
        RECT 39.824 13.676 39.856 13.708 ;
  LAYER M1 ;
        RECT 39.76 11.22 39.792 13.728 ;
  LAYER M3 ;
        RECT 39.76 11.24 39.792 11.272 ;
  LAYER M1 ;
        RECT 39.696 11.22 39.728 13.728 ;
  LAYER M3 ;
        RECT 39.696 13.676 39.728 13.708 ;
  LAYER M1 ;
        RECT 39.632 11.22 39.664 13.728 ;
  LAYER M3 ;
        RECT 39.632 11.24 39.664 11.272 ;
  LAYER M1 ;
        RECT 39.568 11.22 39.6 13.728 ;
  LAYER M3 ;
        RECT 39.568 13.676 39.6 13.708 ;
  LAYER M1 ;
        RECT 39.504 11.22 39.536 13.728 ;
  LAYER M3 ;
        RECT 39.504 11.24 39.536 11.272 ;
  LAYER M1 ;
        RECT 39.44 11.22 39.472 13.728 ;
  LAYER M3 ;
        RECT 39.44 13.676 39.472 13.708 ;
  LAYER M1 ;
        RECT 39.376 11.22 39.408 13.728 ;
  LAYER M3 ;
        RECT 39.376 11.24 39.408 11.272 ;
  LAYER M1 ;
        RECT 39.312 11.22 39.344 13.728 ;
  LAYER M3 ;
        RECT 39.312 13.676 39.344 13.708 ;
  LAYER M1 ;
        RECT 39.248 11.22 39.28 13.728 ;
  LAYER M3 ;
        RECT 39.248 11.24 39.28 11.272 ;
  LAYER M1 ;
        RECT 39.184 11.22 39.216 13.728 ;
  LAYER M3 ;
        RECT 39.184 13.676 39.216 13.708 ;
  LAYER M1 ;
        RECT 39.12 11.22 39.152 13.728 ;
  LAYER M3 ;
        RECT 39.12 11.24 39.152 11.272 ;
  LAYER M1 ;
        RECT 39.056 11.22 39.088 13.728 ;
  LAYER M3 ;
        RECT 39.056 13.676 39.088 13.708 ;
  LAYER M1 ;
        RECT 38.992 11.22 39.024 13.728 ;
  LAYER M3 ;
        RECT 38.992 11.24 39.024 11.272 ;
  LAYER M1 ;
        RECT 38.928 11.22 38.96 13.728 ;
  LAYER M3 ;
        RECT 38.928 13.676 38.96 13.708 ;
  LAYER M1 ;
        RECT 38.864 11.22 38.896 13.728 ;
  LAYER M3 ;
        RECT 38.864 11.24 38.896 11.272 ;
  LAYER M1 ;
        RECT 38.8 11.22 38.832 13.728 ;
  LAYER M3 ;
        RECT 38.8 13.676 38.832 13.708 ;
  LAYER M1 ;
        RECT 38.736 11.22 38.768 13.728 ;
  LAYER M3 ;
        RECT 38.736 11.24 38.768 11.272 ;
  LAYER M1 ;
        RECT 38.672 11.22 38.704 13.728 ;
  LAYER M3 ;
        RECT 38.672 13.676 38.704 13.708 ;
  LAYER M1 ;
        RECT 38.608 11.22 38.64 13.728 ;
  LAYER M3 ;
        RECT 38.608 11.24 38.64 11.272 ;
  LAYER M1 ;
        RECT 38.544 11.22 38.576 13.728 ;
  LAYER M3 ;
        RECT 38.544 13.676 38.576 13.708 ;
  LAYER M1 ;
        RECT 38.48 11.22 38.512 13.728 ;
  LAYER M3 ;
        RECT 40.848 11.304 40.88 11.336 ;
  LAYER M2 ;
        RECT 38.48 11.368 38.512 11.4 ;
  LAYER M2 ;
        RECT 40.848 11.432 40.88 11.464 ;
  LAYER M2 ;
        RECT 38.48 11.496 38.512 11.528 ;
  LAYER M2 ;
        RECT 40.848 11.56 40.88 11.592 ;
  LAYER M2 ;
        RECT 38.48 11.624 38.512 11.656 ;
  LAYER M2 ;
        RECT 40.848 11.688 40.88 11.72 ;
  LAYER M2 ;
        RECT 38.48 11.752 38.512 11.784 ;
  LAYER M2 ;
        RECT 40.848 11.816 40.88 11.848 ;
  LAYER M2 ;
        RECT 38.48 11.88 38.512 11.912 ;
  LAYER M2 ;
        RECT 40.848 11.944 40.88 11.976 ;
  LAYER M2 ;
        RECT 38.48 12.008 38.512 12.04 ;
  LAYER M2 ;
        RECT 40.848 12.072 40.88 12.104 ;
  LAYER M2 ;
        RECT 38.48 12.136 38.512 12.168 ;
  LAYER M2 ;
        RECT 40.848 12.2 40.88 12.232 ;
  LAYER M2 ;
        RECT 38.48 12.264 38.512 12.296 ;
  LAYER M2 ;
        RECT 40.848 12.328 40.88 12.36 ;
  LAYER M2 ;
        RECT 38.48 12.392 38.512 12.424 ;
  LAYER M2 ;
        RECT 40.848 12.456 40.88 12.488 ;
  LAYER M2 ;
        RECT 38.48 12.52 38.512 12.552 ;
  LAYER M2 ;
        RECT 40.848 12.584 40.88 12.616 ;
  LAYER M2 ;
        RECT 38.48 12.648 38.512 12.68 ;
  LAYER M2 ;
        RECT 40.848 12.712 40.88 12.744 ;
  LAYER M2 ;
        RECT 38.48 12.776 38.512 12.808 ;
  LAYER M2 ;
        RECT 40.848 12.84 40.88 12.872 ;
  LAYER M2 ;
        RECT 38.48 12.904 38.512 12.936 ;
  LAYER M2 ;
        RECT 40.848 12.968 40.88 13 ;
  LAYER M2 ;
        RECT 38.48 13.032 38.512 13.064 ;
  LAYER M2 ;
        RECT 40.848 13.096 40.88 13.128 ;
  LAYER M2 ;
        RECT 38.48 13.16 38.512 13.192 ;
  LAYER M2 ;
        RECT 40.848 13.224 40.88 13.256 ;
  LAYER M2 ;
        RECT 38.48 13.288 38.512 13.32 ;
  LAYER M2 ;
        RECT 40.848 13.352 40.88 13.384 ;
  LAYER M2 ;
        RECT 38.48 13.416 38.512 13.448 ;
  LAYER M2 ;
        RECT 40.848 13.48 40.88 13.512 ;
  LAYER M2 ;
        RECT 38.48 13.544 38.512 13.576 ;
  LAYER M2 ;
        RECT 38.432 11.172 40.928 13.776 ;
  LAYER M1 ;
        RECT 37.872 1.896 37.904 4.404 ;
  LAYER M3 ;
        RECT 37.872 4.352 37.904 4.384 ;
  LAYER M1 ;
        RECT 37.808 1.896 37.84 4.404 ;
  LAYER M3 ;
        RECT 37.808 1.916 37.84 1.948 ;
  LAYER M1 ;
        RECT 37.744 1.896 37.776 4.404 ;
  LAYER M3 ;
        RECT 37.744 4.352 37.776 4.384 ;
  LAYER M1 ;
        RECT 37.68 1.896 37.712 4.404 ;
  LAYER M3 ;
        RECT 37.68 1.916 37.712 1.948 ;
  LAYER M1 ;
        RECT 37.616 1.896 37.648 4.404 ;
  LAYER M3 ;
        RECT 37.616 4.352 37.648 4.384 ;
  LAYER M1 ;
        RECT 37.552 1.896 37.584 4.404 ;
  LAYER M3 ;
        RECT 37.552 1.916 37.584 1.948 ;
  LAYER M1 ;
        RECT 37.488 1.896 37.52 4.404 ;
  LAYER M3 ;
        RECT 37.488 4.352 37.52 4.384 ;
  LAYER M1 ;
        RECT 37.424 1.896 37.456 4.404 ;
  LAYER M3 ;
        RECT 37.424 1.916 37.456 1.948 ;
  LAYER M1 ;
        RECT 37.36 1.896 37.392 4.404 ;
  LAYER M3 ;
        RECT 37.36 4.352 37.392 4.384 ;
  LAYER M1 ;
        RECT 37.296 1.896 37.328 4.404 ;
  LAYER M3 ;
        RECT 37.296 1.916 37.328 1.948 ;
  LAYER M1 ;
        RECT 37.232 1.896 37.264 4.404 ;
  LAYER M3 ;
        RECT 37.232 4.352 37.264 4.384 ;
  LAYER M1 ;
        RECT 37.168 1.896 37.2 4.404 ;
  LAYER M3 ;
        RECT 37.168 1.916 37.2 1.948 ;
  LAYER M1 ;
        RECT 37.104 1.896 37.136 4.404 ;
  LAYER M3 ;
        RECT 37.104 4.352 37.136 4.384 ;
  LAYER M1 ;
        RECT 37.04 1.896 37.072 4.404 ;
  LAYER M3 ;
        RECT 37.04 1.916 37.072 1.948 ;
  LAYER M1 ;
        RECT 36.976 1.896 37.008 4.404 ;
  LAYER M3 ;
        RECT 36.976 4.352 37.008 4.384 ;
  LAYER M1 ;
        RECT 36.912 1.896 36.944 4.404 ;
  LAYER M3 ;
        RECT 36.912 1.916 36.944 1.948 ;
  LAYER M1 ;
        RECT 36.848 1.896 36.88 4.404 ;
  LAYER M3 ;
        RECT 36.848 4.352 36.88 4.384 ;
  LAYER M1 ;
        RECT 36.784 1.896 36.816 4.404 ;
  LAYER M3 ;
        RECT 36.784 1.916 36.816 1.948 ;
  LAYER M1 ;
        RECT 36.72 1.896 36.752 4.404 ;
  LAYER M3 ;
        RECT 36.72 4.352 36.752 4.384 ;
  LAYER M1 ;
        RECT 36.656 1.896 36.688 4.404 ;
  LAYER M3 ;
        RECT 36.656 1.916 36.688 1.948 ;
  LAYER M1 ;
        RECT 36.592 1.896 36.624 4.404 ;
  LAYER M3 ;
        RECT 36.592 4.352 36.624 4.384 ;
  LAYER M1 ;
        RECT 36.528 1.896 36.56 4.404 ;
  LAYER M3 ;
        RECT 36.528 1.916 36.56 1.948 ;
  LAYER M1 ;
        RECT 36.464 1.896 36.496 4.404 ;
  LAYER M3 ;
        RECT 36.464 4.352 36.496 4.384 ;
  LAYER M1 ;
        RECT 36.4 1.896 36.432 4.404 ;
  LAYER M3 ;
        RECT 36.4 1.916 36.432 1.948 ;
  LAYER M1 ;
        RECT 36.336 1.896 36.368 4.404 ;
  LAYER M3 ;
        RECT 36.336 4.352 36.368 4.384 ;
  LAYER M1 ;
        RECT 36.272 1.896 36.304 4.404 ;
  LAYER M3 ;
        RECT 36.272 1.916 36.304 1.948 ;
  LAYER M1 ;
        RECT 36.208 1.896 36.24 4.404 ;
  LAYER M3 ;
        RECT 36.208 4.352 36.24 4.384 ;
  LAYER M1 ;
        RECT 36.144 1.896 36.176 4.404 ;
  LAYER M3 ;
        RECT 36.144 1.916 36.176 1.948 ;
  LAYER M1 ;
        RECT 36.08 1.896 36.112 4.404 ;
  LAYER M3 ;
        RECT 36.08 4.352 36.112 4.384 ;
  LAYER M1 ;
        RECT 36.016 1.896 36.048 4.404 ;
  LAYER M3 ;
        RECT 36.016 1.916 36.048 1.948 ;
  LAYER M1 ;
        RECT 35.952 1.896 35.984 4.404 ;
  LAYER M3 ;
        RECT 35.952 4.352 35.984 4.384 ;
  LAYER M1 ;
        RECT 35.888 1.896 35.92 4.404 ;
  LAYER M3 ;
        RECT 35.888 1.916 35.92 1.948 ;
  LAYER M1 ;
        RECT 35.824 1.896 35.856 4.404 ;
  LAYER M3 ;
        RECT 35.824 4.352 35.856 4.384 ;
  LAYER M1 ;
        RECT 35.76 1.896 35.792 4.404 ;
  LAYER M3 ;
        RECT 35.76 1.916 35.792 1.948 ;
  LAYER M1 ;
        RECT 35.696 1.896 35.728 4.404 ;
  LAYER M3 ;
        RECT 35.696 4.352 35.728 4.384 ;
  LAYER M1 ;
        RECT 35.632 1.896 35.664 4.404 ;
  LAYER M3 ;
        RECT 35.632 1.916 35.664 1.948 ;
  LAYER M1 ;
        RECT 35.568 1.896 35.6 4.404 ;
  LAYER M3 ;
        RECT 35.568 4.352 35.6 4.384 ;
  LAYER M1 ;
        RECT 35.504 1.896 35.536 4.404 ;
  LAYER M3 ;
        RECT 37.872 1.98 37.904 2.012 ;
  LAYER M2 ;
        RECT 35.504 2.044 35.536 2.076 ;
  LAYER M2 ;
        RECT 37.872 2.108 37.904 2.14 ;
  LAYER M2 ;
        RECT 35.504 2.172 35.536 2.204 ;
  LAYER M2 ;
        RECT 37.872 2.236 37.904 2.268 ;
  LAYER M2 ;
        RECT 35.504 2.3 35.536 2.332 ;
  LAYER M2 ;
        RECT 37.872 2.364 37.904 2.396 ;
  LAYER M2 ;
        RECT 35.504 2.428 35.536 2.46 ;
  LAYER M2 ;
        RECT 37.872 2.492 37.904 2.524 ;
  LAYER M2 ;
        RECT 35.504 2.556 35.536 2.588 ;
  LAYER M2 ;
        RECT 37.872 2.62 37.904 2.652 ;
  LAYER M2 ;
        RECT 35.504 2.684 35.536 2.716 ;
  LAYER M2 ;
        RECT 37.872 2.748 37.904 2.78 ;
  LAYER M2 ;
        RECT 35.504 2.812 35.536 2.844 ;
  LAYER M2 ;
        RECT 37.872 2.876 37.904 2.908 ;
  LAYER M2 ;
        RECT 35.504 2.94 35.536 2.972 ;
  LAYER M2 ;
        RECT 37.872 3.004 37.904 3.036 ;
  LAYER M2 ;
        RECT 35.504 3.068 35.536 3.1 ;
  LAYER M2 ;
        RECT 37.872 3.132 37.904 3.164 ;
  LAYER M2 ;
        RECT 35.504 3.196 35.536 3.228 ;
  LAYER M2 ;
        RECT 37.872 3.26 37.904 3.292 ;
  LAYER M2 ;
        RECT 35.504 3.324 35.536 3.356 ;
  LAYER M2 ;
        RECT 37.872 3.388 37.904 3.42 ;
  LAYER M2 ;
        RECT 35.504 3.452 35.536 3.484 ;
  LAYER M2 ;
        RECT 37.872 3.516 37.904 3.548 ;
  LAYER M2 ;
        RECT 35.504 3.58 35.536 3.612 ;
  LAYER M2 ;
        RECT 37.872 3.644 37.904 3.676 ;
  LAYER M2 ;
        RECT 35.504 3.708 35.536 3.74 ;
  LAYER M2 ;
        RECT 37.872 3.772 37.904 3.804 ;
  LAYER M2 ;
        RECT 35.504 3.836 35.536 3.868 ;
  LAYER M2 ;
        RECT 37.872 3.9 37.904 3.932 ;
  LAYER M2 ;
        RECT 35.504 3.964 35.536 3.996 ;
  LAYER M2 ;
        RECT 37.872 4.028 37.904 4.06 ;
  LAYER M2 ;
        RECT 35.504 4.092 35.536 4.124 ;
  LAYER M2 ;
        RECT 37.872 4.156 37.904 4.188 ;
  LAYER M2 ;
        RECT 35.504 4.22 35.536 4.252 ;
  LAYER M2 ;
        RECT 35.456 1.848 37.952 4.452 ;
  LAYER M1 ;
        RECT 37.872 5.004 37.904 7.512 ;
  LAYER M3 ;
        RECT 37.872 7.46 37.904 7.492 ;
  LAYER M1 ;
        RECT 37.808 5.004 37.84 7.512 ;
  LAYER M3 ;
        RECT 37.808 5.024 37.84 5.056 ;
  LAYER M1 ;
        RECT 37.744 5.004 37.776 7.512 ;
  LAYER M3 ;
        RECT 37.744 7.46 37.776 7.492 ;
  LAYER M1 ;
        RECT 37.68 5.004 37.712 7.512 ;
  LAYER M3 ;
        RECT 37.68 5.024 37.712 5.056 ;
  LAYER M1 ;
        RECT 37.616 5.004 37.648 7.512 ;
  LAYER M3 ;
        RECT 37.616 7.46 37.648 7.492 ;
  LAYER M1 ;
        RECT 37.552 5.004 37.584 7.512 ;
  LAYER M3 ;
        RECT 37.552 5.024 37.584 5.056 ;
  LAYER M1 ;
        RECT 37.488 5.004 37.52 7.512 ;
  LAYER M3 ;
        RECT 37.488 7.46 37.52 7.492 ;
  LAYER M1 ;
        RECT 37.424 5.004 37.456 7.512 ;
  LAYER M3 ;
        RECT 37.424 5.024 37.456 5.056 ;
  LAYER M1 ;
        RECT 37.36 5.004 37.392 7.512 ;
  LAYER M3 ;
        RECT 37.36 7.46 37.392 7.492 ;
  LAYER M1 ;
        RECT 37.296 5.004 37.328 7.512 ;
  LAYER M3 ;
        RECT 37.296 5.024 37.328 5.056 ;
  LAYER M1 ;
        RECT 37.232 5.004 37.264 7.512 ;
  LAYER M3 ;
        RECT 37.232 7.46 37.264 7.492 ;
  LAYER M1 ;
        RECT 37.168 5.004 37.2 7.512 ;
  LAYER M3 ;
        RECT 37.168 5.024 37.2 5.056 ;
  LAYER M1 ;
        RECT 37.104 5.004 37.136 7.512 ;
  LAYER M3 ;
        RECT 37.104 7.46 37.136 7.492 ;
  LAYER M1 ;
        RECT 37.04 5.004 37.072 7.512 ;
  LAYER M3 ;
        RECT 37.04 5.024 37.072 5.056 ;
  LAYER M1 ;
        RECT 36.976 5.004 37.008 7.512 ;
  LAYER M3 ;
        RECT 36.976 7.46 37.008 7.492 ;
  LAYER M1 ;
        RECT 36.912 5.004 36.944 7.512 ;
  LAYER M3 ;
        RECT 36.912 5.024 36.944 5.056 ;
  LAYER M1 ;
        RECT 36.848 5.004 36.88 7.512 ;
  LAYER M3 ;
        RECT 36.848 7.46 36.88 7.492 ;
  LAYER M1 ;
        RECT 36.784 5.004 36.816 7.512 ;
  LAYER M3 ;
        RECT 36.784 5.024 36.816 5.056 ;
  LAYER M1 ;
        RECT 36.72 5.004 36.752 7.512 ;
  LAYER M3 ;
        RECT 36.72 7.46 36.752 7.492 ;
  LAYER M1 ;
        RECT 36.656 5.004 36.688 7.512 ;
  LAYER M3 ;
        RECT 36.656 5.024 36.688 5.056 ;
  LAYER M1 ;
        RECT 36.592 5.004 36.624 7.512 ;
  LAYER M3 ;
        RECT 36.592 7.46 36.624 7.492 ;
  LAYER M1 ;
        RECT 36.528 5.004 36.56 7.512 ;
  LAYER M3 ;
        RECT 36.528 5.024 36.56 5.056 ;
  LAYER M1 ;
        RECT 36.464 5.004 36.496 7.512 ;
  LAYER M3 ;
        RECT 36.464 7.46 36.496 7.492 ;
  LAYER M1 ;
        RECT 36.4 5.004 36.432 7.512 ;
  LAYER M3 ;
        RECT 36.4 5.024 36.432 5.056 ;
  LAYER M1 ;
        RECT 36.336 5.004 36.368 7.512 ;
  LAYER M3 ;
        RECT 36.336 7.46 36.368 7.492 ;
  LAYER M1 ;
        RECT 36.272 5.004 36.304 7.512 ;
  LAYER M3 ;
        RECT 36.272 5.024 36.304 5.056 ;
  LAYER M1 ;
        RECT 36.208 5.004 36.24 7.512 ;
  LAYER M3 ;
        RECT 36.208 7.46 36.24 7.492 ;
  LAYER M1 ;
        RECT 36.144 5.004 36.176 7.512 ;
  LAYER M3 ;
        RECT 36.144 5.024 36.176 5.056 ;
  LAYER M1 ;
        RECT 36.08 5.004 36.112 7.512 ;
  LAYER M3 ;
        RECT 36.08 7.46 36.112 7.492 ;
  LAYER M1 ;
        RECT 36.016 5.004 36.048 7.512 ;
  LAYER M3 ;
        RECT 36.016 5.024 36.048 5.056 ;
  LAYER M1 ;
        RECT 35.952 5.004 35.984 7.512 ;
  LAYER M3 ;
        RECT 35.952 7.46 35.984 7.492 ;
  LAYER M1 ;
        RECT 35.888 5.004 35.92 7.512 ;
  LAYER M3 ;
        RECT 35.888 5.024 35.92 5.056 ;
  LAYER M1 ;
        RECT 35.824 5.004 35.856 7.512 ;
  LAYER M3 ;
        RECT 35.824 7.46 35.856 7.492 ;
  LAYER M1 ;
        RECT 35.76 5.004 35.792 7.512 ;
  LAYER M3 ;
        RECT 35.76 5.024 35.792 5.056 ;
  LAYER M1 ;
        RECT 35.696 5.004 35.728 7.512 ;
  LAYER M3 ;
        RECT 35.696 7.46 35.728 7.492 ;
  LAYER M1 ;
        RECT 35.632 5.004 35.664 7.512 ;
  LAYER M3 ;
        RECT 35.632 5.024 35.664 5.056 ;
  LAYER M1 ;
        RECT 35.568 5.004 35.6 7.512 ;
  LAYER M3 ;
        RECT 35.568 7.46 35.6 7.492 ;
  LAYER M1 ;
        RECT 35.504 5.004 35.536 7.512 ;
  LAYER M3 ;
        RECT 37.872 5.088 37.904 5.12 ;
  LAYER M2 ;
        RECT 35.504 5.152 35.536 5.184 ;
  LAYER M2 ;
        RECT 37.872 5.216 37.904 5.248 ;
  LAYER M2 ;
        RECT 35.504 5.28 35.536 5.312 ;
  LAYER M2 ;
        RECT 37.872 5.344 37.904 5.376 ;
  LAYER M2 ;
        RECT 35.504 5.408 35.536 5.44 ;
  LAYER M2 ;
        RECT 37.872 5.472 37.904 5.504 ;
  LAYER M2 ;
        RECT 35.504 5.536 35.536 5.568 ;
  LAYER M2 ;
        RECT 37.872 5.6 37.904 5.632 ;
  LAYER M2 ;
        RECT 35.504 5.664 35.536 5.696 ;
  LAYER M2 ;
        RECT 37.872 5.728 37.904 5.76 ;
  LAYER M2 ;
        RECT 35.504 5.792 35.536 5.824 ;
  LAYER M2 ;
        RECT 37.872 5.856 37.904 5.888 ;
  LAYER M2 ;
        RECT 35.504 5.92 35.536 5.952 ;
  LAYER M2 ;
        RECT 37.872 5.984 37.904 6.016 ;
  LAYER M2 ;
        RECT 35.504 6.048 35.536 6.08 ;
  LAYER M2 ;
        RECT 37.872 6.112 37.904 6.144 ;
  LAYER M2 ;
        RECT 35.504 6.176 35.536 6.208 ;
  LAYER M2 ;
        RECT 37.872 6.24 37.904 6.272 ;
  LAYER M2 ;
        RECT 35.504 6.304 35.536 6.336 ;
  LAYER M2 ;
        RECT 37.872 6.368 37.904 6.4 ;
  LAYER M2 ;
        RECT 35.504 6.432 35.536 6.464 ;
  LAYER M2 ;
        RECT 37.872 6.496 37.904 6.528 ;
  LAYER M2 ;
        RECT 35.504 6.56 35.536 6.592 ;
  LAYER M2 ;
        RECT 37.872 6.624 37.904 6.656 ;
  LAYER M2 ;
        RECT 35.504 6.688 35.536 6.72 ;
  LAYER M2 ;
        RECT 37.872 6.752 37.904 6.784 ;
  LAYER M2 ;
        RECT 35.504 6.816 35.536 6.848 ;
  LAYER M2 ;
        RECT 37.872 6.88 37.904 6.912 ;
  LAYER M2 ;
        RECT 35.504 6.944 35.536 6.976 ;
  LAYER M2 ;
        RECT 37.872 7.008 37.904 7.04 ;
  LAYER M2 ;
        RECT 35.504 7.072 35.536 7.104 ;
  LAYER M2 ;
        RECT 37.872 7.136 37.904 7.168 ;
  LAYER M2 ;
        RECT 35.504 7.2 35.536 7.232 ;
  LAYER M2 ;
        RECT 37.872 7.264 37.904 7.296 ;
  LAYER M2 ;
        RECT 35.504 7.328 35.536 7.36 ;
  LAYER M2 ;
        RECT 35.456 4.956 37.952 7.56 ;
  LAYER M1 ;
        RECT 37.872 8.112 37.904 10.62 ;
  LAYER M3 ;
        RECT 37.872 10.568 37.904 10.6 ;
  LAYER M1 ;
        RECT 37.808 8.112 37.84 10.62 ;
  LAYER M3 ;
        RECT 37.808 8.132 37.84 8.164 ;
  LAYER M1 ;
        RECT 37.744 8.112 37.776 10.62 ;
  LAYER M3 ;
        RECT 37.744 10.568 37.776 10.6 ;
  LAYER M1 ;
        RECT 37.68 8.112 37.712 10.62 ;
  LAYER M3 ;
        RECT 37.68 8.132 37.712 8.164 ;
  LAYER M1 ;
        RECT 37.616 8.112 37.648 10.62 ;
  LAYER M3 ;
        RECT 37.616 10.568 37.648 10.6 ;
  LAYER M1 ;
        RECT 37.552 8.112 37.584 10.62 ;
  LAYER M3 ;
        RECT 37.552 8.132 37.584 8.164 ;
  LAYER M1 ;
        RECT 37.488 8.112 37.52 10.62 ;
  LAYER M3 ;
        RECT 37.488 10.568 37.52 10.6 ;
  LAYER M1 ;
        RECT 37.424 8.112 37.456 10.62 ;
  LAYER M3 ;
        RECT 37.424 8.132 37.456 8.164 ;
  LAYER M1 ;
        RECT 37.36 8.112 37.392 10.62 ;
  LAYER M3 ;
        RECT 37.36 10.568 37.392 10.6 ;
  LAYER M1 ;
        RECT 37.296 8.112 37.328 10.62 ;
  LAYER M3 ;
        RECT 37.296 8.132 37.328 8.164 ;
  LAYER M1 ;
        RECT 37.232 8.112 37.264 10.62 ;
  LAYER M3 ;
        RECT 37.232 10.568 37.264 10.6 ;
  LAYER M1 ;
        RECT 37.168 8.112 37.2 10.62 ;
  LAYER M3 ;
        RECT 37.168 8.132 37.2 8.164 ;
  LAYER M1 ;
        RECT 37.104 8.112 37.136 10.62 ;
  LAYER M3 ;
        RECT 37.104 10.568 37.136 10.6 ;
  LAYER M1 ;
        RECT 37.04 8.112 37.072 10.62 ;
  LAYER M3 ;
        RECT 37.04 8.132 37.072 8.164 ;
  LAYER M1 ;
        RECT 36.976 8.112 37.008 10.62 ;
  LAYER M3 ;
        RECT 36.976 10.568 37.008 10.6 ;
  LAYER M1 ;
        RECT 36.912 8.112 36.944 10.62 ;
  LAYER M3 ;
        RECT 36.912 8.132 36.944 8.164 ;
  LAYER M1 ;
        RECT 36.848 8.112 36.88 10.62 ;
  LAYER M3 ;
        RECT 36.848 10.568 36.88 10.6 ;
  LAYER M1 ;
        RECT 36.784 8.112 36.816 10.62 ;
  LAYER M3 ;
        RECT 36.784 8.132 36.816 8.164 ;
  LAYER M1 ;
        RECT 36.72 8.112 36.752 10.62 ;
  LAYER M3 ;
        RECT 36.72 10.568 36.752 10.6 ;
  LAYER M1 ;
        RECT 36.656 8.112 36.688 10.62 ;
  LAYER M3 ;
        RECT 36.656 8.132 36.688 8.164 ;
  LAYER M1 ;
        RECT 36.592 8.112 36.624 10.62 ;
  LAYER M3 ;
        RECT 36.592 10.568 36.624 10.6 ;
  LAYER M1 ;
        RECT 36.528 8.112 36.56 10.62 ;
  LAYER M3 ;
        RECT 36.528 8.132 36.56 8.164 ;
  LAYER M1 ;
        RECT 36.464 8.112 36.496 10.62 ;
  LAYER M3 ;
        RECT 36.464 10.568 36.496 10.6 ;
  LAYER M1 ;
        RECT 36.4 8.112 36.432 10.62 ;
  LAYER M3 ;
        RECT 36.4 8.132 36.432 8.164 ;
  LAYER M1 ;
        RECT 36.336 8.112 36.368 10.62 ;
  LAYER M3 ;
        RECT 36.336 10.568 36.368 10.6 ;
  LAYER M1 ;
        RECT 36.272 8.112 36.304 10.62 ;
  LAYER M3 ;
        RECT 36.272 8.132 36.304 8.164 ;
  LAYER M1 ;
        RECT 36.208 8.112 36.24 10.62 ;
  LAYER M3 ;
        RECT 36.208 10.568 36.24 10.6 ;
  LAYER M1 ;
        RECT 36.144 8.112 36.176 10.62 ;
  LAYER M3 ;
        RECT 36.144 8.132 36.176 8.164 ;
  LAYER M1 ;
        RECT 36.08 8.112 36.112 10.62 ;
  LAYER M3 ;
        RECT 36.08 10.568 36.112 10.6 ;
  LAYER M1 ;
        RECT 36.016 8.112 36.048 10.62 ;
  LAYER M3 ;
        RECT 36.016 8.132 36.048 8.164 ;
  LAYER M1 ;
        RECT 35.952 8.112 35.984 10.62 ;
  LAYER M3 ;
        RECT 35.952 10.568 35.984 10.6 ;
  LAYER M1 ;
        RECT 35.888 8.112 35.92 10.62 ;
  LAYER M3 ;
        RECT 35.888 8.132 35.92 8.164 ;
  LAYER M1 ;
        RECT 35.824 8.112 35.856 10.62 ;
  LAYER M3 ;
        RECT 35.824 10.568 35.856 10.6 ;
  LAYER M1 ;
        RECT 35.76 8.112 35.792 10.62 ;
  LAYER M3 ;
        RECT 35.76 8.132 35.792 8.164 ;
  LAYER M1 ;
        RECT 35.696 8.112 35.728 10.62 ;
  LAYER M3 ;
        RECT 35.696 10.568 35.728 10.6 ;
  LAYER M1 ;
        RECT 35.632 8.112 35.664 10.62 ;
  LAYER M3 ;
        RECT 35.632 8.132 35.664 8.164 ;
  LAYER M1 ;
        RECT 35.568 8.112 35.6 10.62 ;
  LAYER M3 ;
        RECT 35.568 10.568 35.6 10.6 ;
  LAYER M1 ;
        RECT 35.504 8.112 35.536 10.62 ;
  LAYER M3 ;
        RECT 37.872 8.196 37.904 8.228 ;
  LAYER M2 ;
        RECT 35.504 8.26 35.536 8.292 ;
  LAYER M2 ;
        RECT 37.872 8.324 37.904 8.356 ;
  LAYER M2 ;
        RECT 35.504 8.388 35.536 8.42 ;
  LAYER M2 ;
        RECT 37.872 8.452 37.904 8.484 ;
  LAYER M2 ;
        RECT 35.504 8.516 35.536 8.548 ;
  LAYER M2 ;
        RECT 37.872 8.58 37.904 8.612 ;
  LAYER M2 ;
        RECT 35.504 8.644 35.536 8.676 ;
  LAYER M2 ;
        RECT 37.872 8.708 37.904 8.74 ;
  LAYER M2 ;
        RECT 35.504 8.772 35.536 8.804 ;
  LAYER M2 ;
        RECT 37.872 8.836 37.904 8.868 ;
  LAYER M2 ;
        RECT 35.504 8.9 35.536 8.932 ;
  LAYER M2 ;
        RECT 37.872 8.964 37.904 8.996 ;
  LAYER M2 ;
        RECT 35.504 9.028 35.536 9.06 ;
  LAYER M2 ;
        RECT 37.872 9.092 37.904 9.124 ;
  LAYER M2 ;
        RECT 35.504 9.156 35.536 9.188 ;
  LAYER M2 ;
        RECT 37.872 9.22 37.904 9.252 ;
  LAYER M2 ;
        RECT 35.504 9.284 35.536 9.316 ;
  LAYER M2 ;
        RECT 37.872 9.348 37.904 9.38 ;
  LAYER M2 ;
        RECT 35.504 9.412 35.536 9.444 ;
  LAYER M2 ;
        RECT 37.872 9.476 37.904 9.508 ;
  LAYER M2 ;
        RECT 35.504 9.54 35.536 9.572 ;
  LAYER M2 ;
        RECT 37.872 9.604 37.904 9.636 ;
  LAYER M2 ;
        RECT 35.504 9.668 35.536 9.7 ;
  LAYER M2 ;
        RECT 37.872 9.732 37.904 9.764 ;
  LAYER M2 ;
        RECT 35.504 9.796 35.536 9.828 ;
  LAYER M2 ;
        RECT 37.872 9.86 37.904 9.892 ;
  LAYER M2 ;
        RECT 35.504 9.924 35.536 9.956 ;
  LAYER M2 ;
        RECT 37.872 9.988 37.904 10.02 ;
  LAYER M2 ;
        RECT 35.504 10.052 35.536 10.084 ;
  LAYER M2 ;
        RECT 37.872 10.116 37.904 10.148 ;
  LAYER M2 ;
        RECT 35.504 10.18 35.536 10.212 ;
  LAYER M2 ;
        RECT 37.872 10.244 37.904 10.276 ;
  LAYER M2 ;
        RECT 35.504 10.308 35.536 10.34 ;
  LAYER M2 ;
        RECT 37.872 10.372 37.904 10.404 ;
  LAYER M2 ;
        RECT 35.504 10.436 35.536 10.468 ;
  LAYER M2 ;
        RECT 35.456 8.064 37.952 10.668 ;
  LAYER M1 ;
        RECT 37.872 11.22 37.904 13.728 ;
  LAYER M3 ;
        RECT 37.872 13.676 37.904 13.708 ;
  LAYER M1 ;
        RECT 37.808 11.22 37.84 13.728 ;
  LAYER M3 ;
        RECT 37.808 11.24 37.84 11.272 ;
  LAYER M1 ;
        RECT 37.744 11.22 37.776 13.728 ;
  LAYER M3 ;
        RECT 37.744 13.676 37.776 13.708 ;
  LAYER M1 ;
        RECT 37.68 11.22 37.712 13.728 ;
  LAYER M3 ;
        RECT 37.68 11.24 37.712 11.272 ;
  LAYER M1 ;
        RECT 37.616 11.22 37.648 13.728 ;
  LAYER M3 ;
        RECT 37.616 13.676 37.648 13.708 ;
  LAYER M1 ;
        RECT 37.552 11.22 37.584 13.728 ;
  LAYER M3 ;
        RECT 37.552 11.24 37.584 11.272 ;
  LAYER M1 ;
        RECT 37.488 11.22 37.52 13.728 ;
  LAYER M3 ;
        RECT 37.488 13.676 37.52 13.708 ;
  LAYER M1 ;
        RECT 37.424 11.22 37.456 13.728 ;
  LAYER M3 ;
        RECT 37.424 11.24 37.456 11.272 ;
  LAYER M1 ;
        RECT 37.36 11.22 37.392 13.728 ;
  LAYER M3 ;
        RECT 37.36 13.676 37.392 13.708 ;
  LAYER M1 ;
        RECT 37.296 11.22 37.328 13.728 ;
  LAYER M3 ;
        RECT 37.296 11.24 37.328 11.272 ;
  LAYER M1 ;
        RECT 37.232 11.22 37.264 13.728 ;
  LAYER M3 ;
        RECT 37.232 13.676 37.264 13.708 ;
  LAYER M1 ;
        RECT 37.168 11.22 37.2 13.728 ;
  LAYER M3 ;
        RECT 37.168 11.24 37.2 11.272 ;
  LAYER M1 ;
        RECT 37.104 11.22 37.136 13.728 ;
  LAYER M3 ;
        RECT 37.104 13.676 37.136 13.708 ;
  LAYER M1 ;
        RECT 37.04 11.22 37.072 13.728 ;
  LAYER M3 ;
        RECT 37.04 11.24 37.072 11.272 ;
  LAYER M1 ;
        RECT 36.976 11.22 37.008 13.728 ;
  LAYER M3 ;
        RECT 36.976 13.676 37.008 13.708 ;
  LAYER M1 ;
        RECT 36.912 11.22 36.944 13.728 ;
  LAYER M3 ;
        RECT 36.912 11.24 36.944 11.272 ;
  LAYER M1 ;
        RECT 36.848 11.22 36.88 13.728 ;
  LAYER M3 ;
        RECT 36.848 13.676 36.88 13.708 ;
  LAYER M1 ;
        RECT 36.784 11.22 36.816 13.728 ;
  LAYER M3 ;
        RECT 36.784 11.24 36.816 11.272 ;
  LAYER M1 ;
        RECT 36.72 11.22 36.752 13.728 ;
  LAYER M3 ;
        RECT 36.72 13.676 36.752 13.708 ;
  LAYER M1 ;
        RECT 36.656 11.22 36.688 13.728 ;
  LAYER M3 ;
        RECT 36.656 11.24 36.688 11.272 ;
  LAYER M1 ;
        RECT 36.592 11.22 36.624 13.728 ;
  LAYER M3 ;
        RECT 36.592 13.676 36.624 13.708 ;
  LAYER M1 ;
        RECT 36.528 11.22 36.56 13.728 ;
  LAYER M3 ;
        RECT 36.528 11.24 36.56 11.272 ;
  LAYER M1 ;
        RECT 36.464 11.22 36.496 13.728 ;
  LAYER M3 ;
        RECT 36.464 13.676 36.496 13.708 ;
  LAYER M1 ;
        RECT 36.4 11.22 36.432 13.728 ;
  LAYER M3 ;
        RECT 36.4 11.24 36.432 11.272 ;
  LAYER M1 ;
        RECT 36.336 11.22 36.368 13.728 ;
  LAYER M3 ;
        RECT 36.336 13.676 36.368 13.708 ;
  LAYER M1 ;
        RECT 36.272 11.22 36.304 13.728 ;
  LAYER M3 ;
        RECT 36.272 11.24 36.304 11.272 ;
  LAYER M1 ;
        RECT 36.208 11.22 36.24 13.728 ;
  LAYER M3 ;
        RECT 36.208 13.676 36.24 13.708 ;
  LAYER M1 ;
        RECT 36.144 11.22 36.176 13.728 ;
  LAYER M3 ;
        RECT 36.144 11.24 36.176 11.272 ;
  LAYER M1 ;
        RECT 36.08 11.22 36.112 13.728 ;
  LAYER M3 ;
        RECT 36.08 13.676 36.112 13.708 ;
  LAYER M1 ;
        RECT 36.016 11.22 36.048 13.728 ;
  LAYER M3 ;
        RECT 36.016 11.24 36.048 11.272 ;
  LAYER M1 ;
        RECT 35.952 11.22 35.984 13.728 ;
  LAYER M3 ;
        RECT 35.952 13.676 35.984 13.708 ;
  LAYER M1 ;
        RECT 35.888 11.22 35.92 13.728 ;
  LAYER M3 ;
        RECT 35.888 11.24 35.92 11.272 ;
  LAYER M1 ;
        RECT 35.824 11.22 35.856 13.728 ;
  LAYER M3 ;
        RECT 35.824 13.676 35.856 13.708 ;
  LAYER M1 ;
        RECT 35.76 11.22 35.792 13.728 ;
  LAYER M3 ;
        RECT 35.76 11.24 35.792 11.272 ;
  LAYER M1 ;
        RECT 35.696 11.22 35.728 13.728 ;
  LAYER M3 ;
        RECT 35.696 13.676 35.728 13.708 ;
  LAYER M1 ;
        RECT 35.632 11.22 35.664 13.728 ;
  LAYER M3 ;
        RECT 35.632 11.24 35.664 11.272 ;
  LAYER M1 ;
        RECT 35.568 11.22 35.6 13.728 ;
  LAYER M3 ;
        RECT 35.568 13.676 35.6 13.708 ;
  LAYER M1 ;
        RECT 35.504 11.22 35.536 13.728 ;
  LAYER M3 ;
        RECT 37.872 11.304 37.904 11.336 ;
  LAYER M2 ;
        RECT 35.504 11.368 35.536 11.4 ;
  LAYER M2 ;
        RECT 37.872 11.432 37.904 11.464 ;
  LAYER M2 ;
        RECT 35.504 11.496 35.536 11.528 ;
  LAYER M2 ;
        RECT 37.872 11.56 37.904 11.592 ;
  LAYER M2 ;
        RECT 35.504 11.624 35.536 11.656 ;
  LAYER M2 ;
        RECT 37.872 11.688 37.904 11.72 ;
  LAYER M2 ;
        RECT 35.504 11.752 35.536 11.784 ;
  LAYER M2 ;
        RECT 37.872 11.816 37.904 11.848 ;
  LAYER M2 ;
        RECT 35.504 11.88 35.536 11.912 ;
  LAYER M2 ;
        RECT 37.872 11.944 37.904 11.976 ;
  LAYER M2 ;
        RECT 35.504 12.008 35.536 12.04 ;
  LAYER M2 ;
        RECT 37.872 12.072 37.904 12.104 ;
  LAYER M2 ;
        RECT 35.504 12.136 35.536 12.168 ;
  LAYER M2 ;
        RECT 37.872 12.2 37.904 12.232 ;
  LAYER M2 ;
        RECT 35.504 12.264 35.536 12.296 ;
  LAYER M2 ;
        RECT 37.872 12.328 37.904 12.36 ;
  LAYER M2 ;
        RECT 35.504 12.392 35.536 12.424 ;
  LAYER M2 ;
        RECT 37.872 12.456 37.904 12.488 ;
  LAYER M2 ;
        RECT 35.504 12.52 35.536 12.552 ;
  LAYER M2 ;
        RECT 37.872 12.584 37.904 12.616 ;
  LAYER M2 ;
        RECT 35.504 12.648 35.536 12.68 ;
  LAYER M2 ;
        RECT 37.872 12.712 37.904 12.744 ;
  LAYER M2 ;
        RECT 35.504 12.776 35.536 12.808 ;
  LAYER M2 ;
        RECT 37.872 12.84 37.904 12.872 ;
  LAYER M2 ;
        RECT 35.504 12.904 35.536 12.936 ;
  LAYER M2 ;
        RECT 37.872 12.968 37.904 13 ;
  LAYER M2 ;
        RECT 35.504 13.032 35.536 13.064 ;
  LAYER M2 ;
        RECT 37.872 13.096 37.904 13.128 ;
  LAYER M2 ;
        RECT 35.504 13.16 35.536 13.192 ;
  LAYER M2 ;
        RECT 37.872 13.224 37.904 13.256 ;
  LAYER M2 ;
        RECT 35.504 13.288 35.536 13.32 ;
  LAYER M2 ;
        RECT 37.872 13.352 37.904 13.384 ;
  LAYER M2 ;
        RECT 35.504 13.416 35.536 13.448 ;
  LAYER M2 ;
        RECT 37.872 13.48 37.904 13.512 ;
  LAYER M2 ;
        RECT 35.504 13.544 35.536 13.576 ;
  LAYER M2 ;
        RECT 35.456 11.172 37.952 13.776 ;
  LAYER M1 ;
        RECT 34.896 1.896 34.928 4.404 ;
  LAYER M3 ;
        RECT 34.896 4.352 34.928 4.384 ;
  LAYER M1 ;
        RECT 34.832 1.896 34.864 4.404 ;
  LAYER M3 ;
        RECT 34.832 1.916 34.864 1.948 ;
  LAYER M1 ;
        RECT 34.768 1.896 34.8 4.404 ;
  LAYER M3 ;
        RECT 34.768 4.352 34.8 4.384 ;
  LAYER M1 ;
        RECT 34.704 1.896 34.736 4.404 ;
  LAYER M3 ;
        RECT 34.704 1.916 34.736 1.948 ;
  LAYER M1 ;
        RECT 34.64 1.896 34.672 4.404 ;
  LAYER M3 ;
        RECT 34.64 4.352 34.672 4.384 ;
  LAYER M1 ;
        RECT 34.576 1.896 34.608 4.404 ;
  LAYER M3 ;
        RECT 34.576 1.916 34.608 1.948 ;
  LAYER M1 ;
        RECT 34.512 1.896 34.544 4.404 ;
  LAYER M3 ;
        RECT 34.512 4.352 34.544 4.384 ;
  LAYER M1 ;
        RECT 34.448 1.896 34.48 4.404 ;
  LAYER M3 ;
        RECT 34.448 1.916 34.48 1.948 ;
  LAYER M1 ;
        RECT 34.384 1.896 34.416 4.404 ;
  LAYER M3 ;
        RECT 34.384 4.352 34.416 4.384 ;
  LAYER M1 ;
        RECT 34.32 1.896 34.352 4.404 ;
  LAYER M3 ;
        RECT 34.32 1.916 34.352 1.948 ;
  LAYER M1 ;
        RECT 34.256 1.896 34.288 4.404 ;
  LAYER M3 ;
        RECT 34.256 4.352 34.288 4.384 ;
  LAYER M1 ;
        RECT 34.192 1.896 34.224 4.404 ;
  LAYER M3 ;
        RECT 34.192 1.916 34.224 1.948 ;
  LAYER M1 ;
        RECT 34.128 1.896 34.16 4.404 ;
  LAYER M3 ;
        RECT 34.128 4.352 34.16 4.384 ;
  LAYER M1 ;
        RECT 34.064 1.896 34.096 4.404 ;
  LAYER M3 ;
        RECT 34.064 1.916 34.096 1.948 ;
  LAYER M1 ;
        RECT 34 1.896 34.032 4.404 ;
  LAYER M3 ;
        RECT 34 4.352 34.032 4.384 ;
  LAYER M1 ;
        RECT 33.936 1.896 33.968 4.404 ;
  LAYER M3 ;
        RECT 33.936 1.916 33.968 1.948 ;
  LAYER M1 ;
        RECT 33.872 1.896 33.904 4.404 ;
  LAYER M3 ;
        RECT 33.872 4.352 33.904 4.384 ;
  LAYER M1 ;
        RECT 33.808 1.896 33.84 4.404 ;
  LAYER M3 ;
        RECT 33.808 1.916 33.84 1.948 ;
  LAYER M1 ;
        RECT 33.744 1.896 33.776 4.404 ;
  LAYER M3 ;
        RECT 33.744 4.352 33.776 4.384 ;
  LAYER M1 ;
        RECT 33.68 1.896 33.712 4.404 ;
  LAYER M3 ;
        RECT 33.68 1.916 33.712 1.948 ;
  LAYER M1 ;
        RECT 33.616 1.896 33.648 4.404 ;
  LAYER M3 ;
        RECT 33.616 4.352 33.648 4.384 ;
  LAYER M1 ;
        RECT 33.552 1.896 33.584 4.404 ;
  LAYER M3 ;
        RECT 33.552 1.916 33.584 1.948 ;
  LAYER M1 ;
        RECT 33.488 1.896 33.52 4.404 ;
  LAYER M3 ;
        RECT 33.488 4.352 33.52 4.384 ;
  LAYER M1 ;
        RECT 33.424 1.896 33.456 4.404 ;
  LAYER M3 ;
        RECT 33.424 1.916 33.456 1.948 ;
  LAYER M1 ;
        RECT 33.36 1.896 33.392 4.404 ;
  LAYER M3 ;
        RECT 33.36 4.352 33.392 4.384 ;
  LAYER M1 ;
        RECT 33.296 1.896 33.328 4.404 ;
  LAYER M3 ;
        RECT 33.296 1.916 33.328 1.948 ;
  LAYER M1 ;
        RECT 33.232 1.896 33.264 4.404 ;
  LAYER M3 ;
        RECT 33.232 4.352 33.264 4.384 ;
  LAYER M1 ;
        RECT 33.168 1.896 33.2 4.404 ;
  LAYER M3 ;
        RECT 33.168 1.916 33.2 1.948 ;
  LAYER M1 ;
        RECT 33.104 1.896 33.136 4.404 ;
  LAYER M3 ;
        RECT 33.104 4.352 33.136 4.384 ;
  LAYER M1 ;
        RECT 33.04 1.896 33.072 4.404 ;
  LAYER M3 ;
        RECT 33.04 1.916 33.072 1.948 ;
  LAYER M1 ;
        RECT 32.976 1.896 33.008 4.404 ;
  LAYER M3 ;
        RECT 32.976 4.352 33.008 4.384 ;
  LAYER M1 ;
        RECT 32.912 1.896 32.944 4.404 ;
  LAYER M3 ;
        RECT 32.912 1.916 32.944 1.948 ;
  LAYER M1 ;
        RECT 32.848 1.896 32.88 4.404 ;
  LAYER M3 ;
        RECT 32.848 4.352 32.88 4.384 ;
  LAYER M1 ;
        RECT 32.784 1.896 32.816 4.404 ;
  LAYER M3 ;
        RECT 32.784 1.916 32.816 1.948 ;
  LAYER M1 ;
        RECT 32.72 1.896 32.752 4.404 ;
  LAYER M3 ;
        RECT 32.72 4.352 32.752 4.384 ;
  LAYER M1 ;
        RECT 32.656 1.896 32.688 4.404 ;
  LAYER M3 ;
        RECT 32.656 1.916 32.688 1.948 ;
  LAYER M1 ;
        RECT 32.592 1.896 32.624 4.404 ;
  LAYER M3 ;
        RECT 32.592 4.352 32.624 4.384 ;
  LAYER M1 ;
        RECT 32.528 1.896 32.56 4.404 ;
  LAYER M3 ;
        RECT 34.896 1.98 34.928 2.012 ;
  LAYER M2 ;
        RECT 32.528 2.044 32.56 2.076 ;
  LAYER M2 ;
        RECT 34.896 2.108 34.928 2.14 ;
  LAYER M2 ;
        RECT 32.528 2.172 32.56 2.204 ;
  LAYER M2 ;
        RECT 34.896 2.236 34.928 2.268 ;
  LAYER M2 ;
        RECT 32.528 2.3 32.56 2.332 ;
  LAYER M2 ;
        RECT 34.896 2.364 34.928 2.396 ;
  LAYER M2 ;
        RECT 32.528 2.428 32.56 2.46 ;
  LAYER M2 ;
        RECT 34.896 2.492 34.928 2.524 ;
  LAYER M2 ;
        RECT 32.528 2.556 32.56 2.588 ;
  LAYER M2 ;
        RECT 34.896 2.62 34.928 2.652 ;
  LAYER M2 ;
        RECT 32.528 2.684 32.56 2.716 ;
  LAYER M2 ;
        RECT 34.896 2.748 34.928 2.78 ;
  LAYER M2 ;
        RECT 32.528 2.812 32.56 2.844 ;
  LAYER M2 ;
        RECT 34.896 2.876 34.928 2.908 ;
  LAYER M2 ;
        RECT 32.528 2.94 32.56 2.972 ;
  LAYER M2 ;
        RECT 34.896 3.004 34.928 3.036 ;
  LAYER M2 ;
        RECT 32.528 3.068 32.56 3.1 ;
  LAYER M2 ;
        RECT 34.896 3.132 34.928 3.164 ;
  LAYER M2 ;
        RECT 32.528 3.196 32.56 3.228 ;
  LAYER M2 ;
        RECT 34.896 3.26 34.928 3.292 ;
  LAYER M2 ;
        RECT 32.528 3.324 32.56 3.356 ;
  LAYER M2 ;
        RECT 34.896 3.388 34.928 3.42 ;
  LAYER M2 ;
        RECT 32.528 3.452 32.56 3.484 ;
  LAYER M2 ;
        RECT 34.896 3.516 34.928 3.548 ;
  LAYER M2 ;
        RECT 32.528 3.58 32.56 3.612 ;
  LAYER M2 ;
        RECT 34.896 3.644 34.928 3.676 ;
  LAYER M2 ;
        RECT 32.528 3.708 32.56 3.74 ;
  LAYER M2 ;
        RECT 34.896 3.772 34.928 3.804 ;
  LAYER M2 ;
        RECT 32.528 3.836 32.56 3.868 ;
  LAYER M2 ;
        RECT 34.896 3.9 34.928 3.932 ;
  LAYER M2 ;
        RECT 32.528 3.964 32.56 3.996 ;
  LAYER M2 ;
        RECT 34.896 4.028 34.928 4.06 ;
  LAYER M2 ;
        RECT 32.528 4.092 32.56 4.124 ;
  LAYER M2 ;
        RECT 34.896 4.156 34.928 4.188 ;
  LAYER M2 ;
        RECT 32.528 4.22 32.56 4.252 ;
  LAYER M2 ;
        RECT 32.48 1.848 34.976 4.452 ;
  LAYER M1 ;
        RECT 34.896 5.004 34.928 7.512 ;
  LAYER M3 ;
        RECT 34.896 7.46 34.928 7.492 ;
  LAYER M1 ;
        RECT 34.832 5.004 34.864 7.512 ;
  LAYER M3 ;
        RECT 34.832 5.024 34.864 5.056 ;
  LAYER M1 ;
        RECT 34.768 5.004 34.8 7.512 ;
  LAYER M3 ;
        RECT 34.768 7.46 34.8 7.492 ;
  LAYER M1 ;
        RECT 34.704 5.004 34.736 7.512 ;
  LAYER M3 ;
        RECT 34.704 5.024 34.736 5.056 ;
  LAYER M1 ;
        RECT 34.64 5.004 34.672 7.512 ;
  LAYER M3 ;
        RECT 34.64 7.46 34.672 7.492 ;
  LAYER M1 ;
        RECT 34.576 5.004 34.608 7.512 ;
  LAYER M3 ;
        RECT 34.576 5.024 34.608 5.056 ;
  LAYER M1 ;
        RECT 34.512 5.004 34.544 7.512 ;
  LAYER M3 ;
        RECT 34.512 7.46 34.544 7.492 ;
  LAYER M1 ;
        RECT 34.448 5.004 34.48 7.512 ;
  LAYER M3 ;
        RECT 34.448 5.024 34.48 5.056 ;
  LAYER M1 ;
        RECT 34.384 5.004 34.416 7.512 ;
  LAYER M3 ;
        RECT 34.384 7.46 34.416 7.492 ;
  LAYER M1 ;
        RECT 34.32 5.004 34.352 7.512 ;
  LAYER M3 ;
        RECT 34.32 5.024 34.352 5.056 ;
  LAYER M1 ;
        RECT 34.256 5.004 34.288 7.512 ;
  LAYER M3 ;
        RECT 34.256 7.46 34.288 7.492 ;
  LAYER M1 ;
        RECT 34.192 5.004 34.224 7.512 ;
  LAYER M3 ;
        RECT 34.192 5.024 34.224 5.056 ;
  LAYER M1 ;
        RECT 34.128 5.004 34.16 7.512 ;
  LAYER M3 ;
        RECT 34.128 7.46 34.16 7.492 ;
  LAYER M1 ;
        RECT 34.064 5.004 34.096 7.512 ;
  LAYER M3 ;
        RECT 34.064 5.024 34.096 5.056 ;
  LAYER M1 ;
        RECT 34 5.004 34.032 7.512 ;
  LAYER M3 ;
        RECT 34 7.46 34.032 7.492 ;
  LAYER M1 ;
        RECT 33.936 5.004 33.968 7.512 ;
  LAYER M3 ;
        RECT 33.936 5.024 33.968 5.056 ;
  LAYER M1 ;
        RECT 33.872 5.004 33.904 7.512 ;
  LAYER M3 ;
        RECT 33.872 7.46 33.904 7.492 ;
  LAYER M1 ;
        RECT 33.808 5.004 33.84 7.512 ;
  LAYER M3 ;
        RECT 33.808 5.024 33.84 5.056 ;
  LAYER M1 ;
        RECT 33.744 5.004 33.776 7.512 ;
  LAYER M3 ;
        RECT 33.744 7.46 33.776 7.492 ;
  LAYER M1 ;
        RECT 33.68 5.004 33.712 7.512 ;
  LAYER M3 ;
        RECT 33.68 5.024 33.712 5.056 ;
  LAYER M1 ;
        RECT 33.616 5.004 33.648 7.512 ;
  LAYER M3 ;
        RECT 33.616 7.46 33.648 7.492 ;
  LAYER M1 ;
        RECT 33.552 5.004 33.584 7.512 ;
  LAYER M3 ;
        RECT 33.552 5.024 33.584 5.056 ;
  LAYER M1 ;
        RECT 33.488 5.004 33.52 7.512 ;
  LAYER M3 ;
        RECT 33.488 7.46 33.52 7.492 ;
  LAYER M1 ;
        RECT 33.424 5.004 33.456 7.512 ;
  LAYER M3 ;
        RECT 33.424 5.024 33.456 5.056 ;
  LAYER M1 ;
        RECT 33.36 5.004 33.392 7.512 ;
  LAYER M3 ;
        RECT 33.36 7.46 33.392 7.492 ;
  LAYER M1 ;
        RECT 33.296 5.004 33.328 7.512 ;
  LAYER M3 ;
        RECT 33.296 5.024 33.328 5.056 ;
  LAYER M1 ;
        RECT 33.232 5.004 33.264 7.512 ;
  LAYER M3 ;
        RECT 33.232 7.46 33.264 7.492 ;
  LAYER M1 ;
        RECT 33.168 5.004 33.2 7.512 ;
  LAYER M3 ;
        RECT 33.168 5.024 33.2 5.056 ;
  LAYER M1 ;
        RECT 33.104 5.004 33.136 7.512 ;
  LAYER M3 ;
        RECT 33.104 7.46 33.136 7.492 ;
  LAYER M1 ;
        RECT 33.04 5.004 33.072 7.512 ;
  LAYER M3 ;
        RECT 33.04 5.024 33.072 5.056 ;
  LAYER M1 ;
        RECT 32.976 5.004 33.008 7.512 ;
  LAYER M3 ;
        RECT 32.976 7.46 33.008 7.492 ;
  LAYER M1 ;
        RECT 32.912 5.004 32.944 7.512 ;
  LAYER M3 ;
        RECT 32.912 5.024 32.944 5.056 ;
  LAYER M1 ;
        RECT 32.848 5.004 32.88 7.512 ;
  LAYER M3 ;
        RECT 32.848 7.46 32.88 7.492 ;
  LAYER M1 ;
        RECT 32.784 5.004 32.816 7.512 ;
  LAYER M3 ;
        RECT 32.784 5.024 32.816 5.056 ;
  LAYER M1 ;
        RECT 32.72 5.004 32.752 7.512 ;
  LAYER M3 ;
        RECT 32.72 7.46 32.752 7.492 ;
  LAYER M1 ;
        RECT 32.656 5.004 32.688 7.512 ;
  LAYER M3 ;
        RECT 32.656 5.024 32.688 5.056 ;
  LAYER M1 ;
        RECT 32.592 5.004 32.624 7.512 ;
  LAYER M3 ;
        RECT 32.592 7.46 32.624 7.492 ;
  LAYER M1 ;
        RECT 32.528 5.004 32.56 7.512 ;
  LAYER M3 ;
        RECT 34.896 5.088 34.928 5.12 ;
  LAYER M2 ;
        RECT 32.528 5.152 32.56 5.184 ;
  LAYER M2 ;
        RECT 34.896 5.216 34.928 5.248 ;
  LAYER M2 ;
        RECT 32.528 5.28 32.56 5.312 ;
  LAYER M2 ;
        RECT 34.896 5.344 34.928 5.376 ;
  LAYER M2 ;
        RECT 32.528 5.408 32.56 5.44 ;
  LAYER M2 ;
        RECT 34.896 5.472 34.928 5.504 ;
  LAYER M2 ;
        RECT 32.528 5.536 32.56 5.568 ;
  LAYER M2 ;
        RECT 34.896 5.6 34.928 5.632 ;
  LAYER M2 ;
        RECT 32.528 5.664 32.56 5.696 ;
  LAYER M2 ;
        RECT 34.896 5.728 34.928 5.76 ;
  LAYER M2 ;
        RECT 32.528 5.792 32.56 5.824 ;
  LAYER M2 ;
        RECT 34.896 5.856 34.928 5.888 ;
  LAYER M2 ;
        RECT 32.528 5.92 32.56 5.952 ;
  LAYER M2 ;
        RECT 34.896 5.984 34.928 6.016 ;
  LAYER M2 ;
        RECT 32.528 6.048 32.56 6.08 ;
  LAYER M2 ;
        RECT 34.896 6.112 34.928 6.144 ;
  LAYER M2 ;
        RECT 32.528 6.176 32.56 6.208 ;
  LAYER M2 ;
        RECT 34.896 6.24 34.928 6.272 ;
  LAYER M2 ;
        RECT 32.528 6.304 32.56 6.336 ;
  LAYER M2 ;
        RECT 34.896 6.368 34.928 6.4 ;
  LAYER M2 ;
        RECT 32.528 6.432 32.56 6.464 ;
  LAYER M2 ;
        RECT 34.896 6.496 34.928 6.528 ;
  LAYER M2 ;
        RECT 32.528 6.56 32.56 6.592 ;
  LAYER M2 ;
        RECT 34.896 6.624 34.928 6.656 ;
  LAYER M2 ;
        RECT 32.528 6.688 32.56 6.72 ;
  LAYER M2 ;
        RECT 34.896 6.752 34.928 6.784 ;
  LAYER M2 ;
        RECT 32.528 6.816 32.56 6.848 ;
  LAYER M2 ;
        RECT 34.896 6.88 34.928 6.912 ;
  LAYER M2 ;
        RECT 32.528 6.944 32.56 6.976 ;
  LAYER M2 ;
        RECT 34.896 7.008 34.928 7.04 ;
  LAYER M2 ;
        RECT 32.528 7.072 32.56 7.104 ;
  LAYER M2 ;
        RECT 34.896 7.136 34.928 7.168 ;
  LAYER M2 ;
        RECT 32.528 7.2 32.56 7.232 ;
  LAYER M2 ;
        RECT 34.896 7.264 34.928 7.296 ;
  LAYER M2 ;
        RECT 32.528 7.328 32.56 7.36 ;
  LAYER M2 ;
        RECT 32.48 4.956 34.976 7.56 ;
  LAYER M1 ;
        RECT 34.896 8.112 34.928 10.62 ;
  LAYER M3 ;
        RECT 34.896 10.568 34.928 10.6 ;
  LAYER M1 ;
        RECT 34.832 8.112 34.864 10.62 ;
  LAYER M3 ;
        RECT 34.832 8.132 34.864 8.164 ;
  LAYER M1 ;
        RECT 34.768 8.112 34.8 10.62 ;
  LAYER M3 ;
        RECT 34.768 10.568 34.8 10.6 ;
  LAYER M1 ;
        RECT 34.704 8.112 34.736 10.62 ;
  LAYER M3 ;
        RECT 34.704 8.132 34.736 8.164 ;
  LAYER M1 ;
        RECT 34.64 8.112 34.672 10.62 ;
  LAYER M3 ;
        RECT 34.64 10.568 34.672 10.6 ;
  LAYER M1 ;
        RECT 34.576 8.112 34.608 10.62 ;
  LAYER M3 ;
        RECT 34.576 8.132 34.608 8.164 ;
  LAYER M1 ;
        RECT 34.512 8.112 34.544 10.62 ;
  LAYER M3 ;
        RECT 34.512 10.568 34.544 10.6 ;
  LAYER M1 ;
        RECT 34.448 8.112 34.48 10.62 ;
  LAYER M3 ;
        RECT 34.448 8.132 34.48 8.164 ;
  LAYER M1 ;
        RECT 34.384 8.112 34.416 10.62 ;
  LAYER M3 ;
        RECT 34.384 10.568 34.416 10.6 ;
  LAYER M1 ;
        RECT 34.32 8.112 34.352 10.62 ;
  LAYER M3 ;
        RECT 34.32 8.132 34.352 8.164 ;
  LAYER M1 ;
        RECT 34.256 8.112 34.288 10.62 ;
  LAYER M3 ;
        RECT 34.256 10.568 34.288 10.6 ;
  LAYER M1 ;
        RECT 34.192 8.112 34.224 10.62 ;
  LAYER M3 ;
        RECT 34.192 8.132 34.224 8.164 ;
  LAYER M1 ;
        RECT 34.128 8.112 34.16 10.62 ;
  LAYER M3 ;
        RECT 34.128 10.568 34.16 10.6 ;
  LAYER M1 ;
        RECT 34.064 8.112 34.096 10.62 ;
  LAYER M3 ;
        RECT 34.064 8.132 34.096 8.164 ;
  LAYER M1 ;
        RECT 34 8.112 34.032 10.62 ;
  LAYER M3 ;
        RECT 34 10.568 34.032 10.6 ;
  LAYER M1 ;
        RECT 33.936 8.112 33.968 10.62 ;
  LAYER M3 ;
        RECT 33.936 8.132 33.968 8.164 ;
  LAYER M1 ;
        RECT 33.872 8.112 33.904 10.62 ;
  LAYER M3 ;
        RECT 33.872 10.568 33.904 10.6 ;
  LAYER M1 ;
        RECT 33.808 8.112 33.84 10.62 ;
  LAYER M3 ;
        RECT 33.808 8.132 33.84 8.164 ;
  LAYER M1 ;
        RECT 33.744 8.112 33.776 10.62 ;
  LAYER M3 ;
        RECT 33.744 10.568 33.776 10.6 ;
  LAYER M1 ;
        RECT 33.68 8.112 33.712 10.62 ;
  LAYER M3 ;
        RECT 33.68 8.132 33.712 8.164 ;
  LAYER M1 ;
        RECT 33.616 8.112 33.648 10.62 ;
  LAYER M3 ;
        RECT 33.616 10.568 33.648 10.6 ;
  LAYER M1 ;
        RECT 33.552 8.112 33.584 10.62 ;
  LAYER M3 ;
        RECT 33.552 8.132 33.584 8.164 ;
  LAYER M1 ;
        RECT 33.488 8.112 33.52 10.62 ;
  LAYER M3 ;
        RECT 33.488 10.568 33.52 10.6 ;
  LAYER M1 ;
        RECT 33.424 8.112 33.456 10.62 ;
  LAYER M3 ;
        RECT 33.424 8.132 33.456 8.164 ;
  LAYER M1 ;
        RECT 33.36 8.112 33.392 10.62 ;
  LAYER M3 ;
        RECT 33.36 10.568 33.392 10.6 ;
  LAYER M1 ;
        RECT 33.296 8.112 33.328 10.62 ;
  LAYER M3 ;
        RECT 33.296 8.132 33.328 8.164 ;
  LAYER M1 ;
        RECT 33.232 8.112 33.264 10.62 ;
  LAYER M3 ;
        RECT 33.232 10.568 33.264 10.6 ;
  LAYER M1 ;
        RECT 33.168 8.112 33.2 10.62 ;
  LAYER M3 ;
        RECT 33.168 8.132 33.2 8.164 ;
  LAYER M1 ;
        RECT 33.104 8.112 33.136 10.62 ;
  LAYER M3 ;
        RECT 33.104 10.568 33.136 10.6 ;
  LAYER M1 ;
        RECT 33.04 8.112 33.072 10.62 ;
  LAYER M3 ;
        RECT 33.04 8.132 33.072 8.164 ;
  LAYER M1 ;
        RECT 32.976 8.112 33.008 10.62 ;
  LAYER M3 ;
        RECT 32.976 10.568 33.008 10.6 ;
  LAYER M1 ;
        RECT 32.912 8.112 32.944 10.62 ;
  LAYER M3 ;
        RECT 32.912 8.132 32.944 8.164 ;
  LAYER M1 ;
        RECT 32.848 8.112 32.88 10.62 ;
  LAYER M3 ;
        RECT 32.848 10.568 32.88 10.6 ;
  LAYER M1 ;
        RECT 32.784 8.112 32.816 10.62 ;
  LAYER M3 ;
        RECT 32.784 8.132 32.816 8.164 ;
  LAYER M1 ;
        RECT 32.72 8.112 32.752 10.62 ;
  LAYER M3 ;
        RECT 32.72 10.568 32.752 10.6 ;
  LAYER M1 ;
        RECT 32.656 8.112 32.688 10.62 ;
  LAYER M3 ;
        RECT 32.656 8.132 32.688 8.164 ;
  LAYER M1 ;
        RECT 32.592 8.112 32.624 10.62 ;
  LAYER M3 ;
        RECT 32.592 10.568 32.624 10.6 ;
  LAYER M1 ;
        RECT 32.528 8.112 32.56 10.62 ;
  LAYER M3 ;
        RECT 34.896 8.196 34.928 8.228 ;
  LAYER M2 ;
        RECT 32.528 8.26 32.56 8.292 ;
  LAYER M2 ;
        RECT 34.896 8.324 34.928 8.356 ;
  LAYER M2 ;
        RECT 32.528 8.388 32.56 8.42 ;
  LAYER M2 ;
        RECT 34.896 8.452 34.928 8.484 ;
  LAYER M2 ;
        RECT 32.528 8.516 32.56 8.548 ;
  LAYER M2 ;
        RECT 34.896 8.58 34.928 8.612 ;
  LAYER M2 ;
        RECT 32.528 8.644 32.56 8.676 ;
  LAYER M2 ;
        RECT 34.896 8.708 34.928 8.74 ;
  LAYER M2 ;
        RECT 32.528 8.772 32.56 8.804 ;
  LAYER M2 ;
        RECT 34.896 8.836 34.928 8.868 ;
  LAYER M2 ;
        RECT 32.528 8.9 32.56 8.932 ;
  LAYER M2 ;
        RECT 34.896 8.964 34.928 8.996 ;
  LAYER M2 ;
        RECT 32.528 9.028 32.56 9.06 ;
  LAYER M2 ;
        RECT 34.896 9.092 34.928 9.124 ;
  LAYER M2 ;
        RECT 32.528 9.156 32.56 9.188 ;
  LAYER M2 ;
        RECT 34.896 9.22 34.928 9.252 ;
  LAYER M2 ;
        RECT 32.528 9.284 32.56 9.316 ;
  LAYER M2 ;
        RECT 34.896 9.348 34.928 9.38 ;
  LAYER M2 ;
        RECT 32.528 9.412 32.56 9.444 ;
  LAYER M2 ;
        RECT 34.896 9.476 34.928 9.508 ;
  LAYER M2 ;
        RECT 32.528 9.54 32.56 9.572 ;
  LAYER M2 ;
        RECT 34.896 9.604 34.928 9.636 ;
  LAYER M2 ;
        RECT 32.528 9.668 32.56 9.7 ;
  LAYER M2 ;
        RECT 34.896 9.732 34.928 9.764 ;
  LAYER M2 ;
        RECT 32.528 9.796 32.56 9.828 ;
  LAYER M2 ;
        RECT 34.896 9.86 34.928 9.892 ;
  LAYER M2 ;
        RECT 32.528 9.924 32.56 9.956 ;
  LAYER M2 ;
        RECT 34.896 9.988 34.928 10.02 ;
  LAYER M2 ;
        RECT 32.528 10.052 32.56 10.084 ;
  LAYER M2 ;
        RECT 34.896 10.116 34.928 10.148 ;
  LAYER M2 ;
        RECT 32.528 10.18 32.56 10.212 ;
  LAYER M2 ;
        RECT 34.896 10.244 34.928 10.276 ;
  LAYER M2 ;
        RECT 32.528 10.308 32.56 10.34 ;
  LAYER M2 ;
        RECT 34.896 10.372 34.928 10.404 ;
  LAYER M2 ;
        RECT 32.528 10.436 32.56 10.468 ;
  LAYER M2 ;
        RECT 32.48 8.064 34.976 10.668 ;
  LAYER M1 ;
        RECT 34.896 11.22 34.928 13.728 ;
  LAYER M3 ;
        RECT 34.896 13.676 34.928 13.708 ;
  LAYER M1 ;
        RECT 34.832 11.22 34.864 13.728 ;
  LAYER M3 ;
        RECT 34.832 11.24 34.864 11.272 ;
  LAYER M1 ;
        RECT 34.768 11.22 34.8 13.728 ;
  LAYER M3 ;
        RECT 34.768 13.676 34.8 13.708 ;
  LAYER M1 ;
        RECT 34.704 11.22 34.736 13.728 ;
  LAYER M3 ;
        RECT 34.704 11.24 34.736 11.272 ;
  LAYER M1 ;
        RECT 34.64 11.22 34.672 13.728 ;
  LAYER M3 ;
        RECT 34.64 13.676 34.672 13.708 ;
  LAYER M1 ;
        RECT 34.576 11.22 34.608 13.728 ;
  LAYER M3 ;
        RECT 34.576 11.24 34.608 11.272 ;
  LAYER M1 ;
        RECT 34.512 11.22 34.544 13.728 ;
  LAYER M3 ;
        RECT 34.512 13.676 34.544 13.708 ;
  LAYER M1 ;
        RECT 34.448 11.22 34.48 13.728 ;
  LAYER M3 ;
        RECT 34.448 11.24 34.48 11.272 ;
  LAYER M1 ;
        RECT 34.384 11.22 34.416 13.728 ;
  LAYER M3 ;
        RECT 34.384 13.676 34.416 13.708 ;
  LAYER M1 ;
        RECT 34.32 11.22 34.352 13.728 ;
  LAYER M3 ;
        RECT 34.32 11.24 34.352 11.272 ;
  LAYER M1 ;
        RECT 34.256 11.22 34.288 13.728 ;
  LAYER M3 ;
        RECT 34.256 13.676 34.288 13.708 ;
  LAYER M1 ;
        RECT 34.192 11.22 34.224 13.728 ;
  LAYER M3 ;
        RECT 34.192 11.24 34.224 11.272 ;
  LAYER M1 ;
        RECT 34.128 11.22 34.16 13.728 ;
  LAYER M3 ;
        RECT 34.128 13.676 34.16 13.708 ;
  LAYER M1 ;
        RECT 34.064 11.22 34.096 13.728 ;
  LAYER M3 ;
        RECT 34.064 11.24 34.096 11.272 ;
  LAYER M1 ;
        RECT 34 11.22 34.032 13.728 ;
  LAYER M3 ;
        RECT 34 13.676 34.032 13.708 ;
  LAYER M1 ;
        RECT 33.936 11.22 33.968 13.728 ;
  LAYER M3 ;
        RECT 33.936 11.24 33.968 11.272 ;
  LAYER M1 ;
        RECT 33.872 11.22 33.904 13.728 ;
  LAYER M3 ;
        RECT 33.872 13.676 33.904 13.708 ;
  LAYER M1 ;
        RECT 33.808 11.22 33.84 13.728 ;
  LAYER M3 ;
        RECT 33.808 11.24 33.84 11.272 ;
  LAYER M1 ;
        RECT 33.744 11.22 33.776 13.728 ;
  LAYER M3 ;
        RECT 33.744 13.676 33.776 13.708 ;
  LAYER M1 ;
        RECT 33.68 11.22 33.712 13.728 ;
  LAYER M3 ;
        RECT 33.68 11.24 33.712 11.272 ;
  LAYER M1 ;
        RECT 33.616 11.22 33.648 13.728 ;
  LAYER M3 ;
        RECT 33.616 13.676 33.648 13.708 ;
  LAYER M1 ;
        RECT 33.552 11.22 33.584 13.728 ;
  LAYER M3 ;
        RECT 33.552 11.24 33.584 11.272 ;
  LAYER M1 ;
        RECT 33.488 11.22 33.52 13.728 ;
  LAYER M3 ;
        RECT 33.488 13.676 33.52 13.708 ;
  LAYER M1 ;
        RECT 33.424 11.22 33.456 13.728 ;
  LAYER M3 ;
        RECT 33.424 11.24 33.456 11.272 ;
  LAYER M1 ;
        RECT 33.36 11.22 33.392 13.728 ;
  LAYER M3 ;
        RECT 33.36 13.676 33.392 13.708 ;
  LAYER M1 ;
        RECT 33.296 11.22 33.328 13.728 ;
  LAYER M3 ;
        RECT 33.296 11.24 33.328 11.272 ;
  LAYER M1 ;
        RECT 33.232 11.22 33.264 13.728 ;
  LAYER M3 ;
        RECT 33.232 13.676 33.264 13.708 ;
  LAYER M1 ;
        RECT 33.168 11.22 33.2 13.728 ;
  LAYER M3 ;
        RECT 33.168 11.24 33.2 11.272 ;
  LAYER M1 ;
        RECT 33.104 11.22 33.136 13.728 ;
  LAYER M3 ;
        RECT 33.104 13.676 33.136 13.708 ;
  LAYER M1 ;
        RECT 33.04 11.22 33.072 13.728 ;
  LAYER M3 ;
        RECT 33.04 11.24 33.072 11.272 ;
  LAYER M1 ;
        RECT 32.976 11.22 33.008 13.728 ;
  LAYER M3 ;
        RECT 32.976 13.676 33.008 13.708 ;
  LAYER M1 ;
        RECT 32.912 11.22 32.944 13.728 ;
  LAYER M3 ;
        RECT 32.912 11.24 32.944 11.272 ;
  LAYER M1 ;
        RECT 32.848 11.22 32.88 13.728 ;
  LAYER M3 ;
        RECT 32.848 13.676 32.88 13.708 ;
  LAYER M1 ;
        RECT 32.784 11.22 32.816 13.728 ;
  LAYER M3 ;
        RECT 32.784 11.24 32.816 11.272 ;
  LAYER M1 ;
        RECT 32.72 11.22 32.752 13.728 ;
  LAYER M3 ;
        RECT 32.72 13.676 32.752 13.708 ;
  LAYER M1 ;
        RECT 32.656 11.22 32.688 13.728 ;
  LAYER M3 ;
        RECT 32.656 11.24 32.688 11.272 ;
  LAYER M1 ;
        RECT 32.592 11.22 32.624 13.728 ;
  LAYER M3 ;
        RECT 32.592 13.676 32.624 13.708 ;
  LAYER M1 ;
        RECT 32.528 11.22 32.56 13.728 ;
  LAYER M3 ;
        RECT 34.896 11.304 34.928 11.336 ;
  LAYER M2 ;
        RECT 32.528 11.368 32.56 11.4 ;
  LAYER M2 ;
        RECT 34.896 11.432 34.928 11.464 ;
  LAYER M2 ;
        RECT 32.528 11.496 32.56 11.528 ;
  LAYER M2 ;
        RECT 34.896 11.56 34.928 11.592 ;
  LAYER M2 ;
        RECT 32.528 11.624 32.56 11.656 ;
  LAYER M2 ;
        RECT 34.896 11.688 34.928 11.72 ;
  LAYER M2 ;
        RECT 32.528 11.752 32.56 11.784 ;
  LAYER M2 ;
        RECT 34.896 11.816 34.928 11.848 ;
  LAYER M2 ;
        RECT 32.528 11.88 32.56 11.912 ;
  LAYER M2 ;
        RECT 34.896 11.944 34.928 11.976 ;
  LAYER M2 ;
        RECT 32.528 12.008 32.56 12.04 ;
  LAYER M2 ;
        RECT 34.896 12.072 34.928 12.104 ;
  LAYER M2 ;
        RECT 32.528 12.136 32.56 12.168 ;
  LAYER M2 ;
        RECT 34.896 12.2 34.928 12.232 ;
  LAYER M2 ;
        RECT 32.528 12.264 32.56 12.296 ;
  LAYER M2 ;
        RECT 34.896 12.328 34.928 12.36 ;
  LAYER M2 ;
        RECT 32.528 12.392 32.56 12.424 ;
  LAYER M2 ;
        RECT 34.896 12.456 34.928 12.488 ;
  LAYER M2 ;
        RECT 32.528 12.52 32.56 12.552 ;
  LAYER M2 ;
        RECT 34.896 12.584 34.928 12.616 ;
  LAYER M2 ;
        RECT 32.528 12.648 32.56 12.68 ;
  LAYER M2 ;
        RECT 34.896 12.712 34.928 12.744 ;
  LAYER M2 ;
        RECT 32.528 12.776 32.56 12.808 ;
  LAYER M2 ;
        RECT 34.896 12.84 34.928 12.872 ;
  LAYER M2 ;
        RECT 32.528 12.904 32.56 12.936 ;
  LAYER M2 ;
        RECT 34.896 12.968 34.928 13 ;
  LAYER M2 ;
        RECT 32.528 13.032 32.56 13.064 ;
  LAYER M2 ;
        RECT 34.896 13.096 34.928 13.128 ;
  LAYER M2 ;
        RECT 32.528 13.16 32.56 13.192 ;
  LAYER M2 ;
        RECT 34.896 13.224 34.928 13.256 ;
  LAYER M2 ;
        RECT 32.528 13.288 32.56 13.32 ;
  LAYER M2 ;
        RECT 34.896 13.352 34.928 13.384 ;
  LAYER M2 ;
        RECT 32.528 13.416 32.56 13.448 ;
  LAYER M2 ;
        RECT 34.896 13.48 34.928 13.512 ;
  LAYER M2 ;
        RECT 32.528 13.544 32.56 13.576 ;
  LAYER M2 ;
        RECT 32.48 11.172 34.976 13.776 ;
  LAYER M1 ;
        RECT 42.144 0.216 42.176 0.876 ;
  LAYER M1 ;
        RECT 42.224 0.216 42.256 0.876 ;
  LAYER M1 ;
        RECT 42.064 0.656 42.096 0.688 ;
  LAYER M1 ;
        RECT 31.824 0.216 31.856 0.876 ;
  LAYER M1 ;
        RECT 31.744 0.216 31.776 0.876 ;
  LAYER M1 ;
        RECT 31.904 0.656 31.936 0.688 ;
  LAYER M1 ;
        RECT 40.784 0.3 40.816 0.96 ;
  LAYER M1 ;
        RECT 41.424 0.3 41.456 0.96 ;
  LAYER M1 ;
        RECT 40.704 0.3 40.736 0.96 ;
  LAYER M1 ;
        RECT 41.344 0.3 41.376 0.96 ;
  LAYER M1 ;
        RECT 40.864 0.3 40.896 0.96 ;
  LAYER M1 ;
        RECT 41.504 0.488 41.536 0.52 ;
  LAYER M1 ;
        RECT 39.424 0.3 39.456 0.96 ;
  LAYER M1 ;
        RECT 40.064 0.3 40.096 0.96 ;
  LAYER M1 ;
        RECT 39.344 0.3 39.376 0.96 ;
  LAYER M1 ;
        RECT 39.984 0.3 40.016 0.96 ;
  LAYER M1 ;
        RECT 39.504 0.3 39.536 0.96 ;
  LAYER M1 ;
        RECT 40.144 0.488 40.176 0.52 ;
  LAYER M1 ;
        RECT 40.928 24.24 40.96 24.312 ;
  LAYER M2 ;
        RECT 40.908 24.26 40.98 24.292 ;
  LAYER M2 ;
        RECT 38.192 24.26 40.944 24.292 ;
  LAYER M1 ;
        RECT 38.176 24.24 38.208 24.312 ;
  LAYER M2 ;
        RECT 38.156 24.26 38.228 24.292 ;
  LAYER M1 ;
        RECT 37.952 21.132 37.984 21.204 ;
  LAYER M2 ;
        RECT 37.932 21.152 38.004 21.184 ;
  LAYER M1 ;
        RECT 37.952 21.168 37.984 21.336 ;
  LAYER M1 ;
        RECT 37.952 21.3 37.984 21.372 ;
  LAYER M2 ;
        RECT 37.932 21.32 38.004 21.352 ;
  LAYER M2 ;
        RECT 37.968 21.32 38.192 21.352 ;
  LAYER M1 ;
        RECT 38.176 21.3 38.208 21.372 ;
  LAYER M2 ;
        RECT 38.156 21.32 38.228 21.352 ;
  LAYER M1 ;
        RECT 38.176 31.044 38.208 31.116 ;
  LAYER M2 ;
        RECT 38.156 31.064 38.228 31.096 ;
  LAYER M1 ;
        RECT 38.176 30.828 38.208 31.08 ;
  LAYER M1 ;
        RECT 38.176 21.336 38.208 30.828 ;
  LAYER M1 ;
        RECT 43.904 27.348 43.936 27.42 ;
  LAYER M2 ;
        RECT 43.884 27.368 43.956 27.4 ;
  LAYER M2 ;
        RECT 41.168 27.368 43.92 27.4 ;
  LAYER M1 ;
        RECT 41.152 27.348 41.184 27.42 ;
  LAYER M2 ;
        RECT 41.132 27.368 41.204 27.4 ;
  LAYER M1 ;
        RECT 41.152 31.044 41.184 31.116 ;
  LAYER M2 ;
        RECT 41.132 31.064 41.204 31.096 ;
  LAYER M1 ;
        RECT 41.152 30.828 41.184 31.08 ;
  LAYER M1 ;
        RECT 41.152 27.384 41.184 30.828 ;
  LAYER M2 ;
        RECT 38.192 31.064 41.168 31.096 ;
  LAYER M1 ;
        RECT 37.952 24.24 37.984 24.312 ;
  LAYER M2 ;
        RECT 37.932 24.26 38.004 24.292 ;
  LAYER M2 ;
        RECT 35.216 24.26 37.968 24.292 ;
  LAYER M1 ;
        RECT 35.2 24.24 35.232 24.312 ;
  LAYER M2 ;
        RECT 35.18 24.26 35.252 24.292 ;
  LAYER M1 ;
        RECT 37.952 27.348 37.984 27.42 ;
  LAYER M2 ;
        RECT 37.932 27.368 38.004 27.4 ;
  LAYER M2 ;
        RECT 35.216 27.368 37.968 27.4 ;
  LAYER M1 ;
        RECT 35.2 27.348 35.232 27.42 ;
  LAYER M2 ;
        RECT 35.18 27.368 35.252 27.4 ;
  LAYER M1 ;
        RECT 35.2 31.212 35.232 31.284 ;
  LAYER M2 ;
        RECT 35.18 31.232 35.252 31.264 ;
  LAYER M1 ;
        RECT 35.2 30.828 35.232 31.248 ;
  LAYER M1 ;
        RECT 35.2 24.276 35.232 30.828 ;
  LAYER M1 ;
        RECT 43.904 24.24 43.936 24.312 ;
  LAYER M2 ;
        RECT 43.884 24.26 43.956 24.292 ;
  LAYER M1 ;
        RECT 43.904 24.276 43.936 24.444 ;
  LAYER M1 ;
        RECT 43.904 24.408 43.936 24.48 ;
  LAYER M2 ;
        RECT 43.884 24.428 43.956 24.46 ;
  LAYER M2 ;
        RECT 43.92 24.428 44.144 24.46 ;
  LAYER M1 ;
        RECT 44.128 24.408 44.16 24.48 ;
  LAYER M2 ;
        RECT 44.108 24.428 44.18 24.46 ;
  LAYER M1 ;
        RECT 43.904 21.132 43.936 21.204 ;
  LAYER M2 ;
        RECT 43.884 21.152 43.956 21.184 ;
  LAYER M1 ;
        RECT 43.904 21.168 43.936 21.336 ;
  LAYER M1 ;
        RECT 43.904 21.3 43.936 21.372 ;
  LAYER M2 ;
        RECT 43.884 21.32 43.956 21.352 ;
  LAYER M2 ;
        RECT 43.92 21.32 44.144 21.352 ;
  LAYER M1 ;
        RECT 44.128 21.3 44.16 21.372 ;
  LAYER M2 ;
        RECT 44.108 21.32 44.18 21.352 ;
  LAYER M1 ;
        RECT 44.128 31.212 44.16 31.284 ;
  LAYER M2 ;
        RECT 44.108 31.232 44.18 31.264 ;
  LAYER M1 ;
        RECT 44.128 30.828 44.16 31.248 ;
  LAYER M1 ;
        RECT 44.128 21.336 44.16 30.828 ;
  LAYER M2 ;
        RECT 35.216 31.232 44.144 31.264 ;
  LAYER M1 ;
        RECT 40.928 27.348 40.96 27.42 ;
  LAYER M2 ;
        RECT 40.908 27.368 40.98 27.4 ;
  LAYER M2 ;
        RECT 37.968 27.368 40.944 27.4 ;
  LAYER M1 ;
        RECT 37.952 27.348 37.984 27.42 ;
  LAYER M2 ;
        RECT 37.932 27.368 38.004 27.4 ;
  LAYER M1 ;
        RECT 40.928 21.132 40.96 21.204 ;
  LAYER M2 ;
        RECT 40.908 21.152 40.98 21.184 ;
  LAYER M2 ;
        RECT 40.944 21.152 43.92 21.184 ;
  LAYER M1 ;
        RECT 43.904 21.132 43.936 21.204 ;
  LAYER M2 ;
        RECT 43.884 21.152 43.956 21.184 ;
  LAYER M1 ;
        RECT 34.976 30.456 35.008 30.528 ;
  LAYER M2 ;
        RECT 34.956 30.476 35.028 30.508 ;
  LAYER M2 ;
        RECT 32.24 30.476 34.992 30.508 ;
  LAYER M1 ;
        RECT 32.224 30.456 32.256 30.528 ;
  LAYER M2 ;
        RECT 32.204 30.476 32.276 30.508 ;
  LAYER M1 ;
        RECT 34.976 27.348 35.008 27.42 ;
  LAYER M2 ;
        RECT 34.956 27.368 35.028 27.4 ;
  LAYER M2 ;
        RECT 32.24 27.368 34.992 27.4 ;
  LAYER M1 ;
        RECT 32.224 27.348 32.256 27.42 ;
  LAYER M2 ;
        RECT 32.204 27.368 32.276 27.4 ;
  LAYER M1 ;
        RECT 34.976 24.24 35.008 24.312 ;
  LAYER M2 ;
        RECT 34.956 24.26 35.028 24.292 ;
  LAYER M2 ;
        RECT 32.24 24.26 34.992 24.292 ;
  LAYER M1 ;
        RECT 32.224 24.24 32.256 24.312 ;
  LAYER M2 ;
        RECT 32.204 24.26 32.276 24.292 ;
  LAYER M1 ;
        RECT 34.976 21.132 35.008 21.204 ;
  LAYER M2 ;
        RECT 34.956 21.152 35.028 21.184 ;
  LAYER M2 ;
        RECT 32.24 21.152 34.992 21.184 ;
  LAYER M1 ;
        RECT 32.224 21.132 32.256 21.204 ;
  LAYER M2 ;
        RECT 32.204 21.152 32.276 21.184 ;
  LAYER M1 ;
        RECT 34.976 18.024 35.008 18.096 ;
  LAYER M2 ;
        RECT 34.956 18.044 35.028 18.076 ;
  LAYER M2 ;
        RECT 32.24 18.044 34.992 18.076 ;
  LAYER M1 ;
        RECT 32.224 18.024 32.256 18.096 ;
  LAYER M2 ;
        RECT 32.204 18.044 32.276 18.076 ;
  LAYER M1 ;
        RECT 32.224 31.38 32.256 31.452 ;
  LAYER M2 ;
        RECT 32.204 31.4 32.276 31.432 ;
  LAYER M1 ;
        RECT 32.224 30.828 32.256 31.416 ;
  LAYER M1 ;
        RECT 32.224 18.06 32.256 30.828 ;
  LAYER M1 ;
        RECT 46.88 30.456 46.912 30.528 ;
  LAYER M2 ;
        RECT 46.86 30.476 46.932 30.508 ;
  LAYER M1 ;
        RECT 46.88 30.492 46.912 30.66 ;
  LAYER M1 ;
        RECT 46.88 30.624 46.912 30.696 ;
  LAYER M2 ;
        RECT 46.86 30.644 46.932 30.676 ;
  LAYER M2 ;
        RECT 46.896 30.644 47.12 30.676 ;
  LAYER M1 ;
        RECT 47.104 30.624 47.136 30.696 ;
  LAYER M2 ;
        RECT 47.084 30.644 47.156 30.676 ;
  LAYER M1 ;
        RECT 46.88 27.348 46.912 27.42 ;
  LAYER M2 ;
        RECT 46.86 27.368 46.932 27.4 ;
  LAYER M1 ;
        RECT 46.88 27.384 46.912 27.552 ;
  LAYER M1 ;
        RECT 46.88 27.516 46.912 27.588 ;
  LAYER M2 ;
        RECT 46.86 27.536 46.932 27.568 ;
  LAYER M2 ;
        RECT 46.896 27.536 47.12 27.568 ;
  LAYER M1 ;
        RECT 47.104 27.516 47.136 27.588 ;
  LAYER M2 ;
        RECT 47.084 27.536 47.156 27.568 ;
  LAYER M1 ;
        RECT 46.88 24.24 46.912 24.312 ;
  LAYER M2 ;
        RECT 46.86 24.26 46.932 24.292 ;
  LAYER M1 ;
        RECT 46.88 24.276 46.912 24.444 ;
  LAYER M1 ;
        RECT 46.88 24.408 46.912 24.48 ;
  LAYER M2 ;
        RECT 46.86 24.428 46.932 24.46 ;
  LAYER M2 ;
        RECT 46.896 24.428 47.12 24.46 ;
  LAYER M1 ;
        RECT 47.104 24.408 47.136 24.48 ;
  LAYER M2 ;
        RECT 47.084 24.428 47.156 24.46 ;
  LAYER M1 ;
        RECT 46.88 21.132 46.912 21.204 ;
  LAYER M2 ;
        RECT 46.86 21.152 46.932 21.184 ;
  LAYER M1 ;
        RECT 46.88 21.168 46.912 21.336 ;
  LAYER M1 ;
        RECT 46.88 21.3 46.912 21.372 ;
  LAYER M2 ;
        RECT 46.86 21.32 46.932 21.352 ;
  LAYER M2 ;
        RECT 46.896 21.32 47.12 21.352 ;
  LAYER M1 ;
        RECT 47.104 21.3 47.136 21.372 ;
  LAYER M2 ;
        RECT 47.084 21.32 47.156 21.352 ;
  LAYER M1 ;
        RECT 46.88 18.024 46.912 18.096 ;
  LAYER M2 ;
        RECT 46.86 18.044 46.932 18.076 ;
  LAYER M1 ;
        RECT 46.88 18.06 46.912 18.228 ;
  LAYER M1 ;
        RECT 46.88 18.192 46.912 18.264 ;
  LAYER M2 ;
        RECT 46.86 18.212 46.932 18.244 ;
  LAYER M2 ;
        RECT 46.896 18.212 47.12 18.244 ;
  LAYER M1 ;
        RECT 47.104 18.192 47.136 18.264 ;
  LAYER M2 ;
        RECT 47.084 18.212 47.156 18.244 ;
  LAYER M1 ;
        RECT 47.104 31.38 47.136 31.452 ;
  LAYER M2 ;
        RECT 47.084 31.4 47.156 31.432 ;
  LAYER M1 ;
        RECT 47.104 30.828 47.136 31.416 ;
  LAYER M1 ;
        RECT 47.104 18.228 47.136 30.828 ;
  LAYER M2 ;
        RECT 32.24 31.4 47.12 31.432 ;
  LAYER M1 ;
        RECT 37.952 30.456 37.984 30.528 ;
  LAYER M2 ;
        RECT 37.932 30.476 38.004 30.508 ;
  LAYER M2 ;
        RECT 34.992 30.476 37.968 30.508 ;
  LAYER M1 ;
        RECT 34.976 30.456 35.008 30.528 ;
  LAYER M2 ;
        RECT 34.956 30.476 35.028 30.508 ;
  LAYER M1 ;
        RECT 37.952 18.024 37.984 18.096 ;
  LAYER M2 ;
        RECT 37.932 18.044 38.004 18.076 ;
  LAYER M2 ;
        RECT 34.992 18.044 37.968 18.076 ;
  LAYER M1 ;
        RECT 34.976 18.024 35.008 18.096 ;
  LAYER M2 ;
        RECT 34.956 18.044 35.028 18.076 ;
  LAYER M1 ;
        RECT 40.928 18.024 40.96 18.096 ;
  LAYER M2 ;
        RECT 40.908 18.044 40.98 18.076 ;
  LAYER M2 ;
        RECT 37.968 18.044 40.944 18.076 ;
  LAYER M1 ;
        RECT 37.952 18.024 37.984 18.096 ;
  LAYER M2 ;
        RECT 37.932 18.044 38.004 18.076 ;
  LAYER M1 ;
        RECT 43.904 18.024 43.936 18.096 ;
  LAYER M2 ;
        RECT 43.884 18.044 43.956 18.076 ;
  LAYER M2 ;
        RECT 40.944 18.044 43.92 18.076 ;
  LAYER M1 ;
        RECT 40.928 18.024 40.96 18.096 ;
  LAYER M2 ;
        RECT 40.908 18.044 40.98 18.076 ;
  LAYER M1 ;
        RECT 43.904 30.456 43.936 30.528 ;
  LAYER M2 ;
        RECT 43.884 30.476 43.956 30.508 ;
  LAYER M2 ;
        RECT 43.92 30.476 46.896 30.508 ;
  LAYER M1 ;
        RECT 46.88 30.456 46.912 30.528 ;
  LAYER M2 ;
        RECT 46.86 30.476 46.932 30.508 ;
  LAYER M1 ;
        RECT 40.928 30.456 40.96 30.528 ;
  LAYER M2 ;
        RECT 40.908 30.476 40.98 30.508 ;
  LAYER M2 ;
        RECT 40.944 30.476 43.92 30.508 ;
  LAYER M1 ;
        RECT 43.904 30.456 43.936 30.528 ;
  LAYER M2 ;
        RECT 43.884 30.476 43.956 30.508 ;
  LAYER M1 ;
        RECT 38.56 21.804 38.592 21.876 ;
  LAYER M2 ;
        RECT 38.54 21.824 38.612 21.856 ;
  LAYER M2 ;
        RECT 38.352 21.824 38.576 21.856 ;
  LAYER M1 ;
        RECT 38.336 21.804 38.368 21.876 ;
  LAYER M2 ;
        RECT 38.316 21.824 38.388 21.856 ;
  LAYER M1 ;
        RECT 35.584 18.696 35.616 18.768 ;
  LAYER M2 ;
        RECT 35.564 18.716 35.636 18.748 ;
  LAYER M1 ;
        RECT 35.584 18.564 35.616 18.732 ;
  LAYER M1 ;
        RECT 35.584 18.528 35.616 18.6 ;
  LAYER M2 ;
        RECT 35.564 18.548 35.636 18.58 ;
  LAYER M2 ;
        RECT 35.6 18.548 38.352 18.58 ;
  LAYER M1 ;
        RECT 38.336 18.528 38.368 18.6 ;
  LAYER M2 ;
        RECT 38.316 18.548 38.388 18.58 ;
  LAYER M1 ;
        RECT 38.336 15 38.368 15.072 ;
  LAYER M2 ;
        RECT 38.316 15.02 38.388 15.052 ;
  LAYER M1 ;
        RECT 38.336 15.036 38.368 15.288 ;
  LAYER M1 ;
        RECT 38.336 15.288 38.368 21.84 ;
  LAYER M1 ;
        RECT 41.536 24.912 41.568 24.984 ;
  LAYER M2 ;
        RECT 41.516 24.932 41.588 24.964 ;
  LAYER M2 ;
        RECT 41.328 24.932 41.552 24.964 ;
  LAYER M1 ;
        RECT 41.312 24.912 41.344 24.984 ;
  LAYER M2 ;
        RECT 41.292 24.932 41.364 24.964 ;
  LAYER M1 ;
        RECT 41.312 15 41.344 15.072 ;
  LAYER M2 ;
        RECT 41.292 15.02 41.364 15.052 ;
  LAYER M1 ;
        RECT 41.312 15.036 41.344 15.288 ;
  LAYER M1 ;
        RECT 41.312 15.288 41.344 24.948 ;
  LAYER M2 ;
        RECT 38.352 15.02 41.328 15.052 ;
  LAYER M1 ;
        RECT 35.584 21.804 35.616 21.876 ;
  LAYER M2 ;
        RECT 35.564 21.824 35.636 21.856 ;
  LAYER M2 ;
        RECT 35.376 21.824 35.6 21.856 ;
  LAYER M1 ;
        RECT 35.36 21.804 35.392 21.876 ;
  LAYER M2 ;
        RECT 35.34 21.824 35.412 21.856 ;
  LAYER M1 ;
        RECT 35.584 24.912 35.616 24.984 ;
  LAYER M2 ;
        RECT 35.564 24.932 35.636 24.964 ;
  LAYER M2 ;
        RECT 35.376 24.932 35.6 24.964 ;
  LAYER M1 ;
        RECT 35.36 24.912 35.392 24.984 ;
  LAYER M2 ;
        RECT 35.34 24.932 35.412 24.964 ;
  LAYER M1 ;
        RECT 35.36 14.832 35.392 14.904 ;
  LAYER M2 ;
        RECT 35.34 14.852 35.412 14.884 ;
  LAYER M1 ;
        RECT 35.36 14.868 35.392 15.288 ;
  LAYER M1 ;
        RECT 35.36 15.288 35.392 24.948 ;
  LAYER M1 ;
        RECT 41.536 21.804 41.568 21.876 ;
  LAYER M2 ;
        RECT 41.516 21.824 41.588 21.856 ;
  LAYER M1 ;
        RECT 41.536 21.672 41.568 21.84 ;
  LAYER M1 ;
        RECT 41.536 21.636 41.568 21.708 ;
  LAYER M2 ;
        RECT 41.516 21.656 41.588 21.688 ;
  LAYER M2 ;
        RECT 41.552 21.656 44.304 21.688 ;
  LAYER M1 ;
        RECT 44.288 21.636 44.32 21.708 ;
  LAYER M2 ;
        RECT 44.268 21.656 44.34 21.688 ;
  LAYER M1 ;
        RECT 41.536 18.696 41.568 18.768 ;
  LAYER M2 ;
        RECT 41.516 18.716 41.588 18.748 ;
  LAYER M1 ;
        RECT 41.536 18.564 41.568 18.732 ;
  LAYER M1 ;
        RECT 41.536 18.528 41.568 18.6 ;
  LAYER M2 ;
        RECT 41.516 18.548 41.588 18.58 ;
  LAYER M2 ;
        RECT 41.552 18.548 44.304 18.58 ;
  LAYER M1 ;
        RECT 44.288 18.528 44.32 18.6 ;
  LAYER M2 ;
        RECT 44.268 18.548 44.34 18.58 ;
  LAYER M1 ;
        RECT 44.288 14.832 44.32 14.904 ;
  LAYER M2 ;
        RECT 44.268 14.852 44.34 14.884 ;
  LAYER M1 ;
        RECT 44.288 14.868 44.32 15.288 ;
  LAYER M1 ;
        RECT 44.288 15.288 44.32 21.672 ;
  LAYER M2 ;
        RECT 35.376 14.852 44.304 14.884 ;
  LAYER M1 ;
        RECT 38.56 24.912 38.592 24.984 ;
  LAYER M2 ;
        RECT 38.54 24.932 38.612 24.964 ;
  LAYER M2 ;
        RECT 35.6 24.932 38.576 24.964 ;
  LAYER M1 ;
        RECT 35.584 24.912 35.616 24.984 ;
  LAYER M2 ;
        RECT 35.564 24.932 35.636 24.964 ;
  LAYER M1 ;
        RECT 38.56 18.696 38.592 18.768 ;
  LAYER M2 ;
        RECT 38.54 18.716 38.612 18.748 ;
  LAYER M2 ;
        RECT 38.576 18.716 41.552 18.748 ;
  LAYER M1 ;
        RECT 41.536 18.696 41.568 18.768 ;
  LAYER M2 ;
        RECT 41.516 18.716 41.588 18.748 ;
  LAYER M1 ;
        RECT 32.608 28.02 32.64 28.092 ;
  LAYER M2 ;
        RECT 32.588 28.04 32.66 28.072 ;
  LAYER M2 ;
        RECT 32.4 28.04 32.624 28.072 ;
  LAYER M1 ;
        RECT 32.384 28.02 32.416 28.092 ;
  LAYER M2 ;
        RECT 32.364 28.04 32.436 28.072 ;
  LAYER M1 ;
        RECT 32.608 24.912 32.64 24.984 ;
  LAYER M2 ;
        RECT 32.588 24.932 32.66 24.964 ;
  LAYER M2 ;
        RECT 32.4 24.932 32.624 24.964 ;
  LAYER M1 ;
        RECT 32.384 24.912 32.416 24.984 ;
  LAYER M2 ;
        RECT 32.364 24.932 32.436 24.964 ;
  LAYER M1 ;
        RECT 32.608 21.804 32.64 21.876 ;
  LAYER M2 ;
        RECT 32.588 21.824 32.66 21.856 ;
  LAYER M2 ;
        RECT 32.4 21.824 32.624 21.856 ;
  LAYER M1 ;
        RECT 32.384 21.804 32.416 21.876 ;
  LAYER M2 ;
        RECT 32.364 21.824 32.436 21.856 ;
  LAYER M1 ;
        RECT 32.608 18.696 32.64 18.768 ;
  LAYER M2 ;
        RECT 32.588 18.716 32.66 18.748 ;
  LAYER M2 ;
        RECT 32.4 18.716 32.624 18.748 ;
  LAYER M1 ;
        RECT 32.384 18.696 32.416 18.768 ;
  LAYER M2 ;
        RECT 32.364 18.716 32.436 18.748 ;
  LAYER M1 ;
        RECT 32.608 15.588 32.64 15.66 ;
  LAYER M2 ;
        RECT 32.588 15.608 32.66 15.64 ;
  LAYER M2 ;
        RECT 32.4 15.608 32.624 15.64 ;
  LAYER M1 ;
        RECT 32.384 15.588 32.416 15.66 ;
  LAYER M2 ;
        RECT 32.364 15.608 32.436 15.64 ;
  LAYER M1 ;
        RECT 32.384 14.664 32.416 14.736 ;
  LAYER M2 ;
        RECT 32.364 14.684 32.436 14.716 ;
  LAYER M1 ;
        RECT 32.384 14.7 32.416 15.288 ;
  LAYER M1 ;
        RECT 32.384 15.288 32.416 28.056 ;
  LAYER M1 ;
        RECT 44.512 28.02 44.544 28.092 ;
  LAYER M2 ;
        RECT 44.492 28.04 44.564 28.072 ;
  LAYER M1 ;
        RECT 44.512 27.888 44.544 28.056 ;
  LAYER M1 ;
        RECT 44.512 27.852 44.544 27.924 ;
  LAYER M2 ;
        RECT 44.492 27.872 44.564 27.904 ;
  LAYER M2 ;
        RECT 44.528 27.872 47.28 27.904 ;
  LAYER M1 ;
        RECT 47.264 27.852 47.296 27.924 ;
  LAYER M2 ;
        RECT 47.244 27.872 47.316 27.904 ;
  LAYER M1 ;
        RECT 44.512 24.912 44.544 24.984 ;
  LAYER M2 ;
        RECT 44.492 24.932 44.564 24.964 ;
  LAYER M1 ;
        RECT 44.512 24.78 44.544 24.948 ;
  LAYER M1 ;
        RECT 44.512 24.744 44.544 24.816 ;
  LAYER M2 ;
        RECT 44.492 24.764 44.564 24.796 ;
  LAYER M2 ;
        RECT 44.528 24.764 47.28 24.796 ;
  LAYER M1 ;
        RECT 47.264 24.744 47.296 24.816 ;
  LAYER M2 ;
        RECT 47.244 24.764 47.316 24.796 ;
  LAYER M1 ;
        RECT 44.512 21.804 44.544 21.876 ;
  LAYER M2 ;
        RECT 44.492 21.824 44.564 21.856 ;
  LAYER M1 ;
        RECT 44.512 21.672 44.544 21.84 ;
  LAYER M1 ;
        RECT 44.512 21.636 44.544 21.708 ;
  LAYER M2 ;
        RECT 44.492 21.656 44.564 21.688 ;
  LAYER M2 ;
        RECT 44.528 21.656 47.28 21.688 ;
  LAYER M1 ;
        RECT 47.264 21.636 47.296 21.708 ;
  LAYER M2 ;
        RECT 47.244 21.656 47.316 21.688 ;
  LAYER M1 ;
        RECT 44.512 18.696 44.544 18.768 ;
  LAYER M2 ;
        RECT 44.492 18.716 44.564 18.748 ;
  LAYER M1 ;
        RECT 44.512 18.564 44.544 18.732 ;
  LAYER M1 ;
        RECT 44.512 18.528 44.544 18.6 ;
  LAYER M2 ;
        RECT 44.492 18.548 44.564 18.58 ;
  LAYER M2 ;
        RECT 44.528 18.548 47.28 18.58 ;
  LAYER M1 ;
        RECT 47.264 18.528 47.296 18.6 ;
  LAYER M2 ;
        RECT 47.244 18.548 47.316 18.58 ;
  LAYER M1 ;
        RECT 44.512 15.588 44.544 15.66 ;
  LAYER M2 ;
        RECT 44.492 15.608 44.564 15.64 ;
  LAYER M1 ;
        RECT 44.512 15.456 44.544 15.624 ;
  LAYER M1 ;
        RECT 44.512 15.42 44.544 15.492 ;
  LAYER M2 ;
        RECT 44.492 15.44 44.564 15.472 ;
  LAYER M2 ;
        RECT 44.528 15.44 47.28 15.472 ;
  LAYER M1 ;
        RECT 47.264 15.42 47.296 15.492 ;
  LAYER M2 ;
        RECT 47.244 15.44 47.316 15.472 ;
  LAYER M1 ;
        RECT 47.264 14.664 47.296 14.736 ;
  LAYER M2 ;
        RECT 47.244 14.684 47.316 14.716 ;
  LAYER M1 ;
        RECT 47.264 14.7 47.296 15.288 ;
  LAYER M1 ;
        RECT 47.264 15.288 47.296 27.888 ;
  LAYER M2 ;
        RECT 32.4 14.684 47.28 14.716 ;
  LAYER M1 ;
        RECT 35.584 28.02 35.616 28.092 ;
  LAYER M2 ;
        RECT 35.564 28.04 35.636 28.072 ;
  LAYER M2 ;
        RECT 32.624 28.04 35.6 28.072 ;
  LAYER M1 ;
        RECT 32.608 28.02 32.64 28.092 ;
  LAYER M2 ;
        RECT 32.588 28.04 32.66 28.072 ;
  LAYER M1 ;
        RECT 35.584 15.588 35.616 15.66 ;
  LAYER M2 ;
        RECT 35.564 15.608 35.636 15.64 ;
  LAYER M2 ;
        RECT 32.624 15.608 35.6 15.64 ;
  LAYER M1 ;
        RECT 32.608 15.588 32.64 15.66 ;
  LAYER M2 ;
        RECT 32.588 15.608 32.66 15.64 ;
  LAYER M1 ;
        RECT 38.56 15.588 38.592 15.66 ;
  LAYER M2 ;
        RECT 38.54 15.608 38.612 15.64 ;
  LAYER M2 ;
        RECT 35.6 15.608 38.576 15.64 ;
  LAYER M1 ;
        RECT 35.584 15.588 35.616 15.66 ;
  LAYER M2 ;
        RECT 35.564 15.608 35.636 15.64 ;
  LAYER M1 ;
        RECT 41.536 15.588 41.568 15.66 ;
  LAYER M2 ;
        RECT 41.516 15.608 41.588 15.64 ;
  LAYER M2 ;
        RECT 38.576 15.608 41.552 15.64 ;
  LAYER M1 ;
        RECT 38.56 15.588 38.592 15.66 ;
  LAYER M2 ;
        RECT 38.54 15.608 38.612 15.64 ;
  LAYER M1 ;
        RECT 41.536 28.02 41.568 28.092 ;
  LAYER M2 ;
        RECT 41.516 28.04 41.588 28.072 ;
  LAYER M2 ;
        RECT 41.552 28.04 44.528 28.072 ;
  LAYER M1 ;
        RECT 44.512 28.02 44.544 28.092 ;
  LAYER M2 ;
        RECT 44.492 28.04 44.564 28.072 ;
  LAYER M1 ;
        RECT 38.56 28.02 38.592 28.092 ;
  LAYER M2 ;
        RECT 38.54 28.04 38.612 28.072 ;
  LAYER M2 ;
        RECT 38.576 28.04 41.552 28.072 ;
  LAYER M1 ;
        RECT 41.536 28.02 41.568 28.092 ;
  LAYER M2 ;
        RECT 41.516 28.04 41.588 28.072 ;
  LAYER M1 ;
        RECT 32.608 28.02 32.64 30.528 ;
  LAYER M3 ;
        RECT 32.608 28.04 32.64 28.072 ;
  LAYER M1 ;
        RECT 32.672 28.02 32.704 30.528 ;
  LAYER M3 ;
        RECT 32.672 30.476 32.704 30.508 ;
  LAYER M1 ;
        RECT 32.736 28.02 32.768 30.528 ;
  LAYER M3 ;
        RECT 32.736 28.04 32.768 28.072 ;
  LAYER M1 ;
        RECT 32.8 28.02 32.832 30.528 ;
  LAYER M3 ;
        RECT 32.8 30.476 32.832 30.508 ;
  LAYER M1 ;
        RECT 32.864 28.02 32.896 30.528 ;
  LAYER M3 ;
        RECT 32.864 28.04 32.896 28.072 ;
  LAYER M1 ;
        RECT 32.928 28.02 32.96 30.528 ;
  LAYER M3 ;
        RECT 32.928 30.476 32.96 30.508 ;
  LAYER M1 ;
        RECT 32.992 28.02 33.024 30.528 ;
  LAYER M3 ;
        RECT 32.992 28.04 33.024 28.072 ;
  LAYER M1 ;
        RECT 33.056 28.02 33.088 30.528 ;
  LAYER M3 ;
        RECT 33.056 30.476 33.088 30.508 ;
  LAYER M1 ;
        RECT 33.12 28.02 33.152 30.528 ;
  LAYER M3 ;
        RECT 33.12 28.04 33.152 28.072 ;
  LAYER M1 ;
        RECT 33.184 28.02 33.216 30.528 ;
  LAYER M3 ;
        RECT 33.184 30.476 33.216 30.508 ;
  LAYER M1 ;
        RECT 33.248 28.02 33.28 30.528 ;
  LAYER M3 ;
        RECT 33.248 28.04 33.28 28.072 ;
  LAYER M1 ;
        RECT 33.312 28.02 33.344 30.528 ;
  LAYER M3 ;
        RECT 33.312 30.476 33.344 30.508 ;
  LAYER M1 ;
        RECT 33.376 28.02 33.408 30.528 ;
  LAYER M3 ;
        RECT 33.376 28.04 33.408 28.072 ;
  LAYER M1 ;
        RECT 33.44 28.02 33.472 30.528 ;
  LAYER M3 ;
        RECT 33.44 30.476 33.472 30.508 ;
  LAYER M1 ;
        RECT 33.504 28.02 33.536 30.528 ;
  LAYER M3 ;
        RECT 33.504 28.04 33.536 28.072 ;
  LAYER M1 ;
        RECT 33.568 28.02 33.6 30.528 ;
  LAYER M3 ;
        RECT 33.568 30.476 33.6 30.508 ;
  LAYER M1 ;
        RECT 33.632 28.02 33.664 30.528 ;
  LAYER M3 ;
        RECT 33.632 28.04 33.664 28.072 ;
  LAYER M1 ;
        RECT 33.696 28.02 33.728 30.528 ;
  LAYER M3 ;
        RECT 33.696 30.476 33.728 30.508 ;
  LAYER M1 ;
        RECT 33.76 28.02 33.792 30.528 ;
  LAYER M3 ;
        RECT 33.76 28.04 33.792 28.072 ;
  LAYER M1 ;
        RECT 33.824 28.02 33.856 30.528 ;
  LAYER M3 ;
        RECT 33.824 30.476 33.856 30.508 ;
  LAYER M1 ;
        RECT 33.888 28.02 33.92 30.528 ;
  LAYER M3 ;
        RECT 33.888 28.04 33.92 28.072 ;
  LAYER M1 ;
        RECT 33.952 28.02 33.984 30.528 ;
  LAYER M3 ;
        RECT 33.952 30.476 33.984 30.508 ;
  LAYER M1 ;
        RECT 34.016 28.02 34.048 30.528 ;
  LAYER M3 ;
        RECT 34.016 28.04 34.048 28.072 ;
  LAYER M1 ;
        RECT 34.08 28.02 34.112 30.528 ;
  LAYER M3 ;
        RECT 34.08 30.476 34.112 30.508 ;
  LAYER M1 ;
        RECT 34.144 28.02 34.176 30.528 ;
  LAYER M3 ;
        RECT 34.144 28.04 34.176 28.072 ;
  LAYER M1 ;
        RECT 34.208 28.02 34.24 30.528 ;
  LAYER M3 ;
        RECT 34.208 30.476 34.24 30.508 ;
  LAYER M1 ;
        RECT 34.272 28.02 34.304 30.528 ;
  LAYER M3 ;
        RECT 34.272 28.04 34.304 28.072 ;
  LAYER M1 ;
        RECT 34.336 28.02 34.368 30.528 ;
  LAYER M3 ;
        RECT 34.336 30.476 34.368 30.508 ;
  LAYER M1 ;
        RECT 34.4 28.02 34.432 30.528 ;
  LAYER M3 ;
        RECT 34.4 28.04 34.432 28.072 ;
  LAYER M1 ;
        RECT 34.464 28.02 34.496 30.528 ;
  LAYER M3 ;
        RECT 34.464 30.476 34.496 30.508 ;
  LAYER M1 ;
        RECT 34.528 28.02 34.56 30.528 ;
  LAYER M3 ;
        RECT 34.528 28.04 34.56 28.072 ;
  LAYER M1 ;
        RECT 34.592 28.02 34.624 30.528 ;
  LAYER M3 ;
        RECT 34.592 30.476 34.624 30.508 ;
  LAYER M1 ;
        RECT 34.656 28.02 34.688 30.528 ;
  LAYER M3 ;
        RECT 34.656 28.04 34.688 28.072 ;
  LAYER M1 ;
        RECT 34.72 28.02 34.752 30.528 ;
  LAYER M3 ;
        RECT 34.72 30.476 34.752 30.508 ;
  LAYER M1 ;
        RECT 34.784 28.02 34.816 30.528 ;
  LAYER M3 ;
        RECT 34.784 28.04 34.816 28.072 ;
  LAYER M1 ;
        RECT 34.848 28.02 34.88 30.528 ;
  LAYER M3 ;
        RECT 34.848 30.476 34.88 30.508 ;
  LAYER M1 ;
        RECT 34.912 28.02 34.944 30.528 ;
  LAYER M3 ;
        RECT 34.912 28.04 34.944 28.072 ;
  LAYER M1 ;
        RECT 34.976 28.02 35.008 30.528 ;
  LAYER M3 ;
        RECT 32.608 30.412 32.64 30.444 ;
  LAYER M2 ;
        RECT 34.976 30.348 35.008 30.38 ;
  LAYER M2 ;
        RECT 32.608 30.284 32.64 30.316 ;
  LAYER M2 ;
        RECT 34.976 30.22 35.008 30.252 ;
  LAYER M2 ;
        RECT 32.608 30.156 32.64 30.188 ;
  LAYER M2 ;
        RECT 34.976 30.092 35.008 30.124 ;
  LAYER M2 ;
        RECT 32.608 30.028 32.64 30.06 ;
  LAYER M2 ;
        RECT 34.976 29.964 35.008 29.996 ;
  LAYER M2 ;
        RECT 32.608 29.9 32.64 29.932 ;
  LAYER M2 ;
        RECT 34.976 29.836 35.008 29.868 ;
  LAYER M2 ;
        RECT 32.608 29.772 32.64 29.804 ;
  LAYER M2 ;
        RECT 34.976 29.708 35.008 29.74 ;
  LAYER M2 ;
        RECT 32.608 29.644 32.64 29.676 ;
  LAYER M2 ;
        RECT 34.976 29.58 35.008 29.612 ;
  LAYER M2 ;
        RECT 32.608 29.516 32.64 29.548 ;
  LAYER M2 ;
        RECT 34.976 29.452 35.008 29.484 ;
  LAYER M2 ;
        RECT 32.608 29.388 32.64 29.42 ;
  LAYER M2 ;
        RECT 34.976 29.324 35.008 29.356 ;
  LAYER M2 ;
        RECT 32.608 29.26 32.64 29.292 ;
  LAYER M2 ;
        RECT 34.976 29.196 35.008 29.228 ;
  LAYER M2 ;
        RECT 32.608 29.132 32.64 29.164 ;
  LAYER M2 ;
        RECT 34.976 29.068 35.008 29.1 ;
  LAYER M2 ;
        RECT 32.608 29.004 32.64 29.036 ;
  LAYER M2 ;
        RECT 34.976 28.94 35.008 28.972 ;
  LAYER M2 ;
        RECT 32.608 28.876 32.64 28.908 ;
  LAYER M2 ;
        RECT 34.976 28.812 35.008 28.844 ;
  LAYER M2 ;
        RECT 32.608 28.748 32.64 28.78 ;
  LAYER M2 ;
        RECT 34.976 28.684 35.008 28.716 ;
  LAYER M2 ;
        RECT 32.608 28.62 32.64 28.652 ;
  LAYER M2 ;
        RECT 34.976 28.556 35.008 28.588 ;
  LAYER M2 ;
        RECT 32.608 28.492 32.64 28.524 ;
  LAYER M2 ;
        RECT 34.976 28.428 35.008 28.46 ;
  LAYER M2 ;
        RECT 32.608 28.364 32.64 28.396 ;
  LAYER M2 ;
        RECT 34.976 28.3 35.008 28.332 ;
  LAYER M2 ;
        RECT 32.608 28.236 32.64 28.268 ;
  LAYER M2 ;
        RECT 34.976 28.172 35.008 28.204 ;
  LAYER M2 ;
        RECT 32.56 27.972 35.056 30.576 ;
  LAYER M1 ;
        RECT 32.608 24.912 32.64 27.42 ;
  LAYER M3 ;
        RECT 32.608 24.932 32.64 24.964 ;
  LAYER M1 ;
        RECT 32.672 24.912 32.704 27.42 ;
  LAYER M3 ;
        RECT 32.672 27.368 32.704 27.4 ;
  LAYER M1 ;
        RECT 32.736 24.912 32.768 27.42 ;
  LAYER M3 ;
        RECT 32.736 24.932 32.768 24.964 ;
  LAYER M1 ;
        RECT 32.8 24.912 32.832 27.42 ;
  LAYER M3 ;
        RECT 32.8 27.368 32.832 27.4 ;
  LAYER M1 ;
        RECT 32.864 24.912 32.896 27.42 ;
  LAYER M3 ;
        RECT 32.864 24.932 32.896 24.964 ;
  LAYER M1 ;
        RECT 32.928 24.912 32.96 27.42 ;
  LAYER M3 ;
        RECT 32.928 27.368 32.96 27.4 ;
  LAYER M1 ;
        RECT 32.992 24.912 33.024 27.42 ;
  LAYER M3 ;
        RECT 32.992 24.932 33.024 24.964 ;
  LAYER M1 ;
        RECT 33.056 24.912 33.088 27.42 ;
  LAYER M3 ;
        RECT 33.056 27.368 33.088 27.4 ;
  LAYER M1 ;
        RECT 33.12 24.912 33.152 27.42 ;
  LAYER M3 ;
        RECT 33.12 24.932 33.152 24.964 ;
  LAYER M1 ;
        RECT 33.184 24.912 33.216 27.42 ;
  LAYER M3 ;
        RECT 33.184 27.368 33.216 27.4 ;
  LAYER M1 ;
        RECT 33.248 24.912 33.28 27.42 ;
  LAYER M3 ;
        RECT 33.248 24.932 33.28 24.964 ;
  LAYER M1 ;
        RECT 33.312 24.912 33.344 27.42 ;
  LAYER M3 ;
        RECT 33.312 27.368 33.344 27.4 ;
  LAYER M1 ;
        RECT 33.376 24.912 33.408 27.42 ;
  LAYER M3 ;
        RECT 33.376 24.932 33.408 24.964 ;
  LAYER M1 ;
        RECT 33.44 24.912 33.472 27.42 ;
  LAYER M3 ;
        RECT 33.44 27.368 33.472 27.4 ;
  LAYER M1 ;
        RECT 33.504 24.912 33.536 27.42 ;
  LAYER M3 ;
        RECT 33.504 24.932 33.536 24.964 ;
  LAYER M1 ;
        RECT 33.568 24.912 33.6 27.42 ;
  LAYER M3 ;
        RECT 33.568 27.368 33.6 27.4 ;
  LAYER M1 ;
        RECT 33.632 24.912 33.664 27.42 ;
  LAYER M3 ;
        RECT 33.632 24.932 33.664 24.964 ;
  LAYER M1 ;
        RECT 33.696 24.912 33.728 27.42 ;
  LAYER M3 ;
        RECT 33.696 27.368 33.728 27.4 ;
  LAYER M1 ;
        RECT 33.76 24.912 33.792 27.42 ;
  LAYER M3 ;
        RECT 33.76 24.932 33.792 24.964 ;
  LAYER M1 ;
        RECT 33.824 24.912 33.856 27.42 ;
  LAYER M3 ;
        RECT 33.824 27.368 33.856 27.4 ;
  LAYER M1 ;
        RECT 33.888 24.912 33.92 27.42 ;
  LAYER M3 ;
        RECT 33.888 24.932 33.92 24.964 ;
  LAYER M1 ;
        RECT 33.952 24.912 33.984 27.42 ;
  LAYER M3 ;
        RECT 33.952 27.368 33.984 27.4 ;
  LAYER M1 ;
        RECT 34.016 24.912 34.048 27.42 ;
  LAYER M3 ;
        RECT 34.016 24.932 34.048 24.964 ;
  LAYER M1 ;
        RECT 34.08 24.912 34.112 27.42 ;
  LAYER M3 ;
        RECT 34.08 27.368 34.112 27.4 ;
  LAYER M1 ;
        RECT 34.144 24.912 34.176 27.42 ;
  LAYER M3 ;
        RECT 34.144 24.932 34.176 24.964 ;
  LAYER M1 ;
        RECT 34.208 24.912 34.24 27.42 ;
  LAYER M3 ;
        RECT 34.208 27.368 34.24 27.4 ;
  LAYER M1 ;
        RECT 34.272 24.912 34.304 27.42 ;
  LAYER M3 ;
        RECT 34.272 24.932 34.304 24.964 ;
  LAYER M1 ;
        RECT 34.336 24.912 34.368 27.42 ;
  LAYER M3 ;
        RECT 34.336 27.368 34.368 27.4 ;
  LAYER M1 ;
        RECT 34.4 24.912 34.432 27.42 ;
  LAYER M3 ;
        RECT 34.4 24.932 34.432 24.964 ;
  LAYER M1 ;
        RECT 34.464 24.912 34.496 27.42 ;
  LAYER M3 ;
        RECT 34.464 27.368 34.496 27.4 ;
  LAYER M1 ;
        RECT 34.528 24.912 34.56 27.42 ;
  LAYER M3 ;
        RECT 34.528 24.932 34.56 24.964 ;
  LAYER M1 ;
        RECT 34.592 24.912 34.624 27.42 ;
  LAYER M3 ;
        RECT 34.592 27.368 34.624 27.4 ;
  LAYER M1 ;
        RECT 34.656 24.912 34.688 27.42 ;
  LAYER M3 ;
        RECT 34.656 24.932 34.688 24.964 ;
  LAYER M1 ;
        RECT 34.72 24.912 34.752 27.42 ;
  LAYER M3 ;
        RECT 34.72 27.368 34.752 27.4 ;
  LAYER M1 ;
        RECT 34.784 24.912 34.816 27.42 ;
  LAYER M3 ;
        RECT 34.784 24.932 34.816 24.964 ;
  LAYER M1 ;
        RECT 34.848 24.912 34.88 27.42 ;
  LAYER M3 ;
        RECT 34.848 27.368 34.88 27.4 ;
  LAYER M1 ;
        RECT 34.912 24.912 34.944 27.42 ;
  LAYER M3 ;
        RECT 34.912 24.932 34.944 24.964 ;
  LAYER M1 ;
        RECT 34.976 24.912 35.008 27.42 ;
  LAYER M3 ;
        RECT 32.608 27.304 32.64 27.336 ;
  LAYER M2 ;
        RECT 34.976 27.24 35.008 27.272 ;
  LAYER M2 ;
        RECT 32.608 27.176 32.64 27.208 ;
  LAYER M2 ;
        RECT 34.976 27.112 35.008 27.144 ;
  LAYER M2 ;
        RECT 32.608 27.048 32.64 27.08 ;
  LAYER M2 ;
        RECT 34.976 26.984 35.008 27.016 ;
  LAYER M2 ;
        RECT 32.608 26.92 32.64 26.952 ;
  LAYER M2 ;
        RECT 34.976 26.856 35.008 26.888 ;
  LAYER M2 ;
        RECT 32.608 26.792 32.64 26.824 ;
  LAYER M2 ;
        RECT 34.976 26.728 35.008 26.76 ;
  LAYER M2 ;
        RECT 32.608 26.664 32.64 26.696 ;
  LAYER M2 ;
        RECT 34.976 26.6 35.008 26.632 ;
  LAYER M2 ;
        RECT 32.608 26.536 32.64 26.568 ;
  LAYER M2 ;
        RECT 34.976 26.472 35.008 26.504 ;
  LAYER M2 ;
        RECT 32.608 26.408 32.64 26.44 ;
  LAYER M2 ;
        RECT 34.976 26.344 35.008 26.376 ;
  LAYER M2 ;
        RECT 32.608 26.28 32.64 26.312 ;
  LAYER M2 ;
        RECT 34.976 26.216 35.008 26.248 ;
  LAYER M2 ;
        RECT 32.608 26.152 32.64 26.184 ;
  LAYER M2 ;
        RECT 34.976 26.088 35.008 26.12 ;
  LAYER M2 ;
        RECT 32.608 26.024 32.64 26.056 ;
  LAYER M2 ;
        RECT 34.976 25.96 35.008 25.992 ;
  LAYER M2 ;
        RECT 32.608 25.896 32.64 25.928 ;
  LAYER M2 ;
        RECT 34.976 25.832 35.008 25.864 ;
  LAYER M2 ;
        RECT 32.608 25.768 32.64 25.8 ;
  LAYER M2 ;
        RECT 34.976 25.704 35.008 25.736 ;
  LAYER M2 ;
        RECT 32.608 25.64 32.64 25.672 ;
  LAYER M2 ;
        RECT 34.976 25.576 35.008 25.608 ;
  LAYER M2 ;
        RECT 32.608 25.512 32.64 25.544 ;
  LAYER M2 ;
        RECT 34.976 25.448 35.008 25.48 ;
  LAYER M2 ;
        RECT 32.608 25.384 32.64 25.416 ;
  LAYER M2 ;
        RECT 34.976 25.32 35.008 25.352 ;
  LAYER M2 ;
        RECT 32.608 25.256 32.64 25.288 ;
  LAYER M2 ;
        RECT 34.976 25.192 35.008 25.224 ;
  LAYER M2 ;
        RECT 32.608 25.128 32.64 25.16 ;
  LAYER M2 ;
        RECT 34.976 25.064 35.008 25.096 ;
  LAYER M2 ;
        RECT 32.56 24.864 35.056 27.468 ;
  LAYER M1 ;
        RECT 32.608 21.804 32.64 24.312 ;
  LAYER M3 ;
        RECT 32.608 21.824 32.64 21.856 ;
  LAYER M1 ;
        RECT 32.672 21.804 32.704 24.312 ;
  LAYER M3 ;
        RECT 32.672 24.26 32.704 24.292 ;
  LAYER M1 ;
        RECT 32.736 21.804 32.768 24.312 ;
  LAYER M3 ;
        RECT 32.736 21.824 32.768 21.856 ;
  LAYER M1 ;
        RECT 32.8 21.804 32.832 24.312 ;
  LAYER M3 ;
        RECT 32.8 24.26 32.832 24.292 ;
  LAYER M1 ;
        RECT 32.864 21.804 32.896 24.312 ;
  LAYER M3 ;
        RECT 32.864 21.824 32.896 21.856 ;
  LAYER M1 ;
        RECT 32.928 21.804 32.96 24.312 ;
  LAYER M3 ;
        RECT 32.928 24.26 32.96 24.292 ;
  LAYER M1 ;
        RECT 32.992 21.804 33.024 24.312 ;
  LAYER M3 ;
        RECT 32.992 21.824 33.024 21.856 ;
  LAYER M1 ;
        RECT 33.056 21.804 33.088 24.312 ;
  LAYER M3 ;
        RECT 33.056 24.26 33.088 24.292 ;
  LAYER M1 ;
        RECT 33.12 21.804 33.152 24.312 ;
  LAYER M3 ;
        RECT 33.12 21.824 33.152 21.856 ;
  LAYER M1 ;
        RECT 33.184 21.804 33.216 24.312 ;
  LAYER M3 ;
        RECT 33.184 24.26 33.216 24.292 ;
  LAYER M1 ;
        RECT 33.248 21.804 33.28 24.312 ;
  LAYER M3 ;
        RECT 33.248 21.824 33.28 21.856 ;
  LAYER M1 ;
        RECT 33.312 21.804 33.344 24.312 ;
  LAYER M3 ;
        RECT 33.312 24.26 33.344 24.292 ;
  LAYER M1 ;
        RECT 33.376 21.804 33.408 24.312 ;
  LAYER M3 ;
        RECT 33.376 21.824 33.408 21.856 ;
  LAYER M1 ;
        RECT 33.44 21.804 33.472 24.312 ;
  LAYER M3 ;
        RECT 33.44 24.26 33.472 24.292 ;
  LAYER M1 ;
        RECT 33.504 21.804 33.536 24.312 ;
  LAYER M3 ;
        RECT 33.504 21.824 33.536 21.856 ;
  LAYER M1 ;
        RECT 33.568 21.804 33.6 24.312 ;
  LAYER M3 ;
        RECT 33.568 24.26 33.6 24.292 ;
  LAYER M1 ;
        RECT 33.632 21.804 33.664 24.312 ;
  LAYER M3 ;
        RECT 33.632 21.824 33.664 21.856 ;
  LAYER M1 ;
        RECT 33.696 21.804 33.728 24.312 ;
  LAYER M3 ;
        RECT 33.696 24.26 33.728 24.292 ;
  LAYER M1 ;
        RECT 33.76 21.804 33.792 24.312 ;
  LAYER M3 ;
        RECT 33.76 21.824 33.792 21.856 ;
  LAYER M1 ;
        RECT 33.824 21.804 33.856 24.312 ;
  LAYER M3 ;
        RECT 33.824 24.26 33.856 24.292 ;
  LAYER M1 ;
        RECT 33.888 21.804 33.92 24.312 ;
  LAYER M3 ;
        RECT 33.888 21.824 33.92 21.856 ;
  LAYER M1 ;
        RECT 33.952 21.804 33.984 24.312 ;
  LAYER M3 ;
        RECT 33.952 24.26 33.984 24.292 ;
  LAYER M1 ;
        RECT 34.016 21.804 34.048 24.312 ;
  LAYER M3 ;
        RECT 34.016 21.824 34.048 21.856 ;
  LAYER M1 ;
        RECT 34.08 21.804 34.112 24.312 ;
  LAYER M3 ;
        RECT 34.08 24.26 34.112 24.292 ;
  LAYER M1 ;
        RECT 34.144 21.804 34.176 24.312 ;
  LAYER M3 ;
        RECT 34.144 21.824 34.176 21.856 ;
  LAYER M1 ;
        RECT 34.208 21.804 34.24 24.312 ;
  LAYER M3 ;
        RECT 34.208 24.26 34.24 24.292 ;
  LAYER M1 ;
        RECT 34.272 21.804 34.304 24.312 ;
  LAYER M3 ;
        RECT 34.272 21.824 34.304 21.856 ;
  LAYER M1 ;
        RECT 34.336 21.804 34.368 24.312 ;
  LAYER M3 ;
        RECT 34.336 24.26 34.368 24.292 ;
  LAYER M1 ;
        RECT 34.4 21.804 34.432 24.312 ;
  LAYER M3 ;
        RECT 34.4 21.824 34.432 21.856 ;
  LAYER M1 ;
        RECT 34.464 21.804 34.496 24.312 ;
  LAYER M3 ;
        RECT 34.464 24.26 34.496 24.292 ;
  LAYER M1 ;
        RECT 34.528 21.804 34.56 24.312 ;
  LAYER M3 ;
        RECT 34.528 21.824 34.56 21.856 ;
  LAYER M1 ;
        RECT 34.592 21.804 34.624 24.312 ;
  LAYER M3 ;
        RECT 34.592 24.26 34.624 24.292 ;
  LAYER M1 ;
        RECT 34.656 21.804 34.688 24.312 ;
  LAYER M3 ;
        RECT 34.656 21.824 34.688 21.856 ;
  LAYER M1 ;
        RECT 34.72 21.804 34.752 24.312 ;
  LAYER M3 ;
        RECT 34.72 24.26 34.752 24.292 ;
  LAYER M1 ;
        RECT 34.784 21.804 34.816 24.312 ;
  LAYER M3 ;
        RECT 34.784 21.824 34.816 21.856 ;
  LAYER M1 ;
        RECT 34.848 21.804 34.88 24.312 ;
  LAYER M3 ;
        RECT 34.848 24.26 34.88 24.292 ;
  LAYER M1 ;
        RECT 34.912 21.804 34.944 24.312 ;
  LAYER M3 ;
        RECT 34.912 21.824 34.944 21.856 ;
  LAYER M1 ;
        RECT 34.976 21.804 35.008 24.312 ;
  LAYER M3 ;
        RECT 32.608 24.196 32.64 24.228 ;
  LAYER M2 ;
        RECT 34.976 24.132 35.008 24.164 ;
  LAYER M2 ;
        RECT 32.608 24.068 32.64 24.1 ;
  LAYER M2 ;
        RECT 34.976 24.004 35.008 24.036 ;
  LAYER M2 ;
        RECT 32.608 23.94 32.64 23.972 ;
  LAYER M2 ;
        RECT 34.976 23.876 35.008 23.908 ;
  LAYER M2 ;
        RECT 32.608 23.812 32.64 23.844 ;
  LAYER M2 ;
        RECT 34.976 23.748 35.008 23.78 ;
  LAYER M2 ;
        RECT 32.608 23.684 32.64 23.716 ;
  LAYER M2 ;
        RECT 34.976 23.62 35.008 23.652 ;
  LAYER M2 ;
        RECT 32.608 23.556 32.64 23.588 ;
  LAYER M2 ;
        RECT 34.976 23.492 35.008 23.524 ;
  LAYER M2 ;
        RECT 32.608 23.428 32.64 23.46 ;
  LAYER M2 ;
        RECT 34.976 23.364 35.008 23.396 ;
  LAYER M2 ;
        RECT 32.608 23.3 32.64 23.332 ;
  LAYER M2 ;
        RECT 34.976 23.236 35.008 23.268 ;
  LAYER M2 ;
        RECT 32.608 23.172 32.64 23.204 ;
  LAYER M2 ;
        RECT 34.976 23.108 35.008 23.14 ;
  LAYER M2 ;
        RECT 32.608 23.044 32.64 23.076 ;
  LAYER M2 ;
        RECT 34.976 22.98 35.008 23.012 ;
  LAYER M2 ;
        RECT 32.608 22.916 32.64 22.948 ;
  LAYER M2 ;
        RECT 34.976 22.852 35.008 22.884 ;
  LAYER M2 ;
        RECT 32.608 22.788 32.64 22.82 ;
  LAYER M2 ;
        RECT 34.976 22.724 35.008 22.756 ;
  LAYER M2 ;
        RECT 32.608 22.66 32.64 22.692 ;
  LAYER M2 ;
        RECT 34.976 22.596 35.008 22.628 ;
  LAYER M2 ;
        RECT 32.608 22.532 32.64 22.564 ;
  LAYER M2 ;
        RECT 34.976 22.468 35.008 22.5 ;
  LAYER M2 ;
        RECT 32.608 22.404 32.64 22.436 ;
  LAYER M2 ;
        RECT 34.976 22.34 35.008 22.372 ;
  LAYER M2 ;
        RECT 32.608 22.276 32.64 22.308 ;
  LAYER M2 ;
        RECT 34.976 22.212 35.008 22.244 ;
  LAYER M2 ;
        RECT 32.608 22.148 32.64 22.18 ;
  LAYER M2 ;
        RECT 34.976 22.084 35.008 22.116 ;
  LAYER M2 ;
        RECT 32.608 22.02 32.64 22.052 ;
  LAYER M2 ;
        RECT 34.976 21.956 35.008 21.988 ;
  LAYER M2 ;
        RECT 32.56 21.756 35.056 24.36 ;
  LAYER M1 ;
        RECT 32.608 18.696 32.64 21.204 ;
  LAYER M3 ;
        RECT 32.608 18.716 32.64 18.748 ;
  LAYER M1 ;
        RECT 32.672 18.696 32.704 21.204 ;
  LAYER M3 ;
        RECT 32.672 21.152 32.704 21.184 ;
  LAYER M1 ;
        RECT 32.736 18.696 32.768 21.204 ;
  LAYER M3 ;
        RECT 32.736 18.716 32.768 18.748 ;
  LAYER M1 ;
        RECT 32.8 18.696 32.832 21.204 ;
  LAYER M3 ;
        RECT 32.8 21.152 32.832 21.184 ;
  LAYER M1 ;
        RECT 32.864 18.696 32.896 21.204 ;
  LAYER M3 ;
        RECT 32.864 18.716 32.896 18.748 ;
  LAYER M1 ;
        RECT 32.928 18.696 32.96 21.204 ;
  LAYER M3 ;
        RECT 32.928 21.152 32.96 21.184 ;
  LAYER M1 ;
        RECT 32.992 18.696 33.024 21.204 ;
  LAYER M3 ;
        RECT 32.992 18.716 33.024 18.748 ;
  LAYER M1 ;
        RECT 33.056 18.696 33.088 21.204 ;
  LAYER M3 ;
        RECT 33.056 21.152 33.088 21.184 ;
  LAYER M1 ;
        RECT 33.12 18.696 33.152 21.204 ;
  LAYER M3 ;
        RECT 33.12 18.716 33.152 18.748 ;
  LAYER M1 ;
        RECT 33.184 18.696 33.216 21.204 ;
  LAYER M3 ;
        RECT 33.184 21.152 33.216 21.184 ;
  LAYER M1 ;
        RECT 33.248 18.696 33.28 21.204 ;
  LAYER M3 ;
        RECT 33.248 18.716 33.28 18.748 ;
  LAYER M1 ;
        RECT 33.312 18.696 33.344 21.204 ;
  LAYER M3 ;
        RECT 33.312 21.152 33.344 21.184 ;
  LAYER M1 ;
        RECT 33.376 18.696 33.408 21.204 ;
  LAYER M3 ;
        RECT 33.376 18.716 33.408 18.748 ;
  LAYER M1 ;
        RECT 33.44 18.696 33.472 21.204 ;
  LAYER M3 ;
        RECT 33.44 21.152 33.472 21.184 ;
  LAYER M1 ;
        RECT 33.504 18.696 33.536 21.204 ;
  LAYER M3 ;
        RECT 33.504 18.716 33.536 18.748 ;
  LAYER M1 ;
        RECT 33.568 18.696 33.6 21.204 ;
  LAYER M3 ;
        RECT 33.568 21.152 33.6 21.184 ;
  LAYER M1 ;
        RECT 33.632 18.696 33.664 21.204 ;
  LAYER M3 ;
        RECT 33.632 18.716 33.664 18.748 ;
  LAYER M1 ;
        RECT 33.696 18.696 33.728 21.204 ;
  LAYER M3 ;
        RECT 33.696 21.152 33.728 21.184 ;
  LAYER M1 ;
        RECT 33.76 18.696 33.792 21.204 ;
  LAYER M3 ;
        RECT 33.76 18.716 33.792 18.748 ;
  LAYER M1 ;
        RECT 33.824 18.696 33.856 21.204 ;
  LAYER M3 ;
        RECT 33.824 21.152 33.856 21.184 ;
  LAYER M1 ;
        RECT 33.888 18.696 33.92 21.204 ;
  LAYER M3 ;
        RECT 33.888 18.716 33.92 18.748 ;
  LAYER M1 ;
        RECT 33.952 18.696 33.984 21.204 ;
  LAYER M3 ;
        RECT 33.952 21.152 33.984 21.184 ;
  LAYER M1 ;
        RECT 34.016 18.696 34.048 21.204 ;
  LAYER M3 ;
        RECT 34.016 18.716 34.048 18.748 ;
  LAYER M1 ;
        RECT 34.08 18.696 34.112 21.204 ;
  LAYER M3 ;
        RECT 34.08 21.152 34.112 21.184 ;
  LAYER M1 ;
        RECT 34.144 18.696 34.176 21.204 ;
  LAYER M3 ;
        RECT 34.144 18.716 34.176 18.748 ;
  LAYER M1 ;
        RECT 34.208 18.696 34.24 21.204 ;
  LAYER M3 ;
        RECT 34.208 21.152 34.24 21.184 ;
  LAYER M1 ;
        RECT 34.272 18.696 34.304 21.204 ;
  LAYER M3 ;
        RECT 34.272 18.716 34.304 18.748 ;
  LAYER M1 ;
        RECT 34.336 18.696 34.368 21.204 ;
  LAYER M3 ;
        RECT 34.336 21.152 34.368 21.184 ;
  LAYER M1 ;
        RECT 34.4 18.696 34.432 21.204 ;
  LAYER M3 ;
        RECT 34.4 18.716 34.432 18.748 ;
  LAYER M1 ;
        RECT 34.464 18.696 34.496 21.204 ;
  LAYER M3 ;
        RECT 34.464 21.152 34.496 21.184 ;
  LAYER M1 ;
        RECT 34.528 18.696 34.56 21.204 ;
  LAYER M3 ;
        RECT 34.528 18.716 34.56 18.748 ;
  LAYER M1 ;
        RECT 34.592 18.696 34.624 21.204 ;
  LAYER M3 ;
        RECT 34.592 21.152 34.624 21.184 ;
  LAYER M1 ;
        RECT 34.656 18.696 34.688 21.204 ;
  LAYER M3 ;
        RECT 34.656 18.716 34.688 18.748 ;
  LAYER M1 ;
        RECT 34.72 18.696 34.752 21.204 ;
  LAYER M3 ;
        RECT 34.72 21.152 34.752 21.184 ;
  LAYER M1 ;
        RECT 34.784 18.696 34.816 21.204 ;
  LAYER M3 ;
        RECT 34.784 18.716 34.816 18.748 ;
  LAYER M1 ;
        RECT 34.848 18.696 34.88 21.204 ;
  LAYER M3 ;
        RECT 34.848 21.152 34.88 21.184 ;
  LAYER M1 ;
        RECT 34.912 18.696 34.944 21.204 ;
  LAYER M3 ;
        RECT 34.912 18.716 34.944 18.748 ;
  LAYER M1 ;
        RECT 34.976 18.696 35.008 21.204 ;
  LAYER M3 ;
        RECT 32.608 21.088 32.64 21.12 ;
  LAYER M2 ;
        RECT 34.976 21.024 35.008 21.056 ;
  LAYER M2 ;
        RECT 32.608 20.96 32.64 20.992 ;
  LAYER M2 ;
        RECT 34.976 20.896 35.008 20.928 ;
  LAYER M2 ;
        RECT 32.608 20.832 32.64 20.864 ;
  LAYER M2 ;
        RECT 34.976 20.768 35.008 20.8 ;
  LAYER M2 ;
        RECT 32.608 20.704 32.64 20.736 ;
  LAYER M2 ;
        RECT 34.976 20.64 35.008 20.672 ;
  LAYER M2 ;
        RECT 32.608 20.576 32.64 20.608 ;
  LAYER M2 ;
        RECT 34.976 20.512 35.008 20.544 ;
  LAYER M2 ;
        RECT 32.608 20.448 32.64 20.48 ;
  LAYER M2 ;
        RECT 34.976 20.384 35.008 20.416 ;
  LAYER M2 ;
        RECT 32.608 20.32 32.64 20.352 ;
  LAYER M2 ;
        RECT 34.976 20.256 35.008 20.288 ;
  LAYER M2 ;
        RECT 32.608 20.192 32.64 20.224 ;
  LAYER M2 ;
        RECT 34.976 20.128 35.008 20.16 ;
  LAYER M2 ;
        RECT 32.608 20.064 32.64 20.096 ;
  LAYER M2 ;
        RECT 34.976 20 35.008 20.032 ;
  LAYER M2 ;
        RECT 32.608 19.936 32.64 19.968 ;
  LAYER M2 ;
        RECT 34.976 19.872 35.008 19.904 ;
  LAYER M2 ;
        RECT 32.608 19.808 32.64 19.84 ;
  LAYER M2 ;
        RECT 34.976 19.744 35.008 19.776 ;
  LAYER M2 ;
        RECT 32.608 19.68 32.64 19.712 ;
  LAYER M2 ;
        RECT 34.976 19.616 35.008 19.648 ;
  LAYER M2 ;
        RECT 32.608 19.552 32.64 19.584 ;
  LAYER M2 ;
        RECT 34.976 19.488 35.008 19.52 ;
  LAYER M2 ;
        RECT 32.608 19.424 32.64 19.456 ;
  LAYER M2 ;
        RECT 34.976 19.36 35.008 19.392 ;
  LAYER M2 ;
        RECT 32.608 19.296 32.64 19.328 ;
  LAYER M2 ;
        RECT 34.976 19.232 35.008 19.264 ;
  LAYER M2 ;
        RECT 32.608 19.168 32.64 19.2 ;
  LAYER M2 ;
        RECT 34.976 19.104 35.008 19.136 ;
  LAYER M2 ;
        RECT 32.608 19.04 32.64 19.072 ;
  LAYER M2 ;
        RECT 34.976 18.976 35.008 19.008 ;
  LAYER M2 ;
        RECT 32.608 18.912 32.64 18.944 ;
  LAYER M2 ;
        RECT 34.976 18.848 35.008 18.88 ;
  LAYER M2 ;
        RECT 32.56 18.648 35.056 21.252 ;
  LAYER M1 ;
        RECT 32.608 15.588 32.64 18.096 ;
  LAYER M3 ;
        RECT 32.608 15.608 32.64 15.64 ;
  LAYER M1 ;
        RECT 32.672 15.588 32.704 18.096 ;
  LAYER M3 ;
        RECT 32.672 18.044 32.704 18.076 ;
  LAYER M1 ;
        RECT 32.736 15.588 32.768 18.096 ;
  LAYER M3 ;
        RECT 32.736 15.608 32.768 15.64 ;
  LAYER M1 ;
        RECT 32.8 15.588 32.832 18.096 ;
  LAYER M3 ;
        RECT 32.8 18.044 32.832 18.076 ;
  LAYER M1 ;
        RECT 32.864 15.588 32.896 18.096 ;
  LAYER M3 ;
        RECT 32.864 15.608 32.896 15.64 ;
  LAYER M1 ;
        RECT 32.928 15.588 32.96 18.096 ;
  LAYER M3 ;
        RECT 32.928 18.044 32.96 18.076 ;
  LAYER M1 ;
        RECT 32.992 15.588 33.024 18.096 ;
  LAYER M3 ;
        RECT 32.992 15.608 33.024 15.64 ;
  LAYER M1 ;
        RECT 33.056 15.588 33.088 18.096 ;
  LAYER M3 ;
        RECT 33.056 18.044 33.088 18.076 ;
  LAYER M1 ;
        RECT 33.12 15.588 33.152 18.096 ;
  LAYER M3 ;
        RECT 33.12 15.608 33.152 15.64 ;
  LAYER M1 ;
        RECT 33.184 15.588 33.216 18.096 ;
  LAYER M3 ;
        RECT 33.184 18.044 33.216 18.076 ;
  LAYER M1 ;
        RECT 33.248 15.588 33.28 18.096 ;
  LAYER M3 ;
        RECT 33.248 15.608 33.28 15.64 ;
  LAYER M1 ;
        RECT 33.312 15.588 33.344 18.096 ;
  LAYER M3 ;
        RECT 33.312 18.044 33.344 18.076 ;
  LAYER M1 ;
        RECT 33.376 15.588 33.408 18.096 ;
  LAYER M3 ;
        RECT 33.376 15.608 33.408 15.64 ;
  LAYER M1 ;
        RECT 33.44 15.588 33.472 18.096 ;
  LAYER M3 ;
        RECT 33.44 18.044 33.472 18.076 ;
  LAYER M1 ;
        RECT 33.504 15.588 33.536 18.096 ;
  LAYER M3 ;
        RECT 33.504 15.608 33.536 15.64 ;
  LAYER M1 ;
        RECT 33.568 15.588 33.6 18.096 ;
  LAYER M3 ;
        RECT 33.568 18.044 33.6 18.076 ;
  LAYER M1 ;
        RECT 33.632 15.588 33.664 18.096 ;
  LAYER M3 ;
        RECT 33.632 15.608 33.664 15.64 ;
  LAYER M1 ;
        RECT 33.696 15.588 33.728 18.096 ;
  LAYER M3 ;
        RECT 33.696 18.044 33.728 18.076 ;
  LAYER M1 ;
        RECT 33.76 15.588 33.792 18.096 ;
  LAYER M3 ;
        RECT 33.76 15.608 33.792 15.64 ;
  LAYER M1 ;
        RECT 33.824 15.588 33.856 18.096 ;
  LAYER M3 ;
        RECT 33.824 18.044 33.856 18.076 ;
  LAYER M1 ;
        RECT 33.888 15.588 33.92 18.096 ;
  LAYER M3 ;
        RECT 33.888 15.608 33.92 15.64 ;
  LAYER M1 ;
        RECT 33.952 15.588 33.984 18.096 ;
  LAYER M3 ;
        RECT 33.952 18.044 33.984 18.076 ;
  LAYER M1 ;
        RECT 34.016 15.588 34.048 18.096 ;
  LAYER M3 ;
        RECT 34.016 15.608 34.048 15.64 ;
  LAYER M1 ;
        RECT 34.08 15.588 34.112 18.096 ;
  LAYER M3 ;
        RECT 34.08 18.044 34.112 18.076 ;
  LAYER M1 ;
        RECT 34.144 15.588 34.176 18.096 ;
  LAYER M3 ;
        RECT 34.144 15.608 34.176 15.64 ;
  LAYER M1 ;
        RECT 34.208 15.588 34.24 18.096 ;
  LAYER M3 ;
        RECT 34.208 18.044 34.24 18.076 ;
  LAYER M1 ;
        RECT 34.272 15.588 34.304 18.096 ;
  LAYER M3 ;
        RECT 34.272 15.608 34.304 15.64 ;
  LAYER M1 ;
        RECT 34.336 15.588 34.368 18.096 ;
  LAYER M3 ;
        RECT 34.336 18.044 34.368 18.076 ;
  LAYER M1 ;
        RECT 34.4 15.588 34.432 18.096 ;
  LAYER M3 ;
        RECT 34.4 15.608 34.432 15.64 ;
  LAYER M1 ;
        RECT 34.464 15.588 34.496 18.096 ;
  LAYER M3 ;
        RECT 34.464 18.044 34.496 18.076 ;
  LAYER M1 ;
        RECT 34.528 15.588 34.56 18.096 ;
  LAYER M3 ;
        RECT 34.528 15.608 34.56 15.64 ;
  LAYER M1 ;
        RECT 34.592 15.588 34.624 18.096 ;
  LAYER M3 ;
        RECT 34.592 18.044 34.624 18.076 ;
  LAYER M1 ;
        RECT 34.656 15.588 34.688 18.096 ;
  LAYER M3 ;
        RECT 34.656 15.608 34.688 15.64 ;
  LAYER M1 ;
        RECT 34.72 15.588 34.752 18.096 ;
  LAYER M3 ;
        RECT 34.72 18.044 34.752 18.076 ;
  LAYER M1 ;
        RECT 34.784 15.588 34.816 18.096 ;
  LAYER M3 ;
        RECT 34.784 15.608 34.816 15.64 ;
  LAYER M1 ;
        RECT 34.848 15.588 34.88 18.096 ;
  LAYER M3 ;
        RECT 34.848 18.044 34.88 18.076 ;
  LAYER M1 ;
        RECT 34.912 15.588 34.944 18.096 ;
  LAYER M3 ;
        RECT 34.912 15.608 34.944 15.64 ;
  LAYER M1 ;
        RECT 34.976 15.588 35.008 18.096 ;
  LAYER M3 ;
        RECT 32.608 17.98 32.64 18.012 ;
  LAYER M2 ;
        RECT 34.976 17.916 35.008 17.948 ;
  LAYER M2 ;
        RECT 32.608 17.852 32.64 17.884 ;
  LAYER M2 ;
        RECT 34.976 17.788 35.008 17.82 ;
  LAYER M2 ;
        RECT 32.608 17.724 32.64 17.756 ;
  LAYER M2 ;
        RECT 34.976 17.66 35.008 17.692 ;
  LAYER M2 ;
        RECT 32.608 17.596 32.64 17.628 ;
  LAYER M2 ;
        RECT 34.976 17.532 35.008 17.564 ;
  LAYER M2 ;
        RECT 32.608 17.468 32.64 17.5 ;
  LAYER M2 ;
        RECT 34.976 17.404 35.008 17.436 ;
  LAYER M2 ;
        RECT 32.608 17.34 32.64 17.372 ;
  LAYER M2 ;
        RECT 34.976 17.276 35.008 17.308 ;
  LAYER M2 ;
        RECT 32.608 17.212 32.64 17.244 ;
  LAYER M2 ;
        RECT 34.976 17.148 35.008 17.18 ;
  LAYER M2 ;
        RECT 32.608 17.084 32.64 17.116 ;
  LAYER M2 ;
        RECT 34.976 17.02 35.008 17.052 ;
  LAYER M2 ;
        RECT 32.608 16.956 32.64 16.988 ;
  LAYER M2 ;
        RECT 34.976 16.892 35.008 16.924 ;
  LAYER M2 ;
        RECT 32.608 16.828 32.64 16.86 ;
  LAYER M2 ;
        RECT 34.976 16.764 35.008 16.796 ;
  LAYER M2 ;
        RECT 32.608 16.7 32.64 16.732 ;
  LAYER M2 ;
        RECT 34.976 16.636 35.008 16.668 ;
  LAYER M2 ;
        RECT 32.608 16.572 32.64 16.604 ;
  LAYER M2 ;
        RECT 34.976 16.508 35.008 16.54 ;
  LAYER M2 ;
        RECT 32.608 16.444 32.64 16.476 ;
  LAYER M2 ;
        RECT 34.976 16.38 35.008 16.412 ;
  LAYER M2 ;
        RECT 32.608 16.316 32.64 16.348 ;
  LAYER M2 ;
        RECT 34.976 16.252 35.008 16.284 ;
  LAYER M2 ;
        RECT 32.608 16.188 32.64 16.22 ;
  LAYER M2 ;
        RECT 34.976 16.124 35.008 16.156 ;
  LAYER M2 ;
        RECT 32.608 16.06 32.64 16.092 ;
  LAYER M2 ;
        RECT 34.976 15.996 35.008 16.028 ;
  LAYER M2 ;
        RECT 32.608 15.932 32.64 15.964 ;
  LAYER M2 ;
        RECT 34.976 15.868 35.008 15.9 ;
  LAYER M2 ;
        RECT 32.608 15.804 32.64 15.836 ;
  LAYER M2 ;
        RECT 34.976 15.74 35.008 15.772 ;
  LAYER M2 ;
        RECT 32.56 15.54 35.056 18.144 ;
  LAYER M1 ;
        RECT 35.584 28.02 35.616 30.528 ;
  LAYER M3 ;
        RECT 35.584 28.04 35.616 28.072 ;
  LAYER M1 ;
        RECT 35.648 28.02 35.68 30.528 ;
  LAYER M3 ;
        RECT 35.648 30.476 35.68 30.508 ;
  LAYER M1 ;
        RECT 35.712 28.02 35.744 30.528 ;
  LAYER M3 ;
        RECT 35.712 28.04 35.744 28.072 ;
  LAYER M1 ;
        RECT 35.776 28.02 35.808 30.528 ;
  LAYER M3 ;
        RECT 35.776 30.476 35.808 30.508 ;
  LAYER M1 ;
        RECT 35.84 28.02 35.872 30.528 ;
  LAYER M3 ;
        RECT 35.84 28.04 35.872 28.072 ;
  LAYER M1 ;
        RECT 35.904 28.02 35.936 30.528 ;
  LAYER M3 ;
        RECT 35.904 30.476 35.936 30.508 ;
  LAYER M1 ;
        RECT 35.968 28.02 36 30.528 ;
  LAYER M3 ;
        RECT 35.968 28.04 36 28.072 ;
  LAYER M1 ;
        RECT 36.032 28.02 36.064 30.528 ;
  LAYER M3 ;
        RECT 36.032 30.476 36.064 30.508 ;
  LAYER M1 ;
        RECT 36.096 28.02 36.128 30.528 ;
  LAYER M3 ;
        RECT 36.096 28.04 36.128 28.072 ;
  LAYER M1 ;
        RECT 36.16 28.02 36.192 30.528 ;
  LAYER M3 ;
        RECT 36.16 30.476 36.192 30.508 ;
  LAYER M1 ;
        RECT 36.224 28.02 36.256 30.528 ;
  LAYER M3 ;
        RECT 36.224 28.04 36.256 28.072 ;
  LAYER M1 ;
        RECT 36.288 28.02 36.32 30.528 ;
  LAYER M3 ;
        RECT 36.288 30.476 36.32 30.508 ;
  LAYER M1 ;
        RECT 36.352 28.02 36.384 30.528 ;
  LAYER M3 ;
        RECT 36.352 28.04 36.384 28.072 ;
  LAYER M1 ;
        RECT 36.416 28.02 36.448 30.528 ;
  LAYER M3 ;
        RECT 36.416 30.476 36.448 30.508 ;
  LAYER M1 ;
        RECT 36.48 28.02 36.512 30.528 ;
  LAYER M3 ;
        RECT 36.48 28.04 36.512 28.072 ;
  LAYER M1 ;
        RECT 36.544 28.02 36.576 30.528 ;
  LAYER M3 ;
        RECT 36.544 30.476 36.576 30.508 ;
  LAYER M1 ;
        RECT 36.608 28.02 36.64 30.528 ;
  LAYER M3 ;
        RECT 36.608 28.04 36.64 28.072 ;
  LAYER M1 ;
        RECT 36.672 28.02 36.704 30.528 ;
  LAYER M3 ;
        RECT 36.672 30.476 36.704 30.508 ;
  LAYER M1 ;
        RECT 36.736 28.02 36.768 30.528 ;
  LAYER M3 ;
        RECT 36.736 28.04 36.768 28.072 ;
  LAYER M1 ;
        RECT 36.8 28.02 36.832 30.528 ;
  LAYER M3 ;
        RECT 36.8 30.476 36.832 30.508 ;
  LAYER M1 ;
        RECT 36.864 28.02 36.896 30.528 ;
  LAYER M3 ;
        RECT 36.864 28.04 36.896 28.072 ;
  LAYER M1 ;
        RECT 36.928 28.02 36.96 30.528 ;
  LAYER M3 ;
        RECT 36.928 30.476 36.96 30.508 ;
  LAYER M1 ;
        RECT 36.992 28.02 37.024 30.528 ;
  LAYER M3 ;
        RECT 36.992 28.04 37.024 28.072 ;
  LAYER M1 ;
        RECT 37.056 28.02 37.088 30.528 ;
  LAYER M3 ;
        RECT 37.056 30.476 37.088 30.508 ;
  LAYER M1 ;
        RECT 37.12 28.02 37.152 30.528 ;
  LAYER M3 ;
        RECT 37.12 28.04 37.152 28.072 ;
  LAYER M1 ;
        RECT 37.184 28.02 37.216 30.528 ;
  LAYER M3 ;
        RECT 37.184 30.476 37.216 30.508 ;
  LAYER M1 ;
        RECT 37.248 28.02 37.28 30.528 ;
  LAYER M3 ;
        RECT 37.248 28.04 37.28 28.072 ;
  LAYER M1 ;
        RECT 37.312 28.02 37.344 30.528 ;
  LAYER M3 ;
        RECT 37.312 30.476 37.344 30.508 ;
  LAYER M1 ;
        RECT 37.376 28.02 37.408 30.528 ;
  LAYER M3 ;
        RECT 37.376 28.04 37.408 28.072 ;
  LAYER M1 ;
        RECT 37.44 28.02 37.472 30.528 ;
  LAYER M3 ;
        RECT 37.44 30.476 37.472 30.508 ;
  LAYER M1 ;
        RECT 37.504 28.02 37.536 30.528 ;
  LAYER M3 ;
        RECT 37.504 28.04 37.536 28.072 ;
  LAYER M1 ;
        RECT 37.568 28.02 37.6 30.528 ;
  LAYER M3 ;
        RECT 37.568 30.476 37.6 30.508 ;
  LAYER M1 ;
        RECT 37.632 28.02 37.664 30.528 ;
  LAYER M3 ;
        RECT 37.632 28.04 37.664 28.072 ;
  LAYER M1 ;
        RECT 37.696 28.02 37.728 30.528 ;
  LAYER M3 ;
        RECT 37.696 30.476 37.728 30.508 ;
  LAYER M1 ;
        RECT 37.76 28.02 37.792 30.528 ;
  LAYER M3 ;
        RECT 37.76 28.04 37.792 28.072 ;
  LAYER M1 ;
        RECT 37.824 28.02 37.856 30.528 ;
  LAYER M3 ;
        RECT 37.824 30.476 37.856 30.508 ;
  LAYER M1 ;
        RECT 37.888 28.02 37.92 30.528 ;
  LAYER M3 ;
        RECT 37.888 28.04 37.92 28.072 ;
  LAYER M1 ;
        RECT 37.952 28.02 37.984 30.528 ;
  LAYER M3 ;
        RECT 35.584 30.412 35.616 30.444 ;
  LAYER M2 ;
        RECT 37.952 30.348 37.984 30.38 ;
  LAYER M2 ;
        RECT 35.584 30.284 35.616 30.316 ;
  LAYER M2 ;
        RECT 37.952 30.22 37.984 30.252 ;
  LAYER M2 ;
        RECT 35.584 30.156 35.616 30.188 ;
  LAYER M2 ;
        RECT 37.952 30.092 37.984 30.124 ;
  LAYER M2 ;
        RECT 35.584 30.028 35.616 30.06 ;
  LAYER M2 ;
        RECT 37.952 29.964 37.984 29.996 ;
  LAYER M2 ;
        RECT 35.584 29.9 35.616 29.932 ;
  LAYER M2 ;
        RECT 37.952 29.836 37.984 29.868 ;
  LAYER M2 ;
        RECT 35.584 29.772 35.616 29.804 ;
  LAYER M2 ;
        RECT 37.952 29.708 37.984 29.74 ;
  LAYER M2 ;
        RECT 35.584 29.644 35.616 29.676 ;
  LAYER M2 ;
        RECT 37.952 29.58 37.984 29.612 ;
  LAYER M2 ;
        RECT 35.584 29.516 35.616 29.548 ;
  LAYER M2 ;
        RECT 37.952 29.452 37.984 29.484 ;
  LAYER M2 ;
        RECT 35.584 29.388 35.616 29.42 ;
  LAYER M2 ;
        RECT 37.952 29.324 37.984 29.356 ;
  LAYER M2 ;
        RECT 35.584 29.26 35.616 29.292 ;
  LAYER M2 ;
        RECT 37.952 29.196 37.984 29.228 ;
  LAYER M2 ;
        RECT 35.584 29.132 35.616 29.164 ;
  LAYER M2 ;
        RECT 37.952 29.068 37.984 29.1 ;
  LAYER M2 ;
        RECT 35.584 29.004 35.616 29.036 ;
  LAYER M2 ;
        RECT 37.952 28.94 37.984 28.972 ;
  LAYER M2 ;
        RECT 35.584 28.876 35.616 28.908 ;
  LAYER M2 ;
        RECT 37.952 28.812 37.984 28.844 ;
  LAYER M2 ;
        RECT 35.584 28.748 35.616 28.78 ;
  LAYER M2 ;
        RECT 37.952 28.684 37.984 28.716 ;
  LAYER M2 ;
        RECT 35.584 28.62 35.616 28.652 ;
  LAYER M2 ;
        RECT 37.952 28.556 37.984 28.588 ;
  LAYER M2 ;
        RECT 35.584 28.492 35.616 28.524 ;
  LAYER M2 ;
        RECT 37.952 28.428 37.984 28.46 ;
  LAYER M2 ;
        RECT 35.584 28.364 35.616 28.396 ;
  LAYER M2 ;
        RECT 37.952 28.3 37.984 28.332 ;
  LAYER M2 ;
        RECT 35.584 28.236 35.616 28.268 ;
  LAYER M2 ;
        RECT 37.952 28.172 37.984 28.204 ;
  LAYER M2 ;
        RECT 35.536 27.972 38.032 30.576 ;
  LAYER M1 ;
        RECT 35.584 24.912 35.616 27.42 ;
  LAYER M3 ;
        RECT 35.584 24.932 35.616 24.964 ;
  LAYER M1 ;
        RECT 35.648 24.912 35.68 27.42 ;
  LAYER M3 ;
        RECT 35.648 27.368 35.68 27.4 ;
  LAYER M1 ;
        RECT 35.712 24.912 35.744 27.42 ;
  LAYER M3 ;
        RECT 35.712 24.932 35.744 24.964 ;
  LAYER M1 ;
        RECT 35.776 24.912 35.808 27.42 ;
  LAYER M3 ;
        RECT 35.776 27.368 35.808 27.4 ;
  LAYER M1 ;
        RECT 35.84 24.912 35.872 27.42 ;
  LAYER M3 ;
        RECT 35.84 24.932 35.872 24.964 ;
  LAYER M1 ;
        RECT 35.904 24.912 35.936 27.42 ;
  LAYER M3 ;
        RECT 35.904 27.368 35.936 27.4 ;
  LAYER M1 ;
        RECT 35.968 24.912 36 27.42 ;
  LAYER M3 ;
        RECT 35.968 24.932 36 24.964 ;
  LAYER M1 ;
        RECT 36.032 24.912 36.064 27.42 ;
  LAYER M3 ;
        RECT 36.032 27.368 36.064 27.4 ;
  LAYER M1 ;
        RECT 36.096 24.912 36.128 27.42 ;
  LAYER M3 ;
        RECT 36.096 24.932 36.128 24.964 ;
  LAYER M1 ;
        RECT 36.16 24.912 36.192 27.42 ;
  LAYER M3 ;
        RECT 36.16 27.368 36.192 27.4 ;
  LAYER M1 ;
        RECT 36.224 24.912 36.256 27.42 ;
  LAYER M3 ;
        RECT 36.224 24.932 36.256 24.964 ;
  LAYER M1 ;
        RECT 36.288 24.912 36.32 27.42 ;
  LAYER M3 ;
        RECT 36.288 27.368 36.32 27.4 ;
  LAYER M1 ;
        RECT 36.352 24.912 36.384 27.42 ;
  LAYER M3 ;
        RECT 36.352 24.932 36.384 24.964 ;
  LAYER M1 ;
        RECT 36.416 24.912 36.448 27.42 ;
  LAYER M3 ;
        RECT 36.416 27.368 36.448 27.4 ;
  LAYER M1 ;
        RECT 36.48 24.912 36.512 27.42 ;
  LAYER M3 ;
        RECT 36.48 24.932 36.512 24.964 ;
  LAYER M1 ;
        RECT 36.544 24.912 36.576 27.42 ;
  LAYER M3 ;
        RECT 36.544 27.368 36.576 27.4 ;
  LAYER M1 ;
        RECT 36.608 24.912 36.64 27.42 ;
  LAYER M3 ;
        RECT 36.608 24.932 36.64 24.964 ;
  LAYER M1 ;
        RECT 36.672 24.912 36.704 27.42 ;
  LAYER M3 ;
        RECT 36.672 27.368 36.704 27.4 ;
  LAYER M1 ;
        RECT 36.736 24.912 36.768 27.42 ;
  LAYER M3 ;
        RECT 36.736 24.932 36.768 24.964 ;
  LAYER M1 ;
        RECT 36.8 24.912 36.832 27.42 ;
  LAYER M3 ;
        RECT 36.8 27.368 36.832 27.4 ;
  LAYER M1 ;
        RECT 36.864 24.912 36.896 27.42 ;
  LAYER M3 ;
        RECT 36.864 24.932 36.896 24.964 ;
  LAYER M1 ;
        RECT 36.928 24.912 36.96 27.42 ;
  LAYER M3 ;
        RECT 36.928 27.368 36.96 27.4 ;
  LAYER M1 ;
        RECT 36.992 24.912 37.024 27.42 ;
  LAYER M3 ;
        RECT 36.992 24.932 37.024 24.964 ;
  LAYER M1 ;
        RECT 37.056 24.912 37.088 27.42 ;
  LAYER M3 ;
        RECT 37.056 27.368 37.088 27.4 ;
  LAYER M1 ;
        RECT 37.12 24.912 37.152 27.42 ;
  LAYER M3 ;
        RECT 37.12 24.932 37.152 24.964 ;
  LAYER M1 ;
        RECT 37.184 24.912 37.216 27.42 ;
  LAYER M3 ;
        RECT 37.184 27.368 37.216 27.4 ;
  LAYER M1 ;
        RECT 37.248 24.912 37.28 27.42 ;
  LAYER M3 ;
        RECT 37.248 24.932 37.28 24.964 ;
  LAYER M1 ;
        RECT 37.312 24.912 37.344 27.42 ;
  LAYER M3 ;
        RECT 37.312 27.368 37.344 27.4 ;
  LAYER M1 ;
        RECT 37.376 24.912 37.408 27.42 ;
  LAYER M3 ;
        RECT 37.376 24.932 37.408 24.964 ;
  LAYER M1 ;
        RECT 37.44 24.912 37.472 27.42 ;
  LAYER M3 ;
        RECT 37.44 27.368 37.472 27.4 ;
  LAYER M1 ;
        RECT 37.504 24.912 37.536 27.42 ;
  LAYER M3 ;
        RECT 37.504 24.932 37.536 24.964 ;
  LAYER M1 ;
        RECT 37.568 24.912 37.6 27.42 ;
  LAYER M3 ;
        RECT 37.568 27.368 37.6 27.4 ;
  LAYER M1 ;
        RECT 37.632 24.912 37.664 27.42 ;
  LAYER M3 ;
        RECT 37.632 24.932 37.664 24.964 ;
  LAYER M1 ;
        RECT 37.696 24.912 37.728 27.42 ;
  LAYER M3 ;
        RECT 37.696 27.368 37.728 27.4 ;
  LAYER M1 ;
        RECT 37.76 24.912 37.792 27.42 ;
  LAYER M3 ;
        RECT 37.76 24.932 37.792 24.964 ;
  LAYER M1 ;
        RECT 37.824 24.912 37.856 27.42 ;
  LAYER M3 ;
        RECT 37.824 27.368 37.856 27.4 ;
  LAYER M1 ;
        RECT 37.888 24.912 37.92 27.42 ;
  LAYER M3 ;
        RECT 37.888 24.932 37.92 24.964 ;
  LAYER M1 ;
        RECT 37.952 24.912 37.984 27.42 ;
  LAYER M3 ;
        RECT 35.584 27.304 35.616 27.336 ;
  LAYER M2 ;
        RECT 37.952 27.24 37.984 27.272 ;
  LAYER M2 ;
        RECT 35.584 27.176 35.616 27.208 ;
  LAYER M2 ;
        RECT 37.952 27.112 37.984 27.144 ;
  LAYER M2 ;
        RECT 35.584 27.048 35.616 27.08 ;
  LAYER M2 ;
        RECT 37.952 26.984 37.984 27.016 ;
  LAYER M2 ;
        RECT 35.584 26.92 35.616 26.952 ;
  LAYER M2 ;
        RECT 37.952 26.856 37.984 26.888 ;
  LAYER M2 ;
        RECT 35.584 26.792 35.616 26.824 ;
  LAYER M2 ;
        RECT 37.952 26.728 37.984 26.76 ;
  LAYER M2 ;
        RECT 35.584 26.664 35.616 26.696 ;
  LAYER M2 ;
        RECT 37.952 26.6 37.984 26.632 ;
  LAYER M2 ;
        RECT 35.584 26.536 35.616 26.568 ;
  LAYER M2 ;
        RECT 37.952 26.472 37.984 26.504 ;
  LAYER M2 ;
        RECT 35.584 26.408 35.616 26.44 ;
  LAYER M2 ;
        RECT 37.952 26.344 37.984 26.376 ;
  LAYER M2 ;
        RECT 35.584 26.28 35.616 26.312 ;
  LAYER M2 ;
        RECT 37.952 26.216 37.984 26.248 ;
  LAYER M2 ;
        RECT 35.584 26.152 35.616 26.184 ;
  LAYER M2 ;
        RECT 37.952 26.088 37.984 26.12 ;
  LAYER M2 ;
        RECT 35.584 26.024 35.616 26.056 ;
  LAYER M2 ;
        RECT 37.952 25.96 37.984 25.992 ;
  LAYER M2 ;
        RECT 35.584 25.896 35.616 25.928 ;
  LAYER M2 ;
        RECT 37.952 25.832 37.984 25.864 ;
  LAYER M2 ;
        RECT 35.584 25.768 35.616 25.8 ;
  LAYER M2 ;
        RECT 37.952 25.704 37.984 25.736 ;
  LAYER M2 ;
        RECT 35.584 25.64 35.616 25.672 ;
  LAYER M2 ;
        RECT 37.952 25.576 37.984 25.608 ;
  LAYER M2 ;
        RECT 35.584 25.512 35.616 25.544 ;
  LAYER M2 ;
        RECT 37.952 25.448 37.984 25.48 ;
  LAYER M2 ;
        RECT 35.584 25.384 35.616 25.416 ;
  LAYER M2 ;
        RECT 37.952 25.32 37.984 25.352 ;
  LAYER M2 ;
        RECT 35.584 25.256 35.616 25.288 ;
  LAYER M2 ;
        RECT 37.952 25.192 37.984 25.224 ;
  LAYER M2 ;
        RECT 35.584 25.128 35.616 25.16 ;
  LAYER M2 ;
        RECT 37.952 25.064 37.984 25.096 ;
  LAYER M2 ;
        RECT 35.536 24.864 38.032 27.468 ;
  LAYER M1 ;
        RECT 35.584 21.804 35.616 24.312 ;
  LAYER M3 ;
        RECT 35.584 21.824 35.616 21.856 ;
  LAYER M1 ;
        RECT 35.648 21.804 35.68 24.312 ;
  LAYER M3 ;
        RECT 35.648 24.26 35.68 24.292 ;
  LAYER M1 ;
        RECT 35.712 21.804 35.744 24.312 ;
  LAYER M3 ;
        RECT 35.712 21.824 35.744 21.856 ;
  LAYER M1 ;
        RECT 35.776 21.804 35.808 24.312 ;
  LAYER M3 ;
        RECT 35.776 24.26 35.808 24.292 ;
  LAYER M1 ;
        RECT 35.84 21.804 35.872 24.312 ;
  LAYER M3 ;
        RECT 35.84 21.824 35.872 21.856 ;
  LAYER M1 ;
        RECT 35.904 21.804 35.936 24.312 ;
  LAYER M3 ;
        RECT 35.904 24.26 35.936 24.292 ;
  LAYER M1 ;
        RECT 35.968 21.804 36 24.312 ;
  LAYER M3 ;
        RECT 35.968 21.824 36 21.856 ;
  LAYER M1 ;
        RECT 36.032 21.804 36.064 24.312 ;
  LAYER M3 ;
        RECT 36.032 24.26 36.064 24.292 ;
  LAYER M1 ;
        RECT 36.096 21.804 36.128 24.312 ;
  LAYER M3 ;
        RECT 36.096 21.824 36.128 21.856 ;
  LAYER M1 ;
        RECT 36.16 21.804 36.192 24.312 ;
  LAYER M3 ;
        RECT 36.16 24.26 36.192 24.292 ;
  LAYER M1 ;
        RECT 36.224 21.804 36.256 24.312 ;
  LAYER M3 ;
        RECT 36.224 21.824 36.256 21.856 ;
  LAYER M1 ;
        RECT 36.288 21.804 36.32 24.312 ;
  LAYER M3 ;
        RECT 36.288 24.26 36.32 24.292 ;
  LAYER M1 ;
        RECT 36.352 21.804 36.384 24.312 ;
  LAYER M3 ;
        RECT 36.352 21.824 36.384 21.856 ;
  LAYER M1 ;
        RECT 36.416 21.804 36.448 24.312 ;
  LAYER M3 ;
        RECT 36.416 24.26 36.448 24.292 ;
  LAYER M1 ;
        RECT 36.48 21.804 36.512 24.312 ;
  LAYER M3 ;
        RECT 36.48 21.824 36.512 21.856 ;
  LAYER M1 ;
        RECT 36.544 21.804 36.576 24.312 ;
  LAYER M3 ;
        RECT 36.544 24.26 36.576 24.292 ;
  LAYER M1 ;
        RECT 36.608 21.804 36.64 24.312 ;
  LAYER M3 ;
        RECT 36.608 21.824 36.64 21.856 ;
  LAYER M1 ;
        RECT 36.672 21.804 36.704 24.312 ;
  LAYER M3 ;
        RECT 36.672 24.26 36.704 24.292 ;
  LAYER M1 ;
        RECT 36.736 21.804 36.768 24.312 ;
  LAYER M3 ;
        RECT 36.736 21.824 36.768 21.856 ;
  LAYER M1 ;
        RECT 36.8 21.804 36.832 24.312 ;
  LAYER M3 ;
        RECT 36.8 24.26 36.832 24.292 ;
  LAYER M1 ;
        RECT 36.864 21.804 36.896 24.312 ;
  LAYER M3 ;
        RECT 36.864 21.824 36.896 21.856 ;
  LAYER M1 ;
        RECT 36.928 21.804 36.96 24.312 ;
  LAYER M3 ;
        RECT 36.928 24.26 36.96 24.292 ;
  LAYER M1 ;
        RECT 36.992 21.804 37.024 24.312 ;
  LAYER M3 ;
        RECT 36.992 21.824 37.024 21.856 ;
  LAYER M1 ;
        RECT 37.056 21.804 37.088 24.312 ;
  LAYER M3 ;
        RECT 37.056 24.26 37.088 24.292 ;
  LAYER M1 ;
        RECT 37.12 21.804 37.152 24.312 ;
  LAYER M3 ;
        RECT 37.12 21.824 37.152 21.856 ;
  LAYER M1 ;
        RECT 37.184 21.804 37.216 24.312 ;
  LAYER M3 ;
        RECT 37.184 24.26 37.216 24.292 ;
  LAYER M1 ;
        RECT 37.248 21.804 37.28 24.312 ;
  LAYER M3 ;
        RECT 37.248 21.824 37.28 21.856 ;
  LAYER M1 ;
        RECT 37.312 21.804 37.344 24.312 ;
  LAYER M3 ;
        RECT 37.312 24.26 37.344 24.292 ;
  LAYER M1 ;
        RECT 37.376 21.804 37.408 24.312 ;
  LAYER M3 ;
        RECT 37.376 21.824 37.408 21.856 ;
  LAYER M1 ;
        RECT 37.44 21.804 37.472 24.312 ;
  LAYER M3 ;
        RECT 37.44 24.26 37.472 24.292 ;
  LAYER M1 ;
        RECT 37.504 21.804 37.536 24.312 ;
  LAYER M3 ;
        RECT 37.504 21.824 37.536 21.856 ;
  LAYER M1 ;
        RECT 37.568 21.804 37.6 24.312 ;
  LAYER M3 ;
        RECT 37.568 24.26 37.6 24.292 ;
  LAYER M1 ;
        RECT 37.632 21.804 37.664 24.312 ;
  LAYER M3 ;
        RECT 37.632 21.824 37.664 21.856 ;
  LAYER M1 ;
        RECT 37.696 21.804 37.728 24.312 ;
  LAYER M3 ;
        RECT 37.696 24.26 37.728 24.292 ;
  LAYER M1 ;
        RECT 37.76 21.804 37.792 24.312 ;
  LAYER M3 ;
        RECT 37.76 21.824 37.792 21.856 ;
  LAYER M1 ;
        RECT 37.824 21.804 37.856 24.312 ;
  LAYER M3 ;
        RECT 37.824 24.26 37.856 24.292 ;
  LAYER M1 ;
        RECT 37.888 21.804 37.92 24.312 ;
  LAYER M3 ;
        RECT 37.888 21.824 37.92 21.856 ;
  LAYER M1 ;
        RECT 37.952 21.804 37.984 24.312 ;
  LAYER M3 ;
        RECT 35.584 24.196 35.616 24.228 ;
  LAYER M2 ;
        RECT 37.952 24.132 37.984 24.164 ;
  LAYER M2 ;
        RECT 35.584 24.068 35.616 24.1 ;
  LAYER M2 ;
        RECT 37.952 24.004 37.984 24.036 ;
  LAYER M2 ;
        RECT 35.584 23.94 35.616 23.972 ;
  LAYER M2 ;
        RECT 37.952 23.876 37.984 23.908 ;
  LAYER M2 ;
        RECT 35.584 23.812 35.616 23.844 ;
  LAYER M2 ;
        RECT 37.952 23.748 37.984 23.78 ;
  LAYER M2 ;
        RECT 35.584 23.684 35.616 23.716 ;
  LAYER M2 ;
        RECT 37.952 23.62 37.984 23.652 ;
  LAYER M2 ;
        RECT 35.584 23.556 35.616 23.588 ;
  LAYER M2 ;
        RECT 37.952 23.492 37.984 23.524 ;
  LAYER M2 ;
        RECT 35.584 23.428 35.616 23.46 ;
  LAYER M2 ;
        RECT 37.952 23.364 37.984 23.396 ;
  LAYER M2 ;
        RECT 35.584 23.3 35.616 23.332 ;
  LAYER M2 ;
        RECT 37.952 23.236 37.984 23.268 ;
  LAYER M2 ;
        RECT 35.584 23.172 35.616 23.204 ;
  LAYER M2 ;
        RECT 37.952 23.108 37.984 23.14 ;
  LAYER M2 ;
        RECT 35.584 23.044 35.616 23.076 ;
  LAYER M2 ;
        RECT 37.952 22.98 37.984 23.012 ;
  LAYER M2 ;
        RECT 35.584 22.916 35.616 22.948 ;
  LAYER M2 ;
        RECT 37.952 22.852 37.984 22.884 ;
  LAYER M2 ;
        RECT 35.584 22.788 35.616 22.82 ;
  LAYER M2 ;
        RECT 37.952 22.724 37.984 22.756 ;
  LAYER M2 ;
        RECT 35.584 22.66 35.616 22.692 ;
  LAYER M2 ;
        RECT 37.952 22.596 37.984 22.628 ;
  LAYER M2 ;
        RECT 35.584 22.532 35.616 22.564 ;
  LAYER M2 ;
        RECT 37.952 22.468 37.984 22.5 ;
  LAYER M2 ;
        RECT 35.584 22.404 35.616 22.436 ;
  LAYER M2 ;
        RECT 37.952 22.34 37.984 22.372 ;
  LAYER M2 ;
        RECT 35.584 22.276 35.616 22.308 ;
  LAYER M2 ;
        RECT 37.952 22.212 37.984 22.244 ;
  LAYER M2 ;
        RECT 35.584 22.148 35.616 22.18 ;
  LAYER M2 ;
        RECT 37.952 22.084 37.984 22.116 ;
  LAYER M2 ;
        RECT 35.584 22.02 35.616 22.052 ;
  LAYER M2 ;
        RECT 37.952 21.956 37.984 21.988 ;
  LAYER M2 ;
        RECT 35.536 21.756 38.032 24.36 ;
  LAYER M1 ;
        RECT 35.584 18.696 35.616 21.204 ;
  LAYER M3 ;
        RECT 35.584 18.716 35.616 18.748 ;
  LAYER M1 ;
        RECT 35.648 18.696 35.68 21.204 ;
  LAYER M3 ;
        RECT 35.648 21.152 35.68 21.184 ;
  LAYER M1 ;
        RECT 35.712 18.696 35.744 21.204 ;
  LAYER M3 ;
        RECT 35.712 18.716 35.744 18.748 ;
  LAYER M1 ;
        RECT 35.776 18.696 35.808 21.204 ;
  LAYER M3 ;
        RECT 35.776 21.152 35.808 21.184 ;
  LAYER M1 ;
        RECT 35.84 18.696 35.872 21.204 ;
  LAYER M3 ;
        RECT 35.84 18.716 35.872 18.748 ;
  LAYER M1 ;
        RECT 35.904 18.696 35.936 21.204 ;
  LAYER M3 ;
        RECT 35.904 21.152 35.936 21.184 ;
  LAYER M1 ;
        RECT 35.968 18.696 36 21.204 ;
  LAYER M3 ;
        RECT 35.968 18.716 36 18.748 ;
  LAYER M1 ;
        RECT 36.032 18.696 36.064 21.204 ;
  LAYER M3 ;
        RECT 36.032 21.152 36.064 21.184 ;
  LAYER M1 ;
        RECT 36.096 18.696 36.128 21.204 ;
  LAYER M3 ;
        RECT 36.096 18.716 36.128 18.748 ;
  LAYER M1 ;
        RECT 36.16 18.696 36.192 21.204 ;
  LAYER M3 ;
        RECT 36.16 21.152 36.192 21.184 ;
  LAYER M1 ;
        RECT 36.224 18.696 36.256 21.204 ;
  LAYER M3 ;
        RECT 36.224 18.716 36.256 18.748 ;
  LAYER M1 ;
        RECT 36.288 18.696 36.32 21.204 ;
  LAYER M3 ;
        RECT 36.288 21.152 36.32 21.184 ;
  LAYER M1 ;
        RECT 36.352 18.696 36.384 21.204 ;
  LAYER M3 ;
        RECT 36.352 18.716 36.384 18.748 ;
  LAYER M1 ;
        RECT 36.416 18.696 36.448 21.204 ;
  LAYER M3 ;
        RECT 36.416 21.152 36.448 21.184 ;
  LAYER M1 ;
        RECT 36.48 18.696 36.512 21.204 ;
  LAYER M3 ;
        RECT 36.48 18.716 36.512 18.748 ;
  LAYER M1 ;
        RECT 36.544 18.696 36.576 21.204 ;
  LAYER M3 ;
        RECT 36.544 21.152 36.576 21.184 ;
  LAYER M1 ;
        RECT 36.608 18.696 36.64 21.204 ;
  LAYER M3 ;
        RECT 36.608 18.716 36.64 18.748 ;
  LAYER M1 ;
        RECT 36.672 18.696 36.704 21.204 ;
  LAYER M3 ;
        RECT 36.672 21.152 36.704 21.184 ;
  LAYER M1 ;
        RECT 36.736 18.696 36.768 21.204 ;
  LAYER M3 ;
        RECT 36.736 18.716 36.768 18.748 ;
  LAYER M1 ;
        RECT 36.8 18.696 36.832 21.204 ;
  LAYER M3 ;
        RECT 36.8 21.152 36.832 21.184 ;
  LAYER M1 ;
        RECT 36.864 18.696 36.896 21.204 ;
  LAYER M3 ;
        RECT 36.864 18.716 36.896 18.748 ;
  LAYER M1 ;
        RECT 36.928 18.696 36.96 21.204 ;
  LAYER M3 ;
        RECT 36.928 21.152 36.96 21.184 ;
  LAYER M1 ;
        RECT 36.992 18.696 37.024 21.204 ;
  LAYER M3 ;
        RECT 36.992 18.716 37.024 18.748 ;
  LAYER M1 ;
        RECT 37.056 18.696 37.088 21.204 ;
  LAYER M3 ;
        RECT 37.056 21.152 37.088 21.184 ;
  LAYER M1 ;
        RECT 37.12 18.696 37.152 21.204 ;
  LAYER M3 ;
        RECT 37.12 18.716 37.152 18.748 ;
  LAYER M1 ;
        RECT 37.184 18.696 37.216 21.204 ;
  LAYER M3 ;
        RECT 37.184 21.152 37.216 21.184 ;
  LAYER M1 ;
        RECT 37.248 18.696 37.28 21.204 ;
  LAYER M3 ;
        RECT 37.248 18.716 37.28 18.748 ;
  LAYER M1 ;
        RECT 37.312 18.696 37.344 21.204 ;
  LAYER M3 ;
        RECT 37.312 21.152 37.344 21.184 ;
  LAYER M1 ;
        RECT 37.376 18.696 37.408 21.204 ;
  LAYER M3 ;
        RECT 37.376 18.716 37.408 18.748 ;
  LAYER M1 ;
        RECT 37.44 18.696 37.472 21.204 ;
  LAYER M3 ;
        RECT 37.44 21.152 37.472 21.184 ;
  LAYER M1 ;
        RECT 37.504 18.696 37.536 21.204 ;
  LAYER M3 ;
        RECT 37.504 18.716 37.536 18.748 ;
  LAYER M1 ;
        RECT 37.568 18.696 37.6 21.204 ;
  LAYER M3 ;
        RECT 37.568 21.152 37.6 21.184 ;
  LAYER M1 ;
        RECT 37.632 18.696 37.664 21.204 ;
  LAYER M3 ;
        RECT 37.632 18.716 37.664 18.748 ;
  LAYER M1 ;
        RECT 37.696 18.696 37.728 21.204 ;
  LAYER M3 ;
        RECT 37.696 21.152 37.728 21.184 ;
  LAYER M1 ;
        RECT 37.76 18.696 37.792 21.204 ;
  LAYER M3 ;
        RECT 37.76 18.716 37.792 18.748 ;
  LAYER M1 ;
        RECT 37.824 18.696 37.856 21.204 ;
  LAYER M3 ;
        RECT 37.824 21.152 37.856 21.184 ;
  LAYER M1 ;
        RECT 37.888 18.696 37.92 21.204 ;
  LAYER M3 ;
        RECT 37.888 18.716 37.92 18.748 ;
  LAYER M1 ;
        RECT 37.952 18.696 37.984 21.204 ;
  LAYER M3 ;
        RECT 35.584 21.088 35.616 21.12 ;
  LAYER M2 ;
        RECT 37.952 21.024 37.984 21.056 ;
  LAYER M2 ;
        RECT 35.584 20.96 35.616 20.992 ;
  LAYER M2 ;
        RECT 37.952 20.896 37.984 20.928 ;
  LAYER M2 ;
        RECT 35.584 20.832 35.616 20.864 ;
  LAYER M2 ;
        RECT 37.952 20.768 37.984 20.8 ;
  LAYER M2 ;
        RECT 35.584 20.704 35.616 20.736 ;
  LAYER M2 ;
        RECT 37.952 20.64 37.984 20.672 ;
  LAYER M2 ;
        RECT 35.584 20.576 35.616 20.608 ;
  LAYER M2 ;
        RECT 37.952 20.512 37.984 20.544 ;
  LAYER M2 ;
        RECT 35.584 20.448 35.616 20.48 ;
  LAYER M2 ;
        RECT 37.952 20.384 37.984 20.416 ;
  LAYER M2 ;
        RECT 35.584 20.32 35.616 20.352 ;
  LAYER M2 ;
        RECT 37.952 20.256 37.984 20.288 ;
  LAYER M2 ;
        RECT 35.584 20.192 35.616 20.224 ;
  LAYER M2 ;
        RECT 37.952 20.128 37.984 20.16 ;
  LAYER M2 ;
        RECT 35.584 20.064 35.616 20.096 ;
  LAYER M2 ;
        RECT 37.952 20 37.984 20.032 ;
  LAYER M2 ;
        RECT 35.584 19.936 35.616 19.968 ;
  LAYER M2 ;
        RECT 37.952 19.872 37.984 19.904 ;
  LAYER M2 ;
        RECT 35.584 19.808 35.616 19.84 ;
  LAYER M2 ;
        RECT 37.952 19.744 37.984 19.776 ;
  LAYER M2 ;
        RECT 35.584 19.68 35.616 19.712 ;
  LAYER M2 ;
        RECT 37.952 19.616 37.984 19.648 ;
  LAYER M2 ;
        RECT 35.584 19.552 35.616 19.584 ;
  LAYER M2 ;
        RECT 37.952 19.488 37.984 19.52 ;
  LAYER M2 ;
        RECT 35.584 19.424 35.616 19.456 ;
  LAYER M2 ;
        RECT 37.952 19.36 37.984 19.392 ;
  LAYER M2 ;
        RECT 35.584 19.296 35.616 19.328 ;
  LAYER M2 ;
        RECT 37.952 19.232 37.984 19.264 ;
  LAYER M2 ;
        RECT 35.584 19.168 35.616 19.2 ;
  LAYER M2 ;
        RECT 37.952 19.104 37.984 19.136 ;
  LAYER M2 ;
        RECT 35.584 19.04 35.616 19.072 ;
  LAYER M2 ;
        RECT 37.952 18.976 37.984 19.008 ;
  LAYER M2 ;
        RECT 35.584 18.912 35.616 18.944 ;
  LAYER M2 ;
        RECT 37.952 18.848 37.984 18.88 ;
  LAYER M2 ;
        RECT 35.536 18.648 38.032 21.252 ;
  LAYER M1 ;
        RECT 35.584 15.588 35.616 18.096 ;
  LAYER M3 ;
        RECT 35.584 15.608 35.616 15.64 ;
  LAYER M1 ;
        RECT 35.648 15.588 35.68 18.096 ;
  LAYER M3 ;
        RECT 35.648 18.044 35.68 18.076 ;
  LAYER M1 ;
        RECT 35.712 15.588 35.744 18.096 ;
  LAYER M3 ;
        RECT 35.712 15.608 35.744 15.64 ;
  LAYER M1 ;
        RECT 35.776 15.588 35.808 18.096 ;
  LAYER M3 ;
        RECT 35.776 18.044 35.808 18.076 ;
  LAYER M1 ;
        RECT 35.84 15.588 35.872 18.096 ;
  LAYER M3 ;
        RECT 35.84 15.608 35.872 15.64 ;
  LAYER M1 ;
        RECT 35.904 15.588 35.936 18.096 ;
  LAYER M3 ;
        RECT 35.904 18.044 35.936 18.076 ;
  LAYER M1 ;
        RECT 35.968 15.588 36 18.096 ;
  LAYER M3 ;
        RECT 35.968 15.608 36 15.64 ;
  LAYER M1 ;
        RECT 36.032 15.588 36.064 18.096 ;
  LAYER M3 ;
        RECT 36.032 18.044 36.064 18.076 ;
  LAYER M1 ;
        RECT 36.096 15.588 36.128 18.096 ;
  LAYER M3 ;
        RECT 36.096 15.608 36.128 15.64 ;
  LAYER M1 ;
        RECT 36.16 15.588 36.192 18.096 ;
  LAYER M3 ;
        RECT 36.16 18.044 36.192 18.076 ;
  LAYER M1 ;
        RECT 36.224 15.588 36.256 18.096 ;
  LAYER M3 ;
        RECT 36.224 15.608 36.256 15.64 ;
  LAYER M1 ;
        RECT 36.288 15.588 36.32 18.096 ;
  LAYER M3 ;
        RECT 36.288 18.044 36.32 18.076 ;
  LAYER M1 ;
        RECT 36.352 15.588 36.384 18.096 ;
  LAYER M3 ;
        RECT 36.352 15.608 36.384 15.64 ;
  LAYER M1 ;
        RECT 36.416 15.588 36.448 18.096 ;
  LAYER M3 ;
        RECT 36.416 18.044 36.448 18.076 ;
  LAYER M1 ;
        RECT 36.48 15.588 36.512 18.096 ;
  LAYER M3 ;
        RECT 36.48 15.608 36.512 15.64 ;
  LAYER M1 ;
        RECT 36.544 15.588 36.576 18.096 ;
  LAYER M3 ;
        RECT 36.544 18.044 36.576 18.076 ;
  LAYER M1 ;
        RECT 36.608 15.588 36.64 18.096 ;
  LAYER M3 ;
        RECT 36.608 15.608 36.64 15.64 ;
  LAYER M1 ;
        RECT 36.672 15.588 36.704 18.096 ;
  LAYER M3 ;
        RECT 36.672 18.044 36.704 18.076 ;
  LAYER M1 ;
        RECT 36.736 15.588 36.768 18.096 ;
  LAYER M3 ;
        RECT 36.736 15.608 36.768 15.64 ;
  LAYER M1 ;
        RECT 36.8 15.588 36.832 18.096 ;
  LAYER M3 ;
        RECT 36.8 18.044 36.832 18.076 ;
  LAYER M1 ;
        RECT 36.864 15.588 36.896 18.096 ;
  LAYER M3 ;
        RECT 36.864 15.608 36.896 15.64 ;
  LAYER M1 ;
        RECT 36.928 15.588 36.96 18.096 ;
  LAYER M3 ;
        RECT 36.928 18.044 36.96 18.076 ;
  LAYER M1 ;
        RECT 36.992 15.588 37.024 18.096 ;
  LAYER M3 ;
        RECT 36.992 15.608 37.024 15.64 ;
  LAYER M1 ;
        RECT 37.056 15.588 37.088 18.096 ;
  LAYER M3 ;
        RECT 37.056 18.044 37.088 18.076 ;
  LAYER M1 ;
        RECT 37.12 15.588 37.152 18.096 ;
  LAYER M3 ;
        RECT 37.12 15.608 37.152 15.64 ;
  LAYER M1 ;
        RECT 37.184 15.588 37.216 18.096 ;
  LAYER M3 ;
        RECT 37.184 18.044 37.216 18.076 ;
  LAYER M1 ;
        RECT 37.248 15.588 37.28 18.096 ;
  LAYER M3 ;
        RECT 37.248 15.608 37.28 15.64 ;
  LAYER M1 ;
        RECT 37.312 15.588 37.344 18.096 ;
  LAYER M3 ;
        RECT 37.312 18.044 37.344 18.076 ;
  LAYER M1 ;
        RECT 37.376 15.588 37.408 18.096 ;
  LAYER M3 ;
        RECT 37.376 15.608 37.408 15.64 ;
  LAYER M1 ;
        RECT 37.44 15.588 37.472 18.096 ;
  LAYER M3 ;
        RECT 37.44 18.044 37.472 18.076 ;
  LAYER M1 ;
        RECT 37.504 15.588 37.536 18.096 ;
  LAYER M3 ;
        RECT 37.504 15.608 37.536 15.64 ;
  LAYER M1 ;
        RECT 37.568 15.588 37.6 18.096 ;
  LAYER M3 ;
        RECT 37.568 18.044 37.6 18.076 ;
  LAYER M1 ;
        RECT 37.632 15.588 37.664 18.096 ;
  LAYER M3 ;
        RECT 37.632 15.608 37.664 15.64 ;
  LAYER M1 ;
        RECT 37.696 15.588 37.728 18.096 ;
  LAYER M3 ;
        RECT 37.696 18.044 37.728 18.076 ;
  LAYER M1 ;
        RECT 37.76 15.588 37.792 18.096 ;
  LAYER M3 ;
        RECT 37.76 15.608 37.792 15.64 ;
  LAYER M1 ;
        RECT 37.824 15.588 37.856 18.096 ;
  LAYER M3 ;
        RECT 37.824 18.044 37.856 18.076 ;
  LAYER M1 ;
        RECT 37.888 15.588 37.92 18.096 ;
  LAYER M3 ;
        RECT 37.888 15.608 37.92 15.64 ;
  LAYER M1 ;
        RECT 37.952 15.588 37.984 18.096 ;
  LAYER M3 ;
        RECT 35.584 17.98 35.616 18.012 ;
  LAYER M2 ;
        RECT 37.952 17.916 37.984 17.948 ;
  LAYER M2 ;
        RECT 35.584 17.852 35.616 17.884 ;
  LAYER M2 ;
        RECT 37.952 17.788 37.984 17.82 ;
  LAYER M2 ;
        RECT 35.584 17.724 35.616 17.756 ;
  LAYER M2 ;
        RECT 37.952 17.66 37.984 17.692 ;
  LAYER M2 ;
        RECT 35.584 17.596 35.616 17.628 ;
  LAYER M2 ;
        RECT 37.952 17.532 37.984 17.564 ;
  LAYER M2 ;
        RECT 35.584 17.468 35.616 17.5 ;
  LAYER M2 ;
        RECT 37.952 17.404 37.984 17.436 ;
  LAYER M2 ;
        RECT 35.584 17.34 35.616 17.372 ;
  LAYER M2 ;
        RECT 37.952 17.276 37.984 17.308 ;
  LAYER M2 ;
        RECT 35.584 17.212 35.616 17.244 ;
  LAYER M2 ;
        RECT 37.952 17.148 37.984 17.18 ;
  LAYER M2 ;
        RECT 35.584 17.084 35.616 17.116 ;
  LAYER M2 ;
        RECT 37.952 17.02 37.984 17.052 ;
  LAYER M2 ;
        RECT 35.584 16.956 35.616 16.988 ;
  LAYER M2 ;
        RECT 37.952 16.892 37.984 16.924 ;
  LAYER M2 ;
        RECT 35.584 16.828 35.616 16.86 ;
  LAYER M2 ;
        RECT 37.952 16.764 37.984 16.796 ;
  LAYER M2 ;
        RECT 35.584 16.7 35.616 16.732 ;
  LAYER M2 ;
        RECT 37.952 16.636 37.984 16.668 ;
  LAYER M2 ;
        RECT 35.584 16.572 35.616 16.604 ;
  LAYER M2 ;
        RECT 37.952 16.508 37.984 16.54 ;
  LAYER M2 ;
        RECT 35.584 16.444 35.616 16.476 ;
  LAYER M2 ;
        RECT 37.952 16.38 37.984 16.412 ;
  LAYER M2 ;
        RECT 35.584 16.316 35.616 16.348 ;
  LAYER M2 ;
        RECT 37.952 16.252 37.984 16.284 ;
  LAYER M2 ;
        RECT 35.584 16.188 35.616 16.22 ;
  LAYER M2 ;
        RECT 37.952 16.124 37.984 16.156 ;
  LAYER M2 ;
        RECT 35.584 16.06 35.616 16.092 ;
  LAYER M2 ;
        RECT 37.952 15.996 37.984 16.028 ;
  LAYER M2 ;
        RECT 35.584 15.932 35.616 15.964 ;
  LAYER M2 ;
        RECT 37.952 15.868 37.984 15.9 ;
  LAYER M2 ;
        RECT 35.584 15.804 35.616 15.836 ;
  LAYER M2 ;
        RECT 37.952 15.74 37.984 15.772 ;
  LAYER M2 ;
        RECT 35.536 15.54 38.032 18.144 ;
  LAYER M1 ;
        RECT 38.56 28.02 38.592 30.528 ;
  LAYER M3 ;
        RECT 38.56 28.04 38.592 28.072 ;
  LAYER M1 ;
        RECT 38.624 28.02 38.656 30.528 ;
  LAYER M3 ;
        RECT 38.624 30.476 38.656 30.508 ;
  LAYER M1 ;
        RECT 38.688 28.02 38.72 30.528 ;
  LAYER M3 ;
        RECT 38.688 28.04 38.72 28.072 ;
  LAYER M1 ;
        RECT 38.752 28.02 38.784 30.528 ;
  LAYER M3 ;
        RECT 38.752 30.476 38.784 30.508 ;
  LAYER M1 ;
        RECT 38.816 28.02 38.848 30.528 ;
  LAYER M3 ;
        RECT 38.816 28.04 38.848 28.072 ;
  LAYER M1 ;
        RECT 38.88 28.02 38.912 30.528 ;
  LAYER M3 ;
        RECT 38.88 30.476 38.912 30.508 ;
  LAYER M1 ;
        RECT 38.944 28.02 38.976 30.528 ;
  LAYER M3 ;
        RECT 38.944 28.04 38.976 28.072 ;
  LAYER M1 ;
        RECT 39.008 28.02 39.04 30.528 ;
  LAYER M3 ;
        RECT 39.008 30.476 39.04 30.508 ;
  LAYER M1 ;
        RECT 39.072 28.02 39.104 30.528 ;
  LAYER M3 ;
        RECT 39.072 28.04 39.104 28.072 ;
  LAYER M1 ;
        RECT 39.136 28.02 39.168 30.528 ;
  LAYER M3 ;
        RECT 39.136 30.476 39.168 30.508 ;
  LAYER M1 ;
        RECT 39.2 28.02 39.232 30.528 ;
  LAYER M3 ;
        RECT 39.2 28.04 39.232 28.072 ;
  LAYER M1 ;
        RECT 39.264 28.02 39.296 30.528 ;
  LAYER M3 ;
        RECT 39.264 30.476 39.296 30.508 ;
  LAYER M1 ;
        RECT 39.328 28.02 39.36 30.528 ;
  LAYER M3 ;
        RECT 39.328 28.04 39.36 28.072 ;
  LAYER M1 ;
        RECT 39.392 28.02 39.424 30.528 ;
  LAYER M3 ;
        RECT 39.392 30.476 39.424 30.508 ;
  LAYER M1 ;
        RECT 39.456 28.02 39.488 30.528 ;
  LAYER M3 ;
        RECT 39.456 28.04 39.488 28.072 ;
  LAYER M1 ;
        RECT 39.52 28.02 39.552 30.528 ;
  LAYER M3 ;
        RECT 39.52 30.476 39.552 30.508 ;
  LAYER M1 ;
        RECT 39.584 28.02 39.616 30.528 ;
  LAYER M3 ;
        RECT 39.584 28.04 39.616 28.072 ;
  LAYER M1 ;
        RECT 39.648 28.02 39.68 30.528 ;
  LAYER M3 ;
        RECT 39.648 30.476 39.68 30.508 ;
  LAYER M1 ;
        RECT 39.712 28.02 39.744 30.528 ;
  LAYER M3 ;
        RECT 39.712 28.04 39.744 28.072 ;
  LAYER M1 ;
        RECT 39.776 28.02 39.808 30.528 ;
  LAYER M3 ;
        RECT 39.776 30.476 39.808 30.508 ;
  LAYER M1 ;
        RECT 39.84 28.02 39.872 30.528 ;
  LAYER M3 ;
        RECT 39.84 28.04 39.872 28.072 ;
  LAYER M1 ;
        RECT 39.904 28.02 39.936 30.528 ;
  LAYER M3 ;
        RECT 39.904 30.476 39.936 30.508 ;
  LAYER M1 ;
        RECT 39.968 28.02 40 30.528 ;
  LAYER M3 ;
        RECT 39.968 28.04 40 28.072 ;
  LAYER M1 ;
        RECT 40.032 28.02 40.064 30.528 ;
  LAYER M3 ;
        RECT 40.032 30.476 40.064 30.508 ;
  LAYER M1 ;
        RECT 40.096 28.02 40.128 30.528 ;
  LAYER M3 ;
        RECT 40.096 28.04 40.128 28.072 ;
  LAYER M1 ;
        RECT 40.16 28.02 40.192 30.528 ;
  LAYER M3 ;
        RECT 40.16 30.476 40.192 30.508 ;
  LAYER M1 ;
        RECT 40.224 28.02 40.256 30.528 ;
  LAYER M3 ;
        RECT 40.224 28.04 40.256 28.072 ;
  LAYER M1 ;
        RECT 40.288 28.02 40.32 30.528 ;
  LAYER M3 ;
        RECT 40.288 30.476 40.32 30.508 ;
  LAYER M1 ;
        RECT 40.352 28.02 40.384 30.528 ;
  LAYER M3 ;
        RECT 40.352 28.04 40.384 28.072 ;
  LAYER M1 ;
        RECT 40.416 28.02 40.448 30.528 ;
  LAYER M3 ;
        RECT 40.416 30.476 40.448 30.508 ;
  LAYER M1 ;
        RECT 40.48 28.02 40.512 30.528 ;
  LAYER M3 ;
        RECT 40.48 28.04 40.512 28.072 ;
  LAYER M1 ;
        RECT 40.544 28.02 40.576 30.528 ;
  LAYER M3 ;
        RECT 40.544 30.476 40.576 30.508 ;
  LAYER M1 ;
        RECT 40.608 28.02 40.64 30.528 ;
  LAYER M3 ;
        RECT 40.608 28.04 40.64 28.072 ;
  LAYER M1 ;
        RECT 40.672 28.02 40.704 30.528 ;
  LAYER M3 ;
        RECT 40.672 30.476 40.704 30.508 ;
  LAYER M1 ;
        RECT 40.736 28.02 40.768 30.528 ;
  LAYER M3 ;
        RECT 40.736 28.04 40.768 28.072 ;
  LAYER M1 ;
        RECT 40.8 28.02 40.832 30.528 ;
  LAYER M3 ;
        RECT 40.8 30.476 40.832 30.508 ;
  LAYER M1 ;
        RECT 40.864 28.02 40.896 30.528 ;
  LAYER M3 ;
        RECT 40.864 28.04 40.896 28.072 ;
  LAYER M1 ;
        RECT 40.928 28.02 40.96 30.528 ;
  LAYER M3 ;
        RECT 38.56 30.412 38.592 30.444 ;
  LAYER M2 ;
        RECT 40.928 30.348 40.96 30.38 ;
  LAYER M2 ;
        RECT 38.56 30.284 38.592 30.316 ;
  LAYER M2 ;
        RECT 40.928 30.22 40.96 30.252 ;
  LAYER M2 ;
        RECT 38.56 30.156 38.592 30.188 ;
  LAYER M2 ;
        RECT 40.928 30.092 40.96 30.124 ;
  LAYER M2 ;
        RECT 38.56 30.028 38.592 30.06 ;
  LAYER M2 ;
        RECT 40.928 29.964 40.96 29.996 ;
  LAYER M2 ;
        RECT 38.56 29.9 38.592 29.932 ;
  LAYER M2 ;
        RECT 40.928 29.836 40.96 29.868 ;
  LAYER M2 ;
        RECT 38.56 29.772 38.592 29.804 ;
  LAYER M2 ;
        RECT 40.928 29.708 40.96 29.74 ;
  LAYER M2 ;
        RECT 38.56 29.644 38.592 29.676 ;
  LAYER M2 ;
        RECT 40.928 29.58 40.96 29.612 ;
  LAYER M2 ;
        RECT 38.56 29.516 38.592 29.548 ;
  LAYER M2 ;
        RECT 40.928 29.452 40.96 29.484 ;
  LAYER M2 ;
        RECT 38.56 29.388 38.592 29.42 ;
  LAYER M2 ;
        RECT 40.928 29.324 40.96 29.356 ;
  LAYER M2 ;
        RECT 38.56 29.26 38.592 29.292 ;
  LAYER M2 ;
        RECT 40.928 29.196 40.96 29.228 ;
  LAYER M2 ;
        RECT 38.56 29.132 38.592 29.164 ;
  LAYER M2 ;
        RECT 40.928 29.068 40.96 29.1 ;
  LAYER M2 ;
        RECT 38.56 29.004 38.592 29.036 ;
  LAYER M2 ;
        RECT 40.928 28.94 40.96 28.972 ;
  LAYER M2 ;
        RECT 38.56 28.876 38.592 28.908 ;
  LAYER M2 ;
        RECT 40.928 28.812 40.96 28.844 ;
  LAYER M2 ;
        RECT 38.56 28.748 38.592 28.78 ;
  LAYER M2 ;
        RECT 40.928 28.684 40.96 28.716 ;
  LAYER M2 ;
        RECT 38.56 28.62 38.592 28.652 ;
  LAYER M2 ;
        RECT 40.928 28.556 40.96 28.588 ;
  LAYER M2 ;
        RECT 38.56 28.492 38.592 28.524 ;
  LAYER M2 ;
        RECT 40.928 28.428 40.96 28.46 ;
  LAYER M2 ;
        RECT 38.56 28.364 38.592 28.396 ;
  LAYER M2 ;
        RECT 40.928 28.3 40.96 28.332 ;
  LAYER M2 ;
        RECT 38.56 28.236 38.592 28.268 ;
  LAYER M2 ;
        RECT 40.928 28.172 40.96 28.204 ;
  LAYER M2 ;
        RECT 38.512 27.972 41.008 30.576 ;
  LAYER M1 ;
        RECT 38.56 24.912 38.592 27.42 ;
  LAYER M3 ;
        RECT 38.56 24.932 38.592 24.964 ;
  LAYER M1 ;
        RECT 38.624 24.912 38.656 27.42 ;
  LAYER M3 ;
        RECT 38.624 27.368 38.656 27.4 ;
  LAYER M1 ;
        RECT 38.688 24.912 38.72 27.42 ;
  LAYER M3 ;
        RECT 38.688 24.932 38.72 24.964 ;
  LAYER M1 ;
        RECT 38.752 24.912 38.784 27.42 ;
  LAYER M3 ;
        RECT 38.752 27.368 38.784 27.4 ;
  LAYER M1 ;
        RECT 38.816 24.912 38.848 27.42 ;
  LAYER M3 ;
        RECT 38.816 24.932 38.848 24.964 ;
  LAYER M1 ;
        RECT 38.88 24.912 38.912 27.42 ;
  LAYER M3 ;
        RECT 38.88 27.368 38.912 27.4 ;
  LAYER M1 ;
        RECT 38.944 24.912 38.976 27.42 ;
  LAYER M3 ;
        RECT 38.944 24.932 38.976 24.964 ;
  LAYER M1 ;
        RECT 39.008 24.912 39.04 27.42 ;
  LAYER M3 ;
        RECT 39.008 27.368 39.04 27.4 ;
  LAYER M1 ;
        RECT 39.072 24.912 39.104 27.42 ;
  LAYER M3 ;
        RECT 39.072 24.932 39.104 24.964 ;
  LAYER M1 ;
        RECT 39.136 24.912 39.168 27.42 ;
  LAYER M3 ;
        RECT 39.136 27.368 39.168 27.4 ;
  LAYER M1 ;
        RECT 39.2 24.912 39.232 27.42 ;
  LAYER M3 ;
        RECT 39.2 24.932 39.232 24.964 ;
  LAYER M1 ;
        RECT 39.264 24.912 39.296 27.42 ;
  LAYER M3 ;
        RECT 39.264 27.368 39.296 27.4 ;
  LAYER M1 ;
        RECT 39.328 24.912 39.36 27.42 ;
  LAYER M3 ;
        RECT 39.328 24.932 39.36 24.964 ;
  LAYER M1 ;
        RECT 39.392 24.912 39.424 27.42 ;
  LAYER M3 ;
        RECT 39.392 27.368 39.424 27.4 ;
  LAYER M1 ;
        RECT 39.456 24.912 39.488 27.42 ;
  LAYER M3 ;
        RECT 39.456 24.932 39.488 24.964 ;
  LAYER M1 ;
        RECT 39.52 24.912 39.552 27.42 ;
  LAYER M3 ;
        RECT 39.52 27.368 39.552 27.4 ;
  LAYER M1 ;
        RECT 39.584 24.912 39.616 27.42 ;
  LAYER M3 ;
        RECT 39.584 24.932 39.616 24.964 ;
  LAYER M1 ;
        RECT 39.648 24.912 39.68 27.42 ;
  LAYER M3 ;
        RECT 39.648 27.368 39.68 27.4 ;
  LAYER M1 ;
        RECT 39.712 24.912 39.744 27.42 ;
  LAYER M3 ;
        RECT 39.712 24.932 39.744 24.964 ;
  LAYER M1 ;
        RECT 39.776 24.912 39.808 27.42 ;
  LAYER M3 ;
        RECT 39.776 27.368 39.808 27.4 ;
  LAYER M1 ;
        RECT 39.84 24.912 39.872 27.42 ;
  LAYER M3 ;
        RECT 39.84 24.932 39.872 24.964 ;
  LAYER M1 ;
        RECT 39.904 24.912 39.936 27.42 ;
  LAYER M3 ;
        RECT 39.904 27.368 39.936 27.4 ;
  LAYER M1 ;
        RECT 39.968 24.912 40 27.42 ;
  LAYER M3 ;
        RECT 39.968 24.932 40 24.964 ;
  LAYER M1 ;
        RECT 40.032 24.912 40.064 27.42 ;
  LAYER M3 ;
        RECT 40.032 27.368 40.064 27.4 ;
  LAYER M1 ;
        RECT 40.096 24.912 40.128 27.42 ;
  LAYER M3 ;
        RECT 40.096 24.932 40.128 24.964 ;
  LAYER M1 ;
        RECT 40.16 24.912 40.192 27.42 ;
  LAYER M3 ;
        RECT 40.16 27.368 40.192 27.4 ;
  LAYER M1 ;
        RECT 40.224 24.912 40.256 27.42 ;
  LAYER M3 ;
        RECT 40.224 24.932 40.256 24.964 ;
  LAYER M1 ;
        RECT 40.288 24.912 40.32 27.42 ;
  LAYER M3 ;
        RECT 40.288 27.368 40.32 27.4 ;
  LAYER M1 ;
        RECT 40.352 24.912 40.384 27.42 ;
  LAYER M3 ;
        RECT 40.352 24.932 40.384 24.964 ;
  LAYER M1 ;
        RECT 40.416 24.912 40.448 27.42 ;
  LAYER M3 ;
        RECT 40.416 27.368 40.448 27.4 ;
  LAYER M1 ;
        RECT 40.48 24.912 40.512 27.42 ;
  LAYER M3 ;
        RECT 40.48 24.932 40.512 24.964 ;
  LAYER M1 ;
        RECT 40.544 24.912 40.576 27.42 ;
  LAYER M3 ;
        RECT 40.544 27.368 40.576 27.4 ;
  LAYER M1 ;
        RECT 40.608 24.912 40.64 27.42 ;
  LAYER M3 ;
        RECT 40.608 24.932 40.64 24.964 ;
  LAYER M1 ;
        RECT 40.672 24.912 40.704 27.42 ;
  LAYER M3 ;
        RECT 40.672 27.368 40.704 27.4 ;
  LAYER M1 ;
        RECT 40.736 24.912 40.768 27.42 ;
  LAYER M3 ;
        RECT 40.736 24.932 40.768 24.964 ;
  LAYER M1 ;
        RECT 40.8 24.912 40.832 27.42 ;
  LAYER M3 ;
        RECT 40.8 27.368 40.832 27.4 ;
  LAYER M1 ;
        RECT 40.864 24.912 40.896 27.42 ;
  LAYER M3 ;
        RECT 40.864 24.932 40.896 24.964 ;
  LAYER M1 ;
        RECT 40.928 24.912 40.96 27.42 ;
  LAYER M3 ;
        RECT 38.56 27.304 38.592 27.336 ;
  LAYER M2 ;
        RECT 40.928 27.24 40.96 27.272 ;
  LAYER M2 ;
        RECT 38.56 27.176 38.592 27.208 ;
  LAYER M2 ;
        RECT 40.928 27.112 40.96 27.144 ;
  LAYER M2 ;
        RECT 38.56 27.048 38.592 27.08 ;
  LAYER M2 ;
        RECT 40.928 26.984 40.96 27.016 ;
  LAYER M2 ;
        RECT 38.56 26.92 38.592 26.952 ;
  LAYER M2 ;
        RECT 40.928 26.856 40.96 26.888 ;
  LAYER M2 ;
        RECT 38.56 26.792 38.592 26.824 ;
  LAYER M2 ;
        RECT 40.928 26.728 40.96 26.76 ;
  LAYER M2 ;
        RECT 38.56 26.664 38.592 26.696 ;
  LAYER M2 ;
        RECT 40.928 26.6 40.96 26.632 ;
  LAYER M2 ;
        RECT 38.56 26.536 38.592 26.568 ;
  LAYER M2 ;
        RECT 40.928 26.472 40.96 26.504 ;
  LAYER M2 ;
        RECT 38.56 26.408 38.592 26.44 ;
  LAYER M2 ;
        RECT 40.928 26.344 40.96 26.376 ;
  LAYER M2 ;
        RECT 38.56 26.28 38.592 26.312 ;
  LAYER M2 ;
        RECT 40.928 26.216 40.96 26.248 ;
  LAYER M2 ;
        RECT 38.56 26.152 38.592 26.184 ;
  LAYER M2 ;
        RECT 40.928 26.088 40.96 26.12 ;
  LAYER M2 ;
        RECT 38.56 26.024 38.592 26.056 ;
  LAYER M2 ;
        RECT 40.928 25.96 40.96 25.992 ;
  LAYER M2 ;
        RECT 38.56 25.896 38.592 25.928 ;
  LAYER M2 ;
        RECT 40.928 25.832 40.96 25.864 ;
  LAYER M2 ;
        RECT 38.56 25.768 38.592 25.8 ;
  LAYER M2 ;
        RECT 40.928 25.704 40.96 25.736 ;
  LAYER M2 ;
        RECT 38.56 25.64 38.592 25.672 ;
  LAYER M2 ;
        RECT 40.928 25.576 40.96 25.608 ;
  LAYER M2 ;
        RECT 38.56 25.512 38.592 25.544 ;
  LAYER M2 ;
        RECT 40.928 25.448 40.96 25.48 ;
  LAYER M2 ;
        RECT 38.56 25.384 38.592 25.416 ;
  LAYER M2 ;
        RECT 40.928 25.32 40.96 25.352 ;
  LAYER M2 ;
        RECT 38.56 25.256 38.592 25.288 ;
  LAYER M2 ;
        RECT 40.928 25.192 40.96 25.224 ;
  LAYER M2 ;
        RECT 38.56 25.128 38.592 25.16 ;
  LAYER M2 ;
        RECT 40.928 25.064 40.96 25.096 ;
  LAYER M2 ;
        RECT 38.512 24.864 41.008 27.468 ;
  LAYER M1 ;
        RECT 38.56 21.804 38.592 24.312 ;
  LAYER M3 ;
        RECT 38.56 21.824 38.592 21.856 ;
  LAYER M1 ;
        RECT 38.624 21.804 38.656 24.312 ;
  LAYER M3 ;
        RECT 38.624 24.26 38.656 24.292 ;
  LAYER M1 ;
        RECT 38.688 21.804 38.72 24.312 ;
  LAYER M3 ;
        RECT 38.688 21.824 38.72 21.856 ;
  LAYER M1 ;
        RECT 38.752 21.804 38.784 24.312 ;
  LAYER M3 ;
        RECT 38.752 24.26 38.784 24.292 ;
  LAYER M1 ;
        RECT 38.816 21.804 38.848 24.312 ;
  LAYER M3 ;
        RECT 38.816 21.824 38.848 21.856 ;
  LAYER M1 ;
        RECT 38.88 21.804 38.912 24.312 ;
  LAYER M3 ;
        RECT 38.88 24.26 38.912 24.292 ;
  LAYER M1 ;
        RECT 38.944 21.804 38.976 24.312 ;
  LAYER M3 ;
        RECT 38.944 21.824 38.976 21.856 ;
  LAYER M1 ;
        RECT 39.008 21.804 39.04 24.312 ;
  LAYER M3 ;
        RECT 39.008 24.26 39.04 24.292 ;
  LAYER M1 ;
        RECT 39.072 21.804 39.104 24.312 ;
  LAYER M3 ;
        RECT 39.072 21.824 39.104 21.856 ;
  LAYER M1 ;
        RECT 39.136 21.804 39.168 24.312 ;
  LAYER M3 ;
        RECT 39.136 24.26 39.168 24.292 ;
  LAYER M1 ;
        RECT 39.2 21.804 39.232 24.312 ;
  LAYER M3 ;
        RECT 39.2 21.824 39.232 21.856 ;
  LAYER M1 ;
        RECT 39.264 21.804 39.296 24.312 ;
  LAYER M3 ;
        RECT 39.264 24.26 39.296 24.292 ;
  LAYER M1 ;
        RECT 39.328 21.804 39.36 24.312 ;
  LAYER M3 ;
        RECT 39.328 21.824 39.36 21.856 ;
  LAYER M1 ;
        RECT 39.392 21.804 39.424 24.312 ;
  LAYER M3 ;
        RECT 39.392 24.26 39.424 24.292 ;
  LAYER M1 ;
        RECT 39.456 21.804 39.488 24.312 ;
  LAYER M3 ;
        RECT 39.456 21.824 39.488 21.856 ;
  LAYER M1 ;
        RECT 39.52 21.804 39.552 24.312 ;
  LAYER M3 ;
        RECT 39.52 24.26 39.552 24.292 ;
  LAYER M1 ;
        RECT 39.584 21.804 39.616 24.312 ;
  LAYER M3 ;
        RECT 39.584 21.824 39.616 21.856 ;
  LAYER M1 ;
        RECT 39.648 21.804 39.68 24.312 ;
  LAYER M3 ;
        RECT 39.648 24.26 39.68 24.292 ;
  LAYER M1 ;
        RECT 39.712 21.804 39.744 24.312 ;
  LAYER M3 ;
        RECT 39.712 21.824 39.744 21.856 ;
  LAYER M1 ;
        RECT 39.776 21.804 39.808 24.312 ;
  LAYER M3 ;
        RECT 39.776 24.26 39.808 24.292 ;
  LAYER M1 ;
        RECT 39.84 21.804 39.872 24.312 ;
  LAYER M3 ;
        RECT 39.84 21.824 39.872 21.856 ;
  LAYER M1 ;
        RECT 39.904 21.804 39.936 24.312 ;
  LAYER M3 ;
        RECT 39.904 24.26 39.936 24.292 ;
  LAYER M1 ;
        RECT 39.968 21.804 40 24.312 ;
  LAYER M3 ;
        RECT 39.968 21.824 40 21.856 ;
  LAYER M1 ;
        RECT 40.032 21.804 40.064 24.312 ;
  LAYER M3 ;
        RECT 40.032 24.26 40.064 24.292 ;
  LAYER M1 ;
        RECT 40.096 21.804 40.128 24.312 ;
  LAYER M3 ;
        RECT 40.096 21.824 40.128 21.856 ;
  LAYER M1 ;
        RECT 40.16 21.804 40.192 24.312 ;
  LAYER M3 ;
        RECT 40.16 24.26 40.192 24.292 ;
  LAYER M1 ;
        RECT 40.224 21.804 40.256 24.312 ;
  LAYER M3 ;
        RECT 40.224 21.824 40.256 21.856 ;
  LAYER M1 ;
        RECT 40.288 21.804 40.32 24.312 ;
  LAYER M3 ;
        RECT 40.288 24.26 40.32 24.292 ;
  LAYER M1 ;
        RECT 40.352 21.804 40.384 24.312 ;
  LAYER M3 ;
        RECT 40.352 21.824 40.384 21.856 ;
  LAYER M1 ;
        RECT 40.416 21.804 40.448 24.312 ;
  LAYER M3 ;
        RECT 40.416 24.26 40.448 24.292 ;
  LAYER M1 ;
        RECT 40.48 21.804 40.512 24.312 ;
  LAYER M3 ;
        RECT 40.48 21.824 40.512 21.856 ;
  LAYER M1 ;
        RECT 40.544 21.804 40.576 24.312 ;
  LAYER M3 ;
        RECT 40.544 24.26 40.576 24.292 ;
  LAYER M1 ;
        RECT 40.608 21.804 40.64 24.312 ;
  LAYER M3 ;
        RECT 40.608 21.824 40.64 21.856 ;
  LAYER M1 ;
        RECT 40.672 21.804 40.704 24.312 ;
  LAYER M3 ;
        RECT 40.672 24.26 40.704 24.292 ;
  LAYER M1 ;
        RECT 40.736 21.804 40.768 24.312 ;
  LAYER M3 ;
        RECT 40.736 21.824 40.768 21.856 ;
  LAYER M1 ;
        RECT 40.8 21.804 40.832 24.312 ;
  LAYER M3 ;
        RECT 40.8 24.26 40.832 24.292 ;
  LAYER M1 ;
        RECT 40.864 21.804 40.896 24.312 ;
  LAYER M3 ;
        RECT 40.864 21.824 40.896 21.856 ;
  LAYER M1 ;
        RECT 40.928 21.804 40.96 24.312 ;
  LAYER M3 ;
        RECT 38.56 24.196 38.592 24.228 ;
  LAYER M2 ;
        RECT 40.928 24.132 40.96 24.164 ;
  LAYER M2 ;
        RECT 38.56 24.068 38.592 24.1 ;
  LAYER M2 ;
        RECT 40.928 24.004 40.96 24.036 ;
  LAYER M2 ;
        RECT 38.56 23.94 38.592 23.972 ;
  LAYER M2 ;
        RECT 40.928 23.876 40.96 23.908 ;
  LAYER M2 ;
        RECT 38.56 23.812 38.592 23.844 ;
  LAYER M2 ;
        RECT 40.928 23.748 40.96 23.78 ;
  LAYER M2 ;
        RECT 38.56 23.684 38.592 23.716 ;
  LAYER M2 ;
        RECT 40.928 23.62 40.96 23.652 ;
  LAYER M2 ;
        RECT 38.56 23.556 38.592 23.588 ;
  LAYER M2 ;
        RECT 40.928 23.492 40.96 23.524 ;
  LAYER M2 ;
        RECT 38.56 23.428 38.592 23.46 ;
  LAYER M2 ;
        RECT 40.928 23.364 40.96 23.396 ;
  LAYER M2 ;
        RECT 38.56 23.3 38.592 23.332 ;
  LAYER M2 ;
        RECT 40.928 23.236 40.96 23.268 ;
  LAYER M2 ;
        RECT 38.56 23.172 38.592 23.204 ;
  LAYER M2 ;
        RECT 40.928 23.108 40.96 23.14 ;
  LAYER M2 ;
        RECT 38.56 23.044 38.592 23.076 ;
  LAYER M2 ;
        RECT 40.928 22.98 40.96 23.012 ;
  LAYER M2 ;
        RECT 38.56 22.916 38.592 22.948 ;
  LAYER M2 ;
        RECT 40.928 22.852 40.96 22.884 ;
  LAYER M2 ;
        RECT 38.56 22.788 38.592 22.82 ;
  LAYER M2 ;
        RECT 40.928 22.724 40.96 22.756 ;
  LAYER M2 ;
        RECT 38.56 22.66 38.592 22.692 ;
  LAYER M2 ;
        RECT 40.928 22.596 40.96 22.628 ;
  LAYER M2 ;
        RECT 38.56 22.532 38.592 22.564 ;
  LAYER M2 ;
        RECT 40.928 22.468 40.96 22.5 ;
  LAYER M2 ;
        RECT 38.56 22.404 38.592 22.436 ;
  LAYER M2 ;
        RECT 40.928 22.34 40.96 22.372 ;
  LAYER M2 ;
        RECT 38.56 22.276 38.592 22.308 ;
  LAYER M2 ;
        RECT 40.928 22.212 40.96 22.244 ;
  LAYER M2 ;
        RECT 38.56 22.148 38.592 22.18 ;
  LAYER M2 ;
        RECT 40.928 22.084 40.96 22.116 ;
  LAYER M2 ;
        RECT 38.56 22.02 38.592 22.052 ;
  LAYER M2 ;
        RECT 40.928 21.956 40.96 21.988 ;
  LAYER M2 ;
        RECT 38.512 21.756 41.008 24.36 ;
  LAYER M1 ;
        RECT 38.56 18.696 38.592 21.204 ;
  LAYER M3 ;
        RECT 38.56 18.716 38.592 18.748 ;
  LAYER M1 ;
        RECT 38.624 18.696 38.656 21.204 ;
  LAYER M3 ;
        RECT 38.624 21.152 38.656 21.184 ;
  LAYER M1 ;
        RECT 38.688 18.696 38.72 21.204 ;
  LAYER M3 ;
        RECT 38.688 18.716 38.72 18.748 ;
  LAYER M1 ;
        RECT 38.752 18.696 38.784 21.204 ;
  LAYER M3 ;
        RECT 38.752 21.152 38.784 21.184 ;
  LAYER M1 ;
        RECT 38.816 18.696 38.848 21.204 ;
  LAYER M3 ;
        RECT 38.816 18.716 38.848 18.748 ;
  LAYER M1 ;
        RECT 38.88 18.696 38.912 21.204 ;
  LAYER M3 ;
        RECT 38.88 21.152 38.912 21.184 ;
  LAYER M1 ;
        RECT 38.944 18.696 38.976 21.204 ;
  LAYER M3 ;
        RECT 38.944 18.716 38.976 18.748 ;
  LAYER M1 ;
        RECT 39.008 18.696 39.04 21.204 ;
  LAYER M3 ;
        RECT 39.008 21.152 39.04 21.184 ;
  LAYER M1 ;
        RECT 39.072 18.696 39.104 21.204 ;
  LAYER M3 ;
        RECT 39.072 18.716 39.104 18.748 ;
  LAYER M1 ;
        RECT 39.136 18.696 39.168 21.204 ;
  LAYER M3 ;
        RECT 39.136 21.152 39.168 21.184 ;
  LAYER M1 ;
        RECT 39.2 18.696 39.232 21.204 ;
  LAYER M3 ;
        RECT 39.2 18.716 39.232 18.748 ;
  LAYER M1 ;
        RECT 39.264 18.696 39.296 21.204 ;
  LAYER M3 ;
        RECT 39.264 21.152 39.296 21.184 ;
  LAYER M1 ;
        RECT 39.328 18.696 39.36 21.204 ;
  LAYER M3 ;
        RECT 39.328 18.716 39.36 18.748 ;
  LAYER M1 ;
        RECT 39.392 18.696 39.424 21.204 ;
  LAYER M3 ;
        RECT 39.392 21.152 39.424 21.184 ;
  LAYER M1 ;
        RECT 39.456 18.696 39.488 21.204 ;
  LAYER M3 ;
        RECT 39.456 18.716 39.488 18.748 ;
  LAYER M1 ;
        RECT 39.52 18.696 39.552 21.204 ;
  LAYER M3 ;
        RECT 39.52 21.152 39.552 21.184 ;
  LAYER M1 ;
        RECT 39.584 18.696 39.616 21.204 ;
  LAYER M3 ;
        RECT 39.584 18.716 39.616 18.748 ;
  LAYER M1 ;
        RECT 39.648 18.696 39.68 21.204 ;
  LAYER M3 ;
        RECT 39.648 21.152 39.68 21.184 ;
  LAYER M1 ;
        RECT 39.712 18.696 39.744 21.204 ;
  LAYER M3 ;
        RECT 39.712 18.716 39.744 18.748 ;
  LAYER M1 ;
        RECT 39.776 18.696 39.808 21.204 ;
  LAYER M3 ;
        RECT 39.776 21.152 39.808 21.184 ;
  LAYER M1 ;
        RECT 39.84 18.696 39.872 21.204 ;
  LAYER M3 ;
        RECT 39.84 18.716 39.872 18.748 ;
  LAYER M1 ;
        RECT 39.904 18.696 39.936 21.204 ;
  LAYER M3 ;
        RECT 39.904 21.152 39.936 21.184 ;
  LAYER M1 ;
        RECT 39.968 18.696 40 21.204 ;
  LAYER M3 ;
        RECT 39.968 18.716 40 18.748 ;
  LAYER M1 ;
        RECT 40.032 18.696 40.064 21.204 ;
  LAYER M3 ;
        RECT 40.032 21.152 40.064 21.184 ;
  LAYER M1 ;
        RECT 40.096 18.696 40.128 21.204 ;
  LAYER M3 ;
        RECT 40.096 18.716 40.128 18.748 ;
  LAYER M1 ;
        RECT 40.16 18.696 40.192 21.204 ;
  LAYER M3 ;
        RECT 40.16 21.152 40.192 21.184 ;
  LAYER M1 ;
        RECT 40.224 18.696 40.256 21.204 ;
  LAYER M3 ;
        RECT 40.224 18.716 40.256 18.748 ;
  LAYER M1 ;
        RECT 40.288 18.696 40.32 21.204 ;
  LAYER M3 ;
        RECT 40.288 21.152 40.32 21.184 ;
  LAYER M1 ;
        RECT 40.352 18.696 40.384 21.204 ;
  LAYER M3 ;
        RECT 40.352 18.716 40.384 18.748 ;
  LAYER M1 ;
        RECT 40.416 18.696 40.448 21.204 ;
  LAYER M3 ;
        RECT 40.416 21.152 40.448 21.184 ;
  LAYER M1 ;
        RECT 40.48 18.696 40.512 21.204 ;
  LAYER M3 ;
        RECT 40.48 18.716 40.512 18.748 ;
  LAYER M1 ;
        RECT 40.544 18.696 40.576 21.204 ;
  LAYER M3 ;
        RECT 40.544 21.152 40.576 21.184 ;
  LAYER M1 ;
        RECT 40.608 18.696 40.64 21.204 ;
  LAYER M3 ;
        RECT 40.608 18.716 40.64 18.748 ;
  LAYER M1 ;
        RECT 40.672 18.696 40.704 21.204 ;
  LAYER M3 ;
        RECT 40.672 21.152 40.704 21.184 ;
  LAYER M1 ;
        RECT 40.736 18.696 40.768 21.204 ;
  LAYER M3 ;
        RECT 40.736 18.716 40.768 18.748 ;
  LAYER M1 ;
        RECT 40.8 18.696 40.832 21.204 ;
  LAYER M3 ;
        RECT 40.8 21.152 40.832 21.184 ;
  LAYER M1 ;
        RECT 40.864 18.696 40.896 21.204 ;
  LAYER M3 ;
        RECT 40.864 18.716 40.896 18.748 ;
  LAYER M1 ;
        RECT 40.928 18.696 40.96 21.204 ;
  LAYER M3 ;
        RECT 38.56 21.088 38.592 21.12 ;
  LAYER M2 ;
        RECT 40.928 21.024 40.96 21.056 ;
  LAYER M2 ;
        RECT 38.56 20.96 38.592 20.992 ;
  LAYER M2 ;
        RECT 40.928 20.896 40.96 20.928 ;
  LAYER M2 ;
        RECT 38.56 20.832 38.592 20.864 ;
  LAYER M2 ;
        RECT 40.928 20.768 40.96 20.8 ;
  LAYER M2 ;
        RECT 38.56 20.704 38.592 20.736 ;
  LAYER M2 ;
        RECT 40.928 20.64 40.96 20.672 ;
  LAYER M2 ;
        RECT 38.56 20.576 38.592 20.608 ;
  LAYER M2 ;
        RECT 40.928 20.512 40.96 20.544 ;
  LAYER M2 ;
        RECT 38.56 20.448 38.592 20.48 ;
  LAYER M2 ;
        RECT 40.928 20.384 40.96 20.416 ;
  LAYER M2 ;
        RECT 38.56 20.32 38.592 20.352 ;
  LAYER M2 ;
        RECT 40.928 20.256 40.96 20.288 ;
  LAYER M2 ;
        RECT 38.56 20.192 38.592 20.224 ;
  LAYER M2 ;
        RECT 40.928 20.128 40.96 20.16 ;
  LAYER M2 ;
        RECT 38.56 20.064 38.592 20.096 ;
  LAYER M2 ;
        RECT 40.928 20 40.96 20.032 ;
  LAYER M2 ;
        RECT 38.56 19.936 38.592 19.968 ;
  LAYER M2 ;
        RECT 40.928 19.872 40.96 19.904 ;
  LAYER M2 ;
        RECT 38.56 19.808 38.592 19.84 ;
  LAYER M2 ;
        RECT 40.928 19.744 40.96 19.776 ;
  LAYER M2 ;
        RECT 38.56 19.68 38.592 19.712 ;
  LAYER M2 ;
        RECT 40.928 19.616 40.96 19.648 ;
  LAYER M2 ;
        RECT 38.56 19.552 38.592 19.584 ;
  LAYER M2 ;
        RECT 40.928 19.488 40.96 19.52 ;
  LAYER M2 ;
        RECT 38.56 19.424 38.592 19.456 ;
  LAYER M2 ;
        RECT 40.928 19.36 40.96 19.392 ;
  LAYER M2 ;
        RECT 38.56 19.296 38.592 19.328 ;
  LAYER M2 ;
        RECT 40.928 19.232 40.96 19.264 ;
  LAYER M2 ;
        RECT 38.56 19.168 38.592 19.2 ;
  LAYER M2 ;
        RECT 40.928 19.104 40.96 19.136 ;
  LAYER M2 ;
        RECT 38.56 19.04 38.592 19.072 ;
  LAYER M2 ;
        RECT 40.928 18.976 40.96 19.008 ;
  LAYER M2 ;
        RECT 38.56 18.912 38.592 18.944 ;
  LAYER M2 ;
        RECT 40.928 18.848 40.96 18.88 ;
  LAYER M2 ;
        RECT 38.512 18.648 41.008 21.252 ;
  LAYER M1 ;
        RECT 38.56 15.588 38.592 18.096 ;
  LAYER M3 ;
        RECT 38.56 15.608 38.592 15.64 ;
  LAYER M1 ;
        RECT 38.624 15.588 38.656 18.096 ;
  LAYER M3 ;
        RECT 38.624 18.044 38.656 18.076 ;
  LAYER M1 ;
        RECT 38.688 15.588 38.72 18.096 ;
  LAYER M3 ;
        RECT 38.688 15.608 38.72 15.64 ;
  LAYER M1 ;
        RECT 38.752 15.588 38.784 18.096 ;
  LAYER M3 ;
        RECT 38.752 18.044 38.784 18.076 ;
  LAYER M1 ;
        RECT 38.816 15.588 38.848 18.096 ;
  LAYER M3 ;
        RECT 38.816 15.608 38.848 15.64 ;
  LAYER M1 ;
        RECT 38.88 15.588 38.912 18.096 ;
  LAYER M3 ;
        RECT 38.88 18.044 38.912 18.076 ;
  LAYER M1 ;
        RECT 38.944 15.588 38.976 18.096 ;
  LAYER M3 ;
        RECT 38.944 15.608 38.976 15.64 ;
  LAYER M1 ;
        RECT 39.008 15.588 39.04 18.096 ;
  LAYER M3 ;
        RECT 39.008 18.044 39.04 18.076 ;
  LAYER M1 ;
        RECT 39.072 15.588 39.104 18.096 ;
  LAYER M3 ;
        RECT 39.072 15.608 39.104 15.64 ;
  LAYER M1 ;
        RECT 39.136 15.588 39.168 18.096 ;
  LAYER M3 ;
        RECT 39.136 18.044 39.168 18.076 ;
  LAYER M1 ;
        RECT 39.2 15.588 39.232 18.096 ;
  LAYER M3 ;
        RECT 39.2 15.608 39.232 15.64 ;
  LAYER M1 ;
        RECT 39.264 15.588 39.296 18.096 ;
  LAYER M3 ;
        RECT 39.264 18.044 39.296 18.076 ;
  LAYER M1 ;
        RECT 39.328 15.588 39.36 18.096 ;
  LAYER M3 ;
        RECT 39.328 15.608 39.36 15.64 ;
  LAYER M1 ;
        RECT 39.392 15.588 39.424 18.096 ;
  LAYER M3 ;
        RECT 39.392 18.044 39.424 18.076 ;
  LAYER M1 ;
        RECT 39.456 15.588 39.488 18.096 ;
  LAYER M3 ;
        RECT 39.456 15.608 39.488 15.64 ;
  LAYER M1 ;
        RECT 39.52 15.588 39.552 18.096 ;
  LAYER M3 ;
        RECT 39.52 18.044 39.552 18.076 ;
  LAYER M1 ;
        RECT 39.584 15.588 39.616 18.096 ;
  LAYER M3 ;
        RECT 39.584 15.608 39.616 15.64 ;
  LAYER M1 ;
        RECT 39.648 15.588 39.68 18.096 ;
  LAYER M3 ;
        RECT 39.648 18.044 39.68 18.076 ;
  LAYER M1 ;
        RECT 39.712 15.588 39.744 18.096 ;
  LAYER M3 ;
        RECT 39.712 15.608 39.744 15.64 ;
  LAYER M1 ;
        RECT 39.776 15.588 39.808 18.096 ;
  LAYER M3 ;
        RECT 39.776 18.044 39.808 18.076 ;
  LAYER M1 ;
        RECT 39.84 15.588 39.872 18.096 ;
  LAYER M3 ;
        RECT 39.84 15.608 39.872 15.64 ;
  LAYER M1 ;
        RECT 39.904 15.588 39.936 18.096 ;
  LAYER M3 ;
        RECT 39.904 18.044 39.936 18.076 ;
  LAYER M1 ;
        RECT 39.968 15.588 40 18.096 ;
  LAYER M3 ;
        RECT 39.968 15.608 40 15.64 ;
  LAYER M1 ;
        RECT 40.032 15.588 40.064 18.096 ;
  LAYER M3 ;
        RECT 40.032 18.044 40.064 18.076 ;
  LAYER M1 ;
        RECT 40.096 15.588 40.128 18.096 ;
  LAYER M3 ;
        RECT 40.096 15.608 40.128 15.64 ;
  LAYER M1 ;
        RECT 40.16 15.588 40.192 18.096 ;
  LAYER M3 ;
        RECT 40.16 18.044 40.192 18.076 ;
  LAYER M1 ;
        RECT 40.224 15.588 40.256 18.096 ;
  LAYER M3 ;
        RECT 40.224 15.608 40.256 15.64 ;
  LAYER M1 ;
        RECT 40.288 15.588 40.32 18.096 ;
  LAYER M3 ;
        RECT 40.288 18.044 40.32 18.076 ;
  LAYER M1 ;
        RECT 40.352 15.588 40.384 18.096 ;
  LAYER M3 ;
        RECT 40.352 15.608 40.384 15.64 ;
  LAYER M1 ;
        RECT 40.416 15.588 40.448 18.096 ;
  LAYER M3 ;
        RECT 40.416 18.044 40.448 18.076 ;
  LAYER M1 ;
        RECT 40.48 15.588 40.512 18.096 ;
  LAYER M3 ;
        RECT 40.48 15.608 40.512 15.64 ;
  LAYER M1 ;
        RECT 40.544 15.588 40.576 18.096 ;
  LAYER M3 ;
        RECT 40.544 18.044 40.576 18.076 ;
  LAYER M1 ;
        RECT 40.608 15.588 40.64 18.096 ;
  LAYER M3 ;
        RECT 40.608 15.608 40.64 15.64 ;
  LAYER M1 ;
        RECT 40.672 15.588 40.704 18.096 ;
  LAYER M3 ;
        RECT 40.672 18.044 40.704 18.076 ;
  LAYER M1 ;
        RECT 40.736 15.588 40.768 18.096 ;
  LAYER M3 ;
        RECT 40.736 15.608 40.768 15.64 ;
  LAYER M1 ;
        RECT 40.8 15.588 40.832 18.096 ;
  LAYER M3 ;
        RECT 40.8 18.044 40.832 18.076 ;
  LAYER M1 ;
        RECT 40.864 15.588 40.896 18.096 ;
  LAYER M3 ;
        RECT 40.864 15.608 40.896 15.64 ;
  LAYER M1 ;
        RECT 40.928 15.588 40.96 18.096 ;
  LAYER M3 ;
        RECT 38.56 17.98 38.592 18.012 ;
  LAYER M2 ;
        RECT 40.928 17.916 40.96 17.948 ;
  LAYER M2 ;
        RECT 38.56 17.852 38.592 17.884 ;
  LAYER M2 ;
        RECT 40.928 17.788 40.96 17.82 ;
  LAYER M2 ;
        RECT 38.56 17.724 38.592 17.756 ;
  LAYER M2 ;
        RECT 40.928 17.66 40.96 17.692 ;
  LAYER M2 ;
        RECT 38.56 17.596 38.592 17.628 ;
  LAYER M2 ;
        RECT 40.928 17.532 40.96 17.564 ;
  LAYER M2 ;
        RECT 38.56 17.468 38.592 17.5 ;
  LAYER M2 ;
        RECT 40.928 17.404 40.96 17.436 ;
  LAYER M2 ;
        RECT 38.56 17.34 38.592 17.372 ;
  LAYER M2 ;
        RECT 40.928 17.276 40.96 17.308 ;
  LAYER M2 ;
        RECT 38.56 17.212 38.592 17.244 ;
  LAYER M2 ;
        RECT 40.928 17.148 40.96 17.18 ;
  LAYER M2 ;
        RECT 38.56 17.084 38.592 17.116 ;
  LAYER M2 ;
        RECT 40.928 17.02 40.96 17.052 ;
  LAYER M2 ;
        RECT 38.56 16.956 38.592 16.988 ;
  LAYER M2 ;
        RECT 40.928 16.892 40.96 16.924 ;
  LAYER M2 ;
        RECT 38.56 16.828 38.592 16.86 ;
  LAYER M2 ;
        RECT 40.928 16.764 40.96 16.796 ;
  LAYER M2 ;
        RECT 38.56 16.7 38.592 16.732 ;
  LAYER M2 ;
        RECT 40.928 16.636 40.96 16.668 ;
  LAYER M2 ;
        RECT 38.56 16.572 38.592 16.604 ;
  LAYER M2 ;
        RECT 40.928 16.508 40.96 16.54 ;
  LAYER M2 ;
        RECT 38.56 16.444 38.592 16.476 ;
  LAYER M2 ;
        RECT 40.928 16.38 40.96 16.412 ;
  LAYER M2 ;
        RECT 38.56 16.316 38.592 16.348 ;
  LAYER M2 ;
        RECT 40.928 16.252 40.96 16.284 ;
  LAYER M2 ;
        RECT 38.56 16.188 38.592 16.22 ;
  LAYER M2 ;
        RECT 40.928 16.124 40.96 16.156 ;
  LAYER M2 ;
        RECT 38.56 16.06 38.592 16.092 ;
  LAYER M2 ;
        RECT 40.928 15.996 40.96 16.028 ;
  LAYER M2 ;
        RECT 38.56 15.932 38.592 15.964 ;
  LAYER M2 ;
        RECT 40.928 15.868 40.96 15.9 ;
  LAYER M2 ;
        RECT 38.56 15.804 38.592 15.836 ;
  LAYER M2 ;
        RECT 40.928 15.74 40.96 15.772 ;
  LAYER M2 ;
        RECT 38.512 15.54 41.008 18.144 ;
  LAYER M1 ;
        RECT 41.536 28.02 41.568 30.528 ;
  LAYER M3 ;
        RECT 41.536 28.04 41.568 28.072 ;
  LAYER M1 ;
        RECT 41.6 28.02 41.632 30.528 ;
  LAYER M3 ;
        RECT 41.6 30.476 41.632 30.508 ;
  LAYER M1 ;
        RECT 41.664 28.02 41.696 30.528 ;
  LAYER M3 ;
        RECT 41.664 28.04 41.696 28.072 ;
  LAYER M1 ;
        RECT 41.728 28.02 41.76 30.528 ;
  LAYER M3 ;
        RECT 41.728 30.476 41.76 30.508 ;
  LAYER M1 ;
        RECT 41.792 28.02 41.824 30.528 ;
  LAYER M3 ;
        RECT 41.792 28.04 41.824 28.072 ;
  LAYER M1 ;
        RECT 41.856 28.02 41.888 30.528 ;
  LAYER M3 ;
        RECT 41.856 30.476 41.888 30.508 ;
  LAYER M1 ;
        RECT 41.92 28.02 41.952 30.528 ;
  LAYER M3 ;
        RECT 41.92 28.04 41.952 28.072 ;
  LAYER M1 ;
        RECT 41.984 28.02 42.016 30.528 ;
  LAYER M3 ;
        RECT 41.984 30.476 42.016 30.508 ;
  LAYER M1 ;
        RECT 42.048 28.02 42.08 30.528 ;
  LAYER M3 ;
        RECT 42.048 28.04 42.08 28.072 ;
  LAYER M1 ;
        RECT 42.112 28.02 42.144 30.528 ;
  LAYER M3 ;
        RECT 42.112 30.476 42.144 30.508 ;
  LAYER M1 ;
        RECT 42.176 28.02 42.208 30.528 ;
  LAYER M3 ;
        RECT 42.176 28.04 42.208 28.072 ;
  LAYER M1 ;
        RECT 42.24 28.02 42.272 30.528 ;
  LAYER M3 ;
        RECT 42.24 30.476 42.272 30.508 ;
  LAYER M1 ;
        RECT 42.304 28.02 42.336 30.528 ;
  LAYER M3 ;
        RECT 42.304 28.04 42.336 28.072 ;
  LAYER M1 ;
        RECT 42.368 28.02 42.4 30.528 ;
  LAYER M3 ;
        RECT 42.368 30.476 42.4 30.508 ;
  LAYER M1 ;
        RECT 42.432 28.02 42.464 30.528 ;
  LAYER M3 ;
        RECT 42.432 28.04 42.464 28.072 ;
  LAYER M1 ;
        RECT 42.496 28.02 42.528 30.528 ;
  LAYER M3 ;
        RECT 42.496 30.476 42.528 30.508 ;
  LAYER M1 ;
        RECT 42.56 28.02 42.592 30.528 ;
  LAYER M3 ;
        RECT 42.56 28.04 42.592 28.072 ;
  LAYER M1 ;
        RECT 42.624 28.02 42.656 30.528 ;
  LAYER M3 ;
        RECT 42.624 30.476 42.656 30.508 ;
  LAYER M1 ;
        RECT 42.688 28.02 42.72 30.528 ;
  LAYER M3 ;
        RECT 42.688 28.04 42.72 28.072 ;
  LAYER M1 ;
        RECT 42.752 28.02 42.784 30.528 ;
  LAYER M3 ;
        RECT 42.752 30.476 42.784 30.508 ;
  LAYER M1 ;
        RECT 42.816 28.02 42.848 30.528 ;
  LAYER M3 ;
        RECT 42.816 28.04 42.848 28.072 ;
  LAYER M1 ;
        RECT 42.88 28.02 42.912 30.528 ;
  LAYER M3 ;
        RECT 42.88 30.476 42.912 30.508 ;
  LAYER M1 ;
        RECT 42.944 28.02 42.976 30.528 ;
  LAYER M3 ;
        RECT 42.944 28.04 42.976 28.072 ;
  LAYER M1 ;
        RECT 43.008 28.02 43.04 30.528 ;
  LAYER M3 ;
        RECT 43.008 30.476 43.04 30.508 ;
  LAYER M1 ;
        RECT 43.072 28.02 43.104 30.528 ;
  LAYER M3 ;
        RECT 43.072 28.04 43.104 28.072 ;
  LAYER M1 ;
        RECT 43.136 28.02 43.168 30.528 ;
  LAYER M3 ;
        RECT 43.136 30.476 43.168 30.508 ;
  LAYER M1 ;
        RECT 43.2 28.02 43.232 30.528 ;
  LAYER M3 ;
        RECT 43.2 28.04 43.232 28.072 ;
  LAYER M1 ;
        RECT 43.264 28.02 43.296 30.528 ;
  LAYER M3 ;
        RECT 43.264 30.476 43.296 30.508 ;
  LAYER M1 ;
        RECT 43.328 28.02 43.36 30.528 ;
  LAYER M3 ;
        RECT 43.328 28.04 43.36 28.072 ;
  LAYER M1 ;
        RECT 43.392 28.02 43.424 30.528 ;
  LAYER M3 ;
        RECT 43.392 30.476 43.424 30.508 ;
  LAYER M1 ;
        RECT 43.456 28.02 43.488 30.528 ;
  LAYER M3 ;
        RECT 43.456 28.04 43.488 28.072 ;
  LAYER M1 ;
        RECT 43.52 28.02 43.552 30.528 ;
  LAYER M3 ;
        RECT 43.52 30.476 43.552 30.508 ;
  LAYER M1 ;
        RECT 43.584 28.02 43.616 30.528 ;
  LAYER M3 ;
        RECT 43.584 28.04 43.616 28.072 ;
  LAYER M1 ;
        RECT 43.648 28.02 43.68 30.528 ;
  LAYER M3 ;
        RECT 43.648 30.476 43.68 30.508 ;
  LAYER M1 ;
        RECT 43.712 28.02 43.744 30.528 ;
  LAYER M3 ;
        RECT 43.712 28.04 43.744 28.072 ;
  LAYER M1 ;
        RECT 43.776 28.02 43.808 30.528 ;
  LAYER M3 ;
        RECT 43.776 30.476 43.808 30.508 ;
  LAYER M1 ;
        RECT 43.84 28.02 43.872 30.528 ;
  LAYER M3 ;
        RECT 43.84 28.04 43.872 28.072 ;
  LAYER M1 ;
        RECT 43.904 28.02 43.936 30.528 ;
  LAYER M3 ;
        RECT 41.536 30.412 41.568 30.444 ;
  LAYER M2 ;
        RECT 43.904 30.348 43.936 30.38 ;
  LAYER M2 ;
        RECT 41.536 30.284 41.568 30.316 ;
  LAYER M2 ;
        RECT 43.904 30.22 43.936 30.252 ;
  LAYER M2 ;
        RECT 41.536 30.156 41.568 30.188 ;
  LAYER M2 ;
        RECT 43.904 30.092 43.936 30.124 ;
  LAYER M2 ;
        RECT 41.536 30.028 41.568 30.06 ;
  LAYER M2 ;
        RECT 43.904 29.964 43.936 29.996 ;
  LAYER M2 ;
        RECT 41.536 29.9 41.568 29.932 ;
  LAYER M2 ;
        RECT 43.904 29.836 43.936 29.868 ;
  LAYER M2 ;
        RECT 41.536 29.772 41.568 29.804 ;
  LAYER M2 ;
        RECT 43.904 29.708 43.936 29.74 ;
  LAYER M2 ;
        RECT 41.536 29.644 41.568 29.676 ;
  LAYER M2 ;
        RECT 43.904 29.58 43.936 29.612 ;
  LAYER M2 ;
        RECT 41.536 29.516 41.568 29.548 ;
  LAYER M2 ;
        RECT 43.904 29.452 43.936 29.484 ;
  LAYER M2 ;
        RECT 41.536 29.388 41.568 29.42 ;
  LAYER M2 ;
        RECT 43.904 29.324 43.936 29.356 ;
  LAYER M2 ;
        RECT 41.536 29.26 41.568 29.292 ;
  LAYER M2 ;
        RECT 43.904 29.196 43.936 29.228 ;
  LAYER M2 ;
        RECT 41.536 29.132 41.568 29.164 ;
  LAYER M2 ;
        RECT 43.904 29.068 43.936 29.1 ;
  LAYER M2 ;
        RECT 41.536 29.004 41.568 29.036 ;
  LAYER M2 ;
        RECT 43.904 28.94 43.936 28.972 ;
  LAYER M2 ;
        RECT 41.536 28.876 41.568 28.908 ;
  LAYER M2 ;
        RECT 43.904 28.812 43.936 28.844 ;
  LAYER M2 ;
        RECT 41.536 28.748 41.568 28.78 ;
  LAYER M2 ;
        RECT 43.904 28.684 43.936 28.716 ;
  LAYER M2 ;
        RECT 41.536 28.62 41.568 28.652 ;
  LAYER M2 ;
        RECT 43.904 28.556 43.936 28.588 ;
  LAYER M2 ;
        RECT 41.536 28.492 41.568 28.524 ;
  LAYER M2 ;
        RECT 43.904 28.428 43.936 28.46 ;
  LAYER M2 ;
        RECT 41.536 28.364 41.568 28.396 ;
  LAYER M2 ;
        RECT 43.904 28.3 43.936 28.332 ;
  LAYER M2 ;
        RECT 41.536 28.236 41.568 28.268 ;
  LAYER M2 ;
        RECT 43.904 28.172 43.936 28.204 ;
  LAYER M2 ;
        RECT 41.488 27.972 43.984 30.576 ;
  LAYER M1 ;
        RECT 41.536 24.912 41.568 27.42 ;
  LAYER M3 ;
        RECT 41.536 24.932 41.568 24.964 ;
  LAYER M1 ;
        RECT 41.6 24.912 41.632 27.42 ;
  LAYER M3 ;
        RECT 41.6 27.368 41.632 27.4 ;
  LAYER M1 ;
        RECT 41.664 24.912 41.696 27.42 ;
  LAYER M3 ;
        RECT 41.664 24.932 41.696 24.964 ;
  LAYER M1 ;
        RECT 41.728 24.912 41.76 27.42 ;
  LAYER M3 ;
        RECT 41.728 27.368 41.76 27.4 ;
  LAYER M1 ;
        RECT 41.792 24.912 41.824 27.42 ;
  LAYER M3 ;
        RECT 41.792 24.932 41.824 24.964 ;
  LAYER M1 ;
        RECT 41.856 24.912 41.888 27.42 ;
  LAYER M3 ;
        RECT 41.856 27.368 41.888 27.4 ;
  LAYER M1 ;
        RECT 41.92 24.912 41.952 27.42 ;
  LAYER M3 ;
        RECT 41.92 24.932 41.952 24.964 ;
  LAYER M1 ;
        RECT 41.984 24.912 42.016 27.42 ;
  LAYER M3 ;
        RECT 41.984 27.368 42.016 27.4 ;
  LAYER M1 ;
        RECT 42.048 24.912 42.08 27.42 ;
  LAYER M3 ;
        RECT 42.048 24.932 42.08 24.964 ;
  LAYER M1 ;
        RECT 42.112 24.912 42.144 27.42 ;
  LAYER M3 ;
        RECT 42.112 27.368 42.144 27.4 ;
  LAYER M1 ;
        RECT 42.176 24.912 42.208 27.42 ;
  LAYER M3 ;
        RECT 42.176 24.932 42.208 24.964 ;
  LAYER M1 ;
        RECT 42.24 24.912 42.272 27.42 ;
  LAYER M3 ;
        RECT 42.24 27.368 42.272 27.4 ;
  LAYER M1 ;
        RECT 42.304 24.912 42.336 27.42 ;
  LAYER M3 ;
        RECT 42.304 24.932 42.336 24.964 ;
  LAYER M1 ;
        RECT 42.368 24.912 42.4 27.42 ;
  LAYER M3 ;
        RECT 42.368 27.368 42.4 27.4 ;
  LAYER M1 ;
        RECT 42.432 24.912 42.464 27.42 ;
  LAYER M3 ;
        RECT 42.432 24.932 42.464 24.964 ;
  LAYER M1 ;
        RECT 42.496 24.912 42.528 27.42 ;
  LAYER M3 ;
        RECT 42.496 27.368 42.528 27.4 ;
  LAYER M1 ;
        RECT 42.56 24.912 42.592 27.42 ;
  LAYER M3 ;
        RECT 42.56 24.932 42.592 24.964 ;
  LAYER M1 ;
        RECT 42.624 24.912 42.656 27.42 ;
  LAYER M3 ;
        RECT 42.624 27.368 42.656 27.4 ;
  LAYER M1 ;
        RECT 42.688 24.912 42.72 27.42 ;
  LAYER M3 ;
        RECT 42.688 24.932 42.72 24.964 ;
  LAYER M1 ;
        RECT 42.752 24.912 42.784 27.42 ;
  LAYER M3 ;
        RECT 42.752 27.368 42.784 27.4 ;
  LAYER M1 ;
        RECT 42.816 24.912 42.848 27.42 ;
  LAYER M3 ;
        RECT 42.816 24.932 42.848 24.964 ;
  LAYER M1 ;
        RECT 42.88 24.912 42.912 27.42 ;
  LAYER M3 ;
        RECT 42.88 27.368 42.912 27.4 ;
  LAYER M1 ;
        RECT 42.944 24.912 42.976 27.42 ;
  LAYER M3 ;
        RECT 42.944 24.932 42.976 24.964 ;
  LAYER M1 ;
        RECT 43.008 24.912 43.04 27.42 ;
  LAYER M3 ;
        RECT 43.008 27.368 43.04 27.4 ;
  LAYER M1 ;
        RECT 43.072 24.912 43.104 27.42 ;
  LAYER M3 ;
        RECT 43.072 24.932 43.104 24.964 ;
  LAYER M1 ;
        RECT 43.136 24.912 43.168 27.42 ;
  LAYER M3 ;
        RECT 43.136 27.368 43.168 27.4 ;
  LAYER M1 ;
        RECT 43.2 24.912 43.232 27.42 ;
  LAYER M3 ;
        RECT 43.2 24.932 43.232 24.964 ;
  LAYER M1 ;
        RECT 43.264 24.912 43.296 27.42 ;
  LAYER M3 ;
        RECT 43.264 27.368 43.296 27.4 ;
  LAYER M1 ;
        RECT 43.328 24.912 43.36 27.42 ;
  LAYER M3 ;
        RECT 43.328 24.932 43.36 24.964 ;
  LAYER M1 ;
        RECT 43.392 24.912 43.424 27.42 ;
  LAYER M3 ;
        RECT 43.392 27.368 43.424 27.4 ;
  LAYER M1 ;
        RECT 43.456 24.912 43.488 27.42 ;
  LAYER M3 ;
        RECT 43.456 24.932 43.488 24.964 ;
  LAYER M1 ;
        RECT 43.52 24.912 43.552 27.42 ;
  LAYER M3 ;
        RECT 43.52 27.368 43.552 27.4 ;
  LAYER M1 ;
        RECT 43.584 24.912 43.616 27.42 ;
  LAYER M3 ;
        RECT 43.584 24.932 43.616 24.964 ;
  LAYER M1 ;
        RECT 43.648 24.912 43.68 27.42 ;
  LAYER M3 ;
        RECT 43.648 27.368 43.68 27.4 ;
  LAYER M1 ;
        RECT 43.712 24.912 43.744 27.42 ;
  LAYER M3 ;
        RECT 43.712 24.932 43.744 24.964 ;
  LAYER M1 ;
        RECT 43.776 24.912 43.808 27.42 ;
  LAYER M3 ;
        RECT 43.776 27.368 43.808 27.4 ;
  LAYER M1 ;
        RECT 43.84 24.912 43.872 27.42 ;
  LAYER M3 ;
        RECT 43.84 24.932 43.872 24.964 ;
  LAYER M1 ;
        RECT 43.904 24.912 43.936 27.42 ;
  LAYER M3 ;
        RECT 41.536 27.304 41.568 27.336 ;
  LAYER M2 ;
        RECT 43.904 27.24 43.936 27.272 ;
  LAYER M2 ;
        RECT 41.536 27.176 41.568 27.208 ;
  LAYER M2 ;
        RECT 43.904 27.112 43.936 27.144 ;
  LAYER M2 ;
        RECT 41.536 27.048 41.568 27.08 ;
  LAYER M2 ;
        RECT 43.904 26.984 43.936 27.016 ;
  LAYER M2 ;
        RECT 41.536 26.92 41.568 26.952 ;
  LAYER M2 ;
        RECT 43.904 26.856 43.936 26.888 ;
  LAYER M2 ;
        RECT 41.536 26.792 41.568 26.824 ;
  LAYER M2 ;
        RECT 43.904 26.728 43.936 26.76 ;
  LAYER M2 ;
        RECT 41.536 26.664 41.568 26.696 ;
  LAYER M2 ;
        RECT 43.904 26.6 43.936 26.632 ;
  LAYER M2 ;
        RECT 41.536 26.536 41.568 26.568 ;
  LAYER M2 ;
        RECT 43.904 26.472 43.936 26.504 ;
  LAYER M2 ;
        RECT 41.536 26.408 41.568 26.44 ;
  LAYER M2 ;
        RECT 43.904 26.344 43.936 26.376 ;
  LAYER M2 ;
        RECT 41.536 26.28 41.568 26.312 ;
  LAYER M2 ;
        RECT 43.904 26.216 43.936 26.248 ;
  LAYER M2 ;
        RECT 41.536 26.152 41.568 26.184 ;
  LAYER M2 ;
        RECT 43.904 26.088 43.936 26.12 ;
  LAYER M2 ;
        RECT 41.536 26.024 41.568 26.056 ;
  LAYER M2 ;
        RECT 43.904 25.96 43.936 25.992 ;
  LAYER M2 ;
        RECT 41.536 25.896 41.568 25.928 ;
  LAYER M2 ;
        RECT 43.904 25.832 43.936 25.864 ;
  LAYER M2 ;
        RECT 41.536 25.768 41.568 25.8 ;
  LAYER M2 ;
        RECT 43.904 25.704 43.936 25.736 ;
  LAYER M2 ;
        RECT 41.536 25.64 41.568 25.672 ;
  LAYER M2 ;
        RECT 43.904 25.576 43.936 25.608 ;
  LAYER M2 ;
        RECT 41.536 25.512 41.568 25.544 ;
  LAYER M2 ;
        RECT 43.904 25.448 43.936 25.48 ;
  LAYER M2 ;
        RECT 41.536 25.384 41.568 25.416 ;
  LAYER M2 ;
        RECT 43.904 25.32 43.936 25.352 ;
  LAYER M2 ;
        RECT 41.536 25.256 41.568 25.288 ;
  LAYER M2 ;
        RECT 43.904 25.192 43.936 25.224 ;
  LAYER M2 ;
        RECT 41.536 25.128 41.568 25.16 ;
  LAYER M2 ;
        RECT 43.904 25.064 43.936 25.096 ;
  LAYER M2 ;
        RECT 41.488 24.864 43.984 27.468 ;
  LAYER M1 ;
        RECT 41.536 21.804 41.568 24.312 ;
  LAYER M3 ;
        RECT 41.536 21.824 41.568 21.856 ;
  LAYER M1 ;
        RECT 41.6 21.804 41.632 24.312 ;
  LAYER M3 ;
        RECT 41.6 24.26 41.632 24.292 ;
  LAYER M1 ;
        RECT 41.664 21.804 41.696 24.312 ;
  LAYER M3 ;
        RECT 41.664 21.824 41.696 21.856 ;
  LAYER M1 ;
        RECT 41.728 21.804 41.76 24.312 ;
  LAYER M3 ;
        RECT 41.728 24.26 41.76 24.292 ;
  LAYER M1 ;
        RECT 41.792 21.804 41.824 24.312 ;
  LAYER M3 ;
        RECT 41.792 21.824 41.824 21.856 ;
  LAYER M1 ;
        RECT 41.856 21.804 41.888 24.312 ;
  LAYER M3 ;
        RECT 41.856 24.26 41.888 24.292 ;
  LAYER M1 ;
        RECT 41.92 21.804 41.952 24.312 ;
  LAYER M3 ;
        RECT 41.92 21.824 41.952 21.856 ;
  LAYER M1 ;
        RECT 41.984 21.804 42.016 24.312 ;
  LAYER M3 ;
        RECT 41.984 24.26 42.016 24.292 ;
  LAYER M1 ;
        RECT 42.048 21.804 42.08 24.312 ;
  LAYER M3 ;
        RECT 42.048 21.824 42.08 21.856 ;
  LAYER M1 ;
        RECT 42.112 21.804 42.144 24.312 ;
  LAYER M3 ;
        RECT 42.112 24.26 42.144 24.292 ;
  LAYER M1 ;
        RECT 42.176 21.804 42.208 24.312 ;
  LAYER M3 ;
        RECT 42.176 21.824 42.208 21.856 ;
  LAYER M1 ;
        RECT 42.24 21.804 42.272 24.312 ;
  LAYER M3 ;
        RECT 42.24 24.26 42.272 24.292 ;
  LAYER M1 ;
        RECT 42.304 21.804 42.336 24.312 ;
  LAYER M3 ;
        RECT 42.304 21.824 42.336 21.856 ;
  LAYER M1 ;
        RECT 42.368 21.804 42.4 24.312 ;
  LAYER M3 ;
        RECT 42.368 24.26 42.4 24.292 ;
  LAYER M1 ;
        RECT 42.432 21.804 42.464 24.312 ;
  LAYER M3 ;
        RECT 42.432 21.824 42.464 21.856 ;
  LAYER M1 ;
        RECT 42.496 21.804 42.528 24.312 ;
  LAYER M3 ;
        RECT 42.496 24.26 42.528 24.292 ;
  LAYER M1 ;
        RECT 42.56 21.804 42.592 24.312 ;
  LAYER M3 ;
        RECT 42.56 21.824 42.592 21.856 ;
  LAYER M1 ;
        RECT 42.624 21.804 42.656 24.312 ;
  LAYER M3 ;
        RECT 42.624 24.26 42.656 24.292 ;
  LAYER M1 ;
        RECT 42.688 21.804 42.72 24.312 ;
  LAYER M3 ;
        RECT 42.688 21.824 42.72 21.856 ;
  LAYER M1 ;
        RECT 42.752 21.804 42.784 24.312 ;
  LAYER M3 ;
        RECT 42.752 24.26 42.784 24.292 ;
  LAYER M1 ;
        RECT 42.816 21.804 42.848 24.312 ;
  LAYER M3 ;
        RECT 42.816 21.824 42.848 21.856 ;
  LAYER M1 ;
        RECT 42.88 21.804 42.912 24.312 ;
  LAYER M3 ;
        RECT 42.88 24.26 42.912 24.292 ;
  LAYER M1 ;
        RECT 42.944 21.804 42.976 24.312 ;
  LAYER M3 ;
        RECT 42.944 21.824 42.976 21.856 ;
  LAYER M1 ;
        RECT 43.008 21.804 43.04 24.312 ;
  LAYER M3 ;
        RECT 43.008 24.26 43.04 24.292 ;
  LAYER M1 ;
        RECT 43.072 21.804 43.104 24.312 ;
  LAYER M3 ;
        RECT 43.072 21.824 43.104 21.856 ;
  LAYER M1 ;
        RECT 43.136 21.804 43.168 24.312 ;
  LAYER M3 ;
        RECT 43.136 24.26 43.168 24.292 ;
  LAYER M1 ;
        RECT 43.2 21.804 43.232 24.312 ;
  LAYER M3 ;
        RECT 43.2 21.824 43.232 21.856 ;
  LAYER M1 ;
        RECT 43.264 21.804 43.296 24.312 ;
  LAYER M3 ;
        RECT 43.264 24.26 43.296 24.292 ;
  LAYER M1 ;
        RECT 43.328 21.804 43.36 24.312 ;
  LAYER M3 ;
        RECT 43.328 21.824 43.36 21.856 ;
  LAYER M1 ;
        RECT 43.392 21.804 43.424 24.312 ;
  LAYER M3 ;
        RECT 43.392 24.26 43.424 24.292 ;
  LAYER M1 ;
        RECT 43.456 21.804 43.488 24.312 ;
  LAYER M3 ;
        RECT 43.456 21.824 43.488 21.856 ;
  LAYER M1 ;
        RECT 43.52 21.804 43.552 24.312 ;
  LAYER M3 ;
        RECT 43.52 24.26 43.552 24.292 ;
  LAYER M1 ;
        RECT 43.584 21.804 43.616 24.312 ;
  LAYER M3 ;
        RECT 43.584 21.824 43.616 21.856 ;
  LAYER M1 ;
        RECT 43.648 21.804 43.68 24.312 ;
  LAYER M3 ;
        RECT 43.648 24.26 43.68 24.292 ;
  LAYER M1 ;
        RECT 43.712 21.804 43.744 24.312 ;
  LAYER M3 ;
        RECT 43.712 21.824 43.744 21.856 ;
  LAYER M1 ;
        RECT 43.776 21.804 43.808 24.312 ;
  LAYER M3 ;
        RECT 43.776 24.26 43.808 24.292 ;
  LAYER M1 ;
        RECT 43.84 21.804 43.872 24.312 ;
  LAYER M3 ;
        RECT 43.84 21.824 43.872 21.856 ;
  LAYER M1 ;
        RECT 43.904 21.804 43.936 24.312 ;
  LAYER M3 ;
        RECT 41.536 24.196 41.568 24.228 ;
  LAYER M2 ;
        RECT 43.904 24.132 43.936 24.164 ;
  LAYER M2 ;
        RECT 41.536 24.068 41.568 24.1 ;
  LAYER M2 ;
        RECT 43.904 24.004 43.936 24.036 ;
  LAYER M2 ;
        RECT 41.536 23.94 41.568 23.972 ;
  LAYER M2 ;
        RECT 43.904 23.876 43.936 23.908 ;
  LAYER M2 ;
        RECT 41.536 23.812 41.568 23.844 ;
  LAYER M2 ;
        RECT 43.904 23.748 43.936 23.78 ;
  LAYER M2 ;
        RECT 41.536 23.684 41.568 23.716 ;
  LAYER M2 ;
        RECT 43.904 23.62 43.936 23.652 ;
  LAYER M2 ;
        RECT 41.536 23.556 41.568 23.588 ;
  LAYER M2 ;
        RECT 43.904 23.492 43.936 23.524 ;
  LAYER M2 ;
        RECT 41.536 23.428 41.568 23.46 ;
  LAYER M2 ;
        RECT 43.904 23.364 43.936 23.396 ;
  LAYER M2 ;
        RECT 41.536 23.3 41.568 23.332 ;
  LAYER M2 ;
        RECT 43.904 23.236 43.936 23.268 ;
  LAYER M2 ;
        RECT 41.536 23.172 41.568 23.204 ;
  LAYER M2 ;
        RECT 43.904 23.108 43.936 23.14 ;
  LAYER M2 ;
        RECT 41.536 23.044 41.568 23.076 ;
  LAYER M2 ;
        RECT 43.904 22.98 43.936 23.012 ;
  LAYER M2 ;
        RECT 41.536 22.916 41.568 22.948 ;
  LAYER M2 ;
        RECT 43.904 22.852 43.936 22.884 ;
  LAYER M2 ;
        RECT 41.536 22.788 41.568 22.82 ;
  LAYER M2 ;
        RECT 43.904 22.724 43.936 22.756 ;
  LAYER M2 ;
        RECT 41.536 22.66 41.568 22.692 ;
  LAYER M2 ;
        RECT 43.904 22.596 43.936 22.628 ;
  LAYER M2 ;
        RECT 41.536 22.532 41.568 22.564 ;
  LAYER M2 ;
        RECT 43.904 22.468 43.936 22.5 ;
  LAYER M2 ;
        RECT 41.536 22.404 41.568 22.436 ;
  LAYER M2 ;
        RECT 43.904 22.34 43.936 22.372 ;
  LAYER M2 ;
        RECT 41.536 22.276 41.568 22.308 ;
  LAYER M2 ;
        RECT 43.904 22.212 43.936 22.244 ;
  LAYER M2 ;
        RECT 41.536 22.148 41.568 22.18 ;
  LAYER M2 ;
        RECT 43.904 22.084 43.936 22.116 ;
  LAYER M2 ;
        RECT 41.536 22.02 41.568 22.052 ;
  LAYER M2 ;
        RECT 43.904 21.956 43.936 21.988 ;
  LAYER M2 ;
        RECT 41.488 21.756 43.984 24.36 ;
  LAYER M1 ;
        RECT 41.536 18.696 41.568 21.204 ;
  LAYER M3 ;
        RECT 41.536 18.716 41.568 18.748 ;
  LAYER M1 ;
        RECT 41.6 18.696 41.632 21.204 ;
  LAYER M3 ;
        RECT 41.6 21.152 41.632 21.184 ;
  LAYER M1 ;
        RECT 41.664 18.696 41.696 21.204 ;
  LAYER M3 ;
        RECT 41.664 18.716 41.696 18.748 ;
  LAYER M1 ;
        RECT 41.728 18.696 41.76 21.204 ;
  LAYER M3 ;
        RECT 41.728 21.152 41.76 21.184 ;
  LAYER M1 ;
        RECT 41.792 18.696 41.824 21.204 ;
  LAYER M3 ;
        RECT 41.792 18.716 41.824 18.748 ;
  LAYER M1 ;
        RECT 41.856 18.696 41.888 21.204 ;
  LAYER M3 ;
        RECT 41.856 21.152 41.888 21.184 ;
  LAYER M1 ;
        RECT 41.92 18.696 41.952 21.204 ;
  LAYER M3 ;
        RECT 41.92 18.716 41.952 18.748 ;
  LAYER M1 ;
        RECT 41.984 18.696 42.016 21.204 ;
  LAYER M3 ;
        RECT 41.984 21.152 42.016 21.184 ;
  LAYER M1 ;
        RECT 42.048 18.696 42.08 21.204 ;
  LAYER M3 ;
        RECT 42.048 18.716 42.08 18.748 ;
  LAYER M1 ;
        RECT 42.112 18.696 42.144 21.204 ;
  LAYER M3 ;
        RECT 42.112 21.152 42.144 21.184 ;
  LAYER M1 ;
        RECT 42.176 18.696 42.208 21.204 ;
  LAYER M3 ;
        RECT 42.176 18.716 42.208 18.748 ;
  LAYER M1 ;
        RECT 42.24 18.696 42.272 21.204 ;
  LAYER M3 ;
        RECT 42.24 21.152 42.272 21.184 ;
  LAYER M1 ;
        RECT 42.304 18.696 42.336 21.204 ;
  LAYER M3 ;
        RECT 42.304 18.716 42.336 18.748 ;
  LAYER M1 ;
        RECT 42.368 18.696 42.4 21.204 ;
  LAYER M3 ;
        RECT 42.368 21.152 42.4 21.184 ;
  LAYER M1 ;
        RECT 42.432 18.696 42.464 21.204 ;
  LAYER M3 ;
        RECT 42.432 18.716 42.464 18.748 ;
  LAYER M1 ;
        RECT 42.496 18.696 42.528 21.204 ;
  LAYER M3 ;
        RECT 42.496 21.152 42.528 21.184 ;
  LAYER M1 ;
        RECT 42.56 18.696 42.592 21.204 ;
  LAYER M3 ;
        RECT 42.56 18.716 42.592 18.748 ;
  LAYER M1 ;
        RECT 42.624 18.696 42.656 21.204 ;
  LAYER M3 ;
        RECT 42.624 21.152 42.656 21.184 ;
  LAYER M1 ;
        RECT 42.688 18.696 42.72 21.204 ;
  LAYER M3 ;
        RECT 42.688 18.716 42.72 18.748 ;
  LAYER M1 ;
        RECT 42.752 18.696 42.784 21.204 ;
  LAYER M3 ;
        RECT 42.752 21.152 42.784 21.184 ;
  LAYER M1 ;
        RECT 42.816 18.696 42.848 21.204 ;
  LAYER M3 ;
        RECT 42.816 18.716 42.848 18.748 ;
  LAYER M1 ;
        RECT 42.88 18.696 42.912 21.204 ;
  LAYER M3 ;
        RECT 42.88 21.152 42.912 21.184 ;
  LAYER M1 ;
        RECT 42.944 18.696 42.976 21.204 ;
  LAYER M3 ;
        RECT 42.944 18.716 42.976 18.748 ;
  LAYER M1 ;
        RECT 43.008 18.696 43.04 21.204 ;
  LAYER M3 ;
        RECT 43.008 21.152 43.04 21.184 ;
  LAYER M1 ;
        RECT 43.072 18.696 43.104 21.204 ;
  LAYER M3 ;
        RECT 43.072 18.716 43.104 18.748 ;
  LAYER M1 ;
        RECT 43.136 18.696 43.168 21.204 ;
  LAYER M3 ;
        RECT 43.136 21.152 43.168 21.184 ;
  LAYER M1 ;
        RECT 43.2 18.696 43.232 21.204 ;
  LAYER M3 ;
        RECT 43.2 18.716 43.232 18.748 ;
  LAYER M1 ;
        RECT 43.264 18.696 43.296 21.204 ;
  LAYER M3 ;
        RECT 43.264 21.152 43.296 21.184 ;
  LAYER M1 ;
        RECT 43.328 18.696 43.36 21.204 ;
  LAYER M3 ;
        RECT 43.328 18.716 43.36 18.748 ;
  LAYER M1 ;
        RECT 43.392 18.696 43.424 21.204 ;
  LAYER M3 ;
        RECT 43.392 21.152 43.424 21.184 ;
  LAYER M1 ;
        RECT 43.456 18.696 43.488 21.204 ;
  LAYER M3 ;
        RECT 43.456 18.716 43.488 18.748 ;
  LAYER M1 ;
        RECT 43.52 18.696 43.552 21.204 ;
  LAYER M3 ;
        RECT 43.52 21.152 43.552 21.184 ;
  LAYER M1 ;
        RECT 43.584 18.696 43.616 21.204 ;
  LAYER M3 ;
        RECT 43.584 18.716 43.616 18.748 ;
  LAYER M1 ;
        RECT 43.648 18.696 43.68 21.204 ;
  LAYER M3 ;
        RECT 43.648 21.152 43.68 21.184 ;
  LAYER M1 ;
        RECT 43.712 18.696 43.744 21.204 ;
  LAYER M3 ;
        RECT 43.712 18.716 43.744 18.748 ;
  LAYER M1 ;
        RECT 43.776 18.696 43.808 21.204 ;
  LAYER M3 ;
        RECT 43.776 21.152 43.808 21.184 ;
  LAYER M1 ;
        RECT 43.84 18.696 43.872 21.204 ;
  LAYER M3 ;
        RECT 43.84 18.716 43.872 18.748 ;
  LAYER M1 ;
        RECT 43.904 18.696 43.936 21.204 ;
  LAYER M3 ;
        RECT 41.536 21.088 41.568 21.12 ;
  LAYER M2 ;
        RECT 43.904 21.024 43.936 21.056 ;
  LAYER M2 ;
        RECT 41.536 20.96 41.568 20.992 ;
  LAYER M2 ;
        RECT 43.904 20.896 43.936 20.928 ;
  LAYER M2 ;
        RECT 41.536 20.832 41.568 20.864 ;
  LAYER M2 ;
        RECT 43.904 20.768 43.936 20.8 ;
  LAYER M2 ;
        RECT 41.536 20.704 41.568 20.736 ;
  LAYER M2 ;
        RECT 43.904 20.64 43.936 20.672 ;
  LAYER M2 ;
        RECT 41.536 20.576 41.568 20.608 ;
  LAYER M2 ;
        RECT 43.904 20.512 43.936 20.544 ;
  LAYER M2 ;
        RECT 41.536 20.448 41.568 20.48 ;
  LAYER M2 ;
        RECT 43.904 20.384 43.936 20.416 ;
  LAYER M2 ;
        RECT 41.536 20.32 41.568 20.352 ;
  LAYER M2 ;
        RECT 43.904 20.256 43.936 20.288 ;
  LAYER M2 ;
        RECT 41.536 20.192 41.568 20.224 ;
  LAYER M2 ;
        RECT 43.904 20.128 43.936 20.16 ;
  LAYER M2 ;
        RECT 41.536 20.064 41.568 20.096 ;
  LAYER M2 ;
        RECT 43.904 20 43.936 20.032 ;
  LAYER M2 ;
        RECT 41.536 19.936 41.568 19.968 ;
  LAYER M2 ;
        RECT 43.904 19.872 43.936 19.904 ;
  LAYER M2 ;
        RECT 41.536 19.808 41.568 19.84 ;
  LAYER M2 ;
        RECT 43.904 19.744 43.936 19.776 ;
  LAYER M2 ;
        RECT 41.536 19.68 41.568 19.712 ;
  LAYER M2 ;
        RECT 43.904 19.616 43.936 19.648 ;
  LAYER M2 ;
        RECT 41.536 19.552 41.568 19.584 ;
  LAYER M2 ;
        RECT 43.904 19.488 43.936 19.52 ;
  LAYER M2 ;
        RECT 41.536 19.424 41.568 19.456 ;
  LAYER M2 ;
        RECT 43.904 19.36 43.936 19.392 ;
  LAYER M2 ;
        RECT 41.536 19.296 41.568 19.328 ;
  LAYER M2 ;
        RECT 43.904 19.232 43.936 19.264 ;
  LAYER M2 ;
        RECT 41.536 19.168 41.568 19.2 ;
  LAYER M2 ;
        RECT 43.904 19.104 43.936 19.136 ;
  LAYER M2 ;
        RECT 41.536 19.04 41.568 19.072 ;
  LAYER M2 ;
        RECT 43.904 18.976 43.936 19.008 ;
  LAYER M2 ;
        RECT 41.536 18.912 41.568 18.944 ;
  LAYER M2 ;
        RECT 43.904 18.848 43.936 18.88 ;
  LAYER M2 ;
        RECT 41.488 18.648 43.984 21.252 ;
  LAYER M1 ;
        RECT 41.536 15.588 41.568 18.096 ;
  LAYER M3 ;
        RECT 41.536 15.608 41.568 15.64 ;
  LAYER M1 ;
        RECT 41.6 15.588 41.632 18.096 ;
  LAYER M3 ;
        RECT 41.6 18.044 41.632 18.076 ;
  LAYER M1 ;
        RECT 41.664 15.588 41.696 18.096 ;
  LAYER M3 ;
        RECT 41.664 15.608 41.696 15.64 ;
  LAYER M1 ;
        RECT 41.728 15.588 41.76 18.096 ;
  LAYER M3 ;
        RECT 41.728 18.044 41.76 18.076 ;
  LAYER M1 ;
        RECT 41.792 15.588 41.824 18.096 ;
  LAYER M3 ;
        RECT 41.792 15.608 41.824 15.64 ;
  LAYER M1 ;
        RECT 41.856 15.588 41.888 18.096 ;
  LAYER M3 ;
        RECT 41.856 18.044 41.888 18.076 ;
  LAYER M1 ;
        RECT 41.92 15.588 41.952 18.096 ;
  LAYER M3 ;
        RECT 41.92 15.608 41.952 15.64 ;
  LAYER M1 ;
        RECT 41.984 15.588 42.016 18.096 ;
  LAYER M3 ;
        RECT 41.984 18.044 42.016 18.076 ;
  LAYER M1 ;
        RECT 42.048 15.588 42.08 18.096 ;
  LAYER M3 ;
        RECT 42.048 15.608 42.08 15.64 ;
  LAYER M1 ;
        RECT 42.112 15.588 42.144 18.096 ;
  LAYER M3 ;
        RECT 42.112 18.044 42.144 18.076 ;
  LAYER M1 ;
        RECT 42.176 15.588 42.208 18.096 ;
  LAYER M3 ;
        RECT 42.176 15.608 42.208 15.64 ;
  LAYER M1 ;
        RECT 42.24 15.588 42.272 18.096 ;
  LAYER M3 ;
        RECT 42.24 18.044 42.272 18.076 ;
  LAYER M1 ;
        RECT 42.304 15.588 42.336 18.096 ;
  LAYER M3 ;
        RECT 42.304 15.608 42.336 15.64 ;
  LAYER M1 ;
        RECT 42.368 15.588 42.4 18.096 ;
  LAYER M3 ;
        RECT 42.368 18.044 42.4 18.076 ;
  LAYER M1 ;
        RECT 42.432 15.588 42.464 18.096 ;
  LAYER M3 ;
        RECT 42.432 15.608 42.464 15.64 ;
  LAYER M1 ;
        RECT 42.496 15.588 42.528 18.096 ;
  LAYER M3 ;
        RECT 42.496 18.044 42.528 18.076 ;
  LAYER M1 ;
        RECT 42.56 15.588 42.592 18.096 ;
  LAYER M3 ;
        RECT 42.56 15.608 42.592 15.64 ;
  LAYER M1 ;
        RECT 42.624 15.588 42.656 18.096 ;
  LAYER M3 ;
        RECT 42.624 18.044 42.656 18.076 ;
  LAYER M1 ;
        RECT 42.688 15.588 42.72 18.096 ;
  LAYER M3 ;
        RECT 42.688 15.608 42.72 15.64 ;
  LAYER M1 ;
        RECT 42.752 15.588 42.784 18.096 ;
  LAYER M3 ;
        RECT 42.752 18.044 42.784 18.076 ;
  LAYER M1 ;
        RECT 42.816 15.588 42.848 18.096 ;
  LAYER M3 ;
        RECT 42.816 15.608 42.848 15.64 ;
  LAYER M1 ;
        RECT 42.88 15.588 42.912 18.096 ;
  LAYER M3 ;
        RECT 42.88 18.044 42.912 18.076 ;
  LAYER M1 ;
        RECT 42.944 15.588 42.976 18.096 ;
  LAYER M3 ;
        RECT 42.944 15.608 42.976 15.64 ;
  LAYER M1 ;
        RECT 43.008 15.588 43.04 18.096 ;
  LAYER M3 ;
        RECT 43.008 18.044 43.04 18.076 ;
  LAYER M1 ;
        RECT 43.072 15.588 43.104 18.096 ;
  LAYER M3 ;
        RECT 43.072 15.608 43.104 15.64 ;
  LAYER M1 ;
        RECT 43.136 15.588 43.168 18.096 ;
  LAYER M3 ;
        RECT 43.136 18.044 43.168 18.076 ;
  LAYER M1 ;
        RECT 43.2 15.588 43.232 18.096 ;
  LAYER M3 ;
        RECT 43.2 15.608 43.232 15.64 ;
  LAYER M1 ;
        RECT 43.264 15.588 43.296 18.096 ;
  LAYER M3 ;
        RECT 43.264 18.044 43.296 18.076 ;
  LAYER M1 ;
        RECT 43.328 15.588 43.36 18.096 ;
  LAYER M3 ;
        RECT 43.328 15.608 43.36 15.64 ;
  LAYER M1 ;
        RECT 43.392 15.588 43.424 18.096 ;
  LAYER M3 ;
        RECT 43.392 18.044 43.424 18.076 ;
  LAYER M1 ;
        RECT 43.456 15.588 43.488 18.096 ;
  LAYER M3 ;
        RECT 43.456 15.608 43.488 15.64 ;
  LAYER M1 ;
        RECT 43.52 15.588 43.552 18.096 ;
  LAYER M3 ;
        RECT 43.52 18.044 43.552 18.076 ;
  LAYER M1 ;
        RECT 43.584 15.588 43.616 18.096 ;
  LAYER M3 ;
        RECT 43.584 15.608 43.616 15.64 ;
  LAYER M1 ;
        RECT 43.648 15.588 43.68 18.096 ;
  LAYER M3 ;
        RECT 43.648 18.044 43.68 18.076 ;
  LAYER M1 ;
        RECT 43.712 15.588 43.744 18.096 ;
  LAYER M3 ;
        RECT 43.712 15.608 43.744 15.64 ;
  LAYER M1 ;
        RECT 43.776 15.588 43.808 18.096 ;
  LAYER M3 ;
        RECT 43.776 18.044 43.808 18.076 ;
  LAYER M1 ;
        RECT 43.84 15.588 43.872 18.096 ;
  LAYER M3 ;
        RECT 43.84 15.608 43.872 15.64 ;
  LAYER M1 ;
        RECT 43.904 15.588 43.936 18.096 ;
  LAYER M3 ;
        RECT 41.536 17.98 41.568 18.012 ;
  LAYER M2 ;
        RECT 43.904 17.916 43.936 17.948 ;
  LAYER M2 ;
        RECT 41.536 17.852 41.568 17.884 ;
  LAYER M2 ;
        RECT 43.904 17.788 43.936 17.82 ;
  LAYER M2 ;
        RECT 41.536 17.724 41.568 17.756 ;
  LAYER M2 ;
        RECT 43.904 17.66 43.936 17.692 ;
  LAYER M2 ;
        RECT 41.536 17.596 41.568 17.628 ;
  LAYER M2 ;
        RECT 43.904 17.532 43.936 17.564 ;
  LAYER M2 ;
        RECT 41.536 17.468 41.568 17.5 ;
  LAYER M2 ;
        RECT 43.904 17.404 43.936 17.436 ;
  LAYER M2 ;
        RECT 41.536 17.34 41.568 17.372 ;
  LAYER M2 ;
        RECT 43.904 17.276 43.936 17.308 ;
  LAYER M2 ;
        RECT 41.536 17.212 41.568 17.244 ;
  LAYER M2 ;
        RECT 43.904 17.148 43.936 17.18 ;
  LAYER M2 ;
        RECT 41.536 17.084 41.568 17.116 ;
  LAYER M2 ;
        RECT 43.904 17.02 43.936 17.052 ;
  LAYER M2 ;
        RECT 41.536 16.956 41.568 16.988 ;
  LAYER M2 ;
        RECT 43.904 16.892 43.936 16.924 ;
  LAYER M2 ;
        RECT 41.536 16.828 41.568 16.86 ;
  LAYER M2 ;
        RECT 43.904 16.764 43.936 16.796 ;
  LAYER M2 ;
        RECT 41.536 16.7 41.568 16.732 ;
  LAYER M2 ;
        RECT 43.904 16.636 43.936 16.668 ;
  LAYER M2 ;
        RECT 41.536 16.572 41.568 16.604 ;
  LAYER M2 ;
        RECT 43.904 16.508 43.936 16.54 ;
  LAYER M2 ;
        RECT 41.536 16.444 41.568 16.476 ;
  LAYER M2 ;
        RECT 43.904 16.38 43.936 16.412 ;
  LAYER M2 ;
        RECT 41.536 16.316 41.568 16.348 ;
  LAYER M2 ;
        RECT 43.904 16.252 43.936 16.284 ;
  LAYER M2 ;
        RECT 41.536 16.188 41.568 16.22 ;
  LAYER M2 ;
        RECT 43.904 16.124 43.936 16.156 ;
  LAYER M2 ;
        RECT 41.536 16.06 41.568 16.092 ;
  LAYER M2 ;
        RECT 43.904 15.996 43.936 16.028 ;
  LAYER M2 ;
        RECT 41.536 15.932 41.568 15.964 ;
  LAYER M2 ;
        RECT 43.904 15.868 43.936 15.9 ;
  LAYER M2 ;
        RECT 41.536 15.804 41.568 15.836 ;
  LAYER M2 ;
        RECT 43.904 15.74 43.936 15.772 ;
  LAYER M2 ;
        RECT 41.488 15.54 43.984 18.144 ;
  LAYER M1 ;
        RECT 44.512 28.02 44.544 30.528 ;
  LAYER M3 ;
        RECT 44.512 28.04 44.544 28.072 ;
  LAYER M1 ;
        RECT 44.576 28.02 44.608 30.528 ;
  LAYER M3 ;
        RECT 44.576 30.476 44.608 30.508 ;
  LAYER M1 ;
        RECT 44.64 28.02 44.672 30.528 ;
  LAYER M3 ;
        RECT 44.64 28.04 44.672 28.072 ;
  LAYER M1 ;
        RECT 44.704 28.02 44.736 30.528 ;
  LAYER M3 ;
        RECT 44.704 30.476 44.736 30.508 ;
  LAYER M1 ;
        RECT 44.768 28.02 44.8 30.528 ;
  LAYER M3 ;
        RECT 44.768 28.04 44.8 28.072 ;
  LAYER M1 ;
        RECT 44.832 28.02 44.864 30.528 ;
  LAYER M3 ;
        RECT 44.832 30.476 44.864 30.508 ;
  LAYER M1 ;
        RECT 44.896 28.02 44.928 30.528 ;
  LAYER M3 ;
        RECT 44.896 28.04 44.928 28.072 ;
  LAYER M1 ;
        RECT 44.96 28.02 44.992 30.528 ;
  LAYER M3 ;
        RECT 44.96 30.476 44.992 30.508 ;
  LAYER M1 ;
        RECT 45.024 28.02 45.056 30.528 ;
  LAYER M3 ;
        RECT 45.024 28.04 45.056 28.072 ;
  LAYER M1 ;
        RECT 45.088 28.02 45.12 30.528 ;
  LAYER M3 ;
        RECT 45.088 30.476 45.12 30.508 ;
  LAYER M1 ;
        RECT 45.152 28.02 45.184 30.528 ;
  LAYER M3 ;
        RECT 45.152 28.04 45.184 28.072 ;
  LAYER M1 ;
        RECT 45.216 28.02 45.248 30.528 ;
  LAYER M3 ;
        RECT 45.216 30.476 45.248 30.508 ;
  LAYER M1 ;
        RECT 45.28 28.02 45.312 30.528 ;
  LAYER M3 ;
        RECT 45.28 28.04 45.312 28.072 ;
  LAYER M1 ;
        RECT 45.344 28.02 45.376 30.528 ;
  LAYER M3 ;
        RECT 45.344 30.476 45.376 30.508 ;
  LAYER M1 ;
        RECT 45.408 28.02 45.44 30.528 ;
  LAYER M3 ;
        RECT 45.408 28.04 45.44 28.072 ;
  LAYER M1 ;
        RECT 45.472 28.02 45.504 30.528 ;
  LAYER M3 ;
        RECT 45.472 30.476 45.504 30.508 ;
  LAYER M1 ;
        RECT 45.536 28.02 45.568 30.528 ;
  LAYER M3 ;
        RECT 45.536 28.04 45.568 28.072 ;
  LAYER M1 ;
        RECT 45.6 28.02 45.632 30.528 ;
  LAYER M3 ;
        RECT 45.6 30.476 45.632 30.508 ;
  LAYER M1 ;
        RECT 45.664 28.02 45.696 30.528 ;
  LAYER M3 ;
        RECT 45.664 28.04 45.696 28.072 ;
  LAYER M1 ;
        RECT 45.728 28.02 45.76 30.528 ;
  LAYER M3 ;
        RECT 45.728 30.476 45.76 30.508 ;
  LAYER M1 ;
        RECT 45.792 28.02 45.824 30.528 ;
  LAYER M3 ;
        RECT 45.792 28.04 45.824 28.072 ;
  LAYER M1 ;
        RECT 45.856 28.02 45.888 30.528 ;
  LAYER M3 ;
        RECT 45.856 30.476 45.888 30.508 ;
  LAYER M1 ;
        RECT 45.92 28.02 45.952 30.528 ;
  LAYER M3 ;
        RECT 45.92 28.04 45.952 28.072 ;
  LAYER M1 ;
        RECT 45.984 28.02 46.016 30.528 ;
  LAYER M3 ;
        RECT 45.984 30.476 46.016 30.508 ;
  LAYER M1 ;
        RECT 46.048 28.02 46.08 30.528 ;
  LAYER M3 ;
        RECT 46.048 28.04 46.08 28.072 ;
  LAYER M1 ;
        RECT 46.112 28.02 46.144 30.528 ;
  LAYER M3 ;
        RECT 46.112 30.476 46.144 30.508 ;
  LAYER M1 ;
        RECT 46.176 28.02 46.208 30.528 ;
  LAYER M3 ;
        RECT 46.176 28.04 46.208 28.072 ;
  LAYER M1 ;
        RECT 46.24 28.02 46.272 30.528 ;
  LAYER M3 ;
        RECT 46.24 30.476 46.272 30.508 ;
  LAYER M1 ;
        RECT 46.304 28.02 46.336 30.528 ;
  LAYER M3 ;
        RECT 46.304 28.04 46.336 28.072 ;
  LAYER M1 ;
        RECT 46.368 28.02 46.4 30.528 ;
  LAYER M3 ;
        RECT 46.368 30.476 46.4 30.508 ;
  LAYER M1 ;
        RECT 46.432 28.02 46.464 30.528 ;
  LAYER M3 ;
        RECT 46.432 28.04 46.464 28.072 ;
  LAYER M1 ;
        RECT 46.496 28.02 46.528 30.528 ;
  LAYER M3 ;
        RECT 46.496 30.476 46.528 30.508 ;
  LAYER M1 ;
        RECT 46.56 28.02 46.592 30.528 ;
  LAYER M3 ;
        RECT 46.56 28.04 46.592 28.072 ;
  LAYER M1 ;
        RECT 46.624 28.02 46.656 30.528 ;
  LAYER M3 ;
        RECT 46.624 30.476 46.656 30.508 ;
  LAYER M1 ;
        RECT 46.688 28.02 46.72 30.528 ;
  LAYER M3 ;
        RECT 46.688 28.04 46.72 28.072 ;
  LAYER M1 ;
        RECT 46.752 28.02 46.784 30.528 ;
  LAYER M3 ;
        RECT 46.752 30.476 46.784 30.508 ;
  LAYER M1 ;
        RECT 46.816 28.02 46.848 30.528 ;
  LAYER M3 ;
        RECT 46.816 28.04 46.848 28.072 ;
  LAYER M1 ;
        RECT 46.88 28.02 46.912 30.528 ;
  LAYER M3 ;
        RECT 44.512 30.412 44.544 30.444 ;
  LAYER M2 ;
        RECT 46.88 30.348 46.912 30.38 ;
  LAYER M2 ;
        RECT 44.512 30.284 44.544 30.316 ;
  LAYER M2 ;
        RECT 46.88 30.22 46.912 30.252 ;
  LAYER M2 ;
        RECT 44.512 30.156 44.544 30.188 ;
  LAYER M2 ;
        RECT 46.88 30.092 46.912 30.124 ;
  LAYER M2 ;
        RECT 44.512 30.028 44.544 30.06 ;
  LAYER M2 ;
        RECT 46.88 29.964 46.912 29.996 ;
  LAYER M2 ;
        RECT 44.512 29.9 44.544 29.932 ;
  LAYER M2 ;
        RECT 46.88 29.836 46.912 29.868 ;
  LAYER M2 ;
        RECT 44.512 29.772 44.544 29.804 ;
  LAYER M2 ;
        RECT 46.88 29.708 46.912 29.74 ;
  LAYER M2 ;
        RECT 44.512 29.644 44.544 29.676 ;
  LAYER M2 ;
        RECT 46.88 29.58 46.912 29.612 ;
  LAYER M2 ;
        RECT 44.512 29.516 44.544 29.548 ;
  LAYER M2 ;
        RECT 46.88 29.452 46.912 29.484 ;
  LAYER M2 ;
        RECT 44.512 29.388 44.544 29.42 ;
  LAYER M2 ;
        RECT 46.88 29.324 46.912 29.356 ;
  LAYER M2 ;
        RECT 44.512 29.26 44.544 29.292 ;
  LAYER M2 ;
        RECT 46.88 29.196 46.912 29.228 ;
  LAYER M2 ;
        RECT 44.512 29.132 44.544 29.164 ;
  LAYER M2 ;
        RECT 46.88 29.068 46.912 29.1 ;
  LAYER M2 ;
        RECT 44.512 29.004 44.544 29.036 ;
  LAYER M2 ;
        RECT 46.88 28.94 46.912 28.972 ;
  LAYER M2 ;
        RECT 44.512 28.876 44.544 28.908 ;
  LAYER M2 ;
        RECT 46.88 28.812 46.912 28.844 ;
  LAYER M2 ;
        RECT 44.512 28.748 44.544 28.78 ;
  LAYER M2 ;
        RECT 46.88 28.684 46.912 28.716 ;
  LAYER M2 ;
        RECT 44.512 28.62 44.544 28.652 ;
  LAYER M2 ;
        RECT 46.88 28.556 46.912 28.588 ;
  LAYER M2 ;
        RECT 44.512 28.492 44.544 28.524 ;
  LAYER M2 ;
        RECT 46.88 28.428 46.912 28.46 ;
  LAYER M2 ;
        RECT 44.512 28.364 44.544 28.396 ;
  LAYER M2 ;
        RECT 46.88 28.3 46.912 28.332 ;
  LAYER M2 ;
        RECT 44.512 28.236 44.544 28.268 ;
  LAYER M2 ;
        RECT 46.88 28.172 46.912 28.204 ;
  LAYER M2 ;
        RECT 44.464 27.972 46.96 30.576 ;
  LAYER M1 ;
        RECT 44.512 24.912 44.544 27.42 ;
  LAYER M3 ;
        RECT 44.512 24.932 44.544 24.964 ;
  LAYER M1 ;
        RECT 44.576 24.912 44.608 27.42 ;
  LAYER M3 ;
        RECT 44.576 27.368 44.608 27.4 ;
  LAYER M1 ;
        RECT 44.64 24.912 44.672 27.42 ;
  LAYER M3 ;
        RECT 44.64 24.932 44.672 24.964 ;
  LAYER M1 ;
        RECT 44.704 24.912 44.736 27.42 ;
  LAYER M3 ;
        RECT 44.704 27.368 44.736 27.4 ;
  LAYER M1 ;
        RECT 44.768 24.912 44.8 27.42 ;
  LAYER M3 ;
        RECT 44.768 24.932 44.8 24.964 ;
  LAYER M1 ;
        RECT 44.832 24.912 44.864 27.42 ;
  LAYER M3 ;
        RECT 44.832 27.368 44.864 27.4 ;
  LAYER M1 ;
        RECT 44.896 24.912 44.928 27.42 ;
  LAYER M3 ;
        RECT 44.896 24.932 44.928 24.964 ;
  LAYER M1 ;
        RECT 44.96 24.912 44.992 27.42 ;
  LAYER M3 ;
        RECT 44.96 27.368 44.992 27.4 ;
  LAYER M1 ;
        RECT 45.024 24.912 45.056 27.42 ;
  LAYER M3 ;
        RECT 45.024 24.932 45.056 24.964 ;
  LAYER M1 ;
        RECT 45.088 24.912 45.12 27.42 ;
  LAYER M3 ;
        RECT 45.088 27.368 45.12 27.4 ;
  LAYER M1 ;
        RECT 45.152 24.912 45.184 27.42 ;
  LAYER M3 ;
        RECT 45.152 24.932 45.184 24.964 ;
  LAYER M1 ;
        RECT 45.216 24.912 45.248 27.42 ;
  LAYER M3 ;
        RECT 45.216 27.368 45.248 27.4 ;
  LAYER M1 ;
        RECT 45.28 24.912 45.312 27.42 ;
  LAYER M3 ;
        RECT 45.28 24.932 45.312 24.964 ;
  LAYER M1 ;
        RECT 45.344 24.912 45.376 27.42 ;
  LAYER M3 ;
        RECT 45.344 27.368 45.376 27.4 ;
  LAYER M1 ;
        RECT 45.408 24.912 45.44 27.42 ;
  LAYER M3 ;
        RECT 45.408 24.932 45.44 24.964 ;
  LAYER M1 ;
        RECT 45.472 24.912 45.504 27.42 ;
  LAYER M3 ;
        RECT 45.472 27.368 45.504 27.4 ;
  LAYER M1 ;
        RECT 45.536 24.912 45.568 27.42 ;
  LAYER M3 ;
        RECT 45.536 24.932 45.568 24.964 ;
  LAYER M1 ;
        RECT 45.6 24.912 45.632 27.42 ;
  LAYER M3 ;
        RECT 45.6 27.368 45.632 27.4 ;
  LAYER M1 ;
        RECT 45.664 24.912 45.696 27.42 ;
  LAYER M3 ;
        RECT 45.664 24.932 45.696 24.964 ;
  LAYER M1 ;
        RECT 45.728 24.912 45.76 27.42 ;
  LAYER M3 ;
        RECT 45.728 27.368 45.76 27.4 ;
  LAYER M1 ;
        RECT 45.792 24.912 45.824 27.42 ;
  LAYER M3 ;
        RECT 45.792 24.932 45.824 24.964 ;
  LAYER M1 ;
        RECT 45.856 24.912 45.888 27.42 ;
  LAYER M3 ;
        RECT 45.856 27.368 45.888 27.4 ;
  LAYER M1 ;
        RECT 45.92 24.912 45.952 27.42 ;
  LAYER M3 ;
        RECT 45.92 24.932 45.952 24.964 ;
  LAYER M1 ;
        RECT 45.984 24.912 46.016 27.42 ;
  LAYER M3 ;
        RECT 45.984 27.368 46.016 27.4 ;
  LAYER M1 ;
        RECT 46.048 24.912 46.08 27.42 ;
  LAYER M3 ;
        RECT 46.048 24.932 46.08 24.964 ;
  LAYER M1 ;
        RECT 46.112 24.912 46.144 27.42 ;
  LAYER M3 ;
        RECT 46.112 27.368 46.144 27.4 ;
  LAYER M1 ;
        RECT 46.176 24.912 46.208 27.42 ;
  LAYER M3 ;
        RECT 46.176 24.932 46.208 24.964 ;
  LAYER M1 ;
        RECT 46.24 24.912 46.272 27.42 ;
  LAYER M3 ;
        RECT 46.24 27.368 46.272 27.4 ;
  LAYER M1 ;
        RECT 46.304 24.912 46.336 27.42 ;
  LAYER M3 ;
        RECT 46.304 24.932 46.336 24.964 ;
  LAYER M1 ;
        RECT 46.368 24.912 46.4 27.42 ;
  LAYER M3 ;
        RECT 46.368 27.368 46.4 27.4 ;
  LAYER M1 ;
        RECT 46.432 24.912 46.464 27.42 ;
  LAYER M3 ;
        RECT 46.432 24.932 46.464 24.964 ;
  LAYER M1 ;
        RECT 46.496 24.912 46.528 27.42 ;
  LAYER M3 ;
        RECT 46.496 27.368 46.528 27.4 ;
  LAYER M1 ;
        RECT 46.56 24.912 46.592 27.42 ;
  LAYER M3 ;
        RECT 46.56 24.932 46.592 24.964 ;
  LAYER M1 ;
        RECT 46.624 24.912 46.656 27.42 ;
  LAYER M3 ;
        RECT 46.624 27.368 46.656 27.4 ;
  LAYER M1 ;
        RECT 46.688 24.912 46.72 27.42 ;
  LAYER M3 ;
        RECT 46.688 24.932 46.72 24.964 ;
  LAYER M1 ;
        RECT 46.752 24.912 46.784 27.42 ;
  LAYER M3 ;
        RECT 46.752 27.368 46.784 27.4 ;
  LAYER M1 ;
        RECT 46.816 24.912 46.848 27.42 ;
  LAYER M3 ;
        RECT 46.816 24.932 46.848 24.964 ;
  LAYER M1 ;
        RECT 46.88 24.912 46.912 27.42 ;
  LAYER M3 ;
        RECT 44.512 27.304 44.544 27.336 ;
  LAYER M2 ;
        RECT 46.88 27.24 46.912 27.272 ;
  LAYER M2 ;
        RECT 44.512 27.176 44.544 27.208 ;
  LAYER M2 ;
        RECT 46.88 27.112 46.912 27.144 ;
  LAYER M2 ;
        RECT 44.512 27.048 44.544 27.08 ;
  LAYER M2 ;
        RECT 46.88 26.984 46.912 27.016 ;
  LAYER M2 ;
        RECT 44.512 26.92 44.544 26.952 ;
  LAYER M2 ;
        RECT 46.88 26.856 46.912 26.888 ;
  LAYER M2 ;
        RECT 44.512 26.792 44.544 26.824 ;
  LAYER M2 ;
        RECT 46.88 26.728 46.912 26.76 ;
  LAYER M2 ;
        RECT 44.512 26.664 44.544 26.696 ;
  LAYER M2 ;
        RECT 46.88 26.6 46.912 26.632 ;
  LAYER M2 ;
        RECT 44.512 26.536 44.544 26.568 ;
  LAYER M2 ;
        RECT 46.88 26.472 46.912 26.504 ;
  LAYER M2 ;
        RECT 44.512 26.408 44.544 26.44 ;
  LAYER M2 ;
        RECT 46.88 26.344 46.912 26.376 ;
  LAYER M2 ;
        RECT 44.512 26.28 44.544 26.312 ;
  LAYER M2 ;
        RECT 46.88 26.216 46.912 26.248 ;
  LAYER M2 ;
        RECT 44.512 26.152 44.544 26.184 ;
  LAYER M2 ;
        RECT 46.88 26.088 46.912 26.12 ;
  LAYER M2 ;
        RECT 44.512 26.024 44.544 26.056 ;
  LAYER M2 ;
        RECT 46.88 25.96 46.912 25.992 ;
  LAYER M2 ;
        RECT 44.512 25.896 44.544 25.928 ;
  LAYER M2 ;
        RECT 46.88 25.832 46.912 25.864 ;
  LAYER M2 ;
        RECT 44.512 25.768 44.544 25.8 ;
  LAYER M2 ;
        RECT 46.88 25.704 46.912 25.736 ;
  LAYER M2 ;
        RECT 44.512 25.64 44.544 25.672 ;
  LAYER M2 ;
        RECT 46.88 25.576 46.912 25.608 ;
  LAYER M2 ;
        RECT 44.512 25.512 44.544 25.544 ;
  LAYER M2 ;
        RECT 46.88 25.448 46.912 25.48 ;
  LAYER M2 ;
        RECT 44.512 25.384 44.544 25.416 ;
  LAYER M2 ;
        RECT 46.88 25.32 46.912 25.352 ;
  LAYER M2 ;
        RECT 44.512 25.256 44.544 25.288 ;
  LAYER M2 ;
        RECT 46.88 25.192 46.912 25.224 ;
  LAYER M2 ;
        RECT 44.512 25.128 44.544 25.16 ;
  LAYER M2 ;
        RECT 46.88 25.064 46.912 25.096 ;
  LAYER M2 ;
        RECT 44.464 24.864 46.96 27.468 ;
  LAYER M1 ;
        RECT 44.512 21.804 44.544 24.312 ;
  LAYER M3 ;
        RECT 44.512 21.824 44.544 21.856 ;
  LAYER M1 ;
        RECT 44.576 21.804 44.608 24.312 ;
  LAYER M3 ;
        RECT 44.576 24.26 44.608 24.292 ;
  LAYER M1 ;
        RECT 44.64 21.804 44.672 24.312 ;
  LAYER M3 ;
        RECT 44.64 21.824 44.672 21.856 ;
  LAYER M1 ;
        RECT 44.704 21.804 44.736 24.312 ;
  LAYER M3 ;
        RECT 44.704 24.26 44.736 24.292 ;
  LAYER M1 ;
        RECT 44.768 21.804 44.8 24.312 ;
  LAYER M3 ;
        RECT 44.768 21.824 44.8 21.856 ;
  LAYER M1 ;
        RECT 44.832 21.804 44.864 24.312 ;
  LAYER M3 ;
        RECT 44.832 24.26 44.864 24.292 ;
  LAYER M1 ;
        RECT 44.896 21.804 44.928 24.312 ;
  LAYER M3 ;
        RECT 44.896 21.824 44.928 21.856 ;
  LAYER M1 ;
        RECT 44.96 21.804 44.992 24.312 ;
  LAYER M3 ;
        RECT 44.96 24.26 44.992 24.292 ;
  LAYER M1 ;
        RECT 45.024 21.804 45.056 24.312 ;
  LAYER M3 ;
        RECT 45.024 21.824 45.056 21.856 ;
  LAYER M1 ;
        RECT 45.088 21.804 45.12 24.312 ;
  LAYER M3 ;
        RECT 45.088 24.26 45.12 24.292 ;
  LAYER M1 ;
        RECT 45.152 21.804 45.184 24.312 ;
  LAYER M3 ;
        RECT 45.152 21.824 45.184 21.856 ;
  LAYER M1 ;
        RECT 45.216 21.804 45.248 24.312 ;
  LAYER M3 ;
        RECT 45.216 24.26 45.248 24.292 ;
  LAYER M1 ;
        RECT 45.28 21.804 45.312 24.312 ;
  LAYER M3 ;
        RECT 45.28 21.824 45.312 21.856 ;
  LAYER M1 ;
        RECT 45.344 21.804 45.376 24.312 ;
  LAYER M3 ;
        RECT 45.344 24.26 45.376 24.292 ;
  LAYER M1 ;
        RECT 45.408 21.804 45.44 24.312 ;
  LAYER M3 ;
        RECT 45.408 21.824 45.44 21.856 ;
  LAYER M1 ;
        RECT 45.472 21.804 45.504 24.312 ;
  LAYER M3 ;
        RECT 45.472 24.26 45.504 24.292 ;
  LAYER M1 ;
        RECT 45.536 21.804 45.568 24.312 ;
  LAYER M3 ;
        RECT 45.536 21.824 45.568 21.856 ;
  LAYER M1 ;
        RECT 45.6 21.804 45.632 24.312 ;
  LAYER M3 ;
        RECT 45.6 24.26 45.632 24.292 ;
  LAYER M1 ;
        RECT 45.664 21.804 45.696 24.312 ;
  LAYER M3 ;
        RECT 45.664 21.824 45.696 21.856 ;
  LAYER M1 ;
        RECT 45.728 21.804 45.76 24.312 ;
  LAYER M3 ;
        RECT 45.728 24.26 45.76 24.292 ;
  LAYER M1 ;
        RECT 45.792 21.804 45.824 24.312 ;
  LAYER M3 ;
        RECT 45.792 21.824 45.824 21.856 ;
  LAYER M1 ;
        RECT 45.856 21.804 45.888 24.312 ;
  LAYER M3 ;
        RECT 45.856 24.26 45.888 24.292 ;
  LAYER M1 ;
        RECT 45.92 21.804 45.952 24.312 ;
  LAYER M3 ;
        RECT 45.92 21.824 45.952 21.856 ;
  LAYER M1 ;
        RECT 45.984 21.804 46.016 24.312 ;
  LAYER M3 ;
        RECT 45.984 24.26 46.016 24.292 ;
  LAYER M1 ;
        RECT 46.048 21.804 46.08 24.312 ;
  LAYER M3 ;
        RECT 46.048 21.824 46.08 21.856 ;
  LAYER M1 ;
        RECT 46.112 21.804 46.144 24.312 ;
  LAYER M3 ;
        RECT 46.112 24.26 46.144 24.292 ;
  LAYER M1 ;
        RECT 46.176 21.804 46.208 24.312 ;
  LAYER M3 ;
        RECT 46.176 21.824 46.208 21.856 ;
  LAYER M1 ;
        RECT 46.24 21.804 46.272 24.312 ;
  LAYER M3 ;
        RECT 46.24 24.26 46.272 24.292 ;
  LAYER M1 ;
        RECT 46.304 21.804 46.336 24.312 ;
  LAYER M3 ;
        RECT 46.304 21.824 46.336 21.856 ;
  LAYER M1 ;
        RECT 46.368 21.804 46.4 24.312 ;
  LAYER M3 ;
        RECT 46.368 24.26 46.4 24.292 ;
  LAYER M1 ;
        RECT 46.432 21.804 46.464 24.312 ;
  LAYER M3 ;
        RECT 46.432 21.824 46.464 21.856 ;
  LAYER M1 ;
        RECT 46.496 21.804 46.528 24.312 ;
  LAYER M3 ;
        RECT 46.496 24.26 46.528 24.292 ;
  LAYER M1 ;
        RECT 46.56 21.804 46.592 24.312 ;
  LAYER M3 ;
        RECT 46.56 21.824 46.592 21.856 ;
  LAYER M1 ;
        RECT 46.624 21.804 46.656 24.312 ;
  LAYER M3 ;
        RECT 46.624 24.26 46.656 24.292 ;
  LAYER M1 ;
        RECT 46.688 21.804 46.72 24.312 ;
  LAYER M3 ;
        RECT 46.688 21.824 46.72 21.856 ;
  LAYER M1 ;
        RECT 46.752 21.804 46.784 24.312 ;
  LAYER M3 ;
        RECT 46.752 24.26 46.784 24.292 ;
  LAYER M1 ;
        RECT 46.816 21.804 46.848 24.312 ;
  LAYER M3 ;
        RECT 46.816 21.824 46.848 21.856 ;
  LAYER M1 ;
        RECT 46.88 21.804 46.912 24.312 ;
  LAYER M3 ;
        RECT 44.512 24.196 44.544 24.228 ;
  LAYER M2 ;
        RECT 46.88 24.132 46.912 24.164 ;
  LAYER M2 ;
        RECT 44.512 24.068 44.544 24.1 ;
  LAYER M2 ;
        RECT 46.88 24.004 46.912 24.036 ;
  LAYER M2 ;
        RECT 44.512 23.94 44.544 23.972 ;
  LAYER M2 ;
        RECT 46.88 23.876 46.912 23.908 ;
  LAYER M2 ;
        RECT 44.512 23.812 44.544 23.844 ;
  LAYER M2 ;
        RECT 46.88 23.748 46.912 23.78 ;
  LAYER M2 ;
        RECT 44.512 23.684 44.544 23.716 ;
  LAYER M2 ;
        RECT 46.88 23.62 46.912 23.652 ;
  LAYER M2 ;
        RECT 44.512 23.556 44.544 23.588 ;
  LAYER M2 ;
        RECT 46.88 23.492 46.912 23.524 ;
  LAYER M2 ;
        RECT 44.512 23.428 44.544 23.46 ;
  LAYER M2 ;
        RECT 46.88 23.364 46.912 23.396 ;
  LAYER M2 ;
        RECT 44.512 23.3 44.544 23.332 ;
  LAYER M2 ;
        RECT 46.88 23.236 46.912 23.268 ;
  LAYER M2 ;
        RECT 44.512 23.172 44.544 23.204 ;
  LAYER M2 ;
        RECT 46.88 23.108 46.912 23.14 ;
  LAYER M2 ;
        RECT 44.512 23.044 44.544 23.076 ;
  LAYER M2 ;
        RECT 46.88 22.98 46.912 23.012 ;
  LAYER M2 ;
        RECT 44.512 22.916 44.544 22.948 ;
  LAYER M2 ;
        RECT 46.88 22.852 46.912 22.884 ;
  LAYER M2 ;
        RECT 44.512 22.788 44.544 22.82 ;
  LAYER M2 ;
        RECT 46.88 22.724 46.912 22.756 ;
  LAYER M2 ;
        RECT 44.512 22.66 44.544 22.692 ;
  LAYER M2 ;
        RECT 46.88 22.596 46.912 22.628 ;
  LAYER M2 ;
        RECT 44.512 22.532 44.544 22.564 ;
  LAYER M2 ;
        RECT 46.88 22.468 46.912 22.5 ;
  LAYER M2 ;
        RECT 44.512 22.404 44.544 22.436 ;
  LAYER M2 ;
        RECT 46.88 22.34 46.912 22.372 ;
  LAYER M2 ;
        RECT 44.512 22.276 44.544 22.308 ;
  LAYER M2 ;
        RECT 46.88 22.212 46.912 22.244 ;
  LAYER M2 ;
        RECT 44.512 22.148 44.544 22.18 ;
  LAYER M2 ;
        RECT 46.88 22.084 46.912 22.116 ;
  LAYER M2 ;
        RECT 44.512 22.02 44.544 22.052 ;
  LAYER M2 ;
        RECT 46.88 21.956 46.912 21.988 ;
  LAYER M2 ;
        RECT 44.464 21.756 46.96 24.36 ;
  LAYER M1 ;
        RECT 44.512 18.696 44.544 21.204 ;
  LAYER M3 ;
        RECT 44.512 18.716 44.544 18.748 ;
  LAYER M1 ;
        RECT 44.576 18.696 44.608 21.204 ;
  LAYER M3 ;
        RECT 44.576 21.152 44.608 21.184 ;
  LAYER M1 ;
        RECT 44.64 18.696 44.672 21.204 ;
  LAYER M3 ;
        RECT 44.64 18.716 44.672 18.748 ;
  LAYER M1 ;
        RECT 44.704 18.696 44.736 21.204 ;
  LAYER M3 ;
        RECT 44.704 21.152 44.736 21.184 ;
  LAYER M1 ;
        RECT 44.768 18.696 44.8 21.204 ;
  LAYER M3 ;
        RECT 44.768 18.716 44.8 18.748 ;
  LAYER M1 ;
        RECT 44.832 18.696 44.864 21.204 ;
  LAYER M3 ;
        RECT 44.832 21.152 44.864 21.184 ;
  LAYER M1 ;
        RECT 44.896 18.696 44.928 21.204 ;
  LAYER M3 ;
        RECT 44.896 18.716 44.928 18.748 ;
  LAYER M1 ;
        RECT 44.96 18.696 44.992 21.204 ;
  LAYER M3 ;
        RECT 44.96 21.152 44.992 21.184 ;
  LAYER M1 ;
        RECT 45.024 18.696 45.056 21.204 ;
  LAYER M3 ;
        RECT 45.024 18.716 45.056 18.748 ;
  LAYER M1 ;
        RECT 45.088 18.696 45.12 21.204 ;
  LAYER M3 ;
        RECT 45.088 21.152 45.12 21.184 ;
  LAYER M1 ;
        RECT 45.152 18.696 45.184 21.204 ;
  LAYER M3 ;
        RECT 45.152 18.716 45.184 18.748 ;
  LAYER M1 ;
        RECT 45.216 18.696 45.248 21.204 ;
  LAYER M3 ;
        RECT 45.216 21.152 45.248 21.184 ;
  LAYER M1 ;
        RECT 45.28 18.696 45.312 21.204 ;
  LAYER M3 ;
        RECT 45.28 18.716 45.312 18.748 ;
  LAYER M1 ;
        RECT 45.344 18.696 45.376 21.204 ;
  LAYER M3 ;
        RECT 45.344 21.152 45.376 21.184 ;
  LAYER M1 ;
        RECT 45.408 18.696 45.44 21.204 ;
  LAYER M3 ;
        RECT 45.408 18.716 45.44 18.748 ;
  LAYER M1 ;
        RECT 45.472 18.696 45.504 21.204 ;
  LAYER M3 ;
        RECT 45.472 21.152 45.504 21.184 ;
  LAYER M1 ;
        RECT 45.536 18.696 45.568 21.204 ;
  LAYER M3 ;
        RECT 45.536 18.716 45.568 18.748 ;
  LAYER M1 ;
        RECT 45.6 18.696 45.632 21.204 ;
  LAYER M3 ;
        RECT 45.6 21.152 45.632 21.184 ;
  LAYER M1 ;
        RECT 45.664 18.696 45.696 21.204 ;
  LAYER M3 ;
        RECT 45.664 18.716 45.696 18.748 ;
  LAYER M1 ;
        RECT 45.728 18.696 45.76 21.204 ;
  LAYER M3 ;
        RECT 45.728 21.152 45.76 21.184 ;
  LAYER M1 ;
        RECT 45.792 18.696 45.824 21.204 ;
  LAYER M3 ;
        RECT 45.792 18.716 45.824 18.748 ;
  LAYER M1 ;
        RECT 45.856 18.696 45.888 21.204 ;
  LAYER M3 ;
        RECT 45.856 21.152 45.888 21.184 ;
  LAYER M1 ;
        RECT 45.92 18.696 45.952 21.204 ;
  LAYER M3 ;
        RECT 45.92 18.716 45.952 18.748 ;
  LAYER M1 ;
        RECT 45.984 18.696 46.016 21.204 ;
  LAYER M3 ;
        RECT 45.984 21.152 46.016 21.184 ;
  LAYER M1 ;
        RECT 46.048 18.696 46.08 21.204 ;
  LAYER M3 ;
        RECT 46.048 18.716 46.08 18.748 ;
  LAYER M1 ;
        RECT 46.112 18.696 46.144 21.204 ;
  LAYER M3 ;
        RECT 46.112 21.152 46.144 21.184 ;
  LAYER M1 ;
        RECT 46.176 18.696 46.208 21.204 ;
  LAYER M3 ;
        RECT 46.176 18.716 46.208 18.748 ;
  LAYER M1 ;
        RECT 46.24 18.696 46.272 21.204 ;
  LAYER M3 ;
        RECT 46.24 21.152 46.272 21.184 ;
  LAYER M1 ;
        RECT 46.304 18.696 46.336 21.204 ;
  LAYER M3 ;
        RECT 46.304 18.716 46.336 18.748 ;
  LAYER M1 ;
        RECT 46.368 18.696 46.4 21.204 ;
  LAYER M3 ;
        RECT 46.368 21.152 46.4 21.184 ;
  LAYER M1 ;
        RECT 46.432 18.696 46.464 21.204 ;
  LAYER M3 ;
        RECT 46.432 18.716 46.464 18.748 ;
  LAYER M1 ;
        RECT 46.496 18.696 46.528 21.204 ;
  LAYER M3 ;
        RECT 46.496 21.152 46.528 21.184 ;
  LAYER M1 ;
        RECT 46.56 18.696 46.592 21.204 ;
  LAYER M3 ;
        RECT 46.56 18.716 46.592 18.748 ;
  LAYER M1 ;
        RECT 46.624 18.696 46.656 21.204 ;
  LAYER M3 ;
        RECT 46.624 21.152 46.656 21.184 ;
  LAYER M1 ;
        RECT 46.688 18.696 46.72 21.204 ;
  LAYER M3 ;
        RECT 46.688 18.716 46.72 18.748 ;
  LAYER M1 ;
        RECT 46.752 18.696 46.784 21.204 ;
  LAYER M3 ;
        RECT 46.752 21.152 46.784 21.184 ;
  LAYER M1 ;
        RECT 46.816 18.696 46.848 21.204 ;
  LAYER M3 ;
        RECT 46.816 18.716 46.848 18.748 ;
  LAYER M1 ;
        RECT 46.88 18.696 46.912 21.204 ;
  LAYER M3 ;
        RECT 44.512 21.088 44.544 21.12 ;
  LAYER M2 ;
        RECT 46.88 21.024 46.912 21.056 ;
  LAYER M2 ;
        RECT 44.512 20.96 44.544 20.992 ;
  LAYER M2 ;
        RECT 46.88 20.896 46.912 20.928 ;
  LAYER M2 ;
        RECT 44.512 20.832 44.544 20.864 ;
  LAYER M2 ;
        RECT 46.88 20.768 46.912 20.8 ;
  LAYER M2 ;
        RECT 44.512 20.704 44.544 20.736 ;
  LAYER M2 ;
        RECT 46.88 20.64 46.912 20.672 ;
  LAYER M2 ;
        RECT 44.512 20.576 44.544 20.608 ;
  LAYER M2 ;
        RECT 46.88 20.512 46.912 20.544 ;
  LAYER M2 ;
        RECT 44.512 20.448 44.544 20.48 ;
  LAYER M2 ;
        RECT 46.88 20.384 46.912 20.416 ;
  LAYER M2 ;
        RECT 44.512 20.32 44.544 20.352 ;
  LAYER M2 ;
        RECT 46.88 20.256 46.912 20.288 ;
  LAYER M2 ;
        RECT 44.512 20.192 44.544 20.224 ;
  LAYER M2 ;
        RECT 46.88 20.128 46.912 20.16 ;
  LAYER M2 ;
        RECT 44.512 20.064 44.544 20.096 ;
  LAYER M2 ;
        RECT 46.88 20 46.912 20.032 ;
  LAYER M2 ;
        RECT 44.512 19.936 44.544 19.968 ;
  LAYER M2 ;
        RECT 46.88 19.872 46.912 19.904 ;
  LAYER M2 ;
        RECT 44.512 19.808 44.544 19.84 ;
  LAYER M2 ;
        RECT 46.88 19.744 46.912 19.776 ;
  LAYER M2 ;
        RECT 44.512 19.68 44.544 19.712 ;
  LAYER M2 ;
        RECT 46.88 19.616 46.912 19.648 ;
  LAYER M2 ;
        RECT 44.512 19.552 44.544 19.584 ;
  LAYER M2 ;
        RECT 46.88 19.488 46.912 19.52 ;
  LAYER M2 ;
        RECT 44.512 19.424 44.544 19.456 ;
  LAYER M2 ;
        RECT 46.88 19.36 46.912 19.392 ;
  LAYER M2 ;
        RECT 44.512 19.296 44.544 19.328 ;
  LAYER M2 ;
        RECT 46.88 19.232 46.912 19.264 ;
  LAYER M2 ;
        RECT 44.512 19.168 44.544 19.2 ;
  LAYER M2 ;
        RECT 46.88 19.104 46.912 19.136 ;
  LAYER M2 ;
        RECT 44.512 19.04 44.544 19.072 ;
  LAYER M2 ;
        RECT 46.88 18.976 46.912 19.008 ;
  LAYER M2 ;
        RECT 44.512 18.912 44.544 18.944 ;
  LAYER M2 ;
        RECT 46.88 18.848 46.912 18.88 ;
  LAYER M2 ;
        RECT 44.464 18.648 46.96 21.252 ;
  LAYER M1 ;
        RECT 44.512 15.588 44.544 18.096 ;
  LAYER M3 ;
        RECT 44.512 15.608 44.544 15.64 ;
  LAYER M1 ;
        RECT 44.576 15.588 44.608 18.096 ;
  LAYER M3 ;
        RECT 44.576 18.044 44.608 18.076 ;
  LAYER M1 ;
        RECT 44.64 15.588 44.672 18.096 ;
  LAYER M3 ;
        RECT 44.64 15.608 44.672 15.64 ;
  LAYER M1 ;
        RECT 44.704 15.588 44.736 18.096 ;
  LAYER M3 ;
        RECT 44.704 18.044 44.736 18.076 ;
  LAYER M1 ;
        RECT 44.768 15.588 44.8 18.096 ;
  LAYER M3 ;
        RECT 44.768 15.608 44.8 15.64 ;
  LAYER M1 ;
        RECT 44.832 15.588 44.864 18.096 ;
  LAYER M3 ;
        RECT 44.832 18.044 44.864 18.076 ;
  LAYER M1 ;
        RECT 44.896 15.588 44.928 18.096 ;
  LAYER M3 ;
        RECT 44.896 15.608 44.928 15.64 ;
  LAYER M1 ;
        RECT 44.96 15.588 44.992 18.096 ;
  LAYER M3 ;
        RECT 44.96 18.044 44.992 18.076 ;
  LAYER M1 ;
        RECT 45.024 15.588 45.056 18.096 ;
  LAYER M3 ;
        RECT 45.024 15.608 45.056 15.64 ;
  LAYER M1 ;
        RECT 45.088 15.588 45.12 18.096 ;
  LAYER M3 ;
        RECT 45.088 18.044 45.12 18.076 ;
  LAYER M1 ;
        RECT 45.152 15.588 45.184 18.096 ;
  LAYER M3 ;
        RECT 45.152 15.608 45.184 15.64 ;
  LAYER M1 ;
        RECT 45.216 15.588 45.248 18.096 ;
  LAYER M3 ;
        RECT 45.216 18.044 45.248 18.076 ;
  LAYER M1 ;
        RECT 45.28 15.588 45.312 18.096 ;
  LAYER M3 ;
        RECT 45.28 15.608 45.312 15.64 ;
  LAYER M1 ;
        RECT 45.344 15.588 45.376 18.096 ;
  LAYER M3 ;
        RECT 45.344 18.044 45.376 18.076 ;
  LAYER M1 ;
        RECT 45.408 15.588 45.44 18.096 ;
  LAYER M3 ;
        RECT 45.408 15.608 45.44 15.64 ;
  LAYER M1 ;
        RECT 45.472 15.588 45.504 18.096 ;
  LAYER M3 ;
        RECT 45.472 18.044 45.504 18.076 ;
  LAYER M1 ;
        RECT 45.536 15.588 45.568 18.096 ;
  LAYER M3 ;
        RECT 45.536 15.608 45.568 15.64 ;
  LAYER M1 ;
        RECT 45.6 15.588 45.632 18.096 ;
  LAYER M3 ;
        RECT 45.6 18.044 45.632 18.076 ;
  LAYER M1 ;
        RECT 45.664 15.588 45.696 18.096 ;
  LAYER M3 ;
        RECT 45.664 15.608 45.696 15.64 ;
  LAYER M1 ;
        RECT 45.728 15.588 45.76 18.096 ;
  LAYER M3 ;
        RECT 45.728 18.044 45.76 18.076 ;
  LAYER M1 ;
        RECT 45.792 15.588 45.824 18.096 ;
  LAYER M3 ;
        RECT 45.792 15.608 45.824 15.64 ;
  LAYER M1 ;
        RECT 45.856 15.588 45.888 18.096 ;
  LAYER M3 ;
        RECT 45.856 18.044 45.888 18.076 ;
  LAYER M1 ;
        RECT 45.92 15.588 45.952 18.096 ;
  LAYER M3 ;
        RECT 45.92 15.608 45.952 15.64 ;
  LAYER M1 ;
        RECT 45.984 15.588 46.016 18.096 ;
  LAYER M3 ;
        RECT 45.984 18.044 46.016 18.076 ;
  LAYER M1 ;
        RECT 46.048 15.588 46.08 18.096 ;
  LAYER M3 ;
        RECT 46.048 15.608 46.08 15.64 ;
  LAYER M1 ;
        RECT 46.112 15.588 46.144 18.096 ;
  LAYER M3 ;
        RECT 46.112 18.044 46.144 18.076 ;
  LAYER M1 ;
        RECT 46.176 15.588 46.208 18.096 ;
  LAYER M3 ;
        RECT 46.176 15.608 46.208 15.64 ;
  LAYER M1 ;
        RECT 46.24 15.588 46.272 18.096 ;
  LAYER M3 ;
        RECT 46.24 18.044 46.272 18.076 ;
  LAYER M1 ;
        RECT 46.304 15.588 46.336 18.096 ;
  LAYER M3 ;
        RECT 46.304 15.608 46.336 15.64 ;
  LAYER M1 ;
        RECT 46.368 15.588 46.4 18.096 ;
  LAYER M3 ;
        RECT 46.368 18.044 46.4 18.076 ;
  LAYER M1 ;
        RECT 46.432 15.588 46.464 18.096 ;
  LAYER M3 ;
        RECT 46.432 15.608 46.464 15.64 ;
  LAYER M1 ;
        RECT 46.496 15.588 46.528 18.096 ;
  LAYER M3 ;
        RECT 46.496 18.044 46.528 18.076 ;
  LAYER M1 ;
        RECT 46.56 15.588 46.592 18.096 ;
  LAYER M3 ;
        RECT 46.56 15.608 46.592 15.64 ;
  LAYER M1 ;
        RECT 46.624 15.588 46.656 18.096 ;
  LAYER M3 ;
        RECT 46.624 18.044 46.656 18.076 ;
  LAYER M1 ;
        RECT 46.688 15.588 46.72 18.096 ;
  LAYER M3 ;
        RECT 46.688 15.608 46.72 15.64 ;
  LAYER M1 ;
        RECT 46.752 15.588 46.784 18.096 ;
  LAYER M3 ;
        RECT 46.752 18.044 46.784 18.076 ;
  LAYER M1 ;
        RECT 46.816 15.588 46.848 18.096 ;
  LAYER M3 ;
        RECT 46.816 15.608 46.848 15.64 ;
  LAYER M1 ;
        RECT 46.88 15.588 46.912 18.096 ;
  LAYER M3 ;
        RECT 44.512 17.98 44.544 18.012 ;
  LAYER M2 ;
        RECT 46.88 17.916 46.912 17.948 ;
  LAYER M2 ;
        RECT 44.512 17.852 44.544 17.884 ;
  LAYER M2 ;
        RECT 46.88 17.788 46.912 17.82 ;
  LAYER M2 ;
        RECT 44.512 17.724 44.544 17.756 ;
  LAYER M2 ;
        RECT 46.88 17.66 46.912 17.692 ;
  LAYER M2 ;
        RECT 44.512 17.596 44.544 17.628 ;
  LAYER M2 ;
        RECT 46.88 17.532 46.912 17.564 ;
  LAYER M2 ;
        RECT 44.512 17.468 44.544 17.5 ;
  LAYER M2 ;
        RECT 46.88 17.404 46.912 17.436 ;
  LAYER M2 ;
        RECT 44.512 17.34 44.544 17.372 ;
  LAYER M2 ;
        RECT 46.88 17.276 46.912 17.308 ;
  LAYER M2 ;
        RECT 44.512 17.212 44.544 17.244 ;
  LAYER M2 ;
        RECT 46.88 17.148 46.912 17.18 ;
  LAYER M2 ;
        RECT 44.512 17.084 44.544 17.116 ;
  LAYER M2 ;
        RECT 46.88 17.02 46.912 17.052 ;
  LAYER M2 ;
        RECT 44.512 16.956 44.544 16.988 ;
  LAYER M2 ;
        RECT 46.88 16.892 46.912 16.924 ;
  LAYER M2 ;
        RECT 44.512 16.828 44.544 16.86 ;
  LAYER M2 ;
        RECT 46.88 16.764 46.912 16.796 ;
  LAYER M2 ;
        RECT 44.512 16.7 44.544 16.732 ;
  LAYER M2 ;
        RECT 46.88 16.636 46.912 16.668 ;
  LAYER M2 ;
        RECT 44.512 16.572 44.544 16.604 ;
  LAYER M2 ;
        RECT 46.88 16.508 46.912 16.54 ;
  LAYER M2 ;
        RECT 44.512 16.444 44.544 16.476 ;
  LAYER M2 ;
        RECT 46.88 16.38 46.912 16.412 ;
  LAYER M2 ;
        RECT 44.512 16.316 44.544 16.348 ;
  LAYER M2 ;
        RECT 46.88 16.252 46.912 16.284 ;
  LAYER M2 ;
        RECT 44.512 16.188 44.544 16.22 ;
  LAYER M2 ;
        RECT 46.88 16.124 46.912 16.156 ;
  LAYER M2 ;
        RECT 44.512 16.06 44.544 16.092 ;
  LAYER M2 ;
        RECT 46.88 15.996 46.912 16.028 ;
  LAYER M2 ;
        RECT 44.512 15.932 44.544 15.964 ;
  LAYER M2 ;
        RECT 46.88 15.868 46.912 15.9 ;
  LAYER M2 ;
        RECT 44.512 15.804 44.544 15.836 ;
  LAYER M2 ;
        RECT 46.88 15.74 46.912 15.772 ;
  LAYER M2 ;
        RECT 44.464 15.54 46.96 18.144 ;
  LAYER M1 ;
        RECT 22.56 12.816 22.592 12.888 ;
  LAYER M2 ;
        RECT 22.54 12.836 22.612 12.868 ;
  LAYER M2 ;
        RECT 22.576 12.836 25.328 12.868 ;
  LAYER M1 ;
        RECT 25.312 12.816 25.344 12.888 ;
  LAYER M2 ;
        RECT 25.292 12.836 25.364 12.868 ;
  LAYER M1 ;
        RECT 25.536 9.708 25.568 9.78 ;
  LAYER M2 ;
        RECT 25.516 9.728 25.588 9.76 ;
  LAYER M1 ;
        RECT 25.536 9.576 25.568 9.744 ;
  LAYER M1 ;
        RECT 25.536 9.54 25.568 9.612 ;
  LAYER M2 ;
        RECT 25.516 9.56 25.588 9.592 ;
  LAYER M2 ;
        RECT 25.328 9.56 25.552 9.592 ;
  LAYER M1 ;
        RECT 25.312 9.54 25.344 9.612 ;
  LAYER M2 ;
        RECT 25.292 9.56 25.364 9.592 ;
  LAYER M1 ;
        RECT 25.312 6.012 25.344 6.084 ;
  LAYER M2 ;
        RECT 25.292 6.032 25.364 6.064 ;
  LAYER M1 ;
        RECT 25.312 6.048 25.344 6.3 ;
  LAYER M1 ;
        RECT 25.312 6.3 25.344 12.852 ;
  LAYER M1 ;
        RECT 19.584 12.816 19.616 12.888 ;
  LAYER M2 ;
        RECT 19.564 12.836 19.636 12.868 ;
  LAYER M2 ;
        RECT 19.6 12.836 22.352 12.868 ;
  LAYER M1 ;
        RECT 22.336 12.816 22.368 12.888 ;
  LAYER M2 ;
        RECT 22.316 12.836 22.388 12.868 ;
  LAYER M1 ;
        RECT 22.336 6.012 22.368 6.084 ;
  LAYER M2 ;
        RECT 22.316 6.032 22.388 6.064 ;
  LAYER M1 ;
        RECT 22.336 6.048 22.368 6.3 ;
  LAYER M1 ;
        RECT 22.336 6.3 22.368 12.852 ;
  LAYER M2 ;
        RECT 22.352 6.032 25.328 6.064 ;
  LAYER M1 ;
        RECT 25.536 12.816 25.568 12.888 ;
  LAYER M2 ;
        RECT 25.516 12.836 25.588 12.868 ;
  LAYER M2 ;
        RECT 25.552 12.836 28.304 12.868 ;
  LAYER M1 ;
        RECT 28.288 12.816 28.32 12.888 ;
  LAYER M2 ;
        RECT 28.268 12.836 28.34 12.868 ;
  LAYER M1 ;
        RECT 28.288 5.844 28.32 5.916 ;
  LAYER M2 ;
        RECT 28.268 5.864 28.34 5.896 ;
  LAYER M1 ;
        RECT 28.288 5.88 28.32 6.3 ;
  LAYER M1 ;
        RECT 28.288 6.3 28.32 12.852 ;
  LAYER M1 ;
        RECT 19.584 9.708 19.616 9.78 ;
  LAYER M2 ;
        RECT 19.564 9.728 19.636 9.76 ;
  LAYER M1 ;
        RECT 19.584 9.576 19.616 9.744 ;
  LAYER M1 ;
        RECT 19.584 9.54 19.616 9.612 ;
  LAYER M2 ;
        RECT 19.564 9.56 19.636 9.592 ;
  LAYER M2 ;
        RECT 19.376 9.56 19.6 9.592 ;
  LAYER M1 ;
        RECT 19.36 9.54 19.392 9.612 ;
  LAYER M2 ;
        RECT 19.34 9.56 19.412 9.592 ;
  LAYER M1 ;
        RECT 19.36 5.844 19.392 5.916 ;
  LAYER M2 ;
        RECT 19.34 5.864 19.412 5.896 ;
  LAYER M1 ;
        RECT 19.36 5.88 19.392 6.3 ;
  LAYER M1 ;
        RECT 19.36 6.3 19.392 9.576 ;
  LAYER M2 ;
        RECT 19.376 5.864 28.304 5.896 ;
  LAYER M1 ;
        RECT 22.56 9.708 22.592 9.78 ;
  LAYER M2 ;
        RECT 22.54 9.728 22.612 9.76 ;
  LAYER M2 ;
        RECT 19.6 9.728 22.576 9.76 ;
  LAYER M1 ;
        RECT 19.584 9.708 19.616 9.78 ;
  LAYER M2 ;
        RECT 19.564 9.728 19.636 9.76 ;
  LAYER M1 ;
        RECT 28.512 6.6 28.544 6.672 ;
  LAYER M2 ;
        RECT 28.492 6.62 28.564 6.652 ;
  LAYER M2 ;
        RECT 28.528 6.62 31.28 6.652 ;
  LAYER M1 ;
        RECT 31.264 6.6 31.296 6.672 ;
  LAYER M2 ;
        RECT 31.244 6.62 31.316 6.652 ;
  LAYER M1 ;
        RECT 28.512 9.708 28.544 9.78 ;
  LAYER M2 ;
        RECT 28.492 9.728 28.564 9.76 ;
  LAYER M2 ;
        RECT 28.528 9.728 31.28 9.76 ;
  LAYER M1 ;
        RECT 31.264 9.708 31.296 9.78 ;
  LAYER M2 ;
        RECT 31.244 9.728 31.316 9.76 ;
  LAYER M1 ;
        RECT 28.512 12.816 28.544 12.888 ;
  LAYER M2 ;
        RECT 28.492 12.836 28.564 12.868 ;
  LAYER M2 ;
        RECT 28.528 12.836 31.28 12.868 ;
  LAYER M1 ;
        RECT 31.264 12.816 31.296 12.888 ;
  LAYER M2 ;
        RECT 31.244 12.836 31.316 12.868 ;
  LAYER M1 ;
        RECT 28.512 15.924 28.544 15.996 ;
  LAYER M2 ;
        RECT 28.492 15.944 28.564 15.976 ;
  LAYER M2 ;
        RECT 28.528 15.944 31.28 15.976 ;
  LAYER M1 ;
        RECT 31.264 15.924 31.296 15.996 ;
  LAYER M2 ;
        RECT 31.244 15.944 31.316 15.976 ;
  LAYER M1 ;
        RECT 31.264 5.676 31.296 5.748 ;
  LAYER M2 ;
        RECT 31.244 5.696 31.316 5.728 ;
  LAYER M1 ;
        RECT 31.264 5.712 31.296 6.3 ;
  LAYER M1 ;
        RECT 31.264 6.3 31.296 15.96 ;
  LAYER M1 ;
        RECT 16.608 6.6 16.64 6.672 ;
  LAYER M2 ;
        RECT 16.588 6.62 16.66 6.652 ;
  LAYER M1 ;
        RECT 16.608 6.468 16.64 6.636 ;
  LAYER M1 ;
        RECT 16.608 6.432 16.64 6.504 ;
  LAYER M2 ;
        RECT 16.588 6.452 16.66 6.484 ;
  LAYER M2 ;
        RECT 16.4 6.452 16.624 6.484 ;
  LAYER M1 ;
        RECT 16.384 6.432 16.416 6.504 ;
  LAYER M2 ;
        RECT 16.364 6.452 16.436 6.484 ;
  LAYER M1 ;
        RECT 16.608 9.708 16.64 9.78 ;
  LAYER M2 ;
        RECT 16.588 9.728 16.66 9.76 ;
  LAYER M1 ;
        RECT 16.608 9.576 16.64 9.744 ;
  LAYER M1 ;
        RECT 16.608 9.54 16.64 9.612 ;
  LAYER M2 ;
        RECT 16.588 9.56 16.66 9.592 ;
  LAYER M2 ;
        RECT 16.4 9.56 16.624 9.592 ;
  LAYER M1 ;
        RECT 16.384 9.54 16.416 9.612 ;
  LAYER M2 ;
        RECT 16.364 9.56 16.436 9.592 ;
  LAYER M1 ;
        RECT 16.608 12.816 16.64 12.888 ;
  LAYER M2 ;
        RECT 16.588 12.836 16.66 12.868 ;
  LAYER M1 ;
        RECT 16.608 12.684 16.64 12.852 ;
  LAYER M1 ;
        RECT 16.608 12.648 16.64 12.72 ;
  LAYER M2 ;
        RECT 16.588 12.668 16.66 12.7 ;
  LAYER M2 ;
        RECT 16.4 12.668 16.624 12.7 ;
  LAYER M1 ;
        RECT 16.384 12.648 16.416 12.72 ;
  LAYER M2 ;
        RECT 16.364 12.668 16.436 12.7 ;
  LAYER M1 ;
        RECT 16.608 15.924 16.64 15.996 ;
  LAYER M2 ;
        RECT 16.588 15.944 16.66 15.976 ;
  LAYER M1 ;
        RECT 16.608 15.792 16.64 15.96 ;
  LAYER M1 ;
        RECT 16.608 15.756 16.64 15.828 ;
  LAYER M2 ;
        RECT 16.588 15.776 16.66 15.808 ;
  LAYER M2 ;
        RECT 16.4 15.776 16.624 15.808 ;
  LAYER M1 ;
        RECT 16.384 15.756 16.416 15.828 ;
  LAYER M2 ;
        RECT 16.364 15.776 16.436 15.808 ;
  LAYER M1 ;
        RECT 16.384 5.676 16.416 5.748 ;
  LAYER M2 ;
        RECT 16.364 5.696 16.436 5.728 ;
  LAYER M1 ;
        RECT 16.384 5.712 16.416 6.3 ;
  LAYER M1 ;
        RECT 16.384 6.3 16.416 15.792 ;
  LAYER M2 ;
        RECT 16.4 5.696 31.28 5.728 ;
  LAYER M1 ;
        RECT 25.536 6.6 25.568 6.672 ;
  LAYER M2 ;
        RECT 25.516 6.62 25.588 6.652 ;
  LAYER M2 ;
        RECT 25.552 6.62 28.528 6.652 ;
  LAYER M1 ;
        RECT 28.512 6.6 28.544 6.672 ;
  LAYER M2 ;
        RECT 28.492 6.62 28.564 6.652 ;
  LAYER M1 ;
        RECT 25.536 15.924 25.568 15.996 ;
  LAYER M2 ;
        RECT 25.516 15.944 25.588 15.976 ;
  LAYER M2 ;
        RECT 25.552 15.944 28.528 15.976 ;
  LAYER M1 ;
        RECT 28.512 15.924 28.544 15.996 ;
  LAYER M2 ;
        RECT 28.492 15.944 28.564 15.976 ;
  LAYER M1 ;
        RECT 22.56 15.924 22.592 15.996 ;
  LAYER M2 ;
        RECT 22.54 15.944 22.612 15.976 ;
  LAYER M2 ;
        RECT 22.576 15.944 25.552 15.976 ;
  LAYER M1 ;
        RECT 25.536 15.924 25.568 15.996 ;
  LAYER M2 ;
        RECT 25.516 15.944 25.588 15.976 ;
  LAYER M1 ;
        RECT 19.584 15.924 19.616 15.996 ;
  LAYER M2 ;
        RECT 19.564 15.944 19.636 15.976 ;
  LAYER M2 ;
        RECT 19.6 15.944 22.576 15.976 ;
  LAYER M1 ;
        RECT 22.56 15.924 22.592 15.996 ;
  LAYER M2 ;
        RECT 22.54 15.944 22.612 15.976 ;
  LAYER M1 ;
        RECT 19.584 6.6 19.616 6.672 ;
  LAYER M2 ;
        RECT 19.564 6.62 19.636 6.652 ;
  LAYER M2 ;
        RECT 16.624 6.62 19.6 6.652 ;
  LAYER M1 ;
        RECT 16.608 6.6 16.64 6.672 ;
  LAYER M2 ;
        RECT 16.588 6.62 16.66 6.652 ;
  LAYER M1 ;
        RECT 22.56 6.6 22.592 6.672 ;
  LAYER M2 ;
        RECT 22.54 6.62 22.612 6.652 ;
  LAYER M2 ;
        RECT 19.6 6.62 22.576 6.652 ;
  LAYER M1 ;
        RECT 19.584 6.6 19.616 6.672 ;
  LAYER M2 ;
        RECT 19.564 6.62 19.636 6.652 ;
  LAYER M1 ;
        RECT 24.928 15.252 24.96 15.324 ;
  LAYER M2 ;
        RECT 24.908 15.272 24.98 15.304 ;
  LAYER M2 ;
        RECT 24.944 15.272 25.168 15.304 ;
  LAYER M1 ;
        RECT 25.152 15.252 25.184 15.324 ;
  LAYER M2 ;
        RECT 25.132 15.272 25.204 15.304 ;
  LAYER M1 ;
        RECT 27.904 12.144 27.936 12.216 ;
  LAYER M2 ;
        RECT 27.884 12.164 27.956 12.196 ;
  LAYER M1 ;
        RECT 27.904 12.18 27.936 12.348 ;
  LAYER M1 ;
        RECT 27.904 12.312 27.936 12.384 ;
  LAYER M2 ;
        RECT 27.884 12.332 27.956 12.364 ;
  LAYER M2 ;
        RECT 25.168 12.332 27.92 12.364 ;
  LAYER M1 ;
        RECT 25.152 12.312 25.184 12.384 ;
  LAYER M2 ;
        RECT 25.132 12.332 25.204 12.364 ;
  LAYER M1 ;
        RECT 25.152 18.948 25.184 19.02 ;
  LAYER M2 ;
        RECT 25.132 18.968 25.204 19 ;
  LAYER M1 ;
        RECT 25.152 18.732 25.184 18.984 ;
  LAYER M1 ;
        RECT 25.152 12.348 25.184 18.732 ;
  LAYER M1 ;
        RECT 21.952 15.252 21.984 15.324 ;
  LAYER M2 ;
        RECT 21.932 15.272 22.004 15.304 ;
  LAYER M2 ;
        RECT 21.968 15.272 22.192 15.304 ;
  LAYER M1 ;
        RECT 22.176 15.252 22.208 15.324 ;
  LAYER M2 ;
        RECT 22.156 15.272 22.228 15.304 ;
  LAYER M1 ;
        RECT 22.176 18.948 22.208 19.02 ;
  LAYER M2 ;
        RECT 22.156 18.968 22.228 19 ;
  LAYER M1 ;
        RECT 22.176 18.732 22.208 18.984 ;
  LAYER M1 ;
        RECT 22.176 15.288 22.208 18.732 ;
  LAYER M2 ;
        RECT 22.192 18.968 25.168 19 ;
  LAYER M1 ;
        RECT 27.904 15.252 27.936 15.324 ;
  LAYER M2 ;
        RECT 27.884 15.272 27.956 15.304 ;
  LAYER M2 ;
        RECT 27.92 15.272 28.144 15.304 ;
  LAYER M1 ;
        RECT 28.128 15.252 28.16 15.324 ;
  LAYER M2 ;
        RECT 28.108 15.272 28.18 15.304 ;
  LAYER M1 ;
        RECT 28.128 19.116 28.16 19.188 ;
  LAYER M2 ;
        RECT 28.108 19.136 28.18 19.168 ;
  LAYER M1 ;
        RECT 28.128 18.732 28.16 19.152 ;
  LAYER M1 ;
        RECT 28.128 15.288 28.16 18.732 ;
  LAYER M1 ;
        RECT 21.952 12.144 21.984 12.216 ;
  LAYER M2 ;
        RECT 21.932 12.164 22.004 12.196 ;
  LAYER M1 ;
        RECT 21.952 12.18 21.984 12.348 ;
  LAYER M1 ;
        RECT 21.952 12.312 21.984 12.384 ;
  LAYER M2 ;
        RECT 21.932 12.332 22.004 12.364 ;
  LAYER M2 ;
        RECT 19.216 12.332 21.968 12.364 ;
  LAYER M1 ;
        RECT 19.2 12.312 19.232 12.384 ;
  LAYER M2 ;
        RECT 19.18 12.332 19.252 12.364 ;
  LAYER M1 ;
        RECT 19.2 19.116 19.232 19.188 ;
  LAYER M2 ;
        RECT 19.18 19.136 19.252 19.168 ;
  LAYER M1 ;
        RECT 19.2 18.732 19.232 19.152 ;
  LAYER M1 ;
        RECT 19.2 12.348 19.232 18.732 ;
  LAYER M2 ;
        RECT 19.216 19.136 28.144 19.168 ;
  LAYER M1 ;
        RECT 24.928 12.144 24.96 12.216 ;
  LAYER M2 ;
        RECT 24.908 12.164 24.98 12.196 ;
  LAYER M2 ;
        RECT 21.968 12.164 24.944 12.196 ;
  LAYER M1 ;
        RECT 21.952 12.144 21.984 12.216 ;
  LAYER M2 ;
        RECT 21.932 12.164 22.004 12.196 ;
  LAYER M1 ;
        RECT 30.88 9.036 30.912 9.108 ;
  LAYER M2 ;
        RECT 30.86 9.056 30.932 9.088 ;
  LAYER M2 ;
        RECT 30.896 9.056 31.12 9.088 ;
  LAYER M1 ;
        RECT 31.104 9.036 31.136 9.108 ;
  LAYER M2 ;
        RECT 31.084 9.056 31.156 9.088 ;
  LAYER M1 ;
        RECT 30.88 12.144 30.912 12.216 ;
  LAYER M2 ;
        RECT 30.86 12.164 30.932 12.196 ;
  LAYER M2 ;
        RECT 30.896 12.164 31.12 12.196 ;
  LAYER M1 ;
        RECT 31.104 12.144 31.136 12.216 ;
  LAYER M2 ;
        RECT 31.084 12.164 31.156 12.196 ;
  LAYER M1 ;
        RECT 30.88 15.252 30.912 15.324 ;
  LAYER M2 ;
        RECT 30.86 15.272 30.932 15.304 ;
  LAYER M2 ;
        RECT 30.896 15.272 31.12 15.304 ;
  LAYER M1 ;
        RECT 31.104 15.252 31.136 15.324 ;
  LAYER M2 ;
        RECT 31.084 15.272 31.156 15.304 ;
  LAYER M1 ;
        RECT 30.88 18.36 30.912 18.432 ;
  LAYER M2 ;
        RECT 30.86 18.38 30.932 18.412 ;
  LAYER M2 ;
        RECT 30.896 18.38 31.12 18.412 ;
  LAYER M1 ;
        RECT 31.104 18.36 31.136 18.432 ;
  LAYER M2 ;
        RECT 31.084 18.38 31.156 18.412 ;
  LAYER M1 ;
        RECT 31.104 19.284 31.136 19.356 ;
  LAYER M2 ;
        RECT 31.084 19.304 31.156 19.336 ;
  LAYER M1 ;
        RECT 31.104 18.732 31.136 19.32 ;
  LAYER M1 ;
        RECT 31.104 9.072 31.136 18.732 ;
  LAYER M1 ;
        RECT 18.976 9.036 19.008 9.108 ;
  LAYER M2 ;
        RECT 18.956 9.056 19.028 9.088 ;
  LAYER M1 ;
        RECT 18.976 9.072 19.008 9.24 ;
  LAYER M1 ;
        RECT 18.976 9.204 19.008 9.276 ;
  LAYER M2 ;
        RECT 18.956 9.224 19.028 9.256 ;
  LAYER M2 ;
        RECT 16.24 9.224 18.992 9.256 ;
  LAYER M1 ;
        RECT 16.224 9.204 16.256 9.276 ;
  LAYER M2 ;
        RECT 16.204 9.224 16.276 9.256 ;
  LAYER M1 ;
        RECT 18.976 12.144 19.008 12.216 ;
  LAYER M2 ;
        RECT 18.956 12.164 19.028 12.196 ;
  LAYER M1 ;
        RECT 18.976 12.18 19.008 12.348 ;
  LAYER M1 ;
        RECT 18.976 12.312 19.008 12.384 ;
  LAYER M2 ;
        RECT 18.956 12.332 19.028 12.364 ;
  LAYER M2 ;
        RECT 16.24 12.332 18.992 12.364 ;
  LAYER M1 ;
        RECT 16.224 12.312 16.256 12.384 ;
  LAYER M2 ;
        RECT 16.204 12.332 16.276 12.364 ;
  LAYER M1 ;
        RECT 18.976 15.252 19.008 15.324 ;
  LAYER M2 ;
        RECT 18.956 15.272 19.028 15.304 ;
  LAYER M1 ;
        RECT 18.976 15.288 19.008 15.456 ;
  LAYER M1 ;
        RECT 18.976 15.42 19.008 15.492 ;
  LAYER M2 ;
        RECT 18.956 15.44 19.028 15.472 ;
  LAYER M2 ;
        RECT 16.24 15.44 18.992 15.472 ;
  LAYER M1 ;
        RECT 16.224 15.42 16.256 15.492 ;
  LAYER M2 ;
        RECT 16.204 15.44 16.276 15.472 ;
  LAYER M1 ;
        RECT 18.976 18.36 19.008 18.432 ;
  LAYER M2 ;
        RECT 18.956 18.38 19.028 18.412 ;
  LAYER M1 ;
        RECT 18.976 18.396 19.008 18.564 ;
  LAYER M1 ;
        RECT 18.976 18.528 19.008 18.6 ;
  LAYER M2 ;
        RECT 18.956 18.548 19.028 18.58 ;
  LAYER M2 ;
        RECT 16.24 18.548 18.992 18.58 ;
  LAYER M1 ;
        RECT 16.224 18.528 16.256 18.6 ;
  LAYER M2 ;
        RECT 16.204 18.548 16.276 18.58 ;
  LAYER M1 ;
        RECT 16.224 19.284 16.256 19.356 ;
  LAYER M2 ;
        RECT 16.204 19.304 16.276 19.336 ;
  LAYER M1 ;
        RECT 16.224 18.732 16.256 19.32 ;
  LAYER M1 ;
        RECT 16.224 9.24 16.256 18.732 ;
  LAYER M2 ;
        RECT 16.24 19.304 31.12 19.336 ;
  LAYER M1 ;
        RECT 27.904 9.036 27.936 9.108 ;
  LAYER M2 ;
        RECT 27.884 9.056 27.956 9.088 ;
  LAYER M2 ;
        RECT 27.92 9.056 30.896 9.088 ;
  LAYER M1 ;
        RECT 30.88 9.036 30.912 9.108 ;
  LAYER M2 ;
        RECT 30.86 9.056 30.932 9.088 ;
  LAYER M1 ;
        RECT 27.904 18.36 27.936 18.432 ;
  LAYER M2 ;
        RECT 27.884 18.38 27.956 18.412 ;
  LAYER M2 ;
        RECT 27.92 18.38 30.896 18.412 ;
  LAYER M1 ;
        RECT 30.88 18.36 30.912 18.432 ;
  LAYER M2 ;
        RECT 30.86 18.38 30.932 18.412 ;
  LAYER M1 ;
        RECT 24.928 18.36 24.96 18.432 ;
  LAYER M2 ;
        RECT 24.908 18.38 24.98 18.412 ;
  LAYER M2 ;
        RECT 24.944 18.38 27.92 18.412 ;
  LAYER M1 ;
        RECT 27.904 18.36 27.936 18.432 ;
  LAYER M2 ;
        RECT 27.884 18.38 27.956 18.412 ;
  LAYER M1 ;
        RECT 21.952 18.36 21.984 18.432 ;
  LAYER M2 ;
        RECT 21.932 18.38 22.004 18.412 ;
  LAYER M2 ;
        RECT 21.968 18.38 24.944 18.412 ;
  LAYER M1 ;
        RECT 24.928 18.36 24.96 18.432 ;
  LAYER M2 ;
        RECT 24.908 18.38 24.98 18.412 ;
  LAYER M1 ;
        RECT 21.952 9.036 21.984 9.108 ;
  LAYER M2 ;
        RECT 21.932 9.056 22.004 9.088 ;
  LAYER M2 ;
        RECT 18.992 9.056 21.968 9.088 ;
  LAYER M1 ;
        RECT 18.976 9.036 19.008 9.108 ;
  LAYER M2 ;
        RECT 18.956 9.056 19.028 9.088 ;
  LAYER M1 ;
        RECT 24.928 9.036 24.96 9.108 ;
  LAYER M2 ;
        RECT 24.908 9.056 24.98 9.088 ;
  LAYER M2 ;
        RECT 21.968 9.056 24.944 9.088 ;
  LAYER M1 ;
        RECT 21.952 9.036 21.984 9.108 ;
  LAYER M2 ;
        RECT 21.932 9.056 22.004 9.088 ;
  LAYER M1 ;
        RECT 30.88 6.6 30.912 9.108 ;
  LAYER M3 ;
        RECT 30.88 9.056 30.912 9.088 ;
  LAYER M1 ;
        RECT 30.816 6.6 30.848 9.108 ;
  LAYER M3 ;
        RECT 30.816 6.62 30.848 6.652 ;
  LAYER M1 ;
        RECT 30.752 6.6 30.784 9.108 ;
  LAYER M3 ;
        RECT 30.752 9.056 30.784 9.088 ;
  LAYER M1 ;
        RECT 30.688 6.6 30.72 9.108 ;
  LAYER M3 ;
        RECT 30.688 6.62 30.72 6.652 ;
  LAYER M1 ;
        RECT 30.624 6.6 30.656 9.108 ;
  LAYER M3 ;
        RECT 30.624 9.056 30.656 9.088 ;
  LAYER M1 ;
        RECT 30.56 6.6 30.592 9.108 ;
  LAYER M3 ;
        RECT 30.56 6.62 30.592 6.652 ;
  LAYER M1 ;
        RECT 30.496 6.6 30.528 9.108 ;
  LAYER M3 ;
        RECT 30.496 9.056 30.528 9.088 ;
  LAYER M1 ;
        RECT 30.432 6.6 30.464 9.108 ;
  LAYER M3 ;
        RECT 30.432 6.62 30.464 6.652 ;
  LAYER M1 ;
        RECT 30.368 6.6 30.4 9.108 ;
  LAYER M3 ;
        RECT 30.368 9.056 30.4 9.088 ;
  LAYER M1 ;
        RECT 30.304 6.6 30.336 9.108 ;
  LAYER M3 ;
        RECT 30.304 6.62 30.336 6.652 ;
  LAYER M1 ;
        RECT 30.24 6.6 30.272 9.108 ;
  LAYER M3 ;
        RECT 30.24 9.056 30.272 9.088 ;
  LAYER M1 ;
        RECT 30.176 6.6 30.208 9.108 ;
  LAYER M3 ;
        RECT 30.176 6.62 30.208 6.652 ;
  LAYER M1 ;
        RECT 30.112 6.6 30.144 9.108 ;
  LAYER M3 ;
        RECT 30.112 9.056 30.144 9.088 ;
  LAYER M1 ;
        RECT 30.048 6.6 30.08 9.108 ;
  LAYER M3 ;
        RECT 30.048 6.62 30.08 6.652 ;
  LAYER M1 ;
        RECT 29.984 6.6 30.016 9.108 ;
  LAYER M3 ;
        RECT 29.984 9.056 30.016 9.088 ;
  LAYER M1 ;
        RECT 29.92 6.6 29.952 9.108 ;
  LAYER M3 ;
        RECT 29.92 6.62 29.952 6.652 ;
  LAYER M1 ;
        RECT 29.856 6.6 29.888 9.108 ;
  LAYER M3 ;
        RECT 29.856 9.056 29.888 9.088 ;
  LAYER M1 ;
        RECT 29.792 6.6 29.824 9.108 ;
  LAYER M3 ;
        RECT 29.792 6.62 29.824 6.652 ;
  LAYER M1 ;
        RECT 29.728 6.6 29.76 9.108 ;
  LAYER M3 ;
        RECT 29.728 9.056 29.76 9.088 ;
  LAYER M1 ;
        RECT 29.664 6.6 29.696 9.108 ;
  LAYER M3 ;
        RECT 29.664 6.62 29.696 6.652 ;
  LAYER M1 ;
        RECT 29.6 6.6 29.632 9.108 ;
  LAYER M3 ;
        RECT 29.6 9.056 29.632 9.088 ;
  LAYER M1 ;
        RECT 29.536 6.6 29.568 9.108 ;
  LAYER M3 ;
        RECT 29.536 6.62 29.568 6.652 ;
  LAYER M1 ;
        RECT 29.472 6.6 29.504 9.108 ;
  LAYER M3 ;
        RECT 29.472 9.056 29.504 9.088 ;
  LAYER M1 ;
        RECT 29.408 6.6 29.44 9.108 ;
  LAYER M3 ;
        RECT 29.408 6.62 29.44 6.652 ;
  LAYER M1 ;
        RECT 29.344 6.6 29.376 9.108 ;
  LAYER M3 ;
        RECT 29.344 9.056 29.376 9.088 ;
  LAYER M1 ;
        RECT 29.28 6.6 29.312 9.108 ;
  LAYER M3 ;
        RECT 29.28 6.62 29.312 6.652 ;
  LAYER M1 ;
        RECT 29.216 6.6 29.248 9.108 ;
  LAYER M3 ;
        RECT 29.216 9.056 29.248 9.088 ;
  LAYER M1 ;
        RECT 29.152 6.6 29.184 9.108 ;
  LAYER M3 ;
        RECT 29.152 6.62 29.184 6.652 ;
  LAYER M1 ;
        RECT 29.088 6.6 29.12 9.108 ;
  LAYER M3 ;
        RECT 29.088 9.056 29.12 9.088 ;
  LAYER M1 ;
        RECT 29.024 6.6 29.056 9.108 ;
  LAYER M3 ;
        RECT 29.024 6.62 29.056 6.652 ;
  LAYER M1 ;
        RECT 28.96 6.6 28.992 9.108 ;
  LAYER M3 ;
        RECT 28.96 9.056 28.992 9.088 ;
  LAYER M1 ;
        RECT 28.896 6.6 28.928 9.108 ;
  LAYER M3 ;
        RECT 28.896 6.62 28.928 6.652 ;
  LAYER M1 ;
        RECT 28.832 6.6 28.864 9.108 ;
  LAYER M3 ;
        RECT 28.832 9.056 28.864 9.088 ;
  LAYER M1 ;
        RECT 28.768 6.6 28.8 9.108 ;
  LAYER M3 ;
        RECT 28.768 6.62 28.8 6.652 ;
  LAYER M1 ;
        RECT 28.704 6.6 28.736 9.108 ;
  LAYER M3 ;
        RECT 28.704 9.056 28.736 9.088 ;
  LAYER M1 ;
        RECT 28.64 6.6 28.672 9.108 ;
  LAYER M3 ;
        RECT 28.64 6.62 28.672 6.652 ;
  LAYER M1 ;
        RECT 28.576 6.6 28.608 9.108 ;
  LAYER M3 ;
        RECT 28.576 9.056 28.608 9.088 ;
  LAYER M1 ;
        RECT 28.512 6.6 28.544 9.108 ;
  LAYER M3 ;
        RECT 30.88 6.684 30.912 6.716 ;
  LAYER M2 ;
        RECT 28.512 6.748 28.544 6.78 ;
  LAYER M2 ;
        RECT 30.88 6.812 30.912 6.844 ;
  LAYER M2 ;
        RECT 28.512 6.876 28.544 6.908 ;
  LAYER M2 ;
        RECT 30.88 6.94 30.912 6.972 ;
  LAYER M2 ;
        RECT 28.512 7.004 28.544 7.036 ;
  LAYER M2 ;
        RECT 30.88 7.068 30.912 7.1 ;
  LAYER M2 ;
        RECT 28.512 7.132 28.544 7.164 ;
  LAYER M2 ;
        RECT 30.88 7.196 30.912 7.228 ;
  LAYER M2 ;
        RECT 28.512 7.26 28.544 7.292 ;
  LAYER M2 ;
        RECT 30.88 7.324 30.912 7.356 ;
  LAYER M2 ;
        RECT 28.512 7.388 28.544 7.42 ;
  LAYER M2 ;
        RECT 30.88 7.452 30.912 7.484 ;
  LAYER M2 ;
        RECT 28.512 7.516 28.544 7.548 ;
  LAYER M2 ;
        RECT 30.88 7.58 30.912 7.612 ;
  LAYER M2 ;
        RECT 28.512 7.644 28.544 7.676 ;
  LAYER M2 ;
        RECT 30.88 7.708 30.912 7.74 ;
  LAYER M2 ;
        RECT 28.512 7.772 28.544 7.804 ;
  LAYER M2 ;
        RECT 30.88 7.836 30.912 7.868 ;
  LAYER M2 ;
        RECT 28.512 7.9 28.544 7.932 ;
  LAYER M2 ;
        RECT 30.88 7.964 30.912 7.996 ;
  LAYER M2 ;
        RECT 28.512 8.028 28.544 8.06 ;
  LAYER M2 ;
        RECT 30.88 8.092 30.912 8.124 ;
  LAYER M2 ;
        RECT 28.512 8.156 28.544 8.188 ;
  LAYER M2 ;
        RECT 30.88 8.22 30.912 8.252 ;
  LAYER M2 ;
        RECT 28.512 8.284 28.544 8.316 ;
  LAYER M2 ;
        RECT 30.88 8.348 30.912 8.38 ;
  LAYER M2 ;
        RECT 28.512 8.412 28.544 8.444 ;
  LAYER M2 ;
        RECT 30.88 8.476 30.912 8.508 ;
  LAYER M2 ;
        RECT 28.512 8.54 28.544 8.572 ;
  LAYER M2 ;
        RECT 30.88 8.604 30.912 8.636 ;
  LAYER M2 ;
        RECT 28.512 8.668 28.544 8.7 ;
  LAYER M2 ;
        RECT 30.88 8.732 30.912 8.764 ;
  LAYER M2 ;
        RECT 28.512 8.796 28.544 8.828 ;
  LAYER M2 ;
        RECT 30.88 8.86 30.912 8.892 ;
  LAYER M2 ;
        RECT 28.512 8.924 28.544 8.956 ;
  LAYER M2 ;
        RECT 28.464 6.552 30.96 9.156 ;
  LAYER M1 ;
        RECT 30.88 9.708 30.912 12.216 ;
  LAYER M3 ;
        RECT 30.88 12.164 30.912 12.196 ;
  LAYER M1 ;
        RECT 30.816 9.708 30.848 12.216 ;
  LAYER M3 ;
        RECT 30.816 9.728 30.848 9.76 ;
  LAYER M1 ;
        RECT 30.752 9.708 30.784 12.216 ;
  LAYER M3 ;
        RECT 30.752 12.164 30.784 12.196 ;
  LAYER M1 ;
        RECT 30.688 9.708 30.72 12.216 ;
  LAYER M3 ;
        RECT 30.688 9.728 30.72 9.76 ;
  LAYER M1 ;
        RECT 30.624 9.708 30.656 12.216 ;
  LAYER M3 ;
        RECT 30.624 12.164 30.656 12.196 ;
  LAYER M1 ;
        RECT 30.56 9.708 30.592 12.216 ;
  LAYER M3 ;
        RECT 30.56 9.728 30.592 9.76 ;
  LAYER M1 ;
        RECT 30.496 9.708 30.528 12.216 ;
  LAYER M3 ;
        RECT 30.496 12.164 30.528 12.196 ;
  LAYER M1 ;
        RECT 30.432 9.708 30.464 12.216 ;
  LAYER M3 ;
        RECT 30.432 9.728 30.464 9.76 ;
  LAYER M1 ;
        RECT 30.368 9.708 30.4 12.216 ;
  LAYER M3 ;
        RECT 30.368 12.164 30.4 12.196 ;
  LAYER M1 ;
        RECT 30.304 9.708 30.336 12.216 ;
  LAYER M3 ;
        RECT 30.304 9.728 30.336 9.76 ;
  LAYER M1 ;
        RECT 30.24 9.708 30.272 12.216 ;
  LAYER M3 ;
        RECT 30.24 12.164 30.272 12.196 ;
  LAYER M1 ;
        RECT 30.176 9.708 30.208 12.216 ;
  LAYER M3 ;
        RECT 30.176 9.728 30.208 9.76 ;
  LAYER M1 ;
        RECT 30.112 9.708 30.144 12.216 ;
  LAYER M3 ;
        RECT 30.112 12.164 30.144 12.196 ;
  LAYER M1 ;
        RECT 30.048 9.708 30.08 12.216 ;
  LAYER M3 ;
        RECT 30.048 9.728 30.08 9.76 ;
  LAYER M1 ;
        RECT 29.984 9.708 30.016 12.216 ;
  LAYER M3 ;
        RECT 29.984 12.164 30.016 12.196 ;
  LAYER M1 ;
        RECT 29.92 9.708 29.952 12.216 ;
  LAYER M3 ;
        RECT 29.92 9.728 29.952 9.76 ;
  LAYER M1 ;
        RECT 29.856 9.708 29.888 12.216 ;
  LAYER M3 ;
        RECT 29.856 12.164 29.888 12.196 ;
  LAYER M1 ;
        RECT 29.792 9.708 29.824 12.216 ;
  LAYER M3 ;
        RECT 29.792 9.728 29.824 9.76 ;
  LAYER M1 ;
        RECT 29.728 9.708 29.76 12.216 ;
  LAYER M3 ;
        RECT 29.728 12.164 29.76 12.196 ;
  LAYER M1 ;
        RECT 29.664 9.708 29.696 12.216 ;
  LAYER M3 ;
        RECT 29.664 9.728 29.696 9.76 ;
  LAYER M1 ;
        RECT 29.6 9.708 29.632 12.216 ;
  LAYER M3 ;
        RECT 29.6 12.164 29.632 12.196 ;
  LAYER M1 ;
        RECT 29.536 9.708 29.568 12.216 ;
  LAYER M3 ;
        RECT 29.536 9.728 29.568 9.76 ;
  LAYER M1 ;
        RECT 29.472 9.708 29.504 12.216 ;
  LAYER M3 ;
        RECT 29.472 12.164 29.504 12.196 ;
  LAYER M1 ;
        RECT 29.408 9.708 29.44 12.216 ;
  LAYER M3 ;
        RECT 29.408 9.728 29.44 9.76 ;
  LAYER M1 ;
        RECT 29.344 9.708 29.376 12.216 ;
  LAYER M3 ;
        RECT 29.344 12.164 29.376 12.196 ;
  LAYER M1 ;
        RECT 29.28 9.708 29.312 12.216 ;
  LAYER M3 ;
        RECT 29.28 9.728 29.312 9.76 ;
  LAYER M1 ;
        RECT 29.216 9.708 29.248 12.216 ;
  LAYER M3 ;
        RECT 29.216 12.164 29.248 12.196 ;
  LAYER M1 ;
        RECT 29.152 9.708 29.184 12.216 ;
  LAYER M3 ;
        RECT 29.152 9.728 29.184 9.76 ;
  LAYER M1 ;
        RECT 29.088 9.708 29.12 12.216 ;
  LAYER M3 ;
        RECT 29.088 12.164 29.12 12.196 ;
  LAYER M1 ;
        RECT 29.024 9.708 29.056 12.216 ;
  LAYER M3 ;
        RECT 29.024 9.728 29.056 9.76 ;
  LAYER M1 ;
        RECT 28.96 9.708 28.992 12.216 ;
  LAYER M3 ;
        RECT 28.96 12.164 28.992 12.196 ;
  LAYER M1 ;
        RECT 28.896 9.708 28.928 12.216 ;
  LAYER M3 ;
        RECT 28.896 9.728 28.928 9.76 ;
  LAYER M1 ;
        RECT 28.832 9.708 28.864 12.216 ;
  LAYER M3 ;
        RECT 28.832 12.164 28.864 12.196 ;
  LAYER M1 ;
        RECT 28.768 9.708 28.8 12.216 ;
  LAYER M3 ;
        RECT 28.768 9.728 28.8 9.76 ;
  LAYER M1 ;
        RECT 28.704 9.708 28.736 12.216 ;
  LAYER M3 ;
        RECT 28.704 12.164 28.736 12.196 ;
  LAYER M1 ;
        RECT 28.64 9.708 28.672 12.216 ;
  LAYER M3 ;
        RECT 28.64 9.728 28.672 9.76 ;
  LAYER M1 ;
        RECT 28.576 9.708 28.608 12.216 ;
  LAYER M3 ;
        RECT 28.576 12.164 28.608 12.196 ;
  LAYER M1 ;
        RECT 28.512 9.708 28.544 12.216 ;
  LAYER M3 ;
        RECT 30.88 9.792 30.912 9.824 ;
  LAYER M2 ;
        RECT 28.512 9.856 28.544 9.888 ;
  LAYER M2 ;
        RECT 30.88 9.92 30.912 9.952 ;
  LAYER M2 ;
        RECT 28.512 9.984 28.544 10.016 ;
  LAYER M2 ;
        RECT 30.88 10.048 30.912 10.08 ;
  LAYER M2 ;
        RECT 28.512 10.112 28.544 10.144 ;
  LAYER M2 ;
        RECT 30.88 10.176 30.912 10.208 ;
  LAYER M2 ;
        RECT 28.512 10.24 28.544 10.272 ;
  LAYER M2 ;
        RECT 30.88 10.304 30.912 10.336 ;
  LAYER M2 ;
        RECT 28.512 10.368 28.544 10.4 ;
  LAYER M2 ;
        RECT 30.88 10.432 30.912 10.464 ;
  LAYER M2 ;
        RECT 28.512 10.496 28.544 10.528 ;
  LAYER M2 ;
        RECT 30.88 10.56 30.912 10.592 ;
  LAYER M2 ;
        RECT 28.512 10.624 28.544 10.656 ;
  LAYER M2 ;
        RECT 30.88 10.688 30.912 10.72 ;
  LAYER M2 ;
        RECT 28.512 10.752 28.544 10.784 ;
  LAYER M2 ;
        RECT 30.88 10.816 30.912 10.848 ;
  LAYER M2 ;
        RECT 28.512 10.88 28.544 10.912 ;
  LAYER M2 ;
        RECT 30.88 10.944 30.912 10.976 ;
  LAYER M2 ;
        RECT 28.512 11.008 28.544 11.04 ;
  LAYER M2 ;
        RECT 30.88 11.072 30.912 11.104 ;
  LAYER M2 ;
        RECT 28.512 11.136 28.544 11.168 ;
  LAYER M2 ;
        RECT 30.88 11.2 30.912 11.232 ;
  LAYER M2 ;
        RECT 28.512 11.264 28.544 11.296 ;
  LAYER M2 ;
        RECT 30.88 11.328 30.912 11.36 ;
  LAYER M2 ;
        RECT 28.512 11.392 28.544 11.424 ;
  LAYER M2 ;
        RECT 30.88 11.456 30.912 11.488 ;
  LAYER M2 ;
        RECT 28.512 11.52 28.544 11.552 ;
  LAYER M2 ;
        RECT 30.88 11.584 30.912 11.616 ;
  LAYER M2 ;
        RECT 28.512 11.648 28.544 11.68 ;
  LAYER M2 ;
        RECT 30.88 11.712 30.912 11.744 ;
  LAYER M2 ;
        RECT 28.512 11.776 28.544 11.808 ;
  LAYER M2 ;
        RECT 30.88 11.84 30.912 11.872 ;
  LAYER M2 ;
        RECT 28.512 11.904 28.544 11.936 ;
  LAYER M2 ;
        RECT 30.88 11.968 30.912 12 ;
  LAYER M2 ;
        RECT 28.512 12.032 28.544 12.064 ;
  LAYER M2 ;
        RECT 28.464 9.66 30.96 12.264 ;
  LAYER M1 ;
        RECT 30.88 12.816 30.912 15.324 ;
  LAYER M3 ;
        RECT 30.88 15.272 30.912 15.304 ;
  LAYER M1 ;
        RECT 30.816 12.816 30.848 15.324 ;
  LAYER M3 ;
        RECT 30.816 12.836 30.848 12.868 ;
  LAYER M1 ;
        RECT 30.752 12.816 30.784 15.324 ;
  LAYER M3 ;
        RECT 30.752 15.272 30.784 15.304 ;
  LAYER M1 ;
        RECT 30.688 12.816 30.72 15.324 ;
  LAYER M3 ;
        RECT 30.688 12.836 30.72 12.868 ;
  LAYER M1 ;
        RECT 30.624 12.816 30.656 15.324 ;
  LAYER M3 ;
        RECT 30.624 15.272 30.656 15.304 ;
  LAYER M1 ;
        RECT 30.56 12.816 30.592 15.324 ;
  LAYER M3 ;
        RECT 30.56 12.836 30.592 12.868 ;
  LAYER M1 ;
        RECT 30.496 12.816 30.528 15.324 ;
  LAYER M3 ;
        RECT 30.496 15.272 30.528 15.304 ;
  LAYER M1 ;
        RECT 30.432 12.816 30.464 15.324 ;
  LAYER M3 ;
        RECT 30.432 12.836 30.464 12.868 ;
  LAYER M1 ;
        RECT 30.368 12.816 30.4 15.324 ;
  LAYER M3 ;
        RECT 30.368 15.272 30.4 15.304 ;
  LAYER M1 ;
        RECT 30.304 12.816 30.336 15.324 ;
  LAYER M3 ;
        RECT 30.304 12.836 30.336 12.868 ;
  LAYER M1 ;
        RECT 30.24 12.816 30.272 15.324 ;
  LAYER M3 ;
        RECT 30.24 15.272 30.272 15.304 ;
  LAYER M1 ;
        RECT 30.176 12.816 30.208 15.324 ;
  LAYER M3 ;
        RECT 30.176 12.836 30.208 12.868 ;
  LAYER M1 ;
        RECT 30.112 12.816 30.144 15.324 ;
  LAYER M3 ;
        RECT 30.112 15.272 30.144 15.304 ;
  LAYER M1 ;
        RECT 30.048 12.816 30.08 15.324 ;
  LAYER M3 ;
        RECT 30.048 12.836 30.08 12.868 ;
  LAYER M1 ;
        RECT 29.984 12.816 30.016 15.324 ;
  LAYER M3 ;
        RECT 29.984 15.272 30.016 15.304 ;
  LAYER M1 ;
        RECT 29.92 12.816 29.952 15.324 ;
  LAYER M3 ;
        RECT 29.92 12.836 29.952 12.868 ;
  LAYER M1 ;
        RECT 29.856 12.816 29.888 15.324 ;
  LAYER M3 ;
        RECT 29.856 15.272 29.888 15.304 ;
  LAYER M1 ;
        RECT 29.792 12.816 29.824 15.324 ;
  LAYER M3 ;
        RECT 29.792 12.836 29.824 12.868 ;
  LAYER M1 ;
        RECT 29.728 12.816 29.76 15.324 ;
  LAYER M3 ;
        RECT 29.728 15.272 29.76 15.304 ;
  LAYER M1 ;
        RECT 29.664 12.816 29.696 15.324 ;
  LAYER M3 ;
        RECT 29.664 12.836 29.696 12.868 ;
  LAYER M1 ;
        RECT 29.6 12.816 29.632 15.324 ;
  LAYER M3 ;
        RECT 29.6 15.272 29.632 15.304 ;
  LAYER M1 ;
        RECT 29.536 12.816 29.568 15.324 ;
  LAYER M3 ;
        RECT 29.536 12.836 29.568 12.868 ;
  LAYER M1 ;
        RECT 29.472 12.816 29.504 15.324 ;
  LAYER M3 ;
        RECT 29.472 15.272 29.504 15.304 ;
  LAYER M1 ;
        RECT 29.408 12.816 29.44 15.324 ;
  LAYER M3 ;
        RECT 29.408 12.836 29.44 12.868 ;
  LAYER M1 ;
        RECT 29.344 12.816 29.376 15.324 ;
  LAYER M3 ;
        RECT 29.344 15.272 29.376 15.304 ;
  LAYER M1 ;
        RECT 29.28 12.816 29.312 15.324 ;
  LAYER M3 ;
        RECT 29.28 12.836 29.312 12.868 ;
  LAYER M1 ;
        RECT 29.216 12.816 29.248 15.324 ;
  LAYER M3 ;
        RECT 29.216 15.272 29.248 15.304 ;
  LAYER M1 ;
        RECT 29.152 12.816 29.184 15.324 ;
  LAYER M3 ;
        RECT 29.152 12.836 29.184 12.868 ;
  LAYER M1 ;
        RECT 29.088 12.816 29.12 15.324 ;
  LAYER M3 ;
        RECT 29.088 15.272 29.12 15.304 ;
  LAYER M1 ;
        RECT 29.024 12.816 29.056 15.324 ;
  LAYER M3 ;
        RECT 29.024 12.836 29.056 12.868 ;
  LAYER M1 ;
        RECT 28.96 12.816 28.992 15.324 ;
  LAYER M3 ;
        RECT 28.96 15.272 28.992 15.304 ;
  LAYER M1 ;
        RECT 28.896 12.816 28.928 15.324 ;
  LAYER M3 ;
        RECT 28.896 12.836 28.928 12.868 ;
  LAYER M1 ;
        RECT 28.832 12.816 28.864 15.324 ;
  LAYER M3 ;
        RECT 28.832 15.272 28.864 15.304 ;
  LAYER M1 ;
        RECT 28.768 12.816 28.8 15.324 ;
  LAYER M3 ;
        RECT 28.768 12.836 28.8 12.868 ;
  LAYER M1 ;
        RECT 28.704 12.816 28.736 15.324 ;
  LAYER M3 ;
        RECT 28.704 15.272 28.736 15.304 ;
  LAYER M1 ;
        RECT 28.64 12.816 28.672 15.324 ;
  LAYER M3 ;
        RECT 28.64 12.836 28.672 12.868 ;
  LAYER M1 ;
        RECT 28.576 12.816 28.608 15.324 ;
  LAYER M3 ;
        RECT 28.576 15.272 28.608 15.304 ;
  LAYER M1 ;
        RECT 28.512 12.816 28.544 15.324 ;
  LAYER M3 ;
        RECT 30.88 12.9 30.912 12.932 ;
  LAYER M2 ;
        RECT 28.512 12.964 28.544 12.996 ;
  LAYER M2 ;
        RECT 30.88 13.028 30.912 13.06 ;
  LAYER M2 ;
        RECT 28.512 13.092 28.544 13.124 ;
  LAYER M2 ;
        RECT 30.88 13.156 30.912 13.188 ;
  LAYER M2 ;
        RECT 28.512 13.22 28.544 13.252 ;
  LAYER M2 ;
        RECT 30.88 13.284 30.912 13.316 ;
  LAYER M2 ;
        RECT 28.512 13.348 28.544 13.38 ;
  LAYER M2 ;
        RECT 30.88 13.412 30.912 13.444 ;
  LAYER M2 ;
        RECT 28.512 13.476 28.544 13.508 ;
  LAYER M2 ;
        RECT 30.88 13.54 30.912 13.572 ;
  LAYER M2 ;
        RECT 28.512 13.604 28.544 13.636 ;
  LAYER M2 ;
        RECT 30.88 13.668 30.912 13.7 ;
  LAYER M2 ;
        RECT 28.512 13.732 28.544 13.764 ;
  LAYER M2 ;
        RECT 30.88 13.796 30.912 13.828 ;
  LAYER M2 ;
        RECT 28.512 13.86 28.544 13.892 ;
  LAYER M2 ;
        RECT 30.88 13.924 30.912 13.956 ;
  LAYER M2 ;
        RECT 28.512 13.988 28.544 14.02 ;
  LAYER M2 ;
        RECT 30.88 14.052 30.912 14.084 ;
  LAYER M2 ;
        RECT 28.512 14.116 28.544 14.148 ;
  LAYER M2 ;
        RECT 30.88 14.18 30.912 14.212 ;
  LAYER M2 ;
        RECT 28.512 14.244 28.544 14.276 ;
  LAYER M2 ;
        RECT 30.88 14.308 30.912 14.34 ;
  LAYER M2 ;
        RECT 28.512 14.372 28.544 14.404 ;
  LAYER M2 ;
        RECT 30.88 14.436 30.912 14.468 ;
  LAYER M2 ;
        RECT 28.512 14.5 28.544 14.532 ;
  LAYER M2 ;
        RECT 30.88 14.564 30.912 14.596 ;
  LAYER M2 ;
        RECT 28.512 14.628 28.544 14.66 ;
  LAYER M2 ;
        RECT 30.88 14.692 30.912 14.724 ;
  LAYER M2 ;
        RECT 28.512 14.756 28.544 14.788 ;
  LAYER M2 ;
        RECT 30.88 14.82 30.912 14.852 ;
  LAYER M2 ;
        RECT 28.512 14.884 28.544 14.916 ;
  LAYER M2 ;
        RECT 30.88 14.948 30.912 14.98 ;
  LAYER M2 ;
        RECT 28.512 15.012 28.544 15.044 ;
  LAYER M2 ;
        RECT 30.88 15.076 30.912 15.108 ;
  LAYER M2 ;
        RECT 28.512 15.14 28.544 15.172 ;
  LAYER M2 ;
        RECT 28.464 12.768 30.96 15.372 ;
  LAYER M1 ;
        RECT 30.88 15.924 30.912 18.432 ;
  LAYER M3 ;
        RECT 30.88 18.38 30.912 18.412 ;
  LAYER M1 ;
        RECT 30.816 15.924 30.848 18.432 ;
  LAYER M3 ;
        RECT 30.816 15.944 30.848 15.976 ;
  LAYER M1 ;
        RECT 30.752 15.924 30.784 18.432 ;
  LAYER M3 ;
        RECT 30.752 18.38 30.784 18.412 ;
  LAYER M1 ;
        RECT 30.688 15.924 30.72 18.432 ;
  LAYER M3 ;
        RECT 30.688 15.944 30.72 15.976 ;
  LAYER M1 ;
        RECT 30.624 15.924 30.656 18.432 ;
  LAYER M3 ;
        RECT 30.624 18.38 30.656 18.412 ;
  LAYER M1 ;
        RECT 30.56 15.924 30.592 18.432 ;
  LAYER M3 ;
        RECT 30.56 15.944 30.592 15.976 ;
  LAYER M1 ;
        RECT 30.496 15.924 30.528 18.432 ;
  LAYER M3 ;
        RECT 30.496 18.38 30.528 18.412 ;
  LAYER M1 ;
        RECT 30.432 15.924 30.464 18.432 ;
  LAYER M3 ;
        RECT 30.432 15.944 30.464 15.976 ;
  LAYER M1 ;
        RECT 30.368 15.924 30.4 18.432 ;
  LAYER M3 ;
        RECT 30.368 18.38 30.4 18.412 ;
  LAYER M1 ;
        RECT 30.304 15.924 30.336 18.432 ;
  LAYER M3 ;
        RECT 30.304 15.944 30.336 15.976 ;
  LAYER M1 ;
        RECT 30.24 15.924 30.272 18.432 ;
  LAYER M3 ;
        RECT 30.24 18.38 30.272 18.412 ;
  LAYER M1 ;
        RECT 30.176 15.924 30.208 18.432 ;
  LAYER M3 ;
        RECT 30.176 15.944 30.208 15.976 ;
  LAYER M1 ;
        RECT 30.112 15.924 30.144 18.432 ;
  LAYER M3 ;
        RECT 30.112 18.38 30.144 18.412 ;
  LAYER M1 ;
        RECT 30.048 15.924 30.08 18.432 ;
  LAYER M3 ;
        RECT 30.048 15.944 30.08 15.976 ;
  LAYER M1 ;
        RECT 29.984 15.924 30.016 18.432 ;
  LAYER M3 ;
        RECT 29.984 18.38 30.016 18.412 ;
  LAYER M1 ;
        RECT 29.92 15.924 29.952 18.432 ;
  LAYER M3 ;
        RECT 29.92 15.944 29.952 15.976 ;
  LAYER M1 ;
        RECT 29.856 15.924 29.888 18.432 ;
  LAYER M3 ;
        RECT 29.856 18.38 29.888 18.412 ;
  LAYER M1 ;
        RECT 29.792 15.924 29.824 18.432 ;
  LAYER M3 ;
        RECT 29.792 15.944 29.824 15.976 ;
  LAYER M1 ;
        RECT 29.728 15.924 29.76 18.432 ;
  LAYER M3 ;
        RECT 29.728 18.38 29.76 18.412 ;
  LAYER M1 ;
        RECT 29.664 15.924 29.696 18.432 ;
  LAYER M3 ;
        RECT 29.664 15.944 29.696 15.976 ;
  LAYER M1 ;
        RECT 29.6 15.924 29.632 18.432 ;
  LAYER M3 ;
        RECT 29.6 18.38 29.632 18.412 ;
  LAYER M1 ;
        RECT 29.536 15.924 29.568 18.432 ;
  LAYER M3 ;
        RECT 29.536 15.944 29.568 15.976 ;
  LAYER M1 ;
        RECT 29.472 15.924 29.504 18.432 ;
  LAYER M3 ;
        RECT 29.472 18.38 29.504 18.412 ;
  LAYER M1 ;
        RECT 29.408 15.924 29.44 18.432 ;
  LAYER M3 ;
        RECT 29.408 15.944 29.44 15.976 ;
  LAYER M1 ;
        RECT 29.344 15.924 29.376 18.432 ;
  LAYER M3 ;
        RECT 29.344 18.38 29.376 18.412 ;
  LAYER M1 ;
        RECT 29.28 15.924 29.312 18.432 ;
  LAYER M3 ;
        RECT 29.28 15.944 29.312 15.976 ;
  LAYER M1 ;
        RECT 29.216 15.924 29.248 18.432 ;
  LAYER M3 ;
        RECT 29.216 18.38 29.248 18.412 ;
  LAYER M1 ;
        RECT 29.152 15.924 29.184 18.432 ;
  LAYER M3 ;
        RECT 29.152 15.944 29.184 15.976 ;
  LAYER M1 ;
        RECT 29.088 15.924 29.12 18.432 ;
  LAYER M3 ;
        RECT 29.088 18.38 29.12 18.412 ;
  LAYER M1 ;
        RECT 29.024 15.924 29.056 18.432 ;
  LAYER M3 ;
        RECT 29.024 15.944 29.056 15.976 ;
  LAYER M1 ;
        RECT 28.96 15.924 28.992 18.432 ;
  LAYER M3 ;
        RECT 28.96 18.38 28.992 18.412 ;
  LAYER M1 ;
        RECT 28.896 15.924 28.928 18.432 ;
  LAYER M3 ;
        RECT 28.896 15.944 28.928 15.976 ;
  LAYER M1 ;
        RECT 28.832 15.924 28.864 18.432 ;
  LAYER M3 ;
        RECT 28.832 18.38 28.864 18.412 ;
  LAYER M1 ;
        RECT 28.768 15.924 28.8 18.432 ;
  LAYER M3 ;
        RECT 28.768 15.944 28.8 15.976 ;
  LAYER M1 ;
        RECT 28.704 15.924 28.736 18.432 ;
  LAYER M3 ;
        RECT 28.704 18.38 28.736 18.412 ;
  LAYER M1 ;
        RECT 28.64 15.924 28.672 18.432 ;
  LAYER M3 ;
        RECT 28.64 15.944 28.672 15.976 ;
  LAYER M1 ;
        RECT 28.576 15.924 28.608 18.432 ;
  LAYER M3 ;
        RECT 28.576 18.38 28.608 18.412 ;
  LAYER M1 ;
        RECT 28.512 15.924 28.544 18.432 ;
  LAYER M3 ;
        RECT 30.88 16.008 30.912 16.04 ;
  LAYER M2 ;
        RECT 28.512 16.072 28.544 16.104 ;
  LAYER M2 ;
        RECT 30.88 16.136 30.912 16.168 ;
  LAYER M2 ;
        RECT 28.512 16.2 28.544 16.232 ;
  LAYER M2 ;
        RECT 30.88 16.264 30.912 16.296 ;
  LAYER M2 ;
        RECT 28.512 16.328 28.544 16.36 ;
  LAYER M2 ;
        RECT 30.88 16.392 30.912 16.424 ;
  LAYER M2 ;
        RECT 28.512 16.456 28.544 16.488 ;
  LAYER M2 ;
        RECT 30.88 16.52 30.912 16.552 ;
  LAYER M2 ;
        RECT 28.512 16.584 28.544 16.616 ;
  LAYER M2 ;
        RECT 30.88 16.648 30.912 16.68 ;
  LAYER M2 ;
        RECT 28.512 16.712 28.544 16.744 ;
  LAYER M2 ;
        RECT 30.88 16.776 30.912 16.808 ;
  LAYER M2 ;
        RECT 28.512 16.84 28.544 16.872 ;
  LAYER M2 ;
        RECT 30.88 16.904 30.912 16.936 ;
  LAYER M2 ;
        RECT 28.512 16.968 28.544 17 ;
  LAYER M2 ;
        RECT 30.88 17.032 30.912 17.064 ;
  LAYER M2 ;
        RECT 28.512 17.096 28.544 17.128 ;
  LAYER M2 ;
        RECT 30.88 17.16 30.912 17.192 ;
  LAYER M2 ;
        RECT 28.512 17.224 28.544 17.256 ;
  LAYER M2 ;
        RECT 30.88 17.288 30.912 17.32 ;
  LAYER M2 ;
        RECT 28.512 17.352 28.544 17.384 ;
  LAYER M2 ;
        RECT 30.88 17.416 30.912 17.448 ;
  LAYER M2 ;
        RECT 28.512 17.48 28.544 17.512 ;
  LAYER M2 ;
        RECT 30.88 17.544 30.912 17.576 ;
  LAYER M2 ;
        RECT 28.512 17.608 28.544 17.64 ;
  LAYER M2 ;
        RECT 30.88 17.672 30.912 17.704 ;
  LAYER M2 ;
        RECT 28.512 17.736 28.544 17.768 ;
  LAYER M2 ;
        RECT 30.88 17.8 30.912 17.832 ;
  LAYER M2 ;
        RECT 28.512 17.864 28.544 17.896 ;
  LAYER M2 ;
        RECT 30.88 17.928 30.912 17.96 ;
  LAYER M2 ;
        RECT 28.512 17.992 28.544 18.024 ;
  LAYER M2 ;
        RECT 30.88 18.056 30.912 18.088 ;
  LAYER M2 ;
        RECT 28.512 18.12 28.544 18.152 ;
  LAYER M2 ;
        RECT 30.88 18.184 30.912 18.216 ;
  LAYER M2 ;
        RECT 28.512 18.248 28.544 18.28 ;
  LAYER M2 ;
        RECT 28.464 15.876 30.96 18.48 ;
  LAYER M1 ;
        RECT 27.904 6.6 27.936 9.108 ;
  LAYER M3 ;
        RECT 27.904 9.056 27.936 9.088 ;
  LAYER M1 ;
        RECT 27.84 6.6 27.872 9.108 ;
  LAYER M3 ;
        RECT 27.84 6.62 27.872 6.652 ;
  LAYER M1 ;
        RECT 27.776 6.6 27.808 9.108 ;
  LAYER M3 ;
        RECT 27.776 9.056 27.808 9.088 ;
  LAYER M1 ;
        RECT 27.712 6.6 27.744 9.108 ;
  LAYER M3 ;
        RECT 27.712 6.62 27.744 6.652 ;
  LAYER M1 ;
        RECT 27.648 6.6 27.68 9.108 ;
  LAYER M3 ;
        RECT 27.648 9.056 27.68 9.088 ;
  LAYER M1 ;
        RECT 27.584 6.6 27.616 9.108 ;
  LAYER M3 ;
        RECT 27.584 6.62 27.616 6.652 ;
  LAYER M1 ;
        RECT 27.52 6.6 27.552 9.108 ;
  LAYER M3 ;
        RECT 27.52 9.056 27.552 9.088 ;
  LAYER M1 ;
        RECT 27.456 6.6 27.488 9.108 ;
  LAYER M3 ;
        RECT 27.456 6.62 27.488 6.652 ;
  LAYER M1 ;
        RECT 27.392 6.6 27.424 9.108 ;
  LAYER M3 ;
        RECT 27.392 9.056 27.424 9.088 ;
  LAYER M1 ;
        RECT 27.328 6.6 27.36 9.108 ;
  LAYER M3 ;
        RECT 27.328 6.62 27.36 6.652 ;
  LAYER M1 ;
        RECT 27.264 6.6 27.296 9.108 ;
  LAYER M3 ;
        RECT 27.264 9.056 27.296 9.088 ;
  LAYER M1 ;
        RECT 27.2 6.6 27.232 9.108 ;
  LAYER M3 ;
        RECT 27.2 6.62 27.232 6.652 ;
  LAYER M1 ;
        RECT 27.136 6.6 27.168 9.108 ;
  LAYER M3 ;
        RECT 27.136 9.056 27.168 9.088 ;
  LAYER M1 ;
        RECT 27.072 6.6 27.104 9.108 ;
  LAYER M3 ;
        RECT 27.072 6.62 27.104 6.652 ;
  LAYER M1 ;
        RECT 27.008 6.6 27.04 9.108 ;
  LAYER M3 ;
        RECT 27.008 9.056 27.04 9.088 ;
  LAYER M1 ;
        RECT 26.944 6.6 26.976 9.108 ;
  LAYER M3 ;
        RECT 26.944 6.62 26.976 6.652 ;
  LAYER M1 ;
        RECT 26.88 6.6 26.912 9.108 ;
  LAYER M3 ;
        RECT 26.88 9.056 26.912 9.088 ;
  LAYER M1 ;
        RECT 26.816 6.6 26.848 9.108 ;
  LAYER M3 ;
        RECT 26.816 6.62 26.848 6.652 ;
  LAYER M1 ;
        RECT 26.752 6.6 26.784 9.108 ;
  LAYER M3 ;
        RECT 26.752 9.056 26.784 9.088 ;
  LAYER M1 ;
        RECT 26.688 6.6 26.72 9.108 ;
  LAYER M3 ;
        RECT 26.688 6.62 26.72 6.652 ;
  LAYER M1 ;
        RECT 26.624 6.6 26.656 9.108 ;
  LAYER M3 ;
        RECT 26.624 9.056 26.656 9.088 ;
  LAYER M1 ;
        RECT 26.56 6.6 26.592 9.108 ;
  LAYER M3 ;
        RECT 26.56 6.62 26.592 6.652 ;
  LAYER M1 ;
        RECT 26.496 6.6 26.528 9.108 ;
  LAYER M3 ;
        RECT 26.496 9.056 26.528 9.088 ;
  LAYER M1 ;
        RECT 26.432 6.6 26.464 9.108 ;
  LAYER M3 ;
        RECT 26.432 6.62 26.464 6.652 ;
  LAYER M1 ;
        RECT 26.368 6.6 26.4 9.108 ;
  LAYER M3 ;
        RECT 26.368 9.056 26.4 9.088 ;
  LAYER M1 ;
        RECT 26.304 6.6 26.336 9.108 ;
  LAYER M3 ;
        RECT 26.304 6.62 26.336 6.652 ;
  LAYER M1 ;
        RECT 26.24 6.6 26.272 9.108 ;
  LAYER M3 ;
        RECT 26.24 9.056 26.272 9.088 ;
  LAYER M1 ;
        RECT 26.176 6.6 26.208 9.108 ;
  LAYER M3 ;
        RECT 26.176 6.62 26.208 6.652 ;
  LAYER M1 ;
        RECT 26.112 6.6 26.144 9.108 ;
  LAYER M3 ;
        RECT 26.112 9.056 26.144 9.088 ;
  LAYER M1 ;
        RECT 26.048 6.6 26.08 9.108 ;
  LAYER M3 ;
        RECT 26.048 6.62 26.08 6.652 ;
  LAYER M1 ;
        RECT 25.984 6.6 26.016 9.108 ;
  LAYER M3 ;
        RECT 25.984 9.056 26.016 9.088 ;
  LAYER M1 ;
        RECT 25.92 6.6 25.952 9.108 ;
  LAYER M3 ;
        RECT 25.92 6.62 25.952 6.652 ;
  LAYER M1 ;
        RECT 25.856 6.6 25.888 9.108 ;
  LAYER M3 ;
        RECT 25.856 9.056 25.888 9.088 ;
  LAYER M1 ;
        RECT 25.792 6.6 25.824 9.108 ;
  LAYER M3 ;
        RECT 25.792 6.62 25.824 6.652 ;
  LAYER M1 ;
        RECT 25.728 6.6 25.76 9.108 ;
  LAYER M3 ;
        RECT 25.728 9.056 25.76 9.088 ;
  LAYER M1 ;
        RECT 25.664 6.6 25.696 9.108 ;
  LAYER M3 ;
        RECT 25.664 6.62 25.696 6.652 ;
  LAYER M1 ;
        RECT 25.6 6.6 25.632 9.108 ;
  LAYER M3 ;
        RECT 25.6 9.056 25.632 9.088 ;
  LAYER M1 ;
        RECT 25.536 6.6 25.568 9.108 ;
  LAYER M3 ;
        RECT 27.904 6.684 27.936 6.716 ;
  LAYER M2 ;
        RECT 25.536 6.748 25.568 6.78 ;
  LAYER M2 ;
        RECT 27.904 6.812 27.936 6.844 ;
  LAYER M2 ;
        RECT 25.536 6.876 25.568 6.908 ;
  LAYER M2 ;
        RECT 27.904 6.94 27.936 6.972 ;
  LAYER M2 ;
        RECT 25.536 7.004 25.568 7.036 ;
  LAYER M2 ;
        RECT 27.904 7.068 27.936 7.1 ;
  LAYER M2 ;
        RECT 25.536 7.132 25.568 7.164 ;
  LAYER M2 ;
        RECT 27.904 7.196 27.936 7.228 ;
  LAYER M2 ;
        RECT 25.536 7.26 25.568 7.292 ;
  LAYER M2 ;
        RECT 27.904 7.324 27.936 7.356 ;
  LAYER M2 ;
        RECT 25.536 7.388 25.568 7.42 ;
  LAYER M2 ;
        RECT 27.904 7.452 27.936 7.484 ;
  LAYER M2 ;
        RECT 25.536 7.516 25.568 7.548 ;
  LAYER M2 ;
        RECT 27.904 7.58 27.936 7.612 ;
  LAYER M2 ;
        RECT 25.536 7.644 25.568 7.676 ;
  LAYER M2 ;
        RECT 27.904 7.708 27.936 7.74 ;
  LAYER M2 ;
        RECT 25.536 7.772 25.568 7.804 ;
  LAYER M2 ;
        RECT 27.904 7.836 27.936 7.868 ;
  LAYER M2 ;
        RECT 25.536 7.9 25.568 7.932 ;
  LAYER M2 ;
        RECT 27.904 7.964 27.936 7.996 ;
  LAYER M2 ;
        RECT 25.536 8.028 25.568 8.06 ;
  LAYER M2 ;
        RECT 27.904 8.092 27.936 8.124 ;
  LAYER M2 ;
        RECT 25.536 8.156 25.568 8.188 ;
  LAYER M2 ;
        RECT 27.904 8.22 27.936 8.252 ;
  LAYER M2 ;
        RECT 25.536 8.284 25.568 8.316 ;
  LAYER M2 ;
        RECT 27.904 8.348 27.936 8.38 ;
  LAYER M2 ;
        RECT 25.536 8.412 25.568 8.444 ;
  LAYER M2 ;
        RECT 27.904 8.476 27.936 8.508 ;
  LAYER M2 ;
        RECT 25.536 8.54 25.568 8.572 ;
  LAYER M2 ;
        RECT 27.904 8.604 27.936 8.636 ;
  LAYER M2 ;
        RECT 25.536 8.668 25.568 8.7 ;
  LAYER M2 ;
        RECT 27.904 8.732 27.936 8.764 ;
  LAYER M2 ;
        RECT 25.536 8.796 25.568 8.828 ;
  LAYER M2 ;
        RECT 27.904 8.86 27.936 8.892 ;
  LAYER M2 ;
        RECT 25.536 8.924 25.568 8.956 ;
  LAYER M2 ;
        RECT 25.488 6.552 27.984 9.156 ;
  LAYER M1 ;
        RECT 27.904 9.708 27.936 12.216 ;
  LAYER M3 ;
        RECT 27.904 12.164 27.936 12.196 ;
  LAYER M1 ;
        RECT 27.84 9.708 27.872 12.216 ;
  LAYER M3 ;
        RECT 27.84 9.728 27.872 9.76 ;
  LAYER M1 ;
        RECT 27.776 9.708 27.808 12.216 ;
  LAYER M3 ;
        RECT 27.776 12.164 27.808 12.196 ;
  LAYER M1 ;
        RECT 27.712 9.708 27.744 12.216 ;
  LAYER M3 ;
        RECT 27.712 9.728 27.744 9.76 ;
  LAYER M1 ;
        RECT 27.648 9.708 27.68 12.216 ;
  LAYER M3 ;
        RECT 27.648 12.164 27.68 12.196 ;
  LAYER M1 ;
        RECT 27.584 9.708 27.616 12.216 ;
  LAYER M3 ;
        RECT 27.584 9.728 27.616 9.76 ;
  LAYER M1 ;
        RECT 27.52 9.708 27.552 12.216 ;
  LAYER M3 ;
        RECT 27.52 12.164 27.552 12.196 ;
  LAYER M1 ;
        RECT 27.456 9.708 27.488 12.216 ;
  LAYER M3 ;
        RECT 27.456 9.728 27.488 9.76 ;
  LAYER M1 ;
        RECT 27.392 9.708 27.424 12.216 ;
  LAYER M3 ;
        RECT 27.392 12.164 27.424 12.196 ;
  LAYER M1 ;
        RECT 27.328 9.708 27.36 12.216 ;
  LAYER M3 ;
        RECT 27.328 9.728 27.36 9.76 ;
  LAYER M1 ;
        RECT 27.264 9.708 27.296 12.216 ;
  LAYER M3 ;
        RECT 27.264 12.164 27.296 12.196 ;
  LAYER M1 ;
        RECT 27.2 9.708 27.232 12.216 ;
  LAYER M3 ;
        RECT 27.2 9.728 27.232 9.76 ;
  LAYER M1 ;
        RECT 27.136 9.708 27.168 12.216 ;
  LAYER M3 ;
        RECT 27.136 12.164 27.168 12.196 ;
  LAYER M1 ;
        RECT 27.072 9.708 27.104 12.216 ;
  LAYER M3 ;
        RECT 27.072 9.728 27.104 9.76 ;
  LAYER M1 ;
        RECT 27.008 9.708 27.04 12.216 ;
  LAYER M3 ;
        RECT 27.008 12.164 27.04 12.196 ;
  LAYER M1 ;
        RECT 26.944 9.708 26.976 12.216 ;
  LAYER M3 ;
        RECT 26.944 9.728 26.976 9.76 ;
  LAYER M1 ;
        RECT 26.88 9.708 26.912 12.216 ;
  LAYER M3 ;
        RECT 26.88 12.164 26.912 12.196 ;
  LAYER M1 ;
        RECT 26.816 9.708 26.848 12.216 ;
  LAYER M3 ;
        RECT 26.816 9.728 26.848 9.76 ;
  LAYER M1 ;
        RECT 26.752 9.708 26.784 12.216 ;
  LAYER M3 ;
        RECT 26.752 12.164 26.784 12.196 ;
  LAYER M1 ;
        RECT 26.688 9.708 26.72 12.216 ;
  LAYER M3 ;
        RECT 26.688 9.728 26.72 9.76 ;
  LAYER M1 ;
        RECT 26.624 9.708 26.656 12.216 ;
  LAYER M3 ;
        RECT 26.624 12.164 26.656 12.196 ;
  LAYER M1 ;
        RECT 26.56 9.708 26.592 12.216 ;
  LAYER M3 ;
        RECT 26.56 9.728 26.592 9.76 ;
  LAYER M1 ;
        RECT 26.496 9.708 26.528 12.216 ;
  LAYER M3 ;
        RECT 26.496 12.164 26.528 12.196 ;
  LAYER M1 ;
        RECT 26.432 9.708 26.464 12.216 ;
  LAYER M3 ;
        RECT 26.432 9.728 26.464 9.76 ;
  LAYER M1 ;
        RECT 26.368 9.708 26.4 12.216 ;
  LAYER M3 ;
        RECT 26.368 12.164 26.4 12.196 ;
  LAYER M1 ;
        RECT 26.304 9.708 26.336 12.216 ;
  LAYER M3 ;
        RECT 26.304 9.728 26.336 9.76 ;
  LAYER M1 ;
        RECT 26.24 9.708 26.272 12.216 ;
  LAYER M3 ;
        RECT 26.24 12.164 26.272 12.196 ;
  LAYER M1 ;
        RECT 26.176 9.708 26.208 12.216 ;
  LAYER M3 ;
        RECT 26.176 9.728 26.208 9.76 ;
  LAYER M1 ;
        RECT 26.112 9.708 26.144 12.216 ;
  LAYER M3 ;
        RECT 26.112 12.164 26.144 12.196 ;
  LAYER M1 ;
        RECT 26.048 9.708 26.08 12.216 ;
  LAYER M3 ;
        RECT 26.048 9.728 26.08 9.76 ;
  LAYER M1 ;
        RECT 25.984 9.708 26.016 12.216 ;
  LAYER M3 ;
        RECT 25.984 12.164 26.016 12.196 ;
  LAYER M1 ;
        RECT 25.92 9.708 25.952 12.216 ;
  LAYER M3 ;
        RECT 25.92 9.728 25.952 9.76 ;
  LAYER M1 ;
        RECT 25.856 9.708 25.888 12.216 ;
  LAYER M3 ;
        RECT 25.856 12.164 25.888 12.196 ;
  LAYER M1 ;
        RECT 25.792 9.708 25.824 12.216 ;
  LAYER M3 ;
        RECT 25.792 9.728 25.824 9.76 ;
  LAYER M1 ;
        RECT 25.728 9.708 25.76 12.216 ;
  LAYER M3 ;
        RECT 25.728 12.164 25.76 12.196 ;
  LAYER M1 ;
        RECT 25.664 9.708 25.696 12.216 ;
  LAYER M3 ;
        RECT 25.664 9.728 25.696 9.76 ;
  LAYER M1 ;
        RECT 25.6 9.708 25.632 12.216 ;
  LAYER M3 ;
        RECT 25.6 12.164 25.632 12.196 ;
  LAYER M1 ;
        RECT 25.536 9.708 25.568 12.216 ;
  LAYER M3 ;
        RECT 27.904 9.792 27.936 9.824 ;
  LAYER M2 ;
        RECT 25.536 9.856 25.568 9.888 ;
  LAYER M2 ;
        RECT 27.904 9.92 27.936 9.952 ;
  LAYER M2 ;
        RECT 25.536 9.984 25.568 10.016 ;
  LAYER M2 ;
        RECT 27.904 10.048 27.936 10.08 ;
  LAYER M2 ;
        RECT 25.536 10.112 25.568 10.144 ;
  LAYER M2 ;
        RECT 27.904 10.176 27.936 10.208 ;
  LAYER M2 ;
        RECT 25.536 10.24 25.568 10.272 ;
  LAYER M2 ;
        RECT 27.904 10.304 27.936 10.336 ;
  LAYER M2 ;
        RECT 25.536 10.368 25.568 10.4 ;
  LAYER M2 ;
        RECT 27.904 10.432 27.936 10.464 ;
  LAYER M2 ;
        RECT 25.536 10.496 25.568 10.528 ;
  LAYER M2 ;
        RECT 27.904 10.56 27.936 10.592 ;
  LAYER M2 ;
        RECT 25.536 10.624 25.568 10.656 ;
  LAYER M2 ;
        RECT 27.904 10.688 27.936 10.72 ;
  LAYER M2 ;
        RECT 25.536 10.752 25.568 10.784 ;
  LAYER M2 ;
        RECT 27.904 10.816 27.936 10.848 ;
  LAYER M2 ;
        RECT 25.536 10.88 25.568 10.912 ;
  LAYER M2 ;
        RECT 27.904 10.944 27.936 10.976 ;
  LAYER M2 ;
        RECT 25.536 11.008 25.568 11.04 ;
  LAYER M2 ;
        RECT 27.904 11.072 27.936 11.104 ;
  LAYER M2 ;
        RECT 25.536 11.136 25.568 11.168 ;
  LAYER M2 ;
        RECT 27.904 11.2 27.936 11.232 ;
  LAYER M2 ;
        RECT 25.536 11.264 25.568 11.296 ;
  LAYER M2 ;
        RECT 27.904 11.328 27.936 11.36 ;
  LAYER M2 ;
        RECT 25.536 11.392 25.568 11.424 ;
  LAYER M2 ;
        RECT 27.904 11.456 27.936 11.488 ;
  LAYER M2 ;
        RECT 25.536 11.52 25.568 11.552 ;
  LAYER M2 ;
        RECT 27.904 11.584 27.936 11.616 ;
  LAYER M2 ;
        RECT 25.536 11.648 25.568 11.68 ;
  LAYER M2 ;
        RECT 27.904 11.712 27.936 11.744 ;
  LAYER M2 ;
        RECT 25.536 11.776 25.568 11.808 ;
  LAYER M2 ;
        RECT 27.904 11.84 27.936 11.872 ;
  LAYER M2 ;
        RECT 25.536 11.904 25.568 11.936 ;
  LAYER M2 ;
        RECT 27.904 11.968 27.936 12 ;
  LAYER M2 ;
        RECT 25.536 12.032 25.568 12.064 ;
  LAYER M2 ;
        RECT 25.488 9.66 27.984 12.264 ;
  LAYER M1 ;
        RECT 27.904 12.816 27.936 15.324 ;
  LAYER M3 ;
        RECT 27.904 15.272 27.936 15.304 ;
  LAYER M1 ;
        RECT 27.84 12.816 27.872 15.324 ;
  LAYER M3 ;
        RECT 27.84 12.836 27.872 12.868 ;
  LAYER M1 ;
        RECT 27.776 12.816 27.808 15.324 ;
  LAYER M3 ;
        RECT 27.776 15.272 27.808 15.304 ;
  LAYER M1 ;
        RECT 27.712 12.816 27.744 15.324 ;
  LAYER M3 ;
        RECT 27.712 12.836 27.744 12.868 ;
  LAYER M1 ;
        RECT 27.648 12.816 27.68 15.324 ;
  LAYER M3 ;
        RECT 27.648 15.272 27.68 15.304 ;
  LAYER M1 ;
        RECT 27.584 12.816 27.616 15.324 ;
  LAYER M3 ;
        RECT 27.584 12.836 27.616 12.868 ;
  LAYER M1 ;
        RECT 27.52 12.816 27.552 15.324 ;
  LAYER M3 ;
        RECT 27.52 15.272 27.552 15.304 ;
  LAYER M1 ;
        RECT 27.456 12.816 27.488 15.324 ;
  LAYER M3 ;
        RECT 27.456 12.836 27.488 12.868 ;
  LAYER M1 ;
        RECT 27.392 12.816 27.424 15.324 ;
  LAYER M3 ;
        RECT 27.392 15.272 27.424 15.304 ;
  LAYER M1 ;
        RECT 27.328 12.816 27.36 15.324 ;
  LAYER M3 ;
        RECT 27.328 12.836 27.36 12.868 ;
  LAYER M1 ;
        RECT 27.264 12.816 27.296 15.324 ;
  LAYER M3 ;
        RECT 27.264 15.272 27.296 15.304 ;
  LAYER M1 ;
        RECT 27.2 12.816 27.232 15.324 ;
  LAYER M3 ;
        RECT 27.2 12.836 27.232 12.868 ;
  LAYER M1 ;
        RECT 27.136 12.816 27.168 15.324 ;
  LAYER M3 ;
        RECT 27.136 15.272 27.168 15.304 ;
  LAYER M1 ;
        RECT 27.072 12.816 27.104 15.324 ;
  LAYER M3 ;
        RECT 27.072 12.836 27.104 12.868 ;
  LAYER M1 ;
        RECT 27.008 12.816 27.04 15.324 ;
  LAYER M3 ;
        RECT 27.008 15.272 27.04 15.304 ;
  LAYER M1 ;
        RECT 26.944 12.816 26.976 15.324 ;
  LAYER M3 ;
        RECT 26.944 12.836 26.976 12.868 ;
  LAYER M1 ;
        RECT 26.88 12.816 26.912 15.324 ;
  LAYER M3 ;
        RECT 26.88 15.272 26.912 15.304 ;
  LAYER M1 ;
        RECT 26.816 12.816 26.848 15.324 ;
  LAYER M3 ;
        RECT 26.816 12.836 26.848 12.868 ;
  LAYER M1 ;
        RECT 26.752 12.816 26.784 15.324 ;
  LAYER M3 ;
        RECT 26.752 15.272 26.784 15.304 ;
  LAYER M1 ;
        RECT 26.688 12.816 26.72 15.324 ;
  LAYER M3 ;
        RECT 26.688 12.836 26.72 12.868 ;
  LAYER M1 ;
        RECT 26.624 12.816 26.656 15.324 ;
  LAYER M3 ;
        RECT 26.624 15.272 26.656 15.304 ;
  LAYER M1 ;
        RECT 26.56 12.816 26.592 15.324 ;
  LAYER M3 ;
        RECT 26.56 12.836 26.592 12.868 ;
  LAYER M1 ;
        RECT 26.496 12.816 26.528 15.324 ;
  LAYER M3 ;
        RECT 26.496 15.272 26.528 15.304 ;
  LAYER M1 ;
        RECT 26.432 12.816 26.464 15.324 ;
  LAYER M3 ;
        RECT 26.432 12.836 26.464 12.868 ;
  LAYER M1 ;
        RECT 26.368 12.816 26.4 15.324 ;
  LAYER M3 ;
        RECT 26.368 15.272 26.4 15.304 ;
  LAYER M1 ;
        RECT 26.304 12.816 26.336 15.324 ;
  LAYER M3 ;
        RECT 26.304 12.836 26.336 12.868 ;
  LAYER M1 ;
        RECT 26.24 12.816 26.272 15.324 ;
  LAYER M3 ;
        RECT 26.24 15.272 26.272 15.304 ;
  LAYER M1 ;
        RECT 26.176 12.816 26.208 15.324 ;
  LAYER M3 ;
        RECT 26.176 12.836 26.208 12.868 ;
  LAYER M1 ;
        RECT 26.112 12.816 26.144 15.324 ;
  LAYER M3 ;
        RECT 26.112 15.272 26.144 15.304 ;
  LAYER M1 ;
        RECT 26.048 12.816 26.08 15.324 ;
  LAYER M3 ;
        RECT 26.048 12.836 26.08 12.868 ;
  LAYER M1 ;
        RECT 25.984 12.816 26.016 15.324 ;
  LAYER M3 ;
        RECT 25.984 15.272 26.016 15.304 ;
  LAYER M1 ;
        RECT 25.92 12.816 25.952 15.324 ;
  LAYER M3 ;
        RECT 25.92 12.836 25.952 12.868 ;
  LAYER M1 ;
        RECT 25.856 12.816 25.888 15.324 ;
  LAYER M3 ;
        RECT 25.856 15.272 25.888 15.304 ;
  LAYER M1 ;
        RECT 25.792 12.816 25.824 15.324 ;
  LAYER M3 ;
        RECT 25.792 12.836 25.824 12.868 ;
  LAYER M1 ;
        RECT 25.728 12.816 25.76 15.324 ;
  LAYER M3 ;
        RECT 25.728 15.272 25.76 15.304 ;
  LAYER M1 ;
        RECT 25.664 12.816 25.696 15.324 ;
  LAYER M3 ;
        RECT 25.664 12.836 25.696 12.868 ;
  LAYER M1 ;
        RECT 25.6 12.816 25.632 15.324 ;
  LAYER M3 ;
        RECT 25.6 15.272 25.632 15.304 ;
  LAYER M1 ;
        RECT 25.536 12.816 25.568 15.324 ;
  LAYER M3 ;
        RECT 27.904 12.9 27.936 12.932 ;
  LAYER M2 ;
        RECT 25.536 12.964 25.568 12.996 ;
  LAYER M2 ;
        RECT 27.904 13.028 27.936 13.06 ;
  LAYER M2 ;
        RECT 25.536 13.092 25.568 13.124 ;
  LAYER M2 ;
        RECT 27.904 13.156 27.936 13.188 ;
  LAYER M2 ;
        RECT 25.536 13.22 25.568 13.252 ;
  LAYER M2 ;
        RECT 27.904 13.284 27.936 13.316 ;
  LAYER M2 ;
        RECT 25.536 13.348 25.568 13.38 ;
  LAYER M2 ;
        RECT 27.904 13.412 27.936 13.444 ;
  LAYER M2 ;
        RECT 25.536 13.476 25.568 13.508 ;
  LAYER M2 ;
        RECT 27.904 13.54 27.936 13.572 ;
  LAYER M2 ;
        RECT 25.536 13.604 25.568 13.636 ;
  LAYER M2 ;
        RECT 27.904 13.668 27.936 13.7 ;
  LAYER M2 ;
        RECT 25.536 13.732 25.568 13.764 ;
  LAYER M2 ;
        RECT 27.904 13.796 27.936 13.828 ;
  LAYER M2 ;
        RECT 25.536 13.86 25.568 13.892 ;
  LAYER M2 ;
        RECT 27.904 13.924 27.936 13.956 ;
  LAYER M2 ;
        RECT 25.536 13.988 25.568 14.02 ;
  LAYER M2 ;
        RECT 27.904 14.052 27.936 14.084 ;
  LAYER M2 ;
        RECT 25.536 14.116 25.568 14.148 ;
  LAYER M2 ;
        RECT 27.904 14.18 27.936 14.212 ;
  LAYER M2 ;
        RECT 25.536 14.244 25.568 14.276 ;
  LAYER M2 ;
        RECT 27.904 14.308 27.936 14.34 ;
  LAYER M2 ;
        RECT 25.536 14.372 25.568 14.404 ;
  LAYER M2 ;
        RECT 27.904 14.436 27.936 14.468 ;
  LAYER M2 ;
        RECT 25.536 14.5 25.568 14.532 ;
  LAYER M2 ;
        RECT 27.904 14.564 27.936 14.596 ;
  LAYER M2 ;
        RECT 25.536 14.628 25.568 14.66 ;
  LAYER M2 ;
        RECT 27.904 14.692 27.936 14.724 ;
  LAYER M2 ;
        RECT 25.536 14.756 25.568 14.788 ;
  LAYER M2 ;
        RECT 27.904 14.82 27.936 14.852 ;
  LAYER M2 ;
        RECT 25.536 14.884 25.568 14.916 ;
  LAYER M2 ;
        RECT 27.904 14.948 27.936 14.98 ;
  LAYER M2 ;
        RECT 25.536 15.012 25.568 15.044 ;
  LAYER M2 ;
        RECT 27.904 15.076 27.936 15.108 ;
  LAYER M2 ;
        RECT 25.536 15.14 25.568 15.172 ;
  LAYER M2 ;
        RECT 25.488 12.768 27.984 15.372 ;
  LAYER M1 ;
        RECT 27.904 15.924 27.936 18.432 ;
  LAYER M3 ;
        RECT 27.904 18.38 27.936 18.412 ;
  LAYER M1 ;
        RECT 27.84 15.924 27.872 18.432 ;
  LAYER M3 ;
        RECT 27.84 15.944 27.872 15.976 ;
  LAYER M1 ;
        RECT 27.776 15.924 27.808 18.432 ;
  LAYER M3 ;
        RECT 27.776 18.38 27.808 18.412 ;
  LAYER M1 ;
        RECT 27.712 15.924 27.744 18.432 ;
  LAYER M3 ;
        RECT 27.712 15.944 27.744 15.976 ;
  LAYER M1 ;
        RECT 27.648 15.924 27.68 18.432 ;
  LAYER M3 ;
        RECT 27.648 18.38 27.68 18.412 ;
  LAYER M1 ;
        RECT 27.584 15.924 27.616 18.432 ;
  LAYER M3 ;
        RECT 27.584 15.944 27.616 15.976 ;
  LAYER M1 ;
        RECT 27.52 15.924 27.552 18.432 ;
  LAYER M3 ;
        RECT 27.52 18.38 27.552 18.412 ;
  LAYER M1 ;
        RECT 27.456 15.924 27.488 18.432 ;
  LAYER M3 ;
        RECT 27.456 15.944 27.488 15.976 ;
  LAYER M1 ;
        RECT 27.392 15.924 27.424 18.432 ;
  LAYER M3 ;
        RECT 27.392 18.38 27.424 18.412 ;
  LAYER M1 ;
        RECT 27.328 15.924 27.36 18.432 ;
  LAYER M3 ;
        RECT 27.328 15.944 27.36 15.976 ;
  LAYER M1 ;
        RECT 27.264 15.924 27.296 18.432 ;
  LAYER M3 ;
        RECT 27.264 18.38 27.296 18.412 ;
  LAYER M1 ;
        RECT 27.2 15.924 27.232 18.432 ;
  LAYER M3 ;
        RECT 27.2 15.944 27.232 15.976 ;
  LAYER M1 ;
        RECT 27.136 15.924 27.168 18.432 ;
  LAYER M3 ;
        RECT 27.136 18.38 27.168 18.412 ;
  LAYER M1 ;
        RECT 27.072 15.924 27.104 18.432 ;
  LAYER M3 ;
        RECT 27.072 15.944 27.104 15.976 ;
  LAYER M1 ;
        RECT 27.008 15.924 27.04 18.432 ;
  LAYER M3 ;
        RECT 27.008 18.38 27.04 18.412 ;
  LAYER M1 ;
        RECT 26.944 15.924 26.976 18.432 ;
  LAYER M3 ;
        RECT 26.944 15.944 26.976 15.976 ;
  LAYER M1 ;
        RECT 26.88 15.924 26.912 18.432 ;
  LAYER M3 ;
        RECT 26.88 18.38 26.912 18.412 ;
  LAYER M1 ;
        RECT 26.816 15.924 26.848 18.432 ;
  LAYER M3 ;
        RECT 26.816 15.944 26.848 15.976 ;
  LAYER M1 ;
        RECT 26.752 15.924 26.784 18.432 ;
  LAYER M3 ;
        RECT 26.752 18.38 26.784 18.412 ;
  LAYER M1 ;
        RECT 26.688 15.924 26.72 18.432 ;
  LAYER M3 ;
        RECT 26.688 15.944 26.72 15.976 ;
  LAYER M1 ;
        RECT 26.624 15.924 26.656 18.432 ;
  LAYER M3 ;
        RECT 26.624 18.38 26.656 18.412 ;
  LAYER M1 ;
        RECT 26.56 15.924 26.592 18.432 ;
  LAYER M3 ;
        RECT 26.56 15.944 26.592 15.976 ;
  LAYER M1 ;
        RECT 26.496 15.924 26.528 18.432 ;
  LAYER M3 ;
        RECT 26.496 18.38 26.528 18.412 ;
  LAYER M1 ;
        RECT 26.432 15.924 26.464 18.432 ;
  LAYER M3 ;
        RECT 26.432 15.944 26.464 15.976 ;
  LAYER M1 ;
        RECT 26.368 15.924 26.4 18.432 ;
  LAYER M3 ;
        RECT 26.368 18.38 26.4 18.412 ;
  LAYER M1 ;
        RECT 26.304 15.924 26.336 18.432 ;
  LAYER M3 ;
        RECT 26.304 15.944 26.336 15.976 ;
  LAYER M1 ;
        RECT 26.24 15.924 26.272 18.432 ;
  LAYER M3 ;
        RECT 26.24 18.38 26.272 18.412 ;
  LAYER M1 ;
        RECT 26.176 15.924 26.208 18.432 ;
  LAYER M3 ;
        RECT 26.176 15.944 26.208 15.976 ;
  LAYER M1 ;
        RECT 26.112 15.924 26.144 18.432 ;
  LAYER M3 ;
        RECT 26.112 18.38 26.144 18.412 ;
  LAYER M1 ;
        RECT 26.048 15.924 26.08 18.432 ;
  LAYER M3 ;
        RECT 26.048 15.944 26.08 15.976 ;
  LAYER M1 ;
        RECT 25.984 15.924 26.016 18.432 ;
  LAYER M3 ;
        RECT 25.984 18.38 26.016 18.412 ;
  LAYER M1 ;
        RECT 25.92 15.924 25.952 18.432 ;
  LAYER M3 ;
        RECT 25.92 15.944 25.952 15.976 ;
  LAYER M1 ;
        RECT 25.856 15.924 25.888 18.432 ;
  LAYER M3 ;
        RECT 25.856 18.38 25.888 18.412 ;
  LAYER M1 ;
        RECT 25.792 15.924 25.824 18.432 ;
  LAYER M3 ;
        RECT 25.792 15.944 25.824 15.976 ;
  LAYER M1 ;
        RECT 25.728 15.924 25.76 18.432 ;
  LAYER M3 ;
        RECT 25.728 18.38 25.76 18.412 ;
  LAYER M1 ;
        RECT 25.664 15.924 25.696 18.432 ;
  LAYER M3 ;
        RECT 25.664 15.944 25.696 15.976 ;
  LAYER M1 ;
        RECT 25.6 15.924 25.632 18.432 ;
  LAYER M3 ;
        RECT 25.6 18.38 25.632 18.412 ;
  LAYER M1 ;
        RECT 25.536 15.924 25.568 18.432 ;
  LAYER M3 ;
        RECT 27.904 16.008 27.936 16.04 ;
  LAYER M2 ;
        RECT 25.536 16.072 25.568 16.104 ;
  LAYER M2 ;
        RECT 27.904 16.136 27.936 16.168 ;
  LAYER M2 ;
        RECT 25.536 16.2 25.568 16.232 ;
  LAYER M2 ;
        RECT 27.904 16.264 27.936 16.296 ;
  LAYER M2 ;
        RECT 25.536 16.328 25.568 16.36 ;
  LAYER M2 ;
        RECT 27.904 16.392 27.936 16.424 ;
  LAYER M2 ;
        RECT 25.536 16.456 25.568 16.488 ;
  LAYER M2 ;
        RECT 27.904 16.52 27.936 16.552 ;
  LAYER M2 ;
        RECT 25.536 16.584 25.568 16.616 ;
  LAYER M2 ;
        RECT 27.904 16.648 27.936 16.68 ;
  LAYER M2 ;
        RECT 25.536 16.712 25.568 16.744 ;
  LAYER M2 ;
        RECT 27.904 16.776 27.936 16.808 ;
  LAYER M2 ;
        RECT 25.536 16.84 25.568 16.872 ;
  LAYER M2 ;
        RECT 27.904 16.904 27.936 16.936 ;
  LAYER M2 ;
        RECT 25.536 16.968 25.568 17 ;
  LAYER M2 ;
        RECT 27.904 17.032 27.936 17.064 ;
  LAYER M2 ;
        RECT 25.536 17.096 25.568 17.128 ;
  LAYER M2 ;
        RECT 27.904 17.16 27.936 17.192 ;
  LAYER M2 ;
        RECT 25.536 17.224 25.568 17.256 ;
  LAYER M2 ;
        RECT 27.904 17.288 27.936 17.32 ;
  LAYER M2 ;
        RECT 25.536 17.352 25.568 17.384 ;
  LAYER M2 ;
        RECT 27.904 17.416 27.936 17.448 ;
  LAYER M2 ;
        RECT 25.536 17.48 25.568 17.512 ;
  LAYER M2 ;
        RECT 27.904 17.544 27.936 17.576 ;
  LAYER M2 ;
        RECT 25.536 17.608 25.568 17.64 ;
  LAYER M2 ;
        RECT 27.904 17.672 27.936 17.704 ;
  LAYER M2 ;
        RECT 25.536 17.736 25.568 17.768 ;
  LAYER M2 ;
        RECT 27.904 17.8 27.936 17.832 ;
  LAYER M2 ;
        RECT 25.536 17.864 25.568 17.896 ;
  LAYER M2 ;
        RECT 27.904 17.928 27.936 17.96 ;
  LAYER M2 ;
        RECT 25.536 17.992 25.568 18.024 ;
  LAYER M2 ;
        RECT 27.904 18.056 27.936 18.088 ;
  LAYER M2 ;
        RECT 25.536 18.12 25.568 18.152 ;
  LAYER M2 ;
        RECT 27.904 18.184 27.936 18.216 ;
  LAYER M2 ;
        RECT 25.536 18.248 25.568 18.28 ;
  LAYER M2 ;
        RECT 25.488 15.876 27.984 18.48 ;
  LAYER M1 ;
        RECT 24.928 6.6 24.96 9.108 ;
  LAYER M3 ;
        RECT 24.928 9.056 24.96 9.088 ;
  LAYER M1 ;
        RECT 24.864 6.6 24.896 9.108 ;
  LAYER M3 ;
        RECT 24.864 6.62 24.896 6.652 ;
  LAYER M1 ;
        RECT 24.8 6.6 24.832 9.108 ;
  LAYER M3 ;
        RECT 24.8 9.056 24.832 9.088 ;
  LAYER M1 ;
        RECT 24.736 6.6 24.768 9.108 ;
  LAYER M3 ;
        RECT 24.736 6.62 24.768 6.652 ;
  LAYER M1 ;
        RECT 24.672 6.6 24.704 9.108 ;
  LAYER M3 ;
        RECT 24.672 9.056 24.704 9.088 ;
  LAYER M1 ;
        RECT 24.608 6.6 24.64 9.108 ;
  LAYER M3 ;
        RECT 24.608 6.62 24.64 6.652 ;
  LAYER M1 ;
        RECT 24.544 6.6 24.576 9.108 ;
  LAYER M3 ;
        RECT 24.544 9.056 24.576 9.088 ;
  LAYER M1 ;
        RECT 24.48 6.6 24.512 9.108 ;
  LAYER M3 ;
        RECT 24.48 6.62 24.512 6.652 ;
  LAYER M1 ;
        RECT 24.416 6.6 24.448 9.108 ;
  LAYER M3 ;
        RECT 24.416 9.056 24.448 9.088 ;
  LAYER M1 ;
        RECT 24.352 6.6 24.384 9.108 ;
  LAYER M3 ;
        RECT 24.352 6.62 24.384 6.652 ;
  LAYER M1 ;
        RECT 24.288 6.6 24.32 9.108 ;
  LAYER M3 ;
        RECT 24.288 9.056 24.32 9.088 ;
  LAYER M1 ;
        RECT 24.224 6.6 24.256 9.108 ;
  LAYER M3 ;
        RECT 24.224 6.62 24.256 6.652 ;
  LAYER M1 ;
        RECT 24.16 6.6 24.192 9.108 ;
  LAYER M3 ;
        RECT 24.16 9.056 24.192 9.088 ;
  LAYER M1 ;
        RECT 24.096 6.6 24.128 9.108 ;
  LAYER M3 ;
        RECT 24.096 6.62 24.128 6.652 ;
  LAYER M1 ;
        RECT 24.032 6.6 24.064 9.108 ;
  LAYER M3 ;
        RECT 24.032 9.056 24.064 9.088 ;
  LAYER M1 ;
        RECT 23.968 6.6 24 9.108 ;
  LAYER M3 ;
        RECT 23.968 6.62 24 6.652 ;
  LAYER M1 ;
        RECT 23.904 6.6 23.936 9.108 ;
  LAYER M3 ;
        RECT 23.904 9.056 23.936 9.088 ;
  LAYER M1 ;
        RECT 23.84 6.6 23.872 9.108 ;
  LAYER M3 ;
        RECT 23.84 6.62 23.872 6.652 ;
  LAYER M1 ;
        RECT 23.776 6.6 23.808 9.108 ;
  LAYER M3 ;
        RECT 23.776 9.056 23.808 9.088 ;
  LAYER M1 ;
        RECT 23.712 6.6 23.744 9.108 ;
  LAYER M3 ;
        RECT 23.712 6.62 23.744 6.652 ;
  LAYER M1 ;
        RECT 23.648 6.6 23.68 9.108 ;
  LAYER M3 ;
        RECT 23.648 9.056 23.68 9.088 ;
  LAYER M1 ;
        RECT 23.584 6.6 23.616 9.108 ;
  LAYER M3 ;
        RECT 23.584 6.62 23.616 6.652 ;
  LAYER M1 ;
        RECT 23.52 6.6 23.552 9.108 ;
  LAYER M3 ;
        RECT 23.52 9.056 23.552 9.088 ;
  LAYER M1 ;
        RECT 23.456 6.6 23.488 9.108 ;
  LAYER M3 ;
        RECT 23.456 6.62 23.488 6.652 ;
  LAYER M1 ;
        RECT 23.392 6.6 23.424 9.108 ;
  LAYER M3 ;
        RECT 23.392 9.056 23.424 9.088 ;
  LAYER M1 ;
        RECT 23.328 6.6 23.36 9.108 ;
  LAYER M3 ;
        RECT 23.328 6.62 23.36 6.652 ;
  LAYER M1 ;
        RECT 23.264 6.6 23.296 9.108 ;
  LAYER M3 ;
        RECT 23.264 9.056 23.296 9.088 ;
  LAYER M1 ;
        RECT 23.2 6.6 23.232 9.108 ;
  LAYER M3 ;
        RECT 23.2 6.62 23.232 6.652 ;
  LAYER M1 ;
        RECT 23.136 6.6 23.168 9.108 ;
  LAYER M3 ;
        RECT 23.136 9.056 23.168 9.088 ;
  LAYER M1 ;
        RECT 23.072 6.6 23.104 9.108 ;
  LAYER M3 ;
        RECT 23.072 6.62 23.104 6.652 ;
  LAYER M1 ;
        RECT 23.008 6.6 23.04 9.108 ;
  LAYER M3 ;
        RECT 23.008 9.056 23.04 9.088 ;
  LAYER M1 ;
        RECT 22.944 6.6 22.976 9.108 ;
  LAYER M3 ;
        RECT 22.944 6.62 22.976 6.652 ;
  LAYER M1 ;
        RECT 22.88 6.6 22.912 9.108 ;
  LAYER M3 ;
        RECT 22.88 9.056 22.912 9.088 ;
  LAYER M1 ;
        RECT 22.816 6.6 22.848 9.108 ;
  LAYER M3 ;
        RECT 22.816 6.62 22.848 6.652 ;
  LAYER M1 ;
        RECT 22.752 6.6 22.784 9.108 ;
  LAYER M3 ;
        RECT 22.752 9.056 22.784 9.088 ;
  LAYER M1 ;
        RECT 22.688 6.6 22.72 9.108 ;
  LAYER M3 ;
        RECT 22.688 6.62 22.72 6.652 ;
  LAYER M1 ;
        RECT 22.624 6.6 22.656 9.108 ;
  LAYER M3 ;
        RECT 22.624 9.056 22.656 9.088 ;
  LAYER M1 ;
        RECT 22.56 6.6 22.592 9.108 ;
  LAYER M3 ;
        RECT 24.928 6.684 24.96 6.716 ;
  LAYER M2 ;
        RECT 22.56 6.748 22.592 6.78 ;
  LAYER M2 ;
        RECT 24.928 6.812 24.96 6.844 ;
  LAYER M2 ;
        RECT 22.56 6.876 22.592 6.908 ;
  LAYER M2 ;
        RECT 24.928 6.94 24.96 6.972 ;
  LAYER M2 ;
        RECT 22.56 7.004 22.592 7.036 ;
  LAYER M2 ;
        RECT 24.928 7.068 24.96 7.1 ;
  LAYER M2 ;
        RECT 22.56 7.132 22.592 7.164 ;
  LAYER M2 ;
        RECT 24.928 7.196 24.96 7.228 ;
  LAYER M2 ;
        RECT 22.56 7.26 22.592 7.292 ;
  LAYER M2 ;
        RECT 24.928 7.324 24.96 7.356 ;
  LAYER M2 ;
        RECT 22.56 7.388 22.592 7.42 ;
  LAYER M2 ;
        RECT 24.928 7.452 24.96 7.484 ;
  LAYER M2 ;
        RECT 22.56 7.516 22.592 7.548 ;
  LAYER M2 ;
        RECT 24.928 7.58 24.96 7.612 ;
  LAYER M2 ;
        RECT 22.56 7.644 22.592 7.676 ;
  LAYER M2 ;
        RECT 24.928 7.708 24.96 7.74 ;
  LAYER M2 ;
        RECT 22.56 7.772 22.592 7.804 ;
  LAYER M2 ;
        RECT 24.928 7.836 24.96 7.868 ;
  LAYER M2 ;
        RECT 22.56 7.9 22.592 7.932 ;
  LAYER M2 ;
        RECT 24.928 7.964 24.96 7.996 ;
  LAYER M2 ;
        RECT 22.56 8.028 22.592 8.06 ;
  LAYER M2 ;
        RECT 24.928 8.092 24.96 8.124 ;
  LAYER M2 ;
        RECT 22.56 8.156 22.592 8.188 ;
  LAYER M2 ;
        RECT 24.928 8.22 24.96 8.252 ;
  LAYER M2 ;
        RECT 22.56 8.284 22.592 8.316 ;
  LAYER M2 ;
        RECT 24.928 8.348 24.96 8.38 ;
  LAYER M2 ;
        RECT 22.56 8.412 22.592 8.444 ;
  LAYER M2 ;
        RECT 24.928 8.476 24.96 8.508 ;
  LAYER M2 ;
        RECT 22.56 8.54 22.592 8.572 ;
  LAYER M2 ;
        RECT 24.928 8.604 24.96 8.636 ;
  LAYER M2 ;
        RECT 22.56 8.668 22.592 8.7 ;
  LAYER M2 ;
        RECT 24.928 8.732 24.96 8.764 ;
  LAYER M2 ;
        RECT 22.56 8.796 22.592 8.828 ;
  LAYER M2 ;
        RECT 24.928 8.86 24.96 8.892 ;
  LAYER M2 ;
        RECT 22.56 8.924 22.592 8.956 ;
  LAYER M2 ;
        RECT 22.512 6.552 25.008 9.156 ;
  LAYER M1 ;
        RECT 24.928 9.708 24.96 12.216 ;
  LAYER M3 ;
        RECT 24.928 12.164 24.96 12.196 ;
  LAYER M1 ;
        RECT 24.864 9.708 24.896 12.216 ;
  LAYER M3 ;
        RECT 24.864 9.728 24.896 9.76 ;
  LAYER M1 ;
        RECT 24.8 9.708 24.832 12.216 ;
  LAYER M3 ;
        RECT 24.8 12.164 24.832 12.196 ;
  LAYER M1 ;
        RECT 24.736 9.708 24.768 12.216 ;
  LAYER M3 ;
        RECT 24.736 9.728 24.768 9.76 ;
  LAYER M1 ;
        RECT 24.672 9.708 24.704 12.216 ;
  LAYER M3 ;
        RECT 24.672 12.164 24.704 12.196 ;
  LAYER M1 ;
        RECT 24.608 9.708 24.64 12.216 ;
  LAYER M3 ;
        RECT 24.608 9.728 24.64 9.76 ;
  LAYER M1 ;
        RECT 24.544 9.708 24.576 12.216 ;
  LAYER M3 ;
        RECT 24.544 12.164 24.576 12.196 ;
  LAYER M1 ;
        RECT 24.48 9.708 24.512 12.216 ;
  LAYER M3 ;
        RECT 24.48 9.728 24.512 9.76 ;
  LAYER M1 ;
        RECT 24.416 9.708 24.448 12.216 ;
  LAYER M3 ;
        RECT 24.416 12.164 24.448 12.196 ;
  LAYER M1 ;
        RECT 24.352 9.708 24.384 12.216 ;
  LAYER M3 ;
        RECT 24.352 9.728 24.384 9.76 ;
  LAYER M1 ;
        RECT 24.288 9.708 24.32 12.216 ;
  LAYER M3 ;
        RECT 24.288 12.164 24.32 12.196 ;
  LAYER M1 ;
        RECT 24.224 9.708 24.256 12.216 ;
  LAYER M3 ;
        RECT 24.224 9.728 24.256 9.76 ;
  LAYER M1 ;
        RECT 24.16 9.708 24.192 12.216 ;
  LAYER M3 ;
        RECT 24.16 12.164 24.192 12.196 ;
  LAYER M1 ;
        RECT 24.096 9.708 24.128 12.216 ;
  LAYER M3 ;
        RECT 24.096 9.728 24.128 9.76 ;
  LAYER M1 ;
        RECT 24.032 9.708 24.064 12.216 ;
  LAYER M3 ;
        RECT 24.032 12.164 24.064 12.196 ;
  LAYER M1 ;
        RECT 23.968 9.708 24 12.216 ;
  LAYER M3 ;
        RECT 23.968 9.728 24 9.76 ;
  LAYER M1 ;
        RECT 23.904 9.708 23.936 12.216 ;
  LAYER M3 ;
        RECT 23.904 12.164 23.936 12.196 ;
  LAYER M1 ;
        RECT 23.84 9.708 23.872 12.216 ;
  LAYER M3 ;
        RECT 23.84 9.728 23.872 9.76 ;
  LAYER M1 ;
        RECT 23.776 9.708 23.808 12.216 ;
  LAYER M3 ;
        RECT 23.776 12.164 23.808 12.196 ;
  LAYER M1 ;
        RECT 23.712 9.708 23.744 12.216 ;
  LAYER M3 ;
        RECT 23.712 9.728 23.744 9.76 ;
  LAYER M1 ;
        RECT 23.648 9.708 23.68 12.216 ;
  LAYER M3 ;
        RECT 23.648 12.164 23.68 12.196 ;
  LAYER M1 ;
        RECT 23.584 9.708 23.616 12.216 ;
  LAYER M3 ;
        RECT 23.584 9.728 23.616 9.76 ;
  LAYER M1 ;
        RECT 23.52 9.708 23.552 12.216 ;
  LAYER M3 ;
        RECT 23.52 12.164 23.552 12.196 ;
  LAYER M1 ;
        RECT 23.456 9.708 23.488 12.216 ;
  LAYER M3 ;
        RECT 23.456 9.728 23.488 9.76 ;
  LAYER M1 ;
        RECT 23.392 9.708 23.424 12.216 ;
  LAYER M3 ;
        RECT 23.392 12.164 23.424 12.196 ;
  LAYER M1 ;
        RECT 23.328 9.708 23.36 12.216 ;
  LAYER M3 ;
        RECT 23.328 9.728 23.36 9.76 ;
  LAYER M1 ;
        RECT 23.264 9.708 23.296 12.216 ;
  LAYER M3 ;
        RECT 23.264 12.164 23.296 12.196 ;
  LAYER M1 ;
        RECT 23.2 9.708 23.232 12.216 ;
  LAYER M3 ;
        RECT 23.2 9.728 23.232 9.76 ;
  LAYER M1 ;
        RECT 23.136 9.708 23.168 12.216 ;
  LAYER M3 ;
        RECT 23.136 12.164 23.168 12.196 ;
  LAYER M1 ;
        RECT 23.072 9.708 23.104 12.216 ;
  LAYER M3 ;
        RECT 23.072 9.728 23.104 9.76 ;
  LAYER M1 ;
        RECT 23.008 9.708 23.04 12.216 ;
  LAYER M3 ;
        RECT 23.008 12.164 23.04 12.196 ;
  LAYER M1 ;
        RECT 22.944 9.708 22.976 12.216 ;
  LAYER M3 ;
        RECT 22.944 9.728 22.976 9.76 ;
  LAYER M1 ;
        RECT 22.88 9.708 22.912 12.216 ;
  LAYER M3 ;
        RECT 22.88 12.164 22.912 12.196 ;
  LAYER M1 ;
        RECT 22.816 9.708 22.848 12.216 ;
  LAYER M3 ;
        RECT 22.816 9.728 22.848 9.76 ;
  LAYER M1 ;
        RECT 22.752 9.708 22.784 12.216 ;
  LAYER M3 ;
        RECT 22.752 12.164 22.784 12.196 ;
  LAYER M1 ;
        RECT 22.688 9.708 22.72 12.216 ;
  LAYER M3 ;
        RECT 22.688 9.728 22.72 9.76 ;
  LAYER M1 ;
        RECT 22.624 9.708 22.656 12.216 ;
  LAYER M3 ;
        RECT 22.624 12.164 22.656 12.196 ;
  LAYER M1 ;
        RECT 22.56 9.708 22.592 12.216 ;
  LAYER M3 ;
        RECT 24.928 9.792 24.96 9.824 ;
  LAYER M2 ;
        RECT 22.56 9.856 22.592 9.888 ;
  LAYER M2 ;
        RECT 24.928 9.92 24.96 9.952 ;
  LAYER M2 ;
        RECT 22.56 9.984 22.592 10.016 ;
  LAYER M2 ;
        RECT 24.928 10.048 24.96 10.08 ;
  LAYER M2 ;
        RECT 22.56 10.112 22.592 10.144 ;
  LAYER M2 ;
        RECT 24.928 10.176 24.96 10.208 ;
  LAYER M2 ;
        RECT 22.56 10.24 22.592 10.272 ;
  LAYER M2 ;
        RECT 24.928 10.304 24.96 10.336 ;
  LAYER M2 ;
        RECT 22.56 10.368 22.592 10.4 ;
  LAYER M2 ;
        RECT 24.928 10.432 24.96 10.464 ;
  LAYER M2 ;
        RECT 22.56 10.496 22.592 10.528 ;
  LAYER M2 ;
        RECT 24.928 10.56 24.96 10.592 ;
  LAYER M2 ;
        RECT 22.56 10.624 22.592 10.656 ;
  LAYER M2 ;
        RECT 24.928 10.688 24.96 10.72 ;
  LAYER M2 ;
        RECT 22.56 10.752 22.592 10.784 ;
  LAYER M2 ;
        RECT 24.928 10.816 24.96 10.848 ;
  LAYER M2 ;
        RECT 22.56 10.88 22.592 10.912 ;
  LAYER M2 ;
        RECT 24.928 10.944 24.96 10.976 ;
  LAYER M2 ;
        RECT 22.56 11.008 22.592 11.04 ;
  LAYER M2 ;
        RECT 24.928 11.072 24.96 11.104 ;
  LAYER M2 ;
        RECT 22.56 11.136 22.592 11.168 ;
  LAYER M2 ;
        RECT 24.928 11.2 24.96 11.232 ;
  LAYER M2 ;
        RECT 22.56 11.264 22.592 11.296 ;
  LAYER M2 ;
        RECT 24.928 11.328 24.96 11.36 ;
  LAYER M2 ;
        RECT 22.56 11.392 22.592 11.424 ;
  LAYER M2 ;
        RECT 24.928 11.456 24.96 11.488 ;
  LAYER M2 ;
        RECT 22.56 11.52 22.592 11.552 ;
  LAYER M2 ;
        RECT 24.928 11.584 24.96 11.616 ;
  LAYER M2 ;
        RECT 22.56 11.648 22.592 11.68 ;
  LAYER M2 ;
        RECT 24.928 11.712 24.96 11.744 ;
  LAYER M2 ;
        RECT 22.56 11.776 22.592 11.808 ;
  LAYER M2 ;
        RECT 24.928 11.84 24.96 11.872 ;
  LAYER M2 ;
        RECT 22.56 11.904 22.592 11.936 ;
  LAYER M2 ;
        RECT 24.928 11.968 24.96 12 ;
  LAYER M2 ;
        RECT 22.56 12.032 22.592 12.064 ;
  LAYER M2 ;
        RECT 22.512 9.66 25.008 12.264 ;
  LAYER M1 ;
        RECT 24.928 12.816 24.96 15.324 ;
  LAYER M3 ;
        RECT 24.928 15.272 24.96 15.304 ;
  LAYER M1 ;
        RECT 24.864 12.816 24.896 15.324 ;
  LAYER M3 ;
        RECT 24.864 12.836 24.896 12.868 ;
  LAYER M1 ;
        RECT 24.8 12.816 24.832 15.324 ;
  LAYER M3 ;
        RECT 24.8 15.272 24.832 15.304 ;
  LAYER M1 ;
        RECT 24.736 12.816 24.768 15.324 ;
  LAYER M3 ;
        RECT 24.736 12.836 24.768 12.868 ;
  LAYER M1 ;
        RECT 24.672 12.816 24.704 15.324 ;
  LAYER M3 ;
        RECT 24.672 15.272 24.704 15.304 ;
  LAYER M1 ;
        RECT 24.608 12.816 24.64 15.324 ;
  LAYER M3 ;
        RECT 24.608 12.836 24.64 12.868 ;
  LAYER M1 ;
        RECT 24.544 12.816 24.576 15.324 ;
  LAYER M3 ;
        RECT 24.544 15.272 24.576 15.304 ;
  LAYER M1 ;
        RECT 24.48 12.816 24.512 15.324 ;
  LAYER M3 ;
        RECT 24.48 12.836 24.512 12.868 ;
  LAYER M1 ;
        RECT 24.416 12.816 24.448 15.324 ;
  LAYER M3 ;
        RECT 24.416 15.272 24.448 15.304 ;
  LAYER M1 ;
        RECT 24.352 12.816 24.384 15.324 ;
  LAYER M3 ;
        RECT 24.352 12.836 24.384 12.868 ;
  LAYER M1 ;
        RECT 24.288 12.816 24.32 15.324 ;
  LAYER M3 ;
        RECT 24.288 15.272 24.32 15.304 ;
  LAYER M1 ;
        RECT 24.224 12.816 24.256 15.324 ;
  LAYER M3 ;
        RECT 24.224 12.836 24.256 12.868 ;
  LAYER M1 ;
        RECT 24.16 12.816 24.192 15.324 ;
  LAYER M3 ;
        RECT 24.16 15.272 24.192 15.304 ;
  LAYER M1 ;
        RECT 24.096 12.816 24.128 15.324 ;
  LAYER M3 ;
        RECT 24.096 12.836 24.128 12.868 ;
  LAYER M1 ;
        RECT 24.032 12.816 24.064 15.324 ;
  LAYER M3 ;
        RECT 24.032 15.272 24.064 15.304 ;
  LAYER M1 ;
        RECT 23.968 12.816 24 15.324 ;
  LAYER M3 ;
        RECT 23.968 12.836 24 12.868 ;
  LAYER M1 ;
        RECT 23.904 12.816 23.936 15.324 ;
  LAYER M3 ;
        RECT 23.904 15.272 23.936 15.304 ;
  LAYER M1 ;
        RECT 23.84 12.816 23.872 15.324 ;
  LAYER M3 ;
        RECT 23.84 12.836 23.872 12.868 ;
  LAYER M1 ;
        RECT 23.776 12.816 23.808 15.324 ;
  LAYER M3 ;
        RECT 23.776 15.272 23.808 15.304 ;
  LAYER M1 ;
        RECT 23.712 12.816 23.744 15.324 ;
  LAYER M3 ;
        RECT 23.712 12.836 23.744 12.868 ;
  LAYER M1 ;
        RECT 23.648 12.816 23.68 15.324 ;
  LAYER M3 ;
        RECT 23.648 15.272 23.68 15.304 ;
  LAYER M1 ;
        RECT 23.584 12.816 23.616 15.324 ;
  LAYER M3 ;
        RECT 23.584 12.836 23.616 12.868 ;
  LAYER M1 ;
        RECT 23.52 12.816 23.552 15.324 ;
  LAYER M3 ;
        RECT 23.52 15.272 23.552 15.304 ;
  LAYER M1 ;
        RECT 23.456 12.816 23.488 15.324 ;
  LAYER M3 ;
        RECT 23.456 12.836 23.488 12.868 ;
  LAYER M1 ;
        RECT 23.392 12.816 23.424 15.324 ;
  LAYER M3 ;
        RECT 23.392 15.272 23.424 15.304 ;
  LAYER M1 ;
        RECT 23.328 12.816 23.36 15.324 ;
  LAYER M3 ;
        RECT 23.328 12.836 23.36 12.868 ;
  LAYER M1 ;
        RECT 23.264 12.816 23.296 15.324 ;
  LAYER M3 ;
        RECT 23.264 15.272 23.296 15.304 ;
  LAYER M1 ;
        RECT 23.2 12.816 23.232 15.324 ;
  LAYER M3 ;
        RECT 23.2 12.836 23.232 12.868 ;
  LAYER M1 ;
        RECT 23.136 12.816 23.168 15.324 ;
  LAYER M3 ;
        RECT 23.136 15.272 23.168 15.304 ;
  LAYER M1 ;
        RECT 23.072 12.816 23.104 15.324 ;
  LAYER M3 ;
        RECT 23.072 12.836 23.104 12.868 ;
  LAYER M1 ;
        RECT 23.008 12.816 23.04 15.324 ;
  LAYER M3 ;
        RECT 23.008 15.272 23.04 15.304 ;
  LAYER M1 ;
        RECT 22.944 12.816 22.976 15.324 ;
  LAYER M3 ;
        RECT 22.944 12.836 22.976 12.868 ;
  LAYER M1 ;
        RECT 22.88 12.816 22.912 15.324 ;
  LAYER M3 ;
        RECT 22.88 15.272 22.912 15.304 ;
  LAYER M1 ;
        RECT 22.816 12.816 22.848 15.324 ;
  LAYER M3 ;
        RECT 22.816 12.836 22.848 12.868 ;
  LAYER M1 ;
        RECT 22.752 12.816 22.784 15.324 ;
  LAYER M3 ;
        RECT 22.752 15.272 22.784 15.304 ;
  LAYER M1 ;
        RECT 22.688 12.816 22.72 15.324 ;
  LAYER M3 ;
        RECT 22.688 12.836 22.72 12.868 ;
  LAYER M1 ;
        RECT 22.624 12.816 22.656 15.324 ;
  LAYER M3 ;
        RECT 22.624 15.272 22.656 15.304 ;
  LAYER M1 ;
        RECT 22.56 12.816 22.592 15.324 ;
  LAYER M3 ;
        RECT 24.928 12.9 24.96 12.932 ;
  LAYER M2 ;
        RECT 22.56 12.964 22.592 12.996 ;
  LAYER M2 ;
        RECT 24.928 13.028 24.96 13.06 ;
  LAYER M2 ;
        RECT 22.56 13.092 22.592 13.124 ;
  LAYER M2 ;
        RECT 24.928 13.156 24.96 13.188 ;
  LAYER M2 ;
        RECT 22.56 13.22 22.592 13.252 ;
  LAYER M2 ;
        RECT 24.928 13.284 24.96 13.316 ;
  LAYER M2 ;
        RECT 22.56 13.348 22.592 13.38 ;
  LAYER M2 ;
        RECT 24.928 13.412 24.96 13.444 ;
  LAYER M2 ;
        RECT 22.56 13.476 22.592 13.508 ;
  LAYER M2 ;
        RECT 24.928 13.54 24.96 13.572 ;
  LAYER M2 ;
        RECT 22.56 13.604 22.592 13.636 ;
  LAYER M2 ;
        RECT 24.928 13.668 24.96 13.7 ;
  LAYER M2 ;
        RECT 22.56 13.732 22.592 13.764 ;
  LAYER M2 ;
        RECT 24.928 13.796 24.96 13.828 ;
  LAYER M2 ;
        RECT 22.56 13.86 22.592 13.892 ;
  LAYER M2 ;
        RECT 24.928 13.924 24.96 13.956 ;
  LAYER M2 ;
        RECT 22.56 13.988 22.592 14.02 ;
  LAYER M2 ;
        RECT 24.928 14.052 24.96 14.084 ;
  LAYER M2 ;
        RECT 22.56 14.116 22.592 14.148 ;
  LAYER M2 ;
        RECT 24.928 14.18 24.96 14.212 ;
  LAYER M2 ;
        RECT 22.56 14.244 22.592 14.276 ;
  LAYER M2 ;
        RECT 24.928 14.308 24.96 14.34 ;
  LAYER M2 ;
        RECT 22.56 14.372 22.592 14.404 ;
  LAYER M2 ;
        RECT 24.928 14.436 24.96 14.468 ;
  LAYER M2 ;
        RECT 22.56 14.5 22.592 14.532 ;
  LAYER M2 ;
        RECT 24.928 14.564 24.96 14.596 ;
  LAYER M2 ;
        RECT 22.56 14.628 22.592 14.66 ;
  LAYER M2 ;
        RECT 24.928 14.692 24.96 14.724 ;
  LAYER M2 ;
        RECT 22.56 14.756 22.592 14.788 ;
  LAYER M2 ;
        RECT 24.928 14.82 24.96 14.852 ;
  LAYER M2 ;
        RECT 22.56 14.884 22.592 14.916 ;
  LAYER M2 ;
        RECT 24.928 14.948 24.96 14.98 ;
  LAYER M2 ;
        RECT 22.56 15.012 22.592 15.044 ;
  LAYER M2 ;
        RECT 24.928 15.076 24.96 15.108 ;
  LAYER M2 ;
        RECT 22.56 15.14 22.592 15.172 ;
  LAYER M2 ;
        RECT 22.512 12.768 25.008 15.372 ;
  LAYER M1 ;
        RECT 24.928 15.924 24.96 18.432 ;
  LAYER M3 ;
        RECT 24.928 18.38 24.96 18.412 ;
  LAYER M1 ;
        RECT 24.864 15.924 24.896 18.432 ;
  LAYER M3 ;
        RECT 24.864 15.944 24.896 15.976 ;
  LAYER M1 ;
        RECT 24.8 15.924 24.832 18.432 ;
  LAYER M3 ;
        RECT 24.8 18.38 24.832 18.412 ;
  LAYER M1 ;
        RECT 24.736 15.924 24.768 18.432 ;
  LAYER M3 ;
        RECT 24.736 15.944 24.768 15.976 ;
  LAYER M1 ;
        RECT 24.672 15.924 24.704 18.432 ;
  LAYER M3 ;
        RECT 24.672 18.38 24.704 18.412 ;
  LAYER M1 ;
        RECT 24.608 15.924 24.64 18.432 ;
  LAYER M3 ;
        RECT 24.608 15.944 24.64 15.976 ;
  LAYER M1 ;
        RECT 24.544 15.924 24.576 18.432 ;
  LAYER M3 ;
        RECT 24.544 18.38 24.576 18.412 ;
  LAYER M1 ;
        RECT 24.48 15.924 24.512 18.432 ;
  LAYER M3 ;
        RECT 24.48 15.944 24.512 15.976 ;
  LAYER M1 ;
        RECT 24.416 15.924 24.448 18.432 ;
  LAYER M3 ;
        RECT 24.416 18.38 24.448 18.412 ;
  LAYER M1 ;
        RECT 24.352 15.924 24.384 18.432 ;
  LAYER M3 ;
        RECT 24.352 15.944 24.384 15.976 ;
  LAYER M1 ;
        RECT 24.288 15.924 24.32 18.432 ;
  LAYER M3 ;
        RECT 24.288 18.38 24.32 18.412 ;
  LAYER M1 ;
        RECT 24.224 15.924 24.256 18.432 ;
  LAYER M3 ;
        RECT 24.224 15.944 24.256 15.976 ;
  LAYER M1 ;
        RECT 24.16 15.924 24.192 18.432 ;
  LAYER M3 ;
        RECT 24.16 18.38 24.192 18.412 ;
  LAYER M1 ;
        RECT 24.096 15.924 24.128 18.432 ;
  LAYER M3 ;
        RECT 24.096 15.944 24.128 15.976 ;
  LAYER M1 ;
        RECT 24.032 15.924 24.064 18.432 ;
  LAYER M3 ;
        RECT 24.032 18.38 24.064 18.412 ;
  LAYER M1 ;
        RECT 23.968 15.924 24 18.432 ;
  LAYER M3 ;
        RECT 23.968 15.944 24 15.976 ;
  LAYER M1 ;
        RECT 23.904 15.924 23.936 18.432 ;
  LAYER M3 ;
        RECT 23.904 18.38 23.936 18.412 ;
  LAYER M1 ;
        RECT 23.84 15.924 23.872 18.432 ;
  LAYER M3 ;
        RECT 23.84 15.944 23.872 15.976 ;
  LAYER M1 ;
        RECT 23.776 15.924 23.808 18.432 ;
  LAYER M3 ;
        RECT 23.776 18.38 23.808 18.412 ;
  LAYER M1 ;
        RECT 23.712 15.924 23.744 18.432 ;
  LAYER M3 ;
        RECT 23.712 15.944 23.744 15.976 ;
  LAYER M1 ;
        RECT 23.648 15.924 23.68 18.432 ;
  LAYER M3 ;
        RECT 23.648 18.38 23.68 18.412 ;
  LAYER M1 ;
        RECT 23.584 15.924 23.616 18.432 ;
  LAYER M3 ;
        RECT 23.584 15.944 23.616 15.976 ;
  LAYER M1 ;
        RECT 23.52 15.924 23.552 18.432 ;
  LAYER M3 ;
        RECT 23.52 18.38 23.552 18.412 ;
  LAYER M1 ;
        RECT 23.456 15.924 23.488 18.432 ;
  LAYER M3 ;
        RECT 23.456 15.944 23.488 15.976 ;
  LAYER M1 ;
        RECT 23.392 15.924 23.424 18.432 ;
  LAYER M3 ;
        RECT 23.392 18.38 23.424 18.412 ;
  LAYER M1 ;
        RECT 23.328 15.924 23.36 18.432 ;
  LAYER M3 ;
        RECT 23.328 15.944 23.36 15.976 ;
  LAYER M1 ;
        RECT 23.264 15.924 23.296 18.432 ;
  LAYER M3 ;
        RECT 23.264 18.38 23.296 18.412 ;
  LAYER M1 ;
        RECT 23.2 15.924 23.232 18.432 ;
  LAYER M3 ;
        RECT 23.2 15.944 23.232 15.976 ;
  LAYER M1 ;
        RECT 23.136 15.924 23.168 18.432 ;
  LAYER M3 ;
        RECT 23.136 18.38 23.168 18.412 ;
  LAYER M1 ;
        RECT 23.072 15.924 23.104 18.432 ;
  LAYER M3 ;
        RECT 23.072 15.944 23.104 15.976 ;
  LAYER M1 ;
        RECT 23.008 15.924 23.04 18.432 ;
  LAYER M3 ;
        RECT 23.008 18.38 23.04 18.412 ;
  LAYER M1 ;
        RECT 22.944 15.924 22.976 18.432 ;
  LAYER M3 ;
        RECT 22.944 15.944 22.976 15.976 ;
  LAYER M1 ;
        RECT 22.88 15.924 22.912 18.432 ;
  LAYER M3 ;
        RECT 22.88 18.38 22.912 18.412 ;
  LAYER M1 ;
        RECT 22.816 15.924 22.848 18.432 ;
  LAYER M3 ;
        RECT 22.816 15.944 22.848 15.976 ;
  LAYER M1 ;
        RECT 22.752 15.924 22.784 18.432 ;
  LAYER M3 ;
        RECT 22.752 18.38 22.784 18.412 ;
  LAYER M1 ;
        RECT 22.688 15.924 22.72 18.432 ;
  LAYER M3 ;
        RECT 22.688 15.944 22.72 15.976 ;
  LAYER M1 ;
        RECT 22.624 15.924 22.656 18.432 ;
  LAYER M3 ;
        RECT 22.624 18.38 22.656 18.412 ;
  LAYER M1 ;
        RECT 22.56 15.924 22.592 18.432 ;
  LAYER M3 ;
        RECT 24.928 16.008 24.96 16.04 ;
  LAYER M2 ;
        RECT 22.56 16.072 22.592 16.104 ;
  LAYER M2 ;
        RECT 24.928 16.136 24.96 16.168 ;
  LAYER M2 ;
        RECT 22.56 16.2 22.592 16.232 ;
  LAYER M2 ;
        RECT 24.928 16.264 24.96 16.296 ;
  LAYER M2 ;
        RECT 22.56 16.328 22.592 16.36 ;
  LAYER M2 ;
        RECT 24.928 16.392 24.96 16.424 ;
  LAYER M2 ;
        RECT 22.56 16.456 22.592 16.488 ;
  LAYER M2 ;
        RECT 24.928 16.52 24.96 16.552 ;
  LAYER M2 ;
        RECT 22.56 16.584 22.592 16.616 ;
  LAYER M2 ;
        RECT 24.928 16.648 24.96 16.68 ;
  LAYER M2 ;
        RECT 22.56 16.712 22.592 16.744 ;
  LAYER M2 ;
        RECT 24.928 16.776 24.96 16.808 ;
  LAYER M2 ;
        RECT 22.56 16.84 22.592 16.872 ;
  LAYER M2 ;
        RECT 24.928 16.904 24.96 16.936 ;
  LAYER M2 ;
        RECT 22.56 16.968 22.592 17 ;
  LAYER M2 ;
        RECT 24.928 17.032 24.96 17.064 ;
  LAYER M2 ;
        RECT 22.56 17.096 22.592 17.128 ;
  LAYER M2 ;
        RECT 24.928 17.16 24.96 17.192 ;
  LAYER M2 ;
        RECT 22.56 17.224 22.592 17.256 ;
  LAYER M2 ;
        RECT 24.928 17.288 24.96 17.32 ;
  LAYER M2 ;
        RECT 22.56 17.352 22.592 17.384 ;
  LAYER M2 ;
        RECT 24.928 17.416 24.96 17.448 ;
  LAYER M2 ;
        RECT 22.56 17.48 22.592 17.512 ;
  LAYER M2 ;
        RECT 24.928 17.544 24.96 17.576 ;
  LAYER M2 ;
        RECT 22.56 17.608 22.592 17.64 ;
  LAYER M2 ;
        RECT 24.928 17.672 24.96 17.704 ;
  LAYER M2 ;
        RECT 22.56 17.736 22.592 17.768 ;
  LAYER M2 ;
        RECT 24.928 17.8 24.96 17.832 ;
  LAYER M2 ;
        RECT 22.56 17.864 22.592 17.896 ;
  LAYER M2 ;
        RECT 24.928 17.928 24.96 17.96 ;
  LAYER M2 ;
        RECT 22.56 17.992 22.592 18.024 ;
  LAYER M2 ;
        RECT 24.928 18.056 24.96 18.088 ;
  LAYER M2 ;
        RECT 22.56 18.12 22.592 18.152 ;
  LAYER M2 ;
        RECT 24.928 18.184 24.96 18.216 ;
  LAYER M2 ;
        RECT 22.56 18.248 22.592 18.28 ;
  LAYER M2 ;
        RECT 22.512 15.876 25.008 18.48 ;
  LAYER M1 ;
        RECT 21.952 6.6 21.984 9.108 ;
  LAYER M3 ;
        RECT 21.952 9.056 21.984 9.088 ;
  LAYER M1 ;
        RECT 21.888 6.6 21.92 9.108 ;
  LAYER M3 ;
        RECT 21.888 6.62 21.92 6.652 ;
  LAYER M1 ;
        RECT 21.824 6.6 21.856 9.108 ;
  LAYER M3 ;
        RECT 21.824 9.056 21.856 9.088 ;
  LAYER M1 ;
        RECT 21.76 6.6 21.792 9.108 ;
  LAYER M3 ;
        RECT 21.76 6.62 21.792 6.652 ;
  LAYER M1 ;
        RECT 21.696 6.6 21.728 9.108 ;
  LAYER M3 ;
        RECT 21.696 9.056 21.728 9.088 ;
  LAYER M1 ;
        RECT 21.632 6.6 21.664 9.108 ;
  LAYER M3 ;
        RECT 21.632 6.62 21.664 6.652 ;
  LAYER M1 ;
        RECT 21.568 6.6 21.6 9.108 ;
  LAYER M3 ;
        RECT 21.568 9.056 21.6 9.088 ;
  LAYER M1 ;
        RECT 21.504 6.6 21.536 9.108 ;
  LAYER M3 ;
        RECT 21.504 6.62 21.536 6.652 ;
  LAYER M1 ;
        RECT 21.44 6.6 21.472 9.108 ;
  LAYER M3 ;
        RECT 21.44 9.056 21.472 9.088 ;
  LAYER M1 ;
        RECT 21.376 6.6 21.408 9.108 ;
  LAYER M3 ;
        RECT 21.376 6.62 21.408 6.652 ;
  LAYER M1 ;
        RECT 21.312 6.6 21.344 9.108 ;
  LAYER M3 ;
        RECT 21.312 9.056 21.344 9.088 ;
  LAYER M1 ;
        RECT 21.248 6.6 21.28 9.108 ;
  LAYER M3 ;
        RECT 21.248 6.62 21.28 6.652 ;
  LAYER M1 ;
        RECT 21.184 6.6 21.216 9.108 ;
  LAYER M3 ;
        RECT 21.184 9.056 21.216 9.088 ;
  LAYER M1 ;
        RECT 21.12 6.6 21.152 9.108 ;
  LAYER M3 ;
        RECT 21.12 6.62 21.152 6.652 ;
  LAYER M1 ;
        RECT 21.056 6.6 21.088 9.108 ;
  LAYER M3 ;
        RECT 21.056 9.056 21.088 9.088 ;
  LAYER M1 ;
        RECT 20.992 6.6 21.024 9.108 ;
  LAYER M3 ;
        RECT 20.992 6.62 21.024 6.652 ;
  LAYER M1 ;
        RECT 20.928 6.6 20.96 9.108 ;
  LAYER M3 ;
        RECT 20.928 9.056 20.96 9.088 ;
  LAYER M1 ;
        RECT 20.864 6.6 20.896 9.108 ;
  LAYER M3 ;
        RECT 20.864 6.62 20.896 6.652 ;
  LAYER M1 ;
        RECT 20.8 6.6 20.832 9.108 ;
  LAYER M3 ;
        RECT 20.8 9.056 20.832 9.088 ;
  LAYER M1 ;
        RECT 20.736 6.6 20.768 9.108 ;
  LAYER M3 ;
        RECT 20.736 6.62 20.768 6.652 ;
  LAYER M1 ;
        RECT 20.672 6.6 20.704 9.108 ;
  LAYER M3 ;
        RECT 20.672 9.056 20.704 9.088 ;
  LAYER M1 ;
        RECT 20.608 6.6 20.64 9.108 ;
  LAYER M3 ;
        RECT 20.608 6.62 20.64 6.652 ;
  LAYER M1 ;
        RECT 20.544 6.6 20.576 9.108 ;
  LAYER M3 ;
        RECT 20.544 9.056 20.576 9.088 ;
  LAYER M1 ;
        RECT 20.48 6.6 20.512 9.108 ;
  LAYER M3 ;
        RECT 20.48 6.62 20.512 6.652 ;
  LAYER M1 ;
        RECT 20.416 6.6 20.448 9.108 ;
  LAYER M3 ;
        RECT 20.416 9.056 20.448 9.088 ;
  LAYER M1 ;
        RECT 20.352 6.6 20.384 9.108 ;
  LAYER M3 ;
        RECT 20.352 6.62 20.384 6.652 ;
  LAYER M1 ;
        RECT 20.288 6.6 20.32 9.108 ;
  LAYER M3 ;
        RECT 20.288 9.056 20.32 9.088 ;
  LAYER M1 ;
        RECT 20.224 6.6 20.256 9.108 ;
  LAYER M3 ;
        RECT 20.224 6.62 20.256 6.652 ;
  LAYER M1 ;
        RECT 20.16 6.6 20.192 9.108 ;
  LAYER M3 ;
        RECT 20.16 9.056 20.192 9.088 ;
  LAYER M1 ;
        RECT 20.096 6.6 20.128 9.108 ;
  LAYER M3 ;
        RECT 20.096 6.62 20.128 6.652 ;
  LAYER M1 ;
        RECT 20.032 6.6 20.064 9.108 ;
  LAYER M3 ;
        RECT 20.032 9.056 20.064 9.088 ;
  LAYER M1 ;
        RECT 19.968 6.6 20 9.108 ;
  LAYER M3 ;
        RECT 19.968 6.62 20 6.652 ;
  LAYER M1 ;
        RECT 19.904 6.6 19.936 9.108 ;
  LAYER M3 ;
        RECT 19.904 9.056 19.936 9.088 ;
  LAYER M1 ;
        RECT 19.84 6.6 19.872 9.108 ;
  LAYER M3 ;
        RECT 19.84 6.62 19.872 6.652 ;
  LAYER M1 ;
        RECT 19.776 6.6 19.808 9.108 ;
  LAYER M3 ;
        RECT 19.776 9.056 19.808 9.088 ;
  LAYER M1 ;
        RECT 19.712 6.6 19.744 9.108 ;
  LAYER M3 ;
        RECT 19.712 6.62 19.744 6.652 ;
  LAYER M1 ;
        RECT 19.648 6.6 19.68 9.108 ;
  LAYER M3 ;
        RECT 19.648 9.056 19.68 9.088 ;
  LAYER M1 ;
        RECT 19.584 6.6 19.616 9.108 ;
  LAYER M3 ;
        RECT 21.952 6.684 21.984 6.716 ;
  LAYER M2 ;
        RECT 19.584 6.748 19.616 6.78 ;
  LAYER M2 ;
        RECT 21.952 6.812 21.984 6.844 ;
  LAYER M2 ;
        RECT 19.584 6.876 19.616 6.908 ;
  LAYER M2 ;
        RECT 21.952 6.94 21.984 6.972 ;
  LAYER M2 ;
        RECT 19.584 7.004 19.616 7.036 ;
  LAYER M2 ;
        RECT 21.952 7.068 21.984 7.1 ;
  LAYER M2 ;
        RECT 19.584 7.132 19.616 7.164 ;
  LAYER M2 ;
        RECT 21.952 7.196 21.984 7.228 ;
  LAYER M2 ;
        RECT 19.584 7.26 19.616 7.292 ;
  LAYER M2 ;
        RECT 21.952 7.324 21.984 7.356 ;
  LAYER M2 ;
        RECT 19.584 7.388 19.616 7.42 ;
  LAYER M2 ;
        RECT 21.952 7.452 21.984 7.484 ;
  LAYER M2 ;
        RECT 19.584 7.516 19.616 7.548 ;
  LAYER M2 ;
        RECT 21.952 7.58 21.984 7.612 ;
  LAYER M2 ;
        RECT 19.584 7.644 19.616 7.676 ;
  LAYER M2 ;
        RECT 21.952 7.708 21.984 7.74 ;
  LAYER M2 ;
        RECT 19.584 7.772 19.616 7.804 ;
  LAYER M2 ;
        RECT 21.952 7.836 21.984 7.868 ;
  LAYER M2 ;
        RECT 19.584 7.9 19.616 7.932 ;
  LAYER M2 ;
        RECT 21.952 7.964 21.984 7.996 ;
  LAYER M2 ;
        RECT 19.584 8.028 19.616 8.06 ;
  LAYER M2 ;
        RECT 21.952 8.092 21.984 8.124 ;
  LAYER M2 ;
        RECT 19.584 8.156 19.616 8.188 ;
  LAYER M2 ;
        RECT 21.952 8.22 21.984 8.252 ;
  LAYER M2 ;
        RECT 19.584 8.284 19.616 8.316 ;
  LAYER M2 ;
        RECT 21.952 8.348 21.984 8.38 ;
  LAYER M2 ;
        RECT 19.584 8.412 19.616 8.444 ;
  LAYER M2 ;
        RECT 21.952 8.476 21.984 8.508 ;
  LAYER M2 ;
        RECT 19.584 8.54 19.616 8.572 ;
  LAYER M2 ;
        RECT 21.952 8.604 21.984 8.636 ;
  LAYER M2 ;
        RECT 19.584 8.668 19.616 8.7 ;
  LAYER M2 ;
        RECT 21.952 8.732 21.984 8.764 ;
  LAYER M2 ;
        RECT 19.584 8.796 19.616 8.828 ;
  LAYER M2 ;
        RECT 21.952 8.86 21.984 8.892 ;
  LAYER M2 ;
        RECT 19.584 8.924 19.616 8.956 ;
  LAYER M2 ;
        RECT 19.536 6.552 22.032 9.156 ;
  LAYER M1 ;
        RECT 21.952 9.708 21.984 12.216 ;
  LAYER M3 ;
        RECT 21.952 12.164 21.984 12.196 ;
  LAYER M1 ;
        RECT 21.888 9.708 21.92 12.216 ;
  LAYER M3 ;
        RECT 21.888 9.728 21.92 9.76 ;
  LAYER M1 ;
        RECT 21.824 9.708 21.856 12.216 ;
  LAYER M3 ;
        RECT 21.824 12.164 21.856 12.196 ;
  LAYER M1 ;
        RECT 21.76 9.708 21.792 12.216 ;
  LAYER M3 ;
        RECT 21.76 9.728 21.792 9.76 ;
  LAYER M1 ;
        RECT 21.696 9.708 21.728 12.216 ;
  LAYER M3 ;
        RECT 21.696 12.164 21.728 12.196 ;
  LAYER M1 ;
        RECT 21.632 9.708 21.664 12.216 ;
  LAYER M3 ;
        RECT 21.632 9.728 21.664 9.76 ;
  LAYER M1 ;
        RECT 21.568 9.708 21.6 12.216 ;
  LAYER M3 ;
        RECT 21.568 12.164 21.6 12.196 ;
  LAYER M1 ;
        RECT 21.504 9.708 21.536 12.216 ;
  LAYER M3 ;
        RECT 21.504 9.728 21.536 9.76 ;
  LAYER M1 ;
        RECT 21.44 9.708 21.472 12.216 ;
  LAYER M3 ;
        RECT 21.44 12.164 21.472 12.196 ;
  LAYER M1 ;
        RECT 21.376 9.708 21.408 12.216 ;
  LAYER M3 ;
        RECT 21.376 9.728 21.408 9.76 ;
  LAYER M1 ;
        RECT 21.312 9.708 21.344 12.216 ;
  LAYER M3 ;
        RECT 21.312 12.164 21.344 12.196 ;
  LAYER M1 ;
        RECT 21.248 9.708 21.28 12.216 ;
  LAYER M3 ;
        RECT 21.248 9.728 21.28 9.76 ;
  LAYER M1 ;
        RECT 21.184 9.708 21.216 12.216 ;
  LAYER M3 ;
        RECT 21.184 12.164 21.216 12.196 ;
  LAYER M1 ;
        RECT 21.12 9.708 21.152 12.216 ;
  LAYER M3 ;
        RECT 21.12 9.728 21.152 9.76 ;
  LAYER M1 ;
        RECT 21.056 9.708 21.088 12.216 ;
  LAYER M3 ;
        RECT 21.056 12.164 21.088 12.196 ;
  LAYER M1 ;
        RECT 20.992 9.708 21.024 12.216 ;
  LAYER M3 ;
        RECT 20.992 9.728 21.024 9.76 ;
  LAYER M1 ;
        RECT 20.928 9.708 20.96 12.216 ;
  LAYER M3 ;
        RECT 20.928 12.164 20.96 12.196 ;
  LAYER M1 ;
        RECT 20.864 9.708 20.896 12.216 ;
  LAYER M3 ;
        RECT 20.864 9.728 20.896 9.76 ;
  LAYER M1 ;
        RECT 20.8 9.708 20.832 12.216 ;
  LAYER M3 ;
        RECT 20.8 12.164 20.832 12.196 ;
  LAYER M1 ;
        RECT 20.736 9.708 20.768 12.216 ;
  LAYER M3 ;
        RECT 20.736 9.728 20.768 9.76 ;
  LAYER M1 ;
        RECT 20.672 9.708 20.704 12.216 ;
  LAYER M3 ;
        RECT 20.672 12.164 20.704 12.196 ;
  LAYER M1 ;
        RECT 20.608 9.708 20.64 12.216 ;
  LAYER M3 ;
        RECT 20.608 9.728 20.64 9.76 ;
  LAYER M1 ;
        RECT 20.544 9.708 20.576 12.216 ;
  LAYER M3 ;
        RECT 20.544 12.164 20.576 12.196 ;
  LAYER M1 ;
        RECT 20.48 9.708 20.512 12.216 ;
  LAYER M3 ;
        RECT 20.48 9.728 20.512 9.76 ;
  LAYER M1 ;
        RECT 20.416 9.708 20.448 12.216 ;
  LAYER M3 ;
        RECT 20.416 12.164 20.448 12.196 ;
  LAYER M1 ;
        RECT 20.352 9.708 20.384 12.216 ;
  LAYER M3 ;
        RECT 20.352 9.728 20.384 9.76 ;
  LAYER M1 ;
        RECT 20.288 9.708 20.32 12.216 ;
  LAYER M3 ;
        RECT 20.288 12.164 20.32 12.196 ;
  LAYER M1 ;
        RECT 20.224 9.708 20.256 12.216 ;
  LAYER M3 ;
        RECT 20.224 9.728 20.256 9.76 ;
  LAYER M1 ;
        RECT 20.16 9.708 20.192 12.216 ;
  LAYER M3 ;
        RECT 20.16 12.164 20.192 12.196 ;
  LAYER M1 ;
        RECT 20.096 9.708 20.128 12.216 ;
  LAYER M3 ;
        RECT 20.096 9.728 20.128 9.76 ;
  LAYER M1 ;
        RECT 20.032 9.708 20.064 12.216 ;
  LAYER M3 ;
        RECT 20.032 12.164 20.064 12.196 ;
  LAYER M1 ;
        RECT 19.968 9.708 20 12.216 ;
  LAYER M3 ;
        RECT 19.968 9.728 20 9.76 ;
  LAYER M1 ;
        RECT 19.904 9.708 19.936 12.216 ;
  LAYER M3 ;
        RECT 19.904 12.164 19.936 12.196 ;
  LAYER M1 ;
        RECT 19.84 9.708 19.872 12.216 ;
  LAYER M3 ;
        RECT 19.84 9.728 19.872 9.76 ;
  LAYER M1 ;
        RECT 19.776 9.708 19.808 12.216 ;
  LAYER M3 ;
        RECT 19.776 12.164 19.808 12.196 ;
  LAYER M1 ;
        RECT 19.712 9.708 19.744 12.216 ;
  LAYER M3 ;
        RECT 19.712 9.728 19.744 9.76 ;
  LAYER M1 ;
        RECT 19.648 9.708 19.68 12.216 ;
  LAYER M3 ;
        RECT 19.648 12.164 19.68 12.196 ;
  LAYER M1 ;
        RECT 19.584 9.708 19.616 12.216 ;
  LAYER M3 ;
        RECT 21.952 9.792 21.984 9.824 ;
  LAYER M2 ;
        RECT 19.584 9.856 19.616 9.888 ;
  LAYER M2 ;
        RECT 21.952 9.92 21.984 9.952 ;
  LAYER M2 ;
        RECT 19.584 9.984 19.616 10.016 ;
  LAYER M2 ;
        RECT 21.952 10.048 21.984 10.08 ;
  LAYER M2 ;
        RECT 19.584 10.112 19.616 10.144 ;
  LAYER M2 ;
        RECT 21.952 10.176 21.984 10.208 ;
  LAYER M2 ;
        RECT 19.584 10.24 19.616 10.272 ;
  LAYER M2 ;
        RECT 21.952 10.304 21.984 10.336 ;
  LAYER M2 ;
        RECT 19.584 10.368 19.616 10.4 ;
  LAYER M2 ;
        RECT 21.952 10.432 21.984 10.464 ;
  LAYER M2 ;
        RECT 19.584 10.496 19.616 10.528 ;
  LAYER M2 ;
        RECT 21.952 10.56 21.984 10.592 ;
  LAYER M2 ;
        RECT 19.584 10.624 19.616 10.656 ;
  LAYER M2 ;
        RECT 21.952 10.688 21.984 10.72 ;
  LAYER M2 ;
        RECT 19.584 10.752 19.616 10.784 ;
  LAYER M2 ;
        RECT 21.952 10.816 21.984 10.848 ;
  LAYER M2 ;
        RECT 19.584 10.88 19.616 10.912 ;
  LAYER M2 ;
        RECT 21.952 10.944 21.984 10.976 ;
  LAYER M2 ;
        RECT 19.584 11.008 19.616 11.04 ;
  LAYER M2 ;
        RECT 21.952 11.072 21.984 11.104 ;
  LAYER M2 ;
        RECT 19.584 11.136 19.616 11.168 ;
  LAYER M2 ;
        RECT 21.952 11.2 21.984 11.232 ;
  LAYER M2 ;
        RECT 19.584 11.264 19.616 11.296 ;
  LAYER M2 ;
        RECT 21.952 11.328 21.984 11.36 ;
  LAYER M2 ;
        RECT 19.584 11.392 19.616 11.424 ;
  LAYER M2 ;
        RECT 21.952 11.456 21.984 11.488 ;
  LAYER M2 ;
        RECT 19.584 11.52 19.616 11.552 ;
  LAYER M2 ;
        RECT 21.952 11.584 21.984 11.616 ;
  LAYER M2 ;
        RECT 19.584 11.648 19.616 11.68 ;
  LAYER M2 ;
        RECT 21.952 11.712 21.984 11.744 ;
  LAYER M2 ;
        RECT 19.584 11.776 19.616 11.808 ;
  LAYER M2 ;
        RECT 21.952 11.84 21.984 11.872 ;
  LAYER M2 ;
        RECT 19.584 11.904 19.616 11.936 ;
  LAYER M2 ;
        RECT 21.952 11.968 21.984 12 ;
  LAYER M2 ;
        RECT 19.584 12.032 19.616 12.064 ;
  LAYER M2 ;
        RECT 19.536 9.66 22.032 12.264 ;
  LAYER M1 ;
        RECT 21.952 12.816 21.984 15.324 ;
  LAYER M3 ;
        RECT 21.952 15.272 21.984 15.304 ;
  LAYER M1 ;
        RECT 21.888 12.816 21.92 15.324 ;
  LAYER M3 ;
        RECT 21.888 12.836 21.92 12.868 ;
  LAYER M1 ;
        RECT 21.824 12.816 21.856 15.324 ;
  LAYER M3 ;
        RECT 21.824 15.272 21.856 15.304 ;
  LAYER M1 ;
        RECT 21.76 12.816 21.792 15.324 ;
  LAYER M3 ;
        RECT 21.76 12.836 21.792 12.868 ;
  LAYER M1 ;
        RECT 21.696 12.816 21.728 15.324 ;
  LAYER M3 ;
        RECT 21.696 15.272 21.728 15.304 ;
  LAYER M1 ;
        RECT 21.632 12.816 21.664 15.324 ;
  LAYER M3 ;
        RECT 21.632 12.836 21.664 12.868 ;
  LAYER M1 ;
        RECT 21.568 12.816 21.6 15.324 ;
  LAYER M3 ;
        RECT 21.568 15.272 21.6 15.304 ;
  LAYER M1 ;
        RECT 21.504 12.816 21.536 15.324 ;
  LAYER M3 ;
        RECT 21.504 12.836 21.536 12.868 ;
  LAYER M1 ;
        RECT 21.44 12.816 21.472 15.324 ;
  LAYER M3 ;
        RECT 21.44 15.272 21.472 15.304 ;
  LAYER M1 ;
        RECT 21.376 12.816 21.408 15.324 ;
  LAYER M3 ;
        RECT 21.376 12.836 21.408 12.868 ;
  LAYER M1 ;
        RECT 21.312 12.816 21.344 15.324 ;
  LAYER M3 ;
        RECT 21.312 15.272 21.344 15.304 ;
  LAYER M1 ;
        RECT 21.248 12.816 21.28 15.324 ;
  LAYER M3 ;
        RECT 21.248 12.836 21.28 12.868 ;
  LAYER M1 ;
        RECT 21.184 12.816 21.216 15.324 ;
  LAYER M3 ;
        RECT 21.184 15.272 21.216 15.304 ;
  LAYER M1 ;
        RECT 21.12 12.816 21.152 15.324 ;
  LAYER M3 ;
        RECT 21.12 12.836 21.152 12.868 ;
  LAYER M1 ;
        RECT 21.056 12.816 21.088 15.324 ;
  LAYER M3 ;
        RECT 21.056 15.272 21.088 15.304 ;
  LAYER M1 ;
        RECT 20.992 12.816 21.024 15.324 ;
  LAYER M3 ;
        RECT 20.992 12.836 21.024 12.868 ;
  LAYER M1 ;
        RECT 20.928 12.816 20.96 15.324 ;
  LAYER M3 ;
        RECT 20.928 15.272 20.96 15.304 ;
  LAYER M1 ;
        RECT 20.864 12.816 20.896 15.324 ;
  LAYER M3 ;
        RECT 20.864 12.836 20.896 12.868 ;
  LAYER M1 ;
        RECT 20.8 12.816 20.832 15.324 ;
  LAYER M3 ;
        RECT 20.8 15.272 20.832 15.304 ;
  LAYER M1 ;
        RECT 20.736 12.816 20.768 15.324 ;
  LAYER M3 ;
        RECT 20.736 12.836 20.768 12.868 ;
  LAYER M1 ;
        RECT 20.672 12.816 20.704 15.324 ;
  LAYER M3 ;
        RECT 20.672 15.272 20.704 15.304 ;
  LAYER M1 ;
        RECT 20.608 12.816 20.64 15.324 ;
  LAYER M3 ;
        RECT 20.608 12.836 20.64 12.868 ;
  LAYER M1 ;
        RECT 20.544 12.816 20.576 15.324 ;
  LAYER M3 ;
        RECT 20.544 15.272 20.576 15.304 ;
  LAYER M1 ;
        RECT 20.48 12.816 20.512 15.324 ;
  LAYER M3 ;
        RECT 20.48 12.836 20.512 12.868 ;
  LAYER M1 ;
        RECT 20.416 12.816 20.448 15.324 ;
  LAYER M3 ;
        RECT 20.416 15.272 20.448 15.304 ;
  LAYER M1 ;
        RECT 20.352 12.816 20.384 15.324 ;
  LAYER M3 ;
        RECT 20.352 12.836 20.384 12.868 ;
  LAYER M1 ;
        RECT 20.288 12.816 20.32 15.324 ;
  LAYER M3 ;
        RECT 20.288 15.272 20.32 15.304 ;
  LAYER M1 ;
        RECT 20.224 12.816 20.256 15.324 ;
  LAYER M3 ;
        RECT 20.224 12.836 20.256 12.868 ;
  LAYER M1 ;
        RECT 20.16 12.816 20.192 15.324 ;
  LAYER M3 ;
        RECT 20.16 15.272 20.192 15.304 ;
  LAYER M1 ;
        RECT 20.096 12.816 20.128 15.324 ;
  LAYER M3 ;
        RECT 20.096 12.836 20.128 12.868 ;
  LAYER M1 ;
        RECT 20.032 12.816 20.064 15.324 ;
  LAYER M3 ;
        RECT 20.032 15.272 20.064 15.304 ;
  LAYER M1 ;
        RECT 19.968 12.816 20 15.324 ;
  LAYER M3 ;
        RECT 19.968 12.836 20 12.868 ;
  LAYER M1 ;
        RECT 19.904 12.816 19.936 15.324 ;
  LAYER M3 ;
        RECT 19.904 15.272 19.936 15.304 ;
  LAYER M1 ;
        RECT 19.84 12.816 19.872 15.324 ;
  LAYER M3 ;
        RECT 19.84 12.836 19.872 12.868 ;
  LAYER M1 ;
        RECT 19.776 12.816 19.808 15.324 ;
  LAYER M3 ;
        RECT 19.776 15.272 19.808 15.304 ;
  LAYER M1 ;
        RECT 19.712 12.816 19.744 15.324 ;
  LAYER M3 ;
        RECT 19.712 12.836 19.744 12.868 ;
  LAYER M1 ;
        RECT 19.648 12.816 19.68 15.324 ;
  LAYER M3 ;
        RECT 19.648 15.272 19.68 15.304 ;
  LAYER M1 ;
        RECT 19.584 12.816 19.616 15.324 ;
  LAYER M3 ;
        RECT 21.952 12.9 21.984 12.932 ;
  LAYER M2 ;
        RECT 19.584 12.964 19.616 12.996 ;
  LAYER M2 ;
        RECT 21.952 13.028 21.984 13.06 ;
  LAYER M2 ;
        RECT 19.584 13.092 19.616 13.124 ;
  LAYER M2 ;
        RECT 21.952 13.156 21.984 13.188 ;
  LAYER M2 ;
        RECT 19.584 13.22 19.616 13.252 ;
  LAYER M2 ;
        RECT 21.952 13.284 21.984 13.316 ;
  LAYER M2 ;
        RECT 19.584 13.348 19.616 13.38 ;
  LAYER M2 ;
        RECT 21.952 13.412 21.984 13.444 ;
  LAYER M2 ;
        RECT 19.584 13.476 19.616 13.508 ;
  LAYER M2 ;
        RECT 21.952 13.54 21.984 13.572 ;
  LAYER M2 ;
        RECT 19.584 13.604 19.616 13.636 ;
  LAYER M2 ;
        RECT 21.952 13.668 21.984 13.7 ;
  LAYER M2 ;
        RECT 19.584 13.732 19.616 13.764 ;
  LAYER M2 ;
        RECT 21.952 13.796 21.984 13.828 ;
  LAYER M2 ;
        RECT 19.584 13.86 19.616 13.892 ;
  LAYER M2 ;
        RECT 21.952 13.924 21.984 13.956 ;
  LAYER M2 ;
        RECT 19.584 13.988 19.616 14.02 ;
  LAYER M2 ;
        RECT 21.952 14.052 21.984 14.084 ;
  LAYER M2 ;
        RECT 19.584 14.116 19.616 14.148 ;
  LAYER M2 ;
        RECT 21.952 14.18 21.984 14.212 ;
  LAYER M2 ;
        RECT 19.584 14.244 19.616 14.276 ;
  LAYER M2 ;
        RECT 21.952 14.308 21.984 14.34 ;
  LAYER M2 ;
        RECT 19.584 14.372 19.616 14.404 ;
  LAYER M2 ;
        RECT 21.952 14.436 21.984 14.468 ;
  LAYER M2 ;
        RECT 19.584 14.5 19.616 14.532 ;
  LAYER M2 ;
        RECT 21.952 14.564 21.984 14.596 ;
  LAYER M2 ;
        RECT 19.584 14.628 19.616 14.66 ;
  LAYER M2 ;
        RECT 21.952 14.692 21.984 14.724 ;
  LAYER M2 ;
        RECT 19.584 14.756 19.616 14.788 ;
  LAYER M2 ;
        RECT 21.952 14.82 21.984 14.852 ;
  LAYER M2 ;
        RECT 19.584 14.884 19.616 14.916 ;
  LAYER M2 ;
        RECT 21.952 14.948 21.984 14.98 ;
  LAYER M2 ;
        RECT 19.584 15.012 19.616 15.044 ;
  LAYER M2 ;
        RECT 21.952 15.076 21.984 15.108 ;
  LAYER M2 ;
        RECT 19.584 15.14 19.616 15.172 ;
  LAYER M2 ;
        RECT 19.536 12.768 22.032 15.372 ;
  LAYER M1 ;
        RECT 21.952 15.924 21.984 18.432 ;
  LAYER M3 ;
        RECT 21.952 18.38 21.984 18.412 ;
  LAYER M1 ;
        RECT 21.888 15.924 21.92 18.432 ;
  LAYER M3 ;
        RECT 21.888 15.944 21.92 15.976 ;
  LAYER M1 ;
        RECT 21.824 15.924 21.856 18.432 ;
  LAYER M3 ;
        RECT 21.824 18.38 21.856 18.412 ;
  LAYER M1 ;
        RECT 21.76 15.924 21.792 18.432 ;
  LAYER M3 ;
        RECT 21.76 15.944 21.792 15.976 ;
  LAYER M1 ;
        RECT 21.696 15.924 21.728 18.432 ;
  LAYER M3 ;
        RECT 21.696 18.38 21.728 18.412 ;
  LAYER M1 ;
        RECT 21.632 15.924 21.664 18.432 ;
  LAYER M3 ;
        RECT 21.632 15.944 21.664 15.976 ;
  LAYER M1 ;
        RECT 21.568 15.924 21.6 18.432 ;
  LAYER M3 ;
        RECT 21.568 18.38 21.6 18.412 ;
  LAYER M1 ;
        RECT 21.504 15.924 21.536 18.432 ;
  LAYER M3 ;
        RECT 21.504 15.944 21.536 15.976 ;
  LAYER M1 ;
        RECT 21.44 15.924 21.472 18.432 ;
  LAYER M3 ;
        RECT 21.44 18.38 21.472 18.412 ;
  LAYER M1 ;
        RECT 21.376 15.924 21.408 18.432 ;
  LAYER M3 ;
        RECT 21.376 15.944 21.408 15.976 ;
  LAYER M1 ;
        RECT 21.312 15.924 21.344 18.432 ;
  LAYER M3 ;
        RECT 21.312 18.38 21.344 18.412 ;
  LAYER M1 ;
        RECT 21.248 15.924 21.28 18.432 ;
  LAYER M3 ;
        RECT 21.248 15.944 21.28 15.976 ;
  LAYER M1 ;
        RECT 21.184 15.924 21.216 18.432 ;
  LAYER M3 ;
        RECT 21.184 18.38 21.216 18.412 ;
  LAYER M1 ;
        RECT 21.12 15.924 21.152 18.432 ;
  LAYER M3 ;
        RECT 21.12 15.944 21.152 15.976 ;
  LAYER M1 ;
        RECT 21.056 15.924 21.088 18.432 ;
  LAYER M3 ;
        RECT 21.056 18.38 21.088 18.412 ;
  LAYER M1 ;
        RECT 20.992 15.924 21.024 18.432 ;
  LAYER M3 ;
        RECT 20.992 15.944 21.024 15.976 ;
  LAYER M1 ;
        RECT 20.928 15.924 20.96 18.432 ;
  LAYER M3 ;
        RECT 20.928 18.38 20.96 18.412 ;
  LAYER M1 ;
        RECT 20.864 15.924 20.896 18.432 ;
  LAYER M3 ;
        RECT 20.864 15.944 20.896 15.976 ;
  LAYER M1 ;
        RECT 20.8 15.924 20.832 18.432 ;
  LAYER M3 ;
        RECT 20.8 18.38 20.832 18.412 ;
  LAYER M1 ;
        RECT 20.736 15.924 20.768 18.432 ;
  LAYER M3 ;
        RECT 20.736 15.944 20.768 15.976 ;
  LAYER M1 ;
        RECT 20.672 15.924 20.704 18.432 ;
  LAYER M3 ;
        RECT 20.672 18.38 20.704 18.412 ;
  LAYER M1 ;
        RECT 20.608 15.924 20.64 18.432 ;
  LAYER M3 ;
        RECT 20.608 15.944 20.64 15.976 ;
  LAYER M1 ;
        RECT 20.544 15.924 20.576 18.432 ;
  LAYER M3 ;
        RECT 20.544 18.38 20.576 18.412 ;
  LAYER M1 ;
        RECT 20.48 15.924 20.512 18.432 ;
  LAYER M3 ;
        RECT 20.48 15.944 20.512 15.976 ;
  LAYER M1 ;
        RECT 20.416 15.924 20.448 18.432 ;
  LAYER M3 ;
        RECT 20.416 18.38 20.448 18.412 ;
  LAYER M1 ;
        RECT 20.352 15.924 20.384 18.432 ;
  LAYER M3 ;
        RECT 20.352 15.944 20.384 15.976 ;
  LAYER M1 ;
        RECT 20.288 15.924 20.32 18.432 ;
  LAYER M3 ;
        RECT 20.288 18.38 20.32 18.412 ;
  LAYER M1 ;
        RECT 20.224 15.924 20.256 18.432 ;
  LAYER M3 ;
        RECT 20.224 15.944 20.256 15.976 ;
  LAYER M1 ;
        RECT 20.16 15.924 20.192 18.432 ;
  LAYER M3 ;
        RECT 20.16 18.38 20.192 18.412 ;
  LAYER M1 ;
        RECT 20.096 15.924 20.128 18.432 ;
  LAYER M3 ;
        RECT 20.096 15.944 20.128 15.976 ;
  LAYER M1 ;
        RECT 20.032 15.924 20.064 18.432 ;
  LAYER M3 ;
        RECT 20.032 18.38 20.064 18.412 ;
  LAYER M1 ;
        RECT 19.968 15.924 20 18.432 ;
  LAYER M3 ;
        RECT 19.968 15.944 20 15.976 ;
  LAYER M1 ;
        RECT 19.904 15.924 19.936 18.432 ;
  LAYER M3 ;
        RECT 19.904 18.38 19.936 18.412 ;
  LAYER M1 ;
        RECT 19.84 15.924 19.872 18.432 ;
  LAYER M3 ;
        RECT 19.84 15.944 19.872 15.976 ;
  LAYER M1 ;
        RECT 19.776 15.924 19.808 18.432 ;
  LAYER M3 ;
        RECT 19.776 18.38 19.808 18.412 ;
  LAYER M1 ;
        RECT 19.712 15.924 19.744 18.432 ;
  LAYER M3 ;
        RECT 19.712 15.944 19.744 15.976 ;
  LAYER M1 ;
        RECT 19.648 15.924 19.68 18.432 ;
  LAYER M3 ;
        RECT 19.648 18.38 19.68 18.412 ;
  LAYER M1 ;
        RECT 19.584 15.924 19.616 18.432 ;
  LAYER M3 ;
        RECT 21.952 16.008 21.984 16.04 ;
  LAYER M2 ;
        RECT 19.584 16.072 19.616 16.104 ;
  LAYER M2 ;
        RECT 21.952 16.136 21.984 16.168 ;
  LAYER M2 ;
        RECT 19.584 16.2 19.616 16.232 ;
  LAYER M2 ;
        RECT 21.952 16.264 21.984 16.296 ;
  LAYER M2 ;
        RECT 19.584 16.328 19.616 16.36 ;
  LAYER M2 ;
        RECT 21.952 16.392 21.984 16.424 ;
  LAYER M2 ;
        RECT 19.584 16.456 19.616 16.488 ;
  LAYER M2 ;
        RECT 21.952 16.52 21.984 16.552 ;
  LAYER M2 ;
        RECT 19.584 16.584 19.616 16.616 ;
  LAYER M2 ;
        RECT 21.952 16.648 21.984 16.68 ;
  LAYER M2 ;
        RECT 19.584 16.712 19.616 16.744 ;
  LAYER M2 ;
        RECT 21.952 16.776 21.984 16.808 ;
  LAYER M2 ;
        RECT 19.584 16.84 19.616 16.872 ;
  LAYER M2 ;
        RECT 21.952 16.904 21.984 16.936 ;
  LAYER M2 ;
        RECT 19.584 16.968 19.616 17 ;
  LAYER M2 ;
        RECT 21.952 17.032 21.984 17.064 ;
  LAYER M2 ;
        RECT 19.584 17.096 19.616 17.128 ;
  LAYER M2 ;
        RECT 21.952 17.16 21.984 17.192 ;
  LAYER M2 ;
        RECT 19.584 17.224 19.616 17.256 ;
  LAYER M2 ;
        RECT 21.952 17.288 21.984 17.32 ;
  LAYER M2 ;
        RECT 19.584 17.352 19.616 17.384 ;
  LAYER M2 ;
        RECT 21.952 17.416 21.984 17.448 ;
  LAYER M2 ;
        RECT 19.584 17.48 19.616 17.512 ;
  LAYER M2 ;
        RECT 21.952 17.544 21.984 17.576 ;
  LAYER M2 ;
        RECT 19.584 17.608 19.616 17.64 ;
  LAYER M2 ;
        RECT 21.952 17.672 21.984 17.704 ;
  LAYER M2 ;
        RECT 19.584 17.736 19.616 17.768 ;
  LAYER M2 ;
        RECT 21.952 17.8 21.984 17.832 ;
  LAYER M2 ;
        RECT 19.584 17.864 19.616 17.896 ;
  LAYER M2 ;
        RECT 21.952 17.928 21.984 17.96 ;
  LAYER M2 ;
        RECT 19.584 17.992 19.616 18.024 ;
  LAYER M2 ;
        RECT 21.952 18.056 21.984 18.088 ;
  LAYER M2 ;
        RECT 19.584 18.12 19.616 18.152 ;
  LAYER M2 ;
        RECT 21.952 18.184 21.984 18.216 ;
  LAYER M2 ;
        RECT 19.584 18.248 19.616 18.28 ;
  LAYER M2 ;
        RECT 19.536 15.876 22.032 18.48 ;
  LAYER M1 ;
        RECT 18.976 6.6 19.008 9.108 ;
  LAYER M3 ;
        RECT 18.976 9.056 19.008 9.088 ;
  LAYER M1 ;
        RECT 18.912 6.6 18.944 9.108 ;
  LAYER M3 ;
        RECT 18.912 6.62 18.944 6.652 ;
  LAYER M1 ;
        RECT 18.848 6.6 18.88 9.108 ;
  LAYER M3 ;
        RECT 18.848 9.056 18.88 9.088 ;
  LAYER M1 ;
        RECT 18.784 6.6 18.816 9.108 ;
  LAYER M3 ;
        RECT 18.784 6.62 18.816 6.652 ;
  LAYER M1 ;
        RECT 18.72 6.6 18.752 9.108 ;
  LAYER M3 ;
        RECT 18.72 9.056 18.752 9.088 ;
  LAYER M1 ;
        RECT 18.656 6.6 18.688 9.108 ;
  LAYER M3 ;
        RECT 18.656 6.62 18.688 6.652 ;
  LAYER M1 ;
        RECT 18.592 6.6 18.624 9.108 ;
  LAYER M3 ;
        RECT 18.592 9.056 18.624 9.088 ;
  LAYER M1 ;
        RECT 18.528 6.6 18.56 9.108 ;
  LAYER M3 ;
        RECT 18.528 6.62 18.56 6.652 ;
  LAYER M1 ;
        RECT 18.464 6.6 18.496 9.108 ;
  LAYER M3 ;
        RECT 18.464 9.056 18.496 9.088 ;
  LAYER M1 ;
        RECT 18.4 6.6 18.432 9.108 ;
  LAYER M3 ;
        RECT 18.4 6.62 18.432 6.652 ;
  LAYER M1 ;
        RECT 18.336 6.6 18.368 9.108 ;
  LAYER M3 ;
        RECT 18.336 9.056 18.368 9.088 ;
  LAYER M1 ;
        RECT 18.272 6.6 18.304 9.108 ;
  LAYER M3 ;
        RECT 18.272 6.62 18.304 6.652 ;
  LAYER M1 ;
        RECT 18.208 6.6 18.24 9.108 ;
  LAYER M3 ;
        RECT 18.208 9.056 18.24 9.088 ;
  LAYER M1 ;
        RECT 18.144 6.6 18.176 9.108 ;
  LAYER M3 ;
        RECT 18.144 6.62 18.176 6.652 ;
  LAYER M1 ;
        RECT 18.08 6.6 18.112 9.108 ;
  LAYER M3 ;
        RECT 18.08 9.056 18.112 9.088 ;
  LAYER M1 ;
        RECT 18.016 6.6 18.048 9.108 ;
  LAYER M3 ;
        RECT 18.016 6.62 18.048 6.652 ;
  LAYER M1 ;
        RECT 17.952 6.6 17.984 9.108 ;
  LAYER M3 ;
        RECT 17.952 9.056 17.984 9.088 ;
  LAYER M1 ;
        RECT 17.888 6.6 17.92 9.108 ;
  LAYER M3 ;
        RECT 17.888 6.62 17.92 6.652 ;
  LAYER M1 ;
        RECT 17.824 6.6 17.856 9.108 ;
  LAYER M3 ;
        RECT 17.824 9.056 17.856 9.088 ;
  LAYER M1 ;
        RECT 17.76 6.6 17.792 9.108 ;
  LAYER M3 ;
        RECT 17.76 6.62 17.792 6.652 ;
  LAYER M1 ;
        RECT 17.696 6.6 17.728 9.108 ;
  LAYER M3 ;
        RECT 17.696 9.056 17.728 9.088 ;
  LAYER M1 ;
        RECT 17.632 6.6 17.664 9.108 ;
  LAYER M3 ;
        RECT 17.632 6.62 17.664 6.652 ;
  LAYER M1 ;
        RECT 17.568 6.6 17.6 9.108 ;
  LAYER M3 ;
        RECT 17.568 9.056 17.6 9.088 ;
  LAYER M1 ;
        RECT 17.504 6.6 17.536 9.108 ;
  LAYER M3 ;
        RECT 17.504 6.62 17.536 6.652 ;
  LAYER M1 ;
        RECT 17.44 6.6 17.472 9.108 ;
  LAYER M3 ;
        RECT 17.44 9.056 17.472 9.088 ;
  LAYER M1 ;
        RECT 17.376 6.6 17.408 9.108 ;
  LAYER M3 ;
        RECT 17.376 6.62 17.408 6.652 ;
  LAYER M1 ;
        RECT 17.312 6.6 17.344 9.108 ;
  LAYER M3 ;
        RECT 17.312 9.056 17.344 9.088 ;
  LAYER M1 ;
        RECT 17.248 6.6 17.28 9.108 ;
  LAYER M3 ;
        RECT 17.248 6.62 17.28 6.652 ;
  LAYER M1 ;
        RECT 17.184 6.6 17.216 9.108 ;
  LAYER M3 ;
        RECT 17.184 9.056 17.216 9.088 ;
  LAYER M1 ;
        RECT 17.12 6.6 17.152 9.108 ;
  LAYER M3 ;
        RECT 17.12 6.62 17.152 6.652 ;
  LAYER M1 ;
        RECT 17.056 6.6 17.088 9.108 ;
  LAYER M3 ;
        RECT 17.056 9.056 17.088 9.088 ;
  LAYER M1 ;
        RECT 16.992 6.6 17.024 9.108 ;
  LAYER M3 ;
        RECT 16.992 6.62 17.024 6.652 ;
  LAYER M1 ;
        RECT 16.928 6.6 16.96 9.108 ;
  LAYER M3 ;
        RECT 16.928 9.056 16.96 9.088 ;
  LAYER M1 ;
        RECT 16.864 6.6 16.896 9.108 ;
  LAYER M3 ;
        RECT 16.864 6.62 16.896 6.652 ;
  LAYER M1 ;
        RECT 16.8 6.6 16.832 9.108 ;
  LAYER M3 ;
        RECT 16.8 9.056 16.832 9.088 ;
  LAYER M1 ;
        RECT 16.736 6.6 16.768 9.108 ;
  LAYER M3 ;
        RECT 16.736 6.62 16.768 6.652 ;
  LAYER M1 ;
        RECT 16.672 6.6 16.704 9.108 ;
  LAYER M3 ;
        RECT 16.672 9.056 16.704 9.088 ;
  LAYER M1 ;
        RECT 16.608 6.6 16.64 9.108 ;
  LAYER M3 ;
        RECT 18.976 6.684 19.008 6.716 ;
  LAYER M2 ;
        RECT 16.608 6.748 16.64 6.78 ;
  LAYER M2 ;
        RECT 18.976 6.812 19.008 6.844 ;
  LAYER M2 ;
        RECT 16.608 6.876 16.64 6.908 ;
  LAYER M2 ;
        RECT 18.976 6.94 19.008 6.972 ;
  LAYER M2 ;
        RECT 16.608 7.004 16.64 7.036 ;
  LAYER M2 ;
        RECT 18.976 7.068 19.008 7.1 ;
  LAYER M2 ;
        RECT 16.608 7.132 16.64 7.164 ;
  LAYER M2 ;
        RECT 18.976 7.196 19.008 7.228 ;
  LAYER M2 ;
        RECT 16.608 7.26 16.64 7.292 ;
  LAYER M2 ;
        RECT 18.976 7.324 19.008 7.356 ;
  LAYER M2 ;
        RECT 16.608 7.388 16.64 7.42 ;
  LAYER M2 ;
        RECT 18.976 7.452 19.008 7.484 ;
  LAYER M2 ;
        RECT 16.608 7.516 16.64 7.548 ;
  LAYER M2 ;
        RECT 18.976 7.58 19.008 7.612 ;
  LAYER M2 ;
        RECT 16.608 7.644 16.64 7.676 ;
  LAYER M2 ;
        RECT 18.976 7.708 19.008 7.74 ;
  LAYER M2 ;
        RECT 16.608 7.772 16.64 7.804 ;
  LAYER M2 ;
        RECT 18.976 7.836 19.008 7.868 ;
  LAYER M2 ;
        RECT 16.608 7.9 16.64 7.932 ;
  LAYER M2 ;
        RECT 18.976 7.964 19.008 7.996 ;
  LAYER M2 ;
        RECT 16.608 8.028 16.64 8.06 ;
  LAYER M2 ;
        RECT 18.976 8.092 19.008 8.124 ;
  LAYER M2 ;
        RECT 16.608 8.156 16.64 8.188 ;
  LAYER M2 ;
        RECT 18.976 8.22 19.008 8.252 ;
  LAYER M2 ;
        RECT 16.608 8.284 16.64 8.316 ;
  LAYER M2 ;
        RECT 18.976 8.348 19.008 8.38 ;
  LAYER M2 ;
        RECT 16.608 8.412 16.64 8.444 ;
  LAYER M2 ;
        RECT 18.976 8.476 19.008 8.508 ;
  LAYER M2 ;
        RECT 16.608 8.54 16.64 8.572 ;
  LAYER M2 ;
        RECT 18.976 8.604 19.008 8.636 ;
  LAYER M2 ;
        RECT 16.608 8.668 16.64 8.7 ;
  LAYER M2 ;
        RECT 18.976 8.732 19.008 8.764 ;
  LAYER M2 ;
        RECT 16.608 8.796 16.64 8.828 ;
  LAYER M2 ;
        RECT 18.976 8.86 19.008 8.892 ;
  LAYER M2 ;
        RECT 16.608 8.924 16.64 8.956 ;
  LAYER M2 ;
        RECT 16.56 6.552 19.056 9.156 ;
  LAYER M1 ;
        RECT 18.976 9.708 19.008 12.216 ;
  LAYER M3 ;
        RECT 18.976 12.164 19.008 12.196 ;
  LAYER M1 ;
        RECT 18.912 9.708 18.944 12.216 ;
  LAYER M3 ;
        RECT 18.912 9.728 18.944 9.76 ;
  LAYER M1 ;
        RECT 18.848 9.708 18.88 12.216 ;
  LAYER M3 ;
        RECT 18.848 12.164 18.88 12.196 ;
  LAYER M1 ;
        RECT 18.784 9.708 18.816 12.216 ;
  LAYER M3 ;
        RECT 18.784 9.728 18.816 9.76 ;
  LAYER M1 ;
        RECT 18.72 9.708 18.752 12.216 ;
  LAYER M3 ;
        RECT 18.72 12.164 18.752 12.196 ;
  LAYER M1 ;
        RECT 18.656 9.708 18.688 12.216 ;
  LAYER M3 ;
        RECT 18.656 9.728 18.688 9.76 ;
  LAYER M1 ;
        RECT 18.592 9.708 18.624 12.216 ;
  LAYER M3 ;
        RECT 18.592 12.164 18.624 12.196 ;
  LAYER M1 ;
        RECT 18.528 9.708 18.56 12.216 ;
  LAYER M3 ;
        RECT 18.528 9.728 18.56 9.76 ;
  LAYER M1 ;
        RECT 18.464 9.708 18.496 12.216 ;
  LAYER M3 ;
        RECT 18.464 12.164 18.496 12.196 ;
  LAYER M1 ;
        RECT 18.4 9.708 18.432 12.216 ;
  LAYER M3 ;
        RECT 18.4 9.728 18.432 9.76 ;
  LAYER M1 ;
        RECT 18.336 9.708 18.368 12.216 ;
  LAYER M3 ;
        RECT 18.336 12.164 18.368 12.196 ;
  LAYER M1 ;
        RECT 18.272 9.708 18.304 12.216 ;
  LAYER M3 ;
        RECT 18.272 9.728 18.304 9.76 ;
  LAYER M1 ;
        RECT 18.208 9.708 18.24 12.216 ;
  LAYER M3 ;
        RECT 18.208 12.164 18.24 12.196 ;
  LAYER M1 ;
        RECT 18.144 9.708 18.176 12.216 ;
  LAYER M3 ;
        RECT 18.144 9.728 18.176 9.76 ;
  LAYER M1 ;
        RECT 18.08 9.708 18.112 12.216 ;
  LAYER M3 ;
        RECT 18.08 12.164 18.112 12.196 ;
  LAYER M1 ;
        RECT 18.016 9.708 18.048 12.216 ;
  LAYER M3 ;
        RECT 18.016 9.728 18.048 9.76 ;
  LAYER M1 ;
        RECT 17.952 9.708 17.984 12.216 ;
  LAYER M3 ;
        RECT 17.952 12.164 17.984 12.196 ;
  LAYER M1 ;
        RECT 17.888 9.708 17.92 12.216 ;
  LAYER M3 ;
        RECT 17.888 9.728 17.92 9.76 ;
  LAYER M1 ;
        RECT 17.824 9.708 17.856 12.216 ;
  LAYER M3 ;
        RECT 17.824 12.164 17.856 12.196 ;
  LAYER M1 ;
        RECT 17.76 9.708 17.792 12.216 ;
  LAYER M3 ;
        RECT 17.76 9.728 17.792 9.76 ;
  LAYER M1 ;
        RECT 17.696 9.708 17.728 12.216 ;
  LAYER M3 ;
        RECT 17.696 12.164 17.728 12.196 ;
  LAYER M1 ;
        RECT 17.632 9.708 17.664 12.216 ;
  LAYER M3 ;
        RECT 17.632 9.728 17.664 9.76 ;
  LAYER M1 ;
        RECT 17.568 9.708 17.6 12.216 ;
  LAYER M3 ;
        RECT 17.568 12.164 17.6 12.196 ;
  LAYER M1 ;
        RECT 17.504 9.708 17.536 12.216 ;
  LAYER M3 ;
        RECT 17.504 9.728 17.536 9.76 ;
  LAYER M1 ;
        RECT 17.44 9.708 17.472 12.216 ;
  LAYER M3 ;
        RECT 17.44 12.164 17.472 12.196 ;
  LAYER M1 ;
        RECT 17.376 9.708 17.408 12.216 ;
  LAYER M3 ;
        RECT 17.376 9.728 17.408 9.76 ;
  LAYER M1 ;
        RECT 17.312 9.708 17.344 12.216 ;
  LAYER M3 ;
        RECT 17.312 12.164 17.344 12.196 ;
  LAYER M1 ;
        RECT 17.248 9.708 17.28 12.216 ;
  LAYER M3 ;
        RECT 17.248 9.728 17.28 9.76 ;
  LAYER M1 ;
        RECT 17.184 9.708 17.216 12.216 ;
  LAYER M3 ;
        RECT 17.184 12.164 17.216 12.196 ;
  LAYER M1 ;
        RECT 17.12 9.708 17.152 12.216 ;
  LAYER M3 ;
        RECT 17.12 9.728 17.152 9.76 ;
  LAYER M1 ;
        RECT 17.056 9.708 17.088 12.216 ;
  LAYER M3 ;
        RECT 17.056 12.164 17.088 12.196 ;
  LAYER M1 ;
        RECT 16.992 9.708 17.024 12.216 ;
  LAYER M3 ;
        RECT 16.992 9.728 17.024 9.76 ;
  LAYER M1 ;
        RECT 16.928 9.708 16.96 12.216 ;
  LAYER M3 ;
        RECT 16.928 12.164 16.96 12.196 ;
  LAYER M1 ;
        RECT 16.864 9.708 16.896 12.216 ;
  LAYER M3 ;
        RECT 16.864 9.728 16.896 9.76 ;
  LAYER M1 ;
        RECT 16.8 9.708 16.832 12.216 ;
  LAYER M3 ;
        RECT 16.8 12.164 16.832 12.196 ;
  LAYER M1 ;
        RECT 16.736 9.708 16.768 12.216 ;
  LAYER M3 ;
        RECT 16.736 9.728 16.768 9.76 ;
  LAYER M1 ;
        RECT 16.672 9.708 16.704 12.216 ;
  LAYER M3 ;
        RECT 16.672 12.164 16.704 12.196 ;
  LAYER M1 ;
        RECT 16.608 9.708 16.64 12.216 ;
  LAYER M3 ;
        RECT 18.976 9.792 19.008 9.824 ;
  LAYER M2 ;
        RECT 16.608 9.856 16.64 9.888 ;
  LAYER M2 ;
        RECT 18.976 9.92 19.008 9.952 ;
  LAYER M2 ;
        RECT 16.608 9.984 16.64 10.016 ;
  LAYER M2 ;
        RECT 18.976 10.048 19.008 10.08 ;
  LAYER M2 ;
        RECT 16.608 10.112 16.64 10.144 ;
  LAYER M2 ;
        RECT 18.976 10.176 19.008 10.208 ;
  LAYER M2 ;
        RECT 16.608 10.24 16.64 10.272 ;
  LAYER M2 ;
        RECT 18.976 10.304 19.008 10.336 ;
  LAYER M2 ;
        RECT 16.608 10.368 16.64 10.4 ;
  LAYER M2 ;
        RECT 18.976 10.432 19.008 10.464 ;
  LAYER M2 ;
        RECT 16.608 10.496 16.64 10.528 ;
  LAYER M2 ;
        RECT 18.976 10.56 19.008 10.592 ;
  LAYER M2 ;
        RECT 16.608 10.624 16.64 10.656 ;
  LAYER M2 ;
        RECT 18.976 10.688 19.008 10.72 ;
  LAYER M2 ;
        RECT 16.608 10.752 16.64 10.784 ;
  LAYER M2 ;
        RECT 18.976 10.816 19.008 10.848 ;
  LAYER M2 ;
        RECT 16.608 10.88 16.64 10.912 ;
  LAYER M2 ;
        RECT 18.976 10.944 19.008 10.976 ;
  LAYER M2 ;
        RECT 16.608 11.008 16.64 11.04 ;
  LAYER M2 ;
        RECT 18.976 11.072 19.008 11.104 ;
  LAYER M2 ;
        RECT 16.608 11.136 16.64 11.168 ;
  LAYER M2 ;
        RECT 18.976 11.2 19.008 11.232 ;
  LAYER M2 ;
        RECT 16.608 11.264 16.64 11.296 ;
  LAYER M2 ;
        RECT 18.976 11.328 19.008 11.36 ;
  LAYER M2 ;
        RECT 16.608 11.392 16.64 11.424 ;
  LAYER M2 ;
        RECT 18.976 11.456 19.008 11.488 ;
  LAYER M2 ;
        RECT 16.608 11.52 16.64 11.552 ;
  LAYER M2 ;
        RECT 18.976 11.584 19.008 11.616 ;
  LAYER M2 ;
        RECT 16.608 11.648 16.64 11.68 ;
  LAYER M2 ;
        RECT 18.976 11.712 19.008 11.744 ;
  LAYER M2 ;
        RECT 16.608 11.776 16.64 11.808 ;
  LAYER M2 ;
        RECT 18.976 11.84 19.008 11.872 ;
  LAYER M2 ;
        RECT 16.608 11.904 16.64 11.936 ;
  LAYER M2 ;
        RECT 18.976 11.968 19.008 12 ;
  LAYER M2 ;
        RECT 16.608 12.032 16.64 12.064 ;
  LAYER M2 ;
        RECT 16.56 9.66 19.056 12.264 ;
  LAYER M1 ;
        RECT 18.976 12.816 19.008 15.324 ;
  LAYER M3 ;
        RECT 18.976 15.272 19.008 15.304 ;
  LAYER M1 ;
        RECT 18.912 12.816 18.944 15.324 ;
  LAYER M3 ;
        RECT 18.912 12.836 18.944 12.868 ;
  LAYER M1 ;
        RECT 18.848 12.816 18.88 15.324 ;
  LAYER M3 ;
        RECT 18.848 15.272 18.88 15.304 ;
  LAYER M1 ;
        RECT 18.784 12.816 18.816 15.324 ;
  LAYER M3 ;
        RECT 18.784 12.836 18.816 12.868 ;
  LAYER M1 ;
        RECT 18.72 12.816 18.752 15.324 ;
  LAYER M3 ;
        RECT 18.72 15.272 18.752 15.304 ;
  LAYER M1 ;
        RECT 18.656 12.816 18.688 15.324 ;
  LAYER M3 ;
        RECT 18.656 12.836 18.688 12.868 ;
  LAYER M1 ;
        RECT 18.592 12.816 18.624 15.324 ;
  LAYER M3 ;
        RECT 18.592 15.272 18.624 15.304 ;
  LAYER M1 ;
        RECT 18.528 12.816 18.56 15.324 ;
  LAYER M3 ;
        RECT 18.528 12.836 18.56 12.868 ;
  LAYER M1 ;
        RECT 18.464 12.816 18.496 15.324 ;
  LAYER M3 ;
        RECT 18.464 15.272 18.496 15.304 ;
  LAYER M1 ;
        RECT 18.4 12.816 18.432 15.324 ;
  LAYER M3 ;
        RECT 18.4 12.836 18.432 12.868 ;
  LAYER M1 ;
        RECT 18.336 12.816 18.368 15.324 ;
  LAYER M3 ;
        RECT 18.336 15.272 18.368 15.304 ;
  LAYER M1 ;
        RECT 18.272 12.816 18.304 15.324 ;
  LAYER M3 ;
        RECT 18.272 12.836 18.304 12.868 ;
  LAYER M1 ;
        RECT 18.208 12.816 18.24 15.324 ;
  LAYER M3 ;
        RECT 18.208 15.272 18.24 15.304 ;
  LAYER M1 ;
        RECT 18.144 12.816 18.176 15.324 ;
  LAYER M3 ;
        RECT 18.144 12.836 18.176 12.868 ;
  LAYER M1 ;
        RECT 18.08 12.816 18.112 15.324 ;
  LAYER M3 ;
        RECT 18.08 15.272 18.112 15.304 ;
  LAYER M1 ;
        RECT 18.016 12.816 18.048 15.324 ;
  LAYER M3 ;
        RECT 18.016 12.836 18.048 12.868 ;
  LAYER M1 ;
        RECT 17.952 12.816 17.984 15.324 ;
  LAYER M3 ;
        RECT 17.952 15.272 17.984 15.304 ;
  LAYER M1 ;
        RECT 17.888 12.816 17.92 15.324 ;
  LAYER M3 ;
        RECT 17.888 12.836 17.92 12.868 ;
  LAYER M1 ;
        RECT 17.824 12.816 17.856 15.324 ;
  LAYER M3 ;
        RECT 17.824 15.272 17.856 15.304 ;
  LAYER M1 ;
        RECT 17.76 12.816 17.792 15.324 ;
  LAYER M3 ;
        RECT 17.76 12.836 17.792 12.868 ;
  LAYER M1 ;
        RECT 17.696 12.816 17.728 15.324 ;
  LAYER M3 ;
        RECT 17.696 15.272 17.728 15.304 ;
  LAYER M1 ;
        RECT 17.632 12.816 17.664 15.324 ;
  LAYER M3 ;
        RECT 17.632 12.836 17.664 12.868 ;
  LAYER M1 ;
        RECT 17.568 12.816 17.6 15.324 ;
  LAYER M3 ;
        RECT 17.568 15.272 17.6 15.304 ;
  LAYER M1 ;
        RECT 17.504 12.816 17.536 15.324 ;
  LAYER M3 ;
        RECT 17.504 12.836 17.536 12.868 ;
  LAYER M1 ;
        RECT 17.44 12.816 17.472 15.324 ;
  LAYER M3 ;
        RECT 17.44 15.272 17.472 15.304 ;
  LAYER M1 ;
        RECT 17.376 12.816 17.408 15.324 ;
  LAYER M3 ;
        RECT 17.376 12.836 17.408 12.868 ;
  LAYER M1 ;
        RECT 17.312 12.816 17.344 15.324 ;
  LAYER M3 ;
        RECT 17.312 15.272 17.344 15.304 ;
  LAYER M1 ;
        RECT 17.248 12.816 17.28 15.324 ;
  LAYER M3 ;
        RECT 17.248 12.836 17.28 12.868 ;
  LAYER M1 ;
        RECT 17.184 12.816 17.216 15.324 ;
  LAYER M3 ;
        RECT 17.184 15.272 17.216 15.304 ;
  LAYER M1 ;
        RECT 17.12 12.816 17.152 15.324 ;
  LAYER M3 ;
        RECT 17.12 12.836 17.152 12.868 ;
  LAYER M1 ;
        RECT 17.056 12.816 17.088 15.324 ;
  LAYER M3 ;
        RECT 17.056 15.272 17.088 15.304 ;
  LAYER M1 ;
        RECT 16.992 12.816 17.024 15.324 ;
  LAYER M3 ;
        RECT 16.992 12.836 17.024 12.868 ;
  LAYER M1 ;
        RECT 16.928 12.816 16.96 15.324 ;
  LAYER M3 ;
        RECT 16.928 15.272 16.96 15.304 ;
  LAYER M1 ;
        RECT 16.864 12.816 16.896 15.324 ;
  LAYER M3 ;
        RECT 16.864 12.836 16.896 12.868 ;
  LAYER M1 ;
        RECT 16.8 12.816 16.832 15.324 ;
  LAYER M3 ;
        RECT 16.8 15.272 16.832 15.304 ;
  LAYER M1 ;
        RECT 16.736 12.816 16.768 15.324 ;
  LAYER M3 ;
        RECT 16.736 12.836 16.768 12.868 ;
  LAYER M1 ;
        RECT 16.672 12.816 16.704 15.324 ;
  LAYER M3 ;
        RECT 16.672 15.272 16.704 15.304 ;
  LAYER M1 ;
        RECT 16.608 12.816 16.64 15.324 ;
  LAYER M3 ;
        RECT 18.976 12.9 19.008 12.932 ;
  LAYER M2 ;
        RECT 16.608 12.964 16.64 12.996 ;
  LAYER M2 ;
        RECT 18.976 13.028 19.008 13.06 ;
  LAYER M2 ;
        RECT 16.608 13.092 16.64 13.124 ;
  LAYER M2 ;
        RECT 18.976 13.156 19.008 13.188 ;
  LAYER M2 ;
        RECT 16.608 13.22 16.64 13.252 ;
  LAYER M2 ;
        RECT 18.976 13.284 19.008 13.316 ;
  LAYER M2 ;
        RECT 16.608 13.348 16.64 13.38 ;
  LAYER M2 ;
        RECT 18.976 13.412 19.008 13.444 ;
  LAYER M2 ;
        RECT 16.608 13.476 16.64 13.508 ;
  LAYER M2 ;
        RECT 18.976 13.54 19.008 13.572 ;
  LAYER M2 ;
        RECT 16.608 13.604 16.64 13.636 ;
  LAYER M2 ;
        RECT 18.976 13.668 19.008 13.7 ;
  LAYER M2 ;
        RECT 16.608 13.732 16.64 13.764 ;
  LAYER M2 ;
        RECT 18.976 13.796 19.008 13.828 ;
  LAYER M2 ;
        RECT 16.608 13.86 16.64 13.892 ;
  LAYER M2 ;
        RECT 18.976 13.924 19.008 13.956 ;
  LAYER M2 ;
        RECT 16.608 13.988 16.64 14.02 ;
  LAYER M2 ;
        RECT 18.976 14.052 19.008 14.084 ;
  LAYER M2 ;
        RECT 16.608 14.116 16.64 14.148 ;
  LAYER M2 ;
        RECT 18.976 14.18 19.008 14.212 ;
  LAYER M2 ;
        RECT 16.608 14.244 16.64 14.276 ;
  LAYER M2 ;
        RECT 18.976 14.308 19.008 14.34 ;
  LAYER M2 ;
        RECT 16.608 14.372 16.64 14.404 ;
  LAYER M2 ;
        RECT 18.976 14.436 19.008 14.468 ;
  LAYER M2 ;
        RECT 16.608 14.5 16.64 14.532 ;
  LAYER M2 ;
        RECT 18.976 14.564 19.008 14.596 ;
  LAYER M2 ;
        RECT 16.608 14.628 16.64 14.66 ;
  LAYER M2 ;
        RECT 18.976 14.692 19.008 14.724 ;
  LAYER M2 ;
        RECT 16.608 14.756 16.64 14.788 ;
  LAYER M2 ;
        RECT 18.976 14.82 19.008 14.852 ;
  LAYER M2 ;
        RECT 16.608 14.884 16.64 14.916 ;
  LAYER M2 ;
        RECT 18.976 14.948 19.008 14.98 ;
  LAYER M2 ;
        RECT 16.608 15.012 16.64 15.044 ;
  LAYER M2 ;
        RECT 18.976 15.076 19.008 15.108 ;
  LAYER M2 ;
        RECT 16.608 15.14 16.64 15.172 ;
  LAYER M2 ;
        RECT 16.56 12.768 19.056 15.372 ;
  LAYER M1 ;
        RECT 18.976 15.924 19.008 18.432 ;
  LAYER M3 ;
        RECT 18.976 18.38 19.008 18.412 ;
  LAYER M1 ;
        RECT 18.912 15.924 18.944 18.432 ;
  LAYER M3 ;
        RECT 18.912 15.944 18.944 15.976 ;
  LAYER M1 ;
        RECT 18.848 15.924 18.88 18.432 ;
  LAYER M3 ;
        RECT 18.848 18.38 18.88 18.412 ;
  LAYER M1 ;
        RECT 18.784 15.924 18.816 18.432 ;
  LAYER M3 ;
        RECT 18.784 15.944 18.816 15.976 ;
  LAYER M1 ;
        RECT 18.72 15.924 18.752 18.432 ;
  LAYER M3 ;
        RECT 18.72 18.38 18.752 18.412 ;
  LAYER M1 ;
        RECT 18.656 15.924 18.688 18.432 ;
  LAYER M3 ;
        RECT 18.656 15.944 18.688 15.976 ;
  LAYER M1 ;
        RECT 18.592 15.924 18.624 18.432 ;
  LAYER M3 ;
        RECT 18.592 18.38 18.624 18.412 ;
  LAYER M1 ;
        RECT 18.528 15.924 18.56 18.432 ;
  LAYER M3 ;
        RECT 18.528 15.944 18.56 15.976 ;
  LAYER M1 ;
        RECT 18.464 15.924 18.496 18.432 ;
  LAYER M3 ;
        RECT 18.464 18.38 18.496 18.412 ;
  LAYER M1 ;
        RECT 18.4 15.924 18.432 18.432 ;
  LAYER M3 ;
        RECT 18.4 15.944 18.432 15.976 ;
  LAYER M1 ;
        RECT 18.336 15.924 18.368 18.432 ;
  LAYER M3 ;
        RECT 18.336 18.38 18.368 18.412 ;
  LAYER M1 ;
        RECT 18.272 15.924 18.304 18.432 ;
  LAYER M3 ;
        RECT 18.272 15.944 18.304 15.976 ;
  LAYER M1 ;
        RECT 18.208 15.924 18.24 18.432 ;
  LAYER M3 ;
        RECT 18.208 18.38 18.24 18.412 ;
  LAYER M1 ;
        RECT 18.144 15.924 18.176 18.432 ;
  LAYER M3 ;
        RECT 18.144 15.944 18.176 15.976 ;
  LAYER M1 ;
        RECT 18.08 15.924 18.112 18.432 ;
  LAYER M3 ;
        RECT 18.08 18.38 18.112 18.412 ;
  LAYER M1 ;
        RECT 18.016 15.924 18.048 18.432 ;
  LAYER M3 ;
        RECT 18.016 15.944 18.048 15.976 ;
  LAYER M1 ;
        RECT 17.952 15.924 17.984 18.432 ;
  LAYER M3 ;
        RECT 17.952 18.38 17.984 18.412 ;
  LAYER M1 ;
        RECT 17.888 15.924 17.92 18.432 ;
  LAYER M3 ;
        RECT 17.888 15.944 17.92 15.976 ;
  LAYER M1 ;
        RECT 17.824 15.924 17.856 18.432 ;
  LAYER M3 ;
        RECT 17.824 18.38 17.856 18.412 ;
  LAYER M1 ;
        RECT 17.76 15.924 17.792 18.432 ;
  LAYER M3 ;
        RECT 17.76 15.944 17.792 15.976 ;
  LAYER M1 ;
        RECT 17.696 15.924 17.728 18.432 ;
  LAYER M3 ;
        RECT 17.696 18.38 17.728 18.412 ;
  LAYER M1 ;
        RECT 17.632 15.924 17.664 18.432 ;
  LAYER M3 ;
        RECT 17.632 15.944 17.664 15.976 ;
  LAYER M1 ;
        RECT 17.568 15.924 17.6 18.432 ;
  LAYER M3 ;
        RECT 17.568 18.38 17.6 18.412 ;
  LAYER M1 ;
        RECT 17.504 15.924 17.536 18.432 ;
  LAYER M3 ;
        RECT 17.504 15.944 17.536 15.976 ;
  LAYER M1 ;
        RECT 17.44 15.924 17.472 18.432 ;
  LAYER M3 ;
        RECT 17.44 18.38 17.472 18.412 ;
  LAYER M1 ;
        RECT 17.376 15.924 17.408 18.432 ;
  LAYER M3 ;
        RECT 17.376 15.944 17.408 15.976 ;
  LAYER M1 ;
        RECT 17.312 15.924 17.344 18.432 ;
  LAYER M3 ;
        RECT 17.312 18.38 17.344 18.412 ;
  LAYER M1 ;
        RECT 17.248 15.924 17.28 18.432 ;
  LAYER M3 ;
        RECT 17.248 15.944 17.28 15.976 ;
  LAYER M1 ;
        RECT 17.184 15.924 17.216 18.432 ;
  LAYER M3 ;
        RECT 17.184 18.38 17.216 18.412 ;
  LAYER M1 ;
        RECT 17.12 15.924 17.152 18.432 ;
  LAYER M3 ;
        RECT 17.12 15.944 17.152 15.976 ;
  LAYER M1 ;
        RECT 17.056 15.924 17.088 18.432 ;
  LAYER M3 ;
        RECT 17.056 18.38 17.088 18.412 ;
  LAYER M1 ;
        RECT 16.992 15.924 17.024 18.432 ;
  LAYER M3 ;
        RECT 16.992 15.944 17.024 15.976 ;
  LAYER M1 ;
        RECT 16.928 15.924 16.96 18.432 ;
  LAYER M3 ;
        RECT 16.928 18.38 16.96 18.412 ;
  LAYER M1 ;
        RECT 16.864 15.924 16.896 18.432 ;
  LAYER M3 ;
        RECT 16.864 15.944 16.896 15.976 ;
  LAYER M1 ;
        RECT 16.8 15.924 16.832 18.432 ;
  LAYER M3 ;
        RECT 16.8 18.38 16.832 18.412 ;
  LAYER M1 ;
        RECT 16.736 15.924 16.768 18.432 ;
  LAYER M3 ;
        RECT 16.736 15.944 16.768 15.976 ;
  LAYER M1 ;
        RECT 16.672 15.924 16.704 18.432 ;
  LAYER M3 ;
        RECT 16.672 18.38 16.704 18.412 ;
  LAYER M1 ;
        RECT 16.608 15.924 16.64 18.432 ;
  LAYER M3 ;
        RECT 18.976 16.008 19.008 16.04 ;
  LAYER M2 ;
        RECT 16.608 16.072 16.64 16.104 ;
  LAYER M2 ;
        RECT 18.976 16.136 19.008 16.168 ;
  LAYER M2 ;
        RECT 16.608 16.2 16.64 16.232 ;
  LAYER M2 ;
        RECT 18.976 16.264 19.008 16.296 ;
  LAYER M2 ;
        RECT 16.608 16.328 16.64 16.36 ;
  LAYER M2 ;
        RECT 18.976 16.392 19.008 16.424 ;
  LAYER M2 ;
        RECT 16.608 16.456 16.64 16.488 ;
  LAYER M2 ;
        RECT 18.976 16.52 19.008 16.552 ;
  LAYER M2 ;
        RECT 16.608 16.584 16.64 16.616 ;
  LAYER M2 ;
        RECT 18.976 16.648 19.008 16.68 ;
  LAYER M2 ;
        RECT 16.608 16.712 16.64 16.744 ;
  LAYER M2 ;
        RECT 18.976 16.776 19.008 16.808 ;
  LAYER M2 ;
        RECT 16.608 16.84 16.64 16.872 ;
  LAYER M2 ;
        RECT 18.976 16.904 19.008 16.936 ;
  LAYER M2 ;
        RECT 16.608 16.968 16.64 17 ;
  LAYER M2 ;
        RECT 18.976 17.032 19.008 17.064 ;
  LAYER M2 ;
        RECT 16.608 17.096 16.64 17.128 ;
  LAYER M2 ;
        RECT 18.976 17.16 19.008 17.192 ;
  LAYER M2 ;
        RECT 16.608 17.224 16.64 17.256 ;
  LAYER M2 ;
        RECT 18.976 17.288 19.008 17.32 ;
  LAYER M2 ;
        RECT 16.608 17.352 16.64 17.384 ;
  LAYER M2 ;
        RECT 18.976 17.416 19.008 17.448 ;
  LAYER M2 ;
        RECT 16.608 17.48 16.64 17.512 ;
  LAYER M2 ;
        RECT 18.976 17.544 19.008 17.576 ;
  LAYER M2 ;
        RECT 16.608 17.608 16.64 17.64 ;
  LAYER M2 ;
        RECT 18.976 17.672 19.008 17.704 ;
  LAYER M2 ;
        RECT 16.608 17.736 16.64 17.768 ;
  LAYER M2 ;
        RECT 18.976 17.8 19.008 17.832 ;
  LAYER M2 ;
        RECT 16.608 17.864 16.64 17.896 ;
  LAYER M2 ;
        RECT 18.976 17.928 19.008 17.96 ;
  LAYER M2 ;
        RECT 16.608 17.992 16.64 18.024 ;
  LAYER M2 ;
        RECT 18.976 18.056 19.008 18.088 ;
  LAYER M2 ;
        RECT 16.608 18.12 16.64 18.152 ;
  LAYER M2 ;
        RECT 18.976 18.184 19.008 18.216 ;
  LAYER M2 ;
        RECT 16.608 18.248 16.64 18.28 ;
  LAYER M2 ;
        RECT 16.56 15.876 19.056 18.48 ;
  LAYER M1 ;
        RECT 24.928 32.22 24.96 32.292 ;
  LAYER M2 ;
        RECT 24.908 32.24 24.98 32.272 ;
  LAYER M2 ;
        RECT 22.192 32.24 24.944 32.272 ;
  LAYER M1 ;
        RECT 22.176 32.22 22.208 32.292 ;
  LAYER M2 ;
        RECT 22.156 32.24 22.228 32.272 ;
  LAYER M1 ;
        RECT 24.928 29.112 24.96 29.184 ;
  LAYER M2 ;
        RECT 24.908 29.132 24.98 29.164 ;
  LAYER M2 ;
        RECT 22.192 29.132 24.944 29.164 ;
  LAYER M1 ;
        RECT 22.176 29.112 22.208 29.184 ;
  LAYER M2 ;
        RECT 22.156 29.132 22.228 29.164 ;
  LAYER M1 ;
        RECT 21.952 32.22 21.984 32.292 ;
  LAYER M2 ;
        RECT 21.932 32.24 22.004 32.272 ;
  LAYER M1 ;
        RECT 21.952 32.256 21.984 32.424 ;
  LAYER M1 ;
        RECT 21.952 32.388 21.984 32.46 ;
  LAYER M2 ;
        RECT 21.932 32.408 22.004 32.44 ;
  LAYER M2 ;
        RECT 21.968 32.408 22.192 32.44 ;
  LAYER M1 ;
        RECT 22.176 32.388 22.208 32.46 ;
  LAYER M2 ;
        RECT 22.156 32.408 22.228 32.44 ;
  LAYER M1 ;
        RECT 21.952 29.112 21.984 29.184 ;
  LAYER M2 ;
        RECT 21.932 29.132 22.004 29.164 ;
  LAYER M1 ;
        RECT 21.952 29.148 21.984 29.316 ;
  LAYER M1 ;
        RECT 21.952 29.28 21.984 29.352 ;
  LAYER M2 ;
        RECT 21.932 29.3 22.004 29.332 ;
  LAYER M2 ;
        RECT 21.968 29.3 22.192 29.332 ;
  LAYER M1 ;
        RECT 22.176 29.28 22.208 29.352 ;
  LAYER M2 ;
        RECT 22.156 29.3 22.228 29.332 ;
  LAYER M1 ;
        RECT 22.176 39.024 22.208 39.096 ;
  LAYER M2 ;
        RECT 22.156 39.044 22.228 39.076 ;
  LAYER M1 ;
        RECT 22.176 38.808 22.208 39.06 ;
  LAYER M1 ;
        RECT 22.176 29.148 22.208 38.808 ;
  LAYER M1 ;
        RECT 27.904 29.112 27.936 29.184 ;
  LAYER M2 ;
        RECT 27.884 29.132 27.956 29.164 ;
  LAYER M2 ;
        RECT 25.168 29.132 27.92 29.164 ;
  LAYER M1 ;
        RECT 25.152 29.112 25.184 29.184 ;
  LAYER M2 ;
        RECT 25.132 29.132 25.204 29.164 ;
  LAYER M1 ;
        RECT 27.904 32.22 27.936 32.292 ;
  LAYER M2 ;
        RECT 27.884 32.24 27.956 32.272 ;
  LAYER M2 ;
        RECT 25.168 32.24 27.92 32.272 ;
  LAYER M1 ;
        RECT 25.152 32.22 25.184 32.292 ;
  LAYER M2 ;
        RECT 25.132 32.24 25.204 32.272 ;
  LAYER M1 ;
        RECT 25.152 39.024 25.184 39.096 ;
  LAYER M2 ;
        RECT 25.132 39.044 25.204 39.076 ;
  LAYER M1 ;
        RECT 25.152 38.808 25.184 39.06 ;
  LAYER M1 ;
        RECT 25.152 29.148 25.184 38.808 ;
  LAYER M2 ;
        RECT 22.192 39.044 25.168 39.076 ;
  LAYER M1 ;
        RECT 21.952 26.004 21.984 26.076 ;
  LAYER M2 ;
        RECT 21.932 26.024 22.004 26.056 ;
  LAYER M2 ;
        RECT 19.216 26.024 21.968 26.056 ;
  LAYER M1 ;
        RECT 19.2 26.004 19.232 26.076 ;
  LAYER M2 ;
        RECT 19.18 26.024 19.252 26.056 ;
  LAYER M1 ;
        RECT 21.952 35.328 21.984 35.4 ;
  LAYER M2 ;
        RECT 21.932 35.348 22.004 35.38 ;
  LAYER M2 ;
        RECT 19.216 35.348 21.968 35.38 ;
  LAYER M1 ;
        RECT 19.2 35.328 19.232 35.4 ;
  LAYER M2 ;
        RECT 19.18 35.348 19.252 35.38 ;
  LAYER M1 ;
        RECT 19.2 39.192 19.232 39.264 ;
  LAYER M2 ;
        RECT 19.18 39.212 19.252 39.244 ;
  LAYER M1 ;
        RECT 19.2 38.808 19.232 39.228 ;
  LAYER M1 ;
        RECT 19.2 26.04 19.232 38.808 ;
  LAYER M1 ;
        RECT 27.904 35.328 27.936 35.4 ;
  LAYER M2 ;
        RECT 27.884 35.348 27.956 35.38 ;
  LAYER M1 ;
        RECT 27.904 35.364 27.936 35.532 ;
  LAYER M1 ;
        RECT 27.904 35.496 27.936 35.568 ;
  LAYER M2 ;
        RECT 27.884 35.516 27.956 35.548 ;
  LAYER M2 ;
        RECT 27.92 35.516 28.144 35.548 ;
  LAYER M1 ;
        RECT 28.128 35.496 28.16 35.568 ;
  LAYER M2 ;
        RECT 28.108 35.516 28.18 35.548 ;
  LAYER M1 ;
        RECT 27.904 26.004 27.936 26.076 ;
  LAYER M2 ;
        RECT 27.884 26.024 27.956 26.056 ;
  LAYER M1 ;
        RECT 27.904 26.04 27.936 26.208 ;
  LAYER M1 ;
        RECT 27.904 26.172 27.936 26.244 ;
  LAYER M2 ;
        RECT 27.884 26.192 27.956 26.224 ;
  LAYER M2 ;
        RECT 27.92 26.192 28.144 26.224 ;
  LAYER M1 ;
        RECT 28.128 26.172 28.16 26.244 ;
  LAYER M2 ;
        RECT 28.108 26.192 28.18 26.224 ;
  LAYER M1 ;
        RECT 28.128 39.192 28.16 39.264 ;
  LAYER M2 ;
        RECT 28.108 39.212 28.18 39.244 ;
  LAYER M1 ;
        RECT 28.128 38.808 28.16 39.228 ;
  LAYER M1 ;
        RECT 28.128 26.208 28.16 38.808 ;
  LAYER M2 ;
        RECT 19.216 39.212 28.144 39.244 ;
  LAYER M1 ;
        RECT 24.928 35.328 24.96 35.4 ;
  LAYER M2 ;
        RECT 24.908 35.348 24.98 35.38 ;
  LAYER M2 ;
        RECT 24.944 35.348 27.92 35.38 ;
  LAYER M1 ;
        RECT 27.904 35.328 27.936 35.4 ;
  LAYER M2 ;
        RECT 27.884 35.348 27.956 35.38 ;
  LAYER M1 ;
        RECT 24.928 26.004 24.96 26.076 ;
  LAYER M2 ;
        RECT 24.908 26.024 24.98 26.056 ;
  LAYER M2 ;
        RECT 21.968 26.024 24.944 26.056 ;
  LAYER M1 ;
        RECT 21.952 26.004 21.984 26.076 ;
  LAYER M2 ;
        RECT 21.932 26.024 22.004 26.056 ;
  LAYER M1 ;
        RECT 18.976 38.436 19.008 38.508 ;
  LAYER M2 ;
        RECT 18.956 38.456 19.028 38.488 ;
  LAYER M2 ;
        RECT 16.24 38.456 18.992 38.488 ;
  LAYER M1 ;
        RECT 16.224 38.436 16.256 38.508 ;
  LAYER M2 ;
        RECT 16.204 38.456 16.276 38.488 ;
  LAYER M1 ;
        RECT 18.976 35.328 19.008 35.4 ;
  LAYER M2 ;
        RECT 18.956 35.348 19.028 35.38 ;
  LAYER M2 ;
        RECT 16.24 35.348 18.992 35.38 ;
  LAYER M1 ;
        RECT 16.224 35.328 16.256 35.4 ;
  LAYER M2 ;
        RECT 16.204 35.348 16.276 35.38 ;
  LAYER M1 ;
        RECT 18.976 32.22 19.008 32.292 ;
  LAYER M2 ;
        RECT 18.956 32.24 19.028 32.272 ;
  LAYER M2 ;
        RECT 16.24 32.24 18.992 32.272 ;
  LAYER M1 ;
        RECT 16.224 32.22 16.256 32.292 ;
  LAYER M2 ;
        RECT 16.204 32.24 16.276 32.272 ;
  LAYER M1 ;
        RECT 18.976 29.112 19.008 29.184 ;
  LAYER M2 ;
        RECT 18.956 29.132 19.028 29.164 ;
  LAYER M2 ;
        RECT 16.24 29.132 18.992 29.164 ;
  LAYER M1 ;
        RECT 16.224 29.112 16.256 29.184 ;
  LAYER M2 ;
        RECT 16.204 29.132 16.276 29.164 ;
  LAYER M1 ;
        RECT 18.976 26.004 19.008 26.076 ;
  LAYER M2 ;
        RECT 18.956 26.024 19.028 26.056 ;
  LAYER M2 ;
        RECT 16.24 26.024 18.992 26.056 ;
  LAYER M1 ;
        RECT 16.224 26.004 16.256 26.076 ;
  LAYER M2 ;
        RECT 16.204 26.024 16.276 26.056 ;
  LAYER M1 ;
        RECT 18.976 22.896 19.008 22.968 ;
  LAYER M2 ;
        RECT 18.956 22.916 19.028 22.948 ;
  LAYER M2 ;
        RECT 16.24 22.916 18.992 22.948 ;
  LAYER M1 ;
        RECT 16.224 22.896 16.256 22.968 ;
  LAYER M2 ;
        RECT 16.204 22.916 16.276 22.948 ;
  LAYER M1 ;
        RECT 16.224 39.36 16.256 39.432 ;
  LAYER M2 ;
        RECT 16.204 39.38 16.276 39.412 ;
  LAYER M1 ;
        RECT 16.224 38.808 16.256 39.396 ;
  LAYER M1 ;
        RECT 16.224 22.932 16.256 38.808 ;
  LAYER M1 ;
        RECT 30.88 38.436 30.912 38.508 ;
  LAYER M2 ;
        RECT 30.86 38.456 30.932 38.488 ;
  LAYER M1 ;
        RECT 30.88 38.472 30.912 38.64 ;
  LAYER M1 ;
        RECT 30.88 38.604 30.912 38.676 ;
  LAYER M2 ;
        RECT 30.86 38.624 30.932 38.656 ;
  LAYER M2 ;
        RECT 30.896 38.624 31.12 38.656 ;
  LAYER M1 ;
        RECT 31.104 38.604 31.136 38.676 ;
  LAYER M2 ;
        RECT 31.084 38.624 31.156 38.656 ;
  LAYER M1 ;
        RECT 30.88 35.328 30.912 35.4 ;
  LAYER M2 ;
        RECT 30.86 35.348 30.932 35.38 ;
  LAYER M1 ;
        RECT 30.88 35.364 30.912 35.532 ;
  LAYER M1 ;
        RECT 30.88 35.496 30.912 35.568 ;
  LAYER M2 ;
        RECT 30.86 35.516 30.932 35.548 ;
  LAYER M2 ;
        RECT 30.896 35.516 31.12 35.548 ;
  LAYER M1 ;
        RECT 31.104 35.496 31.136 35.568 ;
  LAYER M2 ;
        RECT 31.084 35.516 31.156 35.548 ;
  LAYER M1 ;
        RECT 30.88 32.22 30.912 32.292 ;
  LAYER M2 ;
        RECT 30.86 32.24 30.932 32.272 ;
  LAYER M1 ;
        RECT 30.88 32.256 30.912 32.424 ;
  LAYER M1 ;
        RECT 30.88 32.388 30.912 32.46 ;
  LAYER M2 ;
        RECT 30.86 32.408 30.932 32.44 ;
  LAYER M2 ;
        RECT 30.896 32.408 31.12 32.44 ;
  LAYER M1 ;
        RECT 31.104 32.388 31.136 32.46 ;
  LAYER M2 ;
        RECT 31.084 32.408 31.156 32.44 ;
  LAYER M1 ;
        RECT 30.88 29.112 30.912 29.184 ;
  LAYER M2 ;
        RECT 30.86 29.132 30.932 29.164 ;
  LAYER M1 ;
        RECT 30.88 29.148 30.912 29.316 ;
  LAYER M1 ;
        RECT 30.88 29.28 30.912 29.352 ;
  LAYER M2 ;
        RECT 30.86 29.3 30.932 29.332 ;
  LAYER M2 ;
        RECT 30.896 29.3 31.12 29.332 ;
  LAYER M1 ;
        RECT 31.104 29.28 31.136 29.352 ;
  LAYER M2 ;
        RECT 31.084 29.3 31.156 29.332 ;
  LAYER M1 ;
        RECT 30.88 26.004 30.912 26.076 ;
  LAYER M2 ;
        RECT 30.86 26.024 30.932 26.056 ;
  LAYER M1 ;
        RECT 30.88 26.04 30.912 26.208 ;
  LAYER M1 ;
        RECT 30.88 26.172 30.912 26.244 ;
  LAYER M2 ;
        RECT 30.86 26.192 30.932 26.224 ;
  LAYER M2 ;
        RECT 30.896 26.192 31.12 26.224 ;
  LAYER M1 ;
        RECT 31.104 26.172 31.136 26.244 ;
  LAYER M2 ;
        RECT 31.084 26.192 31.156 26.224 ;
  LAYER M1 ;
        RECT 30.88 22.896 30.912 22.968 ;
  LAYER M2 ;
        RECT 30.86 22.916 30.932 22.948 ;
  LAYER M1 ;
        RECT 30.88 22.932 30.912 23.1 ;
  LAYER M1 ;
        RECT 30.88 23.064 30.912 23.136 ;
  LAYER M2 ;
        RECT 30.86 23.084 30.932 23.116 ;
  LAYER M2 ;
        RECT 30.896 23.084 31.12 23.116 ;
  LAYER M1 ;
        RECT 31.104 23.064 31.136 23.136 ;
  LAYER M2 ;
        RECT 31.084 23.084 31.156 23.116 ;
  LAYER M1 ;
        RECT 31.104 39.36 31.136 39.432 ;
  LAYER M2 ;
        RECT 31.084 39.38 31.156 39.412 ;
  LAYER M1 ;
        RECT 31.104 38.808 31.136 39.396 ;
  LAYER M1 ;
        RECT 31.104 23.1 31.136 38.808 ;
  LAYER M2 ;
        RECT 16.24 39.38 31.12 39.412 ;
  LAYER M1 ;
        RECT 21.952 38.436 21.984 38.508 ;
  LAYER M2 ;
        RECT 21.932 38.456 22.004 38.488 ;
  LAYER M2 ;
        RECT 18.992 38.456 21.968 38.488 ;
  LAYER M1 ;
        RECT 18.976 38.436 19.008 38.508 ;
  LAYER M2 ;
        RECT 18.956 38.456 19.028 38.488 ;
  LAYER M1 ;
        RECT 21.952 22.896 21.984 22.968 ;
  LAYER M2 ;
        RECT 21.932 22.916 22.004 22.948 ;
  LAYER M2 ;
        RECT 18.992 22.916 21.968 22.948 ;
  LAYER M1 ;
        RECT 18.976 22.896 19.008 22.968 ;
  LAYER M2 ;
        RECT 18.956 22.916 19.028 22.948 ;
  LAYER M1 ;
        RECT 24.928 22.896 24.96 22.968 ;
  LAYER M2 ;
        RECT 24.908 22.916 24.98 22.948 ;
  LAYER M2 ;
        RECT 21.968 22.916 24.944 22.948 ;
  LAYER M1 ;
        RECT 21.952 22.896 21.984 22.968 ;
  LAYER M2 ;
        RECT 21.932 22.916 22.004 22.948 ;
  LAYER M1 ;
        RECT 27.904 22.896 27.936 22.968 ;
  LAYER M2 ;
        RECT 27.884 22.916 27.956 22.948 ;
  LAYER M2 ;
        RECT 24.944 22.916 27.92 22.948 ;
  LAYER M1 ;
        RECT 24.928 22.896 24.96 22.968 ;
  LAYER M2 ;
        RECT 24.908 22.916 24.98 22.948 ;
  LAYER M1 ;
        RECT 27.904 38.436 27.936 38.508 ;
  LAYER M2 ;
        RECT 27.884 38.456 27.956 38.488 ;
  LAYER M2 ;
        RECT 27.92 38.456 30.896 38.488 ;
  LAYER M1 ;
        RECT 30.88 38.436 30.912 38.508 ;
  LAYER M2 ;
        RECT 30.86 38.456 30.932 38.488 ;
  LAYER M1 ;
        RECT 24.928 38.436 24.96 38.508 ;
  LAYER M2 ;
        RECT 24.908 38.456 24.98 38.488 ;
  LAYER M2 ;
        RECT 24.944 38.456 27.92 38.488 ;
  LAYER M1 ;
        RECT 27.904 38.436 27.936 38.508 ;
  LAYER M2 ;
        RECT 27.884 38.456 27.956 38.488 ;
  LAYER M1 ;
        RECT 22.56 29.784 22.592 29.856 ;
  LAYER M2 ;
        RECT 22.54 29.804 22.612 29.836 ;
  LAYER M2 ;
        RECT 22.352 29.804 22.576 29.836 ;
  LAYER M1 ;
        RECT 22.336 29.784 22.368 29.856 ;
  LAYER M2 ;
        RECT 22.316 29.804 22.388 29.836 ;
  LAYER M1 ;
        RECT 22.56 26.676 22.592 26.748 ;
  LAYER M2 ;
        RECT 22.54 26.696 22.612 26.728 ;
  LAYER M2 ;
        RECT 22.352 26.696 22.576 26.728 ;
  LAYER M1 ;
        RECT 22.336 26.676 22.368 26.748 ;
  LAYER M2 ;
        RECT 22.316 26.696 22.388 26.728 ;
  LAYER M1 ;
        RECT 19.584 29.784 19.616 29.856 ;
  LAYER M2 ;
        RECT 19.564 29.804 19.636 29.836 ;
  LAYER M1 ;
        RECT 19.584 29.652 19.616 29.82 ;
  LAYER M1 ;
        RECT 19.584 29.616 19.616 29.688 ;
  LAYER M2 ;
        RECT 19.564 29.636 19.636 29.668 ;
  LAYER M2 ;
        RECT 19.6 29.636 22.352 29.668 ;
  LAYER M1 ;
        RECT 22.336 29.616 22.368 29.688 ;
  LAYER M2 ;
        RECT 22.316 29.636 22.388 29.668 ;
  LAYER M1 ;
        RECT 19.584 26.676 19.616 26.748 ;
  LAYER M2 ;
        RECT 19.564 26.696 19.636 26.728 ;
  LAYER M1 ;
        RECT 19.584 26.544 19.616 26.712 ;
  LAYER M1 ;
        RECT 19.584 26.508 19.616 26.58 ;
  LAYER M2 ;
        RECT 19.564 26.528 19.636 26.56 ;
  LAYER M2 ;
        RECT 19.6 26.528 22.352 26.56 ;
  LAYER M1 ;
        RECT 22.336 26.508 22.368 26.58 ;
  LAYER M2 ;
        RECT 22.316 26.528 22.388 26.56 ;
  LAYER M1 ;
        RECT 22.336 19.872 22.368 19.944 ;
  LAYER M2 ;
        RECT 22.316 19.892 22.388 19.924 ;
  LAYER M1 ;
        RECT 22.336 19.908 22.368 20.16 ;
  LAYER M1 ;
        RECT 22.336 20.16 22.368 29.82 ;
  LAYER M1 ;
        RECT 25.536 26.676 25.568 26.748 ;
  LAYER M2 ;
        RECT 25.516 26.696 25.588 26.728 ;
  LAYER M2 ;
        RECT 25.328 26.696 25.552 26.728 ;
  LAYER M1 ;
        RECT 25.312 26.676 25.344 26.748 ;
  LAYER M2 ;
        RECT 25.292 26.696 25.364 26.728 ;
  LAYER M1 ;
        RECT 25.536 29.784 25.568 29.856 ;
  LAYER M2 ;
        RECT 25.516 29.804 25.588 29.836 ;
  LAYER M2 ;
        RECT 25.328 29.804 25.552 29.836 ;
  LAYER M1 ;
        RECT 25.312 29.784 25.344 29.856 ;
  LAYER M2 ;
        RECT 25.292 29.804 25.364 29.836 ;
  LAYER M1 ;
        RECT 25.312 19.872 25.344 19.944 ;
  LAYER M2 ;
        RECT 25.292 19.892 25.364 19.924 ;
  LAYER M1 ;
        RECT 25.312 19.908 25.344 20.16 ;
  LAYER M1 ;
        RECT 25.312 20.16 25.344 29.82 ;
  LAYER M2 ;
        RECT 22.352 19.892 25.328 19.924 ;
  LAYER M1 ;
        RECT 19.584 23.568 19.616 23.64 ;
  LAYER M2 ;
        RECT 19.564 23.588 19.636 23.62 ;
  LAYER M2 ;
        RECT 19.376 23.588 19.6 23.62 ;
  LAYER M1 ;
        RECT 19.36 23.568 19.392 23.64 ;
  LAYER M2 ;
        RECT 19.34 23.588 19.412 23.62 ;
  LAYER M1 ;
        RECT 19.584 32.892 19.616 32.964 ;
  LAYER M2 ;
        RECT 19.564 32.912 19.636 32.944 ;
  LAYER M2 ;
        RECT 19.376 32.912 19.6 32.944 ;
  LAYER M1 ;
        RECT 19.36 32.892 19.392 32.964 ;
  LAYER M2 ;
        RECT 19.34 32.912 19.412 32.944 ;
  LAYER M1 ;
        RECT 19.36 19.704 19.392 19.776 ;
  LAYER M2 ;
        RECT 19.34 19.724 19.412 19.756 ;
  LAYER M1 ;
        RECT 19.36 19.74 19.392 20.16 ;
  LAYER M1 ;
        RECT 19.36 20.16 19.392 32.928 ;
  LAYER M1 ;
        RECT 25.536 32.892 25.568 32.964 ;
  LAYER M2 ;
        RECT 25.516 32.912 25.588 32.944 ;
  LAYER M1 ;
        RECT 25.536 32.76 25.568 32.928 ;
  LAYER M1 ;
        RECT 25.536 32.724 25.568 32.796 ;
  LAYER M2 ;
        RECT 25.516 32.744 25.588 32.776 ;
  LAYER M2 ;
        RECT 25.552 32.744 28.304 32.776 ;
  LAYER M1 ;
        RECT 28.288 32.724 28.32 32.796 ;
  LAYER M2 ;
        RECT 28.268 32.744 28.34 32.776 ;
  LAYER M1 ;
        RECT 25.536 23.568 25.568 23.64 ;
  LAYER M2 ;
        RECT 25.516 23.588 25.588 23.62 ;
  LAYER M1 ;
        RECT 25.536 23.436 25.568 23.604 ;
  LAYER M1 ;
        RECT 25.536 23.4 25.568 23.472 ;
  LAYER M2 ;
        RECT 25.516 23.42 25.588 23.452 ;
  LAYER M2 ;
        RECT 25.552 23.42 28.304 23.452 ;
  LAYER M1 ;
        RECT 28.288 23.4 28.32 23.472 ;
  LAYER M2 ;
        RECT 28.268 23.42 28.34 23.452 ;
  LAYER M1 ;
        RECT 28.288 19.704 28.32 19.776 ;
  LAYER M2 ;
        RECT 28.268 19.724 28.34 19.756 ;
  LAYER M1 ;
        RECT 28.288 19.74 28.32 20.16 ;
  LAYER M1 ;
        RECT 28.288 20.16 28.32 32.76 ;
  LAYER M2 ;
        RECT 19.376 19.724 28.304 19.756 ;
  LAYER M1 ;
        RECT 22.56 32.892 22.592 32.964 ;
  LAYER M2 ;
        RECT 22.54 32.912 22.612 32.944 ;
  LAYER M2 ;
        RECT 22.576 32.912 25.552 32.944 ;
  LAYER M1 ;
        RECT 25.536 32.892 25.568 32.964 ;
  LAYER M2 ;
        RECT 25.516 32.912 25.588 32.944 ;
  LAYER M1 ;
        RECT 22.56 23.568 22.592 23.64 ;
  LAYER M2 ;
        RECT 22.54 23.588 22.612 23.62 ;
  LAYER M2 ;
        RECT 19.6 23.588 22.576 23.62 ;
  LAYER M1 ;
        RECT 19.584 23.568 19.616 23.64 ;
  LAYER M2 ;
        RECT 19.564 23.588 19.636 23.62 ;
  LAYER M1 ;
        RECT 16.608 36 16.64 36.072 ;
  LAYER M2 ;
        RECT 16.588 36.02 16.66 36.052 ;
  LAYER M2 ;
        RECT 16.4 36.02 16.624 36.052 ;
  LAYER M1 ;
        RECT 16.384 36 16.416 36.072 ;
  LAYER M2 ;
        RECT 16.364 36.02 16.436 36.052 ;
  LAYER M1 ;
        RECT 16.608 32.892 16.64 32.964 ;
  LAYER M2 ;
        RECT 16.588 32.912 16.66 32.944 ;
  LAYER M2 ;
        RECT 16.4 32.912 16.624 32.944 ;
  LAYER M1 ;
        RECT 16.384 32.892 16.416 32.964 ;
  LAYER M2 ;
        RECT 16.364 32.912 16.436 32.944 ;
  LAYER M1 ;
        RECT 16.608 29.784 16.64 29.856 ;
  LAYER M2 ;
        RECT 16.588 29.804 16.66 29.836 ;
  LAYER M2 ;
        RECT 16.4 29.804 16.624 29.836 ;
  LAYER M1 ;
        RECT 16.384 29.784 16.416 29.856 ;
  LAYER M2 ;
        RECT 16.364 29.804 16.436 29.836 ;
  LAYER M1 ;
        RECT 16.608 26.676 16.64 26.748 ;
  LAYER M2 ;
        RECT 16.588 26.696 16.66 26.728 ;
  LAYER M2 ;
        RECT 16.4 26.696 16.624 26.728 ;
  LAYER M1 ;
        RECT 16.384 26.676 16.416 26.748 ;
  LAYER M2 ;
        RECT 16.364 26.696 16.436 26.728 ;
  LAYER M1 ;
        RECT 16.608 23.568 16.64 23.64 ;
  LAYER M2 ;
        RECT 16.588 23.588 16.66 23.62 ;
  LAYER M2 ;
        RECT 16.4 23.588 16.624 23.62 ;
  LAYER M1 ;
        RECT 16.384 23.568 16.416 23.64 ;
  LAYER M2 ;
        RECT 16.364 23.588 16.436 23.62 ;
  LAYER M1 ;
        RECT 16.608 20.46 16.64 20.532 ;
  LAYER M2 ;
        RECT 16.588 20.48 16.66 20.512 ;
  LAYER M2 ;
        RECT 16.4 20.48 16.624 20.512 ;
  LAYER M1 ;
        RECT 16.384 20.46 16.416 20.532 ;
  LAYER M2 ;
        RECT 16.364 20.48 16.436 20.512 ;
  LAYER M1 ;
        RECT 16.384 19.536 16.416 19.608 ;
  LAYER M2 ;
        RECT 16.364 19.556 16.436 19.588 ;
  LAYER M1 ;
        RECT 16.384 19.572 16.416 20.16 ;
  LAYER M1 ;
        RECT 16.384 20.16 16.416 36.036 ;
  LAYER M1 ;
        RECT 28.512 36 28.544 36.072 ;
  LAYER M2 ;
        RECT 28.492 36.02 28.564 36.052 ;
  LAYER M1 ;
        RECT 28.512 35.868 28.544 36.036 ;
  LAYER M1 ;
        RECT 28.512 35.832 28.544 35.904 ;
  LAYER M2 ;
        RECT 28.492 35.852 28.564 35.884 ;
  LAYER M2 ;
        RECT 28.528 35.852 31.28 35.884 ;
  LAYER M1 ;
        RECT 31.264 35.832 31.296 35.904 ;
  LAYER M2 ;
        RECT 31.244 35.852 31.316 35.884 ;
  LAYER M1 ;
        RECT 28.512 32.892 28.544 32.964 ;
  LAYER M2 ;
        RECT 28.492 32.912 28.564 32.944 ;
  LAYER M1 ;
        RECT 28.512 32.76 28.544 32.928 ;
  LAYER M1 ;
        RECT 28.512 32.724 28.544 32.796 ;
  LAYER M2 ;
        RECT 28.492 32.744 28.564 32.776 ;
  LAYER M2 ;
        RECT 28.528 32.744 31.28 32.776 ;
  LAYER M1 ;
        RECT 31.264 32.724 31.296 32.796 ;
  LAYER M2 ;
        RECT 31.244 32.744 31.316 32.776 ;
  LAYER M1 ;
        RECT 28.512 29.784 28.544 29.856 ;
  LAYER M2 ;
        RECT 28.492 29.804 28.564 29.836 ;
  LAYER M1 ;
        RECT 28.512 29.652 28.544 29.82 ;
  LAYER M1 ;
        RECT 28.512 29.616 28.544 29.688 ;
  LAYER M2 ;
        RECT 28.492 29.636 28.564 29.668 ;
  LAYER M2 ;
        RECT 28.528 29.636 31.28 29.668 ;
  LAYER M1 ;
        RECT 31.264 29.616 31.296 29.688 ;
  LAYER M2 ;
        RECT 31.244 29.636 31.316 29.668 ;
  LAYER M1 ;
        RECT 28.512 26.676 28.544 26.748 ;
  LAYER M2 ;
        RECT 28.492 26.696 28.564 26.728 ;
  LAYER M1 ;
        RECT 28.512 26.544 28.544 26.712 ;
  LAYER M1 ;
        RECT 28.512 26.508 28.544 26.58 ;
  LAYER M2 ;
        RECT 28.492 26.528 28.564 26.56 ;
  LAYER M2 ;
        RECT 28.528 26.528 31.28 26.56 ;
  LAYER M1 ;
        RECT 31.264 26.508 31.296 26.58 ;
  LAYER M2 ;
        RECT 31.244 26.528 31.316 26.56 ;
  LAYER M1 ;
        RECT 28.512 23.568 28.544 23.64 ;
  LAYER M2 ;
        RECT 28.492 23.588 28.564 23.62 ;
  LAYER M1 ;
        RECT 28.512 23.436 28.544 23.604 ;
  LAYER M1 ;
        RECT 28.512 23.4 28.544 23.472 ;
  LAYER M2 ;
        RECT 28.492 23.42 28.564 23.452 ;
  LAYER M2 ;
        RECT 28.528 23.42 31.28 23.452 ;
  LAYER M1 ;
        RECT 31.264 23.4 31.296 23.472 ;
  LAYER M2 ;
        RECT 31.244 23.42 31.316 23.452 ;
  LAYER M1 ;
        RECT 28.512 20.46 28.544 20.532 ;
  LAYER M2 ;
        RECT 28.492 20.48 28.564 20.512 ;
  LAYER M1 ;
        RECT 28.512 20.328 28.544 20.496 ;
  LAYER M1 ;
        RECT 28.512 20.292 28.544 20.364 ;
  LAYER M2 ;
        RECT 28.492 20.312 28.564 20.344 ;
  LAYER M2 ;
        RECT 28.528 20.312 31.28 20.344 ;
  LAYER M1 ;
        RECT 31.264 20.292 31.296 20.364 ;
  LAYER M2 ;
        RECT 31.244 20.312 31.316 20.344 ;
  LAYER M1 ;
        RECT 31.264 19.536 31.296 19.608 ;
  LAYER M2 ;
        RECT 31.244 19.556 31.316 19.588 ;
  LAYER M1 ;
        RECT 31.264 19.572 31.296 20.16 ;
  LAYER M1 ;
        RECT 31.264 20.16 31.296 35.868 ;
  LAYER M2 ;
        RECT 16.4 19.556 31.28 19.588 ;
  LAYER M1 ;
        RECT 19.584 36 19.616 36.072 ;
  LAYER M2 ;
        RECT 19.564 36.02 19.636 36.052 ;
  LAYER M2 ;
        RECT 16.624 36.02 19.6 36.052 ;
  LAYER M1 ;
        RECT 16.608 36 16.64 36.072 ;
  LAYER M2 ;
        RECT 16.588 36.02 16.66 36.052 ;
  LAYER M1 ;
        RECT 19.584 20.46 19.616 20.532 ;
  LAYER M2 ;
        RECT 19.564 20.48 19.636 20.512 ;
  LAYER M2 ;
        RECT 16.624 20.48 19.6 20.512 ;
  LAYER M1 ;
        RECT 16.608 20.46 16.64 20.532 ;
  LAYER M2 ;
        RECT 16.588 20.48 16.66 20.512 ;
  LAYER M1 ;
        RECT 22.56 20.46 22.592 20.532 ;
  LAYER M2 ;
        RECT 22.54 20.48 22.612 20.512 ;
  LAYER M2 ;
        RECT 19.6 20.48 22.576 20.512 ;
  LAYER M1 ;
        RECT 19.584 20.46 19.616 20.532 ;
  LAYER M2 ;
        RECT 19.564 20.48 19.636 20.512 ;
  LAYER M1 ;
        RECT 25.536 20.46 25.568 20.532 ;
  LAYER M2 ;
        RECT 25.516 20.48 25.588 20.512 ;
  LAYER M2 ;
        RECT 22.576 20.48 25.552 20.512 ;
  LAYER M1 ;
        RECT 22.56 20.46 22.592 20.532 ;
  LAYER M2 ;
        RECT 22.54 20.48 22.612 20.512 ;
  LAYER M1 ;
        RECT 25.536 36 25.568 36.072 ;
  LAYER M2 ;
        RECT 25.516 36.02 25.588 36.052 ;
  LAYER M2 ;
        RECT 25.552 36.02 28.528 36.052 ;
  LAYER M1 ;
        RECT 28.512 36 28.544 36.072 ;
  LAYER M2 ;
        RECT 28.492 36.02 28.564 36.052 ;
  LAYER M1 ;
        RECT 22.56 36 22.592 36.072 ;
  LAYER M2 ;
        RECT 22.54 36.02 22.612 36.052 ;
  LAYER M2 ;
        RECT 22.576 36.02 25.552 36.052 ;
  LAYER M1 ;
        RECT 25.536 36 25.568 36.072 ;
  LAYER M2 ;
        RECT 25.516 36.02 25.588 36.052 ;
  LAYER M1 ;
        RECT 16.608 36 16.64 38.508 ;
  LAYER M3 ;
        RECT 16.608 36.02 16.64 36.052 ;
  LAYER M1 ;
        RECT 16.672 36 16.704 38.508 ;
  LAYER M3 ;
        RECT 16.672 38.456 16.704 38.488 ;
  LAYER M1 ;
        RECT 16.736 36 16.768 38.508 ;
  LAYER M3 ;
        RECT 16.736 36.02 16.768 36.052 ;
  LAYER M1 ;
        RECT 16.8 36 16.832 38.508 ;
  LAYER M3 ;
        RECT 16.8 38.456 16.832 38.488 ;
  LAYER M1 ;
        RECT 16.864 36 16.896 38.508 ;
  LAYER M3 ;
        RECT 16.864 36.02 16.896 36.052 ;
  LAYER M1 ;
        RECT 16.928 36 16.96 38.508 ;
  LAYER M3 ;
        RECT 16.928 38.456 16.96 38.488 ;
  LAYER M1 ;
        RECT 16.992 36 17.024 38.508 ;
  LAYER M3 ;
        RECT 16.992 36.02 17.024 36.052 ;
  LAYER M1 ;
        RECT 17.056 36 17.088 38.508 ;
  LAYER M3 ;
        RECT 17.056 38.456 17.088 38.488 ;
  LAYER M1 ;
        RECT 17.12 36 17.152 38.508 ;
  LAYER M3 ;
        RECT 17.12 36.02 17.152 36.052 ;
  LAYER M1 ;
        RECT 17.184 36 17.216 38.508 ;
  LAYER M3 ;
        RECT 17.184 38.456 17.216 38.488 ;
  LAYER M1 ;
        RECT 17.248 36 17.28 38.508 ;
  LAYER M3 ;
        RECT 17.248 36.02 17.28 36.052 ;
  LAYER M1 ;
        RECT 17.312 36 17.344 38.508 ;
  LAYER M3 ;
        RECT 17.312 38.456 17.344 38.488 ;
  LAYER M1 ;
        RECT 17.376 36 17.408 38.508 ;
  LAYER M3 ;
        RECT 17.376 36.02 17.408 36.052 ;
  LAYER M1 ;
        RECT 17.44 36 17.472 38.508 ;
  LAYER M3 ;
        RECT 17.44 38.456 17.472 38.488 ;
  LAYER M1 ;
        RECT 17.504 36 17.536 38.508 ;
  LAYER M3 ;
        RECT 17.504 36.02 17.536 36.052 ;
  LAYER M1 ;
        RECT 17.568 36 17.6 38.508 ;
  LAYER M3 ;
        RECT 17.568 38.456 17.6 38.488 ;
  LAYER M1 ;
        RECT 17.632 36 17.664 38.508 ;
  LAYER M3 ;
        RECT 17.632 36.02 17.664 36.052 ;
  LAYER M1 ;
        RECT 17.696 36 17.728 38.508 ;
  LAYER M3 ;
        RECT 17.696 38.456 17.728 38.488 ;
  LAYER M1 ;
        RECT 17.76 36 17.792 38.508 ;
  LAYER M3 ;
        RECT 17.76 36.02 17.792 36.052 ;
  LAYER M1 ;
        RECT 17.824 36 17.856 38.508 ;
  LAYER M3 ;
        RECT 17.824 38.456 17.856 38.488 ;
  LAYER M1 ;
        RECT 17.888 36 17.92 38.508 ;
  LAYER M3 ;
        RECT 17.888 36.02 17.92 36.052 ;
  LAYER M1 ;
        RECT 17.952 36 17.984 38.508 ;
  LAYER M3 ;
        RECT 17.952 38.456 17.984 38.488 ;
  LAYER M1 ;
        RECT 18.016 36 18.048 38.508 ;
  LAYER M3 ;
        RECT 18.016 36.02 18.048 36.052 ;
  LAYER M1 ;
        RECT 18.08 36 18.112 38.508 ;
  LAYER M3 ;
        RECT 18.08 38.456 18.112 38.488 ;
  LAYER M1 ;
        RECT 18.144 36 18.176 38.508 ;
  LAYER M3 ;
        RECT 18.144 36.02 18.176 36.052 ;
  LAYER M1 ;
        RECT 18.208 36 18.24 38.508 ;
  LAYER M3 ;
        RECT 18.208 38.456 18.24 38.488 ;
  LAYER M1 ;
        RECT 18.272 36 18.304 38.508 ;
  LAYER M3 ;
        RECT 18.272 36.02 18.304 36.052 ;
  LAYER M1 ;
        RECT 18.336 36 18.368 38.508 ;
  LAYER M3 ;
        RECT 18.336 38.456 18.368 38.488 ;
  LAYER M1 ;
        RECT 18.4 36 18.432 38.508 ;
  LAYER M3 ;
        RECT 18.4 36.02 18.432 36.052 ;
  LAYER M1 ;
        RECT 18.464 36 18.496 38.508 ;
  LAYER M3 ;
        RECT 18.464 38.456 18.496 38.488 ;
  LAYER M1 ;
        RECT 18.528 36 18.56 38.508 ;
  LAYER M3 ;
        RECT 18.528 36.02 18.56 36.052 ;
  LAYER M1 ;
        RECT 18.592 36 18.624 38.508 ;
  LAYER M3 ;
        RECT 18.592 38.456 18.624 38.488 ;
  LAYER M1 ;
        RECT 18.656 36 18.688 38.508 ;
  LAYER M3 ;
        RECT 18.656 36.02 18.688 36.052 ;
  LAYER M1 ;
        RECT 18.72 36 18.752 38.508 ;
  LAYER M3 ;
        RECT 18.72 38.456 18.752 38.488 ;
  LAYER M1 ;
        RECT 18.784 36 18.816 38.508 ;
  LAYER M3 ;
        RECT 18.784 36.02 18.816 36.052 ;
  LAYER M1 ;
        RECT 18.848 36 18.88 38.508 ;
  LAYER M3 ;
        RECT 18.848 38.456 18.88 38.488 ;
  LAYER M1 ;
        RECT 18.912 36 18.944 38.508 ;
  LAYER M3 ;
        RECT 18.912 36.02 18.944 36.052 ;
  LAYER M1 ;
        RECT 18.976 36 19.008 38.508 ;
  LAYER M3 ;
        RECT 16.608 38.392 16.64 38.424 ;
  LAYER M2 ;
        RECT 18.976 38.328 19.008 38.36 ;
  LAYER M2 ;
        RECT 16.608 38.264 16.64 38.296 ;
  LAYER M2 ;
        RECT 18.976 38.2 19.008 38.232 ;
  LAYER M2 ;
        RECT 16.608 38.136 16.64 38.168 ;
  LAYER M2 ;
        RECT 18.976 38.072 19.008 38.104 ;
  LAYER M2 ;
        RECT 16.608 38.008 16.64 38.04 ;
  LAYER M2 ;
        RECT 18.976 37.944 19.008 37.976 ;
  LAYER M2 ;
        RECT 16.608 37.88 16.64 37.912 ;
  LAYER M2 ;
        RECT 18.976 37.816 19.008 37.848 ;
  LAYER M2 ;
        RECT 16.608 37.752 16.64 37.784 ;
  LAYER M2 ;
        RECT 18.976 37.688 19.008 37.72 ;
  LAYER M2 ;
        RECT 16.608 37.624 16.64 37.656 ;
  LAYER M2 ;
        RECT 18.976 37.56 19.008 37.592 ;
  LAYER M2 ;
        RECT 16.608 37.496 16.64 37.528 ;
  LAYER M2 ;
        RECT 18.976 37.432 19.008 37.464 ;
  LAYER M2 ;
        RECT 16.608 37.368 16.64 37.4 ;
  LAYER M2 ;
        RECT 18.976 37.304 19.008 37.336 ;
  LAYER M2 ;
        RECT 16.608 37.24 16.64 37.272 ;
  LAYER M2 ;
        RECT 18.976 37.176 19.008 37.208 ;
  LAYER M2 ;
        RECT 16.608 37.112 16.64 37.144 ;
  LAYER M2 ;
        RECT 18.976 37.048 19.008 37.08 ;
  LAYER M2 ;
        RECT 16.608 36.984 16.64 37.016 ;
  LAYER M2 ;
        RECT 18.976 36.92 19.008 36.952 ;
  LAYER M2 ;
        RECT 16.608 36.856 16.64 36.888 ;
  LAYER M2 ;
        RECT 18.976 36.792 19.008 36.824 ;
  LAYER M2 ;
        RECT 16.608 36.728 16.64 36.76 ;
  LAYER M2 ;
        RECT 18.976 36.664 19.008 36.696 ;
  LAYER M2 ;
        RECT 16.608 36.6 16.64 36.632 ;
  LAYER M2 ;
        RECT 18.976 36.536 19.008 36.568 ;
  LAYER M2 ;
        RECT 16.608 36.472 16.64 36.504 ;
  LAYER M2 ;
        RECT 18.976 36.408 19.008 36.44 ;
  LAYER M2 ;
        RECT 16.608 36.344 16.64 36.376 ;
  LAYER M2 ;
        RECT 18.976 36.28 19.008 36.312 ;
  LAYER M2 ;
        RECT 16.608 36.216 16.64 36.248 ;
  LAYER M2 ;
        RECT 18.976 36.152 19.008 36.184 ;
  LAYER M2 ;
        RECT 16.56 35.952 19.056 38.556 ;
  LAYER M1 ;
        RECT 16.608 32.892 16.64 35.4 ;
  LAYER M3 ;
        RECT 16.608 32.912 16.64 32.944 ;
  LAYER M1 ;
        RECT 16.672 32.892 16.704 35.4 ;
  LAYER M3 ;
        RECT 16.672 35.348 16.704 35.38 ;
  LAYER M1 ;
        RECT 16.736 32.892 16.768 35.4 ;
  LAYER M3 ;
        RECT 16.736 32.912 16.768 32.944 ;
  LAYER M1 ;
        RECT 16.8 32.892 16.832 35.4 ;
  LAYER M3 ;
        RECT 16.8 35.348 16.832 35.38 ;
  LAYER M1 ;
        RECT 16.864 32.892 16.896 35.4 ;
  LAYER M3 ;
        RECT 16.864 32.912 16.896 32.944 ;
  LAYER M1 ;
        RECT 16.928 32.892 16.96 35.4 ;
  LAYER M3 ;
        RECT 16.928 35.348 16.96 35.38 ;
  LAYER M1 ;
        RECT 16.992 32.892 17.024 35.4 ;
  LAYER M3 ;
        RECT 16.992 32.912 17.024 32.944 ;
  LAYER M1 ;
        RECT 17.056 32.892 17.088 35.4 ;
  LAYER M3 ;
        RECT 17.056 35.348 17.088 35.38 ;
  LAYER M1 ;
        RECT 17.12 32.892 17.152 35.4 ;
  LAYER M3 ;
        RECT 17.12 32.912 17.152 32.944 ;
  LAYER M1 ;
        RECT 17.184 32.892 17.216 35.4 ;
  LAYER M3 ;
        RECT 17.184 35.348 17.216 35.38 ;
  LAYER M1 ;
        RECT 17.248 32.892 17.28 35.4 ;
  LAYER M3 ;
        RECT 17.248 32.912 17.28 32.944 ;
  LAYER M1 ;
        RECT 17.312 32.892 17.344 35.4 ;
  LAYER M3 ;
        RECT 17.312 35.348 17.344 35.38 ;
  LAYER M1 ;
        RECT 17.376 32.892 17.408 35.4 ;
  LAYER M3 ;
        RECT 17.376 32.912 17.408 32.944 ;
  LAYER M1 ;
        RECT 17.44 32.892 17.472 35.4 ;
  LAYER M3 ;
        RECT 17.44 35.348 17.472 35.38 ;
  LAYER M1 ;
        RECT 17.504 32.892 17.536 35.4 ;
  LAYER M3 ;
        RECT 17.504 32.912 17.536 32.944 ;
  LAYER M1 ;
        RECT 17.568 32.892 17.6 35.4 ;
  LAYER M3 ;
        RECT 17.568 35.348 17.6 35.38 ;
  LAYER M1 ;
        RECT 17.632 32.892 17.664 35.4 ;
  LAYER M3 ;
        RECT 17.632 32.912 17.664 32.944 ;
  LAYER M1 ;
        RECT 17.696 32.892 17.728 35.4 ;
  LAYER M3 ;
        RECT 17.696 35.348 17.728 35.38 ;
  LAYER M1 ;
        RECT 17.76 32.892 17.792 35.4 ;
  LAYER M3 ;
        RECT 17.76 32.912 17.792 32.944 ;
  LAYER M1 ;
        RECT 17.824 32.892 17.856 35.4 ;
  LAYER M3 ;
        RECT 17.824 35.348 17.856 35.38 ;
  LAYER M1 ;
        RECT 17.888 32.892 17.92 35.4 ;
  LAYER M3 ;
        RECT 17.888 32.912 17.92 32.944 ;
  LAYER M1 ;
        RECT 17.952 32.892 17.984 35.4 ;
  LAYER M3 ;
        RECT 17.952 35.348 17.984 35.38 ;
  LAYER M1 ;
        RECT 18.016 32.892 18.048 35.4 ;
  LAYER M3 ;
        RECT 18.016 32.912 18.048 32.944 ;
  LAYER M1 ;
        RECT 18.08 32.892 18.112 35.4 ;
  LAYER M3 ;
        RECT 18.08 35.348 18.112 35.38 ;
  LAYER M1 ;
        RECT 18.144 32.892 18.176 35.4 ;
  LAYER M3 ;
        RECT 18.144 32.912 18.176 32.944 ;
  LAYER M1 ;
        RECT 18.208 32.892 18.24 35.4 ;
  LAYER M3 ;
        RECT 18.208 35.348 18.24 35.38 ;
  LAYER M1 ;
        RECT 18.272 32.892 18.304 35.4 ;
  LAYER M3 ;
        RECT 18.272 32.912 18.304 32.944 ;
  LAYER M1 ;
        RECT 18.336 32.892 18.368 35.4 ;
  LAYER M3 ;
        RECT 18.336 35.348 18.368 35.38 ;
  LAYER M1 ;
        RECT 18.4 32.892 18.432 35.4 ;
  LAYER M3 ;
        RECT 18.4 32.912 18.432 32.944 ;
  LAYER M1 ;
        RECT 18.464 32.892 18.496 35.4 ;
  LAYER M3 ;
        RECT 18.464 35.348 18.496 35.38 ;
  LAYER M1 ;
        RECT 18.528 32.892 18.56 35.4 ;
  LAYER M3 ;
        RECT 18.528 32.912 18.56 32.944 ;
  LAYER M1 ;
        RECT 18.592 32.892 18.624 35.4 ;
  LAYER M3 ;
        RECT 18.592 35.348 18.624 35.38 ;
  LAYER M1 ;
        RECT 18.656 32.892 18.688 35.4 ;
  LAYER M3 ;
        RECT 18.656 32.912 18.688 32.944 ;
  LAYER M1 ;
        RECT 18.72 32.892 18.752 35.4 ;
  LAYER M3 ;
        RECT 18.72 35.348 18.752 35.38 ;
  LAYER M1 ;
        RECT 18.784 32.892 18.816 35.4 ;
  LAYER M3 ;
        RECT 18.784 32.912 18.816 32.944 ;
  LAYER M1 ;
        RECT 18.848 32.892 18.88 35.4 ;
  LAYER M3 ;
        RECT 18.848 35.348 18.88 35.38 ;
  LAYER M1 ;
        RECT 18.912 32.892 18.944 35.4 ;
  LAYER M3 ;
        RECT 18.912 32.912 18.944 32.944 ;
  LAYER M1 ;
        RECT 18.976 32.892 19.008 35.4 ;
  LAYER M3 ;
        RECT 16.608 35.284 16.64 35.316 ;
  LAYER M2 ;
        RECT 18.976 35.22 19.008 35.252 ;
  LAYER M2 ;
        RECT 16.608 35.156 16.64 35.188 ;
  LAYER M2 ;
        RECT 18.976 35.092 19.008 35.124 ;
  LAYER M2 ;
        RECT 16.608 35.028 16.64 35.06 ;
  LAYER M2 ;
        RECT 18.976 34.964 19.008 34.996 ;
  LAYER M2 ;
        RECT 16.608 34.9 16.64 34.932 ;
  LAYER M2 ;
        RECT 18.976 34.836 19.008 34.868 ;
  LAYER M2 ;
        RECT 16.608 34.772 16.64 34.804 ;
  LAYER M2 ;
        RECT 18.976 34.708 19.008 34.74 ;
  LAYER M2 ;
        RECT 16.608 34.644 16.64 34.676 ;
  LAYER M2 ;
        RECT 18.976 34.58 19.008 34.612 ;
  LAYER M2 ;
        RECT 16.608 34.516 16.64 34.548 ;
  LAYER M2 ;
        RECT 18.976 34.452 19.008 34.484 ;
  LAYER M2 ;
        RECT 16.608 34.388 16.64 34.42 ;
  LAYER M2 ;
        RECT 18.976 34.324 19.008 34.356 ;
  LAYER M2 ;
        RECT 16.608 34.26 16.64 34.292 ;
  LAYER M2 ;
        RECT 18.976 34.196 19.008 34.228 ;
  LAYER M2 ;
        RECT 16.608 34.132 16.64 34.164 ;
  LAYER M2 ;
        RECT 18.976 34.068 19.008 34.1 ;
  LAYER M2 ;
        RECT 16.608 34.004 16.64 34.036 ;
  LAYER M2 ;
        RECT 18.976 33.94 19.008 33.972 ;
  LAYER M2 ;
        RECT 16.608 33.876 16.64 33.908 ;
  LAYER M2 ;
        RECT 18.976 33.812 19.008 33.844 ;
  LAYER M2 ;
        RECT 16.608 33.748 16.64 33.78 ;
  LAYER M2 ;
        RECT 18.976 33.684 19.008 33.716 ;
  LAYER M2 ;
        RECT 16.608 33.62 16.64 33.652 ;
  LAYER M2 ;
        RECT 18.976 33.556 19.008 33.588 ;
  LAYER M2 ;
        RECT 16.608 33.492 16.64 33.524 ;
  LAYER M2 ;
        RECT 18.976 33.428 19.008 33.46 ;
  LAYER M2 ;
        RECT 16.608 33.364 16.64 33.396 ;
  LAYER M2 ;
        RECT 18.976 33.3 19.008 33.332 ;
  LAYER M2 ;
        RECT 16.608 33.236 16.64 33.268 ;
  LAYER M2 ;
        RECT 18.976 33.172 19.008 33.204 ;
  LAYER M2 ;
        RECT 16.608 33.108 16.64 33.14 ;
  LAYER M2 ;
        RECT 18.976 33.044 19.008 33.076 ;
  LAYER M2 ;
        RECT 16.56 32.844 19.056 35.448 ;
  LAYER M1 ;
        RECT 16.608 29.784 16.64 32.292 ;
  LAYER M3 ;
        RECT 16.608 29.804 16.64 29.836 ;
  LAYER M1 ;
        RECT 16.672 29.784 16.704 32.292 ;
  LAYER M3 ;
        RECT 16.672 32.24 16.704 32.272 ;
  LAYER M1 ;
        RECT 16.736 29.784 16.768 32.292 ;
  LAYER M3 ;
        RECT 16.736 29.804 16.768 29.836 ;
  LAYER M1 ;
        RECT 16.8 29.784 16.832 32.292 ;
  LAYER M3 ;
        RECT 16.8 32.24 16.832 32.272 ;
  LAYER M1 ;
        RECT 16.864 29.784 16.896 32.292 ;
  LAYER M3 ;
        RECT 16.864 29.804 16.896 29.836 ;
  LAYER M1 ;
        RECT 16.928 29.784 16.96 32.292 ;
  LAYER M3 ;
        RECT 16.928 32.24 16.96 32.272 ;
  LAYER M1 ;
        RECT 16.992 29.784 17.024 32.292 ;
  LAYER M3 ;
        RECT 16.992 29.804 17.024 29.836 ;
  LAYER M1 ;
        RECT 17.056 29.784 17.088 32.292 ;
  LAYER M3 ;
        RECT 17.056 32.24 17.088 32.272 ;
  LAYER M1 ;
        RECT 17.12 29.784 17.152 32.292 ;
  LAYER M3 ;
        RECT 17.12 29.804 17.152 29.836 ;
  LAYER M1 ;
        RECT 17.184 29.784 17.216 32.292 ;
  LAYER M3 ;
        RECT 17.184 32.24 17.216 32.272 ;
  LAYER M1 ;
        RECT 17.248 29.784 17.28 32.292 ;
  LAYER M3 ;
        RECT 17.248 29.804 17.28 29.836 ;
  LAYER M1 ;
        RECT 17.312 29.784 17.344 32.292 ;
  LAYER M3 ;
        RECT 17.312 32.24 17.344 32.272 ;
  LAYER M1 ;
        RECT 17.376 29.784 17.408 32.292 ;
  LAYER M3 ;
        RECT 17.376 29.804 17.408 29.836 ;
  LAYER M1 ;
        RECT 17.44 29.784 17.472 32.292 ;
  LAYER M3 ;
        RECT 17.44 32.24 17.472 32.272 ;
  LAYER M1 ;
        RECT 17.504 29.784 17.536 32.292 ;
  LAYER M3 ;
        RECT 17.504 29.804 17.536 29.836 ;
  LAYER M1 ;
        RECT 17.568 29.784 17.6 32.292 ;
  LAYER M3 ;
        RECT 17.568 32.24 17.6 32.272 ;
  LAYER M1 ;
        RECT 17.632 29.784 17.664 32.292 ;
  LAYER M3 ;
        RECT 17.632 29.804 17.664 29.836 ;
  LAYER M1 ;
        RECT 17.696 29.784 17.728 32.292 ;
  LAYER M3 ;
        RECT 17.696 32.24 17.728 32.272 ;
  LAYER M1 ;
        RECT 17.76 29.784 17.792 32.292 ;
  LAYER M3 ;
        RECT 17.76 29.804 17.792 29.836 ;
  LAYER M1 ;
        RECT 17.824 29.784 17.856 32.292 ;
  LAYER M3 ;
        RECT 17.824 32.24 17.856 32.272 ;
  LAYER M1 ;
        RECT 17.888 29.784 17.92 32.292 ;
  LAYER M3 ;
        RECT 17.888 29.804 17.92 29.836 ;
  LAYER M1 ;
        RECT 17.952 29.784 17.984 32.292 ;
  LAYER M3 ;
        RECT 17.952 32.24 17.984 32.272 ;
  LAYER M1 ;
        RECT 18.016 29.784 18.048 32.292 ;
  LAYER M3 ;
        RECT 18.016 29.804 18.048 29.836 ;
  LAYER M1 ;
        RECT 18.08 29.784 18.112 32.292 ;
  LAYER M3 ;
        RECT 18.08 32.24 18.112 32.272 ;
  LAYER M1 ;
        RECT 18.144 29.784 18.176 32.292 ;
  LAYER M3 ;
        RECT 18.144 29.804 18.176 29.836 ;
  LAYER M1 ;
        RECT 18.208 29.784 18.24 32.292 ;
  LAYER M3 ;
        RECT 18.208 32.24 18.24 32.272 ;
  LAYER M1 ;
        RECT 18.272 29.784 18.304 32.292 ;
  LAYER M3 ;
        RECT 18.272 29.804 18.304 29.836 ;
  LAYER M1 ;
        RECT 18.336 29.784 18.368 32.292 ;
  LAYER M3 ;
        RECT 18.336 32.24 18.368 32.272 ;
  LAYER M1 ;
        RECT 18.4 29.784 18.432 32.292 ;
  LAYER M3 ;
        RECT 18.4 29.804 18.432 29.836 ;
  LAYER M1 ;
        RECT 18.464 29.784 18.496 32.292 ;
  LAYER M3 ;
        RECT 18.464 32.24 18.496 32.272 ;
  LAYER M1 ;
        RECT 18.528 29.784 18.56 32.292 ;
  LAYER M3 ;
        RECT 18.528 29.804 18.56 29.836 ;
  LAYER M1 ;
        RECT 18.592 29.784 18.624 32.292 ;
  LAYER M3 ;
        RECT 18.592 32.24 18.624 32.272 ;
  LAYER M1 ;
        RECT 18.656 29.784 18.688 32.292 ;
  LAYER M3 ;
        RECT 18.656 29.804 18.688 29.836 ;
  LAYER M1 ;
        RECT 18.72 29.784 18.752 32.292 ;
  LAYER M3 ;
        RECT 18.72 32.24 18.752 32.272 ;
  LAYER M1 ;
        RECT 18.784 29.784 18.816 32.292 ;
  LAYER M3 ;
        RECT 18.784 29.804 18.816 29.836 ;
  LAYER M1 ;
        RECT 18.848 29.784 18.88 32.292 ;
  LAYER M3 ;
        RECT 18.848 32.24 18.88 32.272 ;
  LAYER M1 ;
        RECT 18.912 29.784 18.944 32.292 ;
  LAYER M3 ;
        RECT 18.912 29.804 18.944 29.836 ;
  LAYER M1 ;
        RECT 18.976 29.784 19.008 32.292 ;
  LAYER M3 ;
        RECT 16.608 32.176 16.64 32.208 ;
  LAYER M2 ;
        RECT 18.976 32.112 19.008 32.144 ;
  LAYER M2 ;
        RECT 16.608 32.048 16.64 32.08 ;
  LAYER M2 ;
        RECT 18.976 31.984 19.008 32.016 ;
  LAYER M2 ;
        RECT 16.608 31.92 16.64 31.952 ;
  LAYER M2 ;
        RECT 18.976 31.856 19.008 31.888 ;
  LAYER M2 ;
        RECT 16.608 31.792 16.64 31.824 ;
  LAYER M2 ;
        RECT 18.976 31.728 19.008 31.76 ;
  LAYER M2 ;
        RECT 16.608 31.664 16.64 31.696 ;
  LAYER M2 ;
        RECT 18.976 31.6 19.008 31.632 ;
  LAYER M2 ;
        RECT 16.608 31.536 16.64 31.568 ;
  LAYER M2 ;
        RECT 18.976 31.472 19.008 31.504 ;
  LAYER M2 ;
        RECT 16.608 31.408 16.64 31.44 ;
  LAYER M2 ;
        RECT 18.976 31.344 19.008 31.376 ;
  LAYER M2 ;
        RECT 16.608 31.28 16.64 31.312 ;
  LAYER M2 ;
        RECT 18.976 31.216 19.008 31.248 ;
  LAYER M2 ;
        RECT 16.608 31.152 16.64 31.184 ;
  LAYER M2 ;
        RECT 18.976 31.088 19.008 31.12 ;
  LAYER M2 ;
        RECT 16.608 31.024 16.64 31.056 ;
  LAYER M2 ;
        RECT 18.976 30.96 19.008 30.992 ;
  LAYER M2 ;
        RECT 16.608 30.896 16.64 30.928 ;
  LAYER M2 ;
        RECT 18.976 30.832 19.008 30.864 ;
  LAYER M2 ;
        RECT 16.608 30.768 16.64 30.8 ;
  LAYER M2 ;
        RECT 18.976 30.704 19.008 30.736 ;
  LAYER M2 ;
        RECT 16.608 30.64 16.64 30.672 ;
  LAYER M2 ;
        RECT 18.976 30.576 19.008 30.608 ;
  LAYER M2 ;
        RECT 16.608 30.512 16.64 30.544 ;
  LAYER M2 ;
        RECT 18.976 30.448 19.008 30.48 ;
  LAYER M2 ;
        RECT 16.608 30.384 16.64 30.416 ;
  LAYER M2 ;
        RECT 18.976 30.32 19.008 30.352 ;
  LAYER M2 ;
        RECT 16.608 30.256 16.64 30.288 ;
  LAYER M2 ;
        RECT 18.976 30.192 19.008 30.224 ;
  LAYER M2 ;
        RECT 16.608 30.128 16.64 30.16 ;
  LAYER M2 ;
        RECT 18.976 30.064 19.008 30.096 ;
  LAYER M2 ;
        RECT 16.608 30 16.64 30.032 ;
  LAYER M2 ;
        RECT 18.976 29.936 19.008 29.968 ;
  LAYER M2 ;
        RECT 16.56 29.736 19.056 32.34 ;
  LAYER M1 ;
        RECT 16.608 26.676 16.64 29.184 ;
  LAYER M3 ;
        RECT 16.608 26.696 16.64 26.728 ;
  LAYER M1 ;
        RECT 16.672 26.676 16.704 29.184 ;
  LAYER M3 ;
        RECT 16.672 29.132 16.704 29.164 ;
  LAYER M1 ;
        RECT 16.736 26.676 16.768 29.184 ;
  LAYER M3 ;
        RECT 16.736 26.696 16.768 26.728 ;
  LAYER M1 ;
        RECT 16.8 26.676 16.832 29.184 ;
  LAYER M3 ;
        RECT 16.8 29.132 16.832 29.164 ;
  LAYER M1 ;
        RECT 16.864 26.676 16.896 29.184 ;
  LAYER M3 ;
        RECT 16.864 26.696 16.896 26.728 ;
  LAYER M1 ;
        RECT 16.928 26.676 16.96 29.184 ;
  LAYER M3 ;
        RECT 16.928 29.132 16.96 29.164 ;
  LAYER M1 ;
        RECT 16.992 26.676 17.024 29.184 ;
  LAYER M3 ;
        RECT 16.992 26.696 17.024 26.728 ;
  LAYER M1 ;
        RECT 17.056 26.676 17.088 29.184 ;
  LAYER M3 ;
        RECT 17.056 29.132 17.088 29.164 ;
  LAYER M1 ;
        RECT 17.12 26.676 17.152 29.184 ;
  LAYER M3 ;
        RECT 17.12 26.696 17.152 26.728 ;
  LAYER M1 ;
        RECT 17.184 26.676 17.216 29.184 ;
  LAYER M3 ;
        RECT 17.184 29.132 17.216 29.164 ;
  LAYER M1 ;
        RECT 17.248 26.676 17.28 29.184 ;
  LAYER M3 ;
        RECT 17.248 26.696 17.28 26.728 ;
  LAYER M1 ;
        RECT 17.312 26.676 17.344 29.184 ;
  LAYER M3 ;
        RECT 17.312 29.132 17.344 29.164 ;
  LAYER M1 ;
        RECT 17.376 26.676 17.408 29.184 ;
  LAYER M3 ;
        RECT 17.376 26.696 17.408 26.728 ;
  LAYER M1 ;
        RECT 17.44 26.676 17.472 29.184 ;
  LAYER M3 ;
        RECT 17.44 29.132 17.472 29.164 ;
  LAYER M1 ;
        RECT 17.504 26.676 17.536 29.184 ;
  LAYER M3 ;
        RECT 17.504 26.696 17.536 26.728 ;
  LAYER M1 ;
        RECT 17.568 26.676 17.6 29.184 ;
  LAYER M3 ;
        RECT 17.568 29.132 17.6 29.164 ;
  LAYER M1 ;
        RECT 17.632 26.676 17.664 29.184 ;
  LAYER M3 ;
        RECT 17.632 26.696 17.664 26.728 ;
  LAYER M1 ;
        RECT 17.696 26.676 17.728 29.184 ;
  LAYER M3 ;
        RECT 17.696 29.132 17.728 29.164 ;
  LAYER M1 ;
        RECT 17.76 26.676 17.792 29.184 ;
  LAYER M3 ;
        RECT 17.76 26.696 17.792 26.728 ;
  LAYER M1 ;
        RECT 17.824 26.676 17.856 29.184 ;
  LAYER M3 ;
        RECT 17.824 29.132 17.856 29.164 ;
  LAYER M1 ;
        RECT 17.888 26.676 17.92 29.184 ;
  LAYER M3 ;
        RECT 17.888 26.696 17.92 26.728 ;
  LAYER M1 ;
        RECT 17.952 26.676 17.984 29.184 ;
  LAYER M3 ;
        RECT 17.952 29.132 17.984 29.164 ;
  LAYER M1 ;
        RECT 18.016 26.676 18.048 29.184 ;
  LAYER M3 ;
        RECT 18.016 26.696 18.048 26.728 ;
  LAYER M1 ;
        RECT 18.08 26.676 18.112 29.184 ;
  LAYER M3 ;
        RECT 18.08 29.132 18.112 29.164 ;
  LAYER M1 ;
        RECT 18.144 26.676 18.176 29.184 ;
  LAYER M3 ;
        RECT 18.144 26.696 18.176 26.728 ;
  LAYER M1 ;
        RECT 18.208 26.676 18.24 29.184 ;
  LAYER M3 ;
        RECT 18.208 29.132 18.24 29.164 ;
  LAYER M1 ;
        RECT 18.272 26.676 18.304 29.184 ;
  LAYER M3 ;
        RECT 18.272 26.696 18.304 26.728 ;
  LAYER M1 ;
        RECT 18.336 26.676 18.368 29.184 ;
  LAYER M3 ;
        RECT 18.336 29.132 18.368 29.164 ;
  LAYER M1 ;
        RECT 18.4 26.676 18.432 29.184 ;
  LAYER M3 ;
        RECT 18.4 26.696 18.432 26.728 ;
  LAYER M1 ;
        RECT 18.464 26.676 18.496 29.184 ;
  LAYER M3 ;
        RECT 18.464 29.132 18.496 29.164 ;
  LAYER M1 ;
        RECT 18.528 26.676 18.56 29.184 ;
  LAYER M3 ;
        RECT 18.528 26.696 18.56 26.728 ;
  LAYER M1 ;
        RECT 18.592 26.676 18.624 29.184 ;
  LAYER M3 ;
        RECT 18.592 29.132 18.624 29.164 ;
  LAYER M1 ;
        RECT 18.656 26.676 18.688 29.184 ;
  LAYER M3 ;
        RECT 18.656 26.696 18.688 26.728 ;
  LAYER M1 ;
        RECT 18.72 26.676 18.752 29.184 ;
  LAYER M3 ;
        RECT 18.72 29.132 18.752 29.164 ;
  LAYER M1 ;
        RECT 18.784 26.676 18.816 29.184 ;
  LAYER M3 ;
        RECT 18.784 26.696 18.816 26.728 ;
  LAYER M1 ;
        RECT 18.848 26.676 18.88 29.184 ;
  LAYER M3 ;
        RECT 18.848 29.132 18.88 29.164 ;
  LAYER M1 ;
        RECT 18.912 26.676 18.944 29.184 ;
  LAYER M3 ;
        RECT 18.912 26.696 18.944 26.728 ;
  LAYER M1 ;
        RECT 18.976 26.676 19.008 29.184 ;
  LAYER M3 ;
        RECT 16.608 29.068 16.64 29.1 ;
  LAYER M2 ;
        RECT 18.976 29.004 19.008 29.036 ;
  LAYER M2 ;
        RECT 16.608 28.94 16.64 28.972 ;
  LAYER M2 ;
        RECT 18.976 28.876 19.008 28.908 ;
  LAYER M2 ;
        RECT 16.608 28.812 16.64 28.844 ;
  LAYER M2 ;
        RECT 18.976 28.748 19.008 28.78 ;
  LAYER M2 ;
        RECT 16.608 28.684 16.64 28.716 ;
  LAYER M2 ;
        RECT 18.976 28.62 19.008 28.652 ;
  LAYER M2 ;
        RECT 16.608 28.556 16.64 28.588 ;
  LAYER M2 ;
        RECT 18.976 28.492 19.008 28.524 ;
  LAYER M2 ;
        RECT 16.608 28.428 16.64 28.46 ;
  LAYER M2 ;
        RECT 18.976 28.364 19.008 28.396 ;
  LAYER M2 ;
        RECT 16.608 28.3 16.64 28.332 ;
  LAYER M2 ;
        RECT 18.976 28.236 19.008 28.268 ;
  LAYER M2 ;
        RECT 16.608 28.172 16.64 28.204 ;
  LAYER M2 ;
        RECT 18.976 28.108 19.008 28.14 ;
  LAYER M2 ;
        RECT 16.608 28.044 16.64 28.076 ;
  LAYER M2 ;
        RECT 18.976 27.98 19.008 28.012 ;
  LAYER M2 ;
        RECT 16.608 27.916 16.64 27.948 ;
  LAYER M2 ;
        RECT 18.976 27.852 19.008 27.884 ;
  LAYER M2 ;
        RECT 16.608 27.788 16.64 27.82 ;
  LAYER M2 ;
        RECT 18.976 27.724 19.008 27.756 ;
  LAYER M2 ;
        RECT 16.608 27.66 16.64 27.692 ;
  LAYER M2 ;
        RECT 18.976 27.596 19.008 27.628 ;
  LAYER M2 ;
        RECT 16.608 27.532 16.64 27.564 ;
  LAYER M2 ;
        RECT 18.976 27.468 19.008 27.5 ;
  LAYER M2 ;
        RECT 16.608 27.404 16.64 27.436 ;
  LAYER M2 ;
        RECT 18.976 27.34 19.008 27.372 ;
  LAYER M2 ;
        RECT 16.608 27.276 16.64 27.308 ;
  LAYER M2 ;
        RECT 18.976 27.212 19.008 27.244 ;
  LAYER M2 ;
        RECT 16.608 27.148 16.64 27.18 ;
  LAYER M2 ;
        RECT 18.976 27.084 19.008 27.116 ;
  LAYER M2 ;
        RECT 16.608 27.02 16.64 27.052 ;
  LAYER M2 ;
        RECT 18.976 26.956 19.008 26.988 ;
  LAYER M2 ;
        RECT 16.608 26.892 16.64 26.924 ;
  LAYER M2 ;
        RECT 18.976 26.828 19.008 26.86 ;
  LAYER M2 ;
        RECT 16.56 26.628 19.056 29.232 ;
  LAYER M1 ;
        RECT 16.608 23.568 16.64 26.076 ;
  LAYER M3 ;
        RECT 16.608 23.588 16.64 23.62 ;
  LAYER M1 ;
        RECT 16.672 23.568 16.704 26.076 ;
  LAYER M3 ;
        RECT 16.672 26.024 16.704 26.056 ;
  LAYER M1 ;
        RECT 16.736 23.568 16.768 26.076 ;
  LAYER M3 ;
        RECT 16.736 23.588 16.768 23.62 ;
  LAYER M1 ;
        RECT 16.8 23.568 16.832 26.076 ;
  LAYER M3 ;
        RECT 16.8 26.024 16.832 26.056 ;
  LAYER M1 ;
        RECT 16.864 23.568 16.896 26.076 ;
  LAYER M3 ;
        RECT 16.864 23.588 16.896 23.62 ;
  LAYER M1 ;
        RECT 16.928 23.568 16.96 26.076 ;
  LAYER M3 ;
        RECT 16.928 26.024 16.96 26.056 ;
  LAYER M1 ;
        RECT 16.992 23.568 17.024 26.076 ;
  LAYER M3 ;
        RECT 16.992 23.588 17.024 23.62 ;
  LAYER M1 ;
        RECT 17.056 23.568 17.088 26.076 ;
  LAYER M3 ;
        RECT 17.056 26.024 17.088 26.056 ;
  LAYER M1 ;
        RECT 17.12 23.568 17.152 26.076 ;
  LAYER M3 ;
        RECT 17.12 23.588 17.152 23.62 ;
  LAYER M1 ;
        RECT 17.184 23.568 17.216 26.076 ;
  LAYER M3 ;
        RECT 17.184 26.024 17.216 26.056 ;
  LAYER M1 ;
        RECT 17.248 23.568 17.28 26.076 ;
  LAYER M3 ;
        RECT 17.248 23.588 17.28 23.62 ;
  LAYER M1 ;
        RECT 17.312 23.568 17.344 26.076 ;
  LAYER M3 ;
        RECT 17.312 26.024 17.344 26.056 ;
  LAYER M1 ;
        RECT 17.376 23.568 17.408 26.076 ;
  LAYER M3 ;
        RECT 17.376 23.588 17.408 23.62 ;
  LAYER M1 ;
        RECT 17.44 23.568 17.472 26.076 ;
  LAYER M3 ;
        RECT 17.44 26.024 17.472 26.056 ;
  LAYER M1 ;
        RECT 17.504 23.568 17.536 26.076 ;
  LAYER M3 ;
        RECT 17.504 23.588 17.536 23.62 ;
  LAYER M1 ;
        RECT 17.568 23.568 17.6 26.076 ;
  LAYER M3 ;
        RECT 17.568 26.024 17.6 26.056 ;
  LAYER M1 ;
        RECT 17.632 23.568 17.664 26.076 ;
  LAYER M3 ;
        RECT 17.632 23.588 17.664 23.62 ;
  LAYER M1 ;
        RECT 17.696 23.568 17.728 26.076 ;
  LAYER M3 ;
        RECT 17.696 26.024 17.728 26.056 ;
  LAYER M1 ;
        RECT 17.76 23.568 17.792 26.076 ;
  LAYER M3 ;
        RECT 17.76 23.588 17.792 23.62 ;
  LAYER M1 ;
        RECT 17.824 23.568 17.856 26.076 ;
  LAYER M3 ;
        RECT 17.824 26.024 17.856 26.056 ;
  LAYER M1 ;
        RECT 17.888 23.568 17.92 26.076 ;
  LAYER M3 ;
        RECT 17.888 23.588 17.92 23.62 ;
  LAYER M1 ;
        RECT 17.952 23.568 17.984 26.076 ;
  LAYER M3 ;
        RECT 17.952 26.024 17.984 26.056 ;
  LAYER M1 ;
        RECT 18.016 23.568 18.048 26.076 ;
  LAYER M3 ;
        RECT 18.016 23.588 18.048 23.62 ;
  LAYER M1 ;
        RECT 18.08 23.568 18.112 26.076 ;
  LAYER M3 ;
        RECT 18.08 26.024 18.112 26.056 ;
  LAYER M1 ;
        RECT 18.144 23.568 18.176 26.076 ;
  LAYER M3 ;
        RECT 18.144 23.588 18.176 23.62 ;
  LAYER M1 ;
        RECT 18.208 23.568 18.24 26.076 ;
  LAYER M3 ;
        RECT 18.208 26.024 18.24 26.056 ;
  LAYER M1 ;
        RECT 18.272 23.568 18.304 26.076 ;
  LAYER M3 ;
        RECT 18.272 23.588 18.304 23.62 ;
  LAYER M1 ;
        RECT 18.336 23.568 18.368 26.076 ;
  LAYER M3 ;
        RECT 18.336 26.024 18.368 26.056 ;
  LAYER M1 ;
        RECT 18.4 23.568 18.432 26.076 ;
  LAYER M3 ;
        RECT 18.4 23.588 18.432 23.62 ;
  LAYER M1 ;
        RECT 18.464 23.568 18.496 26.076 ;
  LAYER M3 ;
        RECT 18.464 26.024 18.496 26.056 ;
  LAYER M1 ;
        RECT 18.528 23.568 18.56 26.076 ;
  LAYER M3 ;
        RECT 18.528 23.588 18.56 23.62 ;
  LAYER M1 ;
        RECT 18.592 23.568 18.624 26.076 ;
  LAYER M3 ;
        RECT 18.592 26.024 18.624 26.056 ;
  LAYER M1 ;
        RECT 18.656 23.568 18.688 26.076 ;
  LAYER M3 ;
        RECT 18.656 23.588 18.688 23.62 ;
  LAYER M1 ;
        RECT 18.72 23.568 18.752 26.076 ;
  LAYER M3 ;
        RECT 18.72 26.024 18.752 26.056 ;
  LAYER M1 ;
        RECT 18.784 23.568 18.816 26.076 ;
  LAYER M3 ;
        RECT 18.784 23.588 18.816 23.62 ;
  LAYER M1 ;
        RECT 18.848 23.568 18.88 26.076 ;
  LAYER M3 ;
        RECT 18.848 26.024 18.88 26.056 ;
  LAYER M1 ;
        RECT 18.912 23.568 18.944 26.076 ;
  LAYER M3 ;
        RECT 18.912 23.588 18.944 23.62 ;
  LAYER M1 ;
        RECT 18.976 23.568 19.008 26.076 ;
  LAYER M3 ;
        RECT 16.608 25.96 16.64 25.992 ;
  LAYER M2 ;
        RECT 18.976 25.896 19.008 25.928 ;
  LAYER M2 ;
        RECT 16.608 25.832 16.64 25.864 ;
  LAYER M2 ;
        RECT 18.976 25.768 19.008 25.8 ;
  LAYER M2 ;
        RECT 16.608 25.704 16.64 25.736 ;
  LAYER M2 ;
        RECT 18.976 25.64 19.008 25.672 ;
  LAYER M2 ;
        RECT 16.608 25.576 16.64 25.608 ;
  LAYER M2 ;
        RECT 18.976 25.512 19.008 25.544 ;
  LAYER M2 ;
        RECT 16.608 25.448 16.64 25.48 ;
  LAYER M2 ;
        RECT 18.976 25.384 19.008 25.416 ;
  LAYER M2 ;
        RECT 16.608 25.32 16.64 25.352 ;
  LAYER M2 ;
        RECT 18.976 25.256 19.008 25.288 ;
  LAYER M2 ;
        RECT 16.608 25.192 16.64 25.224 ;
  LAYER M2 ;
        RECT 18.976 25.128 19.008 25.16 ;
  LAYER M2 ;
        RECT 16.608 25.064 16.64 25.096 ;
  LAYER M2 ;
        RECT 18.976 25 19.008 25.032 ;
  LAYER M2 ;
        RECT 16.608 24.936 16.64 24.968 ;
  LAYER M2 ;
        RECT 18.976 24.872 19.008 24.904 ;
  LAYER M2 ;
        RECT 16.608 24.808 16.64 24.84 ;
  LAYER M2 ;
        RECT 18.976 24.744 19.008 24.776 ;
  LAYER M2 ;
        RECT 16.608 24.68 16.64 24.712 ;
  LAYER M2 ;
        RECT 18.976 24.616 19.008 24.648 ;
  LAYER M2 ;
        RECT 16.608 24.552 16.64 24.584 ;
  LAYER M2 ;
        RECT 18.976 24.488 19.008 24.52 ;
  LAYER M2 ;
        RECT 16.608 24.424 16.64 24.456 ;
  LAYER M2 ;
        RECT 18.976 24.36 19.008 24.392 ;
  LAYER M2 ;
        RECT 16.608 24.296 16.64 24.328 ;
  LAYER M2 ;
        RECT 18.976 24.232 19.008 24.264 ;
  LAYER M2 ;
        RECT 16.608 24.168 16.64 24.2 ;
  LAYER M2 ;
        RECT 18.976 24.104 19.008 24.136 ;
  LAYER M2 ;
        RECT 16.608 24.04 16.64 24.072 ;
  LAYER M2 ;
        RECT 18.976 23.976 19.008 24.008 ;
  LAYER M2 ;
        RECT 16.608 23.912 16.64 23.944 ;
  LAYER M2 ;
        RECT 18.976 23.848 19.008 23.88 ;
  LAYER M2 ;
        RECT 16.608 23.784 16.64 23.816 ;
  LAYER M2 ;
        RECT 18.976 23.72 19.008 23.752 ;
  LAYER M2 ;
        RECT 16.56 23.52 19.056 26.124 ;
  LAYER M1 ;
        RECT 16.608 20.46 16.64 22.968 ;
  LAYER M3 ;
        RECT 16.608 20.48 16.64 20.512 ;
  LAYER M1 ;
        RECT 16.672 20.46 16.704 22.968 ;
  LAYER M3 ;
        RECT 16.672 22.916 16.704 22.948 ;
  LAYER M1 ;
        RECT 16.736 20.46 16.768 22.968 ;
  LAYER M3 ;
        RECT 16.736 20.48 16.768 20.512 ;
  LAYER M1 ;
        RECT 16.8 20.46 16.832 22.968 ;
  LAYER M3 ;
        RECT 16.8 22.916 16.832 22.948 ;
  LAYER M1 ;
        RECT 16.864 20.46 16.896 22.968 ;
  LAYER M3 ;
        RECT 16.864 20.48 16.896 20.512 ;
  LAYER M1 ;
        RECT 16.928 20.46 16.96 22.968 ;
  LAYER M3 ;
        RECT 16.928 22.916 16.96 22.948 ;
  LAYER M1 ;
        RECT 16.992 20.46 17.024 22.968 ;
  LAYER M3 ;
        RECT 16.992 20.48 17.024 20.512 ;
  LAYER M1 ;
        RECT 17.056 20.46 17.088 22.968 ;
  LAYER M3 ;
        RECT 17.056 22.916 17.088 22.948 ;
  LAYER M1 ;
        RECT 17.12 20.46 17.152 22.968 ;
  LAYER M3 ;
        RECT 17.12 20.48 17.152 20.512 ;
  LAYER M1 ;
        RECT 17.184 20.46 17.216 22.968 ;
  LAYER M3 ;
        RECT 17.184 22.916 17.216 22.948 ;
  LAYER M1 ;
        RECT 17.248 20.46 17.28 22.968 ;
  LAYER M3 ;
        RECT 17.248 20.48 17.28 20.512 ;
  LAYER M1 ;
        RECT 17.312 20.46 17.344 22.968 ;
  LAYER M3 ;
        RECT 17.312 22.916 17.344 22.948 ;
  LAYER M1 ;
        RECT 17.376 20.46 17.408 22.968 ;
  LAYER M3 ;
        RECT 17.376 20.48 17.408 20.512 ;
  LAYER M1 ;
        RECT 17.44 20.46 17.472 22.968 ;
  LAYER M3 ;
        RECT 17.44 22.916 17.472 22.948 ;
  LAYER M1 ;
        RECT 17.504 20.46 17.536 22.968 ;
  LAYER M3 ;
        RECT 17.504 20.48 17.536 20.512 ;
  LAYER M1 ;
        RECT 17.568 20.46 17.6 22.968 ;
  LAYER M3 ;
        RECT 17.568 22.916 17.6 22.948 ;
  LAYER M1 ;
        RECT 17.632 20.46 17.664 22.968 ;
  LAYER M3 ;
        RECT 17.632 20.48 17.664 20.512 ;
  LAYER M1 ;
        RECT 17.696 20.46 17.728 22.968 ;
  LAYER M3 ;
        RECT 17.696 22.916 17.728 22.948 ;
  LAYER M1 ;
        RECT 17.76 20.46 17.792 22.968 ;
  LAYER M3 ;
        RECT 17.76 20.48 17.792 20.512 ;
  LAYER M1 ;
        RECT 17.824 20.46 17.856 22.968 ;
  LAYER M3 ;
        RECT 17.824 22.916 17.856 22.948 ;
  LAYER M1 ;
        RECT 17.888 20.46 17.92 22.968 ;
  LAYER M3 ;
        RECT 17.888 20.48 17.92 20.512 ;
  LAYER M1 ;
        RECT 17.952 20.46 17.984 22.968 ;
  LAYER M3 ;
        RECT 17.952 22.916 17.984 22.948 ;
  LAYER M1 ;
        RECT 18.016 20.46 18.048 22.968 ;
  LAYER M3 ;
        RECT 18.016 20.48 18.048 20.512 ;
  LAYER M1 ;
        RECT 18.08 20.46 18.112 22.968 ;
  LAYER M3 ;
        RECT 18.08 22.916 18.112 22.948 ;
  LAYER M1 ;
        RECT 18.144 20.46 18.176 22.968 ;
  LAYER M3 ;
        RECT 18.144 20.48 18.176 20.512 ;
  LAYER M1 ;
        RECT 18.208 20.46 18.24 22.968 ;
  LAYER M3 ;
        RECT 18.208 22.916 18.24 22.948 ;
  LAYER M1 ;
        RECT 18.272 20.46 18.304 22.968 ;
  LAYER M3 ;
        RECT 18.272 20.48 18.304 20.512 ;
  LAYER M1 ;
        RECT 18.336 20.46 18.368 22.968 ;
  LAYER M3 ;
        RECT 18.336 22.916 18.368 22.948 ;
  LAYER M1 ;
        RECT 18.4 20.46 18.432 22.968 ;
  LAYER M3 ;
        RECT 18.4 20.48 18.432 20.512 ;
  LAYER M1 ;
        RECT 18.464 20.46 18.496 22.968 ;
  LAYER M3 ;
        RECT 18.464 22.916 18.496 22.948 ;
  LAYER M1 ;
        RECT 18.528 20.46 18.56 22.968 ;
  LAYER M3 ;
        RECT 18.528 20.48 18.56 20.512 ;
  LAYER M1 ;
        RECT 18.592 20.46 18.624 22.968 ;
  LAYER M3 ;
        RECT 18.592 22.916 18.624 22.948 ;
  LAYER M1 ;
        RECT 18.656 20.46 18.688 22.968 ;
  LAYER M3 ;
        RECT 18.656 20.48 18.688 20.512 ;
  LAYER M1 ;
        RECT 18.72 20.46 18.752 22.968 ;
  LAYER M3 ;
        RECT 18.72 22.916 18.752 22.948 ;
  LAYER M1 ;
        RECT 18.784 20.46 18.816 22.968 ;
  LAYER M3 ;
        RECT 18.784 20.48 18.816 20.512 ;
  LAYER M1 ;
        RECT 18.848 20.46 18.88 22.968 ;
  LAYER M3 ;
        RECT 18.848 22.916 18.88 22.948 ;
  LAYER M1 ;
        RECT 18.912 20.46 18.944 22.968 ;
  LAYER M3 ;
        RECT 18.912 20.48 18.944 20.512 ;
  LAYER M1 ;
        RECT 18.976 20.46 19.008 22.968 ;
  LAYER M3 ;
        RECT 16.608 22.852 16.64 22.884 ;
  LAYER M2 ;
        RECT 18.976 22.788 19.008 22.82 ;
  LAYER M2 ;
        RECT 16.608 22.724 16.64 22.756 ;
  LAYER M2 ;
        RECT 18.976 22.66 19.008 22.692 ;
  LAYER M2 ;
        RECT 16.608 22.596 16.64 22.628 ;
  LAYER M2 ;
        RECT 18.976 22.532 19.008 22.564 ;
  LAYER M2 ;
        RECT 16.608 22.468 16.64 22.5 ;
  LAYER M2 ;
        RECT 18.976 22.404 19.008 22.436 ;
  LAYER M2 ;
        RECT 16.608 22.34 16.64 22.372 ;
  LAYER M2 ;
        RECT 18.976 22.276 19.008 22.308 ;
  LAYER M2 ;
        RECT 16.608 22.212 16.64 22.244 ;
  LAYER M2 ;
        RECT 18.976 22.148 19.008 22.18 ;
  LAYER M2 ;
        RECT 16.608 22.084 16.64 22.116 ;
  LAYER M2 ;
        RECT 18.976 22.02 19.008 22.052 ;
  LAYER M2 ;
        RECT 16.608 21.956 16.64 21.988 ;
  LAYER M2 ;
        RECT 18.976 21.892 19.008 21.924 ;
  LAYER M2 ;
        RECT 16.608 21.828 16.64 21.86 ;
  LAYER M2 ;
        RECT 18.976 21.764 19.008 21.796 ;
  LAYER M2 ;
        RECT 16.608 21.7 16.64 21.732 ;
  LAYER M2 ;
        RECT 18.976 21.636 19.008 21.668 ;
  LAYER M2 ;
        RECT 16.608 21.572 16.64 21.604 ;
  LAYER M2 ;
        RECT 18.976 21.508 19.008 21.54 ;
  LAYER M2 ;
        RECT 16.608 21.444 16.64 21.476 ;
  LAYER M2 ;
        RECT 18.976 21.38 19.008 21.412 ;
  LAYER M2 ;
        RECT 16.608 21.316 16.64 21.348 ;
  LAYER M2 ;
        RECT 18.976 21.252 19.008 21.284 ;
  LAYER M2 ;
        RECT 16.608 21.188 16.64 21.22 ;
  LAYER M2 ;
        RECT 18.976 21.124 19.008 21.156 ;
  LAYER M2 ;
        RECT 16.608 21.06 16.64 21.092 ;
  LAYER M2 ;
        RECT 18.976 20.996 19.008 21.028 ;
  LAYER M2 ;
        RECT 16.608 20.932 16.64 20.964 ;
  LAYER M2 ;
        RECT 18.976 20.868 19.008 20.9 ;
  LAYER M2 ;
        RECT 16.608 20.804 16.64 20.836 ;
  LAYER M2 ;
        RECT 18.976 20.74 19.008 20.772 ;
  LAYER M2 ;
        RECT 16.608 20.676 16.64 20.708 ;
  LAYER M2 ;
        RECT 18.976 20.612 19.008 20.644 ;
  LAYER M2 ;
        RECT 16.56 20.412 19.056 23.016 ;
  LAYER M1 ;
        RECT 19.584 36 19.616 38.508 ;
  LAYER M3 ;
        RECT 19.584 36.02 19.616 36.052 ;
  LAYER M1 ;
        RECT 19.648 36 19.68 38.508 ;
  LAYER M3 ;
        RECT 19.648 38.456 19.68 38.488 ;
  LAYER M1 ;
        RECT 19.712 36 19.744 38.508 ;
  LAYER M3 ;
        RECT 19.712 36.02 19.744 36.052 ;
  LAYER M1 ;
        RECT 19.776 36 19.808 38.508 ;
  LAYER M3 ;
        RECT 19.776 38.456 19.808 38.488 ;
  LAYER M1 ;
        RECT 19.84 36 19.872 38.508 ;
  LAYER M3 ;
        RECT 19.84 36.02 19.872 36.052 ;
  LAYER M1 ;
        RECT 19.904 36 19.936 38.508 ;
  LAYER M3 ;
        RECT 19.904 38.456 19.936 38.488 ;
  LAYER M1 ;
        RECT 19.968 36 20 38.508 ;
  LAYER M3 ;
        RECT 19.968 36.02 20 36.052 ;
  LAYER M1 ;
        RECT 20.032 36 20.064 38.508 ;
  LAYER M3 ;
        RECT 20.032 38.456 20.064 38.488 ;
  LAYER M1 ;
        RECT 20.096 36 20.128 38.508 ;
  LAYER M3 ;
        RECT 20.096 36.02 20.128 36.052 ;
  LAYER M1 ;
        RECT 20.16 36 20.192 38.508 ;
  LAYER M3 ;
        RECT 20.16 38.456 20.192 38.488 ;
  LAYER M1 ;
        RECT 20.224 36 20.256 38.508 ;
  LAYER M3 ;
        RECT 20.224 36.02 20.256 36.052 ;
  LAYER M1 ;
        RECT 20.288 36 20.32 38.508 ;
  LAYER M3 ;
        RECT 20.288 38.456 20.32 38.488 ;
  LAYER M1 ;
        RECT 20.352 36 20.384 38.508 ;
  LAYER M3 ;
        RECT 20.352 36.02 20.384 36.052 ;
  LAYER M1 ;
        RECT 20.416 36 20.448 38.508 ;
  LAYER M3 ;
        RECT 20.416 38.456 20.448 38.488 ;
  LAYER M1 ;
        RECT 20.48 36 20.512 38.508 ;
  LAYER M3 ;
        RECT 20.48 36.02 20.512 36.052 ;
  LAYER M1 ;
        RECT 20.544 36 20.576 38.508 ;
  LAYER M3 ;
        RECT 20.544 38.456 20.576 38.488 ;
  LAYER M1 ;
        RECT 20.608 36 20.64 38.508 ;
  LAYER M3 ;
        RECT 20.608 36.02 20.64 36.052 ;
  LAYER M1 ;
        RECT 20.672 36 20.704 38.508 ;
  LAYER M3 ;
        RECT 20.672 38.456 20.704 38.488 ;
  LAYER M1 ;
        RECT 20.736 36 20.768 38.508 ;
  LAYER M3 ;
        RECT 20.736 36.02 20.768 36.052 ;
  LAYER M1 ;
        RECT 20.8 36 20.832 38.508 ;
  LAYER M3 ;
        RECT 20.8 38.456 20.832 38.488 ;
  LAYER M1 ;
        RECT 20.864 36 20.896 38.508 ;
  LAYER M3 ;
        RECT 20.864 36.02 20.896 36.052 ;
  LAYER M1 ;
        RECT 20.928 36 20.96 38.508 ;
  LAYER M3 ;
        RECT 20.928 38.456 20.96 38.488 ;
  LAYER M1 ;
        RECT 20.992 36 21.024 38.508 ;
  LAYER M3 ;
        RECT 20.992 36.02 21.024 36.052 ;
  LAYER M1 ;
        RECT 21.056 36 21.088 38.508 ;
  LAYER M3 ;
        RECT 21.056 38.456 21.088 38.488 ;
  LAYER M1 ;
        RECT 21.12 36 21.152 38.508 ;
  LAYER M3 ;
        RECT 21.12 36.02 21.152 36.052 ;
  LAYER M1 ;
        RECT 21.184 36 21.216 38.508 ;
  LAYER M3 ;
        RECT 21.184 38.456 21.216 38.488 ;
  LAYER M1 ;
        RECT 21.248 36 21.28 38.508 ;
  LAYER M3 ;
        RECT 21.248 36.02 21.28 36.052 ;
  LAYER M1 ;
        RECT 21.312 36 21.344 38.508 ;
  LAYER M3 ;
        RECT 21.312 38.456 21.344 38.488 ;
  LAYER M1 ;
        RECT 21.376 36 21.408 38.508 ;
  LAYER M3 ;
        RECT 21.376 36.02 21.408 36.052 ;
  LAYER M1 ;
        RECT 21.44 36 21.472 38.508 ;
  LAYER M3 ;
        RECT 21.44 38.456 21.472 38.488 ;
  LAYER M1 ;
        RECT 21.504 36 21.536 38.508 ;
  LAYER M3 ;
        RECT 21.504 36.02 21.536 36.052 ;
  LAYER M1 ;
        RECT 21.568 36 21.6 38.508 ;
  LAYER M3 ;
        RECT 21.568 38.456 21.6 38.488 ;
  LAYER M1 ;
        RECT 21.632 36 21.664 38.508 ;
  LAYER M3 ;
        RECT 21.632 36.02 21.664 36.052 ;
  LAYER M1 ;
        RECT 21.696 36 21.728 38.508 ;
  LAYER M3 ;
        RECT 21.696 38.456 21.728 38.488 ;
  LAYER M1 ;
        RECT 21.76 36 21.792 38.508 ;
  LAYER M3 ;
        RECT 21.76 36.02 21.792 36.052 ;
  LAYER M1 ;
        RECT 21.824 36 21.856 38.508 ;
  LAYER M3 ;
        RECT 21.824 38.456 21.856 38.488 ;
  LAYER M1 ;
        RECT 21.888 36 21.92 38.508 ;
  LAYER M3 ;
        RECT 21.888 36.02 21.92 36.052 ;
  LAYER M1 ;
        RECT 21.952 36 21.984 38.508 ;
  LAYER M3 ;
        RECT 19.584 38.392 19.616 38.424 ;
  LAYER M2 ;
        RECT 21.952 38.328 21.984 38.36 ;
  LAYER M2 ;
        RECT 19.584 38.264 19.616 38.296 ;
  LAYER M2 ;
        RECT 21.952 38.2 21.984 38.232 ;
  LAYER M2 ;
        RECT 19.584 38.136 19.616 38.168 ;
  LAYER M2 ;
        RECT 21.952 38.072 21.984 38.104 ;
  LAYER M2 ;
        RECT 19.584 38.008 19.616 38.04 ;
  LAYER M2 ;
        RECT 21.952 37.944 21.984 37.976 ;
  LAYER M2 ;
        RECT 19.584 37.88 19.616 37.912 ;
  LAYER M2 ;
        RECT 21.952 37.816 21.984 37.848 ;
  LAYER M2 ;
        RECT 19.584 37.752 19.616 37.784 ;
  LAYER M2 ;
        RECT 21.952 37.688 21.984 37.72 ;
  LAYER M2 ;
        RECT 19.584 37.624 19.616 37.656 ;
  LAYER M2 ;
        RECT 21.952 37.56 21.984 37.592 ;
  LAYER M2 ;
        RECT 19.584 37.496 19.616 37.528 ;
  LAYER M2 ;
        RECT 21.952 37.432 21.984 37.464 ;
  LAYER M2 ;
        RECT 19.584 37.368 19.616 37.4 ;
  LAYER M2 ;
        RECT 21.952 37.304 21.984 37.336 ;
  LAYER M2 ;
        RECT 19.584 37.24 19.616 37.272 ;
  LAYER M2 ;
        RECT 21.952 37.176 21.984 37.208 ;
  LAYER M2 ;
        RECT 19.584 37.112 19.616 37.144 ;
  LAYER M2 ;
        RECT 21.952 37.048 21.984 37.08 ;
  LAYER M2 ;
        RECT 19.584 36.984 19.616 37.016 ;
  LAYER M2 ;
        RECT 21.952 36.92 21.984 36.952 ;
  LAYER M2 ;
        RECT 19.584 36.856 19.616 36.888 ;
  LAYER M2 ;
        RECT 21.952 36.792 21.984 36.824 ;
  LAYER M2 ;
        RECT 19.584 36.728 19.616 36.76 ;
  LAYER M2 ;
        RECT 21.952 36.664 21.984 36.696 ;
  LAYER M2 ;
        RECT 19.584 36.6 19.616 36.632 ;
  LAYER M2 ;
        RECT 21.952 36.536 21.984 36.568 ;
  LAYER M2 ;
        RECT 19.584 36.472 19.616 36.504 ;
  LAYER M2 ;
        RECT 21.952 36.408 21.984 36.44 ;
  LAYER M2 ;
        RECT 19.584 36.344 19.616 36.376 ;
  LAYER M2 ;
        RECT 21.952 36.28 21.984 36.312 ;
  LAYER M2 ;
        RECT 19.584 36.216 19.616 36.248 ;
  LAYER M2 ;
        RECT 21.952 36.152 21.984 36.184 ;
  LAYER M2 ;
        RECT 19.536 35.952 22.032 38.556 ;
  LAYER M1 ;
        RECT 19.584 32.892 19.616 35.4 ;
  LAYER M3 ;
        RECT 19.584 32.912 19.616 32.944 ;
  LAYER M1 ;
        RECT 19.648 32.892 19.68 35.4 ;
  LAYER M3 ;
        RECT 19.648 35.348 19.68 35.38 ;
  LAYER M1 ;
        RECT 19.712 32.892 19.744 35.4 ;
  LAYER M3 ;
        RECT 19.712 32.912 19.744 32.944 ;
  LAYER M1 ;
        RECT 19.776 32.892 19.808 35.4 ;
  LAYER M3 ;
        RECT 19.776 35.348 19.808 35.38 ;
  LAYER M1 ;
        RECT 19.84 32.892 19.872 35.4 ;
  LAYER M3 ;
        RECT 19.84 32.912 19.872 32.944 ;
  LAYER M1 ;
        RECT 19.904 32.892 19.936 35.4 ;
  LAYER M3 ;
        RECT 19.904 35.348 19.936 35.38 ;
  LAYER M1 ;
        RECT 19.968 32.892 20 35.4 ;
  LAYER M3 ;
        RECT 19.968 32.912 20 32.944 ;
  LAYER M1 ;
        RECT 20.032 32.892 20.064 35.4 ;
  LAYER M3 ;
        RECT 20.032 35.348 20.064 35.38 ;
  LAYER M1 ;
        RECT 20.096 32.892 20.128 35.4 ;
  LAYER M3 ;
        RECT 20.096 32.912 20.128 32.944 ;
  LAYER M1 ;
        RECT 20.16 32.892 20.192 35.4 ;
  LAYER M3 ;
        RECT 20.16 35.348 20.192 35.38 ;
  LAYER M1 ;
        RECT 20.224 32.892 20.256 35.4 ;
  LAYER M3 ;
        RECT 20.224 32.912 20.256 32.944 ;
  LAYER M1 ;
        RECT 20.288 32.892 20.32 35.4 ;
  LAYER M3 ;
        RECT 20.288 35.348 20.32 35.38 ;
  LAYER M1 ;
        RECT 20.352 32.892 20.384 35.4 ;
  LAYER M3 ;
        RECT 20.352 32.912 20.384 32.944 ;
  LAYER M1 ;
        RECT 20.416 32.892 20.448 35.4 ;
  LAYER M3 ;
        RECT 20.416 35.348 20.448 35.38 ;
  LAYER M1 ;
        RECT 20.48 32.892 20.512 35.4 ;
  LAYER M3 ;
        RECT 20.48 32.912 20.512 32.944 ;
  LAYER M1 ;
        RECT 20.544 32.892 20.576 35.4 ;
  LAYER M3 ;
        RECT 20.544 35.348 20.576 35.38 ;
  LAYER M1 ;
        RECT 20.608 32.892 20.64 35.4 ;
  LAYER M3 ;
        RECT 20.608 32.912 20.64 32.944 ;
  LAYER M1 ;
        RECT 20.672 32.892 20.704 35.4 ;
  LAYER M3 ;
        RECT 20.672 35.348 20.704 35.38 ;
  LAYER M1 ;
        RECT 20.736 32.892 20.768 35.4 ;
  LAYER M3 ;
        RECT 20.736 32.912 20.768 32.944 ;
  LAYER M1 ;
        RECT 20.8 32.892 20.832 35.4 ;
  LAYER M3 ;
        RECT 20.8 35.348 20.832 35.38 ;
  LAYER M1 ;
        RECT 20.864 32.892 20.896 35.4 ;
  LAYER M3 ;
        RECT 20.864 32.912 20.896 32.944 ;
  LAYER M1 ;
        RECT 20.928 32.892 20.96 35.4 ;
  LAYER M3 ;
        RECT 20.928 35.348 20.96 35.38 ;
  LAYER M1 ;
        RECT 20.992 32.892 21.024 35.4 ;
  LAYER M3 ;
        RECT 20.992 32.912 21.024 32.944 ;
  LAYER M1 ;
        RECT 21.056 32.892 21.088 35.4 ;
  LAYER M3 ;
        RECT 21.056 35.348 21.088 35.38 ;
  LAYER M1 ;
        RECT 21.12 32.892 21.152 35.4 ;
  LAYER M3 ;
        RECT 21.12 32.912 21.152 32.944 ;
  LAYER M1 ;
        RECT 21.184 32.892 21.216 35.4 ;
  LAYER M3 ;
        RECT 21.184 35.348 21.216 35.38 ;
  LAYER M1 ;
        RECT 21.248 32.892 21.28 35.4 ;
  LAYER M3 ;
        RECT 21.248 32.912 21.28 32.944 ;
  LAYER M1 ;
        RECT 21.312 32.892 21.344 35.4 ;
  LAYER M3 ;
        RECT 21.312 35.348 21.344 35.38 ;
  LAYER M1 ;
        RECT 21.376 32.892 21.408 35.4 ;
  LAYER M3 ;
        RECT 21.376 32.912 21.408 32.944 ;
  LAYER M1 ;
        RECT 21.44 32.892 21.472 35.4 ;
  LAYER M3 ;
        RECT 21.44 35.348 21.472 35.38 ;
  LAYER M1 ;
        RECT 21.504 32.892 21.536 35.4 ;
  LAYER M3 ;
        RECT 21.504 32.912 21.536 32.944 ;
  LAYER M1 ;
        RECT 21.568 32.892 21.6 35.4 ;
  LAYER M3 ;
        RECT 21.568 35.348 21.6 35.38 ;
  LAYER M1 ;
        RECT 21.632 32.892 21.664 35.4 ;
  LAYER M3 ;
        RECT 21.632 32.912 21.664 32.944 ;
  LAYER M1 ;
        RECT 21.696 32.892 21.728 35.4 ;
  LAYER M3 ;
        RECT 21.696 35.348 21.728 35.38 ;
  LAYER M1 ;
        RECT 21.76 32.892 21.792 35.4 ;
  LAYER M3 ;
        RECT 21.76 32.912 21.792 32.944 ;
  LAYER M1 ;
        RECT 21.824 32.892 21.856 35.4 ;
  LAYER M3 ;
        RECT 21.824 35.348 21.856 35.38 ;
  LAYER M1 ;
        RECT 21.888 32.892 21.92 35.4 ;
  LAYER M3 ;
        RECT 21.888 32.912 21.92 32.944 ;
  LAYER M1 ;
        RECT 21.952 32.892 21.984 35.4 ;
  LAYER M3 ;
        RECT 19.584 35.284 19.616 35.316 ;
  LAYER M2 ;
        RECT 21.952 35.22 21.984 35.252 ;
  LAYER M2 ;
        RECT 19.584 35.156 19.616 35.188 ;
  LAYER M2 ;
        RECT 21.952 35.092 21.984 35.124 ;
  LAYER M2 ;
        RECT 19.584 35.028 19.616 35.06 ;
  LAYER M2 ;
        RECT 21.952 34.964 21.984 34.996 ;
  LAYER M2 ;
        RECT 19.584 34.9 19.616 34.932 ;
  LAYER M2 ;
        RECT 21.952 34.836 21.984 34.868 ;
  LAYER M2 ;
        RECT 19.584 34.772 19.616 34.804 ;
  LAYER M2 ;
        RECT 21.952 34.708 21.984 34.74 ;
  LAYER M2 ;
        RECT 19.584 34.644 19.616 34.676 ;
  LAYER M2 ;
        RECT 21.952 34.58 21.984 34.612 ;
  LAYER M2 ;
        RECT 19.584 34.516 19.616 34.548 ;
  LAYER M2 ;
        RECT 21.952 34.452 21.984 34.484 ;
  LAYER M2 ;
        RECT 19.584 34.388 19.616 34.42 ;
  LAYER M2 ;
        RECT 21.952 34.324 21.984 34.356 ;
  LAYER M2 ;
        RECT 19.584 34.26 19.616 34.292 ;
  LAYER M2 ;
        RECT 21.952 34.196 21.984 34.228 ;
  LAYER M2 ;
        RECT 19.584 34.132 19.616 34.164 ;
  LAYER M2 ;
        RECT 21.952 34.068 21.984 34.1 ;
  LAYER M2 ;
        RECT 19.584 34.004 19.616 34.036 ;
  LAYER M2 ;
        RECT 21.952 33.94 21.984 33.972 ;
  LAYER M2 ;
        RECT 19.584 33.876 19.616 33.908 ;
  LAYER M2 ;
        RECT 21.952 33.812 21.984 33.844 ;
  LAYER M2 ;
        RECT 19.584 33.748 19.616 33.78 ;
  LAYER M2 ;
        RECT 21.952 33.684 21.984 33.716 ;
  LAYER M2 ;
        RECT 19.584 33.62 19.616 33.652 ;
  LAYER M2 ;
        RECT 21.952 33.556 21.984 33.588 ;
  LAYER M2 ;
        RECT 19.584 33.492 19.616 33.524 ;
  LAYER M2 ;
        RECT 21.952 33.428 21.984 33.46 ;
  LAYER M2 ;
        RECT 19.584 33.364 19.616 33.396 ;
  LAYER M2 ;
        RECT 21.952 33.3 21.984 33.332 ;
  LAYER M2 ;
        RECT 19.584 33.236 19.616 33.268 ;
  LAYER M2 ;
        RECT 21.952 33.172 21.984 33.204 ;
  LAYER M2 ;
        RECT 19.584 33.108 19.616 33.14 ;
  LAYER M2 ;
        RECT 21.952 33.044 21.984 33.076 ;
  LAYER M2 ;
        RECT 19.536 32.844 22.032 35.448 ;
  LAYER M1 ;
        RECT 19.584 29.784 19.616 32.292 ;
  LAYER M3 ;
        RECT 19.584 29.804 19.616 29.836 ;
  LAYER M1 ;
        RECT 19.648 29.784 19.68 32.292 ;
  LAYER M3 ;
        RECT 19.648 32.24 19.68 32.272 ;
  LAYER M1 ;
        RECT 19.712 29.784 19.744 32.292 ;
  LAYER M3 ;
        RECT 19.712 29.804 19.744 29.836 ;
  LAYER M1 ;
        RECT 19.776 29.784 19.808 32.292 ;
  LAYER M3 ;
        RECT 19.776 32.24 19.808 32.272 ;
  LAYER M1 ;
        RECT 19.84 29.784 19.872 32.292 ;
  LAYER M3 ;
        RECT 19.84 29.804 19.872 29.836 ;
  LAYER M1 ;
        RECT 19.904 29.784 19.936 32.292 ;
  LAYER M3 ;
        RECT 19.904 32.24 19.936 32.272 ;
  LAYER M1 ;
        RECT 19.968 29.784 20 32.292 ;
  LAYER M3 ;
        RECT 19.968 29.804 20 29.836 ;
  LAYER M1 ;
        RECT 20.032 29.784 20.064 32.292 ;
  LAYER M3 ;
        RECT 20.032 32.24 20.064 32.272 ;
  LAYER M1 ;
        RECT 20.096 29.784 20.128 32.292 ;
  LAYER M3 ;
        RECT 20.096 29.804 20.128 29.836 ;
  LAYER M1 ;
        RECT 20.16 29.784 20.192 32.292 ;
  LAYER M3 ;
        RECT 20.16 32.24 20.192 32.272 ;
  LAYER M1 ;
        RECT 20.224 29.784 20.256 32.292 ;
  LAYER M3 ;
        RECT 20.224 29.804 20.256 29.836 ;
  LAYER M1 ;
        RECT 20.288 29.784 20.32 32.292 ;
  LAYER M3 ;
        RECT 20.288 32.24 20.32 32.272 ;
  LAYER M1 ;
        RECT 20.352 29.784 20.384 32.292 ;
  LAYER M3 ;
        RECT 20.352 29.804 20.384 29.836 ;
  LAYER M1 ;
        RECT 20.416 29.784 20.448 32.292 ;
  LAYER M3 ;
        RECT 20.416 32.24 20.448 32.272 ;
  LAYER M1 ;
        RECT 20.48 29.784 20.512 32.292 ;
  LAYER M3 ;
        RECT 20.48 29.804 20.512 29.836 ;
  LAYER M1 ;
        RECT 20.544 29.784 20.576 32.292 ;
  LAYER M3 ;
        RECT 20.544 32.24 20.576 32.272 ;
  LAYER M1 ;
        RECT 20.608 29.784 20.64 32.292 ;
  LAYER M3 ;
        RECT 20.608 29.804 20.64 29.836 ;
  LAYER M1 ;
        RECT 20.672 29.784 20.704 32.292 ;
  LAYER M3 ;
        RECT 20.672 32.24 20.704 32.272 ;
  LAYER M1 ;
        RECT 20.736 29.784 20.768 32.292 ;
  LAYER M3 ;
        RECT 20.736 29.804 20.768 29.836 ;
  LAYER M1 ;
        RECT 20.8 29.784 20.832 32.292 ;
  LAYER M3 ;
        RECT 20.8 32.24 20.832 32.272 ;
  LAYER M1 ;
        RECT 20.864 29.784 20.896 32.292 ;
  LAYER M3 ;
        RECT 20.864 29.804 20.896 29.836 ;
  LAYER M1 ;
        RECT 20.928 29.784 20.96 32.292 ;
  LAYER M3 ;
        RECT 20.928 32.24 20.96 32.272 ;
  LAYER M1 ;
        RECT 20.992 29.784 21.024 32.292 ;
  LAYER M3 ;
        RECT 20.992 29.804 21.024 29.836 ;
  LAYER M1 ;
        RECT 21.056 29.784 21.088 32.292 ;
  LAYER M3 ;
        RECT 21.056 32.24 21.088 32.272 ;
  LAYER M1 ;
        RECT 21.12 29.784 21.152 32.292 ;
  LAYER M3 ;
        RECT 21.12 29.804 21.152 29.836 ;
  LAYER M1 ;
        RECT 21.184 29.784 21.216 32.292 ;
  LAYER M3 ;
        RECT 21.184 32.24 21.216 32.272 ;
  LAYER M1 ;
        RECT 21.248 29.784 21.28 32.292 ;
  LAYER M3 ;
        RECT 21.248 29.804 21.28 29.836 ;
  LAYER M1 ;
        RECT 21.312 29.784 21.344 32.292 ;
  LAYER M3 ;
        RECT 21.312 32.24 21.344 32.272 ;
  LAYER M1 ;
        RECT 21.376 29.784 21.408 32.292 ;
  LAYER M3 ;
        RECT 21.376 29.804 21.408 29.836 ;
  LAYER M1 ;
        RECT 21.44 29.784 21.472 32.292 ;
  LAYER M3 ;
        RECT 21.44 32.24 21.472 32.272 ;
  LAYER M1 ;
        RECT 21.504 29.784 21.536 32.292 ;
  LAYER M3 ;
        RECT 21.504 29.804 21.536 29.836 ;
  LAYER M1 ;
        RECT 21.568 29.784 21.6 32.292 ;
  LAYER M3 ;
        RECT 21.568 32.24 21.6 32.272 ;
  LAYER M1 ;
        RECT 21.632 29.784 21.664 32.292 ;
  LAYER M3 ;
        RECT 21.632 29.804 21.664 29.836 ;
  LAYER M1 ;
        RECT 21.696 29.784 21.728 32.292 ;
  LAYER M3 ;
        RECT 21.696 32.24 21.728 32.272 ;
  LAYER M1 ;
        RECT 21.76 29.784 21.792 32.292 ;
  LAYER M3 ;
        RECT 21.76 29.804 21.792 29.836 ;
  LAYER M1 ;
        RECT 21.824 29.784 21.856 32.292 ;
  LAYER M3 ;
        RECT 21.824 32.24 21.856 32.272 ;
  LAYER M1 ;
        RECT 21.888 29.784 21.92 32.292 ;
  LAYER M3 ;
        RECT 21.888 29.804 21.92 29.836 ;
  LAYER M1 ;
        RECT 21.952 29.784 21.984 32.292 ;
  LAYER M3 ;
        RECT 19.584 32.176 19.616 32.208 ;
  LAYER M2 ;
        RECT 21.952 32.112 21.984 32.144 ;
  LAYER M2 ;
        RECT 19.584 32.048 19.616 32.08 ;
  LAYER M2 ;
        RECT 21.952 31.984 21.984 32.016 ;
  LAYER M2 ;
        RECT 19.584 31.92 19.616 31.952 ;
  LAYER M2 ;
        RECT 21.952 31.856 21.984 31.888 ;
  LAYER M2 ;
        RECT 19.584 31.792 19.616 31.824 ;
  LAYER M2 ;
        RECT 21.952 31.728 21.984 31.76 ;
  LAYER M2 ;
        RECT 19.584 31.664 19.616 31.696 ;
  LAYER M2 ;
        RECT 21.952 31.6 21.984 31.632 ;
  LAYER M2 ;
        RECT 19.584 31.536 19.616 31.568 ;
  LAYER M2 ;
        RECT 21.952 31.472 21.984 31.504 ;
  LAYER M2 ;
        RECT 19.584 31.408 19.616 31.44 ;
  LAYER M2 ;
        RECT 21.952 31.344 21.984 31.376 ;
  LAYER M2 ;
        RECT 19.584 31.28 19.616 31.312 ;
  LAYER M2 ;
        RECT 21.952 31.216 21.984 31.248 ;
  LAYER M2 ;
        RECT 19.584 31.152 19.616 31.184 ;
  LAYER M2 ;
        RECT 21.952 31.088 21.984 31.12 ;
  LAYER M2 ;
        RECT 19.584 31.024 19.616 31.056 ;
  LAYER M2 ;
        RECT 21.952 30.96 21.984 30.992 ;
  LAYER M2 ;
        RECT 19.584 30.896 19.616 30.928 ;
  LAYER M2 ;
        RECT 21.952 30.832 21.984 30.864 ;
  LAYER M2 ;
        RECT 19.584 30.768 19.616 30.8 ;
  LAYER M2 ;
        RECT 21.952 30.704 21.984 30.736 ;
  LAYER M2 ;
        RECT 19.584 30.64 19.616 30.672 ;
  LAYER M2 ;
        RECT 21.952 30.576 21.984 30.608 ;
  LAYER M2 ;
        RECT 19.584 30.512 19.616 30.544 ;
  LAYER M2 ;
        RECT 21.952 30.448 21.984 30.48 ;
  LAYER M2 ;
        RECT 19.584 30.384 19.616 30.416 ;
  LAYER M2 ;
        RECT 21.952 30.32 21.984 30.352 ;
  LAYER M2 ;
        RECT 19.584 30.256 19.616 30.288 ;
  LAYER M2 ;
        RECT 21.952 30.192 21.984 30.224 ;
  LAYER M2 ;
        RECT 19.584 30.128 19.616 30.16 ;
  LAYER M2 ;
        RECT 21.952 30.064 21.984 30.096 ;
  LAYER M2 ;
        RECT 19.584 30 19.616 30.032 ;
  LAYER M2 ;
        RECT 21.952 29.936 21.984 29.968 ;
  LAYER M2 ;
        RECT 19.536 29.736 22.032 32.34 ;
  LAYER M1 ;
        RECT 19.584 26.676 19.616 29.184 ;
  LAYER M3 ;
        RECT 19.584 26.696 19.616 26.728 ;
  LAYER M1 ;
        RECT 19.648 26.676 19.68 29.184 ;
  LAYER M3 ;
        RECT 19.648 29.132 19.68 29.164 ;
  LAYER M1 ;
        RECT 19.712 26.676 19.744 29.184 ;
  LAYER M3 ;
        RECT 19.712 26.696 19.744 26.728 ;
  LAYER M1 ;
        RECT 19.776 26.676 19.808 29.184 ;
  LAYER M3 ;
        RECT 19.776 29.132 19.808 29.164 ;
  LAYER M1 ;
        RECT 19.84 26.676 19.872 29.184 ;
  LAYER M3 ;
        RECT 19.84 26.696 19.872 26.728 ;
  LAYER M1 ;
        RECT 19.904 26.676 19.936 29.184 ;
  LAYER M3 ;
        RECT 19.904 29.132 19.936 29.164 ;
  LAYER M1 ;
        RECT 19.968 26.676 20 29.184 ;
  LAYER M3 ;
        RECT 19.968 26.696 20 26.728 ;
  LAYER M1 ;
        RECT 20.032 26.676 20.064 29.184 ;
  LAYER M3 ;
        RECT 20.032 29.132 20.064 29.164 ;
  LAYER M1 ;
        RECT 20.096 26.676 20.128 29.184 ;
  LAYER M3 ;
        RECT 20.096 26.696 20.128 26.728 ;
  LAYER M1 ;
        RECT 20.16 26.676 20.192 29.184 ;
  LAYER M3 ;
        RECT 20.16 29.132 20.192 29.164 ;
  LAYER M1 ;
        RECT 20.224 26.676 20.256 29.184 ;
  LAYER M3 ;
        RECT 20.224 26.696 20.256 26.728 ;
  LAYER M1 ;
        RECT 20.288 26.676 20.32 29.184 ;
  LAYER M3 ;
        RECT 20.288 29.132 20.32 29.164 ;
  LAYER M1 ;
        RECT 20.352 26.676 20.384 29.184 ;
  LAYER M3 ;
        RECT 20.352 26.696 20.384 26.728 ;
  LAYER M1 ;
        RECT 20.416 26.676 20.448 29.184 ;
  LAYER M3 ;
        RECT 20.416 29.132 20.448 29.164 ;
  LAYER M1 ;
        RECT 20.48 26.676 20.512 29.184 ;
  LAYER M3 ;
        RECT 20.48 26.696 20.512 26.728 ;
  LAYER M1 ;
        RECT 20.544 26.676 20.576 29.184 ;
  LAYER M3 ;
        RECT 20.544 29.132 20.576 29.164 ;
  LAYER M1 ;
        RECT 20.608 26.676 20.64 29.184 ;
  LAYER M3 ;
        RECT 20.608 26.696 20.64 26.728 ;
  LAYER M1 ;
        RECT 20.672 26.676 20.704 29.184 ;
  LAYER M3 ;
        RECT 20.672 29.132 20.704 29.164 ;
  LAYER M1 ;
        RECT 20.736 26.676 20.768 29.184 ;
  LAYER M3 ;
        RECT 20.736 26.696 20.768 26.728 ;
  LAYER M1 ;
        RECT 20.8 26.676 20.832 29.184 ;
  LAYER M3 ;
        RECT 20.8 29.132 20.832 29.164 ;
  LAYER M1 ;
        RECT 20.864 26.676 20.896 29.184 ;
  LAYER M3 ;
        RECT 20.864 26.696 20.896 26.728 ;
  LAYER M1 ;
        RECT 20.928 26.676 20.96 29.184 ;
  LAYER M3 ;
        RECT 20.928 29.132 20.96 29.164 ;
  LAYER M1 ;
        RECT 20.992 26.676 21.024 29.184 ;
  LAYER M3 ;
        RECT 20.992 26.696 21.024 26.728 ;
  LAYER M1 ;
        RECT 21.056 26.676 21.088 29.184 ;
  LAYER M3 ;
        RECT 21.056 29.132 21.088 29.164 ;
  LAYER M1 ;
        RECT 21.12 26.676 21.152 29.184 ;
  LAYER M3 ;
        RECT 21.12 26.696 21.152 26.728 ;
  LAYER M1 ;
        RECT 21.184 26.676 21.216 29.184 ;
  LAYER M3 ;
        RECT 21.184 29.132 21.216 29.164 ;
  LAYER M1 ;
        RECT 21.248 26.676 21.28 29.184 ;
  LAYER M3 ;
        RECT 21.248 26.696 21.28 26.728 ;
  LAYER M1 ;
        RECT 21.312 26.676 21.344 29.184 ;
  LAYER M3 ;
        RECT 21.312 29.132 21.344 29.164 ;
  LAYER M1 ;
        RECT 21.376 26.676 21.408 29.184 ;
  LAYER M3 ;
        RECT 21.376 26.696 21.408 26.728 ;
  LAYER M1 ;
        RECT 21.44 26.676 21.472 29.184 ;
  LAYER M3 ;
        RECT 21.44 29.132 21.472 29.164 ;
  LAYER M1 ;
        RECT 21.504 26.676 21.536 29.184 ;
  LAYER M3 ;
        RECT 21.504 26.696 21.536 26.728 ;
  LAYER M1 ;
        RECT 21.568 26.676 21.6 29.184 ;
  LAYER M3 ;
        RECT 21.568 29.132 21.6 29.164 ;
  LAYER M1 ;
        RECT 21.632 26.676 21.664 29.184 ;
  LAYER M3 ;
        RECT 21.632 26.696 21.664 26.728 ;
  LAYER M1 ;
        RECT 21.696 26.676 21.728 29.184 ;
  LAYER M3 ;
        RECT 21.696 29.132 21.728 29.164 ;
  LAYER M1 ;
        RECT 21.76 26.676 21.792 29.184 ;
  LAYER M3 ;
        RECT 21.76 26.696 21.792 26.728 ;
  LAYER M1 ;
        RECT 21.824 26.676 21.856 29.184 ;
  LAYER M3 ;
        RECT 21.824 29.132 21.856 29.164 ;
  LAYER M1 ;
        RECT 21.888 26.676 21.92 29.184 ;
  LAYER M3 ;
        RECT 21.888 26.696 21.92 26.728 ;
  LAYER M1 ;
        RECT 21.952 26.676 21.984 29.184 ;
  LAYER M3 ;
        RECT 19.584 29.068 19.616 29.1 ;
  LAYER M2 ;
        RECT 21.952 29.004 21.984 29.036 ;
  LAYER M2 ;
        RECT 19.584 28.94 19.616 28.972 ;
  LAYER M2 ;
        RECT 21.952 28.876 21.984 28.908 ;
  LAYER M2 ;
        RECT 19.584 28.812 19.616 28.844 ;
  LAYER M2 ;
        RECT 21.952 28.748 21.984 28.78 ;
  LAYER M2 ;
        RECT 19.584 28.684 19.616 28.716 ;
  LAYER M2 ;
        RECT 21.952 28.62 21.984 28.652 ;
  LAYER M2 ;
        RECT 19.584 28.556 19.616 28.588 ;
  LAYER M2 ;
        RECT 21.952 28.492 21.984 28.524 ;
  LAYER M2 ;
        RECT 19.584 28.428 19.616 28.46 ;
  LAYER M2 ;
        RECT 21.952 28.364 21.984 28.396 ;
  LAYER M2 ;
        RECT 19.584 28.3 19.616 28.332 ;
  LAYER M2 ;
        RECT 21.952 28.236 21.984 28.268 ;
  LAYER M2 ;
        RECT 19.584 28.172 19.616 28.204 ;
  LAYER M2 ;
        RECT 21.952 28.108 21.984 28.14 ;
  LAYER M2 ;
        RECT 19.584 28.044 19.616 28.076 ;
  LAYER M2 ;
        RECT 21.952 27.98 21.984 28.012 ;
  LAYER M2 ;
        RECT 19.584 27.916 19.616 27.948 ;
  LAYER M2 ;
        RECT 21.952 27.852 21.984 27.884 ;
  LAYER M2 ;
        RECT 19.584 27.788 19.616 27.82 ;
  LAYER M2 ;
        RECT 21.952 27.724 21.984 27.756 ;
  LAYER M2 ;
        RECT 19.584 27.66 19.616 27.692 ;
  LAYER M2 ;
        RECT 21.952 27.596 21.984 27.628 ;
  LAYER M2 ;
        RECT 19.584 27.532 19.616 27.564 ;
  LAYER M2 ;
        RECT 21.952 27.468 21.984 27.5 ;
  LAYER M2 ;
        RECT 19.584 27.404 19.616 27.436 ;
  LAYER M2 ;
        RECT 21.952 27.34 21.984 27.372 ;
  LAYER M2 ;
        RECT 19.584 27.276 19.616 27.308 ;
  LAYER M2 ;
        RECT 21.952 27.212 21.984 27.244 ;
  LAYER M2 ;
        RECT 19.584 27.148 19.616 27.18 ;
  LAYER M2 ;
        RECT 21.952 27.084 21.984 27.116 ;
  LAYER M2 ;
        RECT 19.584 27.02 19.616 27.052 ;
  LAYER M2 ;
        RECT 21.952 26.956 21.984 26.988 ;
  LAYER M2 ;
        RECT 19.584 26.892 19.616 26.924 ;
  LAYER M2 ;
        RECT 21.952 26.828 21.984 26.86 ;
  LAYER M2 ;
        RECT 19.536 26.628 22.032 29.232 ;
  LAYER M1 ;
        RECT 19.584 23.568 19.616 26.076 ;
  LAYER M3 ;
        RECT 19.584 23.588 19.616 23.62 ;
  LAYER M1 ;
        RECT 19.648 23.568 19.68 26.076 ;
  LAYER M3 ;
        RECT 19.648 26.024 19.68 26.056 ;
  LAYER M1 ;
        RECT 19.712 23.568 19.744 26.076 ;
  LAYER M3 ;
        RECT 19.712 23.588 19.744 23.62 ;
  LAYER M1 ;
        RECT 19.776 23.568 19.808 26.076 ;
  LAYER M3 ;
        RECT 19.776 26.024 19.808 26.056 ;
  LAYER M1 ;
        RECT 19.84 23.568 19.872 26.076 ;
  LAYER M3 ;
        RECT 19.84 23.588 19.872 23.62 ;
  LAYER M1 ;
        RECT 19.904 23.568 19.936 26.076 ;
  LAYER M3 ;
        RECT 19.904 26.024 19.936 26.056 ;
  LAYER M1 ;
        RECT 19.968 23.568 20 26.076 ;
  LAYER M3 ;
        RECT 19.968 23.588 20 23.62 ;
  LAYER M1 ;
        RECT 20.032 23.568 20.064 26.076 ;
  LAYER M3 ;
        RECT 20.032 26.024 20.064 26.056 ;
  LAYER M1 ;
        RECT 20.096 23.568 20.128 26.076 ;
  LAYER M3 ;
        RECT 20.096 23.588 20.128 23.62 ;
  LAYER M1 ;
        RECT 20.16 23.568 20.192 26.076 ;
  LAYER M3 ;
        RECT 20.16 26.024 20.192 26.056 ;
  LAYER M1 ;
        RECT 20.224 23.568 20.256 26.076 ;
  LAYER M3 ;
        RECT 20.224 23.588 20.256 23.62 ;
  LAYER M1 ;
        RECT 20.288 23.568 20.32 26.076 ;
  LAYER M3 ;
        RECT 20.288 26.024 20.32 26.056 ;
  LAYER M1 ;
        RECT 20.352 23.568 20.384 26.076 ;
  LAYER M3 ;
        RECT 20.352 23.588 20.384 23.62 ;
  LAYER M1 ;
        RECT 20.416 23.568 20.448 26.076 ;
  LAYER M3 ;
        RECT 20.416 26.024 20.448 26.056 ;
  LAYER M1 ;
        RECT 20.48 23.568 20.512 26.076 ;
  LAYER M3 ;
        RECT 20.48 23.588 20.512 23.62 ;
  LAYER M1 ;
        RECT 20.544 23.568 20.576 26.076 ;
  LAYER M3 ;
        RECT 20.544 26.024 20.576 26.056 ;
  LAYER M1 ;
        RECT 20.608 23.568 20.64 26.076 ;
  LAYER M3 ;
        RECT 20.608 23.588 20.64 23.62 ;
  LAYER M1 ;
        RECT 20.672 23.568 20.704 26.076 ;
  LAYER M3 ;
        RECT 20.672 26.024 20.704 26.056 ;
  LAYER M1 ;
        RECT 20.736 23.568 20.768 26.076 ;
  LAYER M3 ;
        RECT 20.736 23.588 20.768 23.62 ;
  LAYER M1 ;
        RECT 20.8 23.568 20.832 26.076 ;
  LAYER M3 ;
        RECT 20.8 26.024 20.832 26.056 ;
  LAYER M1 ;
        RECT 20.864 23.568 20.896 26.076 ;
  LAYER M3 ;
        RECT 20.864 23.588 20.896 23.62 ;
  LAYER M1 ;
        RECT 20.928 23.568 20.96 26.076 ;
  LAYER M3 ;
        RECT 20.928 26.024 20.96 26.056 ;
  LAYER M1 ;
        RECT 20.992 23.568 21.024 26.076 ;
  LAYER M3 ;
        RECT 20.992 23.588 21.024 23.62 ;
  LAYER M1 ;
        RECT 21.056 23.568 21.088 26.076 ;
  LAYER M3 ;
        RECT 21.056 26.024 21.088 26.056 ;
  LAYER M1 ;
        RECT 21.12 23.568 21.152 26.076 ;
  LAYER M3 ;
        RECT 21.12 23.588 21.152 23.62 ;
  LAYER M1 ;
        RECT 21.184 23.568 21.216 26.076 ;
  LAYER M3 ;
        RECT 21.184 26.024 21.216 26.056 ;
  LAYER M1 ;
        RECT 21.248 23.568 21.28 26.076 ;
  LAYER M3 ;
        RECT 21.248 23.588 21.28 23.62 ;
  LAYER M1 ;
        RECT 21.312 23.568 21.344 26.076 ;
  LAYER M3 ;
        RECT 21.312 26.024 21.344 26.056 ;
  LAYER M1 ;
        RECT 21.376 23.568 21.408 26.076 ;
  LAYER M3 ;
        RECT 21.376 23.588 21.408 23.62 ;
  LAYER M1 ;
        RECT 21.44 23.568 21.472 26.076 ;
  LAYER M3 ;
        RECT 21.44 26.024 21.472 26.056 ;
  LAYER M1 ;
        RECT 21.504 23.568 21.536 26.076 ;
  LAYER M3 ;
        RECT 21.504 23.588 21.536 23.62 ;
  LAYER M1 ;
        RECT 21.568 23.568 21.6 26.076 ;
  LAYER M3 ;
        RECT 21.568 26.024 21.6 26.056 ;
  LAYER M1 ;
        RECT 21.632 23.568 21.664 26.076 ;
  LAYER M3 ;
        RECT 21.632 23.588 21.664 23.62 ;
  LAYER M1 ;
        RECT 21.696 23.568 21.728 26.076 ;
  LAYER M3 ;
        RECT 21.696 26.024 21.728 26.056 ;
  LAYER M1 ;
        RECT 21.76 23.568 21.792 26.076 ;
  LAYER M3 ;
        RECT 21.76 23.588 21.792 23.62 ;
  LAYER M1 ;
        RECT 21.824 23.568 21.856 26.076 ;
  LAYER M3 ;
        RECT 21.824 26.024 21.856 26.056 ;
  LAYER M1 ;
        RECT 21.888 23.568 21.92 26.076 ;
  LAYER M3 ;
        RECT 21.888 23.588 21.92 23.62 ;
  LAYER M1 ;
        RECT 21.952 23.568 21.984 26.076 ;
  LAYER M3 ;
        RECT 19.584 25.96 19.616 25.992 ;
  LAYER M2 ;
        RECT 21.952 25.896 21.984 25.928 ;
  LAYER M2 ;
        RECT 19.584 25.832 19.616 25.864 ;
  LAYER M2 ;
        RECT 21.952 25.768 21.984 25.8 ;
  LAYER M2 ;
        RECT 19.584 25.704 19.616 25.736 ;
  LAYER M2 ;
        RECT 21.952 25.64 21.984 25.672 ;
  LAYER M2 ;
        RECT 19.584 25.576 19.616 25.608 ;
  LAYER M2 ;
        RECT 21.952 25.512 21.984 25.544 ;
  LAYER M2 ;
        RECT 19.584 25.448 19.616 25.48 ;
  LAYER M2 ;
        RECT 21.952 25.384 21.984 25.416 ;
  LAYER M2 ;
        RECT 19.584 25.32 19.616 25.352 ;
  LAYER M2 ;
        RECT 21.952 25.256 21.984 25.288 ;
  LAYER M2 ;
        RECT 19.584 25.192 19.616 25.224 ;
  LAYER M2 ;
        RECT 21.952 25.128 21.984 25.16 ;
  LAYER M2 ;
        RECT 19.584 25.064 19.616 25.096 ;
  LAYER M2 ;
        RECT 21.952 25 21.984 25.032 ;
  LAYER M2 ;
        RECT 19.584 24.936 19.616 24.968 ;
  LAYER M2 ;
        RECT 21.952 24.872 21.984 24.904 ;
  LAYER M2 ;
        RECT 19.584 24.808 19.616 24.84 ;
  LAYER M2 ;
        RECT 21.952 24.744 21.984 24.776 ;
  LAYER M2 ;
        RECT 19.584 24.68 19.616 24.712 ;
  LAYER M2 ;
        RECT 21.952 24.616 21.984 24.648 ;
  LAYER M2 ;
        RECT 19.584 24.552 19.616 24.584 ;
  LAYER M2 ;
        RECT 21.952 24.488 21.984 24.52 ;
  LAYER M2 ;
        RECT 19.584 24.424 19.616 24.456 ;
  LAYER M2 ;
        RECT 21.952 24.36 21.984 24.392 ;
  LAYER M2 ;
        RECT 19.584 24.296 19.616 24.328 ;
  LAYER M2 ;
        RECT 21.952 24.232 21.984 24.264 ;
  LAYER M2 ;
        RECT 19.584 24.168 19.616 24.2 ;
  LAYER M2 ;
        RECT 21.952 24.104 21.984 24.136 ;
  LAYER M2 ;
        RECT 19.584 24.04 19.616 24.072 ;
  LAYER M2 ;
        RECT 21.952 23.976 21.984 24.008 ;
  LAYER M2 ;
        RECT 19.584 23.912 19.616 23.944 ;
  LAYER M2 ;
        RECT 21.952 23.848 21.984 23.88 ;
  LAYER M2 ;
        RECT 19.584 23.784 19.616 23.816 ;
  LAYER M2 ;
        RECT 21.952 23.72 21.984 23.752 ;
  LAYER M2 ;
        RECT 19.536 23.52 22.032 26.124 ;
  LAYER M1 ;
        RECT 19.584 20.46 19.616 22.968 ;
  LAYER M3 ;
        RECT 19.584 20.48 19.616 20.512 ;
  LAYER M1 ;
        RECT 19.648 20.46 19.68 22.968 ;
  LAYER M3 ;
        RECT 19.648 22.916 19.68 22.948 ;
  LAYER M1 ;
        RECT 19.712 20.46 19.744 22.968 ;
  LAYER M3 ;
        RECT 19.712 20.48 19.744 20.512 ;
  LAYER M1 ;
        RECT 19.776 20.46 19.808 22.968 ;
  LAYER M3 ;
        RECT 19.776 22.916 19.808 22.948 ;
  LAYER M1 ;
        RECT 19.84 20.46 19.872 22.968 ;
  LAYER M3 ;
        RECT 19.84 20.48 19.872 20.512 ;
  LAYER M1 ;
        RECT 19.904 20.46 19.936 22.968 ;
  LAYER M3 ;
        RECT 19.904 22.916 19.936 22.948 ;
  LAYER M1 ;
        RECT 19.968 20.46 20 22.968 ;
  LAYER M3 ;
        RECT 19.968 20.48 20 20.512 ;
  LAYER M1 ;
        RECT 20.032 20.46 20.064 22.968 ;
  LAYER M3 ;
        RECT 20.032 22.916 20.064 22.948 ;
  LAYER M1 ;
        RECT 20.096 20.46 20.128 22.968 ;
  LAYER M3 ;
        RECT 20.096 20.48 20.128 20.512 ;
  LAYER M1 ;
        RECT 20.16 20.46 20.192 22.968 ;
  LAYER M3 ;
        RECT 20.16 22.916 20.192 22.948 ;
  LAYER M1 ;
        RECT 20.224 20.46 20.256 22.968 ;
  LAYER M3 ;
        RECT 20.224 20.48 20.256 20.512 ;
  LAYER M1 ;
        RECT 20.288 20.46 20.32 22.968 ;
  LAYER M3 ;
        RECT 20.288 22.916 20.32 22.948 ;
  LAYER M1 ;
        RECT 20.352 20.46 20.384 22.968 ;
  LAYER M3 ;
        RECT 20.352 20.48 20.384 20.512 ;
  LAYER M1 ;
        RECT 20.416 20.46 20.448 22.968 ;
  LAYER M3 ;
        RECT 20.416 22.916 20.448 22.948 ;
  LAYER M1 ;
        RECT 20.48 20.46 20.512 22.968 ;
  LAYER M3 ;
        RECT 20.48 20.48 20.512 20.512 ;
  LAYER M1 ;
        RECT 20.544 20.46 20.576 22.968 ;
  LAYER M3 ;
        RECT 20.544 22.916 20.576 22.948 ;
  LAYER M1 ;
        RECT 20.608 20.46 20.64 22.968 ;
  LAYER M3 ;
        RECT 20.608 20.48 20.64 20.512 ;
  LAYER M1 ;
        RECT 20.672 20.46 20.704 22.968 ;
  LAYER M3 ;
        RECT 20.672 22.916 20.704 22.948 ;
  LAYER M1 ;
        RECT 20.736 20.46 20.768 22.968 ;
  LAYER M3 ;
        RECT 20.736 20.48 20.768 20.512 ;
  LAYER M1 ;
        RECT 20.8 20.46 20.832 22.968 ;
  LAYER M3 ;
        RECT 20.8 22.916 20.832 22.948 ;
  LAYER M1 ;
        RECT 20.864 20.46 20.896 22.968 ;
  LAYER M3 ;
        RECT 20.864 20.48 20.896 20.512 ;
  LAYER M1 ;
        RECT 20.928 20.46 20.96 22.968 ;
  LAYER M3 ;
        RECT 20.928 22.916 20.96 22.948 ;
  LAYER M1 ;
        RECT 20.992 20.46 21.024 22.968 ;
  LAYER M3 ;
        RECT 20.992 20.48 21.024 20.512 ;
  LAYER M1 ;
        RECT 21.056 20.46 21.088 22.968 ;
  LAYER M3 ;
        RECT 21.056 22.916 21.088 22.948 ;
  LAYER M1 ;
        RECT 21.12 20.46 21.152 22.968 ;
  LAYER M3 ;
        RECT 21.12 20.48 21.152 20.512 ;
  LAYER M1 ;
        RECT 21.184 20.46 21.216 22.968 ;
  LAYER M3 ;
        RECT 21.184 22.916 21.216 22.948 ;
  LAYER M1 ;
        RECT 21.248 20.46 21.28 22.968 ;
  LAYER M3 ;
        RECT 21.248 20.48 21.28 20.512 ;
  LAYER M1 ;
        RECT 21.312 20.46 21.344 22.968 ;
  LAYER M3 ;
        RECT 21.312 22.916 21.344 22.948 ;
  LAYER M1 ;
        RECT 21.376 20.46 21.408 22.968 ;
  LAYER M3 ;
        RECT 21.376 20.48 21.408 20.512 ;
  LAYER M1 ;
        RECT 21.44 20.46 21.472 22.968 ;
  LAYER M3 ;
        RECT 21.44 22.916 21.472 22.948 ;
  LAYER M1 ;
        RECT 21.504 20.46 21.536 22.968 ;
  LAYER M3 ;
        RECT 21.504 20.48 21.536 20.512 ;
  LAYER M1 ;
        RECT 21.568 20.46 21.6 22.968 ;
  LAYER M3 ;
        RECT 21.568 22.916 21.6 22.948 ;
  LAYER M1 ;
        RECT 21.632 20.46 21.664 22.968 ;
  LAYER M3 ;
        RECT 21.632 20.48 21.664 20.512 ;
  LAYER M1 ;
        RECT 21.696 20.46 21.728 22.968 ;
  LAYER M3 ;
        RECT 21.696 22.916 21.728 22.948 ;
  LAYER M1 ;
        RECT 21.76 20.46 21.792 22.968 ;
  LAYER M3 ;
        RECT 21.76 20.48 21.792 20.512 ;
  LAYER M1 ;
        RECT 21.824 20.46 21.856 22.968 ;
  LAYER M3 ;
        RECT 21.824 22.916 21.856 22.948 ;
  LAYER M1 ;
        RECT 21.888 20.46 21.92 22.968 ;
  LAYER M3 ;
        RECT 21.888 20.48 21.92 20.512 ;
  LAYER M1 ;
        RECT 21.952 20.46 21.984 22.968 ;
  LAYER M3 ;
        RECT 19.584 22.852 19.616 22.884 ;
  LAYER M2 ;
        RECT 21.952 22.788 21.984 22.82 ;
  LAYER M2 ;
        RECT 19.584 22.724 19.616 22.756 ;
  LAYER M2 ;
        RECT 21.952 22.66 21.984 22.692 ;
  LAYER M2 ;
        RECT 19.584 22.596 19.616 22.628 ;
  LAYER M2 ;
        RECT 21.952 22.532 21.984 22.564 ;
  LAYER M2 ;
        RECT 19.584 22.468 19.616 22.5 ;
  LAYER M2 ;
        RECT 21.952 22.404 21.984 22.436 ;
  LAYER M2 ;
        RECT 19.584 22.34 19.616 22.372 ;
  LAYER M2 ;
        RECT 21.952 22.276 21.984 22.308 ;
  LAYER M2 ;
        RECT 19.584 22.212 19.616 22.244 ;
  LAYER M2 ;
        RECT 21.952 22.148 21.984 22.18 ;
  LAYER M2 ;
        RECT 19.584 22.084 19.616 22.116 ;
  LAYER M2 ;
        RECT 21.952 22.02 21.984 22.052 ;
  LAYER M2 ;
        RECT 19.584 21.956 19.616 21.988 ;
  LAYER M2 ;
        RECT 21.952 21.892 21.984 21.924 ;
  LAYER M2 ;
        RECT 19.584 21.828 19.616 21.86 ;
  LAYER M2 ;
        RECT 21.952 21.764 21.984 21.796 ;
  LAYER M2 ;
        RECT 19.584 21.7 19.616 21.732 ;
  LAYER M2 ;
        RECT 21.952 21.636 21.984 21.668 ;
  LAYER M2 ;
        RECT 19.584 21.572 19.616 21.604 ;
  LAYER M2 ;
        RECT 21.952 21.508 21.984 21.54 ;
  LAYER M2 ;
        RECT 19.584 21.444 19.616 21.476 ;
  LAYER M2 ;
        RECT 21.952 21.38 21.984 21.412 ;
  LAYER M2 ;
        RECT 19.584 21.316 19.616 21.348 ;
  LAYER M2 ;
        RECT 21.952 21.252 21.984 21.284 ;
  LAYER M2 ;
        RECT 19.584 21.188 19.616 21.22 ;
  LAYER M2 ;
        RECT 21.952 21.124 21.984 21.156 ;
  LAYER M2 ;
        RECT 19.584 21.06 19.616 21.092 ;
  LAYER M2 ;
        RECT 21.952 20.996 21.984 21.028 ;
  LAYER M2 ;
        RECT 19.584 20.932 19.616 20.964 ;
  LAYER M2 ;
        RECT 21.952 20.868 21.984 20.9 ;
  LAYER M2 ;
        RECT 19.584 20.804 19.616 20.836 ;
  LAYER M2 ;
        RECT 21.952 20.74 21.984 20.772 ;
  LAYER M2 ;
        RECT 19.584 20.676 19.616 20.708 ;
  LAYER M2 ;
        RECT 21.952 20.612 21.984 20.644 ;
  LAYER M2 ;
        RECT 19.536 20.412 22.032 23.016 ;
  LAYER M1 ;
        RECT 22.56 36 22.592 38.508 ;
  LAYER M3 ;
        RECT 22.56 36.02 22.592 36.052 ;
  LAYER M1 ;
        RECT 22.624 36 22.656 38.508 ;
  LAYER M3 ;
        RECT 22.624 38.456 22.656 38.488 ;
  LAYER M1 ;
        RECT 22.688 36 22.72 38.508 ;
  LAYER M3 ;
        RECT 22.688 36.02 22.72 36.052 ;
  LAYER M1 ;
        RECT 22.752 36 22.784 38.508 ;
  LAYER M3 ;
        RECT 22.752 38.456 22.784 38.488 ;
  LAYER M1 ;
        RECT 22.816 36 22.848 38.508 ;
  LAYER M3 ;
        RECT 22.816 36.02 22.848 36.052 ;
  LAYER M1 ;
        RECT 22.88 36 22.912 38.508 ;
  LAYER M3 ;
        RECT 22.88 38.456 22.912 38.488 ;
  LAYER M1 ;
        RECT 22.944 36 22.976 38.508 ;
  LAYER M3 ;
        RECT 22.944 36.02 22.976 36.052 ;
  LAYER M1 ;
        RECT 23.008 36 23.04 38.508 ;
  LAYER M3 ;
        RECT 23.008 38.456 23.04 38.488 ;
  LAYER M1 ;
        RECT 23.072 36 23.104 38.508 ;
  LAYER M3 ;
        RECT 23.072 36.02 23.104 36.052 ;
  LAYER M1 ;
        RECT 23.136 36 23.168 38.508 ;
  LAYER M3 ;
        RECT 23.136 38.456 23.168 38.488 ;
  LAYER M1 ;
        RECT 23.2 36 23.232 38.508 ;
  LAYER M3 ;
        RECT 23.2 36.02 23.232 36.052 ;
  LAYER M1 ;
        RECT 23.264 36 23.296 38.508 ;
  LAYER M3 ;
        RECT 23.264 38.456 23.296 38.488 ;
  LAYER M1 ;
        RECT 23.328 36 23.36 38.508 ;
  LAYER M3 ;
        RECT 23.328 36.02 23.36 36.052 ;
  LAYER M1 ;
        RECT 23.392 36 23.424 38.508 ;
  LAYER M3 ;
        RECT 23.392 38.456 23.424 38.488 ;
  LAYER M1 ;
        RECT 23.456 36 23.488 38.508 ;
  LAYER M3 ;
        RECT 23.456 36.02 23.488 36.052 ;
  LAYER M1 ;
        RECT 23.52 36 23.552 38.508 ;
  LAYER M3 ;
        RECT 23.52 38.456 23.552 38.488 ;
  LAYER M1 ;
        RECT 23.584 36 23.616 38.508 ;
  LAYER M3 ;
        RECT 23.584 36.02 23.616 36.052 ;
  LAYER M1 ;
        RECT 23.648 36 23.68 38.508 ;
  LAYER M3 ;
        RECT 23.648 38.456 23.68 38.488 ;
  LAYER M1 ;
        RECT 23.712 36 23.744 38.508 ;
  LAYER M3 ;
        RECT 23.712 36.02 23.744 36.052 ;
  LAYER M1 ;
        RECT 23.776 36 23.808 38.508 ;
  LAYER M3 ;
        RECT 23.776 38.456 23.808 38.488 ;
  LAYER M1 ;
        RECT 23.84 36 23.872 38.508 ;
  LAYER M3 ;
        RECT 23.84 36.02 23.872 36.052 ;
  LAYER M1 ;
        RECT 23.904 36 23.936 38.508 ;
  LAYER M3 ;
        RECT 23.904 38.456 23.936 38.488 ;
  LAYER M1 ;
        RECT 23.968 36 24 38.508 ;
  LAYER M3 ;
        RECT 23.968 36.02 24 36.052 ;
  LAYER M1 ;
        RECT 24.032 36 24.064 38.508 ;
  LAYER M3 ;
        RECT 24.032 38.456 24.064 38.488 ;
  LAYER M1 ;
        RECT 24.096 36 24.128 38.508 ;
  LAYER M3 ;
        RECT 24.096 36.02 24.128 36.052 ;
  LAYER M1 ;
        RECT 24.16 36 24.192 38.508 ;
  LAYER M3 ;
        RECT 24.16 38.456 24.192 38.488 ;
  LAYER M1 ;
        RECT 24.224 36 24.256 38.508 ;
  LAYER M3 ;
        RECT 24.224 36.02 24.256 36.052 ;
  LAYER M1 ;
        RECT 24.288 36 24.32 38.508 ;
  LAYER M3 ;
        RECT 24.288 38.456 24.32 38.488 ;
  LAYER M1 ;
        RECT 24.352 36 24.384 38.508 ;
  LAYER M3 ;
        RECT 24.352 36.02 24.384 36.052 ;
  LAYER M1 ;
        RECT 24.416 36 24.448 38.508 ;
  LAYER M3 ;
        RECT 24.416 38.456 24.448 38.488 ;
  LAYER M1 ;
        RECT 24.48 36 24.512 38.508 ;
  LAYER M3 ;
        RECT 24.48 36.02 24.512 36.052 ;
  LAYER M1 ;
        RECT 24.544 36 24.576 38.508 ;
  LAYER M3 ;
        RECT 24.544 38.456 24.576 38.488 ;
  LAYER M1 ;
        RECT 24.608 36 24.64 38.508 ;
  LAYER M3 ;
        RECT 24.608 36.02 24.64 36.052 ;
  LAYER M1 ;
        RECT 24.672 36 24.704 38.508 ;
  LAYER M3 ;
        RECT 24.672 38.456 24.704 38.488 ;
  LAYER M1 ;
        RECT 24.736 36 24.768 38.508 ;
  LAYER M3 ;
        RECT 24.736 36.02 24.768 36.052 ;
  LAYER M1 ;
        RECT 24.8 36 24.832 38.508 ;
  LAYER M3 ;
        RECT 24.8 38.456 24.832 38.488 ;
  LAYER M1 ;
        RECT 24.864 36 24.896 38.508 ;
  LAYER M3 ;
        RECT 24.864 36.02 24.896 36.052 ;
  LAYER M1 ;
        RECT 24.928 36 24.96 38.508 ;
  LAYER M3 ;
        RECT 22.56 38.392 22.592 38.424 ;
  LAYER M2 ;
        RECT 24.928 38.328 24.96 38.36 ;
  LAYER M2 ;
        RECT 22.56 38.264 22.592 38.296 ;
  LAYER M2 ;
        RECT 24.928 38.2 24.96 38.232 ;
  LAYER M2 ;
        RECT 22.56 38.136 22.592 38.168 ;
  LAYER M2 ;
        RECT 24.928 38.072 24.96 38.104 ;
  LAYER M2 ;
        RECT 22.56 38.008 22.592 38.04 ;
  LAYER M2 ;
        RECT 24.928 37.944 24.96 37.976 ;
  LAYER M2 ;
        RECT 22.56 37.88 22.592 37.912 ;
  LAYER M2 ;
        RECT 24.928 37.816 24.96 37.848 ;
  LAYER M2 ;
        RECT 22.56 37.752 22.592 37.784 ;
  LAYER M2 ;
        RECT 24.928 37.688 24.96 37.72 ;
  LAYER M2 ;
        RECT 22.56 37.624 22.592 37.656 ;
  LAYER M2 ;
        RECT 24.928 37.56 24.96 37.592 ;
  LAYER M2 ;
        RECT 22.56 37.496 22.592 37.528 ;
  LAYER M2 ;
        RECT 24.928 37.432 24.96 37.464 ;
  LAYER M2 ;
        RECT 22.56 37.368 22.592 37.4 ;
  LAYER M2 ;
        RECT 24.928 37.304 24.96 37.336 ;
  LAYER M2 ;
        RECT 22.56 37.24 22.592 37.272 ;
  LAYER M2 ;
        RECT 24.928 37.176 24.96 37.208 ;
  LAYER M2 ;
        RECT 22.56 37.112 22.592 37.144 ;
  LAYER M2 ;
        RECT 24.928 37.048 24.96 37.08 ;
  LAYER M2 ;
        RECT 22.56 36.984 22.592 37.016 ;
  LAYER M2 ;
        RECT 24.928 36.92 24.96 36.952 ;
  LAYER M2 ;
        RECT 22.56 36.856 22.592 36.888 ;
  LAYER M2 ;
        RECT 24.928 36.792 24.96 36.824 ;
  LAYER M2 ;
        RECT 22.56 36.728 22.592 36.76 ;
  LAYER M2 ;
        RECT 24.928 36.664 24.96 36.696 ;
  LAYER M2 ;
        RECT 22.56 36.6 22.592 36.632 ;
  LAYER M2 ;
        RECT 24.928 36.536 24.96 36.568 ;
  LAYER M2 ;
        RECT 22.56 36.472 22.592 36.504 ;
  LAYER M2 ;
        RECT 24.928 36.408 24.96 36.44 ;
  LAYER M2 ;
        RECT 22.56 36.344 22.592 36.376 ;
  LAYER M2 ;
        RECT 24.928 36.28 24.96 36.312 ;
  LAYER M2 ;
        RECT 22.56 36.216 22.592 36.248 ;
  LAYER M2 ;
        RECT 24.928 36.152 24.96 36.184 ;
  LAYER M2 ;
        RECT 22.512 35.952 25.008 38.556 ;
  LAYER M1 ;
        RECT 22.56 32.892 22.592 35.4 ;
  LAYER M3 ;
        RECT 22.56 32.912 22.592 32.944 ;
  LAYER M1 ;
        RECT 22.624 32.892 22.656 35.4 ;
  LAYER M3 ;
        RECT 22.624 35.348 22.656 35.38 ;
  LAYER M1 ;
        RECT 22.688 32.892 22.72 35.4 ;
  LAYER M3 ;
        RECT 22.688 32.912 22.72 32.944 ;
  LAYER M1 ;
        RECT 22.752 32.892 22.784 35.4 ;
  LAYER M3 ;
        RECT 22.752 35.348 22.784 35.38 ;
  LAYER M1 ;
        RECT 22.816 32.892 22.848 35.4 ;
  LAYER M3 ;
        RECT 22.816 32.912 22.848 32.944 ;
  LAYER M1 ;
        RECT 22.88 32.892 22.912 35.4 ;
  LAYER M3 ;
        RECT 22.88 35.348 22.912 35.38 ;
  LAYER M1 ;
        RECT 22.944 32.892 22.976 35.4 ;
  LAYER M3 ;
        RECT 22.944 32.912 22.976 32.944 ;
  LAYER M1 ;
        RECT 23.008 32.892 23.04 35.4 ;
  LAYER M3 ;
        RECT 23.008 35.348 23.04 35.38 ;
  LAYER M1 ;
        RECT 23.072 32.892 23.104 35.4 ;
  LAYER M3 ;
        RECT 23.072 32.912 23.104 32.944 ;
  LAYER M1 ;
        RECT 23.136 32.892 23.168 35.4 ;
  LAYER M3 ;
        RECT 23.136 35.348 23.168 35.38 ;
  LAYER M1 ;
        RECT 23.2 32.892 23.232 35.4 ;
  LAYER M3 ;
        RECT 23.2 32.912 23.232 32.944 ;
  LAYER M1 ;
        RECT 23.264 32.892 23.296 35.4 ;
  LAYER M3 ;
        RECT 23.264 35.348 23.296 35.38 ;
  LAYER M1 ;
        RECT 23.328 32.892 23.36 35.4 ;
  LAYER M3 ;
        RECT 23.328 32.912 23.36 32.944 ;
  LAYER M1 ;
        RECT 23.392 32.892 23.424 35.4 ;
  LAYER M3 ;
        RECT 23.392 35.348 23.424 35.38 ;
  LAYER M1 ;
        RECT 23.456 32.892 23.488 35.4 ;
  LAYER M3 ;
        RECT 23.456 32.912 23.488 32.944 ;
  LAYER M1 ;
        RECT 23.52 32.892 23.552 35.4 ;
  LAYER M3 ;
        RECT 23.52 35.348 23.552 35.38 ;
  LAYER M1 ;
        RECT 23.584 32.892 23.616 35.4 ;
  LAYER M3 ;
        RECT 23.584 32.912 23.616 32.944 ;
  LAYER M1 ;
        RECT 23.648 32.892 23.68 35.4 ;
  LAYER M3 ;
        RECT 23.648 35.348 23.68 35.38 ;
  LAYER M1 ;
        RECT 23.712 32.892 23.744 35.4 ;
  LAYER M3 ;
        RECT 23.712 32.912 23.744 32.944 ;
  LAYER M1 ;
        RECT 23.776 32.892 23.808 35.4 ;
  LAYER M3 ;
        RECT 23.776 35.348 23.808 35.38 ;
  LAYER M1 ;
        RECT 23.84 32.892 23.872 35.4 ;
  LAYER M3 ;
        RECT 23.84 32.912 23.872 32.944 ;
  LAYER M1 ;
        RECT 23.904 32.892 23.936 35.4 ;
  LAYER M3 ;
        RECT 23.904 35.348 23.936 35.38 ;
  LAYER M1 ;
        RECT 23.968 32.892 24 35.4 ;
  LAYER M3 ;
        RECT 23.968 32.912 24 32.944 ;
  LAYER M1 ;
        RECT 24.032 32.892 24.064 35.4 ;
  LAYER M3 ;
        RECT 24.032 35.348 24.064 35.38 ;
  LAYER M1 ;
        RECT 24.096 32.892 24.128 35.4 ;
  LAYER M3 ;
        RECT 24.096 32.912 24.128 32.944 ;
  LAYER M1 ;
        RECT 24.16 32.892 24.192 35.4 ;
  LAYER M3 ;
        RECT 24.16 35.348 24.192 35.38 ;
  LAYER M1 ;
        RECT 24.224 32.892 24.256 35.4 ;
  LAYER M3 ;
        RECT 24.224 32.912 24.256 32.944 ;
  LAYER M1 ;
        RECT 24.288 32.892 24.32 35.4 ;
  LAYER M3 ;
        RECT 24.288 35.348 24.32 35.38 ;
  LAYER M1 ;
        RECT 24.352 32.892 24.384 35.4 ;
  LAYER M3 ;
        RECT 24.352 32.912 24.384 32.944 ;
  LAYER M1 ;
        RECT 24.416 32.892 24.448 35.4 ;
  LAYER M3 ;
        RECT 24.416 35.348 24.448 35.38 ;
  LAYER M1 ;
        RECT 24.48 32.892 24.512 35.4 ;
  LAYER M3 ;
        RECT 24.48 32.912 24.512 32.944 ;
  LAYER M1 ;
        RECT 24.544 32.892 24.576 35.4 ;
  LAYER M3 ;
        RECT 24.544 35.348 24.576 35.38 ;
  LAYER M1 ;
        RECT 24.608 32.892 24.64 35.4 ;
  LAYER M3 ;
        RECT 24.608 32.912 24.64 32.944 ;
  LAYER M1 ;
        RECT 24.672 32.892 24.704 35.4 ;
  LAYER M3 ;
        RECT 24.672 35.348 24.704 35.38 ;
  LAYER M1 ;
        RECT 24.736 32.892 24.768 35.4 ;
  LAYER M3 ;
        RECT 24.736 32.912 24.768 32.944 ;
  LAYER M1 ;
        RECT 24.8 32.892 24.832 35.4 ;
  LAYER M3 ;
        RECT 24.8 35.348 24.832 35.38 ;
  LAYER M1 ;
        RECT 24.864 32.892 24.896 35.4 ;
  LAYER M3 ;
        RECT 24.864 32.912 24.896 32.944 ;
  LAYER M1 ;
        RECT 24.928 32.892 24.96 35.4 ;
  LAYER M3 ;
        RECT 22.56 35.284 22.592 35.316 ;
  LAYER M2 ;
        RECT 24.928 35.22 24.96 35.252 ;
  LAYER M2 ;
        RECT 22.56 35.156 22.592 35.188 ;
  LAYER M2 ;
        RECT 24.928 35.092 24.96 35.124 ;
  LAYER M2 ;
        RECT 22.56 35.028 22.592 35.06 ;
  LAYER M2 ;
        RECT 24.928 34.964 24.96 34.996 ;
  LAYER M2 ;
        RECT 22.56 34.9 22.592 34.932 ;
  LAYER M2 ;
        RECT 24.928 34.836 24.96 34.868 ;
  LAYER M2 ;
        RECT 22.56 34.772 22.592 34.804 ;
  LAYER M2 ;
        RECT 24.928 34.708 24.96 34.74 ;
  LAYER M2 ;
        RECT 22.56 34.644 22.592 34.676 ;
  LAYER M2 ;
        RECT 24.928 34.58 24.96 34.612 ;
  LAYER M2 ;
        RECT 22.56 34.516 22.592 34.548 ;
  LAYER M2 ;
        RECT 24.928 34.452 24.96 34.484 ;
  LAYER M2 ;
        RECT 22.56 34.388 22.592 34.42 ;
  LAYER M2 ;
        RECT 24.928 34.324 24.96 34.356 ;
  LAYER M2 ;
        RECT 22.56 34.26 22.592 34.292 ;
  LAYER M2 ;
        RECT 24.928 34.196 24.96 34.228 ;
  LAYER M2 ;
        RECT 22.56 34.132 22.592 34.164 ;
  LAYER M2 ;
        RECT 24.928 34.068 24.96 34.1 ;
  LAYER M2 ;
        RECT 22.56 34.004 22.592 34.036 ;
  LAYER M2 ;
        RECT 24.928 33.94 24.96 33.972 ;
  LAYER M2 ;
        RECT 22.56 33.876 22.592 33.908 ;
  LAYER M2 ;
        RECT 24.928 33.812 24.96 33.844 ;
  LAYER M2 ;
        RECT 22.56 33.748 22.592 33.78 ;
  LAYER M2 ;
        RECT 24.928 33.684 24.96 33.716 ;
  LAYER M2 ;
        RECT 22.56 33.62 22.592 33.652 ;
  LAYER M2 ;
        RECT 24.928 33.556 24.96 33.588 ;
  LAYER M2 ;
        RECT 22.56 33.492 22.592 33.524 ;
  LAYER M2 ;
        RECT 24.928 33.428 24.96 33.46 ;
  LAYER M2 ;
        RECT 22.56 33.364 22.592 33.396 ;
  LAYER M2 ;
        RECT 24.928 33.3 24.96 33.332 ;
  LAYER M2 ;
        RECT 22.56 33.236 22.592 33.268 ;
  LAYER M2 ;
        RECT 24.928 33.172 24.96 33.204 ;
  LAYER M2 ;
        RECT 22.56 33.108 22.592 33.14 ;
  LAYER M2 ;
        RECT 24.928 33.044 24.96 33.076 ;
  LAYER M2 ;
        RECT 22.512 32.844 25.008 35.448 ;
  LAYER M1 ;
        RECT 22.56 29.784 22.592 32.292 ;
  LAYER M3 ;
        RECT 22.56 29.804 22.592 29.836 ;
  LAYER M1 ;
        RECT 22.624 29.784 22.656 32.292 ;
  LAYER M3 ;
        RECT 22.624 32.24 22.656 32.272 ;
  LAYER M1 ;
        RECT 22.688 29.784 22.72 32.292 ;
  LAYER M3 ;
        RECT 22.688 29.804 22.72 29.836 ;
  LAYER M1 ;
        RECT 22.752 29.784 22.784 32.292 ;
  LAYER M3 ;
        RECT 22.752 32.24 22.784 32.272 ;
  LAYER M1 ;
        RECT 22.816 29.784 22.848 32.292 ;
  LAYER M3 ;
        RECT 22.816 29.804 22.848 29.836 ;
  LAYER M1 ;
        RECT 22.88 29.784 22.912 32.292 ;
  LAYER M3 ;
        RECT 22.88 32.24 22.912 32.272 ;
  LAYER M1 ;
        RECT 22.944 29.784 22.976 32.292 ;
  LAYER M3 ;
        RECT 22.944 29.804 22.976 29.836 ;
  LAYER M1 ;
        RECT 23.008 29.784 23.04 32.292 ;
  LAYER M3 ;
        RECT 23.008 32.24 23.04 32.272 ;
  LAYER M1 ;
        RECT 23.072 29.784 23.104 32.292 ;
  LAYER M3 ;
        RECT 23.072 29.804 23.104 29.836 ;
  LAYER M1 ;
        RECT 23.136 29.784 23.168 32.292 ;
  LAYER M3 ;
        RECT 23.136 32.24 23.168 32.272 ;
  LAYER M1 ;
        RECT 23.2 29.784 23.232 32.292 ;
  LAYER M3 ;
        RECT 23.2 29.804 23.232 29.836 ;
  LAYER M1 ;
        RECT 23.264 29.784 23.296 32.292 ;
  LAYER M3 ;
        RECT 23.264 32.24 23.296 32.272 ;
  LAYER M1 ;
        RECT 23.328 29.784 23.36 32.292 ;
  LAYER M3 ;
        RECT 23.328 29.804 23.36 29.836 ;
  LAYER M1 ;
        RECT 23.392 29.784 23.424 32.292 ;
  LAYER M3 ;
        RECT 23.392 32.24 23.424 32.272 ;
  LAYER M1 ;
        RECT 23.456 29.784 23.488 32.292 ;
  LAYER M3 ;
        RECT 23.456 29.804 23.488 29.836 ;
  LAYER M1 ;
        RECT 23.52 29.784 23.552 32.292 ;
  LAYER M3 ;
        RECT 23.52 32.24 23.552 32.272 ;
  LAYER M1 ;
        RECT 23.584 29.784 23.616 32.292 ;
  LAYER M3 ;
        RECT 23.584 29.804 23.616 29.836 ;
  LAYER M1 ;
        RECT 23.648 29.784 23.68 32.292 ;
  LAYER M3 ;
        RECT 23.648 32.24 23.68 32.272 ;
  LAYER M1 ;
        RECT 23.712 29.784 23.744 32.292 ;
  LAYER M3 ;
        RECT 23.712 29.804 23.744 29.836 ;
  LAYER M1 ;
        RECT 23.776 29.784 23.808 32.292 ;
  LAYER M3 ;
        RECT 23.776 32.24 23.808 32.272 ;
  LAYER M1 ;
        RECT 23.84 29.784 23.872 32.292 ;
  LAYER M3 ;
        RECT 23.84 29.804 23.872 29.836 ;
  LAYER M1 ;
        RECT 23.904 29.784 23.936 32.292 ;
  LAYER M3 ;
        RECT 23.904 32.24 23.936 32.272 ;
  LAYER M1 ;
        RECT 23.968 29.784 24 32.292 ;
  LAYER M3 ;
        RECT 23.968 29.804 24 29.836 ;
  LAYER M1 ;
        RECT 24.032 29.784 24.064 32.292 ;
  LAYER M3 ;
        RECT 24.032 32.24 24.064 32.272 ;
  LAYER M1 ;
        RECT 24.096 29.784 24.128 32.292 ;
  LAYER M3 ;
        RECT 24.096 29.804 24.128 29.836 ;
  LAYER M1 ;
        RECT 24.16 29.784 24.192 32.292 ;
  LAYER M3 ;
        RECT 24.16 32.24 24.192 32.272 ;
  LAYER M1 ;
        RECT 24.224 29.784 24.256 32.292 ;
  LAYER M3 ;
        RECT 24.224 29.804 24.256 29.836 ;
  LAYER M1 ;
        RECT 24.288 29.784 24.32 32.292 ;
  LAYER M3 ;
        RECT 24.288 32.24 24.32 32.272 ;
  LAYER M1 ;
        RECT 24.352 29.784 24.384 32.292 ;
  LAYER M3 ;
        RECT 24.352 29.804 24.384 29.836 ;
  LAYER M1 ;
        RECT 24.416 29.784 24.448 32.292 ;
  LAYER M3 ;
        RECT 24.416 32.24 24.448 32.272 ;
  LAYER M1 ;
        RECT 24.48 29.784 24.512 32.292 ;
  LAYER M3 ;
        RECT 24.48 29.804 24.512 29.836 ;
  LAYER M1 ;
        RECT 24.544 29.784 24.576 32.292 ;
  LAYER M3 ;
        RECT 24.544 32.24 24.576 32.272 ;
  LAYER M1 ;
        RECT 24.608 29.784 24.64 32.292 ;
  LAYER M3 ;
        RECT 24.608 29.804 24.64 29.836 ;
  LAYER M1 ;
        RECT 24.672 29.784 24.704 32.292 ;
  LAYER M3 ;
        RECT 24.672 32.24 24.704 32.272 ;
  LAYER M1 ;
        RECT 24.736 29.784 24.768 32.292 ;
  LAYER M3 ;
        RECT 24.736 29.804 24.768 29.836 ;
  LAYER M1 ;
        RECT 24.8 29.784 24.832 32.292 ;
  LAYER M3 ;
        RECT 24.8 32.24 24.832 32.272 ;
  LAYER M1 ;
        RECT 24.864 29.784 24.896 32.292 ;
  LAYER M3 ;
        RECT 24.864 29.804 24.896 29.836 ;
  LAYER M1 ;
        RECT 24.928 29.784 24.96 32.292 ;
  LAYER M3 ;
        RECT 22.56 32.176 22.592 32.208 ;
  LAYER M2 ;
        RECT 24.928 32.112 24.96 32.144 ;
  LAYER M2 ;
        RECT 22.56 32.048 22.592 32.08 ;
  LAYER M2 ;
        RECT 24.928 31.984 24.96 32.016 ;
  LAYER M2 ;
        RECT 22.56 31.92 22.592 31.952 ;
  LAYER M2 ;
        RECT 24.928 31.856 24.96 31.888 ;
  LAYER M2 ;
        RECT 22.56 31.792 22.592 31.824 ;
  LAYER M2 ;
        RECT 24.928 31.728 24.96 31.76 ;
  LAYER M2 ;
        RECT 22.56 31.664 22.592 31.696 ;
  LAYER M2 ;
        RECT 24.928 31.6 24.96 31.632 ;
  LAYER M2 ;
        RECT 22.56 31.536 22.592 31.568 ;
  LAYER M2 ;
        RECT 24.928 31.472 24.96 31.504 ;
  LAYER M2 ;
        RECT 22.56 31.408 22.592 31.44 ;
  LAYER M2 ;
        RECT 24.928 31.344 24.96 31.376 ;
  LAYER M2 ;
        RECT 22.56 31.28 22.592 31.312 ;
  LAYER M2 ;
        RECT 24.928 31.216 24.96 31.248 ;
  LAYER M2 ;
        RECT 22.56 31.152 22.592 31.184 ;
  LAYER M2 ;
        RECT 24.928 31.088 24.96 31.12 ;
  LAYER M2 ;
        RECT 22.56 31.024 22.592 31.056 ;
  LAYER M2 ;
        RECT 24.928 30.96 24.96 30.992 ;
  LAYER M2 ;
        RECT 22.56 30.896 22.592 30.928 ;
  LAYER M2 ;
        RECT 24.928 30.832 24.96 30.864 ;
  LAYER M2 ;
        RECT 22.56 30.768 22.592 30.8 ;
  LAYER M2 ;
        RECT 24.928 30.704 24.96 30.736 ;
  LAYER M2 ;
        RECT 22.56 30.64 22.592 30.672 ;
  LAYER M2 ;
        RECT 24.928 30.576 24.96 30.608 ;
  LAYER M2 ;
        RECT 22.56 30.512 22.592 30.544 ;
  LAYER M2 ;
        RECT 24.928 30.448 24.96 30.48 ;
  LAYER M2 ;
        RECT 22.56 30.384 22.592 30.416 ;
  LAYER M2 ;
        RECT 24.928 30.32 24.96 30.352 ;
  LAYER M2 ;
        RECT 22.56 30.256 22.592 30.288 ;
  LAYER M2 ;
        RECT 24.928 30.192 24.96 30.224 ;
  LAYER M2 ;
        RECT 22.56 30.128 22.592 30.16 ;
  LAYER M2 ;
        RECT 24.928 30.064 24.96 30.096 ;
  LAYER M2 ;
        RECT 22.56 30 22.592 30.032 ;
  LAYER M2 ;
        RECT 24.928 29.936 24.96 29.968 ;
  LAYER M2 ;
        RECT 22.512 29.736 25.008 32.34 ;
  LAYER M1 ;
        RECT 22.56 26.676 22.592 29.184 ;
  LAYER M3 ;
        RECT 22.56 26.696 22.592 26.728 ;
  LAYER M1 ;
        RECT 22.624 26.676 22.656 29.184 ;
  LAYER M3 ;
        RECT 22.624 29.132 22.656 29.164 ;
  LAYER M1 ;
        RECT 22.688 26.676 22.72 29.184 ;
  LAYER M3 ;
        RECT 22.688 26.696 22.72 26.728 ;
  LAYER M1 ;
        RECT 22.752 26.676 22.784 29.184 ;
  LAYER M3 ;
        RECT 22.752 29.132 22.784 29.164 ;
  LAYER M1 ;
        RECT 22.816 26.676 22.848 29.184 ;
  LAYER M3 ;
        RECT 22.816 26.696 22.848 26.728 ;
  LAYER M1 ;
        RECT 22.88 26.676 22.912 29.184 ;
  LAYER M3 ;
        RECT 22.88 29.132 22.912 29.164 ;
  LAYER M1 ;
        RECT 22.944 26.676 22.976 29.184 ;
  LAYER M3 ;
        RECT 22.944 26.696 22.976 26.728 ;
  LAYER M1 ;
        RECT 23.008 26.676 23.04 29.184 ;
  LAYER M3 ;
        RECT 23.008 29.132 23.04 29.164 ;
  LAYER M1 ;
        RECT 23.072 26.676 23.104 29.184 ;
  LAYER M3 ;
        RECT 23.072 26.696 23.104 26.728 ;
  LAYER M1 ;
        RECT 23.136 26.676 23.168 29.184 ;
  LAYER M3 ;
        RECT 23.136 29.132 23.168 29.164 ;
  LAYER M1 ;
        RECT 23.2 26.676 23.232 29.184 ;
  LAYER M3 ;
        RECT 23.2 26.696 23.232 26.728 ;
  LAYER M1 ;
        RECT 23.264 26.676 23.296 29.184 ;
  LAYER M3 ;
        RECT 23.264 29.132 23.296 29.164 ;
  LAYER M1 ;
        RECT 23.328 26.676 23.36 29.184 ;
  LAYER M3 ;
        RECT 23.328 26.696 23.36 26.728 ;
  LAYER M1 ;
        RECT 23.392 26.676 23.424 29.184 ;
  LAYER M3 ;
        RECT 23.392 29.132 23.424 29.164 ;
  LAYER M1 ;
        RECT 23.456 26.676 23.488 29.184 ;
  LAYER M3 ;
        RECT 23.456 26.696 23.488 26.728 ;
  LAYER M1 ;
        RECT 23.52 26.676 23.552 29.184 ;
  LAYER M3 ;
        RECT 23.52 29.132 23.552 29.164 ;
  LAYER M1 ;
        RECT 23.584 26.676 23.616 29.184 ;
  LAYER M3 ;
        RECT 23.584 26.696 23.616 26.728 ;
  LAYER M1 ;
        RECT 23.648 26.676 23.68 29.184 ;
  LAYER M3 ;
        RECT 23.648 29.132 23.68 29.164 ;
  LAYER M1 ;
        RECT 23.712 26.676 23.744 29.184 ;
  LAYER M3 ;
        RECT 23.712 26.696 23.744 26.728 ;
  LAYER M1 ;
        RECT 23.776 26.676 23.808 29.184 ;
  LAYER M3 ;
        RECT 23.776 29.132 23.808 29.164 ;
  LAYER M1 ;
        RECT 23.84 26.676 23.872 29.184 ;
  LAYER M3 ;
        RECT 23.84 26.696 23.872 26.728 ;
  LAYER M1 ;
        RECT 23.904 26.676 23.936 29.184 ;
  LAYER M3 ;
        RECT 23.904 29.132 23.936 29.164 ;
  LAYER M1 ;
        RECT 23.968 26.676 24 29.184 ;
  LAYER M3 ;
        RECT 23.968 26.696 24 26.728 ;
  LAYER M1 ;
        RECT 24.032 26.676 24.064 29.184 ;
  LAYER M3 ;
        RECT 24.032 29.132 24.064 29.164 ;
  LAYER M1 ;
        RECT 24.096 26.676 24.128 29.184 ;
  LAYER M3 ;
        RECT 24.096 26.696 24.128 26.728 ;
  LAYER M1 ;
        RECT 24.16 26.676 24.192 29.184 ;
  LAYER M3 ;
        RECT 24.16 29.132 24.192 29.164 ;
  LAYER M1 ;
        RECT 24.224 26.676 24.256 29.184 ;
  LAYER M3 ;
        RECT 24.224 26.696 24.256 26.728 ;
  LAYER M1 ;
        RECT 24.288 26.676 24.32 29.184 ;
  LAYER M3 ;
        RECT 24.288 29.132 24.32 29.164 ;
  LAYER M1 ;
        RECT 24.352 26.676 24.384 29.184 ;
  LAYER M3 ;
        RECT 24.352 26.696 24.384 26.728 ;
  LAYER M1 ;
        RECT 24.416 26.676 24.448 29.184 ;
  LAYER M3 ;
        RECT 24.416 29.132 24.448 29.164 ;
  LAYER M1 ;
        RECT 24.48 26.676 24.512 29.184 ;
  LAYER M3 ;
        RECT 24.48 26.696 24.512 26.728 ;
  LAYER M1 ;
        RECT 24.544 26.676 24.576 29.184 ;
  LAYER M3 ;
        RECT 24.544 29.132 24.576 29.164 ;
  LAYER M1 ;
        RECT 24.608 26.676 24.64 29.184 ;
  LAYER M3 ;
        RECT 24.608 26.696 24.64 26.728 ;
  LAYER M1 ;
        RECT 24.672 26.676 24.704 29.184 ;
  LAYER M3 ;
        RECT 24.672 29.132 24.704 29.164 ;
  LAYER M1 ;
        RECT 24.736 26.676 24.768 29.184 ;
  LAYER M3 ;
        RECT 24.736 26.696 24.768 26.728 ;
  LAYER M1 ;
        RECT 24.8 26.676 24.832 29.184 ;
  LAYER M3 ;
        RECT 24.8 29.132 24.832 29.164 ;
  LAYER M1 ;
        RECT 24.864 26.676 24.896 29.184 ;
  LAYER M3 ;
        RECT 24.864 26.696 24.896 26.728 ;
  LAYER M1 ;
        RECT 24.928 26.676 24.96 29.184 ;
  LAYER M3 ;
        RECT 22.56 29.068 22.592 29.1 ;
  LAYER M2 ;
        RECT 24.928 29.004 24.96 29.036 ;
  LAYER M2 ;
        RECT 22.56 28.94 22.592 28.972 ;
  LAYER M2 ;
        RECT 24.928 28.876 24.96 28.908 ;
  LAYER M2 ;
        RECT 22.56 28.812 22.592 28.844 ;
  LAYER M2 ;
        RECT 24.928 28.748 24.96 28.78 ;
  LAYER M2 ;
        RECT 22.56 28.684 22.592 28.716 ;
  LAYER M2 ;
        RECT 24.928 28.62 24.96 28.652 ;
  LAYER M2 ;
        RECT 22.56 28.556 22.592 28.588 ;
  LAYER M2 ;
        RECT 24.928 28.492 24.96 28.524 ;
  LAYER M2 ;
        RECT 22.56 28.428 22.592 28.46 ;
  LAYER M2 ;
        RECT 24.928 28.364 24.96 28.396 ;
  LAYER M2 ;
        RECT 22.56 28.3 22.592 28.332 ;
  LAYER M2 ;
        RECT 24.928 28.236 24.96 28.268 ;
  LAYER M2 ;
        RECT 22.56 28.172 22.592 28.204 ;
  LAYER M2 ;
        RECT 24.928 28.108 24.96 28.14 ;
  LAYER M2 ;
        RECT 22.56 28.044 22.592 28.076 ;
  LAYER M2 ;
        RECT 24.928 27.98 24.96 28.012 ;
  LAYER M2 ;
        RECT 22.56 27.916 22.592 27.948 ;
  LAYER M2 ;
        RECT 24.928 27.852 24.96 27.884 ;
  LAYER M2 ;
        RECT 22.56 27.788 22.592 27.82 ;
  LAYER M2 ;
        RECT 24.928 27.724 24.96 27.756 ;
  LAYER M2 ;
        RECT 22.56 27.66 22.592 27.692 ;
  LAYER M2 ;
        RECT 24.928 27.596 24.96 27.628 ;
  LAYER M2 ;
        RECT 22.56 27.532 22.592 27.564 ;
  LAYER M2 ;
        RECT 24.928 27.468 24.96 27.5 ;
  LAYER M2 ;
        RECT 22.56 27.404 22.592 27.436 ;
  LAYER M2 ;
        RECT 24.928 27.34 24.96 27.372 ;
  LAYER M2 ;
        RECT 22.56 27.276 22.592 27.308 ;
  LAYER M2 ;
        RECT 24.928 27.212 24.96 27.244 ;
  LAYER M2 ;
        RECT 22.56 27.148 22.592 27.18 ;
  LAYER M2 ;
        RECT 24.928 27.084 24.96 27.116 ;
  LAYER M2 ;
        RECT 22.56 27.02 22.592 27.052 ;
  LAYER M2 ;
        RECT 24.928 26.956 24.96 26.988 ;
  LAYER M2 ;
        RECT 22.56 26.892 22.592 26.924 ;
  LAYER M2 ;
        RECT 24.928 26.828 24.96 26.86 ;
  LAYER M2 ;
        RECT 22.512 26.628 25.008 29.232 ;
  LAYER M1 ;
        RECT 22.56 23.568 22.592 26.076 ;
  LAYER M3 ;
        RECT 22.56 23.588 22.592 23.62 ;
  LAYER M1 ;
        RECT 22.624 23.568 22.656 26.076 ;
  LAYER M3 ;
        RECT 22.624 26.024 22.656 26.056 ;
  LAYER M1 ;
        RECT 22.688 23.568 22.72 26.076 ;
  LAYER M3 ;
        RECT 22.688 23.588 22.72 23.62 ;
  LAYER M1 ;
        RECT 22.752 23.568 22.784 26.076 ;
  LAYER M3 ;
        RECT 22.752 26.024 22.784 26.056 ;
  LAYER M1 ;
        RECT 22.816 23.568 22.848 26.076 ;
  LAYER M3 ;
        RECT 22.816 23.588 22.848 23.62 ;
  LAYER M1 ;
        RECT 22.88 23.568 22.912 26.076 ;
  LAYER M3 ;
        RECT 22.88 26.024 22.912 26.056 ;
  LAYER M1 ;
        RECT 22.944 23.568 22.976 26.076 ;
  LAYER M3 ;
        RECT 22.944 23.588 22.976 23.62 ;
  LAYER M1 ;
        RECT 23.008 23.568 23.04 26.076 ;
  LAYER M3 ;
        RECT 23.008 26.024 23.04 26.056 ;
  LAYER M1 ;
        RECT 23.072 23.568 23.104 26.076 ;
  LAYER M3 ;
        RECT 23.072 23.588 23.104 23.62 ;
  LAYER M1 ;
        RECT 23.136 23.568 23.168 26.076 ;
  LAYER M3 ;
        RECT 23.136 26.024 23.168 26.056 ;
  LAYER M1 ;
        RECT 23.2 23.568 23.232 26.076 ;
  LAYER M3 ;
        RECT 23.2 23.588 23.232 23.62 ;
  LAYER M1 ;
        RECT 23.264 23.568 23.296 26.076 ;
  LAYER M3 ;
        RECT 23.264 26.024 23.296 26.056 ;
  LAYER M1 ;
        RECT 23.328 23.568 23.36 26.076 ;
  LAYER M3 ;
        RECT 23.328 23.588 23.36 23.62 ;
  LAYER M1 ;
        RECT 23.392 23.568 23.424 26.076 ;
  LAYER M3 ;
        RECT 23.392 26.024 23.424 26.056 ;
  LAYER M1 ;
        RECT 23.456 23.568 23.488 26.076 ;
  LAYER M3 ;
        RECT 23.456 23.588 23.488 23.62 ;
  LAYER M1 ;
        RECT 23.52 23.568 23.552 26.076 ;
  LAYER M3 ;
        RECT 23.52 26.024 23.552 26.056 ;
  LAYER M1 ;
        RECT 23.584 23.568 23.616 26.076 ;
  LAYER M3 ;
        RECT 23.584 23.588 23.616 23.62 ;
  LAYER M1 ;
        RECT 23.648 23.568 23.68 26.076 ;
  LAYER M3 ;
        RECT 23.648 26.024 23.68 26.056 ;
  LAYER M1 ;
        RECT 23.712 23.568 23.744 26.076 ;
  LAYER M3 ;
        RECT 23.712 23.588 23.744 23.62 ;
  LAYER M1 ;
        RECT 23.776 23.568 23.808 26.076 ;
  LAYER M3 ;
        RECT 23.776 26.024 23.808 26.056 ;
  LAYER M1 ;
        RECT 23.84 23.568 23.872 26.076 ;
  LAYER M3 ;
        RECT 23.84 23.588 23.872 23.62 ;
  LAYER M1 ;
        RECT 23.904 23.568 23.936 26.076 ;
  LAYER M3 ;
        RECT 23.904 26.024 23.936 26.056 ;
  LAYER M1 ;
        RECT 23.968 23.568 24 26.076 ;
  LAYER M3 ;
        RECT 23.968 23.588 24 23.62 ;
  LAYER M1 ;
        RECT 24.032 23.568 24.064 26.076 ;
  LAYER M3 ;
        RECT 24.032 26.024 24.064 26.056 ;
  LAYER M1 ;
        RECT 24.096 23.568 24.128 26.076 ;
  LAYER M3 ;
        RECT 24.096 23.588 24.128 23.62 ;
  LAYER M1 ;
        RECT 24.16 23.568 24.192 26.076 ;
  LAYER M3 ;
        RECT 24.16 26.024 24.192 26.056 ;
  LAYER M1 ;
        RECT 24.224 23.568 24.256 26.076 ;
  LAYER M3 ;
        RECT 24.224 23.588 24.256 23.62 ;
  LAYER M1 ;
        RECT 24.288 23.568 24.32 26.076 ;
  LAYER M3 ;
        RECT 24.288 26.024 24.32 26.056 ;
  LAYER M1 ;
        RECT 24.352 23.568 24.384 26.076 ;
  LAYER M3 ;
        RECT 24.352 23.588 24.384 23.62 ;
  LAYER M1 ;
        RECT 24.416 23.568 24.448 26.076 ;
  LAYER M3 ;
        RECT 24.416 26.024 24.448 26.056 ;
  LAYER M1 ;
        RECT 24.48 23.568 24.512 26.076 ;
  LAYER M3 ;
        RECT 24.48 23.588 24.512 23.62 ;
  LAYER M1 ;
        RECT 24.544 23.568 24.576 26.076 ;
  LAYER M3 ;
        RECT 24.544 26.024 24.576 26.056 ;
  LAYER M1 ;
        RECT 24.608 23.568 24.64 26.076 ;
  LAYER M3 ;
        RECT 24.608 23.588 24.64 23.62 ;
  LAYER M1 ;
        RECT 24.672 23.568 24.704 26.076 ;
  LAYER M3 ;
        RECT 24.672 26.024 24.704 26.056 ;
  LAYER M1 ;
        RECT 24.736 23.568 24.768 26.076 ;
  LAYER M3 ;
        RECT 24.736 23.588 24.768 23.62 ;
  LAYER M1 ;
        RECT 24.8 23.568 24.832 26.076 ;
  LAYER M3 ;
        RECT 24.8 26.024 24.832 26.056 ;
  LAYER M1 ;
        RECT 24.864 23.568 24.896 26.076 ;
  LAYER M3 ;
        RECT 24.864 23.588 24.896 23.62 ;
  LAYER M1 ;
        RECT 24.928 23.568 24.96 26.076 ;
  LAYER M3 ;
        RECT 22.56 25.96 22.592 25.992 ;
  LAYER M2 ;
        RECT 24.928 25.896 24.96 25.928 ;
  LAYER M2 ;
        RECT 22.56 25.832 22.592 25.864 ;
  LAYER M2 ;
        RECT 24.928 25.768 24.96 25.8 ;
  LAYER M2 ;
        RECT 22.56 25.704 22.592 25.736 ;
  LAYER M2 ;
        RECT 24.928 25.64 24.96 25.672 ;
  LAYER M2 ;
        RECT 22.56 25.576 22.592 25.608 ;
  LAYER M2 ;
        RECT 24.928 25.512 24.96 25.544 ;
  LAYER M2 ;
        RECT 22.56 25.448 22.592 25.48 ;
  LAYER M2 ;
        RECT 24.928 25.384 24.96 25.416 ;
  LAYER M2 ;
        RECT 22.56 25.32 22.592 25.352 ;
  LAYER M2 ;
        RECT 24.928 25.256 24.96 25.288 ;
  LAYER M2 ;
        RECT 22.56 25.192 22.592 25.224 ;
  LAYER M2 ;
        RECT 24.928 25.128 24.96 25.16 ;
  LAYER M2 ;
        RECT 22.56 25.064 22.592 25.096 ;
  LAYER M2 ;
        RECT 24.928 25 24.96 25.032 ;
  LAYER M2 ;
        RECT 22.56 24.936 22.592 24.968 ;
  LAYER M2 ;
        RECT 24.928 24.872 24.96 24.904 ;
  LAYER M2 ;
        RECT 22.56 24.808 22.592 24.84 ;
  LAYER M2 ;
        RECT 24.928 24.744 24.96 24.776 ;
  LAYER M2 ;
        RECT 22.56 24.68 22.592 24.712 ;
  LAYER M2 ;
        RECT 24.928 24.616 24.96 24.648 ;
  LAYER M2 ;
        RECT 22.56 24.552 22.592 24.584 ;
  LAYER M2 ;
        RECT 24.928 24.488 24.96 24.52 ;
  LAYER M2 ;
        RECT 22.56 24.424 22.592 24.456 ;
  LAYER M2 ;
        RECT 24.928 24.36 24.96 24.392 ;
  LAYER M2 ;
        RECT 22.56 24.296 22.592 24.328 ;
  LAYER M2 ;
        RECT 24.928 24.232 24.96 24.264 ;
  LAYER M2 ;
        RECT 22.56 24.168 22.592 24.2 ;
  LAYER M2 ;
        RECT 24.928 24.104 24.96 24.136 ;
  LAYER M2 ;
        RECT 22.56 24.04 22.592 24.072 ;
  LAYER M2 ;
        RECT 24.928 23.976 24.96 24.008 ;
  LAYER M2 ;
        RECT 22.56 23.912 22.592 23.944 ;
  LAYER M2 ;
        RECT 24.928 23.848 24.96 23.88 ;
  LAYER M2 ;
        RECT 22.56 23.784 22.592 23.816 ;
  LAYER M2 ;
        RECT 24.928 23.72 24.96 23.752 ;
  LAYER M2 ;
        RECT 22.512 23.52 25.008 26.124 ;
  LAYER M1 ;
        RECT 22.56 20.46 22.592 22.968 ;
  LAYER M3 ;
        RECT 22.56 20.48 22.592 20.512 ;
  LAYER M1 ;
        RECT 22.624 20.46 22.656 22.968 ;
  LAYER M3 ;
        RECT 22.624 22.916 22.656 22.948 ;
  LAYER M1 ;
        RECT 22.688 20.46 22.72 22.968 ;
  LAYER M3 ;
        RECT 22.688 20.48 22.72 20.512 ;
  LAYER M1 ;
        RECT 22.752 20.46 22.784 22.968 ;
  LAYER M3 ;
        RECT 22.752 22.916 22.784 22.948 ;
  LAYER M1 ;
        RECT 22.816 20.46 22.848 22.968 ;
  LAYER M3 ;
        RECT 22.816 20.48 22.848 20.512 ;
  LAYER M1 ;
        RECT 22.88 20.46 22.912 22.968 ;
  LAYER M3 ;
        RECT 22.88 22.916 22.912 22.948 ;
  LAYER M1 ;
        RECT 22.944 20.46 22.976 22.968 ;
  LAYER M3 ;
        RECT 22.944 20.48 22.976 20.512 ;
  LAYER M1 ;
        RECT 23.008 20.46 23.04 22.968 ;
  LAYER M3 ;
        RECT 23.008 22.916 23.04 22.948 ;
  LAYER M1 ;
        RECT 23.072 20.46 23.104 22.968 ;
  LAYER M3 ;
        RECT 23.072 20.48 23.104 20.512 ;
  LAYER M1 ;
        RECT 23.136 20.46 23.168 22.968 ;
  LAYER M3 ;
        RECT 23.136 22.916 23.168 22.948 ;
  LAYER M1 ;
        RECT 23.2 20.46 23.232 22.968 ;
  LAYER M3 ;
        RECT 23.2 20.48 23.232 20.512 ;
  LAYER M1 ;
        RECT 23.264 20.46 23.296 22.968 ;
  LAYER M3 ;
        RECT 23.264 22.916 23.296 22.948 ;
  LAYER M1 ;
        RECT 23.328 20.46 23.36 22.968 ;
  LAYER M3 ;
        RECT 23.328 20.48 23.36 20.512 ;
  LAYER M1 ;
        RECT 23.392 20.46 23.424 22.968 ;
  LAYER M3 ;
        RECT 23.392 22.916 23.424 22.948 ;
  LAYER M1 ;
        RECT 23.456 20.46 23.488 22.968 ;
  LAYER M3 ;
        RECT 23.456 20.48 23.488 20.512 ;
  LAYER M1 ;
        RECT 23.52 20.46 23.552 22.968 ;
  LAYER M3 ;
        RECT 23.52 22.916 23.552 22.948 ;
  LAYER M1 ;
        RECT 23.584 20.46 23.616 22.968 ;
  LAYER M3 ;
        RECT 23.584 20.48 23.616 20.512 ;
  LAYER M1 ;
        RECT 23.648 20.46 23.68 22.968 ;
  LAYER M3 ;
        RECT 23.648 22.916 23.68 22.948 ;
  LAYER M1 ;
        RECT 23.712 20.46 23.744 22.968 ;
  LAYER M3 ;
        RECT 23.712 20.48 23.744 20.512 ;
  LAYER M1 ;
        RECT 23.776 20.46 23.808 22.968 ;
  LAYER M3 ;
        RECT 23.776 22.916 23.808 22.948 ;
  LAYER M1 ;
        RECT 23.84 20.46 23.872 22.968 ;
  LAYER M3 ;
        RECT 23.84 20.48 23.872 20.512 ;
  LAYER M1 ;
        RECT 23.904 20.46 23.936 22.968 ;
  LAYER M3 ;
        RECT 23.904 22.916 23.936 22.948 ;
  LAYER M1 ;
        RECT 23.968 20.46 24 22.968 ;
  LAYER M3 ;
        RECT 23.968 20.48 24 20.512 ;
  LAYER M1 ;
        RECT 24.032 20.46 24.064 22.968 ;
  LAYER M3 ;
        RECT 24.032 22.916 24.064 22.948 ;
  LAYER M1 ;
        RECT 24.096 20.46 24.128 22.968 ;
  LAYER M3 ;
        RECT 24.096 20.48 24.128 20.512 ;
  LAYER M1 ;
        RECT 24.16 20.46 24.192 22.968 ;
  LAYER M3 ;
        RECT 24.16 22.916 24.192 22.948 ;
  LAYER M1 ;
        RECT 24.224 20.46 24.256 22.968 ;
  LAYER M3 ;
        RECT 24.224 20.48 24.256 20.512 ;
  LAYER M1 ;
        RECT 24.288 20.46 24.32 22.968 ;
  LAYER M3 ;
        RECT 24.288 22.916 24.32 22.948 ;
  LAYER M1 ;
        RECT 24.352 20.46 24.384 22.968 ;
  LAYER M3 ;
        RECT 24.352 20.48 24.384 20.512 ;
  LAYER M1 ;
        RECT 24.416 20.46 24.448 22.968 ;
  LAYER M3 ;
        RECT 24.416 22.916 24.448 22.948 ;
  LAYER M1 ;
        RECT 24.48 20.46 24.512 22.968 ;
  LAYER M3 ;
        RECT 24.48 20.48 24.512 20.512 ;
  LAYER M1 ;
        RECT 24.544 20.46 24.576 22.968 ;
  LAYER M3 ;
        RECT 24.544 22.916 24.576 22.948 ;
  LAYER M1 ;
        RECT 24.608 20.46 24.64 22.968 ;
  LAYER M3 ;
        RECT 24.608 20.48 24.64 20.512 ;
  LAYER M1 ;
        RECT 24.672 20.46 24.704 22.968 ;
  LAYER M3 ;
        RECT 24.672 22.916 24.704 22.948 ;
  LAYER M1 ;
        RECT 24.736 20.46 24.768 22.968 ;
  LAYER M3 ;
        RECT 24.736 20.48 24.768 20.512 ;
  LAYER M1 ;
        RECT 24.8 20.46 24.832 22.968 ;
  LAYER M3 ;
        RECT 24.8 22.916 24.832 22.948 ;
  LAYER M1 ;
        RECT 24.864 20.46 24.896 22.968 ;
  LAYER M3 ;
        RECT 24.864 20.48 24.896 20.512 ;
  LAYER M1 ;
        RECT 24.928 20.46 24.96 22.968 ;
  LAYER M3 ;
        RECT 22.56 22.852 22.592 22.884 ;
  LAYER M2 ;
        RECT 24.928 22.788 24.96 22.82 ;
  LAYER M2 ;
        RECT 22.56 22.724 22.592 22.756 ;
  LAYER M2 ;
        RECT 24.928 22.66 24.96 22.692 ;
  LAYER M2 ;
        RECT 22.56 22.596 22.592 22.628 ;
  LAYER M2 ;
        RECT 24.928 22.532 24.96 22.564 ;
  LAYER M2 ;
        RECT 22.56 22.468 22.592 22.5 ;
  LAYER M2 ;
        RECT 24.928 22.404 24.96 22.436 ;
  LAYER M2 ;
        RECT 22.56 22.34 22.592 22.372 ;
  LAYER M2 ;
        RECT 24.928 22.276 24.96 22.308 ;
  LAYER M2 ;
        RECT 22.56 22.212 22.592 22.244 ;
  LAYER M2 ;
        RECT 24.928 22.148 24.96 22.18 ;
  LAYER M2 ;
        RECT 22.56 22.084 22.592 22.116 ;
  LAYER M2 ;
        RECT 24.928 22.02 24.96 22.052 ;
  LAYER M2 ;
        RECT 22.56 21.956 22.592 21.988 ;
  LAYER M2 ;
        RECT 24.928 21.892 24.96 21.924 ;
  LAYER M2 ;
        RECT 22.56 21.828 22.592 21.86 ;
  LAYER M2 ;
        RECT 24.928 21.764 24.96 21.796 ;
  LAYER M2 ;
        RECT 22.56 21.7 22.592 21.732 ;
  LAYER M2 ;
        RECT 24.928 21.636 24.96 21.668 ;
  LAYER M2 ;
        RECT 22.56 21.572 22.592 21.604 ;
  LAYER M2 ;
        RECT 24.928 21.508 24.96 21.54 ;
  LAYER M2 ;
        RECT 22.56 21.444 22.592 21.476 ;
  LAYER M2 ;
        RECT 24.928 21.38 24.96 21.412 ;
  LAYER M2 ;
        RECT 22.56 21.316 22.592 21.348 ;
  LAYER M2 ;
        RECT 24.928 21.252 24.96 21.284 ;
  LAYER M2 ;
        RECT 22.56 21.188 22.592 21.22 ;
  LAYER M2 ;
        RECT 24.928 21.124 24.96 21.156 ;
  LAYER M2 ;
        RECT 22.56 21.06 22.592 21.092 ;
  LAYER M2 ;
        RECT 24.928 20.996 24.96 21.028 ;
  LAYER M2 ;
        RECT 22.56 20.932 22.592 20.964 ;
  LAYER M2 ;
        RECT 24.928 20.868 24.96 20.9 ;
  LAYER M2 ;
        RECT 22.56 20.804 22.592 20.836 ;
  LAYER M2 ;
        RECT 24.928 20.74 24.96 20.772 ;
  LAYER M2 ;
        RECT 22.56 20.676 22.592 20.708 ;
  LAYER M2 ;
        RECT 24.928 20.612 24.96 20.644 ;
  LAYER M2 ;
        RECT 22.512 20.412 25.008 23.016 ;
  LAYER M1 ;
        RECT 25.536 36 25.568 38.508 ;
  LAYER M3 ;
        RECT 25.536 36.02 25.568 36.052 ;
  LAYER M1 ;
        RECT 25.6 36 25.632 38.508 ;
  LAYER M3 ;
        RECT 25.6 38.456 25.632 38.488 ;
  LAYER M1 ;
        RECT 25.664 36 25.696 38.508 ;
  LAYER M3 ;
        RECT 25.664 36.02 25.696 36.052 ;
  LAYER M1 ;
        RECT 25.728 36 25.76 38.508 ;
  LAYER M3 ;
        RECT 25.728 38.456 25.76 38.488 ;
  LAYER M1 ;
        RECT 25.792 36 25.824 38.508 ;
  LAYER M3 ;
        RECT 25.792 36.02 25.824 36.052 ;
  LAYER M1 ;
        RECT 25.856 36 25.888 38.508 ;
  LAYER M3 ;
        RECT 25.856 38.456 25.888 38.488 ;
  LAYER M1 ;
        RECT 25.92 36 25.952 38.508 ;
  LAYER M3 ;
        RECT 25.92 36.02 25.952 36.052 ;
  LAYER M1 ;
        RECT 25.984 36 26.016 38.508 ;
  LAYER M3 ;
        RECT 25.984 38.456 26.016 38.488 ;
  LAYER M1 ;
        RECT 26.048 36 26.08 38.508 ;
  LAYER M3 ;
        RECT 26.048 36.02 26.08 36.052 ;
  LAYER M1 ;
        RECT 26.112 36 26.144 38.508 ;
  LAYER M3 ;
        RECT 26.112 38.456 26.144 38.488 ;
  LAYER M1 ;
        RECT 26.176 36 26.208 38.508 ;
  LAYER M3 ;
        RECT 26.176 36.02 26.208 36.052 ;
  LAYER M1 ;
        RECT 26.24 36 26.272 38.508 ;
  LAYER M3 ;
        RECT 26.24 38.456 26.272 38.488 ;
  LAYER M1 ;
        RECT 26.304 36 26.336 38.508 ;
  LAYER M3 ;
        RECT 26.304 36.02 26.336 36.052 ;
  LAYER M1 ;
        RECT 26.368 36 26.4 38.508 ;
  LAYER M3 ;
        RECT 26.368 38.456 26.4 38.488 ;
  LAYER M1 ;
        RECT 26.432 36 26.464 38.508 ;
  LAYER M3 ;
        RECT 26.432 36.02 26.464 36.052 ;
  LAYER M1 ;
        RECT 26.496 36 26.528 38.508 ;
  LAYER M3 ;
        RECT 26.496 38.456 26.528 38.488 ;
  LAYER M1 ;
        RECT 26.56 36 26.592 38.508 ;
  LAYER M3 ;
        RECT 26.56 36.02 26.592 36.052 ;
  LAYER M1 ;
        RECT 26.624 36 26.656 38.508 ;
  LAYER M3 ;
        RECT 26.624 38.456 26.656 38.488 ;
  LAYER M1 ;
        RECT 26.688 36 26.72 38.508 ;
  LAYER M3 ;
        RECT 26.688 36.02 26.72 36.052 ;
  LAYER M1 ;
        RECT 26.752 36 26.784 38.508 ;
  LAYER M3 ;
        RECT 26.752 38.456 26.784 38.488 ;
  LAYER M1 ;
        RECT 26.816 36 26.848 38.508 ;
  LAYER M3 ;
        RECT 26.816 36.02 26.848 36.052 ;
  LAYER M1 ;
        RECT 26.88 36 26.912 38.508 ;
  LAYER M3 ;
        RECT 26.88 38.456 26.912 38.488 ;
  LAYER M1 ;
        RECT 26.944 36 26.976 38.508 ;
  LAYER M3 ;
        RECT 26.944 36.02 26.976 36.052 ;
  LAYER M1 ;
        RECT 27.008 36 27.04 38.508 ;
  LAYER M3 ;
        RECT 27.008 38.456 27.04 38.488 ;
  LAYER M1 ;
        RECT 27.072 36 27.104 38.508 ;
  LAYER M3 ;
        RECT 27.072 36.02 27.104 36.052 ;
  LAYER M1 ;
        RECT 27.136 36 27.168 38.508 ;
  LAYER M3 ;
        RECT 27.136 38.456 27.168 38.488 ;
  LAYER M1 ;
        RECT 27.2 36 27.232 38.508 ;
  LAYER M3 ;
        RECT 27.2 36.02 27.232 36.052 ;
  LAYER M1 ;
        RECT 27.264 36 27.296 38.508 ;
  LAYER M3 ;
        RECT 27.264 38.456 27.296 38.488 ;
  LAYER M1 ;
        RECT 27.328 36 27.36 38.508 ;
  LAYER M3 ;
        RECT 27.328 36.02 27.36 36.052 ;
  LAYER M1 ;
        RECT 27.392 36 27.424 38.508 ;
  LAYER M3 ;
        RECT 27.392 38.456 27.424 38.488 ;
  LAYER M1 ;
        RECT 27.456 36 27.488 38.508 ;
  LAYER M3 ;
        RECT 27.456 36.02 27.488 36.052 ;
  LAYER M1 ;
        RECT 27.52 36 27.552 38.508 ;
  LAYER M3 ;
        RECT 27.52 38.456 27.552 38.488 ;
  LAYER M1 ;
        RECT 27.584 36 27.616 38.508 ;
  LAYER M3 ;
        RECT 27.584 36.02 27.616 36.052 ;
  LAYER M1 ;
        RECT 27.648 36 27.68 38.508 ;
  LAYER M3 ;
        RECT 27.648 38.456 27.68 38.488 ;
  LAYER M1 ;
        RECT 27.712 36 27.744 38.508 ;
  LAYER M3 ;
        RECT 27.712 36.02 27.744 36.052 ;
  LAYER M1 ;
        RECT 27.776 36 27.808 38.508 ;
  LAYER M3 ;
        RECT 27.776 38.456 27.808 38.488 ;
  LAYER M1 ;
        RECT 27.84 36 27.872 38.508 ;
  LAYER M3 ;
        RECT 27.84 36.02 27.872 36.052 ;
  LAYER M1 ;
        RECT 27.904 36 27.936 38.508 ;
  LAYER M3 ;
        RECT 25.536 38.392 25.568 38.424 ;
  LAYER M2 ;
        RECT 27.904 38.328 27.936 38.36 ;
  LAYER M2 ;
        RECT 25.536 38.264 25.568 38.296 ;
  LAYER M2 ;
        RECT 27.904 38.2 27.936 38.232 ;
  LAYER M2 ;
        RECT 25.536 38.136 25.568 38.168 ;
  LAYER M2 ;
        RECT 27.904 38.072 27.936 38.104 ;
  LAYER M2 ;
        RECT 25.536 38.008 25.568 38.04 ;
  LAYER M2 ;
        RECT 27.904 37.944 27.936 37.976 ;
  LAYER M2 ;
        RECT 25.536 37.88 25.568 37.912 ;
  LAYER M2 ;
        RECT 27.904 37.816 27.936 37.848 ;
  LAYER M2 ;
        RECT 25.536 37.752 25.568 37.784 ;
  LAYER M2 ;
        RECT 27.904 37.688 27.936 37.72 ;
  LAYER M2 ;
        RECT 25.536 37.624 25.568 37.656 ;
  LAYER M2 ;
        RECT 27.904 37.56 27.936 37.592 ;
  LAYER M2 ;
        RECT 25.536 37.496 25.568 37.528 ;
  LAYER M2 ;
        RECT 27.904 37.432 27.936 37.464 ;
  LAYER M2 ;
        RECT 25.536 37.368 25.568 37.4 ;
  LAYER M2 ;
        RECT 27.904 37.304 27.936 37.336 ;
  LAYER M2 ;
        RECT 25.536 37.24 25.568 37.272 ;
  LAYER M2 ;
        RECT 27.904 37.176 27.936 37.208 ;
  LAYER M2 ;
        RECT 25.536 37.112 25.568 37.144 ;
  LAYER M2 ;
        RECT 27.904 37.048 27.936 37.08 ;
  LAYER M2 ;
        RECT 25.536 36.984 25.568 37.016 ;
  LAYER M2 ;
        RECT 27.904 36.92 27.936 36.952 ;
  LAYER M2 ;
        RECT 25.536 36.856 25.568 36.888 ;
  LAYER M2 ;
        RECT 27.904 36.792 27.936 36.824 ;
  LAYER M2 ;
        RECT 25.536 36.728 25.568 36.76 ;
  LAYER M2 ;
        RECT 27.904 36.664 27.936 36.696 ;
  LAYER M2 ;
        RECT 25.536 36.6 25.568 36.632 ;
  LAYER M2 ;
        RECT 27.904 36.536 27.936 36.568 ;
  LAYER M2 ;
        RECT 25.536 36.472 25.568 36.504 ;
  LAYER M2 ;
        RECT 27.904 36.408 27.936 36.44 ;
  LAYER M2 ;
        RECT 25.536 36.344 25.568 36.376 ;
  LAYER M2 ;
        RECT 27.904 36.28 27.936 36.312 ;
  LAYER M2 ;
        RECT 25.536 36.216 25.568 36.248 ;
  LAYER M2 ;
        RECT 27.904 36.152 27.936 36.184 ;
  LAYER M2 ;
        RECT 25.488 35.952 27.984 38.556 ;
  LAYER M1 ;
        RECT 25.536 32.892 25.568 35.4 ;
  LAYER M3 ;
        RECT 25.536 32.912 25.568 32.944 ;
  LAYER M1 ;
        RECT 25.6 32.892 25.632 35.4 ;
  LAYER M3 ;
        RECT 25.6 35.348 25.632 35.38 ;
  LAYER M1 ;
        RECT 25.664 32.892 25.696 35.4 ;
  LAYER M3 ;
        RECT 25.664 32.912 25.696 32.944 ;
  LAYER M1 ;
        RECT 25.728 32.892 25.76 35.4 ;
  LAYER M3 ;
        RECT 25.728 35.348 25.76 35.38 ;
  LAYER M1 ;
        RECT 25.792 32.892 25.824 35.4 ;
  LAYER M3 ;
        RECT 25.792 32.912 25.824 32.944 ;
  LAYER M1 ;
        RECT 25.856 32.892 25.888 35.4 ;
  LAYER M3 ;
        RECT 25.856 35.348 25.888 35.38 ;
  LAYER M1 ;
        RECT 25.92 32.892 25.952 35.4 ;
  LAYER M3 ;
        RECT 25.92 32.912 25.952 32.944 ;
  LAYER M1 ;
        RECT 25.984 32.892 26.016 35.4 ;
  LAYER M3 ;
        RECT 25.984 35.348 26.016 35.38 ;
  LAYER M1 ;
        RECT 26.048 32.892 26.08 35.4 ;
  LAYER M3 ;
        RECT 26.048 32.912 26.08 32.944 ;
  LAYER M1 ;
        RECT 26.112 32.892 26.144 35.4 ;
  LAYER M3 ;
        RECT 26.112 35.348 26.144 35.38 ;
  LAYER M1 ;
        RECT 26.176 32.892 26.208 35.4 ;
  LAYER M3 ;
        RECT 26.176 32.912 26.208 32.944 ;
  LAYER M1 ;
        RECT 26.24 32.892 26.272 35.4 ;
  LAYER M3 ;
        RECT 26.24 35.348 26.272 35.38 ;
  LAYER M1 ;
        RECT 26.304 32.892 26.336 35.4 ;
  LAYER M3 ;
        RECT 26.304 32.912 26.336 32.944 ;
  LAYER M1 ;
        RECT 26.368 32.892 26.4 35.4 ;
  LAYER M3 ;
        RECT 26.368 35.348 26.4 35.38 ;
  LAYER M1 ;
        RECT 26.432 32.892 26.464 35.4 ;
  LAYER M3 ;
        RECT 26.432 32.912 26.464 32.944 ;
  LAYER M1 ;
        RECT 26.496 32.892 26.528 35.4 ;
  LAYER M3 ;
        RECT 26.496 35.348 26.528 35.38 ;
  LAYER M1 ;
        RECT 26.56 32.892 26.592 35.4 ;
  LAYER M3 ;
        RECT 26.56 32.912 26.592 32.944 ;
  LAYER M1 ;
        RECT 26.624 32.892 26.656 35.4 ;
  LAYER M3 ;
        RECT 26.624 35.348 26.656 35.38 ;
  LAYER M1 ;
        RECT 26.688 32.892 26.72 35.4 ;
  LAYER M3 ;
        RECT 26.688 32.912 26.72 32.944 ;
  LAYER M1 ;
        RECT 26.752 32.892 26.784 35.4 ;
  LAYER M3 ;
        RECT 26.752 35.348 26.784 35.38 ;
  LAYER M1 ;
        RECT 26.816 32.892 26.848 35.4 ;
  LAYER M3 ;
        RECT 26.816 32.912 26.848 32.944 ;
  LAYER M1 ;
        RECT 26.88 32.892 26.912 35.4 ;
  LAYER M3 ;
        RECT 26.88 35.348 26.912 35.38 ;
  LAYER M1 ;
        RECT 26.944 32.892 26.976 35.4 ;
  LAYER M3 ;
        RECT 26.944 32.912 26.976 32.944 ;
  LAYER M1 ;
        RECT 27.008 32.892 27.04 35.4 ;
  LAYER M3 ;
        RECT 27.008 35.348 27.04 35.38 ;
  LAYER M1 ;
        RECT 27.072 32.892 27.104 35.4 ;
  LAYER M3 ;
        RECT 27.072 32.912 27.104 32.944 ;
  LAYER M1 ;
        RECT 27.136 32.892 27.168 35.4 ;
  LAYER M3 ;
        RECT 27.136 35.348 27.168 35.38 ;
  LAYER M1 ;
        RECT 27.2 32.892 27.232 35.4 ;
  LAYER M3 ;
        RECT 27.2 32.912 27.232 32.944 ;
  LAYER M1 ;
        RECT 27.264 32.892 27.296 35.4 ;
  LAYER M3 ;
        RECT 27.264 35.348 27.296 35.38 ;
  LAYER M1 ;
        RECT 27.328 32.892 27.36 35.4 ;
  LAYER M3 ;
        RECT 27.328 32.912 27.36 32.944 ;
  LAYER M1 ;
        RECT 27.392 32.892 27.424 35.4 ;
  LAYER M3 ;
        RECT 27.392 35.348 27.424 35.38 ;
  LAYER M1 ;
        RECT 27.456 32.892 27.488 35.4 ;
  LAYER M3 ;
        RECT 27.456 32.912 27.488 32.944 ;
  LAYER M1 ;
        RECT 27.52 32.892 27.552 35.4 ;
  LAYER M3 ;
        RECT 27.52 35.348 27.552 35.38 ;
  LAYER M1 ;
        RECT 27.584 32.892 27.616 35.4 ;
  LAYER M3 ;
        RECT 27.584 32.912 27.616 32.944 ;
  LAYER M1 ;
        RECT 27.648 32.892 27.68 35.4 ;
  LAYER M3 ;
        RECT 27.648 35.348 27.68 35.38 ;
  LAYER M1 ;
        RECT 27.712 32.892 27.744 35.4 ;
  LAYER M3 ;
        RECT 27.712 32.912 27.744 32.944 ;
  LAYER M1 ;
        RECT 27.776 32.892 27.808 35.4 ;
  LAYER M3 ;
        RECT 27.776 35.348 27.808 35.38 ;
  LAYER M1 ;
        RECT 27.84 32.892 27.872 35.4 ;
  LAYER M3 ;
        RECT 27.84 32.912 27.872 32.944 ;
  LAYER M1 ;
        RECT 27.904 32.892 27.936 35.4 ;
  LAYER M3 ;
        RECT 25.536 35.284 25.568 35.316 ;
  LAYER M2 ;
        RECT 27.904 35.22 27.936 35.252 ;
  LAYER M2 ;
        RECT 25.536 35.156 25.568 35.188 ;
  LAYER M2 ;
        RECT 27.904 35.092 27.936 35.124 ;
  LAYER M2 ;
        RECT 25.536 35.028 25.568 35.06 ;
  LAYER M2 ;
        RECT 27.904 34.964 27.936 34.996 ;
  LAYER M2 ;
        RECT 25.536 34.9 25.568 34.932 ;
  LAYER M2 ;
        RECT 27.904 34.836 27.936 34.868 ;
  LAYER M2 ;
        RECT 25.536 34.772 25.568 34.804 ;
  LAYER M2 ;
        RECT 27.904 34.708 27.936 34.74 ;
  LAYER M2 ;
        RECT 25.536 34.644 25.568 34.676 ;
  LAYER M2 ;
        RECT 27.904 34.58 27.936 34.612 ;
  LAYER M2 ;
        RECT 25.536 34.516 25.568 34.548 ;
  LAYER M2 ;
        RECT 27.904 34.452 27.936 34.484 ;
  LAYER M2 ;
        RECT 25.536 34.388 25.568 34.42 ;
  LAYER M2 ;
        RECT 27.904 34.324 27.936 34.356 ;
  LAYER M2 ;
        RECT 25.536 34.26 25.568 34.292 ;
  LAYER M2 ;
        RECT 27.904 34.196 27.936 34.228 ;
  LAYER M2 ;
        RECT 25.536 34.132 25.568 34.164 ;
  LAYER M2 ;
        RECT 27.904 34.068 27.936 34.1 ;
  LAYER M2 ;
        RECT 25.536 34.004 25.568 34.036 ;
  LAYER M2 ;
        RECT 27.904 33.94 27.936 33.972 ;
  LAYER M2 ;
        RECT 25.536 33.876 25.568 33.908 ;
  LAYER M2 ;
        RECT 27.904 33.812 27.936 33.844 ;
  LAYER M2 ;
        RECT 25.536 33.748 25.568 33.78 ;
  LAYER M2 ;
        RECT 27.904 33.684 27.936 33.716 ;
  LAYER M2 ;
        RECT 25.536 33.62 25.568 33.652 ;
  LAYER M2 ;
        RECT 27.904 33.556 27.936 33.588 ;
  LAYER M2 ;
        RECT 25.536 33.492 25.568 33.524 ;
  LAYER M2 ;
        RECT 27.904 33.428 27.936 33.46 ;
  LAYER M2 ;
        RECT 25.536 33.364 25.568 33.396 ;
  LAYER M2 ;
        RECT 27.904 33.3 27.936 33.332 ;
  LAYER M2 ;
        RECT 25.536 33.236 25.568 33.268 ;
  LAYER M2 ;
        RECT 27.904 33.172 27.936 33.204 ;
  LAYER M2 ;
        RECT 25.536 33.108 25.568 33.14 ;
  LAYER M2 ;
        RECT 27.904 33.044 27.936 33.076 ;
  LAYER M2 ;
        RECT 25.488 32.844 27.984 35.448 ;
  LAYER M1 ;
        RECT 25.536 29.784 25.568 32.292 ;
  LAYER M3 ;
        RECT 25.536 29.804 25.568 29.836 ;
  LAYER M1 ;
        RECT 25.6 29.784 25.632 32.292 ;
  LAYER M3 ;
        RECT 25.6 32.24 25.632 32.272 ;
  LAYER M1 ;
        RECT 25.664 29.784 25.696 32.292 ;
  LAYER M3 ;
        RECT 25.664 29.804 25.696 29.836 ;
  LAYER M1 ;
        RECT 25.728 29.784 25.76 32.292 ;
  LAYER M3 ;
        RECT 25.728 32.24 25.76 32.272 ;
  LAYER M1 ;
        RECT 25.792 29.784 25.824 32.292 ;
  LAYER M3 ;
        RECT 25.792 29.804 25.824 29.836 ;
  LAYER M1 ;
        RECT 25.856 29.784 25.888 32.292 ;
  LAYER M3 ;
        RECT 25.856 32.24 25.888 32.272 ;
  LAYER M1 ;
        RECT 25.92 29.784 25.952 32.292 ;
  LAYER M3 ;
        RECT 25.92 29.804 25.952 29.836 ;
  LAYER M1 ;
        RECT 25.984 29.784 26.016 32.292 ;
  LAYER M3 ;
        RECT 25.984 32.24 26.016 32.272 ;
  LAYER M1 ;
        RECT 26.048 29.784 26.08 32.292 ;
  LAYER M3 ;
        RECT 26.048 29.804 26.08 29.836 ;
  LAYER M1 ;
        RECT 26.112 29.784 26.144 32.292 ;
  LAYER M3 ;
        RECT 26.112 32.24 26.144 32.272 ;
  LAYER M1 ;
        RECT 26.176 29.784 26.208 32.292 ;
  LAYER M3 ;
        RECT 26.176 29.804 26.208 29.836 ;
  LAYER M1 ;
        RECT 26.24 29.784 26.272 32.292 ;
  LAYER M3 ;
        RECT 26.24 32.24 26.272 32.272 ;
  LAYER M1 ;
        RECT 26.304 29.784 26.336 32.292 ;
  LAYER M3 ;
        RECT 26.304 29.804 26.336 29.836 ;
  LAYER M1 ;
        RECT 26.368 29.784 26.4 32.292 ;
  LAYER M3 ;
        RECT 26.368 32.24 26.4 32.272 ;
  LAYER M1 ;
        RECT 26.432 29.784 26.464 32.292 ;
  LAYER M3 ;
        RECT 26.432 29.804 26.464 29.836 ;
  LAYER M1 ;
        RECT 26.496 29.784 26.528 32.292 ;
  LAYER M3 ;
        RECT 26.496 32.24 26.528 32.272 ;
  LAYER M1 ;
        RECT 26.56 29.784 26.592 32.292 ;
  LAYER M3 ;
        RECT 26.56 29.804 26.592 29.836 ;
  LAYER M1 ;
        RECT 26.624 29.784 26.656 32.292 ;
  LAYER M3 ;
        RECT 26.624 32.24 26.656 32.272 ;
  LAYER M1 ;
        RECT 26.688 29.784 26.72 32.292 ;
  LAYER M3 ;
        RECT 26.688 29.804 26.72 29.836 ;
  LAYER M1 ;
        RECT 26.752 29.784 26.784 32.292 ;
  LAYER M3 ;
        RECT 26.752 32.24 26.784 32.272 ;
  LAYER M1 ;
        RECT 26.816 29.784 26.848 32.292 ;
  LAYER M3 ;
        RECT 26.816 29.804 26.848 29.836 ;
  LAYER M1 ;
        RECT 26.88 29.784 26.912 32.292 ;
  LAYER M3 ;
        RECT 26.88 32.24 26.912 32.272 ;
  LAYER M1 ;
        RECT 26.944 29.784 26.976 32.292 ;
  LAYER M3 ;
        RECT 26.944 29.804 26.976 29.836 ;
  LAYER M1 ;
        RECT 27.008 29.784 27.04 32.292 ;
  LAYER M3 ;
        RECT 27.008 32.24 27.04 32.272 ;
  LAYER M1 ;
        RECT 27.072 29.784 27.104 32.292 ;
  LAYER M3 ;
        RECT 27.072 29.804 27.104 29.836 ;
  LAYER M1 ;
        RECT 27.136 29.784 27.168 32.292 ;
  LAYER M3 ;
        RECT 27.136 32.24 27.168 32.272 ;
  LAYER M1 ;
        RECT 27.2 29.784 27.232 32.292 ;
  LAYER M3 ;
        RECT 27.2 29.804 27.232 29.836 ;
  LAYER M1 ;
        RECT 27.264 29.784 27.296 32.292 ;
  LAYER M3 ;
        RECT 27.264 32.24 27.296 32.272 ;
  LAYER M1 ;
        RECT 27.328 29.784 27.36 32.292 ;
  LAYER M3 ;
        RECT 27.328 29.804 27.36 29.836 ;
  LAYER M1 ;
        RECT 27.392 29.784 27.424 32.292 ;
  LAYER M3 ;
        RECT 27.392 32.24 27.424 32.272 ;
  LAYER M1 ;
        RECT 27.456 29.784 27.488 32.292 ;
  LAYER M3 ;
        RECT 27.456 29.804 27.488 29.836 ;
  LAYER M1 ;
        RECT 27.52 29.784 27.552 32.292 ;
  LAYER M3 ;
        RECT 27.52 32.24 27.552 32.272 ;
  LAYER M1 ;
        RECT 27.584 29.784 27.616 32.292 ;
  LAYER M3 ;
        RECT 27.584 29.804 27.616 29.836 ;
  LAYER M1 ;
        RECT 27.648 29.784 27.68 32.292 ;
  LAYER M3 ;
        RECT 27.648 32.24 27.68 32.272 ;
  LAYER M1 ;
        RECT 27.712 29.784 27.744 32.292 ;
  LAYER M3 ;
        RECT 27.712 29.804 27.744 29.836 ;
  LAYER M1 ;
        RECT 27.776 29.784 27.808 32.292 ;
  LAYER M3 ;
        RECT 27.776 32.24 27.808 32.272 ;
  LAYER M1 ;
        RECT 27.84 29.784 27.872 32.292 ;
  LAYER M3 ;
        RECT 27.84 29.804 27.872 29.836 ;
  LAYER M1 ;
        RECT 27.904 29.784 27.936 32.292 ;
  LAYER M3 ;
        RECT 25.536 32.176 25.568 32.208 ;
  LAYER M2 ;
        RECT 27.904 32.112 27.936 32.144 ;
  LAYER M2 ;
        RECT 25.536 32.048 25.568 32.08 ;
  LAYER M2 ;
        RECT 27.904 31.984 27.936 32.016 ;
  LAYER M2 ;
        RECT 25.536 31.92 25.568 31.952 ;
  LAYER M2 ;
        RECT 27.904 31.856 27.936 31.888 ;
  LAYER M2 ;
        RECT 25.536 31.792 25.568 31.824 ;
  LAYER M2 ;
        RECT 27.904 31.728 27.936 31.76 ;
  LAYER M2 ;
        RECT 25.536 31.664 25.568 31.696 ;
  LAYER M2 ;
        RECT 27.904 31.6 27.936 31.632 ;
  LAYER M2 ;
        RECT 25.536 31.536 25.568 31.568 ;
  LAYER M2 ;
        RECT 27.904 31.472 27.936 31.504 ;
  LAYER M2 ;
        RECT 25.536 31.408 25.568 31.44 ;
  LAYER M2 ;
        RECT 27.904 31.344 27.936 31.376 ;
  LAYER M2 ;
        RECT 25.536 31.28 25.568 31.312 ;
  LAYER M2 ;
        RECT 27.904 31.216 27.936 31.248 ;
  LAYER M2 ;
        RECT 25.536 31.152 25.568 31.184 ;
  LAYER M2 ;
        RECT 27.904 31.088 27.936 31.12 ;
  LAYER M2 ;
        RECT 25.536 31.024 25.568 31.056 ;
  LAYER M2 ;
        RECT 27.904 30.96 27.936 30.992 ;
  LAYER M2 ;
        RECT 25.536 30.896 25.568 30.928 ;
  LAYER M2 ;
        RECT 27.904 30.832 27.936 30.864 ;
  LAYER M2 ;
        RECT 25.536 30.768 25.568 30.8 ;
  LAYER M2 ;
        RECT 27.904 30.704 27.936 30.736 ;
  LAYER M2 ;
        RECT 25.536 30.64 25.568 30.672 ;
  LAYER M2 ;
        RECT 27.904 30.576 27.936 30.608 ;
  LAYER M2 ;
        RECT 25.536 30.512 25.568 30.544 ;
  LAYER M2 ;
        RECT 27.904 30.448 27.936 30.48 ;
  LAYER M2 ;
        RECT 25.536 30.384 25.568 30.416 ;
  LAYER M2 ;
        RECT 27.904 30.32 27.936 30.352 ;
  LAYER M2 ;
        RECT 25.536 30.256 25.568 30.288 ;
  LAYER M2 ;
        RECT 27.904 30.192 27.936 30.224 ;
  LAYER M2 ;
        RECT 25.536 30.128 25.568 30.16 ;
  LAYER M2 ;
        RECT 27.904 30.064 27.936 30.096 ;
  LAYER M2 ;
        RECT 25.536 30 25.568 30.032 ;
  LAYER M2 ;
        RECT 27.904 29.936 27.936 29.968 ;
  LAYER M2 ;
        RECT 25.488 29.736 27.984 32.34 ;
  LAYER M1 ;
        RECT 25.536 26.676 25.568 29.184 ;
  LAYER M3 ;
        RECT 25.536 26.696 25.568 26.728 ;
  LAYER M1 ;
        RECT 25.6 26.676 25.632 29.184 ;
  LAYER M3 ;
        RECT 25.6 29.132 25.632 29.164 ;
  LAYER M1 ;
        RECT 25.664 26.676 25.696 29.184 ;
  LAYER M3 ;
        RECT 25.664 26.696 25.696 26.728 ;
  LAYER M1 ;
        RECT 25.728 26.676 25.76 29.184 ;
  LAYER M3 ;
        RECT 25.728 29.132 25.76 29.164 ;
  LAYER M1 ;
        RECT 25.792 26.676 25.824 29.184 ;
  LAYER M3 ;
        RECT 25.792 26.696 25.824 26.728 ;
  LAYER M1 ;
        RECT 25.856 26.676 25.888 29.184 ;
  LAYER M3 ;
        RECT 25.856 29.132 25.888 29.164 ;
  LAYER M1 ;
        RECT 25.92 26.676 25.952 29.184 ;
  LAYER M3 ;
        RECT 25.92 26.696 25.952 26.728 ;
  LAYER M1 ;
        RECT 25.984 26.676 26.016 29.184 ;
  LAYER M3 ;
        RECT 25.984 29.132 26.016 29.164 ;
  LAYER M1 ;
        RECT 26.048 26.676 26.08 29.184 ;
  LAYER M3 ;
        RECT 26.048 26.696 26.08 26.728 ;
  LAYER M1 ;
        RECT 26.112 26.676 26.144 29.184 ;
  LAYER M3 ;
        RECT 26.112 29.132 26.144 29.164 ;
  LAYER M1 ;
        RECT 26.176 26.676 26.208 29.184 ;
  LAYER M3 ;
        RECT 26.176 26.696 26.208 26.728 ;
  LAYER M1 ;
        RECT 26.24 26.676 26.272 29.184 ;
  LAYER M3 ;
        RECT 26.24 29.132 26.272 29.164 ;
  LAYER M1 ;
        RECT 26.304 26.676 26.336 29.184 ;
  LAYER M3 ;
        RECT 26.304 26.696 26.336 26.728 ;
  LAYER M1 ;
        RECT 26.368 26.676 26.4 29.184 ;
  LAYER M3 ;
        RECT 26.368 29.132 26.4 29.164 ;
  LAYER M1 ;
        RECT 26.432 26.676 26.464 29.184 ;
  LAYER M3 ;
        RECT 26.432 26.696 26.464 26.728 ;
  LAYER M1 ;
        RECT 26.496 26.676 26.528 29.184 ;
  LAYER M3 ;
        RECT 26.496 29.132 26.528 29.164 ;
  LAYER M1 ;
        RECT 26.56 26.676 26.592 29.184 ;
  LAYER M3 ;
        RECT 26.56 26.696 26.592 26.728 ;
  LAYER M1 ;
        RECT 26.624 26.676 26.656 29.184 ;
  LAYER M3 ;
        RECT 26.624 29.132 26.656 29.164 ;
  LAYER M1 ;
        RECT 26.688 26.676 26.72 29.184 ;
  LAYER M3 ;
        RECT 26.688 26.696 26.72 26.728 ;
  LAYER M1 ;
        RECT 26.752 26.676 26.784 29.184 ;
  LAYER M3 ;
        RECT 26.752 29.132 26.784 29.164 ;
  LAYER M1 ;
        RECT 26.816 26.676 26.848 29.184 ;
  LAYER M3 ;
        RECT 26.816 26.696 26.848 26.728 ;
  LAYER M1 ;
        RECT 26.88 26.676 26.912 29.184 ;
  LAYER M3 ;
        RECT 26.88 29.132 26.912 29.164 ;
  LAYER M1 ;
        RECT 26.944 26.676 26.976 29.184 ;
  LAYER M3 ;
        RECT 26.944 26.696 26.976 26.728 ;
  LAYER M1 ;
        RECT 27.008 26.676 27.04 29.184 ;
  LAYER M3 ;
        RECT 27.008 29.132 27.04 29.164 ;
  LAYER M1 ;
        RECT 27.072 26.676 27.104 29.184 ;
  LAYER M3 ;
        RECT 27.072 26.696 27.104 26.728 ;
  LAYER M1 ;
        RECT 27.136 26.676 27.168 29.184 ;
  LAYER M3 ;
        RECT 27.136 29.132 27.168 29.164 ;
  LAYER M1 ;
        RECT 27.2 26.676 27.232 29.184 ;
  LAYER M3 ;
        RECT 27.2 26.696 27.232 26.728 ;
  LAYER M1 ;
        RECT 27.264 26.676 27.296 29.184 ;
  LAYER M3 ;
        RECT 27.264 29.132 27.296 29.164 ;
  LAYER M1 ;
        RECT 27.328 26.676 27.36 29.184 ;
  LAYER M3 ;
        RECT 27.328 26.696 27.36 26.728 ;
  LAYER M1 ;
        RECT 27.392 26.676 27.424 29.184 ;
  LAYER M3 ;
        RECT 27.392 29.132 27.424 29.164 ;
  LAYER M1 ;
        RECT 27.456 26.676 27.488 29.184 ;
  LAYER M3 ;
        RECT 27.456 26.696 27.488 26.728 ;
  LAYER M1 ;
        RECT 27.52 26.676 27.552 29.184 ;
  LAYER M3 ;
        RECT 27.52 29.132 27.552 29.164 ;
  LAYER M1 ;
        RECT 27.584 26.676 27.616 29.184 ;
  LAYER M3 ;
        RECT 27.584 26.696 27.616 26.728 ;
  LAYER M1 ;
        RECT 27.648 26.676 27.68 29.184 ;
  LAYER M3 ;
        RECT 27.648 29.132 27.68 29.164 ;
  LAYER M1 ;
        RECT 27.712 26.676 27.744 29.184 ;
  LAYER M3 ;
        RECT 27.712 26.696 27.744 26.728 ;
  LAYER M1 ;
        RECT 27.776 26.676 27.808 29.184 ;
  LAYER M3 ;
        RECT 27.776 29.132 27.808 29.164 ;
  LAYER M1 ;
        RECT 27.84 26.676 27.872 29.184 ;
  LAYER M3 ;
        RECT 27.84 26.696 27.872 26.728 ;
  LAYER M1 ;
        RECT 27.904 26.676 27.936 29.184 ;
  LAYER M3 ;
        RECT 25.536 29.068 25.568 29.1 ;
  LAYER M2 ;
        RECT 27.904 29.004 27.936 29.036 ;
  LAYER M2 ;
        RECT 25.536 28.94 25.568 28.972 ;
  LAYER M2 ;
        RECT 27.904 28.876 27.936 28.908 ;
  LAYER M2 ;
        RECT 25.536 28.812 25.568 28.844 ;
  LAYER M2 ;
        RECT 27.904 28.748 27.936 28.78 ;
  LAYER M2 ;
        RECT 25.536 28.684 25.568 28.716 ;
  LAYER M2 ;
        RECT 27.904 28.62 27.936 28.652 ;
  LAYER M2 ;
        RECT 25.536 28.556 25.568 28.588 ;
  LAYER M2 ;
        RECT 27.904 28.492 27.936 28.524 ;
  LAYER M2 ;
        RECT 25.536 28.428 25.568 28.46 ;
  LAYER M2 ;
        RECT 27.904 28.364 27.936 28.396 ;
  LAYER M2 ;
        RECT 25.536 28.3 25.568 28.332 ;
  LAYER M2 ;
        RECT 27.904 28.236 27.936 28.268 ;
  LAYER M2 ;
        RECT 25.536 28.172 25.568 28.204 ;
  LAYER M2 ;
        RECT 27.904 28.108 27.936 28.14 ;
  LAYER M2 ;
        RECT 25.536 28.044 25.568 28.076 ;
  LAYER M2 ;
        RECT 27.904 27.98 27.936 28.012 ;
  LAYER M2 ;
        RECT 25.536 27.916 25.568 27.948 ;
  LAYER M2 ;
        RECT 27.904 27.852 27.936 27.884 ;
  LAYER M2 ;
        RECT 25.536 27.788 25.568 27.82 ;
  LAYER M2 ;
        RECT 27.904 27.724 27.936 27.756 ;
  LAYER M2 ;
        RECT 25.536 27.66 25.568 27.692 ;
  LAYER M2 ;
        RECT 27.904 27.596 27.936 27.628 ;
  LAYER M2 ;
        RECT 25.536 27.532 25.568 27.564 ;
  LAYER M2 ;
        RECT 27.904 27.468 27.936 27.5 ;
  LAYER M2 ;
        RECT 25.536 27.404 25.568 27.436 ;
  LAYER M2 ;
        RECT 27.904 27.34 27.936 27.372 ;
  LAYER M2 ;
        RECT 25.536 27.276 25.568 27.308 ;
  LAYER M2 ;
        RECT 27.904 27.212 27.936 27.244 ;
  LAYER M2 ;
        RECT 25.536 27.148 25.568 27.18 ;
  LAYER M2 ;
        RECT 27.904 27.084 27.936 27.116 ;
  LAYER M2 ;
        RECT 25.536 27.02 25.568 27.052 ;
  LAYER M2 ;
        RECT 27.904 26.956 27.936 26.988 ;
  LAYER M2 ;
        RECT 25.536 26.892 25.568 26.924 ;
  LAYER M2 ;
        RECT 27.904 26.828 27.936 26.86 ;
  LAYER M2 ;
        RECT 25.488 26.628 27.984 29.232 ;
  LAYER M1 ;
        RECT 25.536 23.568 25.568 26.076 ;
  LAYER M3 ;
        RECT 25.536 23.588 25.568 23.62 ;
  LAYER M1 ;
        RECT 25.6 23.568 25.632 26.076 ;
  LAYER M3 ;
        RECT 25.6 26.024 25.632 26.056 ;
  LAYER M1 ;
        RECT 25.664 23.568 25.696 26.076 ;
  LAYER M3 ;
        RECT 25.664 23.588 25.696 23.62 ;
  LAYER M1 ;
        RECT 25.728 23.568 25.76 26.076 ;
  LAYER M3 ;
        RECT 25.728 26.024 25.76 26.056 ;
  LAYER M1 ;
        RECT 25.792 23.568 25.824 26.076 ;
  LAYER M3 ;
        RECT 25.792 23.588 25.824 23.62 ;
  LAYER M1 ;
        RECT 25.856 23.568 25.888 26.076 ;
  LAYER M3 ;
        RECT 25.856 26.024 25.888 26.056 ;
  LAYER M1 ;
        RECT 25.92 23.568 25.952 26.076 ;
  LAYER M3 ;
        RECT 25.92 23.588 25.952 23.62 ;
  LAYER M1 ;
        RECT 25.984 23.568 26.016 26.076 ;
  LAYER M3 ;
        RECT 25.984 26.024 26.016 26.056 ;
  LAYER M1 ;
        RECT 26.048 23.568 26.08 26.076 ;
  LAYER M3 ;
        RECT 26.048 23.588 26.08 23.62 ;
  LAYER M1 ;
        RECT 26.112 23.568 26.144 26.076 ;
  LAYER M3 ;
        RECT 26.112 26.024 26.144 26.056 ;
  LAYER M1 ;
        RECT 26.176 23.568 26.208 26.076 ;
  LAYER M3 ;
        RECT 26.176 23.588 26.208 23.62 ;
  LAYER M1 ;
        RECT 26.24 23.568 26.272 26.076 ;
  LAYER M3 ;
        RECT 26.24 26.024 26.272 26.056 ;
  LAYER M1 ;
        RECT 26.304 23.568 26.336 26.076 ;
  LAYER M3 ;
        RECT 26.304 23.588 26.336 23.62 ;
  LAYER M1 ;
        RECT 26.368 23.568 26.4 26.076 ;
  LAYER M3 ;
        RECT 26.368 26.024 26.4 26.056 ;
  LAYER M1 ;
        RECT 26.432 23.568 26.464 26.076 ;
  LAYER M3 ;
        RECT 26.432 23.588 26.464 23.62 ;
  LAYER M1 ;
        RECT 26.496 23.568 26.528 26.076 ;
  LAYER M3 ;
        RECT 26.496 26.024 26.528 26.056 ;
  LAYER M1 ;
        RECT 26.56 23.568 26.592 26.076 ;
  LAYER M3 ;
        RECT 26.56 23.588 26.592 23.62 ;
  LAYER M1 ;
        RECT 26.624 23.568 26.656 26.076 ;
  LAYER M3 ;
        RECT 26.624 26.024 26.656 26.056 ;
  LAYER M1 ;
        RECT 26.688 23.568 26.72 26.076 ;
  LAYER M3 ;
        RECT 26.688 23.588 26.72 23.62 ;
  LAYER M1 ;
        RECT 26.752 23.568 26.784 26.076 ;
  LAYER M3 ;
        RECT 26.752 26.024 26.784 26.056 ;
  LAYER M1 ;
        RECT 26.816 23.568 26.848 26.076 ;
  LAYER M3 ;
        RECT 26.816 23.588 26.848 23.62 ;
  LAYER M1 ;
        RECT 26.88 23.568 26.912 26.076 ;
  LAYER M3 ;
        RECT 26.88 26.024 26.912 26.056 ;
  LAYER M1 ;
        RECT 26.944 23.568 26.976 26.076 ;
  LAYER M3 ;
        RECT 26.944 23.588 26.976 23.62 ;
  LAYER M1 ;
        RECT 27.008 23.568 27.04 26.076 ;
  LAYER M3 ;
        RECT 27.008 26.024 27.04 26.056 ;
  LAYER M1 ;
        RECT 27.072 23.568 27.104 26.076 ;
  LAYER M3 ;
        RECT 27.072 23.588 27.104 23.62 ;
  LAYER M1 ;
        RECT 27.136 23.568 27.168 26.076 ;
  LAYER M3 ;
        RECT 27.136 26.024 27.168 26.056 ;
  LAYER M1 ;
        RECT 27.2 23.568 27.232 26.076 ;
  LAYER M3 ;
        RECT 27.2 23.588 27.232 23.62 ;
  LAYER M1 ;
        RECT 27.264 23.568 27.296 26.076 ;
  LAYER M3 ;
        RECT 27.264 26.024 27.296 26.056 ;
  LAYER M1 ;
        RECT 27.328 23.568 27.36 26.076 ;
  LAYER M3 ;
        RECT 27.328 23.588 27.36 23.62 ;
  LAYER M1 ;
        RECT 27.392 23.568 27.424 26.076 ;
  LAYER M3 ;
        RECT 27.392 26.024 27.424 26.056 ;
  LAYER M1 ;
        RECT 27.456 23.568 27.488 26.076 ;
  LAYER M3 ;
        RECT 27.456 23.588 27.488 23.62 ;
  LAYER M1 ;
        RECT 27.52 23.568 27.552 26.076 ;
  LAYER M3 ;
        RECT 27.52 26.024 27.552 26.056 ;
  LAYER M1 ;
        RECT 27.584 23.568 27.616 26.076 ;
  LAYER M3 ;
        RECT 27.584 23.588 27.616 23.62 ;
  LAYER M1 ;
        RECT 27.648 23.568 27.68 26.076 ;
  LAYER M3 ;
        RECT 27.648 26.024 27.68 26.056 ;
  LAYER M1 ;
        RECT 27.712 23.568 27.744 26.076 ;
  LAYER M3 ;
        RECT 27.712 23.588 27.744 23.62 ;
  LAYER M1 ;
        RECT 27.776 23.568 27.808 26.076 ;
  LAYER M3 ;
        RECT 27.776 26.024 27.808 26.056 ;
  LAYER M1 ;
        RECT 27.84 23.568 27.872 26.076 ;
  LAYER M3 ;
        RECT 27.84 23.588 27.872 23.62 ;
  LAYER M1 ;
        RECT 27.904 23.568 27.936 26.076 ;
  LAYER M3 ;
        RECT 25.536 25.96 25.568 25.992 ;
  LAYER M2 ;
        RECT 27.904 25.896 27.936 25.928 ;
  LAYER M2 ;
        RECT 25.536 25.832 25.568 25.864 ;
  LAYER M2 ;
        RECT 27.904 25.768 27.936 25.8 ;
  LAYER M2 ;
        RECT 25.536 25.704 25.568 25.736 ;
  LAYER M2 ;
        RECT 27.904 25.64 27.936 25.672 ;
  LAYER M2 ;
        RECT 25.536 25.576 25.568 25.608 ;
  LAYER M2 ;
        RECT 27.904 25.512 27.936 25.544 ;
  LAYER M2 ;
        RECT 25.536 25.448 25.568 25.48 ;
  LAYER M2 ;
        RECT 27.904 25.384 27.936 25.416 ;
  LAYER M2 ;
        RECT 25.536 25.32 25.568 25.352 ;
  LAYER M2 ;
        RECT 27.904 25.256 27.936 25.288 ;
  LAYER M2 ;
        RECT 25.536 25.192 25.568 25.224 ;
  LAYER M2 ;
        RECT 27.904 25.128 27.936 25.16 ;
  LAYER M2 ;
        RECT 25.536 25.064 25.568 25.096 ;
  LAYER M2 ;
        RECT 27.904 25 27.936 25.032 ;
  LAYER M2 ;
        RECT 25.536 24.936 25.568 24.968 ;
  LAYER M2 ;
        RECT 27.904 24.872 27.936 24.904 ;
  LAYER M2 ;
        RECT 25.536 24.808 25.568 24.84 ;
  LAYER M2 ;
        RECT 27.904 24.744 27.936 24.776 ;
  LAYER M2 ;
        RECT 25.536 24.68 25.568 24.712 ;
  LAYER M2 ;
        RECT 27.904 24.616 27.936 24.648 ;
  LAYER M2 ;
        RECT 25.536 24.552 25.568 24.584 ;
  LAYER M2 ;
        RECT 27.904 24.488 27.936 24.52 ;
  LAYER M2 ;
        RECT 25.536 24.424 25.568 24.456 ;
  LAYER M2 ;
        RECT 27.904 24.36 27.936 24.392 ;
  LAYER M2 ;
        RECT 25.536 24.296 25.568 24.328 ;
  LAYER M2 ;
        RECT 27.904 24.232 27.936 24.264 ;
  LAYER M2 ;
        RECT 25.536 24.168 25.568 24.2 ;
  LAYER M2 ;
        RECT 27.904 24.104 27.936 24.136 ;
  LAYER M2 ;
        RECT 25.536 24.04 25.568 24.072 ;
  LAYER M2 ;
        RECT 27.904 23.976 27.936 24.008 ;
  LAYER M2 ;
        RECT 25.536 23.912 25.568 23.944 ;
  LAYER M2 ;
        RECT 27.904 23.848 27.936 23.88 ;
  LAYER M2 ;
        RECT 25.536 23.784 25.568 23.816 ;
  LAYER M2 ;
        RECT 27.904 23.72 27.936 23.752 ;
  LAYER M2 ;
        RECT 25.488 23.52 27.984 26.124 ;
  LAYER M1 ;
        RECT 25.536 20.46 25.568 22.968 ;
  LAYER M3 ;
        RECT 25.536 20.48 25.568 20.512 ;
  LAYER M1 ;
        RECT 25.6 20.46 25.632 22.968 ;
  LAYER M3 ;
        RECT 25.6 22.916 25.632 22.948 ;
  LAYER M1 ;
        RECT 25.664 20.46 25.696 22.968 ;
  LAYER M3 ;
        RECT 25.664 20.48 25.696 20.512 ;
  LAYER M1 ;
        RECT 25.728 20.46 25.76 22.968 ;
  LAYER M3 ;
        RECT 25.728 22.916 25.76 22.948 ;
  LAYER M1 ;
        RECT 25.792 20.46 25.824 22.968 ;
  LAYER M3 ;
        RECT 25.792 20.48 25.824 20.512 ;
  LAYER M1 ;
        RECT 25.856 20.46 25.888 22.968 ;
  LAYER M3 ;
        RECT 25.856 22.916 25.888 22.948 ;
  LAYER M1 ;
        RECT 25.92 20.46 25.952 22.968 ;
  LAYER M3 ;
        RECT 25.92 20.48 25.952 20.512 ;
  LAYER M1 ;
        RECT 25.984 20.46 26.016 22.968 ;
  LAYER M3 ;
        RECT 25.984 22.916 26.016 22.948 ;
  LAYER M1 ;
        RECT 26.048 20.46 26.08 22.968 ;
  LAYER M3 ;
        RECT 26.048 20.48 26.08 20.512 ;
  LAYER M1 ;
        RECT 26.112 20.46 26.144 22.968 ;
  LAYER M3 ;
        RECT 26.112 22.916 26.144 22.948 ;
  LAYER M1 ;
        RECT 26.176 20.46 26.208 22.968 ;
  LAYER M3 ;
        RECT 26.176 20.48 26.208 20.512 ;
  LAYER M1 ;
        RECT 26.24 20.46 26.272 22.968 ;
  LAYER M3 ;
        RECT 26.24 22.916 26.272 22.948 ;
  LAYER M1 ;
        RECT 26.304 20.46 26.336 22.968 ;
  LAYER M3 ;
        RECT 26.304 20.48 26.336 20.512 ;
  LAYER M1 ;
        RECT 26.368 20.46 26.4 22.968 ;
  LAYER M3 ;
        RECT 26.368 22.916 26.4 22.948 ;
  LAYER M1 ;
        RECT 26.432 20.46 26.464 22.968 ;
  LAYER M3 ;
        RECT 26.432 20.48 26.464 20.512 ;
  LAYER M1 ;
        RECT 26.496 20.46 26.528 22.968 ;
  LAYER M3 ;
        RECT 26.496 22.916 26.528 22.948 ;
  LAYER M1 ;
        RECT 26.56 20.46 26.592 22.968 ;
  LAYER M3 ;
        RECT 26.56 20.48 26.592 20.512 ;
  LAYER M1 ;
        RECT 26.624 20.46 26.656 22.968 ;
  LAYER M3 ;
        RECT 26.624 22.916 26.656 22.948 ;
  LAYER M1 ;
        RECT 26.688 20.46 26.72 22.968 ;
  LAYER M3 ;
        RECT 26.688 20.48 26.72 20.512 ;
  LAYER M1 ;
        RECT 26.752 20.46 26.784 22.968 ;
  LAYER M3 ;
        RECT 26.752 22.916 26.784 22.948 ;
  LAYER M1 ;
        RECT 26.816 20.46 26.848 22.968 ;
  LAYER M3 ;
        RECT 26.816 20.48 26.848 20.512 ;
  LAYER M1 ;
        RECT 26.88 20.46 26.912 22.968 ;
  LAYER M3 ;
        RECT 26.88 22.916 26.912 22.948 ;
  LAYER M1 ;
        RECT 26.944 20.46 26.976 22.968 ;
  LAYER M3 ;
        RECT 26.944 20.48 26.976 20.512 ;
  LAYER M1 ;
        RECT 27.008 20.46 27.04 22.968 ;
  LAYER M3 ;
        RECT 27.008 22.916 27.04 22.948 ;
  LAYER M1 ;
        RECT 27.072 20.46 27.104 22.968 ;
  LAYER M3 ;
        RECT 27.072 20.48 27.104 20.512 ;
  LAYER M1 ;
        RECT 27.136 20.46 27.168 22.968 ;
  LAYER M3 ;
        RECT 27.136 22.916 27.168 22.948 ;
  LAYER M1 ;
        RECT 27.2 20.46 27.232 22.968 ;
  LAYER M3 ;
        RECT 27.2 20.48 27.232 20.512 ;
  LAYER M1 ;
        RECT 27.264 20.46 27.296 22.968 ;
  LAYER M3 ;
        RECT 27.264 22.916 27.296 22.948 ;
  LAYER M1 ;
        RECT 27.328 20.46 27.36 22.968 ;
  LAYER M3 ;
        RECT 27.328 20.48 27.36 20.512 ;
  LAYER M1 ;
        RECT 27.392 20.46 27.424 22.968 ;
  LAYER M3 ;
        RECT 27.392 22.916 27.424 22.948 ;
  LAYER M1 ;
        RECT 27.456 20.46 27.488 22.968 ;
  LAYER M3 ;
        RECT 27.456 20.48 27.488 20.512 ;
  LAYER M1 ;
        RECT 27.52 20.46 27.552 22.968 ;
  LAYER M3 ;
        RECT 27.52 22.916 27.552 22.948 ;
  LAYER M1 ;
        RECT 27.584 20.46 27.616 22.968 ;
  LAYER M3 ;
        RECT 27.584 20.48 27.616 20.512 ;
  LAYER M1 ;
        RECT 27.648 20.46 27.68 22.968 ;
  LAYER M3 ;
        RECT 27.648 22.916 27.68 22.948 ;
  LAYER M1 ;
        RECT 27.712 20.46 27.744 22.968 ;
  LAYER M3 ;
        RECT 27.712 20.48 27.744 20.512 ;
  LAYER M1 ;
        RECT 27.776 20.46 27.808 22.968 ;
  LAYER M3 ;
        RECT 27.776 22.916 27.808 22.948 ;
  LAYER M1 ;
        RECT 27.84 20.46 27.872 22.968 ;
  LAYER M3 ;
        RECT 27.84 20.48 27.872 20.512 ;
  LAYER M1 ;
        RECT 27.904 20.46 27.936 22.968 ;
  LAYER M3 ;
        RECT 25.536 22.852 25.568 22.884 ;
  LAYER M2 ;
        RECT 27.904 22.788 27.936 22.82 ;
  LAYER M2 ;
        RECT 25.536 22.724 25.568 22.756 ;
  LAYER M2 ;
        RECT 27.904 22.66 27.936 22.692 ;
  LAYER M2 ;
        RECT 25.536 22.596 25.568 22.628 ;
  LAYER M2 ;
        RECT 27.904 22.532 27.936 22.564 ;
  LAYER M2 ;
        RECT 25.536 22.468 25.568 22.5 ;
  LAYER M2 ;
        RECT 27.904 22.404 27.936 22.436 ;
  LAYER M2 ;
        RECT 25.536 22.34 25.568 22.372 ;
  LAYER M2 ;
        RECT 27.904 22.276 27.936 22.308 ;
  LAYER M2 ;
        RECT 25.536 22.212 25.568 22.244 ;
  LAYER M2 ;
        RECT 27.904 22.148 27.936 22.18 ;
  LAYER M2 ;
        RECT 25.536 22.084 25.568 22.116 ;
  LAYER M2 ;
        RECT 27.904 22.02 27.936 22.052 ;
  LAYER M2 ;
        RECT 25.536 21.956 25.568 21.988 ;
  LAYER M2 ;
        RECT 27.904 21.892 27.936 21.924 ;
  LAYER M2 ;
        RECT 25.536 21.828 25.568 21.86 ;
  LAYER M2 ;
        RECT 27.904 21.764 27.936 21.796 ;
  LAYER M2 ;
        RECT 25.536 21.7 25.568 21.732 ;
  LAYER M2 ;
        RECT 27.904 21.636 27.936 21.668 ;
  LAYER M2 ;
        RECT 25.536 21.572 25.568 21.604 ;
  LAYER M2 ;
        RECT 27.904 21.508 27.936 21.54 ;
  LAYER M2 ;
        RECT 25.536 21.444 25.568 21.476 ;
  LAYER M2 ;
        RECT 27.904 21.38 27.936 21.412 ;
  LAYER M2 ;
        RECT 25.536 21.316 25.568 21.348 ;
  LAYER M2 ;
        RECT 27.904 21.252 27.936 21.284 ;
  LAYER M2 ;
        RECT 25.536 21.188 25.568 21.22 ;
  LAYER M2 ;
        RECT 27.904 21.124 27.936 21.156 ;
  LAYER M2 ;
        RECT 25.536 21.06 25.568 21.092 ;
  LAYER M2 ;
        RECT 27.904 20.996 27.936 21.028 ;
  LAYER M2 ;
        RECT 25.536 20.932 25.568 20.964 ;
  LAYER M2 ;
        RECT 27.904 20.868 27.936 20.9 ;
  LAYER M2 ;
        RECT 25.536 20.804 25.568 20.836 ;
  LAYER M2 ;
        RECT 27.904 20.74 27.936 20.772 ;
  LAYER M2 ;
        RECT 25.536 20.676 25.568 20.708 ;
  LAYER M2 ;
        RECT 27.904 20.612 27.936 20.644 ;
  LAYER M2 ;
        RECT 25.488 20.412 27.984 23.016 ;
  LAYER M1 ;
        RECT 28.512 36 28.544 38.508 ;
  LAYER M3 ;
        RECT 28.512 36.02 28.544 36.052 ;
  LAYER M1 ;
        RECT 28.576 36 28.608 38.508 ;
  LAYER M3 ;
        RECT 28.576 38.456 28.608 38.488 ;
  LAYER M1 ;
        RECT 28.64 36 28.672 38.508 ;
  LAYER M3 ;
        RECT 28.64 36.02 28.672 36.052 ;
  LAYER M1 ;
        RECT 28.704 36 28.736 38.508 ;
  LAYER M3 ;
        RECT 28.704 38.456 28.736 38.488 ;
  LAYER M1 ;
        RECT 28.768 36 28.8 38.508 ;
  LAYER M3 ;
        RECT 28.768 36.02 28.8 36.052 ;
  LAYER M1 ;
        RECT 28.832 36 28.864 38.508 ;
  LAYER M3 ;
        RECT 28.832 38.456 28.864 38.488 ;
  LAYER M1 ;
        RECT 28.896 36 28.928 38.508 ;
  LAYER M3 ;
        RECT 28.896 36.02 28.928 36.052 ;
  LAYER M1 ;
        RECT 28.96 36 28.992 38.508 ;
  LAYER M3 ;
        RECT 28.96 38.456 28.992 38.488 ;
  LAYER M1 ;
        RECT 29.024 36 29.056 38.508 ;
  LAYER M3 ;
        RECT 29.024 36.02 29.056 36.052 ;
  LAYER M1 ;
        RECT 29.088 36 29.12 38.508 ;
  LAYER M3 ;
        RECT 29.088 38.456 29.12 38.488 ;
  LAYER M1 ;
        RECT 29.152 36 29.184 38.508 ;
  LAYER M3 ;
        RECT 29.152 36.02 29.184 36.052 ;
  LAYER M1 ;
        RECT 29.216 36 29.248 38.508 ;
  LAYER M3 ;
        RECT 29.216 38.456 29.248 38.488 ;
  LAYER M1 ;
        RECT 29.28 36 29.312 38.508 ;
  LAYER M3 ;
        RECT 29.28 36.02 29.312 36.052 ;
  LAYER M1 ;
        RECT 29.344 36 29.376 38.508 ;
  LAYER M3 ;
        RECT 29.344 38.456 29.376 38.488 ;
  LAYER M1 ;
        RECT 29.408 36 29.44 38.508 ;
  LAYER M3 ;
        RECT 29.408 36.02 29.44 36.052 ;
  LAYER M1 ;
        RECT 29.472 36 29.504 38.508 ;
  LAYER M3 ;
        RECT 29.472 38.456 29.504 38.488 ;
  LAYER M1 ;
        RECT 29.536 36 29.568 38.508 ;
  LAYER M3 ;
        RECT 29.536 36.02 29.568 36.052 ;
  LAYER M1 ;
        RECT 29.6 36 29.632 38.508 ;
  LAYER M3 ;
        RECT 29.6 38.456 29.632 38.488 ;
  LAYER M1 ;
        RECT 29.664 36 29.696 38.508 ;
  LAYER M3 ;
        RECT 29.664 36.02 29.696 36.052 ;
  LAYER M1 ;
        RECT 29.728 36 29.76 38.508 ;
  LAYER M3 ;
        RECT 29.728 38.456 29.76 38.488 ;
  LAYER M1 ;
        RECT 29.792 36 29.824 38.508 ;
  LAYER M3 ;
        RECT 29.792 36.02 29.824 36.052 ;
  LAYER M1 ;
        RECT 29.856 36 29.888 38.508 ;
  LAYER M3 ;
        RECT 29.856 38.456 29.888 38.488 ;
  LAYER M1 ;
        RECT 29.92 36 29.952 38.508 ;
  LAYER M3 ;
        RECT 29.92 36.02 29.952 36.052 ;
  LAYER M1 ;
        RECT 29.984 36 30.016 38.508 ;
  LAYER M3 ;
        RECT 29.984 38.456 30.016 38.488 ;
  LAYER M1 ;
        RECT 30.048 36 30.08 38.508 ;
  LAYER M3 ;
        RECT 30.048 36.02 30.08 36.052 ;
  LAYER M1 ;
        RECT 30.112 36 30.144 38.508 ;
  LAYER M3 ;
        RECT 30.112 38.456 30.144 38.488 ;
  LAYER M1 ;
        RECT 30.176 36 30.208 38.508 ;
  LAYER M3 ;
        RECT 30.176 36.02 30.208 36.052 ;
  LAYER M1 ;
        RECT 30.24 36 30.272 38.508 ;
  LAYER M3 ;
        RECT 30.24 38.456 30.272 38.488 ;
  LAYER M1 ;
        RECT 30.304 36 30.336 38.508 ;
  LAYER M3 ;
        RECT 30.304 36.02 30.336 36.052 ;
  LAYER M1 ;
        RECT 30.368 36 30.4 38.508 ;
  LAYER M3 ;
        RECT 30.368 38.456 30.4 38.488 ;
  LAYER M1 ;
        RECT 30.432 36 30.464 38.508 ;
  LAYER M3 ;
        RECT 30.432 36.02 30.464 36.052 ;
  LAYER M1 ;
        RECT 30.496 36 30.528 38.508 ;
  LAYER M3 ;
        RECT 30.496 38.456 30.528 38.488 ;
  LAYER M1 ;
        RECT 30.56 36 30.592 38.508 ;
  LAYER M3 ;
        RECT 30.56 36.02 30.592 36.052 ;
  LAYER M1 ;
        RECT 30.624 36 30.656 38.508 ;
  LAYER M3 ;
        RECT 30.624 38.456 30.656 38.488 ;
  LAYER M1 ;
        RECT 30.688 36 30.72 38.508 ;
  LAYER M3 ;
        RECT 30.688 36.02 30.72 36.052 ;
  LAYER M1 ;
        RECT 30.752 36 30.784 38.508 ;
  LAYER M3 ;
        RECT 30.752 38.456 30.784 38.488 ;
  LAYER M1 ;
        RECT 30.816 36 30.848 38.508 ;
  LAYER M3 ;
        RECT 30.816 36.02 30.848 36.052 ;
  LAYER M1 ;
        RECT 30.88 36 30.912 38.508 ;
  LAYER M3 ;
        RECT 28.512 38.392 28.544 38.424 ;
  LAYER M2 ;
        RECT 30.88 38.328 30.912 38.36 ;
  LAYER M2 ;
        RECT 28.512 38.264 28.544 38.296 ;
  LAYER M2 ;
        RECT 30.88 38.2 30.912 38.232 ;
  LAYER M2 ;
        RECT 28.512 38.136 28.544 38.168 ;
  LAYER M2 ;
        RECT 30.88 38.072 30.912 38.104 ;
  LAYER M2 ;
        RECT 28.512 38.008 28.544 38.04 ;
  LAYER M2 ;
        RECT 30.88 37.944 30.912 37.976 ;
  LAYER M2 ;
        RECT 28.512 37.88 28.544 37.912 ;
  LAYER M2 ;
        RECT 30.88 37.816 30.912 37.848 ;
  LAYER M2 ;
        RECT 28.512 37.752 28.544 37.784 ;
  LAYER M2 ;
        RECT 30.88 37.688 30.912 37.72 ;
  LAYER M2 ;
        RECT 28.512 37.624 28.544 37.656 ;
  LAYER M2 ;
        RECT 30.88 37.56 30.912 37.592 ;
  LAYER M2 ;
        RECT 28.512 37.496 28.544 37.528 ;
  LAYER M2 ;
        RECT 30.88 37.432 30.912 37.464 ;
  LAYER M2 ;
        RECT 28.512 37.368 28.544 37.4 ;
  LAYER M2 ;
        RECT 30.88 37.304 30.912 37.336 ;
  LAYER M2 ;
        RECT 28.512 37.24 28.544 37.272 ;
  LAYER M2 ;
        RECT 30.88 37.176 30.912 37.208 ;
  LAYER M2 ;
        RECT 28.512 37.112 28.544 37.144 ;
  LAYER M2 ;
        RECT 30.88 37.048 30.912 37.08 ;
  LAYER M2 ;
        RECT 28.512 36.984 28.544 37.016 ;
  LAYER M2 ;
        RECT 30.88 36.92 30.912 36.952 ;
  LAYER M2 ;
        RECT 28.512 36.856 28.544 36.888 ;
  LAYER M2 ;
        RECT 30.88 36.792 30.912 36.824 ;
  LAYER M2 ;
        RECT 28.512 36.728 28.544 36.76 ;
  LAYER M2 ;
        RECT 30.88 36.664 30.912 36.696 ;
  LAYER M2 ;
        RECT 28.512 36.6 28.544 36.632 ;
  LAYER M2 ;
        RECT 30.88 36.536 30.912 36.568 ;
  LAYER M2 ;
        RECT 28.512 36.472 28.544 36.504 ;
  LAYER M2 ;
        RECT 30.88 36.408 30.912 36.44 ;
  LAYER M2 ;
        RECT 28.512 36.344 28.544 36.376 ;
  LAYER M2 ;
        RECT 30.88 36.28 30.912 36.312 ;
  LAYER M2 ;
        RECT 28.512 36.216 28.544 36.248 ;
  LAYER M2 ;
        RECT 30.88 36.152 30.912 36.184 ;
  LAYER M2 ;
        RECT 28.464 35.952 30.96 38.556 ;
  LAYER M1 ;
        RECT 28.512 32.892 28.544 35.4 ;
  LAYER M3 ;
        RECT 28.512 32.912 28.544 32.944 ;
  LAYER M1 ;
        RECT 28.576 32.892 28.608 35.4 ;
  LAYER M3 ;
        RECT 28.576 35.348 28.608 35.38 ;
  LAYER M1 ;
        RECT 28.64 32.892 28.672 35.4 ;
  LAYER M3 ;
        RECT 28.64 32.912 28.672 32.944 ;
  LAYER M1 ;
        RECT 28.704 32.892 28.736 35.4 ;
  LAYER M3 ;
        RECT 28.704 35.348 28.736 35.38 ;
  LAYER M1 ;
        RECT 28.768 32.892 28.8 35.4 ;
  LAYER M3 ;
        RECT 28.768 32.912 28.8 32.944 ;
  LAYER M1 ;
        RECT 28.832 32.892 28.864 35.4 ;
  LAYER M3 ;
        RECT 28.832 35.348 28.864 35.38 ;
  LAYER M1 ;
        RECT 28.896 32.892 28.928 35.4 ;
  LAYER M3 ;
        RECT 28.896 32.912 28.928 32.944 ;
  LAYER M1 ;
        RECT 28.96 32.892 28.992 35.4 ;
  LAYER M3 ;
        RECT 28.96 35.348 28.992 35.38 ;
  LAYER M1 ;
        RECT 29.024 32.892 29.056 35.4 ;
  LAYER M3 ;
        RECT 29.024 32.912 29.056 32.944 ;
  LAYER M1 ;
        RECT 29.088 32.892 29.12 35.4 ;
  LAYER M3 ;
        RECT 29.088 35.348 29.12 35.38 ;
  LAYER M1 ;
        RECT 29.152 32.892 29.184 35.4 ;
  LAYER M3 ;
        RECT 29.152 32.912 29.184 32.944 ;
  LAYER M1 ;
        RECT 29.216 32.892 29.248 35.4 ;
  LAYER M3 ;
        RECT 29.216 35.348 29.248 35.38 ;
  LAYER M1 ;
        RECT 29.28 32.892 29.312 35.4 ;
  LAYER M3 ;
        RECT 29.28 32.912 29.312 32.944 ;
  LAYER M1 ;
        RECT 29.344 32.892 29.376 35.4 ;
  LAYER M3 ;
        RECT 29.344 35.348 29.376 35.38 ;
  LAYER M1 ;
        RECT 29.408 32.892 29.44 35.4 ;
  LAYER M3 ;
        RECT 29.408 32.912 29.44 32.944 ;
  LAYER M1 ;
        RECT 29.472 32.892 29.504 35.4 ;
  LAYER M3 ;
        RECT 29.472 35.348 29.504 35.38 ;
  LAYER M1 ;
        RECT 29.536 32.892 29.568 35.4 ;
  LAYER M3 ;
        RECT 29.536 32.912 29.568 32.944 ;
  LAYER M1 ;
        RECT 29.6 32.892 29.632 35.4 ;
  LAYER M3 ;
        RECT 29.6 35.348 29.632 35.38 ;
  LAYER M1 ;
        RECT 29.664 32.892 29.696 35.4 ;
  LAYER M3 ;
        RECT 29.664 32.912 29.696 32.944 ;
  LAYER M1 ;
        RECT 29.728 32.892 29.76 35.4 ;
  LAYER M3 ;
        RECT 29.728 35.348 29.76 35.38 ;
  LAYER M1 ;
        RECT 29.792 32.892 29.824 35.4 ;
  LAYER M3 ;
        RECT 29.792 32.912 29.824 32.944 ;
  LAYER M1 ;
        RECT 29.856 32.892 29.888 35.4 ;
  LAYER M3 ;
        RECT 29.856 35.348 29.888 35.38 ;
  LAYER M1 ;
        RECT 29.92 32.892 29.952 35.4 ;
  LAYER M3 ;
        RECT 29.92 32.912 29.952 32.944 ;
  LAYER M1 ;
        RECT 29.984 32.892 30.016 35.4 ;
  LAYER M3 ;
        RECT 29.984 35.348 30.016 35.38 ;
  LAYER M1 ;
        RECT 30.048 32.892 30.08 35.4 ;
  LAYER M3 ;
        RECT 30.048 32.912 30.08 32.944 ;
  LAYER M1 ;
        RECT 30.112 32.892 30.144 35.4 ;
  LAYER M3 ;
        RECT 30.112 35.348 30.144 35.38 ;
  LAYER M1 ;
        RECT 30.176 32.892 30.208 35.4 ;
  LAYER M3 ;
        RECT 30.176 32.912 30.208 32.944 ;
  LAYER M1 ;
        RECT 30.24 32.892 30.272 35.4 ;
  LAYER M3 ;
        RECT 30.24 35.348 30.272 35.38 ;
  LAYER M1 ;
        RECT 30.304 32.892 30.336 35.4 ;
  LAYER M3 ;
        RECT 30.304 32.912 30.336 32.944 ;
  LAYER M1 ;
        RECT 30.368 32.892 30.4 35.4 ;
  LAYER M3 ;
        RECT 30.368 35.348 30.4 35.38 ;
  LAYER M1 ;
        RECT 30.432 32.892 30.464 35.4 ;
  LAYER M3 ;
        RECT 30.432 32.912 30.464 32.944 ;
  LAYER M1 ;
        RECT 30.496 32.892 30.528 35.4 ;
  LAYER M3 ;
        RECT 30.496 35.348 30.528 35.38 ;
  LAYER M1 ;
        RECT 30.56 32.892 30.592 35.4 ;
  LAYER M3 ;
        RECT 30.56 32.912 30.592 32.944 ;
  LAYER M1 ;
        RECT 30.624 32.892 30.656 35.4 ;
  LAYER M3 ;
        RECT 30.624 35.348 30.656 35.38 ;
  LAYER M1 ;
        RECT 30.688 32.892 30.72 35.4 ;
  LAYER M3 ;
        RECT 30.688 32.912 30.72 32.944 ;
  LAYER M1 ;
        RECT 30.752 32.892 30.784 35.4 ;
  LAYER M3 ;
        RECT 30.752 35.348 30.784 35.38 ;
  LAYER M1 ;
        RECT 30.816 32.892 30.848 35.4 ;
  LAYER M3 ;
        RECT 30.816 32.912 30.848 32.944 ;
  LAYER M1 ;
        RECT 30.88 32.892 30.912 35.4 ;
  LAYER M3 ;
        RECT 28.512 35.284 28.544 35.316 ;
  LAYER M2 ;
        RECT 30.88 35.22 30.912 35.252 ;
  LAYER M2 ;
        RECT 28.512 35.156 28.544 35.188 ;
  LAYER M2 ;
        RECT 30.88 35.092 30.912 35.124 ;
  LAYER M2 ;
        RECT 28.512 35.028 28.544 35.06 ;
  LAYER M2 ;
        RECT 30.88 34.964 30.912 34.996 ;
  LAYER M2 ;
        RECT 28.512 34.9 28.544 34.932 ;
  LAYER M2 ;
        RECT 30.88 34.836 30.912 34.868 ;
  LAYER M2 ;
        RECT 28.512 34.772 28.544 34.804 ;
  LAYER M2 ;
        RECT 30.88 34.708 30.912 34.74 ;
  LAYER M2 ;
        RECT 28.512 34.644 28.544 34.676 ;
  LAYER M2 ;
        RECT 30.88 34.58 30.912 34.612 ;
  LAYER M2 ;
        RECT 28.512 34.516 28.544 34.548 ;
  LAYER M2 ;
        RECT 30.88 34.452 30.912 34.484 ;
  LAYER M2 ;
        RECT 28.512 34.388 28.544 34.42 ;
  LAYER M2 ;
        RECT 30.88 34.324 30.912 34.356 ;
  LAYER M2 ;
        RECT 28.512 34.26 28.544 34.292 ;
  LAYER M2 ;
        RECT 30.88 34.196 30.912 34.228 ;
  LAYER M2 ;
        RECT 28.512 34.132 28.544 34.164 ;
  LAYER M2 ;
        RECT 30.88 34.068 30.912 34.1 ;
  LAYER M2 ;
        RECT 28.512 34.004 28.544 34.036 ;
  LAYER M2 ;
        RECT 30.88 33.94 30.912 33.972 ;
  LAYER M2 ;
        RECT 28.512 33.876 28.544 33.908 ;
  LAYER M2 ;
        RECT 30.88 33.812 30.912 33.844 ;
  LAYER M2 ;
        RECT 28.512 33.748 28.544 33.78 ;
  LAYER M2 ;
        RECT 30.88 33.684 30.912 33.716 ;
  LAYER M2 ;
        RECT 28.512 33.62 28.544 33.652 ;
  LAYER M2 ;
        RECT 30.88 33.556 30.912 33.588 ;
  LAYER M2 ;
        RECT 28.512 33.492 28.544 33.524 ;
  LAYER M2 ;
        RECT 30.88 33.428 30.912 33.46 ;
  LAYER M2 ;
        RECT 28.512 33.364 28.544 33.396 ;
  LAYER M2 ;
        RECT 30.88 33.3 30.912 33.332 ;
  LAYER M2 ;
        RECT 28.512 33.236 28.544 33.268 ;
  LAYER M2 ;
        RECT 30.88 33.172 30.912 33.204 ;
  LAYER M2 ;
        RECT 28.512 33.108 28.544 33.14 ;
  LAYER M2 ;
        RECT 30.88 33.044 30.912 33.076 ;
  LAYER M2 ;
        RECT 28.464 32.844 30.96 35.448 ;
  LAYER M1 ;
        RECT 28.512 29.784 28.544 32.292 ;
  LAYER M3 ;
        RECT 28.512 29.804 28.544 29.836 ;
  LAYER M1 ;
        RECT 28.576 29.784 28.608 32.292 ;
  LAYER M3 ;
        RECT 28.576 32.24 28.608 32.272 ;
  LAYER M1 ;
        RECT 28.64 29.784 28.672 32.292 ;
  LAYER M3 ;
        RECT 28.64 29.804 28.672 29.836 ;
  LAYER M1 ;
        RECT 28.704 29.784 28.736 32.292 ;
  LAYER M3 ;
        RECT 28.704 32.24 28.736 32.272 ;
  LAYER M1 ;
        RECT 28.768 29.784 28.8 32.292 ;
  LAYER M3 ;
        RECT 28.768 29.804 28.8 29.836 ;
  LAYER M1 ;
        RECT 28.832 29.784 28.864 32.292 ;
  LAYER M3 ;
        RECT 28.832 32.24 28.864 32.272 ;
  LAYER M1 ;
        RECT 28.896 29.784 28.928 32.292 ;
  LAYER M3 ;
        RECT 28.896 29.804 28.928 29.836 ;
  LAYER M1 ;
        RECT 28.96 29.784 28.992 32.292 ;
  LAYER M3 ;
        RECT 28.96 32.24 28.992 32.272 ;
  LAYER M1 ;
        RECT 29.024 29.784 29.056 32.292 ;
  LAYER M3 ;
        RECT 29.024 29.804 29.056 29.836 ;
  LAYER M1 ;
        RECT 29.088 29.784 29.12 32.292 ;
  LAYER M3 ;
        RECT 29.088 32.24 29.12 32.272 ;
  LAYER M1 ;
        RECT 29.152 29.784 29.184 32.292 ;
  LAYER M3 ;
        RECT 29.152 29.804 29.184 29.836 ;
  LAYER M1 ;
        RECT 29.216 29.784 29.248 32.292 ;
  LAYER M3 ;
        RECT 29.216 32.24 29.248 32.272 ;
  LAYER M1 ;
        RECT 29.28 29.784 29.312 32.292 ;
  LAYER M3 ;
        RECT 29.28 29.804 29.312 29.836 ;
  LAYER M1 ;
        RECT 29.344 29.784 29.376 32.292 ;
  LAYER M3 ;
        RECT 29.344 32.24 29.376 32.272 ;
  LAYER M1 ;
        RECT 29.408 29.784 29.44 32.292 ;
  LAYER M3 ;
        RECT 29.408 29.804 29.44 29.836 ;
  LAYER M1 ;
        RECT 29.472 29.784 29.504 32.292 ;
  LAYER M3 ;
        RECT 29.472 32.24 29.504 32.272 ;
  LAYER M1 ;
        RECT 29.536 29.784 29.568 32.292 ;
  LAYER M3 ;
        RECT 29.536 29.804 29.568 29.836 ;
  LAYER M1 ;
        RECT 29.6 29.784 29.632 32.292 ;
  LAYER M3 ;
        RECT 29.6 32.24 29.632 32.272 ;
  LAYER M1 ;
        RECT 29.664 29.784 29.696 32.292 ;
  LAYER M3 ;
        RECT 29.664 29.804 29.696 29.836 ;
  LAYER M1 ;
        RECT 29.728 29.784 29.76 32.292 ;
  LAYER M3 ;
        RECT 29.728 32.24 29.76 32.272 ;
  LAYER M1 ;
        RECT 29.792 29.784 29.824 32.292 ;
  LAYER M3 ;
        RECT 29.792 29.804 29.824 29.836 ;
  LAYER M1 ;
        RECT 29.856 29.784 29.888 32.292 ;
  LAYER M3 ;
        RECT 29.856 32.24 29.888 32.272 ;
  LAYER M1 ;
        RECT 29.92 29.784 29.952 32.292 ;
  LAYER M3 ;
        RECT 29.92 29.804 29.952 29.836 ;
  LAYER M1 ;
        RECT 29.984 29.784 30.016 32.292 ;
  LAYER M3 ;
        RECT 29.984 32.24 30.016 32.272 ;
  LAYER M1 ;
        RECT 30.048 29.784 30.08 32.292 ;
  LAYER M3 ;
        RECT 30.048 29.804 30.08 29.836 ;
  LAYER M1 ;
        RECT 30.112 29.784 30.144 32.292 ;
  LAYER M3 ;
        RECT 30.112 32.24 30.144 32.272 ;
  LAYER M1 ;
        RECT 30.176 29.784 30.208 32.292 ;
  LAYER M3 ;
        RECT 30.176 29.804 30.208 29.836 ;
  LAYER M1 ;
        RECT 30.24 29.784 30.272 32.292 ;
  LAYER M3 ;
        RECT 30.24 32.24 30.272 32.272 ;
  LAYER M1 ;
        RECT 30.304 29.784 30.336 32.292 ;
  LAYER M3 ;
        RECT 30.304 29.804 30.336 29.836 ;
  LAYER M1 ;
        RECT 30.368 29.784 30.4 32.292 ;
  LAYER M3 ;
        RECT 30.368 32.24 30.4 32.272 ;
  LAYER M1 ;
        RECT 30.432 29.784 30.464 32.292 ;
  LAYER M3 ;
        RECT 30.432 29.804 30.464 29.836 ;
  LAYER M1 ;
        RECT 30.496 29.784 30.528 32.292 ;
  LAYER M3 ;
        RECT 30.496 32.24 30.528 32.272 ;
  LAYER M1 ;
        RECT 30.56 29.784 30.592 32.292 ;
  LAYER M3 ;
        RECT 30.56 29.804 30.592 29.836 ;
  LAYER M1 ;
        RECT 30.624 29.784 30.656 32.292 ;
  LAYER M3 ;
        RECT 30.624 32.24 30.656 32.272 ;
  LAYER M1 ;
        RECT 30.688 29.784 30.72 32.292 ;
  LAYER M3 ;
        RECT 30.688 29.804 30.72 29.836 ;
  LAYER M1 ;
        RECT 30.752 29.784 30.784 32.292 ;
  LAYER M3 ;
        RECT 30.752 32.24 30.784 32.272 ;
  LAYER M1 ;
        RECT 30.816 29.784 30.848 32.292 ;
  LAYER M3 ;
        RECT 30.816 29.804 30.848 29.836 ;
  LAYER M1 ;
        RECT 30.88 29.784 30.912 32.292 ;
  LAYER M3 ;
        RECT 28.512 32.176 28.544 32.208 ;
  LAYER M2 ;
        RECT 30.88 32.112 30.912 32.144 ;
  LAYER M2 ;
        RECT 28.512 32.048 28.544 32.08 ;
  LAYER M2 ;
        RECT 30.88 31.984 30.912 32.016 ;
  LAYER M2 ;
        RECT 28.512 31.92 28.544 31.952 ;
  LAYER M2 ;
        RECT 30.88 31.856 30.912 31.888 ;
  LAYER M2 ;
        RECT 28.512 31.792 28.544 31.824 ;
  LAYER M2 ;
        RECT 30.88 31.728 30.912 31.76 ;
  LAYER M2 ;
        RECT 28.512 31.664 28.544 31.696 ;
  LAYER M2 ;
        RECT 30.88 31.6 30.912 31.632 ;
  LAYER M2 ;
        RECT 28.512 31.536 28.544 31.568 ;
  LAYER M2 ;
        RECT 30.88 31.472 30.912 31.504 ;
  LAYER M2 ;
        RECT 28.512 31.408 28.544 31.44 ;
  LAYER M2 ;
        RECT 30.88 31.344 30.912 31.376 ;
  LAYER M2 ;
        RECT 28.512 31.28 28.544 31.312 ;
  LAYER M2 ;
        RECT 30.88 31.216 30.912 31.248 ;
  LAYER M2 ;
        RECT 28.512 31.152 28.544 31.184 ;
  LAYER M2 ;
        RECT 30.88 31.088 30.912 31.12 ;
  LAYER M2 ;
        RECT 28.512 31.024 28.544 31.056 ;
  LAYER M2 ;
        RECT 30.88 30.96 30.912 30.992 ;
  LAYER M2 ;
        RECT 28.512 30.896 28.544 30.928 ;
  LAYER M2 ;
        RECT 30.88 30.832 30.912 30.864 ;
  LAYER M2 ;
        RECT 28.512 30.768 28.544 30.8 ;
  LAYER M2 ;
        RECT 30.88 30.704 30.912 30.736 ;
  LAYER M2 ;
        RECT 28.512 30.64 28.544 30.672 ;
  LAYER M2 ;
        RECT 30.88 30.576 30.912 30.608 ;
  LAYER M2 ;
        RECT 28.512 30.512 28.544 30.544 ;
  LAYER M2 ;
        RECT 30.88 30.448 30.912 30.48 ;
  LAYER M2 ;
        RECT 28.512 30.384 28.544 30.416 ;
  LAYER M2 ;
        RECT 30.88 30.32 30.912 30.352 ;
  LAYER M2 ;
        RECT 28.512 30.256 28.544 30.288 ;
  LAYER M2 ;
        RECT 30.88 30.192 30.912 30.224 ;
  LAYER M2 ;
        RECT 28.512 30.128 28.544 30.16 ;
  LAYER M2 ;
        RECT 30.88 30.064 30.912 30.096 ;
  LAYER M2 ;
        RECT 28.512 30 28.544 30.032 ;
  LAYER M2 ;
        RECT 30.88 29.936 30.912 29.968 ;
  LAYER M2 ;
        RECT 28.464 29.736 30.96 32.34 ;
  LAYER M1 ;
        RECT 28.512 26.676 28.544 29.184 ;
  LAYER M3 ;
        RECT 28.512 26.696 28.544 26.728 ;
  LAYER M1 ;
        RECT 28.576 26.676 28.608 29.184 ;
  LAYER M3 ;
        RECT 28.576 29.132 28.608 29.164 ;
  LAYER M1 ;
        RECT 28.64 26.676 28.672 29.184 ;
  LAYER M3 ;
        RECT 28.64 26.696 28.672 26.728 ;
  LAYER M1 ;
        RECT 28.704 26.676 28.736 29.184 ;
  LAYER M3 ;
        RECT 28.704 29.132 28.736 29.164 ;
  LAYER M1 ;
        RECT 28.768 26.676 28.8 29.184 ;
  LAYER M3 ;
        RECT 28.768 26.696 28.8 26.728 ;
  LAYER M1 ;
        RECT 28.832 26.676 28.864 29.184 ;
  LAYER M3 ;
        RECT 28.832 29.132 28.864 29.164 ;
  LAYER M1 ;
        RECT 28.896 26.676 28.928 29.184 ;
  LAYER M3 ;
        RECT 28.896 26.696 28.928 26.728 ;
  LAYER M1 ;
        RECT 28.96 26.676 28.992 29.184 ;
  LAYER M3 ;
        RECT 28.96 29.132 28.992 29.164 ;
  LAYER M1 ;
        RECT 29.024 26.676 29.056 29.184 ;
  LAYER M3 ;
        RECT 29.024 26.696 29.056 26.728 ;
  LAYER M1 ;
        RECT 29.088 26.676 29.12 29.184 ;
  LAYER M3 ;
        RECT 29.088 29.132 29.12 29.164 ;
  LAYER M1 ;
        RECT 29.152 26.676 29.184 29.184 ;
  LAYER M3 ;
        RECT 29.152 26.696 29.184 26.728 ;
  LAYER M1 ;
        RECT 29.216 26.676 29.248 29.184 ;
  LAYER M3 ;
        RECT 29.216 29.132 29.248 29.164 ;
  LAYER M1 ;
        RECT 29.28 26.676 29.312 29.184 ;
  LAYER M3 ;
        RECT 29.28 26.696 29.312 26.728 ;
  LAYER M1 ;
        RECT 29.344 26.676 29.376 29.184 ;
  LAYER M3 ;
        RECT 29.344 29.132 29.376 29.164 ;
  LAYER M1 ;
        RECT 29.408 26.676 29.44 29.184 ;
  LAYER M3 ;
        RECT 29.408 26.696 29.44 26.728 ;
  LAYER M1 ;
        RECT 29.472 26.676 29.504 29.184 ;
  LAYER M3 ;
        RECT 29.472 29.132 29.504 29.164 ;
  LAYER M1 ;
        RECT 29.536 26.676 29.568 29.184 ;
  LAYER M3 ;
        RECT 29.536 26.696 29.568 26.728 ;
  LAYER M1 ;
        RECT 29.6 26.676 29.632 29.184 ;
  LAYER M3 ;
        RECT 29.6 29.132 29.632 29.164 ;
  LAYER M1 ;
        RECT 29.664 26.676 29.696 29.184 ;
  LAYER M3 ;
        RECT 29.664 26.696 29.696 26.728 ;
  LAYER M1 ;
        RECT 29.728 26.676 29.76 29.184 ;
  LAYER M3 ;
        RECT 29.728 29.132 29.76 29.164 ;
  LAYER M1 ;
        RECT 29.792 26.676 29.824 29.184 ;
  LAYER M3 ;
        RECT 29.792 26.696 29.824 26.728 ;
  LAYER M1 ;
        RECT 29.856 26.676 29.888 29.184 ;
  LAYER M3 ;
        RECT 29.856 29.132 29.888 29.164 ;
  LAYER M1 ;
        RECT 29.92 26.676 29.952 29.184 ;
  LAYER M3 ;
        RECT 29.92 26.696 29.952 26.728 ;
  LAYER M1 ;
        RECT 29.984 26.676 30.016 29.184 ;
  LAYER M3 ;
        RECT 29.984 29.132 30.016 29.164 ;
  LAYER M1 ;
        RECT 30.048 26.676 30.08 29.184 ;
  LAYER M3 ;
        RECT 30.048 26.696 30.08 26.728 ;
  LAYER M1 ;
        RECT 30.112 26.676 30.144 29.184 ;
  LAYER M3 ;
        RECT 30.112 29.132 30.144 29.164 ;
  LAYER M1 ;
        RECT 30.176 26.676 30.208 29.184 ;
  LAYER M3 ;
        RECT 30.176 26.696 30.208 26.728 ;
  LAYER M1 ;
        RECT 30.24 26.676 30.272 29.184 ;
  LAYER M3 ;
        RECT 30.24 29.132 30.272 29.164 ;
  LAYER M1 ;
        RECT 30.304 26.676 30.336 29.184 ;
  LAYER M3 ;
        RECT 30.304 26.696 30.336 26.728 ;
  LAYER M1 ;
        RECT 30.368 26.676 30.4 29.184 ;
  LAYER M3 ;
        RECT 30.368 29.132 30.4 29.164 ;
  LAYER M1 ;
        RECT 30.432 26.676 30.464 29.184 ;
  LAYER M3 ;
        RECT 30.432 26.696 30.464 26.728 ;
  LAYER M1 ;
        RECT 30.496 26.676 30.528 29.184 ;
  LAYER M3 ;
        RECT 30.496 29.132 30.528 29.164 ;
  LAYER M1 ;
        RECT 30.56 26.676 30.592 29.184 ;
  LAYER M3 ;
        RECT 30.56 26.696 30.592 26.728 ;
  LAYER M1 ;
        RECT 30.624 26.676 30.656 29.184 ;
  LAYER M3 ;
        RECT 30.624 29.132 30.656 29.164 ;
  LAYER M1 ;
        RECT 30.688 26.676 30.72 29.184 ;
  LAYER M3 ;
        RECT 30.688 26.696 30.72 26.728 ;
  LAYER M1 ;
        RECT 30.752 26.676 30.784 29.184 ;
  LAYER M3 ;
        RECT 30.752 29.132 30.784 29.164 ;
  LAYER M1 ;
        RECT 30.816 26.676 30.848 29.184 ;
  LAYER M3 ;
        RECT 30.816 26.696 30.848 26.728 ;
  LAYER M1 ;
        RECT 30.88 26.676 30.912 29.184 ;
  LAYER M3 ;
        RECT 28.512 29.068 28.544 29.1 ;
  LAYER M2 ;
        RECT 30.88 29.004 30.912 29.036 ;
  LAYER M2 ;
        RECT 28.512 28.94 28.544 28.972 ;
  LAYER M2 ;
        RECT 30.88 28.876 30.912 28.908 ;
  LAYER M2 ;
        RECT 28.512 28.812 28.544 28.844 ;
  LAYER M2 ;
        RECT 30.88 28.748 30.912 28.78 ;
  LAYER M2 ;
        RECT 28.512 28.684 28.544 28.716 ;
  LAYER M2 ;
        RECT 30.88 28.62 30.912 28.652 ;
  LAYER M2 ;
        RECT 28.512 28.556 28.544 28.588 ;
  LAYER M2 ;
        RECT 30.88 28.492 30.912 28.524 ;
  LAYER M2 ;
        RECT 28.512 28.428 28.544 28.46 ;
  LAYER M2 ;
        RECT 30.88 28.364 30.912 28.396 ;
  LAYER M2 ;
        RECT 28.512 28.3 28.544 28.332 ;
  LAYER M2 ;
        RECT 30.88 28.236 30.912 28.268 ;
  LAYER M2 ;
        RECT 28.512 28.172 28.544 28.204 ;
  LAYER M2 ;
        RECT 30.88 28.108 30.912 28.14 ;
  LAYER M2 ;
        RECT 28.512 28.044 28.544 28.076 ;
  LAYER M2 ;
        RECT 30.88 27.98 30.912 28.012 ;
  LAYER M2 ;
        RECT 28.512 27.916 28.544 27.948 ;
  LAYER M2 ;
        RECT 30.88 27.852 30.912 27.884 ;
  LAYER M2 ;
        RECT 28.512 27.788 28.544 27.82 ;
  LAYER M2 ;
        RECT 30.88 27.724 30.912 27.756 ;
  LAYER M2 ;
        RECT 28.512 27.66 28.544 27.692 ;
  LAYER M2 ;
        RECT 30.88 27.596 30.912 27.628 ;
  LAYER M2 ;
        RECT 28.512 27.532 28.544 27.564 ;
  LAYER M2 ;
        RECT 30.88 27.468 30.912 27.5 ;
  LAYER M2 ;
        RECT 28.512 27.404 28.544 27.436 ;
  LAYER M2 ;
        RECT 30.88 27.34 30.912 27.372 ;
  LAYER M2 ;
        RECT 28.512 27.276 28.544 27.308 ;
  LAYER M2 ;
        RECT 30.88 27.212 30.912 27.244 ;
  LAYER M2 ;
        RECT 28.512 27.148 28.544 27.18 ;
  LAYER M2 ;
        RECT 30.88 27.084 30.912 27.116 ;
  LAYER M2 ;
        RECT 28.512 27.02 28.544 27.052 ;
  LAYER M2 ;
        RECT 30.88 26.956 30.912 26.988 ;
  LAYER M2 ;
        RECT 28.512 26.892 28.544 26.924 ;
  LAYER M2 ;
        RECT 30.88 26.828 30.912 26.86 ;
  LAYER M2 ;
        RECT 28.464 26.628 30.96 29.232 ;
  LAYER M1 ;
        RECT 28.512 23.568 28.544 26.076 ;
  LAYER M3 ;
        RECT 28.512 23.588 28.544 23.62 ;
  LAYER M1 ;
        RECT 28.576 23.568 28.608 26.076 ;
  LAYER M3 ;
        RECT 28.576 26.024 28.608 26.056 ;
  LAYER M1 ;
        RECT 28.64 23.568 28.672 26.076 ;
  LAYER M3 ;
        RECT 28.64 23.588 28.672 23.62 ;
  LAYER M1 ;
        RECT 28.704 23.568 28.736 26.076 ;
  LAYER M3 ;
        RECT 28.704 26.024 28.736 26.056 ;
  LAYER M1 ;
        RECT 28.768 23.568 28.8 26.076 ;
  LAYER M3 ;
        RECT 28.768 23.588 28.8 23.62 ;
  LAYER M1 ;
        RECT 28.832 23.568 28.864 26.076 ;
  LAYER M3 ;
        RECT 28.832 26.024 28.864 26.056 ;
  LAYER M1 ;
        RECT 28.896 23.568 28.928 26.076 ;
  LAYER M3 ;
        RECT 28.896 23.588 28.928 23.62 ;
  LAYER M1 ;
        RECT 28.96 23.568 28.992 26.076 ;
  LAYER M3 ;
        RECT 28.96 26.024 28.992 26.056 ;
  LAYER M1 ;
        RECT 29.024 23.568 29.056 26.076 ;
  LAYER M3 ;
        RECT 29.024 23.588 29.056 23.62 ;
  LAYER M1 ;
        RECT 29.088 23.568 29.12 26.076 ;
  LAYER M3 ;
        RECT 29.088 26.024 29.12 26.056 ;
  LAYER M1 ;
        RECT 29.152 23.568 29.184 26.076 ;
  LAYER M3 ;
        RECT 29.152 23.588 29.184 23.62 ;
  LAYER M1 ;
        RECT 29.216 23.568 29.248 26.076 ;
  LAYER M3 ;
        RECT 29.216 26.024 29.248 26.056 ;
  LAYER M1 ;
        RECT 29.28 23.568 29.312 26.076 ;
  LAYER M3 ;
        RECT 29.28 23.588 29.312 23.62 ;
  LAYER M1 ;
        RECT 29.344 23.568 29.376 26.076 ;
  LAYER M3 ;
        RECT 29.344 26.024 29.376 26.056 ;
  LAYER M1 ;
        RECT 29.408 23.568 29.44 26.076 ;
  LAYER M3 ;
        RECT 29.408 23.588 29.44 23.62 ;
  LAYER M1 ;
        RECT 29.472 23.568 29.504 26.076 ;
  LAYER M3 ;
        RECT 29.472 26.024 29.504 26.056 ;
  LAYER M1 ;
        RECT 29.536 23.568 29.568 26.076 ;
  LAYER M3 ;
        RECT 29.536 23.588 29.568 23.62 ;
  LAYER M1 ;
        RECT 29.6 23.568 29.632 26.076 ;
  LAYER M3 ;
        RECT 29.6 26.024 29.632 26.056 ;
  LAYER M1 ;
        RECT 29.664 23.568 29.696 26.076 ;
  LAYER M3 ;
        RECT 29.664 23.588 29.696 23.62 ;
  LAYER M1 ;
        RECT 29.728 23.568 29.76 26.076 ;
  LAYER M3 ;
        RECT 29.728 26.024 29.76 26.056 ;
  LAYER M1 ;
        RECT 29.792 23.568 29.824 26.076 ;
  LAYER M3 ;
        RECT 29.792 23.588 29.824 23.62 ;
  LAYER M1 ;
        RECT 29.856 23.568 29.888 26.076 ;
  LAYER M3 ;
        RECT 29.856 26.024 29.888 26.056 ;
  LAYER M1 ;
        RECT 29.92 23.568 29.952 26.076 ;
  LAYER M3 ;
        RECT 29.92 23.588 29.952 23.62 ;
  LAYER M1 ;
        RECT 29.984 23.568 30.016 26.076 ;
  LAYER M3 ;
        RECT 29.984 26.024 30.016 26.056 ;
  LAYER M1 ;
        RECT 30.048 23.568 30.08 26.076 ;
  LAYER M3 ;
        RECT 30.048 23.588 30.08 23.62 ;
  LAYER M1 ;
        RECT 30.112 23.568 30.144 26.076 ;
  LAYER M3 ;
        RECT 30.112 26.024 30.144 26.056 ;
  LAYER M1 ;
        RECT 30.176 23.568 30.208 26.076 ;
  LAYER M3 ;
        RECT 30.176 23.588 30.208 23.62 ;
  LAYER M1 ;
        RECT 30.24 23.568 30.272 26.076 ;
  LAYER M3 ;
        RECT 30.24 26.024 30.272 26.056 ;
  LAYER M1 ;
        RECT 30.304 23.568 30.336 26.076 ;
  LAYER M3 ;
        RECT 30.304 23.588 30.336 23.62 ;
  LAYER M1 ;
        RECT 30.368 23.568 30.4 26.076 ;
  LAYER M3 ;
        RECT 30.368 26.024 30.4 26.056 ;
  LAYER M1 ;
        RECT 30.432 23.568 30.464 26.076 ;
  LAYER M3 ;
        RECT 30.432 23.588 30.464 23.62 ;
  LAYER M1 ;
        RECT 30.496 23.568 30.528 26.076 ;
  LAYER M3 ;
        RECT 30.496 26.024 30.528 26.056 ;
  LAYER M1 ;
        RECT 30.56 23.568 30.592 26.076 ;
  LAYER M3 ;
        RECT 30.56 23.588 30.592 23.62 ;
  LAYER M1 ;
        RECT 30.624 23.568 30.656 26.076 ;
  LAYER M3 ;
        RECT 30.624 26.024 30.656 26.056 ;
  LAYER M1 ;
        RECT 30.688 23.568 30.72 26.076 ;
  LAYER M3 ;
        RECT 30.688 23.588 30.72 23.62 ;
  LAYER M1 ;
        RECT 30.752 23.568 30.784 26.076 ;
  LAYER M3 ;
        RECT 30.752 26.024 30.784 26.056 ;
  LAYER M1 ;
        RECT 30.816 23.568 30.848 26.076 ;
  LAYER M3 ;
        RECT 30.816 23.588 30.848 23.62 ;
  LAYER M1 ;
        RECT 30.88 23.568 30.912 26.076 ;
  LAYER M3 ;
        RECT 28.512 25.96 28.544 25.992 ;
  LAYER M2 ;
        RECT 30.88 25.896 30.912 25.928 ;
  LAYER M2 ;
        RECT 28.512 25.832 28.544 25.864 ;
  LAYER M2 ;
        RECT 30.88 25.768 30.912 25.8 ;
  LAYER M2 ;
        RECT 28.512 25.704 28.544 25.736 ;
  LAYER M2 ;
        RECT 30.88 25.64 30.912 25.672 ;
  LAYER M2 ;
        RECT 28.512 25.576 28.544 25.608 ;
  LAYER M2 ;
        RECT 30.88 25.512 30.912 25.544 ;
  LAYER M2 ;
        RECT 28.512 25.448 28.544 25.48 ;
  LAYER M2 ;
        RECT 30.88 25.384 30.912 25.416 ;
  LAYER M2 ;
        RECT 28.512 25.32 28.544 25.352 ;
  LAYER M2 ;
        RECT 30.88 25.256 30.912 25.288 ;
  LAYER M2 ;
        RECT 28.512 25.192 28.544 25.224 ;
  LAYER M2 ;
        RECT 30.88 25.128 30.912 25.16 ;
  LAYER M2 ;
        RECT 28.512 25.064 28.544 25.096 ;
  LAYER M2 ;
        RECT 30.88 25 30.912 25.032 ;
  LAYER M2 ;
        RECT 28.512 24.936 28.544 24.968 ;
  LAYER M2 ;
        RECT 30.88 24.872 30.912 24.904 ;
  LAYER M2 ;
        RECT 28.512 24.808 28.544 24.84 ;
  LAYER M2 ;
        RECT 30.88 24.744 30.912 24.776 ;
  LAYER M2 ;
        RECT 28.512 24.68 28.544 24.712 ;
  LAYER M2 ;
        RECT 30.88 24.616 30.912 24.648 ;
  LAYER M2 ;
        RECT 28.512 24.552 28.544 24.584 ;
  LAYER M2 ;
        RECT 30.88 24.488 30.912 24.52 ;
  LAYER M2 ;
        RECT 28.512 24.424 28.544 24.456 ;
  LAYER M2 ;
        RECT 30.88 24.36 30.912 24.392 ;
  LAYER M2 ;
        RECT 28.512 24.296 28.544 24.328 ;
  LAYER M2 ;
        RECT 30.88 24.232 30.912 24.264 ;
  LAYER M2 ;
        RECT 28.512 24.168 28.544 24.2 ;
  LAYER M2 ;
        RECT 30.88 24.104 30.912 24.136 ;
  LAYER M2 ;
        RECT 28.512 24.04 28.544 24.072 ;
  LAYER M2 ;
        RECT 30.88 23.976 30.912 24.008 ;
  LAYER M2 ;
        RECT 28.512 23.912 28.544 23.944 ;
  LAYER M2 ;
        RECT 30.88 23.848 30.912 23.88 ;
  LAYER M2 ;
        RECT 28.512 23.784 28.544 23.816 ;
  LAYER M2 ;
        RECT 30.88 23.72 30.912 23.752 ;
  LAYER M2 ;
        RECT 28.464 23.52 30.96 26.124 ;
  LAYER M1 ;
        RECT 28.512 20.46 28.544 22.968 ;
  LAYER M3 ;
        RECT 28.512 20.48 28.544 20.512 ;
  LAYER M1 ;
        RECT 28.576 20.46 28.608 22.968 ;
  LAYER M3 ;
        RECT 28.576 22.916 28.608 22.948 ;
  LAYER M1 ;
        RECT 28.64 20.46 28.672 22.968 ;
  LAYER M3 ;
        RECT 28.64 20.48 28.672 20.512 ;
  LAYER M1 ;
        RECT 28.704 20.46 28.736 22.968 ;
  LAYER M3 ;
        RECT 28.704 22.916 28.736 22.948 ;
  LAYER M1 ;
        RECT 28.768 20.46 28.8 22.968 ;
  LAYER M3 ;
        RECT 28.768 20.48 28.8 20.512 ;
  LAYER M1 ;
        RECT 28.832 20.46 28.864 22.968 ;
  LAYER M3 ;
        RECT 28.832 22.916 28.864 22.948 ;
  LAYER M1 ;
        RECT 28.896 20.46 28.928 22.968 ;
  LAYER M3 ;
        RECT 28.896 20.48 28.928 20.512 ;
  LAYER M1 ;
        RECT 28.96 20.46 28.992 22.968 ;
  LAYER M3 ;
        RECT 28.96 22.916 28.992 22.948 ;
  LAYER M1 ;
        RECT 29.024 20.46 29.056 22.968 ;
  LAYER M3 ;
        RECT 29.024 20.48 29.056 20.512 ;
  LAYER M1 ;
        RECT 29.088 20.46 29.12 22.968 ;
  LAYER M3 ;
        RECT 29.088 22.916 29.12 22.948 ;
  LAYER M1 ;
        RECT 29.152 20.46 29.184 22.968 ;
  LAYER M3 ;
        RECT 29.152 20.48 29.184 20.512 ;
  LAYER M1 ;
        RECT 29.216 20.46 29.248 22.968 ;
  LAYER M3 ;
        RECT 29.216 22.916 29.248 22.948 ;
  LAYER M1 ;
        RECT 29.28 20.46 29.312 22.968 ;
  LAYER M3 ;
        RECT 29.28 20.48 29.312 20.512 ;
  LAYER M1 ;
        RECT 29.344 20.46 29.376 22.968 ;
  LAYER M3 ;
        RECT 29.344 22.916 29.376 22.948 ;
  LAYER M1 ;
        RECT 29.408 20.46 29.44 22.968 ;
  LAYER M3 ;
        RECT 29.408 20.48 29.44 20.512 ;
  LAYER M1 ;
        RECT 29.472 20.46 29.504 22.968 ;
  LAYER M3 ;
        RECT 29.472 22.916 29.504 22.948 ;
  LAYER M1 ;
        RECT 29.536 20.46 29.568 22.968 ;
  LAYER M3 ;
        RECT 29.536 20.48 29.568 20.512 ;
  LAYER M1 ;
        RECT 29.6 20.46 29.632 22.968 ;
  LAYER M3 ;
        RECT 29.6 22.916 29.632 22.948 ;
  LAYER M1 ;
        RECT 29.664 20.46 29.696 22.968 ;
  LAYER M3 ;
        RECT 29.664 20.48 29.696 20.512 ;
  LAYER M1 ;
        RECT 29.728 20.46 29.76 22.968 ;
  LAYER M3 ;
        RECT 29.728 22.916 29.76 22.948 ;
  LAYER M1 ;
        RECT 29.792 20.46 29.824 22.968 ;
  LAYER M3 ;
        RECT 29.792 20.48 29.824 20.512 ;
  LAYER M1 ;
        RECT 29.856 20.46 29.888 22.968 ;
  LAYER M3 ;
        RECT 29.856 22.916 29.888 22.948 ;
  LAYER M1 ;
        RECT 29.92 20.46 29.952 22.968 ;
  LAYER M3 ;
        RECT 29.92 20.48 29.952 20.512 ;
  LAYER M1 ;
        RECT 29.984 20.46 30.016 22.968 ;
  LAYER M3 ;
        RECT 29.984 22.916 30.016 22.948 ;
  LAYER M1 ;
        RECT 30.048 20.46 30.08 22.968 ;
  LAYER M3 ;
        RECT 30.048 20.48 30.08 20.512 ;
  LAYER M1 ;
        RECT 30.112 20.46 30.144 22.968 ;
  LAYER M3 ;
        RECT 30.112 22.916 30.144 22.948 ;
  LAYER M1 ;
        RECT 30.176 20.46 30.208 22.968 ;
  LAYER M3 ;
        RECT 30.176 20.48 30.208 20.512 ;
  LAYER M1 ;
        RECT 30.24 20.46 30.272 22.968 ;
  LAYER M3 ;
        RECT 30.24 22.916 30.272 22.948 ;
  LAYER M1 ;
        RECT 30.304 20.46 30.336 22.968 ;
  LAYER M3 ;
        RECT 30.304 20.48 30.336 20.512 ;
  LAYER M1 ;
        RECT 30.368 20.46 30.4 22.968 ;
  LAYER M3 ;
        RECT 30.368 22.916 30.4 22.948 ;
  LAYER M1 ;
        RECT 30.432 20.46 30.464 22.968 ;
  LAYER M3 ;
        RECT 30.432 20.48 30.464 20.512 ;
  LAYER M1 ;
        RECT 30.496 20.46 30.528 22.968 ;
  LAYER M3 ;
        RECT 30.496 22.916 30.528 22.948 ;
  LAYER M1 ;
        RECT 30.56 20.46 30.592 22.968 ;
  LAYER M3 ;
        RECT 30.56 20.48 30.592 20.512 ;
  LAYER M1 ;
        RECT 30.624 20.46 30.656 22.968 ;
  LAYER M3 ;
        RECT 30.624 22.916 30.656 22.948 ;
  LAYER M1 ;
        RECT 30.688 20.46 30.72 22.968 ;
  LAYER M3 ;
        RECT 30.688 20.48 30.72 20.512 ;
  LAYER M1 ;
        RECT 30.752 20.46 30.784 22.968 ;
  LAYER M3 ;
        RECT 30.752 22.916 30.784 22.948 ;
  LAYER M1 ;
        RECT 30.816 20.46 30.848 22.968 ;
  LAYER M3 ;
        RECT 30.816 20.48 30.848 20.512 ;
  LAYER M1 ;
        RECT 30.88 20.46 30.912 22.968 ;
  LAYER M3 ;
        RECT 28.512 22.852 28.544 22.884 ;
  LAYER M2 ;
        RECT 30.88 22.788 30.912 22.82 ;
  LAYER M2 ;
        RECT 28.512 22.724 28.544 22.756 ;
  LAYER M2 ;
        RECT 30.88 22.66 30.912 22.692 ;
  LAYER M2 ;
        RECT 28.512 22.596 28.544 22.628 ;
  LAYER M2 ;
        RECT 30.88 22.532 30.912 22.564 ;
  LAYER M2 ;
        RECT 28.512 22.468 28.544 22.5 ;
  LAYER M2 ;
        RECT 30.88 22.404 30.912 22.436 ;
  LAYER M2 ;
        RECT 28.512 22.34 28.544 22.372 ;
  LAYER M2 ;
        RECT 30.88 22.276 30.912 22.308 ;
  LAYER M2 ;
        RECT 28.512 22.212 28.544 22.244 ;
  LAYER M2 ;
        RECT 30.88 22.148 30.912 22.18 ;
  LAYER M2 ;
        RECT 28.512 22.084 28.544 22.116 ;
  LAYER M2 ;
        RECT 30.88 22.02 30.912 22.052 ;
  LAYER M2 ;
        RECT 28.512 21.956 28.544 21.988 ;
  LAYER M2 ;
        RECT 30.88 21.892 30.912 21.924 ;
  LAYER M2 ;
        RECT 28.512 21.828 28.544 21.86 ;
  LAYER M2 ;
        RECT 30.88 21.764 30.912 21.796 ;
  LAYER M2 ;
        RECT 28.512 21.7 28.544 21.732 ;
  LAYER M2 ;
        RECT 30.88 21.636 30.912 21.668 ;
  LAYER M2 ;
        RECT 28.512 21.572 28.544 21.604 ;
  LAYER M2 ;
        RECT 30.88 21.508 30.912 21.54 ;
  LAYER M2 ;
        RECT 28.512 21.444 28.544 21.476 ;
  LAYER M2 ;
        RECT 30.88 21.38 30.912 21.412 ;
  LAYER M2 ;
        RECT 28.512 21.316 28.544 21.348 ;
  LAYER M2 ;
        RECT 30.88 21.252 30.912 21.284 ;
  LAYER M2 ;
        RECT 28.512 21.188 28.544 21.22 ;
  LAYER M2 ;
        RECT 30.88 21.124 30.912 21.156 ;
  LAYER M2 ;
        RECT 28.512 21.06 28.544 21.092 ;
  LAYER M2 ;
        RECT 30.88 20.996 30.912 21.028 ;
  LAYER M2 ;
        RECT 28.512 20.932 28.544 20.964 ;
  LAYER M2 ;
        RECT 30.88 20.868 30.912 20.9 ;
  LAYER M2 ;
        RECT 28.512 20.804 28.544 20.836 ;
  LAYER M2 ;
        RECT 30.88 20.74 30.912 20.772 ;
  LAYER M2 ;
        RECT 28.512 20.676 28.544 20.708 ;
  LAYER M2 ;
        RECT 30.88 20.612 30.912 20.644 ;
  LAYER M2 ;
        RECT 28.464 20.412 30.96 23.016 ;
  END 
END switched_capacitor_filter
