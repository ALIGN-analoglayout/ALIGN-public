MACRO switched_capacitor_combination
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_combination 0 0 ;
  SIZE 16 BY 31.416 ;
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.684 0.32 10.756 0.352 ;
      LAYER M2 ;
        RECT 9.964 0.488 10.036 0.52 ;
      LAYER M2 ;
        RECT 8.604 0.488 8.676 0.52 ;
      LAYER M2 ;
        RECT 10.24 0.32 10.72 0.352 ;
      LAYER M3 ;
        RECT 10.22 0.316 10.26 0.356 ;
      LAYER M4 ;
        RECT 10.08 0.316 10.24 0.356 ;
      LAYER M5 ;
        RECT 10.048 0.336 10.112 0.504 ;
      LAYER M4 ;
        RECT 10.08 0.484 10.24 0.524 ;
      LAYER M3 ;
        RECT 10.22 0.484 10.26 0.524 ;
      LAYER M2 ;
        RECT 10 0.488 10.24 0.52 ;
      LAYER M2 ;
        RECT 8.64 0.488 10.08 0.52 ;
    END
  END phi2
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.764 0.152 10.836 0.184 ;
      LAYER M2 ;
        RECT 10.044 0.656 10.116 0.688 ;
      LAYER M2 ;
        RECT 8.684 0.656 8.756 0.688 ;
      LAYER M2 ;
        RECT 10.08 0.152 10.8 0.184 ;
      LAYER M3 ;
        RECT 10.06 0.168 10.1 0.672 ;
      LAYER M2 ;
        RECT 10.064 0.656 10.096 0.688 ;
      LAYER M2 ;
        RECT 8.88 0.656 10.08 0.688 ;
      LAYER M3 ;
        RECT 8.86 0.652 8.9 0.692 ;
      LAYER M4 ;
        RECT 8.72 0.652 8.88 0.692 ;
      LAYER M3 ;
        RECT 8.7 0.652 8.74 0.692 ;
      LAYER M2 ;
        RECT 8.704 0.656 8.736 0.688 ;
    END
  END agnd
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 0.32 0.436 0.352 ;
      LAYER M2 ;
        RECT 9.324 0.572 9.396 0.604 ;
      LAYER M2 ;
        RECT 7.964 0.572 8.036 0.604 ;
      LAYER M2 ;
        RECT 0.4 0.32 7.6 0.352 ;
      LAYER M3 ;
        RECT 7.58 0.336 7.62 0.588 ;
      LAYER M4 ;
        RECT 7.6 0.568 7.76 0.608 ;
      LAYER M3 ;
        RECT 7.74 0.568 7.78 0.608 ;
      LAYER M2 ;
        RECT 7.76 0.572 8 0.604 ;
      LAYER M2 ;
        RECT 7.92 0.572 9.36 0.604 ;
    END
  END phi1
  PIN Vin
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 0.152 0.356 0.184 ;
    END
  END Vin
  PIN Vin_ota
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.404 0.74 9.476 0.772 ;
      LAYER M1 ;
        RECT 3.76 31.128 3.792 31.2 ;
      LAYER M2 ;
        RECT 3.74 31.148 3.812 31.18 ;
      LAYER M1 ;
        RECT 12.688 31.128 12.72 31.2 ;
      LAYER M2 ;
        RECT 12.668 31.148 12.74 31.18 ;
      LAYER M2 ;
        RECT 3.776 31.148 12.704 31.18 ;
      LAYER M2 ;
        RECT 9.44 0.74 9.68 0.772 ;
      LAYER M3 ;
        RECT 9.66 0.756 9.7 30.996 ;
      LAYER M4 ;
        RECT 9.36 30.976 9.68 31.016 ;
      LAYER M5 ;
        RECT 9.328 30.996 9.392 31.164 ;
      LAYER M4 ;
        RECT 9.34 31.144 9.38 31.184 ;
      LAYER M3 ;
        RECT 9.34 31.144 9.38 31.184 ;
      LAYER M2 ;
        RECT 9.344 31.148 9.376 31.18 ;
    END
  END Vin_ota
  PIN Voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.044 0.74 8.116 0.772 ;
      LAYER M1 ;
        RECT 3.92 14.748 3.952 14.82 ;
      LAYER M2 ;
        RECT 3.9 14.768 3.972 14.8 ;
      LAYER M1 ;
        RECT 12.848 14.748 12.88 14.82 ;
      LAYER M2 ;
        RECT 12.828 14.768 12.9 14.8 ;
      LAYER M2 ;
        RECT 3.936 14.768 12.864 14.8 ;
      LAYER M2 ;
        RECT 8.064 0.74 8.096 0.772 ;
      LAYER M3 ;
        RECT 8.06 0.756 8.1 1.512 ;
      LAYER M4 ;
        RECT 8.08 1.492 8.24 1.532 ;
      LAYER M3 ;
        RECT 8.22 1.512 8.26 14.616 ;
      LAYER M4 ;
        RECT 7.92 14.596 8.24 14.636 ;
      LAYER M5 ;
        RECT 7.888 14.616 7.952 14.784 ;
      LAYER M4 ;
        RECT 7.9 14.764 7.94 14.804 ;
      LAYER M3 ;
        RECT 7.9 14.764 7.94 14.804 ;
      LAYER M2 ;
        RECT 7.904 14.768 7.936 14.8 ;
    END
  END Voutn
  OBS 
  LAYER M1 ;
        RECT 9.632 14.16 9.664 14.232 ;
  LAYER M2 ;
        RECT 9.612 14.18 9.684 14.212 ;
  LAYER M1 ;
        RECT 6.656 14.16 6.688 14.232 ;
  LAYER M2 ;
        RECT 6.636 14.18 6.708 14.212 ;
  LAYER M2 ;
        RECT 6.672 14.18 9.648 14.212 ;
  LAYER M2 ;
        RECT 9.244 0.824 9.956 0.856 ;
  LAYER M1 ;
        RECT 6.736 30.96 6.768 31.032 ;
  LAYER M2 ;
        RECT 6.716 30.98 6.788 31.012 ;
  LAYER M1 ;
        RECT 9.712 30.96 9.744 31.032 ;
  LAYER M2 ;
        RECT 9.692 30.98 9.764 31.012 ;
  LAYER M2 ;
        RECT 6.752 30.98 9.728 31.012 ;
  LAYER M2 ;
        RECT 9.504 14.18 9.536 14.212 ;
  LAYER M3 ;
        RECT 9.5 0.84 9.54 14.196 ;
  LAYER M2 ;
        RECT 9.504 0.824 9.536 0.856 ;
  LAYER M2 ;
        RECT 7.184 14.18 7.216 14.212 ;
  LAYER M3 ;
        RECT 7.18 14.196 7.22 17.724 ;
  LAYER M4 ;
        RECT 7.18 17.704 7.22 17.744 ;
  LAYER M5 ;
        RECT 7.168 17.724 7.232 30.996 ;
  LAYER M4 ;
        RECT 7.18 30.976 7.22 31.016 ;
  LAYER M3 ;
        RECT 7.18 30.976 7.22 31.016 ;
  LAYER M2 ;
        RECT 7.184 30.98 7.216 31.012 ;
  LAYER M1 ;
        RECT 9.792 1.224 9.824 1.296 ;
  LAYER M2 ;
        RECT 9.772 1.244 9.844 1.276 ;
  LAYER M1 ;
        RECT 6.816 1.224 6.848 1.296 ;
  LAYER M2 ;
        RECT 6.796 1.244 6.868 1.276 ;
  LAYER M2 ;
        RECT 6.832 1.244 9.808 1.276 ;
  LAYER M2 ;
        RECT 10.604 0.236 10.676 0.268 ;
  LAYER M2 ;
        RECT 0.444 0.236 0.516 0.268 ;
  LAYER M2 ;
        RECT 9.84 1.244 10.32 1.276 ;
  LAYER M3 ;
        RECT 10.3 0.252 10.34 1.26 ;
  LAYER M4 ;
        RECT 10.32 0.232 10.64 0.272 ;
  LAYER M3 ;
        RECT 10.62 0.232 10.66 0.272 ;
  LAYER M2 ;
        RECT 10.624 0.236 10.656 0.268 ;
  LAYER M2 ;
        RECT 0.8 1.244 6.8 1.276 ;
  LAYER M3 ;
        RECT 0.78 0.252 0.82 1.26 ;
  LAYER M4 ;
        RECT 0.48 0.232 0.8 0.272 ;
  LAYER M3 ;
        RECT 0.46 0.232 0.5 0.272 ;
  LAYER M2 ;
        RECT 0.464 0.236 0.496 0.268 ;
  LAYER M2 ;
        RECT 7.884 0.824 8.596 0.856 ;
  LAYER M1 ;
        RECT 6.896 14.916 6.928 14.988 ;
  LAYER M2 ;
        RECT 6.876 14.936 6.948 14.968 ;
  LAYER M1 ;
        RECT 9.872 14.916 9.904 14.988 ;
  LAYER M2 ;
        RECT 9.852 14.936 9.924 14.968 ;
  LAYER M2 ;
        RECT 6.912 14.936 9.888 14.968 ;
  LAYER M2 ;
        RECT 8.544 0.824 8.576 0.856 ;
  LAYER M3 ;
        RECT 8.54 0.84 8.58 14.952 ;
  LAYER M2 ;
        RECT 8.544 14.936 8.576 14.968 ;
  LAYER M1 ;
        RECT 7.04 4.92 7.072 4.992 ;
  LAYER M2 ;
        RECT 7.02 4.94 7.092 4.972 ;
  LAYER M2 ;
        RECT 7.056 4.94 9.808 4.972 ;
  LAYER M1 ;
        RECT 9.792 4.92 9.824 4.992 ;
  LAYER M2 ;
        RECT 9.772 4.94 9.844 4.972 ;
  LAYER M1 ;
        RECT 7.04 8.028 7.072 8.1 ;
  LAYER M2 ;
        RECT 7.02 8.048 7.092 8.08 ;
  LAYER M2 ;
        RECT 7.056 8.048 9.808 8.08 ;
  LAYER M1 ;
        RECT 9.792 8.028 9.824 8.1 ;
  LAYER M2 ;
        RECT 9.772 8.048 9.844 8.08 ;
  LAYER M1 ;
        RECT 10.016 4.92 10.048 4.992 ;
  LAYER M2 ;
        RECT 9.996 4.94 10.068 4.972 ;
  LAYER M1 ;
        RECT 10.016 4.788 10.048 4.956 ;
  LAYER M1 ;
        RECT 10.016 4.752 10.048 4.824 ;
  LAYER M2 ;
        RECT 9.996 4.772 10.068 4.804 ;
  LAYER M2 ;
        RECT 9.808 4.772 10.032 4.804 ;
  LAYER M1 ;
        RECT 9.792 4.752 9.824 4.824 ;
  LAYER M2 ;
        RECT 9.772 4.772 9.844 4.804 ;
  LAYER M1 ;
        RECT 10.016 8.028 10.048 8.1 ;
  LAYER M2 ;
        RECT 9.996 8.048 10.068 8.08 ;
  LAYER M1 ;
        RECT 10.016 7.896 10.048 8.064 ;
  LAYER M1 ;
        RECT 10.016 7.86 10.048 7.932 ;
  LAYER M2 ;
        RECT 9.996 7.88 10.068 7.912 ;
  LAYER M2 ;
        RECT 9.808 7.88 10.032 7.912 ;
  LAYER M1 ;
        RECT 9.792 7.86 9.824 7.932 ;
  LAYER M2 ;
        RECT 9.772 7.88 9.844 7.912 ;
  LAYER M1 ;
        RECT 9.792 1.224 9.824 1.296 ;
  LAYER M2 ;
        RECT 9.772 1.244 9.844 1.276 ;
  LAYER M1 ;
        RECT 9.792 1.26 9.824 1.512 ;
  LAYER M1 ;
        RECT 9.792 1.512 9.824 8.064 ;
  LAYER M1 ;
        RECT 4.064 8.028 4.096 8.1 ;
  LAYER M2 ;
        RECT 4.044 8.048 4.116 8.08 ;
  LAYER M2 ;
        RECT 4.08 8.048 6.832 8.08 ;
  LAYER M1 ;
        RECT 6.816 8.028 6.848 8.1 ;
  LAYER M2 ;
        RECT 6.796 8.048 6.868 8.08 ;
  LAYER M1 ;
        RECT 4.064 4.92 4.096 4.992 ;
  LAYER M2 ;
        RECT 4.044 4.94 4.116 4.972 ;
  LAYER M2 ;
        RECT 4.08 4.94 6.832 4.972 ;
  LAYER M1 ;
        RECT 6.816 4.92 6.848 4.992 ;
  LAYER M2 ;
        RECT 6.796 4.94 6.868 4.972 ;
  LAYER M1 ;
        RECT 6.816 1.224 6.848 1.296 ;
  LAYER M2 ;
        RECT 6.796 1.244 6.868 1.276 ;
  LAYER M1 ;
        RECT 6.816 1.26 6.848 1.512 ;
  LAYER M1 ;
        RECT 6.816 1.512 6.848 8.064 ;
  LAYER M2 ;
        RECT 6.832 1.244 9.808 1.276 ;
  LAYER M1 ;
        RECT 12.992 1.812 13.024 1.884 ;
  LAYER M2 ;
        RECT 12.972 1.832 13.044 1.864 ;
  LAYER M1 ;
        RECT 12.992 1.68 13.024 1.848 ;
  LAYER M1 ;
        RECT 12.992 1.644 13.024 1.716 ;
  LAYER M2 ;
        RECT 12.972 1.664 13.044 1.696 ;
  LAYER M2 ;
        RECT 12.784 1.664 13.008 1.696 ;
  LAYER M1 ;
        RECT 12.768 1.644 12.8 1.716 ;
  LAYER M2 ;
        RECT 12.748 1.664 12.82 1.696 ;
  LAYER M1 ;
        RECT 12.992 4.92 13.024 4.992 ;
  LAYER M2 ;
        RECT 12.972 4.94 13.044 4.972 ;
  LAYER M1 ;
        RECT 12.992 4.788 13.024 4.956 ;
  LAYER M1 ;
        RECT 12.992 4.752 13.024 4.824 ;
  LAYER M2 ;
        RECT 12.972 4.772 13.044 4.804 ;
  LAYER M2 ;
        RECT 12.784 4.772 13.008 4.804 ;
  LAYER M1 ;
        RECT 12.768 4.752 12.8 4.824 ;
  LAYER M2 ;
        RECT 12.748 4.772 12.82 4.804 ;
  LAYER M1 ;
        RECT 12.992 8.028 13.024 8.1 ;
  LAYER M2 ;
        RECT 12.972 8.048 13.044 8.08 ;
  LAYER M1 ;
        RECT 12.992 7.896 13.024 8.064 ;
  LAYER M1 ;
        RECT 12.992 7.86 13.024 7.932 ;
  LAYER M2 ;
        RECT 12.972 7.88 13.044 7.912 ;
  LAYER M2 ;
        RECT 12.784 7.88 13.008 7.912 ;
  LAYER M1 ;
        RECT 12.768 7.86 12.8 7.932 ;
  LAYER M2 ;
        RECT 12.748 7.88 12.82 7.912 ;
  LAYER M1 ;
        RECT 12.992 11.136 13.024 11.208 ;
  LAYER M2 ;
        RECT 12.972 11.156 13.044 11.188 ;
  LAYER M1 ;
        RECT 12.992 11.004 13.024 11.172 ;
  LAYER M1 ;
        RECT 12.992 10.968 13.024 11.04 ;
  LAYER M2 ;
        RECT 12.972 10.988 13.044 11.02 ;
  LAYER M2 ;
        RECT 12.784 10.988 13.008 11.02 ;
  LAYER M1 ;
        RECT 12.768 10.968 12.8 11.04 ;
  LAYER M2 ;
        RECT 12.748 10.988 12.82 11.02 ;
  LAYER M1 ;
        RECT 10.016 1.812 10.048 1.884 ;
  LAYER M2 ;
        RECT 9.996 1.832 10.068 1.864 ;
  LAYER M2 ;
        RECT 10.032 1.832 12.784 1.864 ;
  LAYER M1 ;
        RECT 12.768 1.812 12.8 1.884 ;
  LAYER M2 ;
        RECT 12.748 1.832 12.82 1.864 ;
  LAYER M1 ;
        RECT 10.016 11.136 10.048 11.208 ;
  LAYER M2 ;
        RECT 9.996 11.156 10.068 11.188 ;
  LAYER M2 ;
        RECT 10.032 11.156 12.784 11.188 ;
  LAYER M1 ;
        RECT 12.768 11.136 12.8 11.208 ;
  LAYER M2 ;
        RECT 12.748 11.156 12.82 11.188 ;
  LAYER M1 ;
        RECT 12.768 1.056 12.8 1.128 ;
  LAYER M2 ;
        RECT 12.748 1.076 12.82 1.108 ;
  LAYER M1 ;
        RECT 12.768 1.092 12.8 1.512 ;
  LAYER M1 ;
        RECT 12.768 1.512 12.8 11.172 ;
  LAYER M1 ;
        RECT 4.064 1.812 4.096 1.884 ;
  LAYER M2 ;
        RECT 4.044 1.832 4.116 1.864 ;
  LAYER M1 ;
        RECT 4.064 1.68 4.096 1.848 ;
  LAYER M1 ;
        RECT 4.064 1.644 4.096 1.716 ;
  LAYER M2 ;
        RECT 4.044 1.664 4.116 1.696 ;
  LAYER M2 ;
        RECT 3.856 1.664 4.08 1.696 ;
  LAYER M1 ;
        RECT 3.84 1.644 3.872 1.716 ;
  LAYER M2 ;
        RECT 3.82 1.664 3.892 1.696 ;
  LAYER M1 ;
        RECT 4.064 11.136 4.096 11.208 ;
  LAYER M2 ;
        RECT 4.044 11.156 4.116 11.188 ;
  LAYER M1 ;
        RECT 4.064 11.004 4.096 11.172 ;
  LAYER M1 ;
        RECT 4.064 10.968 4.096 11.04 ;
  LAYER M2 ;
        RECT 4.044 10.988 4.116 11.02 ;
  LAYER M2 ;
        RECT 3.856 10.988 4.08 11.02 ;
  LAYER M1 ;
        RECT 3.84 10.968 3.872 11.04 ;
  LAYER M2 ;
        RECT 3.82 10.988 3.892 11.02 ;
  LAYER M1 ;
        RECT 1.088 1.812 1.12 1.884 ;
  LAYER M2 ;
        RECT 1.068 1.832 1.14 1.864 ;
  LAYER M2 ;
        RECT 1.104 1.832 3.856 1.864 ;
  LAYER M1 ;
        RECT 3.84 1.812 3.872 1.884 ;
  LAYER M2 ;
        RECT 3.82 1.832 3.892 1.864 ;
  LAYER M1 ;
        RECT 1.088 4.92 1.12 4.992 ;
  LAYER M2 ;
        RECT 1.068 4.94 1.14 4.972 ;
  LAYER M2 ;
        RECT 1.104 4.94 3.856 4.972 ;
  LAYER M1 ;
        RECT 3.84 4.92 3.872 4.992 ;
  LAYER M2 ;
        RECT 3.82 4.94 3.892 4.972 ;
  LAYER M1 ;
        RECT 1.088 8.028 1.12 8.1 ;
  LAYER M2 ;
        RECT 1.068 8.048 1.14 8.08 ;
  LAYER M2 ;
        RECT 1.104 8.048 3.856 8.08 ;
  LAYER M1 ;
        RECT 3.84 8.028 3.872 8.1 ;
  LAYER M2 ;
        RECT 3.82 8.048 3.892 8.08 ;
  LAYER M1 ;
        RECT 1.088 11.136 1.12 11.208 ;
  LAYER M2 ;
        RECT 1.068 11.156 1.14 11.188 ;
  LAYER M2 ;
        RECT 1.104 11.156 3.856 11.188 ;
  LAYER M1 ;
        RECT 3.84 11.136 3.872 11.208 ;
  LAYER M2 ;
        RECT 3.82 11.156 3.892 11.188 ;
  LAYER M1 ;
        RECT 3.84 1.056 3.872 1.128 ;
  LAYER M2 ;
        RECT 3.82 1.076 3.892 1.108 ;
  LAYER M1 ;
        RECT 3.84 1.092 3.872 1.512 ;
  LAYER M1 ;
        RECT 3.84 1.512 3.872 11.172 ;
  LAYER M2 ;
        RECT 3.856 1.076 12.784 1.108 ;
  LAYER M1 ;
        RECT 7.04 11.136 7.072 11.208 ;
  LAYER M2 ;
        RECT 7.02 11.156 7.092 11.188 ;
  LAYER M2 ;
        RECT 7.056 11.156 10.032 11.188 ;
  LAYER M1 ;
        RECT 10.016 11.136 10.048 11.208 ;
  LAYER M2 ;
        RECT 9.996 11.156 10.068 11.188 ;
  LAYER M1 ;
        RECT 7.04 1.812 7.072 1.884 ;
  LAYER M2 ;
        RECT 7.02 1.832 7.092 1.864 ;
  LAYER M2 ;
        RECT 4.08 1.832 7.056 1.864 ;
  LAYER M1 ;
        RECT 4.064 1.812 4.096 1.884 ;
  LAYER M2 ;
        RECT 4.044 1.832 4.116 1.864 ;
  LAYER M1 ;
        RECT 9.408 7.356 9.44 7.428 ;
  LAYER M2 ;
        RECT 9.388 7.376 9.46 7.408 ;
  LAYER M2 ;
        RECT 9.424 7.376 9.648 7.408 ;
  LAYER M1 ;
        RECT 9.632 7.356 9.664 7.428 ;
  LAYER M2 ;
        RECT 9.612 7.376 9.684 7.408 ;
  LAYER M1 ;
        RECT 9.408 10.464 9.44 10.536 ;
  LAYER M2 ;
        RECT 9.388 10.484 9.46 10.516 ;
  LAYER M2 ;
        RECT 9.424 10.484 9.648 10.516 ;
  LAYER M1 ;
        RECT 9.632 10.464 9.664 10.536 ;
  LAYER M2 ;
        RECT 9.612 10.484 9.684 10.516 ;
  LAYER M1 ;
        RECT 12.384 7.356 12.416 7.428 ;
  LAYER M2 ;
        RECT 12.364 7.376 12.436 7.408 ;
  LAYER M1 ;
        RECT 12.384 7.392 12.416 7.56 ;
  LAYER M1 ;
        RECT 12.384 7.524 12.416 7.596 ;
  LAYER M2 ;
        RECT 12.364 7.544 12.436 7.576 ;
  LAYER M2 ;
        RECT 9.648 7.544 12.4 7.576 ;
  LAYER M1 ;
        RECT 9.632 7.524 9.664 7.596 ;
  LAYER M2 ;
        RECT 9.612 7.544 9.684 7.576 ;
  LAYER M1 ;
        RECT 12.384 10.464 12.416 10.536 ;
  LAYER M2 ;
        RECT 12.364 10.484 12.436 10.516 ;
  LAYER M1 ;
        RECT 12.384 10.5 12.416 10.668 ;
  LAYER M1 ;
        RECT 12.384 10.632 12.416 10.704 ;
  LAYER M2 ;
        RECT 12.364 10.652 12.436 10.684 ;
  LAYER M2 ;
        RECT 9.648 10.652 12.4 10.684 ;
  LAYER M1 ;
        RECT 9.632 10.632 9.664 10.704 ;
  LAYER M2 ;
        RECT 9.612 10.652 9.684 10.684 ;
  LAYER M1 ;
        RECT 9.632 14.16 9.664 14.232 ;
  LAYER M2 ;
        RECT 9.612 14.18 9.684 14.212 ;
  LAYER M1 ;
        RECT 9.632 13.944 9.664 14.196 ;
  LAYER M1 ;
        RECT 9.632 7.392 9.664 13.944 ;
  LAYER M1 ;
        RECT 6.432 10.464 6.464 10.536 ;
  LAYER M2 ;
        RECT 6.412 10.484 6.484 10.516 ;
  LAYER M2 ;
        RECT 6.448 10.484 6.672 10.516 ;
  LAYER M1 ;
        RECT 6.656 10.464 6.688 10.536 ;
  LAYER M2 ;
        RECT 6.636 10.484 6.708 10.516 ;
  LAYER M1 ;
        RECT 6.432 7.356 6.464 7.428 ;
  LAYER M2 ;
        RECT 6.412 7.376 6.484 7.408 ;
  LAYER M2 ;
        RECT 6.448 7.376 6.672 7.408 ;
  LAYER M1 ;
        RECT 6.656 7.356 6.688 7.428 ;
  LAYER M2 ;
        RECT 6.636 7.376 6.708 7.408 ;
  LAYER M1 ;
        RECT 6.656 14.16 6.688 14.232 ;
  LAYER M2 ;
        RECT 6.636 14.18 6.708 14.212 ;
  LAYER M1 ;
        RECT 6.656 13.944 6.688 14.196 ;
  LAYER M1 ;
        RECT 6.656 7.392 6.688 13.944 ;
  LAYER M2 ;
        RECT 6.672 14.18 9.648 14.212 ;
  LAYER M1 ;
        RECT 15.36 4.248 15.392 4.32 ;
  LAYER M2 ;
        RECT 15.34 4.268 15.412 4.3 ;
  LAYER M2 ;
        RECT 15.376 4.268 15.76 4.3 ;
  LAYER M1 ;
        RECT 15.744 4.248 15.776 4.32 ;
  LAYER M2 ;
        RECT 15.724 4.268 15.796 4.3 ;
  LAYER M1 ;
        RECT 15.36 7.356 15.392 7.428 ;
  LAYER M2 ;
        RECT 15.34 7.376 15.412 7.408 ;
  LAYER M2 ;
        RECT 15.376 7.376 15.76 7.408 ;
  LAYER M1 ;
        RECT 15.744 7.356 15.776 7.428 ;
  LAYER M2 ;
        RECT 15.724 7.376 15.796 7.408 ;
  LAYER M1 ;
        RECT 15.36 10.464 15.392 10.536 ;
  LAYER M2 ;
        RECT 15.34 10.484 15.412 10.516 ;
  LAYER M2 ;
        RECT 15.376 10.484 15.76 10.516 ;
  LAYER M1 ;
        RECT 15.744 10.464 15.776 10.536 ;
  LAYER M2 ;
        RECT 15.724 10.484 15.796 10.516 ;
  LAYER M1 ;
        RECT 15.36 13.572 15.392 13.644 ;
  LAYER M2 ;
        RECT 15.34 13.592 15.412 13.624 ;
  LAYER M2 ;
        RECT 15.376 13.592 15.76 13.624 ;
  LAYER M1 ;
        RECT 15.744 13.572 15.776 13.644 ;
  LAYER M2 ;
        RECT 15.724 13.592 15.796 13.624 ;
  LAYER M1 ;
        RECT 15.744 14.328 15.776 14.4 ;
  LAYER M2 ;
        RECT 15.724 14.348 15.796 14.38 ;
  LAYER M1 ;
        RECT 15.744 13.944 15.776 14.364 ;
  LAYER M1 ;
        RECT 15.744 4.284 15.776 13.944 ;
  LAYER M1 ;
        RECT 3.456 4.248 3.488 4.32 ;
  LAYER M2 ;
        RECT 3.436 4.268 3.508 4.3 ;
  LAYER M1 ;
        RECT 3.456 4.284 3.488 4.452 ;
  LAYER M1 ;
        RECT 3.456 4.416 3.488 4.488 ;
  LAYER M2 ;
        RECT 3.436 4.436 3.508 4.468 ;
  LAYER M2 ;
        RECT 0.88 4.436 3.472 4.468 ;
  LAYER M1 ;
        RECT 0.864 4.416 0.896 4.488 ;
  LAYER M2 ;
        RECT 0.844 4.436 0.916 4.468 ;
  LAYER M1 ;
        RECT 3.456 7.356 3.488 7.428 ;
  LAYER M2 ;
        RECT 3.436 7.376 3.508 7.408 ;
  LAYER M1 ;
        RECT 3.456 7.392 3.488 7.56 ;
  LAYER M1 ;
        RECT 3.456 7.524 3.488 7.596 ;
  LAYER M2 ;
        RECT 3.436 7.544 3.508 7.576 ;
  LAYER M2 ;
        RECT 0.88 7.544 3.472 7.576 ;
  LAYER M1 ;
        RECT 0.864 7.524 0.896 7.596 ;
  LAYER M2 ;
        RECT 0.844 7.544 0.916 7.576 ;
  LAYER M1 ;
        RECT 3.456 10.464 3.488 10.536 ;
  LAYER M2 ;
        RECT 3.436 10.484 3.508 10.516 ;
  LAYER M1 ;
        RECT 3.456 10.5 3.488 10.668 ;
  LAYER M1 ;
        RECT 3.456 10.632 3.488 10.704 ;
  LAYER M2 ;
        RECT 3.436 10.652 3.508 10.684 ;
  LAYER M2 ;
        RECT 0.88 10.652 3.472 10.684 ;
  LAYER M1 ;
        RECT 0.864 10.632 0.896 10.704 ;
  LAYER M2 ;
        RECT 0.844 10.652 0.916 10.684 ;
  LAYER M1 ;
        RECT 3.456 13.572 3.488 13.644 ;
  LAYER M2 ;
        RECT 3.436 13.592 3.508 13.624 ;
  LAYER M1 ;
        RECT 3.456 13.608 3.488 13.776 ;
  LAYER M1 ;
        RECT 3.456 13.74 3.488 13.812 ;
  LAYER M2 ;
        RECT 3.436 13.76 3.508 13.792 ;
  LAYER M2 ;
        RECT 0.88 13.76 3.472 13.792 ;
  LAYER M1 ;
        RECT 0.864 13.74 0.896 13.812 ;
  LAYER M2 ;
        RECT 0.844 13.76 0.916 13.792 ;
  LAYER M1 ;
        RECT 0.864 14.328 0.896 14.4 ;
  LAYER M2 ;
        RECT 0.844 14.348 0.916 14.38 ;
  LAYER M1 ;
        RECT 0.864 13.944 0.896 14.364 ;
  LAYER M1 ;
        RECT 0.864 4.452 0.896 13.944 ;
  LAYER M2 ;
        RECT 0.88 14.348 15.76 14.38 ;
  LAYER M1 ;
        RECT 12.384 4.248 12.416 4.32 ;
  LAYER M2 ;
        RECT 12.364 4.268 12.436 4.3 ;
  LAYER M2 ;
        RECT 12.4 4.268 15.376 4.3 ;
  LAYER M1 ;
        RECT 15.36 4.248 15.392 4.32 ;
  LAYER M2 ;
        RECT 15.34 4.268 15.412 4.3 ;
  LAYER M1 ;
        RECT 12.384 13.572 12.416 13.644 ;
  LAYER M2 ;
        RECT 12.364 13.592 12.436 13.624 ;
  LAYER M2 ;
        RECT 12.4 13.592 15.376 13.624 ;
  LAYER M1 ;
        RECT 15.36 13.572 15.392 13.644 ;
  LAYER M2 ;
        RECT 15.34 13.592 15.412 13.624 ;
  LAYER M1 ;
        RECT 9.408 13.572 9.44 13.644 ;
  LAYER M2 ;
        RECT 9.388 13.592 9.46 13.624 ;
  LAYER M2 ;
        RECT 9.424 13.592 12.4 13.624 ;
  LAYER M1 ;
        RECT 12.384 13.572 12.416 13.644 ;
  LAYER M2 ;
        RECT 12.364 13.592 12.436 13.624 ;
  LAYER M1 ;
        RECT 6.432 13.572 6.464 13.644 ;
  LAYER M2 ;
        RECT 6.412 13.592 6.484 13.624 ;
  LAYER M2 ;
        RECT 6.448 13.592 9.424 13.624 ;
  LAYER M1 ;
        RECT 9.408 13.572 9.44 13.644 ;
  LAYER M2 ;
        RECT 9.388 13.592 9.46 13.624 ;
  LAYER M1 ;
        RECT 6.432 4.248 6.464 4.32 ;
  LAYER M2 ;
        RECT 6.412 4.268 6.484 4.3 ;
  LAYER M2 ;
        RECT 3.472 4.268 6.448 4.3 ;
  LAYER M1 ;
        RECT 3.456 4.248 3.488 4.32 ;
  LAYER M2 ;
        RECT 3.436 4.268 3.508 4.3 ;
  LAYER M1 ;
        RECT 9.408 4.248 9.44 4.32 ;
  LAYER M2 ;
        RECT 9.388 4.268 9.46 4.3 ;
  LAYER M2 ;
        RECT 6.448 4.268 9.424 4.3 ;
  LAYER M1 ;
        RECT 6.432 4.248 6.464 4.32 ;
  LAYER M2 ;
        RECT 6.412 4.268 6.484 4.3 ;
  LAYER M1 ;
        RECT 15.36 1.812 15.392 4.32 ;
  LAYER M3 ;
        RECT 15.36 4.268 15.392 4.3 ;
  LAYER M1 ;
        RECT 15.296 1.812 15.328 4.32 ;
  LAYER M3 ;
        RECT 15.296 1.832 15.328 1.864 ;
  LAYER M1 ;
        RECT 15.232 1.812 15.264 4.32 ;
  LAYER M3 ;
        RECT 15.232 4.268 15.264 4.3 ;
  LAYER M1 ;
        RECT 15.168 1.812 15.2 4.32 ;
  LAYER M3 ;
        RECT 15.168 1.832 15.2 1.864 ;
  LAYER M1 ;
        RECT 15.104 1.812 15.136 4.32 ;
  LAYER M3 ;
        RECT 15.104 4.268 15.136 4.3 ;
  LAYER M1 ;
        RECT 15.04 1.812 15.072 4.32 ;
  LAYER M3 ;
        RECT 15.04 1.832 15.072 1.864 ;
  LAYER M1 ;
        RECT 14.976 1.812 15.008 4.32 ;
  LAYER M3 ;
        RECT 14.976 4.268 15.008 4.3 ;
  LAYER M1 ;
        RECT 14.912 1.812 14.944 4.32 ;
  LAYER M3 ;
        RECT 14.912 1.832 14.944 1.864 ;
  LAYER M1 ;
        RECT 14.848 1.812 14.88 4.32 ;
  LAYER M3 ;
        RECT 14.848 4.268 14.88 4.3 ;
  LAYER M1 ;
        RECT 14.784 1.812 14.816 4.32 ;
  LAYER M3 ;
        RECT 14.784 1.832 14.816 1.864 ;
  LAYER M1 ;
        RECT 14.72 1.812 14.752 4.32 ;
  LAYER M3 ;
        RECT 14.72 4.268 14.752 4.3 ;
  LAYER M1 ;
        RECT 14.656 1.812 14.688 4.32 ;
  LAYER M3 ;
        RECT 14.656 1.832 14.688 1.864 ;
  LAYER M1 ;
        RECT 14.592 1.812 14.624 4.32 ;
  LAYER M3 ;
        RECT 14.592 4.268 14.624 4.3 ;
  LAYER M1 ;
        RECT 14.528 1.812 14.56 4.32 ;
  LAYER M3 ;
        RECT 14.528 1.832 14.56 1.864 ;
  LAYER M1 ;
        RECT 14.464 1.812 14.496 4.32 ;
  LAYER M3 ;
        RECT 14.464 4.268 14.496 4.3 ;
  LAYER M1 ;
        RECT 14.4 1.812 14.432 4.32 ;
  LAYER M3 ;
        RECT 14.4 1.832 14.432 1.864 ;
  LAYER M1 ;
        RECT 14.336 1.812 14.368 4.32 ;
  LAYER M3 ;
        RECT 14.336 4.268 14.368 4.3 ;
  LAYER M1 ;
        RECT 14.272 1.812 14.304 4.32 ;
  LAYER M3 ;
        RECT 14.272 1.832 14.304 1.864 ;
  LAYER M1 ;
        RECT 14.208 1.812 14.24 4.32 ;
  LAYER M3 ;
        RECT 14.208 4.268 14.24 4.3 ;
  LAYER M1 ;
        RECT 14.144 1.812 14.176 4.32 ;
  LAYER M3 ;
        RECT 14.144 1.832 14.176 1.864 ;
  LAYER M1 ;
        RECT 14.08 1.812 14.112 4.32 ;
  LAYER M3 ;
        RECT 14.08 4.268 14.112 4.3 ;
  LAYER M1 ;
        RECT 14.016 1.812 14.048 4.32 ;
  LAYER M3 ;
        RECT 14.016 1.832 14.048 1.864 ;
  LAYER M1 ;
        RECT 13.952 1.812 13.984 4.32 ;
  LAYER M3 ;
        RECT 13.952 4.268 13.984 4.3 ;
  LAYER M1 ;
        RECT 13.888 1.812 13.92 4.32 ;
  LAYER M3 ;
        RECT 13.888 1.832 13.92 1.864 ;
  LAYER M1 ;
        RECT 13.824 1.812 13.856 4.32 ;
  LAYER M3 ;
        RECT 13.824 4.268 13.856 4.3 ;
  LAYER M1 ;
        RECT 13.76 1.812 13.792 4.32 ;
  LAYER M3 ;
        RECT 13.76 1.832 13.792 1.864 ;
  LAYER M1 ;
        RECT 13.696 1.812 13.728 4.32 ;
  LAYER M3 ;
        RECT 13.696 4.268 13.728 4.3 ;
  LAYER M1 ;
        RECT 13.632 1.812 13.664 4.32 ;
  LAYER M3 ;
        RECT 13.632 1.832 13.664 1.864 ;
  LAYER M1 ;
        RECT 13.568 1.812 13.6 4.32 ;
  LAYER M3 ;
        RECT 13.568 4.268 13.6 4.3 ;
  LAYER M1 ;
        RECT 13.504 1.812 13.536 4.32 ;
  LAYER M3 ;
        RECT 13.504 1.832 13.536 1.864 ;
  LAYER M1 ;
        RECT 13.44 1.812 13.472 4.32 ;
  LAYER M3 ;
        RECT 13.44 4.268 13.472 4.3 ;
  LAYER M1 ;
        RECT 13.376 1.812 13.408 4.32 ;
  LAYER M3 ;
        RECT 13.376 1.832 13.408 1.864 ;
  LAYER M1 ;
        RECT 13.312 1.812 13.344 4.32 ;
  LAYER M3 ;
        RECT 13.312 4.268 13.344 4.3 ;
  LAYER M1 ;
        RECT 13.248 1.812 13.28 4.32 ;
  LAYER M3 ;
        RECT 13.248 1.832 13.28 1.864 ;
  LAYER M1 ;
        RECT 13.184 1.812 13.216 4.32 ;
  LAYER M3 ;
        RECT 13.184 4.268 13.216 4.3 ;
  LAYER M1 ;
        RECT 13.12 1.812 13.152 4.32 ;
  LAYER M3 ;
        RECT 13.12 1.832 13.152 1.864 ;
  LAYER M1 ;
        RECT 13.056 1.812 13.088 4.32 ;
  LAYER M3 ;
        RECT 13.056 4.268 13.088 4.3 ;
  LAYER M1 ;
        RECT 12.992 1.812 13.024 4.32 ;
  LAYER M3 ;
        RECT 15.36 1.896 15.392 1.928 ;
  LAYER M2 ;
        RECT 12.992 1.96 13.024 1.992 ;
  LAYER M2 ;
        RECT 15.36 2.024 15.392 2.056 ;
  LAYER M2 ;
        RECT 12.992 2.088 13.024 2.12 ;
  LAYER M2 ;
        RECT 15.36 2.152 15.392 2.184 ;
  LAYER M2 ;
        RECT 12.992 2.216 13.024 2.248 ;
  LAYER M2 ;
        RECT 15.36 2.28 15.392 2.312 ;
  LAYER M2 ;
        RECT 12.992 2.344 13.024 2.376 ;
  LAYER M2 ;
        RECT 15.36 2.408 15.392 2.44 ;
  LAYER M2 ;
        RECT 12.992 2.472 13.024 2.504 ;
  LAYER M2 ;
        RECT 15.36 2.536 15.392 2.568 ;
  LAYER M2 ;
        RECT 12.992 2.6 13.024 2.632 ;
  LAYER M2 ;
        RECT 15.36 2.664 15.392 2.696 ;
  LAYER M2 ;
        RECT 12.992 2.728 13.024 2.76 ;
  LAYER M2 ;
        RECT 15.36 2.792 15.392 2.824 ;
  LAYER M2 ;
        RECT 12.992 2.856 13.024 2.888 ;
  LAYER M2 ;
        RECT 15.36 2.92 15.392 2.952 ;
  LAYER M2 ;
        RECT 12.992 2.984 13.024 3.016 ;
  LAYER M2 ;
        RECT 15.36 3.048 15.392 3.08 ;
  LAYER M2 ;
        RECT 12.992 3.112 13.024 3.144 ;
  LAYER M2 ;
        RECT 15.36 3.176 15.392 3.208 ;
  LAYER M2 ;
        RECT 12.992 3.24 13.024 3.272 ;
  LAYER M2 ;
        RECT 15.36 3.304 15.392 3.336 ;
  LAYER M2 ;
        RECT 12.992 3.368 13.024 3.4 ;
  LAYER M2 ;
        RECT 15.36 3.432 15.392 3.464 ;
  LAYER M2 ;
        RECT 12.992 3.496 13.024 3.528 ;
  LAYER M2 ;
        RECT 15.36 3.56 15.392 3.592 ;
  LAYER M2 ;
        RECT 12.992 3.624 13.024 3.656 ;
  LAYER M2 ;
        RECT 15.36 3.688 15.392 3.72 ;
  LAYER M2 ;
        RECT 12.992 3.752 13.024 3.784 ;
  LAYER M2 ;
        RECT 15.36 3.816 15.392 3.848 ;
  LAYER M2 ;
        RECT 12.992 3.88 13.024 3.912 ;
  LAYER M2 ;
        RECT 15.36 3.944 15.392 3.976 ;
  LAYER M2 ;
        RECT 12.992 4.008 13.024 4.04 ;
  LAYER M2 ;
        RECT 15.36 4.072 15.392 4.104 ;
  LAYER M2 ;
        RECT 12.992 4.136 13.024 4.168 ;
  LAYER M2 ;
        RECT 12.944 1.764 15.44 4.368 ;
  LAYER M1 ;
        RECT 15.36 4.92 15.392 7.428 ;
  LAYER M3 ;
        RECT 15.36 7.376 15.392 7.408 ;
  LAYER M1 ;
        RECT 15.296 4.92 15.328 7.428 ;
  LAYER M3 ;
        RECT 15.296 4.94 15.328 4.972 ;
  LAYER M1 ;
        RECT 15.232 4.92 15.264 7.428 ;
  LAYER M3 ;
        RECT 15.232 7.376 15.264 7.408 ;
  LAYER M1 ;
        RECT 15.168 4.92 15.2 7.428 ;
  LAYER M3 ;
        RECT 15.168 4.94 15.2 4.972 ;
  LAYER M1 ;
        RECT 15.104 4.92 15.136 7.428 ;
  LAYER M3 ;
        RECT 15.104 7.376 15.136 7.408 ;
  LAYER M1 ;
        RECT 15.04 4.92 15.072 7.428 ;
  LAYER M3 ;
        RECT 15.04 4.94 15.072 4.972 ;
  LAYER M1 ;
        RECT 14.976 4.92 15.008 7.428 ;
  LAYER M3 ;
        RECT 14.976 7.376 15.008 7.408 ;
  LAYER M1 ;
        RECT 14.912 4.92 14.944 7.428 ;
  LAYER M3 ;
        RECT 14.912 4.94 14.944 4.972 ;
  LAYER M1 ;
        RECT 14.848 4.92 14.88 7.428 ;
  LAYER M3 ;
        RECT 14.848 7.376 14.88 7.408 ;
  LAYER M1 ;
        RECT 14.784 4.92 14.816 7.428 ;
  LAYER M3 ;
        RECT 14.784 4.94 14.816 4.972 ;
  LAYER M1 ;
        RECT 14.72 4.92 14.752 7.428 ;
  LAYER M3 ;
        RECT 14.72 7.376 14.752 7.408 ;
  LAYER M1 ;
        RECT 14.656 4.92 14.688 7.428 ;
  LAYER M3 ;
        RECT 14.656 4.94 14.688 4.972 ;
  LAYER M1 ;
        RECT 14.592 4.92 14.624 7.428 ;
  LAYER M3 ;
        RECT 14.592 7.376 14.624 7.408 ;
  LAYER M1 ;
        RECT 14.528 4.92 14.56 7.428 ;
  LAYER M3 ;
        RECT 14.528 4.94 14.56 4.972 ;
  LAYER M1 ;
        RECT 14.464 4.92 14.496 7.428 ;
  LAYER M3 ;
        RECT 14.464 7.376 14.496 7.408 ;
  LAYER M1 ;
        RECT 14.4 4.92 14.432 7.428 ;
  LAYER M3 ;
        RECT 14.4 4.94 14.432 4.972 ;
  LAYER M1 ;
        RECT 14.336 4.92 14.368 7.428 ;
  LAYER M3 ;
        RECT 14.336 7.376 14.368 7.408 ;
  LAYER M1 ;
        RECT 14.272 4.92 14.304 7.428 ;
  LAYER M3 ;
        RECT 14.272 4.94 14.304 4.972 ;
  LAYER M1 ;
        RECT 14.208 4.92 14.24 7.428 ;
  LAYER M3 ;
        RECT 14.208 7.376 14.24 7.408 ;
  LAYER M1 ;
        RECT 14.144 4.92 14.176 7.428 ;
  LAYER M3 ;
        RECT 14.144 4.94 14.176 4.972 ;
  LAYER M1 ;
        RECT 14.08 4.92 14.112 7.428 ;
  LAYER M3 ;
        RECT 14.08 7.376 14.112 7.408 ;
  LAYER M1 ;
        RECT 14.016 4.92 14.048 7.428 ;
  LAYER M3 ;
        RECT 14.016 4.94 14.048 4.972 ;
  LAYER M1 ;
        RECT 13.952 4.92 13.984 7.428 ;
  LAYER M3 ;
        RECT 13.952 7.376 13.984 7.408 ;
  LAYER M1 ;
        RECT 13.888 4.92 13.92 7.428 ;
  LAYER M3 ;
        RECT 13.888 4.94 13.92 4.972 ;
  LAYER M1 ;
        RECT 13.824 4.92 13.856 7.428 ;
  LAYER M3 ;
        RECT 13.824 7.376 13.856 7.408 ;
  LAYER M1 ;
        RECT 13.76 4.92 13.792 7.428 ;
  LAYER M3 ;
        RECT 13.76 4.94 13.792 4.972 ;
  LAYER M1 ;
        RECT 13.696 4.92 13.728 7.428 ;
  LAYER M3 ;
        RECT 13.696 7.376 13.728 7.408 ;
  LAYER M1 ;
        RECT 13.632 4.92 13.664 7.428 ;
  LAYER M3 ;
        RECT 13.632 4.94 13.664 4.972 ;
  LAYER M1 ;
        RECT 13.568 4.92 13.6 7.428 ;
  LAYER M3 ;
        RECT 13.568 7.376 13.6 7.408 ;
  LAYER M1 ;
        RECT 13.504 4.92 13.536 7.428 ;
  LAYER M3 ;
        RECT 13.504 4.94 13.536 4.972 ;
  LAYER M1 ;
        RECT 13.44 4.92 13.472 7.428 ;
  LAYER M3 ;
        RECT 13.44 7.376 13.472 7.408 ;
  LAYER M1 ;
        RECT 13.376 4.92 13.408 7.428 ;
  LAYER M3 ;
        RECT 13.376 4.94 13.408 4.972 ;
  LAYER M1 ;
        RECT 13.312 4.92 13.344 7.428 ;
  LAYER M3 ;
        RECT 13.312 7.376 13.344 7.408 ;
  LAYER M1 ;
        RECT 13.248 4.92 13.28 7.428 ;
  LAYER M3 ;
        RECT 13.248 4.94 13.28 4.972 ;
  LAYER M1 ;
        RECT 13.184 4.92 13.216 7.428 ;
  LAYER M3 ;
        RECT 13.184 7.376 13.216 7.408 ;
  LAYER M1 ;
        RECT 13.12 4.92 13.152 7.428 ;
  LAYER M3 ;
        RECT 13.12 4.94 13.152 4.972 ;
  LAYER M1 ;
        RECT 13.056 4.92 13.088 7.428 ;
  LAYER M3 ;
        RECT 13.056 7.376 13.088 7.408 ;
  LAYER M1 ;
        RECT 12.992 4.92 13.024 7.428 ;
  LAYER M3 ;
        RECT 15.36 5.004 15.392 5.036 ;
  LAYER M2 ;
        RECT 12.992 5.068 13.024 5.1 ;
  LAYER M2 ;
        RECT 15.36 5.132 15.392 5.164 ;
  LAYER M2 ;
        RECT 12.992 5.196 13.024 5.228 ;
  LAYER M2 ;
        RECT 15.36 5.26 15.392 5.292 ;
  LAYER M2 ;
        RECT 12.992 5.324 13.024 5.356 ;
  LAYER M2 ;
        RECT 15.36 5.388 15.392 5.42 ;
  LAYER M2 ;
        RECT 12.992 5.452 13.024 5.484 ;
  LAYER M2 ;
        RECT 15.36 5.516 15.392 5.548 ;
  LAYER M2 ;
        RECT 12.992 5.58 13.024 5.612 ;
  LAYER M2 ;
        RECT 15.36 5.644 15.392 5.676 ;
  LAYER M2 ;
        RECT 12.992 5.708 13.024 5.74 ;
  LAYER M2 ;
        RECT 15.36 5.772 15.392 5.804 ;
  LAYER M2 ;
        RECT 12.992 5.836 13.024 5.868 ;
  LAYER M2 ;
        RECT 15.36 5.9 15.392 5.932 ;
  LAYER M2 ;
        RECT 12.992 5.964 13.024 5.996 ;
  LAYER M2 ;
        RECT 15.36 6.028 15.392 6.06 ;
  LAYER M2 ;
        RECT 12.992 6.092 13.024 6.124 ;
  LAYER M2 ;
        RECT 15.36 6.156 15.392 6.188 ;
  LAYER M2 ;
        RECT 12.992 6.22 13.024 6.252 ;
  LAYER M2 ;
        RECT 15.36 6.284 15.392 6.316 ;
  LAYER M2 ;
        RECT 12.992 6.348 13.024 6.38 ;
  LAYER M2 ;
        RECT 15.36 6.412 15.392 6.444 ;
  LAYER M2 ;
        RECT 12.992 6.476 13.024 6.508 ;
  LAYER M2 ;
        RECT 15.36 6.54 15.392 6.572 ;
  LAYER M2 ;
        RECT 12.992 6.604 13.024 6.636 ;
  LAYER M2 ;
        RECT 15.36 6.668 15.392 6.7 ;
  LAYER M2 ;
        RECT 12.992 6.732 13.024 6.764 ;
  LAYER M2 ;
        RECT 15.36 6.796 15.392 6.828 ;
  LAYER M2 ;
        RECT 12.992 6.86 13.024 6.892 ;
  LAYER M2 ;
        RECT 15.36 6.924 15.392 6.956 ;
  LAYER M2 ;
        RECT 12.992 6.988 13.024 7.02 ;
  LAYER M2 ;
        RECT 15.36 7.052 15.392 7.084 ;
  LAYER M2 ;
        RECT 12.992 7.116 13.024 7.148 ;
  LAYER M2 ;
        RECT 15.36 7.18 15.392 7.212 ;
  LAYER M2 ;
        RECT 12.992 7.244 13.024 7.276 ;
  LAYER M2 ;
        RECT 12.944 4.872 15.44 7.476 ;
  LAYER M1 ;
        RECT 15.36 8.028 15.392 10.536 ;
  LAYER M3 ;
        RECT 15.36 10.484 15.392 10.516 ;
  LAYER M1 ;
        RECT 15.296 8.028 15.328 10.536 ;
  LAYER M3 ;
        RECT 15.296 8.048 15.328 8.08 ;
  LAYER M1 ;
        RECT 15.232 8.028 15.264 10.536 ;
  LAYER M3 ;
        RECT 15.232 10.484 15.264 10.516 ;
  LAYER M1 ;
        RECT 15.168 8.028 15.2 10.536 ;
  LAYER M3 ;
        RECT 15.168 8.048 15.2 8.08 ;
  LAYER M1 ;
        RECT 15.104 8.028 15.136 10.536 ;
  LAYER M3 ;
        RECT 15.104 10.484 15.136 10.516 ;
  LAYER M1 ;
        RECT 15.04 8.028 15.072 10.536 ;
  LAYER M3 ;
        RECT 15.04 8.048 15.072 8.08 ;
  LAYER M1 ;
        RECT 14.976 8.028 15.008 10.536 ;
  LAYER M3 ;
        RECT 14.976 10.484 15.008 10.516 ;
  LAYER M1 ;
        RECT 14.912 8.028 14.944 10.536 ;
  LAYER M3 ;
        RECT 14.912 8.048 14.944 8.08 ;
  LAYER M1 ;
        RECT 14.848 8.028 14.88 10.536 ;
  LAYER M3 ;
        RECT 14.848 10.484 14.88 10.516 ;
  LAYER M1 ;
        RECT 14.784 8.028 14.816 10.536 ;
  LAYER M3 ;
        RECT 14.784 8.048 14.816 8.08 ;
  LAYER M1 ;
        RECT 14.72 8.028 14.752 10.536 ;
  LAYER M3 ;
        RECT 14.72 10.484 14.752 10.516 ;
  LAYER M1 ;
        RECT 14.656 8.028 14.688 10.536 ;
  LAYER M3 ;
        RECT 14.656 8.048 14.688 8.08 ;
  LAYER M1 ;
        RECT 14.592 8.028 14.624 10.536 ;
  LAYER M3 ;
        RECT 14.592 10.484 14.624 10.516 ;
  LAYER M1 ;
        RECT 14.528 8.028 14.56 10.536 ;
  LAYER M3 ;
        RECT 14.528 8.048 14.56 8.08 ;
  LAYER M1 ;
        RECT 14.464 8.028 14.496 10.536 ;
  LAYER M3 ;
        RECT 14.464 10.484 14.496 10.516 ;
  LAYER M1 ;
        RECT 14.4 8.028 14.432 10.536 ;
  LAYER M3 ;
        RECT 14.4 8.048 14.432 8.08 ;
  LAYER M1 ;
        RECT 14.336 8.028 14.368 10.536 ;
  LAYER M3 ;
        RECT 14.336 10.484 14.368 10.516 ;
  LAYER M1 ;
        RECT 14.272 8.028 14.304 10.536 ;
  LAYER M3 ;
        RECT 14.272 8.048 14.304 8.08 ;
  LAYER M1 ;
        RECT 14.208 8.028 14.24 10.536 ;
  LAYER M3 ;
        RECT 14.208 10.484 14.24 10.516 ;
  LAYER M1 ;
        RECT 14.144 8.028 14.176 10.536 ;
  LAYER M3 ;
        RECT 14.144 8.048 14.176 8.08 ;
  LAYER M1 ;
        RECT 14.08 8.028 14.112 10.536 ;
  LAYER M3 ;
        RECT 14.08 10.484 14.112 10.516 ;
  LAYER M1 ;
        RECT 14.016 8.028 14.048 10.536 ;
  LAYER M3 ;
        RECT 14.016 8.048 14.048 8.08 ;
  LAYER M1 ;
        RECT 13.952 8.028 13.984 10.536 ;
  LAYER M3 ;
        RECT 13.952 10.484 13.984 10.516 ;
  LAYER M1 ;
        RECT 13.888 8.028 13.92 10.536 ;
  LAYER M3 ;
        RECT 13.888 8.048 13.92 8.08 ;
  LAYER M1 ;
        RECT 13.824 8.028 13.856 10.536 ;
  LAYER M3 ;
        RECT 13.824 10.484 13.856 10.516 ;
  LAYER M1 ;
        RECT 13.76 8.028 13.792 10.536 ;
  LAYER M3 ;
        RECT 13.76 8.048 13.792 8.08 ;
  LAYER M1 ;
        RECT 13.696 8.028 13.728 10.536 ;
  LAYER M3 ;
        RECT 13.696 10.484 13.728 10.516 ;
  LAYER M1 ;
        RECT 13.632 8.028 13.664 10.536 ;
  LAYER M3 ;
        RECT 13.632 8.048 13.664 8.08 ;
  LAYER M1 ;
        RECT 13.568 8.028 13.6 10.536 ;
  LAYER M3 ;
        RECT 13.568 10.484 13.6 10.516 ;
  LAYER M1 ;
        RECT 13.504 8.028 13.536 10.536 ;
  LAYER M3 ;
        RECT 13.504 8.048 13.536 8.08 ;
  LAYER M1 ;
        RECT 13.44 8.028 13.472 10.536 ;
  LAYER M3 ;
        RECT 13.44 10.484 13.472 10.516 ;
  LAYER M1 ;
        RECT 13.376 8.028 13.408 10.536 ;
  LAYER M3 ;
        RECT 13.376 8.048 13.408 8.08 ;
  LAYER M1 ;
        RECT 13.312 8.028 13.344 10.536 ;
  LAYER M3 ;
        RECT 13.312 10.484 13.344 10.516 ;
  LAYER M1 ;
        RECT 13.248 8.028 13.28 10.536 ;
  LAYER M3 ;
        RECT 13.248 8.048 13.28 8.08 ;
  LAYER M1 ;
        RECT 13.184 8.028 13.216 10.536 ;
  LAYER M3 ;
        RECT 13.184 10.484 13.216 10.516 ;
  LAYER M1 ;
        RECT 13.12 8.028 13.152 10.536 ;
  LAYER M3 ;
        RECT 13.12 8.048 13.152 8.08 ;
  LAYER M1 ;
        RECT 13.056 8.028 13.088 10.536 ;
  LAYER M3 ;
        RECT 13.056 10.484 13.088 10.516 ;
  LAYER M1 ;
        RECT 12.992 8.028 13.024 10.536 ;
  LAYER M3 ;
        RECT 15.36 8.112 15.392 8.144 ;
  LAYER M2 ;
        RECT 12.992 8.176 13.024 8.208 ;
  LAYER M2 ;
        RECT 15.36 8.24 15.392 8.272 ;
  LAYER M2 ;
        RECT 12.992 8.304 13.024 8.336 ;
  LAYER M2 ;
        RECT 15.36 8.368 15.392 8.4 ;
  LAYER M2 ;
        RECT 12.992 8.432 13.024 8.464 ;
  LAYER M2 ;
        RECT 15.36 8.496 15.392 8.528 ;
  LAYER M2 ;
        RECT 12.992 8.56 13.024 8.592 ;
  LAYER M2 ;
        RECT 15.36 8.624 15.392 8.656 ;
  LAYER M2 ;
        RECT 12.992 8.688 13.024 8.72 ;
  LAYER M2 ;
        RECT 15.36 8.752 15.392 8.784 ;
  LAYER M2 ;
        RECT 12.992 8.816 13.024 8.848 ;
  LAYER M2 ;
        RECT 15.36 8.88 15.392 8.912 ;
  LAYER M2 ;
        RECT 12.992 8.944 13.024 8.976 ;
  LAYER M2 ;
        RECT 15.36 9.008 15.392 9.04 ;
  LAYER M2 ;
        RECT 12.992 9.072 13.024 9.104 ;
  LAYER M2 ;
        RECT 15.36 9.136 15.392 9.168 ;
  LAYER M2 ;
        RECT 12.992 9.2 13.024 9.232 ;
  LAYER M2 ;
        RECT 15.36 9.264 15.392 9.296 ;
  LAYER M2 ;
        RECT 12.992 9.328 13.024 9.36 ;
  LAYER M2 ;
        RECT 15.36 9.392 15.392 9.424 ;
  LAYER M2 ;
        RECT 12.992 9.456 13.024 9.488 ;
  LAYER M2 ;
        RECT 15.36 9.52 15.392 9.552 ;
  LAYER M2 ;
        RECT 12.992 9.584 13.024 9.616 ;
  LAYER M2 ;
        RECT 15.36 9.648 15.392 9.68 ;
  LAYER M2 ;
        RECT 12.992 9.712 13.024 9.744 ;
  LAYER M2 ;
        RECT 15.36 9.776 15.392 9.808 ;
  LAYER M2 ;
        RECT 12.992 9.84 13.024 9.872 ;
  LAYER M2 ;
        RECT 15.36 9.904 15.392 9.936 ;
  LAYER M2 ;
        RECT 12.992 9.968 13.024 10 ;
  LAYER M2 ;
        RECT 15.36 10.032 15.392 10.064 ;
  LAYER M2 ;
        RECT 12.992 10.096 13.024 10.128 ;
  LAYER M2 ;
        RECT 15.36 10.16 15.392 10.192 ;
  LAYER M2 ;
        RECT 12.992 10.224 13.024 10.256 ;
  LAYER M2 ;
        RECT 15.36 10.288 15.392 10.32 ;
  LAYER M2 ;
        RECT 12.992 10.352 13.024 10.384 ;
  LAYER M2 ;
        RECT 12.944 7.98 15.44 10.584 ;
  LAYER M1 ;
        RECT 15.36 11.136 15.392 13.644 ;
  LAYER M3 ;
        RECT 15.36 13.592 15.392 13.624 ;
  LAYER M1 ;
        RECT 15.296 11.136 15.328 13.644 ;
  LAYER M3 ;
        RECT 15.296 11.156 15.328 11.188 ;
  LAYER M1 ;
        RECT 15.232 11.136 15.264 13.644 ;
  LAYER M3 ;
        RECT 15.232 13.592 15.264 13.624 ;
  LAYER M1 ;
        RECT 15.168 11.136 15.2 13.644 ;
  LAYER M3 ;
        RECT 15.168 11.156 15.2 11.188 ;
  LAYER M1 ;
        RECT 15.104 11.136 15.136 13.644 ;
  LAYER M3 ;
        RECT 15.104 13.592 15.136 13.624 ;
  LAYER M1 ;
        RECT 15.04 11.136 15.072 13.644 ;
  LAYER M3 ;
        RECT 15.04 11.156 15.072 11.188 ;
  LAYER M1 ;
        RECT 14.976 11.136 15.008 13.644 ;
  LAYER M3 ;
        RECT 14.976 13.592 15.008 13.624 ;
  LAYER M1 ;
        RECT 14.912 11.136 14.944 13.644 ;
  LAYER M3 ;
        RECT 14.912 11.156 14.944 11.188 ;
  LAYER M1 ;
        RECT 14.848 11.136 14.88 13.644 ;
  LAYER M3 ;
        RECT 14.848 13.592 14.88 13.624 ;
  LAYER M1 ;
        RECT 14.784 11.136 14.816 13.644 ;
  LAYER M3 ;
        RECT 14.784 11.156 14.816 11.188 ;
  LAYER M1 ;
        RECT 14.72 11.136 14.752 13.644 ;
  LAYER M3 ;
        RECT 14.72 13.592 14.752 13.624 ;
  LAYER M1 ;
        RECT 14.656 11.136 14.688 13.644 ;
  LAYER M3 ;
        RECT 14.656 11.156 14.688 11.188 ;
  LAYER M1 ;
        RECT 14.592 11.136 14.624 13.644 ;
  LAYER M3 ;
        RECT 14.592 13.592 14.624 13.624 ;
  LAYER M1 ;
        RECT 14.528 11.136 14.56 13.644 ;
  LAYER M3 ;
        RECT 14.528 11.156 14.56 11.188 ;
  LAYER M1 ;
        RECT 14.464 11.136 14.496 13.644 ;
  LAYER M3 ;
        RECT 14.464 13.592 14.496 13.624 ;
  LAYER M1 ;
        RECT 14.4 11.136 14.432 13.644 ;
  LAYER M3 ;
        RECT 14.4 11.156 14.432 11.188 ;
  LAYER M1 ;
        RECT 14.336 11.136 14.368 13.644 ;
  LAYER M3 ;
        RECT 14.336 13.592 14.368 13.624 ;
  LAYER M1 ;
        RECT 14.272 11.136 14.304 13.644 ;
  LAYER M3 ;
        RECT 14.272 11.156 14.304 11.188 ;
  LAYER M1 ;
        RECT 14.208 11.136 14.24 13.644 ;
  LAYER M3 ;
        RECT 14.208 13.592 14.24 13.624 ;
  LAYER M1 ;
        RECT 14.144 11.136 14.176 13.644 ;
  LAYER M3 ;
        RECT 14.144 11.156 14.176 11.188 ;
  LAYER M1 ;
        RECT 14.08 11.136 14.112 13.644 ;
  LAYER M3 ;
        RECT 14.08 13.592 14.112 13.624 ;
  LAYER M1 ;
        RECT 14.016 11.136 14.048 13.644 ;
  LAYER M3 ;
        RECT 14.016 11.156 14.048 11.188 ;
  LAYER M1 ;
        RECT 13.952 11.136 13.984 13.644 ;
  LAYER M3 ;
        RECT 13.952 13.592 13.984 13.624 ;
  LAYER M1 ;
        RECT 13.888 11.136 13.92 13.644 ;
  LAYER M3 ;
        RECT 13.888 11.156 13.92 11.188 ;
  LAYER M1 ;
        RECT 13.824 11.136 13.856 13.644 ;
  LAYER M3 ;
        RECT 13.824 13.592 13.856 13.624 ;
  LAYER M1 ;
        RECT 13.76 11.136 13.792 13.644 ;
  LAYER M3 ;
        RECT 13.76 11.156 13.792 11.188 ;
  LAYER M1 ;
        RECT 13.696 11.136 13.728 13.644 ;
  LAYER M3 ;
        RECT 13.696 13.592 13.728 13.624 ;
  LAYER M1 ;
        RECT 13.632 11.136 13.664 13.644 ;
  LAYER M3 ;
        RECT 13.632 11.156 13.664 11.188 ;
  LAYER M1 ;
        RECT 13.568 11.136 13.6 13.644 ;
  LAYER M3 ;
        RECT 13.568 13.592 13.6 13.624 ;
  LAYER M1 ;
        RECT 13.504 11.136 13.536 13.644 ;
  LAYER M3 ;
        RECT 13.504 11.156 13.536 11.188 ;
  LAYER M1 ;
        RECT 13.44 11.136 13.472 13.644 ;
  LAYER M3 ;
        RECT 13.44 13.592 13.472 13.624 ;
  LAYER M1 ;
        RECT 13.376 11.136 13.408 13.644 ;
  LAYER M3 ;
        RECT 13.376 11.156 13.408 11.188 ;
  LAYER M1 ;
        RECT 13.312 11.136 13.344 13.644 ;
  LAYER M3 ;
        RECT 13.312 13.592 13.344 13.624 ;
  LAYER M1 ;
        RECT 13.248 11.136 13.28 13.644 ;
  LAYER M3 ;
        RECT 13.248 11.156 13.28 11.188 ;
  LAYER M1 ;
        RECT 13.184 11.136 13.216 13.644 ;
  LAYER M3 ;
        RECT 13.184 13.592 13.216 13.624 ;
  LAYER M1 ;
        RECT 13.12 11.136 13.152 13.644 ;
  LAYER M3 ;
        RECT 13.12 11.156 13.152 11.188 ;
  LAYER M1 ;
        RECT 13.056 11.136 13.088 13.644 ;
  LAYER M3 ;
        RECT 13.056 13.592 13.088 13.624 ;
  LAYER M1 ;
        RECT 12.992 11.136 13.024 13.644 ;
  LAYER M3 ;
        RECT 15.36 11.22 15.392 11.252 ;
  LAYER M2 ;
        RECT 12.992 11.284 13.024 11.316 ;
  LAYER M2 ;
        RECT 15.36 11.348 15.392 11.38 ;
  LAYER M2 ;
        RECT 12.992 11.412 13.024 11.444 ;
  LAYER M2 ;
        RECT 15.36 11.476 15.392 11.508 ;
  LAYER M2 ;
        RECT 12.992 11.54 13.024 11.572 ;
  LAYER M2 ;
        RECT 15.36 11.604 15.392 11.636 ;
  LAYER M2 ;
        RECT 12.992 11.668 13.024 11.7 ;
  LAYER M2 ;
        RECT 15.36 11.732 15.392 11.764 ;
  LAYER M2 ;
        RECT 12.992 11.796 13.024 11.828 ;
  LAYER M2 ;
        RECT 15.36 11.86 15.392 11.892 ;
  LAYER M2 ;
        RECT 12.992 11.924 13.024 11.956 ;
  LAYER M2 ;
        RECT 15.36 11.988 15.392 12.02 ;
  LAYER M2 ;
        RECT 12.992 12.052 13.024 12.084 ;
  LAYER M2 ;
        RECT 15.36 12.116 15.392 12.148 ;
  LAYER M2 ;
        RECT 12.992 12.18 13.024 12.212 ;
  LAYER M2 ;
        RECT 15.36 12.244 15.392 12.276 ;
  LAYER M2 ;
        RECT 12.992 12.308 13.024 12.34 ;
  LAYER M2 ;
        RECT 15.36 12.372 15.392 12.404 ;
  LAYER M2 ;
        RECT 12.992 12.436 13.024 12.468 ;
  LAYER M2 ;
        RECT 15.36 12.5 15.392 12.532 ;
  LAYER M2 ;
        RECT 12.992 12.564 13.024 12.596 ;
  LAYER M2 ;
        RECT 15.36 12.628 15.392 12.66 ;
  LAYER M2 ;
        RECT 12.992 12.692 13.024 12.724 ;
  LAYER M2 ;
        RECT 15.36 12.756 15.392 12.788 ;
  LAYER M2 ;
        RECT 12.992 12.82 13.024 12.852 ;
  LAYER M2 ;
        RECT 15.36 12.884 15.392 12.916 ;
  LAYER M2 ;
        RECT 12.992 12.948 13.024 12.98 ;
  LAYER M2 ;
        RECT 15.36 13.012 15.392 13.044 ;
  LAYER M2 ;
        RECT 12.992 13.076 13.024 13.108 ;
  LAYER M2 ;
        RECT 15.36 13.14 15.392 13.172 ;
  LAYER M2 ;
        RECT 12.992 13.204 13.024 13.236 ;
  LAYER M2 ;
        RECT 15.36 13.268 15.392 13.3 ;
  LAYER M2 ;
        RECT 12.992 13.332 13.024 13.364 ;
  LAYER M2 ;
        RECT 15.36 13.396 15.392 13.428 ;
  LAYER M2 ;
        RECT 12.992 13.46 13.024 13.492 ;
  LAYER M2 ;
        RECT 12.944 11.088 15.44 13.692 ;
  LAYER M1 ;
        RECT 12.384 1.812 12.416 4.32 ;
  LAYER M3 ;
        RECT 12.384 4.268 12.416 4.3 ;
  LAYER M1 ;
        RECT 12.32 1.812 12.352 4.32 ;
  LAYER M3 ;
        RECT 12.32 1.832 12.352 1.864 ;
  LAYER M1 ;
        RECT 12.256 1.812 12.288 4.32 ;
  LAYER M3 ;
        RECT 12.256 4.268 12.288 4.3 ;
  LAYER M1 ;
        RECT 12.192 1.812 12.224 4.32 ;
  LAYER M3 ;
        RECT 12.192 1.832 12.224 1.864 ;
  LAYER M1 ;
        RECT 12.128 1.812 12.16 4.32 ;
  LAYER M3 ;
        RECT 12.128 4.268 12.16 4.3 ;
  LAYER M1 ;
        RECT 12.064 1.812 12.096 4.32 ;
  LAYER M3 ;
        RECT 12.064 1.832 12.096 1.864 ;
  LAYER M1 ;
        RECT 12 1.812 12.032 4.32 ;
  LAYER M3 ;
        RECT 12 4.268 12.032 4.3 ;
  LAYER M1 ;
        RECT 11.936 1.812 11.968 4.32 ;
  LAYER M3 ;
        RECT 11.936 1.832 11.968 1.864 ;
  LAYER M1 ;
        RECT 11.872 1.812 11.904 4.32 ;
  LAYER M3 ;
        RECT 11.872 4.268 11.904 4.3 ;
  LAYER M1 ;
        RECT 11.808 1.812 11.84 4.32 ;
  LAYER M3 ;
        RECT 11.808 1.832 11.84 1.864 ;
  LAYER M1 ;
        RECT 11.744 1.812 11.776 4.32 ;
  LAYER M3 ;
        RECT 11.744 4.268 11.776 4.3 ;
  LAYER M1 ;
        RECT 11.68 1.812 11.712 4.32 ;
  LAYER M3 ;
        RECT 11.68 1.832 11.712 1.864 ;
  LAYER M1 ;
        RECT 11.616 1.812 11.648 4.32 ;
  LAYER M3 ;
        RECT 11.616 4.268 11.648 4.3 ;
  LAYER M1 ;
        RECT 11.552 1.812 11.584 4.32 ;
  LAYER M3 ;
        RECT 11.552 1.832 11.584 1.864 ;
  LAYER M1 ;
        RECT 11.488 1.812 11.52 4.32 ;
  LAYER M3 ;
        RECT 11.488 4.268 11.52 4.3 ;
  LAYER M1 ;
        RECT 11.424 1.812 11.456 4.32 ;
  LAYER M3 ;
        RECT 11.424 1.832 11.456 1.864 ;
  LAYER M1 ;
        RECT 11.36 1.812 11.392 4.32 ;
  LAYER M3 ;
        RECT 11.36 4.268 11.392 4.3 ;
  LAYER M1 ;
        RECT 11.296 1.812 11.328 4.32 ;
  LAYER M3 ;
        RECT 11.296 1.832 11.328 1.864 ;
  LAYER M1 ;
        RECT 11.232 1.812 11.264 4.32 ;
  LAYER M3 ;
        RECT 11.232 4.268 11.264 4.3 ;
  LAYER M1 ;
        RECT 11.168 1.812 11.2 4.32 ;
  LAYER M3 ;
        RECT 11.168 1.832 11.2 1.864 ;
  LAYER M1 ;
        RECT 11.104 1.812 11.136 4.32 ;
  LAYER M3 ;
        RECT 11.104 4.268 11.136 4.3 ;
  LAYER M1 ;
        RECT 11.04 1.812 11.072 4.32 ;
  LAYER M3 ;
        RECT 11.04 1.832 11.072 1.864 ;
  LAYER M1 ;
        RECT 10.976 1.812 11.008 4.32 ;
  LAYER M3 ;
        RECT 10.976 4.268 11.008 4.3 ;
  LAYER M1 ;
        RECT 10.912 1.812 10.944 4.32 ;
  LAYER M3 ;
        RECT 10.912 1.832 10.944 1.864 ;
  LAYER M1 ;
        RECT 10.848 1.812 10.88 4.32 ;
  LAYER M3 ;
        RECT 10.848 4.268 10.88 4.3 ;
  LAYER M1 ;
        RECT 10.784 1.812 10.816 4.32 ;
  LAYER M3 ;
        RECT 10.784 1.832 10.816 1.864 ;
  LAYER M1 ;
        RECT 10.72 1.812 10.752 4.32 ;
  LAYER M3 ;
        RECT 10.72 4.268 10.752 4.3 ;
  LAYER M1 ;
        RECT 10.656 1.812 10.688 4.32 ;
  LAYER M3 ;
        RECT 10.656 1.832 10.688 1.864 ;
  LAYER M1 ;
        RECT 10.592 1.812 10.624 4.32 ;
  LAYER M3 ;
        RECT 10.592 4.268 10.624 4.3 ;
  LAYER M1 ;
        RECT 10.528 1.812 10.56 4.32 ;
  LAYER M3 ;
        RECT 10.528 1.832 10.56 1.864 ;
  LAYER M1 ;
        RECT 10.464 1.812 10.496 4.32 ;
  LAYER M3 ;
        RECT 10.464 4.268 10.496 4.3 ;
  LAYER M1 ;
        RECT 10.4 1.812 10.432 4.32 ;
  LAYER M3 ;
        RECT 10.4 1.832 10.432 1.864 ;
  LAYER M1 ;
        RECT 10.336 1.812 10.368 4.32 ;
  LAYER M3 ;
        RECT 10.336 4.268 10.368 4.3 ;
  LAYER M1 ;
        RECT 10.272 1.812 10.304 4.32 ;
  LAYER M3 ;
        RECT 10.272 1.832 10.304 1.864 ;
  LAYER M1 ;
        RECT 10.208 1.812 10.24 4.32 ;
  LAYER M3 ;
        RECT 10.208 4.268 10.24 4.3 ;
  LAYER M1 ;
        RECT 10.144 1.812 10.176 4.32 ;
  LAYER M3 ;
        RECT 10.144 1.832 10.176 1.864 ;
  LAYER M1 ;
        RECT 10.08 1.812 10.112 4.32 ;
  LAYER M3 ;
        RECT 10.08 4.268 10.112 4.3 ;
  LAYER M1 ;
        RECT 10.016 1.812 10.048 4.32 ;
  LAYER M3 ;
        RECT 12.384 1.896 12.416 1.928 ;
  LAYER M2 ;
        RECT 10.016 1.96 10.048 1.992 ;
  LAYER M2 ;
        RECT 12.384 2.024 12.416 2.056 ;
  LAYER M2 ;
        RECT 10.016 2.088 10.048 2.12 ;
  LAYER M2 ;
        RECT 12.384 2.152 12.416 2.184 ;
  LAYER M2 ;
        RECT 10.016 2.216 10.048 2.248 ;
  LAYER M2 ;
        RECT 12.384 2.28 12.416 2.312 ;
  LAYER M2 ;
        RECT 10.016 2.344 10.048 2.376 ;
  LAYER M2 ;
        RECT 12.384 2.408 12.416 2.44 ;
  LAYER M2 ;
        RECT 10.016 2.472 10.048 2.504 ;
  LAYER M2 ;
        RECT 12.384 2.536 12.416 2.568 ;
  LAYER M2 ;
        RECT 10.016 2.6 10.048 2.632 ;
  LAYER M2 ;
        RECT 12.384 2.664 12.416 2.696 ;
  LAYER M2 ;
        RECT 10.016 2.728 10.048 2.76 ;
  LAYER M2 ;
        RECT 12.384 2.792 12.416 2.824 ;
  LAYER M2 ;
        RECT 10.016 2.856 10.048 2.888 ;
  LAYER M2 ;
        RECT 12.384 2.92 12.416 2.952 ;
  LAYER M2 ;
        RECT 10.016 2.984 10.048 3.016 ;
  LAYER M2 ;
        RECT 12.384 3.048 12.416 3.08 ;
  LAYER M2 ;
        RECT 10.016 3.112 10.048 3.144 ;
  LAYER M2 ;
        RECT 12.384 3.176 12.416 3.208 ;
  LAYER M2 ;
        RECT 10.016 3.24 10.048 3.272 ;
  LAYER M2 ;
        RECT 12.384 3.304 12.416 3.336 ;
  LAYER M2 ;
        RECT 10.016 3.368 10.048 3.4 ;
  LAYER M2 ;
        RECT 12.384 3.432 12.416 3.464 ;
  LAYER M2 ;
        RECT 10.016 3.496 10.048 3.528 ;
  LAYER M2 ;
        RECT 12.384 3.56 12.416 3.592 ;
  LAYER M2 ;
        RECT 10.016 3.624 10.048 3.656 ;
  LAYER M2 ;
        RECT 12.384 3.688 12.416 3.72 ;
  LAYER M2 ;
        RECT 10.016 3.752 10.048 3.784 ;
  LAYER M2 ;
        RECT 12.384 3.816 12.416 3.848 ;
  LAYER M2 ;
        RECT 10.016 3.88 10.048 3.912 ;
  LAYER M2 ;
        RECT 12.384 3.944 12.416 3.976 ;
  LAYER M2 ;
        RECT 10.016 4.008 10.048 4.04 ;
  LAYER M2 ;
        RECT 12.384 4.072 12.416 4.104 ;
  LAYER M2 ;
        RECT 10.016 4.136 10.048 4.168 ;
  LAYER M2 ;
        RECT 9.968 1.764 12.464 4.368 ;
  LAYER M1 ;
        RECT 12.384 4.92 12.416 7.428 ;
  LAYER M3 ;
        RECT 12.384 7.376 12.416 7.408 ;
  LAYER M1 ;
        RECT 12.32 4.92 12.352 7.428 ;
  LAYER M3 ;
        RECT 12.32 4.94 12.352 4.972 ;
  LAYER M1 ;
        RECT 12.256 4.92 12.288 7.428 ;
  LAYER M3 ;
        RECT 12.256 7.376 12.288 7.408 ;
  LAYER M1 ;
        RECT 12.192 4.92 12.224 7.428 ;
  LAYER M3 ;
        RECT 12.192 4.94 12.224 4.972 ;
  LAYER M1 ;
        RECT 12.128 4.92 12.16 7.428 ;
  LAYER M3 ;
        RECT 12.128 7.376 12.16 7.408 ;
  LAYER M1 ;
        RECT 12.064 4.92 12.096 7.428 ;
  LAYER M3 ;
        RECT 12.064 4.94 12.096 4.972 ;
  LAYER M1 ;
        RECT 12 4.92 12.032 7.428 ;
  LAYER M3 ;
        RECT 12 7.376 12.032 7.408 ;
  LAYER M1 ;
        RECT 11.936 4.92 11.968 7.428 ;
  LAYER M3 ;
        RECT 11.936 4.94 11.968 4.972 ;
  LAYER M1 ;
        RECT 11.872 4.92 11.904 7.428 ;
  LAYER M3 ;
        RECT 11.872 7.376 11.904 7.408 ;
  LAYER M1 ;
        RECT 11.808 4.92 11.84 7.428 ;
  LAYER M3 ;
        RECT 11.808 4.94 11.84 4.972 ;
  LAYER M1 ;
        RECT 11.744 4.92 11.776 7.428 ;
  LAYER M3 ;
        RECT 11.744 7.376 11.776 7.408 ;
  LAYER M1 ;
        RECT 11.68 4.92 11.712 7.428 ;
  LAYER M3 ;
        RECT 11.68 4.94 11.712 4.972 ;
  LAYER M1 ;
        RECT 11.616 4.92 11.648 7.428 ;
  LAYER M3 ;
        RECT 11.616 7.376 11.648 7.408 ;
  LAYER M1 ;
        RECT 11.552 4.92 11.584 7.428 ;
  LAYER M3 ;
        RECT 11.552 4.94 11.584 4.972 ;
  LAYER M1 ;
        RECT 11.488 4.92 11.52 7.428 ;
  LAYER M3 ;
        RECT 11.488 7.376 11.52 7.408 ;
  LAYER M1 ;
        RECT 11.424 4.92 11.456 7.428 ;
  LAYER M3 ;
        RECT 11.424 4.94 11.456 4.972 ;
  LAYER M1 ;
        RECT 11.36 4.92 11.392 7.428 ;
  LAYER M3 ;
        RECT 11.36 7.376 11.392 7.408 ;
  LAYER M1 ;
        RECT 11.296 4.92 11.328 7.428 ;
  LAYER M3 ;
        RECT 11.296 4.94 11.328 4.972 ;
  LAYER M1 ;
        RECT 11.232 4.92 11.264 7.428 ;
  LAYER M3 ;
        RECT 11.232 7.376 11.264 7.408 ;
  LAYER M1 ;
        RECT 11.168 4.92 11.2 7.428 ;
  LAYER M3 ;
        RECT 11.168 4.94 11.2 4.972 ;
  LAYER M1 ;
        RECT 11.104 4.92 11.136 7.428 ;
  LAYER M3 ;
        RECT 11.104 7.376 11.136 7.408 ;
  LAYER M1 ;
        RECT 11.04 4.92 11.072 7.428 ;
  LAYER M3 ;
        RECT 11.04 4.94 11.072 4.972 ;
  LAYER M1 ;
        RECT 10.976 4.92 11.008 7.428 ;
  LAYER M3 ;
        RECT 10.976 7.376 11.008 7.408 ;
  LAYER M1 ;
        RECT 10.912 4.92 10.944 7.428 ;
  LAYER M3 ;
        RECT 10.912 4.94 10.944 4.972 ;
  LAYER M1 ;
        RECT 10.848 4.92 10.88 7.428 ;
  LAYER M3 ;
        RECT 10.848 7.376 10.88 7.408 ;
  LAYER M1 ;
        RECT 10.784 4.92 10.816 7.428 ;
  LAYER M3 ;
        RECT 10.784 4.94 10.816 4.972 ;
  LAYER M1 ;
        RECT 10.72 4.92 10.752 7.428 ;
  LAYER M3 ;
        RECT 10.72 7.376 10.752 7.408 ;
  LAYER M1 ;
        RECT 10.656 4.92 10.688 7.428 ;
  LAYER M3 ;
        RECT 10.656 4.94 10.688 4.972 ;
  LAYER M1 ;
        RECT 10.592 4.92 10.624 7.428 ;
  LAYER M3 ;
        RECT 10.592 7.376 10.624 7.408 ;
  LAYER M1 ;
        RECT 10.528 4.92 10.56 7.428 ;
  LAYER M3 ;
        RECT 10.528 4.94 10.56 4.972 ;
  LAYER M1 ;
        RECT 10.464 4.92 10.496 7.428 ;
  LAYER M3 ;
        RECT 10.464 7.376 10.496 7.408 ;
  LAYER M1 ;
        RECT 10.4 4.92 10.432 7.428 ;
  LAYER M3 ;
        RECT 10.4 4.94 10.432 4.972 ;
  LAYER M1 ;
        RECT 10.336 4.92 10.368 7.428 ;
  LAYER M3 ;
        RECT 10.336 7.376 10.368 7.408 ;
  LAYER M1 ;
        RECT 10.272 4.92 10.304 7.428 ;
  LAYER M3 ;
        RECT 10.272 4.94 10.304 4.972 ;
  LAYER M1 ;
        RECT 10.208 4.92 10.24 7.428 ;
  LAYER M3 ;
        RECT 10.208 7.376 10.24 7.408 ;
  LAYER M1 ;
        RECT 10.144 4.92 10.176 7.428 ;
  LAYER M3 ;
        RECT 10.144 4.94 10.176 4.972 ;
  LAYER M1 ;
        RECT 10.08 4.92 10.112 7.428 ;
  LAYER M3 ;
        RECT 10.08 7.376 10.112 7.408 ;
  LAYER M1 ;
        RECT 10.016 4.92 10.048 7.428 ;
  LAYER M3 ;
        RECT 12.384 5.004 12.416 5.036 ;
  LAYER M2 ;
        RECT 10.016 5.068 10.048 5.1 ;
  LAYER M2 ;
        RECT 12.384 5.132 12.416 5.164 ;
  LAYER M2 ;
        RECT 10.016 5.196 10.048 5.228 ;
  LAYER M2 ;
        RECT 12.384 5.26 12.416 5.292 ;
  LAYER M2 ;
        RECT 10.016 5.324 10.048 5.356 ;
  LAYER M2 ;
        RECT 12.384 5.388 12.416 5.42 ;
  LAYER M2 ;
        RECT 10.016 5.452 10.048 5.484 ;
  LAYER M2 ;
        RECT 12.384 5.516 12.416 5.548 ;
  LAYER M2 ;
        RECT 10.016 5.58 10.048 5.612 ;
  LAYER M2 ;
        RECT 12.384 5.644 12.416 5.676 ;
  LAYER M2 ;
        RECT 10.016 5.708 10.048 5.74 ;
  LAYER M2 ;
        RECT 12.384 5.772 12.416 5.804 ;
  LAYER M2 ;
        RECT 10.016 5.836 10.048 5.868 ;
  LAYER M2 ;
        RECT 12.384 5.9 12.416 5.932 ;
  LAYER M2 ;
        RECT 10.016 5.964 10.048 5.996 ;
  LAYER M2 ;
        RECT 12.384 6.028 12.416 6.06 ;
  LAYER M2 ;
        RECT 10.016 6.092 10.048 6.124 ;
  LAYER M2 ;
        RECT 12.384 6.156 12.416 6.188 ;
  LAYER M2 ;
        RECT 10.016 6.22 10.048 6.252 ;
  LAYER M2 ;
        RECT 12.384 6.284 12.416 6.316 ;
  LAYER M2 ;
        RECT 10.016 6.348 10.048 6.38 ;
  LAYER M2 ;
        RECT 12.384 6.412 12.416 6.444 ;
  LAYER M2 ;
        RECT 10.016 6.476 10.048 6.508 ;
  LAYER M2 ;
        RECT 12.384 6.54 12.416 6.572 ;
  LAYER M2 ;
        RECT 10.016 6.604 10.048 6.636 ;
  LAYER M2 ;
        RECT 12.384 6.668 12.416 6.7 ;
  LAYER M2 ;
        RECT 10.016 6.732 10.048 6.764 ;
  LAYER M2 ;
        RECT 12.384 6.796 12.416 6.828 ;
  LAYER M2 ;
        RECT 10.016 6.86 10.048 6.892 ;
  LAYER M2 ;
        RECT 12.384 6.924 12.416 6.956 ;
  LAYER M2 ;
        RECT 10.016 6.988 10.048 7.02 ;
  LAYER M2 ;
        RECT 12.384 7.052 12.416 7.084 ;
  LAYER M2 ;
        RECT 10.016 7.116 10.048 7.148 ;
  LAYER M2 ;
        RECT 12.384 7.18 12.416 7.212 ;
  LAYER M2 ;
        RECT 10.016 7.244 10.048 7.276 ;
  LAYER M2 ;
        RECT 9.968 4.872 12.464 7.476 ;
  LAYER M1 ;
        RECT 12.384 8.028 12.416 10.536 ;
  LAYER M3 ;
        RECT 12.384 10.484 12.416 10.516 ;
  LAYER M1 ;
        RECT 12.32 8.028 12.352 10.536 ;
  LAYER M3 ;
        RECT 12.32 8.048 12.352 8.08 ;
  LAYER M1 ;
        RECT 12.256 8.028 12.288 10.536 ;
  LAYER M3 ;
        RECT 12.256 10.484 12.288 10.516 ;
  LAYER M1 ;
        RECT 12.192 8.028 12.224 10.536 ;
  LAYER M3 ;
        RECT 12.192 8.048 12.224 8.08 ;
  LAYER M1 ;
        RECT 12.128 8.028 12.16 10.536 ;
  LAYER M3 ;
        RECT 12.128 10.484 12.16 10.516 ;
  LAYER M1 ;
        RECT 12.064 8.028 12.096 10.536 ;
  LAYER M3 ;
        RECT 12.064 8.048 12.096 8.08 ;
  LAYER M1 ;
        RECT 12 8.028 12.032 10.536 ;
  LAYER M3 ;
        RECT 12 10.484 12.032 10.516 ;
  LAYER M1 ;
        RECT 11.936 8.028 11.968 10.536 ;
  LAYER M3 ;
        RECT 11.936 8.048 11.968 8.08 ;
  LAYER M1 ;
        RECT 11.872 8.028 11.904 10.536 ;
  LAYER M3 ;
        RECT 11.872 10.484 11.904 10.516 ;
  LAYER M1 ;
        RECT 11.808 8.028 11.84 10.536 ;
  LAYER M3 ;
        RECT 11.808 8.048 11.84 8.08 ;
  LAYER M1 ;
        RECT 11.744 8.028 11.776 10.536 ;
  LAYER M3 ;
        RECT 11.744 10.484 11.776 10.516 ;
  LAYER M1 ;
        RECT 11.68 8.028 11.712 10.536 ;
  LAYER M3 ;
        RECT 11.68 8.048 11.712 8.08 ;
  LAYER M1 ;
        RECT 11.616 8.028 11.648 10.536 ;
  LAYER M3 ;
        RECT 11.616 10.484 11.648 10.516 ;
  LAYER M1 ;
        RECT 11.552 8.028 11.584 10.536 ;
  LAYER M3 ;
        RECT 11.552 8.048 11.584 8.08 ;
  LAYER M1 ;
        RECT 11.488 8.028 11.52 10.536 ;
  LAYER M3 ;
        RECT 11.488 10.484 11.52 10.516 ;
  LAYER M1 ;
        RECT 11.424 8.028 11.456 10.536 ;
  LAYER M3 ;
        RECT 11.424 8.048 11.456 8.08 ;
  LAYER M1 ;
        RECT 11.36 8.028 11.392 10.536 ;
  LAYER M3 ;
        RECT 11.36 10.484 11.392 10.516 ;
  LAYER M1 ;
        RECT 11.296 8.028 11.328 10.536 ;
  LAYER M3 ;
        RECT 11.296 8.048 11.328 8.08 ;
  LAYER M1 ;
        RECT 11.232 8.028 11.264 10.536 ;
  LAYER M3 ;
        RECT 11.232 10.484 11.264 10.516 ;
  LAYER M1 ;
        RECT 11.168 8.028 11.2 10.536 ;
  LAYER M3 ;
        RECT 11.168 8.048 11.2 8.08 ;
  LAYER M1 ;
        RECT 11.104 8.028 11.136 10.536 ;
  LAYER M3 ;
        RECT 11.104 10.484 11.136 10.516 ;
  LAYER M1 ;
        RECT 11.04 8.028 11.072 10.536 ;
  LAYER M3 ;
        RECT 11.04 8.048 11.072 8.08 ;
  LAYER M1 ;
        RECT 10.976 8.028 11.008 10.536 ;
  LAYER M3 ;
        RECT 10.976 10.484 11.008 10.516 ;
  LAYER M1 ;
        RECT 10.912 8.028 10.944 10.536 ;
  LAYER M3 ;
        RECT 10.912 8.048 10.944 8.08 ;
  LAYER M1 ;
        RECT 10.848 8.028 10.88 10.536 ;
  LAYER M3 ;
        RECT 10.848 10.484 10.88 10.516 ;
  LAYER M1 ;
        RECT 10.784 8.028 10.816 10.536 ;
  LAYER M3 ;
        RECT 10.784 8.048 10.816 8.08 ;
  LAYER M1 ;
        RECT 10.72 8.028 10.752 10.536 ;
  LAYER M3 ;
        RECT 10.72 10.484 10.752 10.516 ;
  LAYER M1 ;
        RECT 10.656 8.028 10.688 10.536 ;
  LAYER M3 ;
        RECT 10.656 8.048 10.688 8.08 ;
  LAYER M1 ;
        RECT 10.592 8.028 10.624 10.536 ;
  LAYER M3 ;
        RECT 10.592 10.484 10.624 10.516 ;
  LAYER M1 ;
        RECT 10.528 8.028 10.56 10.536 ;
  LAYER M3 ;
        RECT 10.528 8.048 10.56 8.08 ;
  LAYER M1 ;
        RECT 10.464 8.028 10.496 10.536 ;
  LAYER M3 ;
        RECT 10.464 10.484 10.496 10.516 ;
  LAYER M1 ;
        RECT 10.4 8.028 10.432 10.536 ;
  LAYER M3 ;
        RECT 10.4 8.048 10.432 8.08 ;
  LAYER M1 ;
        RECT 10.336 8.028 10.368 10.536 ;
  LAYER M3 ;
        RECT 10.336 10.484 10.368 10.516 ;
  LAYER M1 ;
        RECT 10.272 8.028 10.304 10.536 ;
  LAYER M3 ;
        RECT 10.272 8.048 10.304 8.08 ;
  LAYER M1 ;
        RECT 10.208 8.028 10.24 10.536 ;
  LAYER M3 ;
        RECT 10.208 10.484 10.24 10.516 ;
  LAYER M1 ;
        RECT 10.144 8.028 10.176 10.536 ;
  LAYER M3 ;
        RECT 10.144 8.048 10.176 8.08 ;
  LAYER M1 ;
        RECT 10.08 8.028 10.112 10.536 ;
  LAYER M3 ;
        RECT 10.08 10.484 10.112 10.516 ;
  LAYER M1 ;
        RECT 10.016 8.028 10.048 10.536 ;
  LAYER M3 ;
        RECT 12.384 8.112 12.416 8.144 ;
  LAYER M2 ;
        RECT 10.016 8.176 10.048 8.208 ;
  LAYER M2 ;
        RECT 12.384 8.24 12.416 8.272 ;
  LAYER M2 ;
        RECT 10.016 8.304 10.048 8.336 ;
  LAYER M2 ;
        RECT 12.384 8.368 12.416 8.4 ;
  LAYER M2 ;
        RECT 10.016 8.432 10.048 8.464 ;
  LAYER M2 ;
        RECT 12.384 8.496 12.416 8.528 ;
  LAYER M2 ;
        RECT 10.016 8.56 10.048 8.592 ;
  LAYER M2 ;
        RECT 12.384 8.624 12.416 8.656 ;
  LAYER M2 ;
        RECT 10.016 8.688 10.048 8.72 ;
  LAYER M2 ;
        RECT 12.384 8.752 12.416 8.784 ;
  LAYER M2 ;
        RECT 10.016 8.816 10.048 8.848 ;
  LAYER M2 ;
        RECT 12.384 8.88 12.416 8.912 ;
  LAYER M2 ;
        RECT 10.016 8.944 10.048 8.976 ;
  LAYER M2 ;
        RECT 12.384 9.008 12.416 9.04 ;
  LAYER M2 ;
        RECT 10.016 9.072 10.048 9.104 ;
  LAYER M2 ;
        RECT 12.384 9.136 12.416 9.168 ;
  LAYER M2 ;
        RECT 10.016 9.2 10.048 9.232 ;
  LAYER M2 ;
        RECT 12.384 9.264 12.416 9.296 ;
  LAYER M2 ;
        RECT 10.016 9.328 10.048 9.36 ;
  LAYER M2 ;
        RECT 12.384 9.392 12.416 9.424 ;
  LAYER M2 ;
        RECT 10.016 9.456 10.048 9.488 ;
  LAYER M2 ;
        RECT 12.384 9.52 12.416 9.552 ;
  LAYER M2 ;
        RECT 10.016 9.584 10.048 9.616 ;
  LAYER M2 ;
        RECT 12.384 9.648 12.416 9.68 ;
  LAYER M2 ;
        RECT 10.016 9.712 10.048 9.744 ;
  LAYER M2 ;
        RECT 12.384 9.776 12.416 9.808 ;
  LAYER M2 ;
        RECT 10.016 9.84 10.048 9.872 ;
  LAYER M2 ;
        RECT 12.384 9.904 12.416 9.936 ;
  LAYER M2 ;
        RECT 10.016 9.968 10.048 10 ;
  LAYER M2 ;
        RECT 12.384 10.032 12.416 10.064 ;
  LAYER M2 ;
        RECT 10.016 10.096 10.048 10.128 ;
  LAYER M2 ;
        RECT 12.384 10.16 12.416 10.192 ;
  LAYER M2 ;
        RECT 10.016 10.224 10.048 10.256 ;
  LAYER M2 ;
        RECT 12.384 10.288 12.416 10.32 ;
  LAYER M2 ;
        RECT 10.016 10.352 10.048 10.384 ;
  LAYER M2 ;
        RECT 9.968 7.98 12.464 10.584 ;
  LAYER M1 ;
        RECT 12.384 11.136 12.416 13.644 ;
  LAYER M3 ;
        RECT 12.384 13.592 12.416 13.624 ;
  LAYER M1 ;
        RECT 12.32 11.136 12.352 13.644 ;
  LAYER M3 ;
        RECT 12.32 11.156 12.352 11.188 ;
  LAYER M1 ;
        RECT 12.256 11.136 12.288 13.644 ;
  LAYER M3 ;
        RECT 12.256 13.592 12.288 13.624 ;
  LAYER M1 ;
        RECT 12.192 11.136 12.224 13.644 ;
  LAYER M3 ;
        RECT 12.192 11.156 12.224 11.188 ;
  LAYER M1 ;
        RECT 12.128 11.136 12.16 13.644 ;
  LAYER M3 ;
        RECT 12.128 13.592 12.16 13.624 ;
  LAYER M1 ;
        RECT 12.064 11.136 12.096 13.644 ;
  LAYER M3 ;
        RECT 12.064 11.156 12.096 11.188 ;
  LAYER M1 ;
        RECT 12 11.136 12.032 13.644 ;
  LAYER M3 ;
        RECT 12 13.592 12.032 13.624 ;
  LAYER M1 ;
        RECT 11.936 11.136 11.968 13.644 ;
  LAYER M3 ;
        RECT 11.936 11.156 11.968 11.188 ;
  LAYER M1 ;
        RECT 11.872 11.136 11.904 13.644 ;
  LAYER M3 ;
        RECT 11.872 13.592 11.904 13.624 ;
  LAYER M1 ;
        RECT 11.808 11.136 11.84 13.644 ;
  LAYER M3 ;
        RECT 11.808 11.156 11.84 11.188 ;
  LAYER M1 ;
        RECT 11.744 11.136 11.776 13.644 ;
  LAYER M3 ;
        RECT 11.744 13.592 11.776 13.624 ;
  LAYER M1 ;
        RECT 11.68 11.136 11.712 13.644 ;
  LAYER M3 ;
        RECT 11.68 11.156 11.712 11.188 ;
  LAYER M1 ;
        RECT 11.616 11.136 11.648 13.644 ;
  LAYER M3 ;
        RECT 11.616 13.592 11.648 13.624 ;
  LAYER M1 ;
        RECT 11.552 11.136 11.584 13.644 ;
  LAYER M3 ;
        RECT 11.552 11.156 11.584 11.188 ;
  LAYER M1 ;
        RECT 11.488 11.136 11.52 13.644 ;
  LAYER M3 ;
        RECT 11.488 13.592 11.52 13.624 ;
  LAYER M1 ;
        RECT 11.424 11.136 11.456 13.644 ;
  LAYER M3 ;
        RECT 11.424 11.156 11.456 11.188 ;
  LAYER M1 ;
        RECT 11.36 11.136 11.392 13.644 ;
  LAYER M3 ;
        RECT 11.36 13.592 11.392 13.624 ;
  LAYER M1 ;
        RECT 11.296 11.136 11.328 13.644 ;
  LAYER M3 ;
        RECT 11.296 11.156 11.328 11.188 ;
  LAYER M1 ;
        RECT 11.232 11.136 11.264 13.644 ;
  LAYER M3 ;
        RECT 11.232 13.592 11.264 13.624 ;
  LAYER M1 ;
        RECT 11.168 11.136 11.2 13.644 ;
  LAYER M3 ;
        RECT 11.168 11.156 11.2 11.188 ;
  LAYER M1 ;
        RECT 11.104 11.136 11.136 13.644 ;
  LAYER M3 ;
        RECT 11.104 13.592 11.136 13.624 ;
  LAYER M1 ;
        RECT 11.04 11.136 11.072 13.644 ;
  LAYER M3 ;
        RECT 11.04 11.156 11.072 11.188 ;
  LAYER M1 ;
        RECT 10.976 11.136 11.008 13.644 ;
  LAYER M3 ;
        RECT 10.976 13.592 11.008 13.624 ;
  LAYER M1 ;
        RECT 10.912 11.136 10.944 13.644 ;
  LAYER M3 ;
        RECT 10.912 11.156 10.944 11.188 ;
  LAYER M1 ;
        RECT 10.848 11.136 10.88 13.644 ;
  LAYER M3 ;
        RECT 10.848 13.592 10.88 13.624 ;
  LAYER M1 ;
        RECT 10.784 11.136 10.816 13.644 ;
  LAYER M3 ;
        RECT 10.784 11.156 10.816 11.188 ;
  LAYER M1 ;
        RECT 10.72 11.136 10.752 13.644 ;
  LAYER M3 ;
        RECT 10.72 13.592 10.752 13.624 ;
  LAYER M1 ;
        RECT 10.656 11.136 10.688 13.644 ;
  LAYER M3 ;
        RECT 10.656 11.156 10.688 11.188 ;
  LAYER M1 ;
        RECT 10.592 11.136 10.624 13.644 ;
  LAYER M3 ;
        RECT 10.592 13.592 10.624 13.624 ;
  LAYER M1 ;
        RECT 10.528 11.136 10.56 13.644 ;
  LAYER M3 ;
        RECT 10.528 11.156 10.56 11.188 ;
  LAYER M1 ;
        RECT 10.464 11.136 10.496 13.644 ;
  LAYER M3 ;
        RECT 10.464 13.592 10.496 13.624 ;
  LAYER M1 ;
        RECT 10.4 11.136 10.432 13.644 ;
  LAYER M3 ;
        RECT 10.4 11.156 10.432 11.188 ;
  LAYER M1 ;
        RECT 10.336 11.136 10.368 13.644 ;
  LAYER M3 ;
        RECT 10.336 13.592 10.368 13.624 ;
  LAYER M1 ;
        RECT 10.272 11.136 10.304 13.644 ;
  LAYER M3 ;
        RECT 10.272 11.156 10.304 11.188 ;
  LAYER M1 ;
        RECT 10.208 11.136 10.24 13.644 ;
  LAYER M3 ;
        RECT 10.208 13.592 10.24 13.624 ;
  LAYER M1 ;
        RECT 10.144 11.136 10.176 13.644 ;
  LAYER M3 ;
        RECT 10.144 11.156 10.176 11.188 ;
  LAYER M1 ;
        RECT 10.08 11.136 10.112 13.644 ;
  LAYER M3 ;
        RECT 10.08 13.592 10.112 13.624 ;
  LAYER M1 ;
        RECT 10.016 11.136 10.048 13.644 ;
  LAYER M3 ;
        RECT 12.384 11.22 12.416 11.252 ;
  LAYER M2 ;
        RECT 10.016 11.284 10.048 11.316 ;
  LAYER M2 ;
        RECT 12.384 11.348 12.416 11.38 ;
  LAYER M2 ;
        RECT 10.016 11.412 10.048 11.444 ;
  LAYER M2 ;
        RECT 12.384 11.476 12.416 11.508 ;
  LAYER M2 ;
        RECT 10.016 11.54 10.048 11.572 ;
  LAYER M2 ;
        RECT 12.384 11.604 12.416 11.636 ;
  LAYER M2 ;
        RECT 10.016 11.668 10.048 11.7 ;
  LAYER M2 ;
        RECT 12.384 11.732 12.416 11.764 ;
  LAYER M2 ;
        RECT 10.016 11.796 10.048 11.828 ;
  LAYER M2 ;
        RECT 12.384 11.86 12.416 11.892 ;
  LAYER M2 ;
        RECT 10.016 11.924 10.048 11.956 ;
  LAYER M2 ;
        RECT 12.384 11.988 12.416 12.02 ;
  LAYER M2 ;
        RECT 10.016 12.052 10.048 12.084 ;
  LAYER M2 ;
        RECT 12.384 12.116 12.416 12.148 ;
  LAYER M2 ;
        RECT 10.016 12.18 10.048 12.212 ;
  LAYER M2 ;
        RECT 12.384 12.244 12.416 12.276 ;
  LAYER M2 ;
        RECT 10.016 12.308 10.048 12.34 ;
  LAYER M2 ;
        RECT 12.384 12.372 12.416 12.404 ;
  LAYER M2 ;
        RECT 10.016 12.436 10.048 12.468 ;
  LAYER M2 ;
        RECT 12.384 12.5 12.416 12.532 ;
  LAYER M2 ;
        RECT 10.016 12.564 10.048 12.596 ;
  LAYER M2 ;
        RECT 12.384 12.628 12.416 12.66 ;
  LAYER M2 ;
        RECT 10.016 12.692 10.048 12.724 ;
  LAYER M2 ;
        RECT 12.384 12.756 12.416 12.788 ;
  LAYER M2 ;
        RECT 10.016 12.82 10.048 12.852 ;
  LAYER M2 ;
        RECT 12.384 12.884 12.416 12.916 ;
  LAYER M2 ;
        RECT 10.016 12.948 10.048 12.98 ;
  LAYER M2 ;
        RECT 12.384 13.012 12.416 13.044 ;
  LAYER M2 ;
        RECT 10.016 13.076 10.048 13.108 ;
  LAYER M2 ;
        RECT 12.384 13.14 12.416 13.172 ;
  LAYER M2 ;
        RECT 10.016 13.204 10.048 13.236 ;
  LAYER M2 ;
        RECT 12.384 13.268 12.416 13.3 ;
  LAYER M2 ;
        RECT 10.016 13.332 10.048 13.364 ;
  LAYER M2 ;
        RECT 12.384 13.396 12.416 13.428 ;
  LAYER M2 ;
        RECT 10.016 13.46 10.048 13.492 ;
  LAYER M2 ;
        RECT 9.968 11.088 12.464 13.692 ;
  LAYER M1 ;
        RECT 9.408 1.812 9.44 4.32 ;
  LAYER M3 ;
        RECT 9.408 4.268 9.44 4.3 ;
  LAYER M1 ;
        RECT 9.344 1.812 9.376 4.32 ;
  LAYER M3 ;
        RECT 9.344 1.832 9.376 1.864 ;
  LAYER M1 ;
        RECT 9.28 1.812 9.312 4.32 ;
  LAYER M3 ;
        RECT 9.28 4.268 9.312 4.3 ;
  LAYER M1 ;
        RECT 9.216 1.812 9.248 4.32 ;
  LAYER M3 ;
        RECT 9.216 1.832 9.248 1.864 ;
  LAYER M1 ;
        RECT 9.152 1.812 9.184 4.32 ;
  LAYER M3 ;
        RECT 9.152 4.268 9.184 4.3 ;
  LAYER M1 ;
        RECT 9.088 1.812 9.12 4.32 ;
  LAYER M3 ;
        RECT 9.088 1.832 9.12 1.864 ;
  LAYER M1 ;
        RECT 9.024 1.812 9.056 4.32 ;
  LAYER M3 ;
        RECT 9.024 4.268 9.056 4.3 ;
  LAYER M1 ;
        RECT 8.96 1.812 8.992 4.32 ;
  LAYER M3 ;
        RECT 8.96 1.832 8.992 1.864 ;
  LAYER M1 ;
        RECT 8.896 1.812 8.928 4.32 ;
  LAYER M3 ;
        RECT 8.896 4.268 8.928 4.3 ;
  LAYER M1 ;
        RECT 8.832 1.812 8.864 4.32 ;
  LAYER M3 ;
        RECT 8.832 1.832 8.864 1.864 ;
  LAYER M1 ;
        RECT 8.768 1.812 8.8 4.32 ;
  LAYER M3 ;
        RECT 8.768 4.268 8.8 4.3 ;
  LAYER M1 ;
        RECT 8.704 1.812 8.736 4.32 ;
  LAYER M3 ;
        RECT 8.704 1.832 8.736 1.864 ;
  LAYER M1 ;
        RECT 8.64 1.812 8.672 4.32 ;
  LAYER M3 ;
        RECT 8.64 4.268 8.672 4.3 ;
  LAYER M1 ;
        RECT 8.576 1.812 8.608 4.32 ;
  LAYER M3 ;
        RECT 8.576 1.832 8.608 1.864 ;
  LAYER M1 ;
        RECT 8.512 1.812 8.544 4.32 ;
  LAYER M3 ;
        RECT 8.512 4.268 8.544 4.3 ;
  LAYER M1 ;
        RECT 8.448 1.812 8.48 4.32 ;
  LAYER M3 ;
        RECT 8.448 1.832 8.48 1.864 ;
  LAYER M1 ;
        RECT 8.384 1.812 8.416 4.32 ;
  LAYER M3 ;
        RECT 8.384 4.268 8.416 4.3 ;
  LAYER M1 ;
        RECT 8.32 1.812 8.352 4.32 ;
  LAYER M3 ;
        RECT 8.32 1.832 8.352 1.864 ;
  LAYER M1 ;
        RECT 8.256 1.812 8.288 4.32 ;
  LAYER M3 ;
        RECT 8.256 4.268 8.288 4.3 ;
  LAYER M1 ;
        RECT 8.192 1.812 8.224 4.32 ;
  LAYER M3 ;
        RECT 8.192 1.832 8.224 1.864 ;
  LAYER M1 ;
        RECT 8.128 1.812 8.16 4.32 ;
  LAYER M3 ;
        RECT 8.128 4.268 8.16 4.3 ;
  LAYER M1 ;
        RECT 8.064 1.812 8.096 4.32 ;
  LAYER M3 ;
        RECT 8.064 1.832 8.096 1.864 ;
  LAYER M1 ;
        RECT 8 1.812 8.032 4.32 ;
  LAYER M3 ;
        RECT 8 4.268 8.032 4.3 ;
  LAYER M1 ;
        RECT 7.936 1.812 7.968 4.32 ;
  LAYER M3 ;
        RECT 7.936 1.832 7.968 1.864 ;
  LAYER M1 ;
        RECT 7.872 1.812 7.904 4.32 ;
  LAYER M3 ;
        RECT 7.872 4.268 7.904 4.3 ;
  LAYER M1 ;
        RECT 7.808 1.812 7.84 4.32 ;
  LAYER M3 ;
        RECT 7.808 1.832 7.84 1.864 ;
  LAYER M1 ;
        RECT 7.744 1.812 7.776 4.32 ;
  LAYER M3 ;
        RECT 7.744 4.268 7.776 4.3 ;
  LAYER M1 ;
        RECT 7.68 1.812 7.712 4.32 ;
  LAYER M3 ;
        RECT 7.68 1.832 7.712 1.864 ;
  LAYER M1 ;
        RECT 7.616 1.812 7.648 4.32 ;
  LAYER M3 ;
        RECT 7.616 4.268 7.648 4.3 ;
  LAYER M1 ;
        RECT 7.552 1.812 7.584 4.32 ;
  LAYER M3 ;
        RECT 7.552 1.832 7.584 1.864 ;
  LAYER M1 ;
        RECT 7.488 1.812 7.52 4.32 ;
  LAYER M3 ;
        RECT 7.488 4.268 7.52 4.3 ;
  LAYER M1 ;
        RECT 7.424 1.812 7.456 4.32 ;
  LAYER M3 ;
        RECT 7.424 1.832 7.456 1.864 ;
  LAYER M1 ;
        RECT 7.36 1.812 7.392 4.32 ;
  LAYER M3 ;
        RECT 7.36 4.268 7.392 4.3 ;
  LAYER M1 ;
        RECT 7.296 1.812 7.328 4.32 ;
  LAYER M3 ;
        RECT 7.296 1.832 7.328 1.864 ;
  LAYER M1 ;
        RECT 7.232 1.812 7.264 4.32 ;
  LAYER M3 ;
        RECT 7.232 4.268 7.264 4.3 ;
  LAYER M1 ;
        RECT 7.168 1.812 7.2 4.32 ;
  LAYER M3 ;
        RECT 7.168 1.832 7.2 1.864 ;
  LAYER M1 ;
        RECT 7.104 1.812 7.136 4.32 ;
  LAYER M3 ;
        RECT 7.104 4.268 7.136 4.3 ;
  LAYER M1 ;
        RECT 7.04 1.812 7.072 4.32 ;
  LAYER M3 ;
        RECT 9.408 1.896 9.44 1.928 ;
  LAYER M2 ;
        RECT 7.04 1.96 7.072 1.992 ;
  LAYER M2 ;
        RECT 9.408 2.024 9.44 2.056 ;
  LAYER M2 ;
        RECT 7.04 2.088 7.072 2.12 ;
  LAYER M2 ;
        RECT 9.408 2.152 9.44 2.184 ;
  LAYER M2 ;
        RECT 7.04 2.216 7.072 2.248 ;
  LAYER M2 ;
        RECT 9.408 2.28 9.44 2.312 ;
  LAYER M2 ;
        RECT 7.04 2.344 7.072 2.376 ;
  LAYER M2 ;
        RECT 9.408 2.408 9.44 2.44 ;
  LAYER M2 ;
        RECT 7.04 2.472 7.072 2.504 ;
  LAYER M2 ;
        RECT 9.408 2.536 9.44 2.568 ;
  LAYER M2 ;
        RECT 7.04 2.6 7.072 2.632 ;
  LAYER M2 ;
        RECT 9.408 2.664 9.44 2.696 ;
  LAYER M2 ;
        RECT 7.04 2.728 7.072 2.76 ;
  LAYER M2 ;
        RECT 9.408 2.792 9.44 2.824 ;
  LAYER M2 ;
        RECT 7.04 2.856 7.072 2.888 ;
  LAYER M2 ;
        RECT 9.408 2.92 9.44 2.952 ;
  LAYER M2 ;
        RECT 7.04 2.984 7.072 3.016 ;
  LAYER M2 ;
        RECT 9.408 3.048 9.44 3.08 ;
  LAYER M2 ;
        RECT 7.04 3.112 7.072 3.144 ;
  LAYER M2 ;
        RECT 9.408 3.176 9.44 3.208 ;
  LAYER M2 ;
        RECT 7.04 3.24 7.072 3.272 ;
  LAYER M2 ;
        RECT 9.408 3.304 9.44 3.336 ;
  LAYER M2 ;
        RECT 7.04 3.368 7.072 3.4 ;
  LAYER M2 ;
        RECT 9.408 3.432 9.44 3.464 ;
  LAYER M2 ;
        RECT 7.04 3.496 7.072 3.528 ;
  LAYER M2 ;
        RECT 9.408 3.56 9.44 3.592 ;
  LAYER M2 ;
        RECT 7.04 3.624 7.072 3.656 ;
  LAYER M2 ;
        RECT 9.408 3.688 9.44 3.72 ;
  LAYER M2 ;
        RECT 7.04 3.752 7.072 3.784 ;
  LAYER M2 ;
        RECT 9.408 3.816 9.44 3.848 ;
  LAYER M2 ;
        RECT 7.04 3.88 7.072 3.912 ;
  LAYER M2 ;
        RECT 9.408 3.944 9.44 3.976 ;
  LAYER M2 ;
        RECT 7.04 4.008 7.072 4.04 ;
  LAYER M2 ;
        RECT 9.408 4.072 9.44 4.104 ;
  LAYER M2 ;
        RECT 7.04 4.136 7.072 4.168 ;
  LAYER M2 ;
        RECT 6.992 1.764 9.488 4.368 ;
  LAYER M1 ;
        RECT 9.408 4.92 9.44 7.428 ;
  LAYER M3 ;
        RECT 9.408 7.376 9.44 7.408 ;
  LAYER M1 ;
        RECT 9.344 4.92 9.376 7.428 ;
  LAYER M3 ;
        RECT 9.344 4.94 9.376 4.972 ;
  LAYER M1 ;
        RECT 9.28 4.92 9.312 7.428 ;
  LAYER M3 ;
        RECT 9.28 7.376 9.312 7.408 ;
  LAYER M1 ;
        RECT 9.216 4.92 9.248 7.428 ;
  LAYER M3 ;
        RECT 9.216 4.94 9.248 4.972 ;
  LAYER M1 ;
        RECT 9.152 4.92 9.184 7.428 ;
  LAYER M3 ;
        RECT 9.152 7.376 9.184 7.408 ;
  LAYER M1 ;
        RECT 9.088 4.92 9.12 7.428 ;
  LAYER M3 ;
        RECT 9.088 4.94 9.12 4.972 ;
  LAYER M1 ;
        RECT 9.024 4.92 9.056 7.428 ;
  LAYER M3 ;
        RECT 9.024 7.376 9.056 7.408 ;
  LAYER M1 ;
        RECT 8.96 4.92 8.992 7.428 ;
  LAYER M3 ;
        RECT 8.96 4.94 8.992 4.972 ;
  LAYER M1 ;
        RECT 8.896 4.92 8.928 7.428 ;
  LAYER M3 ;
        RECT 8.896 7.376 8.928 7.408 ;
  LAYER M1 ;
        RECT 8.832 4.92 8.864 7.428 ;
  LAYER M3 ;
        RECT 8.832 4.94 8.864 4.972 ;
  LAYER M1 ;
        RECT 8.768 4.92 8.8 7.428 ;
  LAYER M3 ;
        RECT 8.768 7.376 8.8 7.408 ;
  LAYER M1 ;
        RECT 8.704 4.92 8.736 7.428 ;
  LAYER M3 ;
        RECT 8.704 4.94 8.736 4.972 ;
  LAYER M1 ;
        RECT 8.64 4.92 8.672 7.428 ;
  LAYER M3 ;
        RECT 8.64 7.376 8.672 7.408 ;
  LAYER M1 ;
        RECT 8.576 4.92 8.608 7.428 ;
  LAYER M3 ;
        RECT 8.576 4.94 8.608 4.972 ;
  LAYER M1 ;
        RECT 8.512 4.92 8.544 7.428 ;
  LAYER M3 ;
        RECT 8.512 7.376 8.544 7.408 ;
  LAYER M1 ;
        RECT 8.448 4.92 8.48 7.428 ;
  LAYER M3 ;
        RECT 8.448 4.94 8.48 4.972 ;
  LAYER M1 ;
        RECT 8.384 4.92 8.416 7.428 ;
  LAYER M3 ;
        RECT 8.384 7.376 8.416 7.408 ;
  LAYER M1 ;
        RECT 8.32 4.92 8.352 7.428 ;
  LAYER M3 ;
        RECT 8.32 4.94 8.352 4.972 ;
  LAYER M1 ;
        RECT 8.256 4.92 8.288 7.428 ;
  LAYER M3 ;
        RECT 8.256 7.376 8.288 7.408 ;
  LAYER M1 ;
        RECT 8.192 4.92 8.224 7.428 ;
  LAYER M3 ;
        RECT 8.192 4.94 8.224 4.972 ;
  LAYER M1 ;
        RECT 8.128 4.92 8.16 7.428 ;
  LAYER M3 ;
        RECT 8.128 7.376 8.16 7.408 ;
  LAYER M1 ;
        RECT 8.064 4.92 8.096 7.428 ;
  LAYER M3 ;
        RECT 8.064 4.94 8.096 4.972 ;
  LAYER M1 ;
        RECT 8 4.92 8.032 7.428 ;
  LAYER M3 ;
        RECT 8 7.376 8.032 7.408 ;
  LAYER M1 ;
        RECT 7.936 4.92 7.968 7.428 ;
  LAYER M3 ;
        RECT 7.936 4.94 7.968 4.972 ;
  LAYER M1 ;
        RECT 7.872 4.92 7.904 7.428 ;
  LAYER M3 ;
        RECT 7.872 7.376 7.904 7.408 ;
  LAYER M1 ;
        RECT 7.808 4.92 7.84 7.428 ;
  LAYER M3 ;
        RECT 7.808 4.94 7.84 4.972 ;
  LAYER M1 ;
        RECT 7.744 4.92 7.776 7.428 ;
  LAYER M3 ;
        RECT 7.744 7.376 7.776 7.408 ;
  LAYER M1 ;
        RECT 7.68 4.92 7.712 7.428 ;
  LAYER M3 ;
        RECT 7.68 4.94 7.712 4.972 ;
  LAYER M1 ;
        RECT 7.616 4.92 7.648 7.428 ;
  LAYER M3 ;
        RECT 7.616 7.376 7.648 7.408 ;
  LAYER M1 ;
        RECT 7.552 4.92 7.584 7.428 ;
  LAYER M3 ;
        RECT 7.552 4.94 7.584 4.972 ;
  LAYER M1 ;
        RECT 7.488 4.92 7.52 7.428 ;
  LAYER M3 ;
        RECT 7.488 7.376 7.52 7.408 ;
  LAYER M1 ;
        RECT 7.424 4.92 7.456 7.428 ;
  LAYER M3 ;
        RECT 7.424 4.94 7.456 4.972 ;
  LAYER M1 ;
        RECT 7.36 4.92 7.392 7.428 ;
  LAYER M3 ;
        RECT 7.36 7.376 7.392 7.408 ;
  LAYER M1 ;
        RECT 7.296 4.92 7.328 7.428 ;
  LAYER M3 ;
        RECT 7.296 4.94 7.328 4.972 ;
  LAYER M1 ;
        RECT 7.232 4.92 7.264 7.428 ;
  LAYER M3 ;
        RECT 7.232 7.376 7.264 7.408 ;
  LAYER M1 ;
        RECT 7.168 4.92 7.2 7.428 ;
  LAYER M3 ;
        RECT 7.168 4.94 7.2 4.972 ;
  LAYER M1 ;
        RECT 7.104 4.92 7.136 7.428 ;
  LAYER M3 ;
        RECT 7.104 7.376 7.136 7.408 ;
  LAYER M1 ;
        RECT 7.04 4.92 7.072 7.428 ;
  LAYER M3 ;
        RECT 9.408 5.004 9.44 5.036 ;
  LAYER M2 ;
        RECT 7.04 5.068 7.072 5.1 ;
  LAYER M2 ;
        RECT 9.408 5.132 9.44 5.164 ;
  LAYER M2 ;
        RECT 7.04 5.196 7.072 5.228 ;
  LAYER M2 ;
        RECT 9.408 5.26 9.44 5.292 ;
  LAYER M2 ;
        RECT 7.04 5.324 7.072 5.356 ;
  LAYER M2 ;
        RECT 9.408 5.388 9.44 5.42 ;
  LAYER M2 ;
        RECT 7.04 5.452 7.072 5.484 ;
  LAYER M2 ;
        RECT 9.408 5.516 9.44 5.548 ;
  LAYER M2 ;
        RECT 7.04 5.58 7.072 5.612 ;
  LAYER M2 ;
        RECT 9.408 5.644 9.44 5.676 ;
  LAYER M2 ;
        RECT 7.04 5.708 7.072 5.74 ;
  LAYER M2 ;
        RECT 9.408 5.772 9.44 5.804 ;
  LAYER M2 ;
        RECT 7.04 5.836 7.072 5.868 ;
  LAYER M2 ;
        RECT 9.408 5.9 9.44 5.932 ;
  LAYER M2 ;
        RECT 7.04 5.964 7.072 5.996 ;
  LAYER M2 ;
        RECT 9.408 6.028 9.44 6.06 ;
  LAYER M2 ;
        RECT 7.04 6.092 7.072 6.124 ;
  LAYER M2 ;
        RECT 9.408 6.156 9.44 6.188 ;
  LAYER M2 ;
        RECT 7.04 6.22 7.072 6.252 ;
  LAYER M2 ;
        RECT 9.408 6.284 9.44 6.316 ;
  LAYER M2 ;
        RECT 7.04 6.348 7.072 6.38 ;
  LAYER M2 ;
        RECT 9.408 6.412 9.44 6.444 ;
  LAYER M2 ;
        RECT 7.04 6.476 7.072 6.508 ;
  LAYER M2 ;
        RECT 9.408 6.54 9.44 6.572 ;
  LAYER M2 ;
        RECT 7.04 6.604 7.072 6.636 ;
  LAYER M2 ;
        RECT 9.408 6.668 9.44 6.7 ;
  LAYER M2 ;
        RECT 7.04 6.732 7.072 6.764 ;
  LAYER M2 ;
        RECT 9.408 6.796 9.44 6.828 ;
  LAYER M2 ;
        RECT 7.04 6.86 7.072 6.892 ;
  LAYER M2 ;
        RECT 9.408 6.924 9.44 6.956 ;
  LAYER M2 ;
        RECT 7.04 6.988 7.072 7.02 ;
  LAYER M2 ;
        RECT 9.408 7.052 9.44 7.084 ;
  LAYER M2 ;
        RECT 7.04 7.116 7.072 7.148 ;
  LAYER M2 ;
        RECT 9.408 7.18 9.44 7.212 ;
  LAYER M2 ;
        RECT 7.04 7.244 7.072 7.276 ;
  LAYER M2 ;
        RECT 6.992 4.872 9.488 7.476 ;
  LAYER M1 ;
        RECT 9.408 8.028 9.44 10.536 ;
  LAYER M3 ;
        RECT 9.408 10.484 9.44 10.516 ;
  LAYER M1 ;
        RECT 9.344 8.028 9.376 10.536 ;
  LAYER M3 ;
        RECT 9.344 8.048 9.376 8.08 ;
  LAYER M1 ;
        RECT 9.28 8.028 9.312 10.536 ;
  LAYER M3 ;
        RECT 9.28 10.484 9.312 10.516 ;
  LAYER M1 ;
        RECT 9.216 8.028 9.248 10.536 ;
  LAYER M3 ;
        RECT 9.216 8.048 9.248 8.08 ;
  LAYER M1 ;
        RECT 9.152 8.028 9.184 10.536 ;
  LAYER M3 ;
        RECT 9.152 10.484 9.184 10.516 ;
  LAYER M1 ;
        RECT 9.088 8.028 9.12 10.536 ;
  LAYER M3 ;
        RECT 9.088 8.048 9.12 8.08 ;
  LAYER M1 ;
        RECT 9.024 8.028 9.056 10.536 ;
  LAYER M3 ;
        RECT 9.024 10.484 9.056 10.516 ;
  LAYER M1 ;
        RECT 8.96 8.028 8.992 10.536 ;
  LAYER M3 ;
        RECT 8.96 8.048 8.992 8.08 ;
  LAYER M1 ;
        RECT 8.896 8.028 8.928 10.536 ;
  LAYER M3 ;
        RECT 8.896 10.484 8.928 10.516 ;
  LAYER M1 ;
        RECT 8.832 8.028 8.864 10.536 ;
  LAYER M3 ;
        RECT 8.832 8.048 8.864 8.08 ;
  LAYER M1 ;
        RECT 8.768 8.028 8.8 10.536 ;
  LAYER M3 ;
        RECT 8.768 10.484 8.8 10.516 ;
  LAYER M1 ;
        RECT 8.704 8.028 8.736 10.536 ;
  LAYER M3 ;
        RECT 8.704 8.048 8.736 8.08 ;
  LAYER M1 ;
        RECT 8.64 8.028 8.672 10.536 ;
  LAYER M3 ;
        RECT 8.64 10.484 8.672 10.516 ;
  LAYER M1 ;
        RECT 8.576 8.028 8.608 10.536 ;
  LAYER M3 ;
        RECT 8.576 8.048 8.608 8.08 ;
  LAYER M1 ;
        RECT 8.512 8.028 8.544 10.536 ;
  LAYER M3 ;
        RECT 8.512 10.484 8.544 10.516 ;
  LAYER M1 ;
        RECT 8.448 8.028 8.48 10.536 ;
  LAYER M3 ;
        RECT 8.448 8.048 8.48 8.08 ;
  LAYER M1 ;
        RECT 8.384 8.028 8.416 10.536 ;
  LAYER M3 ;
        RECT 8.384 10.484 8.416 10.516 ;
  LAYER M1 ;
        RECT 8.32 8.028 8.352 10.536 ;
  LAYER M3 ;
        RECT 8.32 8.048 8.352 8.08 ;
  LAYER M1 ;
        RECT 8.256 8.028 8.288 10.536 ;
  LAYER M3 ;
        RECT 8.256 10.484 8.288 10.516 ;
  LAYER M1 ;
        RECT 8.192 8.028 8.224 10.536 ;
  LAYER M3 ;
        RECT 8.192 8.048 8.224 8.08 ;
  LAYER M1 ;
        RECT 8.128 8.028 8.16 10.536 ;
  LAYER M3 ;
        RECT 8.128 10.484 8.16 10.516 ;
  LAYER M1 ;
        RECT 8.064 8.028 8.096 10.536 ;
  LAYER M3 ;
        RECT 8.064 8.048 8.096 8.08 ;
  LAYER M1 ;
        RECT 8 8.028 8.032 10.536 ;
  LAYER M3 ;
        RECT 8 10.484 8.032 10.516 ;
  LAYER M1 ;
        RECT 7.936 8.028 7.968 10.536 ;
  LAYER M3 ;
        RECT 7.936 8.048 7.968 8.08 ;
  LAYER M1 ;
        RECT 7.872 8.028 7.904 10.536 ;
  LAYER M3 ;
        RECT 7.872 10.484 7.904 10.516 ;
  LAYER M1 ;
        RECT 7.808 8.028 7.84 10.536 ;
  LAYER M3 ;
        RECT 7.808 8.048 7.84 8.08 ;
  LAYER M1 ;
        RECT 7.744 8.028 7.776 10.536 ;
  LAYER M3 ;
        RECT 7.744 10.484 7.776 10.516 ;
  LAYER M1 ;
        RECT 7.68 8.028 7.712 10.536 ;
  LAYER M3 ;
        RECT 7.68 8.048 7.712 8.08 ;
  LAYER M1 ;
        RECT 7.616 8.028 7.648 10.536 ;
  LAYER M3 ;
        RECT 7.616 10.484 7.648 10.516 ;
  LAYER M1 ;
        RECT 7.552 8.028 7.584 10.536 ;
  LAYER M3 ;
        RECT 7.552 8.048 7.584 8.08 ;
  LAYER M1 ;
        RECT 7.488 8.028 7.52 10.536 ;
  LAYER M3 ;
        RECT 7.488 10.484 7.52 10.516 ;
  LAYER M1 ;
        RECT 7.424 8.028 7.456 10.536 ;
  LAYER M3 ;
        RECT 7.424 8.048 7.456 8.08 ;
  LAYER M1 ;
        RECT 7.36 8.028 7.392 10.536 ;
  LAYER M3 ;
        RECT 7.36 10.484 7.392 10.516 ;
  LAYER M1 ;
        RECT 7.296 8.028 7.328 10.536 ;
  LAYER M3 ;
        RECT 7.296 8.048 7.328 8.08 ;
  LAYER M1 ;
        RECT 7.232 8.028 7.264 10.536 ;
  LAYER M3 ;
        RECT 7.232 10.484 7.264 10.516 ;
  LAYER M1 ;
        RECT 7.168 8.028 7.2 10.536 ;
  LAYER M3 ;
        RECT 7.168 8.048 7.2 8.08 ;
  LAYER M1 ;
        RECT 7.104 8.028 7.136 10.536 ;
  LAYER M3 ;
        RECT 7.104 10.484 7.136 10.516 ;
  LAYER M1 ;
        RECT 7.04 8.028 7.072 10.536 ;
  LAYER M3 ;
        RECT 9.408 8.112 9.44 8.144 ;
  LAYER M2 ;
        RECT 7.04 8.176 7.072 8.208 ;
  LAYER M2 ;
        RECT 9.408 8.24 9.44 8.272 ;
  LAYER M2 ;
        RECT 7.04 8.304 7.072 8.336 ;
  LAYER M2 ;
        RECT 9.408 8.368 9.44 8.4 ;
  LAYER M2 ;
        RECT 7.04 8.432 7.072 8.464 ;
  LAYER M2 ;
        RECT 9.408 8.496 9.44 8.528 ;
  LAYER M2 ;
        RECT 7.04 8.56 7.072 8.592 ;
  LAYER M2 ;
        RECT 9.408 8.624 9.44 8.656 ;
  LAYER M2 ;
        RECT 7.04 8.688 7.072 8.72 ;
  LAYER M2 ;
        RECT 9.408 8.752 9.44 8.784 ;
  LAYER M2 ;
        RECT 7.04 8.816 7.072 8.848 ;
  LAYER M2 ;
        RECT 9.408 8.88 9.44 8.912 ;
  LAYER M2 ;
        RECT 7.04 8.944 7.072 8.976 ;
  LAYER M2 ;
        RECT 9.408 9.008 9.44 9.04 ;
  LAYER M2 ;
        RECT 7.04 9.072 7.072 9.104 ;
  LAYER M2 ;
        RECT 9.408 9.136 9.44 9.168 ;
  LAYER M2 ;
        RECT 7.04 9.2 7.072 9.232 ;
  LAYER M2 ;
        RECT 9.408 9.264 9.44 9.296 ;
  LAYER M2 ;
        RECT 7.04 9.328 7.072 9.36 ;
  LAYER M2 ;
        RECT 9.408 9.392 9.44 9.424 ;
  LAYER M2 ;
        RECT 7.04 9.456 7.072 9.488 ;
  LAYER M2 ;
        RECT 9.408 9.52 9.44 9.552 ;
  LAYER M2 ;
        RECT 7.04 9.584 7.072 9.616 ;
  LAYER M2 ;
        RECT 9.408 9.648 9.44 9.68 ;
  LAYER M2 ;
        RECT 7.04 9.712 7.072 9.744 ;
  LAYER M2 ;
        RECT 9.408 9.776 9.44 9.808 ;
  LAYER M2 ;
        RECT 7.04 9.84 7.072 9.872 ;
  LAYER M2 ;
        RECT 9.408 9.904 9.44 9.936 ;
  LAYER M2 ;
        RECT 7.04 9.968 7.072 10 ;
  LAYER M2 ;
        RECT 9.408 10.032 9.44 10.064 ;
  LAYER M2 ;
        RECT 7.04 10.096 7.072 10.128 ;
  LAYER M2 ;
        RECT 9.408 10.16 9.44 10.192 ;
  LAYER M2 ;
        RECT 7.04 10.224 7.072 10.256 ;
  LAYER M2 ;
        RECT 9.408 10.288 9.44 10.32 ;
  LAYER M2 ;
        RECT 7.04 10.352 7.072 10.384 ;
  LAYER M2 ;
        RECT 6.992 7.98 9.488 10.584 ;
  LAYER M1 ;
        RECT 9.408 11.136 9.44 13.644 ;
  LAYER M3 ;
        RECT 9.408 13.592 9.44 13.624 ;
  LAYER M1 ;
        RECT 9.344 11.136 9.376 13.644 ;
  LAYER M3 ;
        RECT 9.344 11.156 9.376 11.188 ;
  LAYER M1 ;
        RECT 9.28 11.136 9.312 13.644 ;
  LAYER M3 ;
        RECT 9.28 13.592 9.312 13.624 ;
  LAYER M1 ;
        RECT 9.216 11.136 9.248 13.644 ;
  LAYER M3 ;
        RECT 9.216 11.156 9.248 11.188 ;
  LAYER M1 ;
        RECT 9.152 11.136 9.184 13.644 ;
  LAYER M3 ;
        RECT 9.152 13.592 9.184 13.624 ;
  LAYER M1 ;
        RECT 9.088 11.136 9.12 13.644 ;
  LAYER M3 ;
        RECT 9.088 11.156 9.12 11.188 ;
  LAYER M1 ;
        RECT 9.024 11.136 9.056 13.644 ;
  LAYER M3 ;
        RECT 9.024 13.592 9.056 13.624 ;
  LAYER M1 ;
        RECT 8.96 11.136 8.992 13.644 ;
  LAYER M3 ;
        RECT 8.96 11.156 8.992 11.188 ;
  LAYER M1 ;
        RECT 8.896 11.136 8.928 13.644 ;
  LAYER M3 ;
        RECT 8.896 13.592 8.928 13.624 ;
  LAYER M1 ;
        RECT 8.832 11.136 8.864 13.644 ;
  LAYER M3 ;
        RECT 8.832 11.156 8.864 11.188 ;
  LAYER M1 ;
        RECT 8.768 11.136 8.8 13.644 ;
  LAYER M3 ;
        RECT 8.768 13.592 8.8 13.624 ;
  LAYER M1 ;
        RECT 8.704 11.136 8.736 13.644 ;
  LAYER M3 ;
        RECT 8.704 11.156 8.736 11.188 ;
  LAYER M1 ;
        RECT 8.64 11.136 8.672 13.644 ;
  LAYER M3 ;
        RECT 8.64 13.592 8.672 13.624 ;
  LAYER M1 ;
        RECT 8.576 11.136 8.608 13.644 ;
  LAYER M3 ;
        RECT 8.576 11.156 8.608 11.188 ;
  LAYER M1 ;
        RECT 8.512 11.136 8.544 13.644 ;
  LAYER M3 ;
        RECT 8.512 13.592 8.544 13.624 ;
  LAYER M1 ;
        RECT 8.448 11.136 8.48 13.644 ;
  LAYER M3 ;
        RECT 8.448 11.156 8.48 11.188 ;
  LAYER M1 ;
        RECT 8.384 11.136 8.416 13.644 ;
  LAYER M3 ;
        RECT 8.384 13.592 8.416 13.624 ;
  LAYER M1 ;
        RECT 8.32 11.136 8.352 13.644 ;
  LAYER M3 ;
        RECT 8.32 11.156 8.352 11.188 ;
  LAYER M1 ;
        RECT 8.256 11.136 8.288 13.644 ;
  LAYER M3 ;
        RECT 8.256 13.592 8.288 13.624 ;
  LAYER M1 ;
        RECT 8.192 11.136 8.224 13.644 ;
  LAYER M3 ;
        RECT 8.192 11.156 8.224 11.188 ;
  LAYER M1 ;
        RECT 8.128 11.136 8.16 13.644 ;
  LAYER M3 ;
        RECT 8.128 13.592 8.16 13.624 ;
  LAYER M1 ;
        RECT 8.064 11.136 8.096 13.644 ;
  LAYER M3 ;
        RECT 8.064 11.156 8.096 11.188 ;
  LAYER M1 ;
        RECT 8 11.136 8.032 13.644 ;
  LAYER M3 ;
        RECT 8 13.592 8.032 13.624 ;
  LAYER M1 ;
        RECT 7.936 11.136 7.968 13.644 ;
  LAYER M3 ;
        RECT 7.936 11.156 7.968 11.188 ;
  LAYER M1 ;
        RECT 7.872 11.136 7.904 13.644 ;
  LAYER M3 ;
        RECT 7.872 13.592 7.904 13.624 ;
  LAYER M1 ;
        RECT 7.808 11.136 7.84 13.644 ;
  LAYER M3 ;
        RECT 7.808 11.156 7.84 11.188 ;
  LAYER M1 ;
        RECT 7.744 11.136 7.776 13.644 ;
  LAYER M3 ;
        RECT 7.744 13.592 7.776 13.624 ;
  LAYER M1 ;
        RECT 7.68 11.136 7.712 13.644 ;
  LAYER M3 ;
        RECT 7.68 11.156 7.712 11.188 ;
  LAYER M1 ;
        RECT 7.616 11.136 7.648 13.644 ;
  LAYER M3 ;
        RECT 7.616 13.592 7.648 13.624 ;
  LAYER M1 ;
        RECT 7.552 11.136 7.584 13.644 ;
  LAYER M3 ;
        RECT 7.552 11.156 7.584 11.188 ;
  LAYER M1 ;
        RECT 7.488 11.136 7.52 13.644 ;
  LAYER M3 ;
        RECT 7.488 13.592 7.52 13.624 ;
  LAYER M1 ;
        RECT 7.424 11.136 7.456 13.644 ;
  LAYER M3 ;
        RECT 7.424 11.156 7.456 11.188 ;
  LAYER M1 ;
        RECT 7.36 11.136 7.392 13.644 ;
  LAYER M3 ;
        RECT 7.36 13.592 7.392 13.624 ;
  LAYER M1 ;
        RECT 7.296 11.136 7.328 13.644 ;
  LAYER M3 ;
        RECT 7.296 11.156 7.328 11.188 ;
  LAYER M1 ;
        RECT 7.232 11.136 7.264 13.644 ;
  LAYER M3 ;
        RECT 7.232 13.592 7.264 13.624 ;
  LAYER M1 ;
        RECT 7.168 11.136 7.2 13.644 ;
  LAYER M3 ;
        RECT 7.168 11.156 7.2 11.188 ;
  LAYER M1 ;
        RECT 7.104 11.136 7.136 13.644 ;
  LAYER M3 ;
        RECT 7.104 13.592 7.136 13.624 ;
  LAYER M1 ;
        RECT 7.04 11.136 7.072 13.644 ;
  LAYER M3 ;
        RECT 9.408 11.22 9.44 11.252 ;
  LAYER M2 ;
        RECT 7.04 11.284 7.072 11.316 ;
  LAYER M2 ;
        RECT 9.408 11.348 9.44 11.38 ;
  LAYER M2 ;
        RECT 7.04 11.412 7.072 11.444 ;
  LAYER M2 ;
        RECT 9.408 11.476 9.44 11.508 ;
  LAYER M2 ;
        RECT 7.04 11.54 7.072 11.572 ;
  LAYER M2 ;
        RECT 9.408 11.604 9.44 11.636 ;
  LAYER M2 ;
        RECT 7.04 11.668 7.072 11.7 ;
  LAYER M2 ;
        RECT 9.408 11.732 9.44 11.764 ;
  LAYER M2 ;
        RECT 7.04 11.796 7.072 11.828 ;
  LAYER M2 ;
        RECT 9.408 11.86 9.44 11.892 ;
  LAYER M2 ;
        RECT 7.04 11.924 7.072 11.956 ;
  LAYER M2 ;
        RECT 9.408 11.988 9.44 12.02 ;
  LAYER M2 ;
        RECT 7.04 12.052 7.072 12.084 ;
  LAYER M2 ;
        RECT 9.408 12.116 9.44 12.148 ;
  LAYER M2 ;
        RECT 7.04 12.18 7.072 12.212 ;
  LAYER M2 ;
        RECT 9.408 12.244 9.44 12.276 ;
  LAYER M2 ;
        RECT 7.04 12.308 7.072 12.34 ;
  LAYER M2 ;
        RECT 9.408 12.372 9.44 12.404 ;
  LAYER M2 ;
        RECT 7.04 12.436 7.072 12.468 ;
  LAYER M2 ;
        RECT 9.408 12.5 9.44 12.532 ;
  LAYER M2 ;
        RECT 7.04 12.564 7.072 12.596 ;
  LAYER M2 ;
        RECT 9.408 12.628 9.44 12.66 ;
  LAYER M2 ;
        RECT 7.04 12.692 7.072 12.724 ;
  LAYER M2 ;
        RECT 9.408 12.756 9.44 12.788 ;
  LAYER M2 ;
        RECT 7.04 12.82 7.072 12.852 ;
  LAYER M2 ;
        RECT 9.408 12.884 9.44 12.916 ;
  LAYER M2 ;
        RECT 7.04 12.948 7.072 12.98 ;
  LAYER M2 ;
        RECT 9.408 13.012 9.44 13.044 ;
  LAYER M2 ;
        RECT 7.04 13.076 7.072 13.108 ;
  LAYER M2 ;
        RECT 9.408 13.14 9.44 13.172 ;
  LAYER M2 ;
        RECT 7.04 13.204 7.072 13.236 ;
  LAYER M2 ;
        RECT 9.408 13.268 9.44 13.3 ;
  LAYER M2 ;
        RECT 7.04 13.332 7.072 13.364 ;
  LAYER M2 ;
        RECT 9.408 13.396 9.44 13.428 ;
  LAYER M2 ;
        RECT 7.04 13.46 7.072 13.492 ;
  LAYER M2 ;
        RECT 6.992 11.088 9.488 13.692 ;
  LAYER M1 ;
        RECT 6.432 1.812 6.464 4.32 ;
  LAYER M3 ;
        RECT 6.432 4.268 6.464 4.3 ;
  LAYER M1 ;
        RECT 6.368 1.812 6.4 4.32 ;
  LAYER M3 ;
        RECT 6.368 1.832 6.4 1.864 ;
  LAYER M1 ;
        RECT 6.304 1.812 6.336 4.32 ;
  LAYER M3 ;
        RECT 6.304 4.268 6.336 4.3 ;
  LAYER M1 ;
        RECT 6.24 1.812 6.272 4.32 ;
  LAYER M3 ;
        RECT 6.24 1.832 6.272 1.864 ;
  LAYER M1 ;
        RECT 6.176 1.812 6.208 4.32 ;
  LAYER M3 ;
        RECT 6.176 4.268 6.208 4.3 ;
  LAYER M1 ;
        RECT 6.112 1.812 6.144 4.32 ;
  LAYER M3 ;
        RECT 6.112 1.832 6.144 1.864 ;
  LAYER M1 ;
        RECT 6.048 1.812 6.08 4.32 ;
  LAYER M3 ;
        RECT 6.048 4.268 6.08 4.3 ;
  LAYER M1 ;
        RECT 5.984 1.812 6.016 4.32 ;
  LAYER M3 ;
        RECT 5.984 1.832 6.016 1.864 ;
  LAYER M1 ;
        RECT 5.92 1.812 5.952 4.32 ;
  LAYER M3 ;
        RECT 5.92 4.268 5.952 4.3 ;
  LAYER M1 ;
        RECT 5.856 1.812 5.888 4.32 ;
  LAYER M3 ;
        RECT 5.856 1.832 5.888 1.864 ;
  LAYER M1 ;
        RECT 5.792 1.812 5.824 4.32 ;
  LAYER M3 ;
        RECT 5.792 4.268 5.824 4.3 ;
  LAYER M1 ;
        RECT 5.728 1.812 5.76 4.32 ;
  LAYER M3 ;
        RECT 5.728 1.832 5.76 1.864 ;
  LAYER M1 ;
        RECT 5.664 1.812 5.696 4.32 ;
  LAYER M3 ;
        RECT 5.664 4.268 5.696 4.3 ;
  LAYER M1 ;
        RECT 5.6 1.812 5.632 4.32 ;
  LAYER M3 ;
        RECT 5.6 1.832 5.632 1.864 ;
  LAYER M1 ;
        RECT 5.536 1.812 5.568 4.32 ;
  LAYER M3 ;
        RECT 5.536 4.268 5.568 4.3 ;
  LAYER M1 ;
        RECT 5.472 1.812 5.504 4.32 ;
  LAYER M3 ;
        RECT 5.472 1.832 5.504 1.864 ;
  LAYER M1 ;
        RECT 5.408 1.812 5.44 4.32 ;
  LAYER M3 ;
        RECT 5.408 4.268 5.44 4.3 ;
  LAYER M1 ;
        RECT 5.344 1.812 5.376 4.32 ;
  LAYER M3 ;
        RECT 5.344 1.832 5.376 1.864 ;
  LAYER M1 ;
        RECT 5.28 1.812 5.312 4.32 ;
  LAYER M3 ;
        RECT 5.28 4.268 5.312 4.3 ;
  LAYER M1 ;
        RECT 5.216 1.812 5.248 4.32 ;
  LAYER M3 ;
        RECT 5.216 1.832 5.248 1.864 ;
  LAYER M1 ;
        RECT 5.152 1.812 5.184 4.32 ;
  LAYER M3 ;
        RECT 5.152 4.268 5.184 4.3 ;
  LAYER M1 ;
        RECT 5.088 1.812 5.12 4.32 ;
  LAYER M3 ;
        RECT 5.088 1.832 5.12 1.864 ;
  LAYER M1 ;
        RECT 5.024 1.812 5.056 4.32 ;
  LAYER M3 ;
        RECT 5.024 4.268 5.056 4.3 ;
  LAYER M1 ;
        RECT 4.96 1.812 4.992 4.32 ;
  LAYER M3 ;
        RECT 4.96 1.832 4.992 1.864 ;
  LAYER M1 ;
        RECT 4.896 1.812 4.928 4.32 ;
  LAYER M3 ;
        RECT 4.896 4.268 4.928 4.3 ;
  LAYER M1 ;
        RECT 4.832 1.812 4.864 4.32 ;
  LAYER M3 ;
        RECT 4.832 1.832 4.864 1.864 ;
  LAYER M1 ;
        RECT 4.768 1.812 4.8 4.32 ;
  LAYER M3 ;
        RECT 4.768 4.268 4.8 4.3 ;
  LAYER M1 ;
        RECT 4.704 1.812 4.736 4.32 ;
  LAYER M3 ;
        RECT 4.704 1.832 4.736 1.864 ;
  LAYER M1 ;
        RECT 4.64 1.812 4.672 4.32 ;
  LAYER M3 ;
        RECT 4.64 4.268 4.672 4.3 ;
  LAYER M1 ;
        RECT 4.576 1.812 4.608 4.32 ;
  LAYER M3 ;
        RECT 4.576 1.832 4.608 1.864 ;
  LAYER M1 ;
        RECT 4.512 1.812 4.544 4.32 ;
  LAYER M3 ;
        RECT 4.512 4.268 4.544 4.3 ;
  LAYER M1 ;
        RECT 4.448 1.812 4.48 4.32 ;
  LAYER M3 ;
        RECT 4.448 1.832 4.48 1.864 ;
  LAYER M1 ;
        RECT 4.384 1.812 4.416 4.32 ;
  LAYER M3 ;
        RECT 4.384 4.268 4.416 4.3 ;
  LAYER M1 ;
        RECT 4.32 1.812 4.352 4.32 ;
  LAYER M3 ;
        RECT 4.32 1.832 4.352 1.864 ;
  LAYER M1 ;
        RECT 4.256 1.812 4.288 4.32 ;
  LAYER M3 ;
        RECT 4.256 4.268 4.288 4.3 ;
  LAYER M1 ;
        RECT 4.192 1.812 4.224 4.32 ;
  LAYER M3 ;
        RECT 4.192 1.832 4.224 1.864 ;
  LAYER M1 ;
        RECT 4.128 1.812 4.16 4.32 ;
  LAYER M3 ;
        RECT 4.128 4.268 4.16 4.3 ;
  LAYER M1 ;
        RECT 4.064 1.812 4.096 4.32 ;
  LAYER M3 ;
        RECT 6.432 1.896 6.464 1.928 ;
  LAYER M2 ;
        RECT 4.064 1.96 4.096 1.992 ;
  LAYER M2 ;
        RECT 6.432 2.024 6.464 2.056 ;
  LAYER M2 ;
        RECT 4.064 2.088 4.096 2.12 ;
  LAYER M2 ;
        RECT 6.432 2.152 6.464 2.184 ;
  LAYER M2 ;
        RECT 4.064 2.216 4.096 2.248 ;
  LAYER M2 ;
        RECT 6.432 2.28 6.464 2.312 ;
  LAYER M2 ;
        RECT 4.064 2.344 4.096 2.376 ;
  LAYER M2 ;
        RECT 6.432 2.408 6.464 2.44 ;
  LAYER M2 ;
        RECT 4.064 2.472 4.096 2.504 ;
  LAYER M2 ;
        RECT 6.432 2.536 6.464 2.568 ;
  LAYER M2 ;
        RECT 4.064 2.6 4.096 2.632 ;
  LAYER M2 ;
        RECT 6.432 2.664 6.464 2.696 ;
  LAYER M2 ;
        RECT 4.064 2.728 4.096 2.76 ;
  LAYER M2 ;
        RECT 6.432 2.792 6.464 2.824 ;
  LAYER M2 ;
        RECT 4.064 2.856 4.096 2.888 ;
  LAYER M2 ;
        RECT 6.432 2.92 6.464 2.952 ;
  LAYER M2 ;
        RECT 4.064 2.984 4.096 3.016 ;
  LAYER M2 ;
        RECT 6.432 3.048 6.464 3.08 ;
  LAYER M2 ;
        RECT 4.064 3.112 4.096 3.144 ;
  LAYER M2 ;
        RECT 6.432 3.176 6.464 3.208 ;
  LAYER M2 ;
        RECT 4.064 3.24 4.096 3.272 ;
  LAYER M2 ;
        RECT 6.432 3.304 6.464 3.336 ;
  LAYER M2 ;
        RECT 4.064 3.368 4.096 3.4 ;
  LAYER M2 ;
        RECT 6.432 3.432 6.464 3.464 ;
  LAYER M2 ;
        RECT 4.064 3.496 4.096 3.528 ;
  LAYER M2 ;
        RECT 6.432 3.56 6.464 3.592 ;
  LAYER M2 ;
        RECT 4.064 3.624 4.096 3.656 ;
  LAYER M2 ;
        RECT 6.432 3.688 6.464 3.72 ;
  LAYER M2 ;
        RECT 4.064 3.752 4.096 3.784 ;
  LAYER M2 ;
        RECT 6.432 3.816 6.464 3.848 ;
  LAYER M2 ;
        RECT 4.064 3.88 4.096 3.912 ;
  LAYER M2 ;
        RECT 6.432 3.944 6.464 3.976 ;
  LAYER M2 ;
        RECT 4.064 4.008 4.096 4.04 ;
  LAYER M2 ;
        RECT 6.432 4.072 6.464 4.104 ;
  LAYER M2 ;
        RECT 4.064 4.136 4.096 4.168 ;
  LAYER M2 ;
        RECT 4.016 1.764 6.512 4.368 ;
  LAYER M1 ;
        RECT 6.432 4.92 6.464 7.428 ;
  LAYER M3 ;
        RECT 6.432 7.376 6.464 7.408 ;
  LAYER M1 ;
        RECT 6.368 4.92 6.4 7.428 ;
  LAYER M3 ;
        RECT 6.368 4.94 6.4 4.972 ;
  LAYER M1 ;
        RECT 6.304 4.92 6.336 7.428 ;
  LAYER M3 ;
        RECT 6.304 7.376 6.336 7.408 ;
  LAYER M1 ;
        RECT 6.24 4.92 6.272 7.428 ;
  LAYER M3 ;
        RECT 6.24 4.94 6.272 4.972 ;
  LAYER M1 ;
        RECT 6.176 4.92 6.208 7.428 ;
  LAYER M3 ;
        RECT 6.176 7.376 6.208 7.408 ;
  LAYER M1 ;
        RECT 6.112 4.92 6.144 7.428 ;
  LAYER M3 ;
        RECT 6.112 4.94 6.144 4.972 ;
  LAYER M1 ;
        RECT 6.048 4.92 6.08 7.428 ;
  LAYER M3 ;
        RECT 6.048 7.376 6.08 7.408 ;
  LAYER M1 ;
        RECT 5.984 4.92 6.016 7.428 ;
  LAYER M3 ;
        RECT 5.984 4.94 6.016 4.972 ;
  LAYER M1 ;
        RECT 5.92 4.92 5.952 7.428 ;
  LAYER M3 ;
        RECT 5.92 7.376 5.952 7.408 ;
  LAYER M1 ;
        RECT 5.856 4.92 5.888 7.428 ;
  LAYER M3 ;
        RECT 5.856 4.94 5.888 4.972 ;
  LAYER M1 ;
        RECT 5.792 4.92 5.824 7.428 ;
  LAYER M3 ;
        RECT 5.792 7.376 5.824 7.408 ;
  LAYER M1 ;
        RECT 5.728 4.92 5.76 7.428 ;
  LAYER M3 ;
        RECT 5.728 4.94 5.76 4.972 ;
  LAYER M1 ;
        RECT 5.664 4.92 5.696 7.428 ;
  LAYER M3 ;
        RECT 5.664 7.376 5.696 7.408 ;
  LAYER M1 ;
        RECT 5.6 4.92 5.632 7.428 ;
  LAYER M3 ;
        RECT 5.6 4.94 5.632 4.972 ;
  LAYER M1 ;
        RECT 5.536 4.92 5.568 7.428 ;
  LAYER M3 ;
        RECT 5.536 7.376 5.568 7.408 ;
  LAYER M1 ;
        RECT 5.472 4.92 5.504 7.428 ;
  LAYER M3 ;
        RECT 5.472 4.94 5.504 4.972 ;
  LAYER M1 ;
        RECT 5.408 4.92 5.44 7.428 ;
  LAYER M3 ;
        RECT 5.408 7.376 5.44 7.408 ;
  LAYER M1 ;
        RECT 5.344 4.92 5.376 7.428 ;
  LAYER M3 ;
        RECT 5.344 4.94 5.376 4.972 ;
  LAYER M1 ;
        RECT 5.28 4.92 5.312 7.428 ;
  LAYER M3 ;
        RECT 5.28 7.376 5.312 7.408 ;
  LAYER M1 ;
        RECT 5.216 4.92 5.248 7.428 ;
  LAYER M3 ;
        RECT 5.216 4.94 5.248 4.972 ;
  LAYER M1 ;
        RECT 5.152 4.92 5.184 7.428 ;
  LAYER M3 ;
        RECT 5.152 7.376 5.184 7.408 ;
  LAYER M1 ;
        RECT 5.088 4.92 5.12 7.428 ;
  LAYER M3 ;
        RECT 5.088 4.94 5.12 4.972 ;
  LAYER M1 ;
        RECT 5.024 4.92 5.056 7.428 ;
  LAYER M3 ;
        RECT 5.024 7.376 5.056 7.408 ;
  LAYER M1 ;
        RECT 4.96 4.92 4.992 7.428 ;
  LAYER M3 ;
        RECT 4.96 4.94 4.992 4.972 ;
  LAYER M1 ;
        RECT 4.896 4.92 4.928 7.428 ;
  LAYER M3 ;
        RECT 4.896 7.376 4.928 7.408 ;
  LAYER M1 ;
        RECT 4.832 4.92 4.864 7.428 ;
  LAYER M3 ;
        RECT 4.832 4.94 4.864 4.972 ;
  LAYER M1 ;
        RECT 4.768 4.92 4.8 7.428 ;
  LAYER M3 ;
        RECT 4.768 7.376 4.8 7.408 ;
  LAYER M1 ;
        RECT 4.704 4.92 4.736 7.428 ;
  LAYER M3 ;
        RECT 4.704 4.94 4.736 4.972 ;
  LAYER M1 ;
        RECT 4.64 4.92 4.672 7.428 ;
  LAYER M3 ;
        RECT 4.64 7.376 4.672 7.408 ;
  LAYER M1 ;
        RECT 4.576 4.92 4.608 7.428 ;
  LAYER M3 ;
        RECT 4.576 4.94 4.608 4.972 ;
  LAYER M1 ;
        RECT 4.512 4.92 4.544 7.428 ;
  LAYER M3 ;
        RECT 4.512 7.376 4.544 7.408 ;
  LAYER M1 ;
        RECT 4.448 4.92 4.48 7.428 ;
  LAYER M3 ;
        RECT 4.448 4.94 4.48 4.972 ;
  LAYER M1 ;
        RECT 4.384 4.92 4.416 7.428 ;
  LAYER M3 ;
        RECT 4.384 7.376 4.416 7.408 ;
  LAYER M1 ;
        RECT 4.32 4.92 4.352 7.428 ;
  LAYER M3 ;
        RECT 4.32 4.94 4.352 4.972 ;
  LAYER M1 ;
        RECT 4.256 4.92 4.288 7.428 ;
  LAYER M3 ;
        RECT 4.256 7.376 4.288 7.408 ;
  LAYER M1 ;
        RECT 4.192 4.92 4.224 7.428 ;
  LAYER M3 ;
        RECT 4.192 4.94 4.224 4.972 ;
  LAYER M1 ;
        RECT 4.128 4.92 4.16 7.428 ;
  LAYER M3 ;
        RECT 4.128 7.376 4.16 7.408 ;
  LAYER M1 ;
        RECT 4.064 4.92 4.096 7.428 ;
  LAYER M3 ;
        RECT 6.432 5.004 6.464 5.036 ;
  LAYER M2 ;
        RECT 4.064 5.068 4.096 5.1 ;
  LAYER M2 ;
        RECT 6.432 5.132 6.464 5.164 ;
  LAYER M2 ;
        RECT 4.064 5.196 4.096 5.228 ;
  LAYER M2 ;
        RECT 6.432 5.26 6.464 5.292 ;
  LAYER M2 ;
        RECT 4.064 5.324 4.096 5.356 ;
  LAYER M2 ;
        RECT 6.432 5.388 6.464 5.42 ;
  LAYER M2 ;
        RECT 4.064 5.452 4.096 5.484 ;
  LAYER M2 ;
        RECT 6.432 5.516 6.464 5.548 ;
  LAYER M2 ;
        RECT 4.064 5.58 4.096 5.612 ;
  LAYER M2 ;
        RECT 6.432 5.644 6.464 5.676 ;
  LAYER M2 ;
        RECT 4.064 5.708 4.096 5.74 ;
  LAYER M2 ;
        RECT 6.432 5.772 6.464 5.804 ;
  LAYER M2 ;
        RECT 4.064 5.836 4.096 5.868 ;
  LAYER M2 ;
        RECT 6.432 5.9 6.464 5.932 ;
  LAYER M2 ;
        RECT 4.064 5.964 4.096 5.996 ;
  LAYER M2 ;
        RECT 6.432 6.028 6.464 6.06 ;
  LAYER M2 ;
        RECT 4.064 6.092 4.096 6.124 ;
  LAYER M2 ;
        RECT 6.432 6.156 6.464 6.188 ;
  LAYER M2 ;
        RECT 4.064 6.22 4.096 6.252 ;
  LAYER M2 ;
        RECT 6.432 6.284 6.464 6.316 ;
  LAYER M2 ;
        RECT 4.064 6.348 4.096 6.38 ;
  LAYER M2 ;
        RECT 6.432 6.412 6.464 6.444 ;
  LAYER M2 ;
        RECT 4.064 6.476 4.096 6.508 ;
  LAYER M2 ;
        RECT 6.432 6.54 6.464 6.572 ;
  LAYER M2 ;
        RECT 4.064 6.604 4.096 6.636 ;
  LAYER M2 ;
        RECT 6.432 6.668 6.464 6.7 ;
  LAYER M2 ;
        RECT 4.064 6.732 4.096 6.764 ;
  LAYER M2 ;
        RECT 6.432 6.796 6.464 6.828 ;
  LAYER M2 ;
        RECT 4.064 6.86 4.096 6.892 ;
  LAYER M2 ;
        RECT 6.432 6.924 6.464 6.956 ;
  LAYER M2 ;
        RECT 4.064 6.988 4.096 7.02 ;
  LAYER M2 ;
        RECT 6.432 7.052 6.464 7.084 ;
  LAYER M2 ;
        RECT 4.064 7.116 4.096 7.148 ;
  LAYER M2 ;
        RECT 6.432 7.18 6.464 7.212 ;
  LAYER M2 ;
        RECT 4.064 7.244 4.096 7.276 ;
  LAYER M2 ;
        RECT 4.016 4.872 6.512 7.476 ;
  LAYER M1 ;
        RECT 6.432 8.028 6.464 10.536 ;
  LAYER M3 ;
        RECT 6.432 10.484 6.464 10.516 ;
  LAYER M1 ;
        RECT 6.368 8.028 6.4 10.536 ;
  LAYER M3 ;
        RECT 6.368 8.048 6.4 8.08 ;
  LAYER M1 ;
        RECT 6.304 8.028 6.336 10.536 ;
  LAYER M3 ;
        RECT 6.304 10.484 6.336 10.516 ;
  LAYER M1 ;
        RECT 6.24 8.028 6.272 10.536 ;
  LAYER M3 ;
        RECT 6.24 8.048 6.272 8.08 ;
  LAYER M1 ;
        RECT 6.176 8.028 6.208 10.536 ;
  LAYER M3 ;
        RECT 6.176 10.484 6.208 10.516 ;
  LAYER M1 ;
        RECT 6.112 8.028 6.144 10.536 ;
  LAYER M3 ;
        RECT 6.112 8.048 6.144 8.08 ;
  LAYER M1 ;
        RECT 6.048 8.028 6.08 10.536 ;
  LAYER M3 ;
        RECT 6.048 10.484 6.08 10.516 ;
  LAYER M1 ;
        RECT 5.984 8.028 6.016 10.536 ;
  LAYER M3 ;
        RECT 5.984 8.048 6.016 8.08 ;
  LAYER M1 ;
        RECT 5.92 8.028 5.952 10.536 ;
  LAYER M3 ;
        RECT 5.92 10.484 5.952 10.516 ;
  LAYER M1 ;
        RECT 5.856 8.028 5.888 10.536 ;
  LAYER M3 ;
        RECT 5.856 8.048 5.888 8.08 ;
  LAYER M1 ;
        RECT 5.792 8.028 5.824 10.536 ;
  LAYER M3 ;
        RECT 5.792 10.484 5.824 10.516 ;
  LAYER M1 ;
        RECT 5.728 8.028 5.76 10.536 ;
  LAYER M3 ;
        RECT 5.728 8.048 5.76 8.08 ;
  LAYER M1 ;
        RECT 5.664 8.028 5.696 10.536 ;
  LAYER M3 ;
        RECT 5.664 10.484 5.696 10.516 ;
  LAYER M1 ;
        RECT 5.6 8.028 5.632 10.536 ;
  LAYER M3 ;
        RECT 5.6 8.048 5.632 8.08 ;
  LAYER M1 ;
        RECT 5.536 8.028 5.568 10.536 ;
  LAYER M3 ;
        RECT 5.536 10.484 5.568 10.516 ;
  LAYER M1 ;
        RECT 5.472 8.028 5.504 10.536 ;
  LAYER M3 ;
        RECT 5.472 8.048 5.504 8.08 ;
  LAYER M1 ;
        RECT 5.408 8.028 5.44 10.536 ;
  LAYER M3 ;
        RECT 5.408 10.484 5.44 10.516 ;
  LAYER M1 ;
        RECT 5.344 8.028 5.376 10.536 ;
  LAYER M3 ;
        RECT 5.344 8.048 5.376 8.08 ;
  LAYER M1 ;
        RECT 5.28 8.028 5.312 10.536 ;
  LAYER M3 ;
        RECT 5.28 10.484 5.312 10.516 ;
  LAYER M1 ;
        RECT 5.216 8.028 5.248 10.536 ;
  LAYER M3 ;
        RECT 5.216 8.048 5.248 8.08 ;
  LAYER M1 ;
        RECT 5.152 8.028 5.184 10.536 ;
  LAYER M3 ;
        RECT 5.152 10.484 5.184 10.516 ;
  LAYER M1 ;
        RECT 5.088 8.028 5.12 10.536 ;
  LAYER M3 ;
        RECT 5.088 8.048 5.12 8.08 ;
  LAYER M1 ;
        RECT 5.024 8.028 5.056 10.536 ;
  LAYER M3 ;
        RECT 5.024 10.484 5.056 10.516 ;
  LAYER M1 ;
        RECT 4.96 8.028 4.992 10.536 ;
  LAYER M3 ;
        RECT 4.96 8.048 4.992 8.08 ;
  LAYER M1 ;
        RECT 4.896 8.028 4.928 10.536 ;
  LAYER M3 ;
        RECT 4.896 10.484 4.928 10.516 ;
  LAYER M1 ;
        RECT 4.832 8.028 4.864 10.536 ;
  LAYER M3 ;
        RECT 4.832 8.048 4.864 8.08 ;
  LAYER M1 ;
        RECT 4.768 8.028 4.8 10.536 ;
  LAYER M3 ;
        RECT 4.768 10.484 4.8 10.516 ;
  LAYER M1 ;
        RECT 4.704 8.028 4.736 10.536 ;
  LAYER M3 ;
        RECT 4.704 8.048 4.736 8.08 ;
  LAYER M1 ;
        RECT 4.64 8.028 4.672 10.536 ;
  LAYER M3 ;
        RECT 4.64 10.484 4.672 10.516 ;
  LAYER M1 ;
        RECT 4.576 8.028 4.608 10.536 ;
  LAYER M3 ;
        RECT 4.576 8.048 4.608 8.08 ;
  LAYER M1 ;
        RECT 4.512 8.028 4.544 10.536 ;
  LAYER M3 ;
        RECT 4.512 10.484 4.544 10.516 ;
  LAYER M1 ;
        RECT 4.448 8.028 4.48 10.536 ;
  LAYER M3 ;
        RECT 4.448 8.048 4.48 8.08 ;
  LAYER M1 ;
        RECT 4.384 8.028 4.416 10.536 ;
  LAYER M3 ;
        RECT 4.384 10.484 4.416 10.516 ;
  LAYER M1 ;
        RECT 4.32 8.028 4.352 10.536 ;
  LAYER M3 ;
        RECT 4.32 8.048 4.352 8.08 ;
  LAYER M1 ;
        RECT 4.256 8.028 4.288 10.536 ;
  LAYER M3 ;
        RECT 4.256 10.484 4.288 10.516 ;
  LAYER M1 ;
        RECT 4.192 8.028 4.224 10.536 ;
  LAYER M3 ;
        RECT 4.192 8.048 4.224 8.08 ;
  LAYER M1 ;
        RECT 4.128 8.028 4.16 10.536 ;
  LAYER M3 ;
        RECT 4.128 10.484 4.16 10.516 ;
  LAYER M1 ;
        RECT 4.064 8.028 4.096 10.536 ;
  LAYER M3 ;
        RECT 6.432 8.112 6.464 8.144 ;
  LAYER M2 ;
        RECT 4.064 8.176 4.096 8.208 ;
  LAYER M2 ;
        RECT 6.432 8.24 6.464 8.272 ;
  LAYER M2 ;
        RECT 4.064 8.304 4.096 8.336 ;
  LAYER M2 ;
        RECT 6.432 8.368 6.464 8.4 ;
  LAYER M2 ;
        RECT 4.064 8.432 4.096 8.464 ;
  LAYER M2 ;
        RECT 6.432 8.496 6.464 8.528 ;
  LAYER M2 ;
        RECT 4.064 8.56 4.096 8.592 ;
  LAYER M2 ;
        RECT 6.432 8.624 6.464 8.656 ;
  LAYER M2 ;
        RECT 4.064 8.688 4.096 8.72 ;
  LAYER M2 ;
        RECT 6.432 8.752 6.464 8.784 ;
  LAYER M2 ;
        RECT 4.064 8.816 4.096 8.848 ;
  LAYER M2 ;
        RECT 6.432 8.88 6.464 8.912 ;
  LAYER M2 ;
        RECT 4.064 8.944 4.096 8.976 ;
  LAYER M2 ;
        RECT 6.432 9.008 6.464 9.04 ;
  LAYER M2 ;
        RECT 4.064 9.072 4.096 9.104 ;
  LAYER M2 ;
        RECT 6.432 9.136 6.464 9.168 ;
  LAYER M2 ;
        RECT 4.064 9.2 4.096 9.232 ;
  LAYER M2 ;
        RECT 6.432 9.264 6.464 9.296 ;
  LAYER M2 ;
        RECT 4.064 9.328 4.096 9.36 ;
  LAYER M2 ;
        RECT 6.432 9.392 6.464 9.424 ;
  LAYER M2 ;
        RECT 4.064 9.456 4.096 9.488 ;
  LAYER M2 ;
        RECT 6.432 9.52 6.464 9.552 ;
  LAYER M2 ;
        RECT 4.064 9.584 4.096 9.616 ;
  LAYER M2 ;
        RECT 6.432 9.648 6.464 9.68 ;
  LAYER M2 ;
        RECT 4.064 9.712 4.096 9.744 ;
  LAYER M2 ;
        RECT 6.432 9.776 6.464 9.808 ;
  LAYER M2 ;
        RECT 4.064 9.84 4.096 9.872 ;
  LAYER M2 ;
        RECT 6.432 9.904 6.464 9.936 ;
  LAYER M2 ;
        RECT 4.064 9.968 4.096 10 ;
  LAYER M2 ;
        RECT 6.432 10.032 6.464 10.064 ;
  LAYER M2 ;
        RECT 4.064 10.096 4.096 10.128 ;
  LAYER M2 ;
        RECT 6.432 10.16 6.464 10.192 ;
  LAYER M2 ;
        RECT 4.064 10.224 4.096 10.256 ;
  LAYER M2 ;
        RECT 6.432 10.288 6.464 10.32 ;
  LAYER M2 ;
        RECT 4.064 10.352 4.096 10.384 ;
  LAYER M2 ;
        RECT 4.016 7.98 6.512 10.584 ;
  LAYER M1 ;
        RECT 6.432 11.136 6.464 13.644 ;
  LAYER M3 ;
        RECT 6.432 13.592 6.464 13.624 ;
  LAYER M1 ;
        RECT 6.368 11.136 6.4 13.644 ;
  LAYER M3 ;
        RECT 6.368 11.156 6.4 11.188 ;
  LAYER M1 ;
        RECT 6.304 11.136 6.336 13.644 ;
  LAYER M3 ;
        RECT 6.304 13.592 6.336 13.624 ;
  LAYER M1 ;
        RECT 6.24 11.136 6.272 13.644 ;
  LAYER M3 ;
        RECT 6.24 11.156 6.272 11.188 ;
  LAYER M1 ;
        RECT 6.176 11.136 6.208 13.644 ;
  LAYER M3 ;
        RECT 6.176 13.592 6.208 13.624 ;
  LAYER M1 ;
        RECT 6.112 11.136 6.144 13.644 ;
  LAYER M3 ;
        RECT 6.112 11.156 6.144 11.188 ;
  LAYER M1 ;
        RECT 6.048 11.136 6.08 13.644 ;
  LAYER M3 ;
        RECT 6.048 13.592 6.08 13.624 ;
  LAYER M1 ;
        RECT 5.984 11.136 6.016 13.644 ;
  LAYER M3 ;
        RECT 5.984 11.156 6.016 11.188 ;
  LAYER M1 ;
        RECT 5.92 11.136 5.952 13.644 ;
  LAYER M3 ;
        RECT 5.92 13.592 5.952 13.624 ;
  LAYER M1 ;
        RECT 5.856 11.136 5.888 13.644 ;
  LAYER M3 ;
        RECT 5.856 11.156 5.888 11.188 ;
  LAYER M1 ;
        RECT 5.792 11.136 5.824 13.644 ;
  LAYER M3 ;
        RECT 5.792 13.592 5.824 13.624 ;
  LAYER M1 ;
        RECT 5.728 11.136 5.76 13.644 ;
  LAYER M3 ;
        RECT 5.728 11.156 5.76 11.188 ;
  LAYER M1 ;
        RECT 5.664 11.136 5.696 13.644 ;
  LAYER M3 ;
        RECT 5.664 13.592 5.696 13.624 ;
  LAYER M1 ;
        RECT 5.6 11.136 5.632 13.644 ;
  LAYER M3 ;
        RECT 5.6 11.156 5.632 11.188 ;
  LAYER M1 ;
        RECT 5.536 11.136 5.568 13.644 ;
  LAYER M3 ;
        RECT 5.536 13.592 5.568 13.624 ;
  LAYER M1 ;
        RECT 5.472 11.136 5.504 13.644 ;
  LAYER M3 ;
        RECT 5.472 11.156 5.504 11.188 ;
  LAYER M1 ;
        RECT 5.408 11.136 5.44 13.644 ;
  LAYER M3 ;
        RECT 5.408 13.592 5.44 13.624 ;
  LAYER M1 ;
        RECT 5.344 11.136 5.376 13.644 ;
  LAYER M3 ;
        RECT 5.344 11.156 5.376 11.188 ;
  LAYER M1 ;
        RECT 5.28 11.136 5.312 13.644 ;
  LAYER M3 ;
        RECT 5.28 13.592 5.312 13.624 ;
  LAYER M1 ;
        RECT 5.216 11.136 5.248 13.644 ;
  LAYER M3 ;
        RECT 5.216 11.156 5.248 11.188 ;
  LAYER M1 ;
        RECT 5.152 11.136 5.184 13.644 ;
  LAYER M3 ;
        RECT 5.152 13.592 5.184 13.624 ;
  LAYER M1 ;
        RECT 5.088 11.136 5.12 13.644 ;
  LAYER M3 ;
        RECT 5.088 11.156 5.12 11.188 ;
  LAYER M1 ;
        RECT 5.024 11.136 5.056 13.644 ;
  LAYER M3 ;
        RECT 5.024 13.592 5.056 13.624 ;
  LAYER M1 ;
        RECT 4.96 11.136 4.992 13.644 ;
  LAYER M3 ;
        RECT 4.96 11.156 4.992 11.188 ;
  LAYER M1 ;
        RECT 4.896 11.136 4.928 13.644 ;
  LAYER M3 ;
        RECT 4.896 13.592 4.928 13.624 ;
  LAYER M1 ;
        RECT 4.832 11.136 4.864 13.644 ;
  LAYER M3 ;
        RECT 4.832 11.156 4.864 11.188 ;
  LAYER M1 ;
        RECT 4.768 11.136 4.8 13.644 ;
  LAYER M3 ;
        RECT 4.768 13.592 4.8 13.624 ;
  LAYER M1 ;
        RECT 4.704 11.136 4.736 13.644 ;
  LAYER M3 ;
        RECT 4.704 11.156 4.736 11.188 ;
  LAYER M1 ;
        RECT 4.64 11.136 4.672 13.644 ;
  LAYER M3 ;
        RECT 4.64 13.592 4.672 13.624 ;
  LAYER M1 ;
        RECT 4.576 11.136 4.608 13.644 ;
  LAYER M3 ;
        RECT 4.576 11.156 4.608 11.188 ;
  LAYER M1 ;
        RECT 4.512 11.136 4.544 13.644 ;
  LAYER M3 ;
        RECT 4.512 13.592 4.544 13.624 ;
  LAYER M1 ;
        RECT 4.448 11.136 4.48 13.644 ;
  LAYER M3 ;
        RECT 4.448 11.156 4.48 11.188 ;
  LAYER M1 ;
        RECT 4.384 11.136 4.416 13.644 ;
  LAYER M3 ;
        RECT 4.384 13.592 4.416 13.624 ;
  LAYER M1 ;
        RECT 4.32 11.136 4.352 13.644 ;
  LAYER M3 ;
        RECT 4.32 11.156 4.352 11.188 ;
  LAYER M1 ;
        RECT 4.256 11.136 4.288 13.644 ;
  LAYER M3 ;
        RECT 4.256 13.592 4.288 13.624 ;
  LAYER M1 ;
        RECT 4.192 11.136 4.224 13.644 ;
  LAYER M3 ;
        RECT 4.192 11.156 4.224 11.188 ;
  LAYER M1 ;
        RECT 4.128 11.136 4.16 13.644 ;
  LAYER M3 ;
        RECT 4.128 13.592 4.16 13.624 ;
  LAYER M1 ;
        RECT 4.064 11.136 4.096 13.644 ;
  LAYER M3 ;
        RECT 6.432 11.22 6.464 11.252 ;
  LAYER M2 ;
        RECT 4.064 11.284 4.096 11.316 ;
  LAYER M2 ;
        RECT 6.432 11.348 6.464 11.38 ;
  LAYER M2 ;
        RECT 4.064 11.412 4.096 11.444 ;
  LAYER M2 ;
        RECT 6.432 11.476 6.464 11.508 ;
  LAYER M2 ;
        RECT 4.064 11.54 4.096 11.572 ;
  LAYER M2 ;
        RECT 6.432 11.604 6.464 11.636 ;
  LAYER M2 ;
        RECT 4.064 11.668 4.096 11.7 ;
  LAYER M2 ;
        RECT 6.432 11.732 6.464 11.764 ;
  LAYER M2 ;
        RECT 4.064 11.796 4.096 11.828 ;
  LAYER M2 ;
        RECT 6.432 11.86 6.464 11.892 ;
  LAYER M2 ;
        RECT 4.064 11.924 4.096 11.956 ;
  LAYER M2 ;
        RECT 6.432 11.988 6.464 12.02 ;
  LAYER M2 ;
        RECT 4.064 12.052 4.096 12.084 ;
  LAYER M2 ;
        RECT 6.432 12.116 6.464 12.148 ;
  LAYER M2 ;
        RECT 4.064 12.18 4.096 12.212 ;
  LAYER M2 ;
        RECT 6.432 12.244 6.464 12.276 ;
  LAYER M2 ;
        RECT 4.064 12.308 4.096 12.34 ;
  LAYER M2 ;
        RECT 6.432 12.372 6.464 12.404 ;
  LAYER M2 ;
        RECT 4.064 12.436 4.096 12.468 ;
  LAYER M2 ;
        RECT 6.432 12.5 6.464 12.532 ;
  LAYER M2 ;
        RECT 4.064 12.564 4.096 12.596 ;
  LAYER M2 ;
        RECT 6.432 12.628 6.464 12.66 ;
  LAYER M2 ;
        RECT 4.064 12.692 4.096 12.724 ;
  LAYER M2 ;
        RECT 6.432 12.756 6.464 12.788 ;
  LAYER M2 ;
        RECT 4.064 12.82 4.096 12.852 ;
  LAYER M2 ;
        RECT 6.432 12.884 6.464 12.916 ;
  LAYER M2 ;
        RECT 4.064 12.948 4.096 12.98 ;
  LAYER M2 ;
        RECT 6.432 13.012 6.464 13.044 ;
  LAYER M2 ;
        RECT 4.064 13.076 4.096 13.108 ;
  LAYER M2 ;
        RECT 6.432 13.14 6.464 13.172 ;
  LAYER M2 ;
        RECT 4.064 13.204 4.096 13.236 ;
  LAYER M2 ;
        RECT 6.432 13.268 6.464 13.3 ;
  LAYER M2 ;
        RECT 4.064 13.332 4.096 13.364 ;
  LAYER M2 ;
        RECT 6.432 13.396 6.464 13.428 ;
  LAYER M2 ;
        RECT 4.064 13.46 4.096 13.492 ;
  LAYER M2 ;
        RECT 4.016 11.088 6.512 13.692 ;
  LAYER M1 ;
        RECT 3.456 1.812 3.488 4.32 ;
  LAYER M3 ;
        RECT 3.456 4.268 3.488 4.3 ;
  LAYER M1 ;
        RECT 3.392 1.812 3.424 4.32 ;
  LAYER M3 ;
        RECT 3.392 1.832 3.424 1.864 ;
  LAYER M1 ;
        RECT 3.328 1.812 3.36 4.32 ;
  LAYER M3 ;
        RECT 3.328 4.268 3.36 4.3 ;
  LAYER M1 ;
        RECT 3.264 1.812 3.296 4.32 ;
  LAYER M3 ;
        RECT 3.264 1.832 3.296 1.864 ;
  LAYER M1 ;
        RECT 3.2 1.812 3.232 4.32 ;
  LAYER M3 ;
        RECT 3.2 4.268 3.232 4.3 ;
  LAYER M1 ;
        RECT 3.136 1.812 3.168 4.32 ;
  LAYER M3 ;
        RECT 3.136 1.832 3.168 1.864 ;
  LAYER M1 ;
        RECT 3.072 1.812 3.104 4.32 ;
  LAYER M3 ;
        RECT 3.072 4.268 3.104 4.3 ;
  LAYER M1 ;
        RECT 3.008 1.812 3.04 4.32 ;
  LAYER M3 ;
        RECT 3.008 1.832 3.04 1.864 ;
  LAYER M1 ;
        RECT 2.944 1.812 2.976 4.32 ;
  LAYER M3 ;
        RECT 2.944 4.268 2.976 4.3 ;
  LAYER M1 ;
        RECT 2.88 1.812 2.912 4.32 ;
  LAYER M3 ;
        RECT 2.88 1.832 2.912 1.864 ;
  LAYER M1 ;
        RECT 2.816 1.812 2.848 4.32 ;
  LAYER M3 ;
        RECT 2.816 4.268 2.848 4.3 ;
  LAYER M1 ;
        RECT 2.752 1.812 2.784 4.32 ;
  LAYER M3 ;
        RECT 2.752 1.832 2.784 1.864 ;
  LAYER M1 ;
        RECT 2.688 1.812 2.72 4.32 ;
  LAYER M3 ;
        RECT 2.688 4.268 2.72 4.3 ;
  LAYER M1 ;
        RECT 2.624 1.812 2.656 4.32 ;
  LAYER M3 ;
        RECT 2.624 1.832 2.656 1.864 ;
  LAYER M1 ;
        RECT 2.56 1.812 2.592 4.32 ;
  LAYER M3 ;
        RECT 2.56 4.268 2.592 4.3 ;
  LAYER M1 ;
        RECT 2.496 1.812 2.528 4.32 ;
  LAYER M3 ;
        RECT 2.496 1.832 2.528 1.864 ;
  LAYER M1 ;
        RECT 2.432 1.812 2.464 4.32 ;
  LAYER M3 ;
        RECT 2.432 4.268 2.464 4.3 ;
  LAYER M1 ;
        RECT 2.368 1.812 2.4 4.32 ;
  LAYER M3 ;
        RECT 2.368 1.832 2.4 1.864 ;
  LAYER M1 ;
        RECT 2.304 1.812 2.336 4.32 ;
  LAYER M3 ;
        RECT 2.304 4.268 2.336 4.3 ;
  LAYER M1 ;
        RECT 2.24 1.812 2.272 4.32 ;
  LAYER M3 ;
        RECT 2.24 1.832 2.272 1.864 ;
  LAYER M1 ;
        RECT 2.176 1.812 2.208 4.32 ;
  LAYER M3 ;
        RECT 2.176 4.268 2.208 4.3 ;
  LAYER M1 ;
        RECT 2.112 1.812 2.144 4.32 ;
  LAYER M3 ;
        RECT 2.112 1.832 2.144 1.864 ;
  LAYER M1 ;
        RECT 2.048 1.812 2.08 4.32 ;
  LAYER M3 ;
        RECT 2.048 4.268 2.08 4.3 ;
  LAYER M1 ;
        RECT 1.984 1.812 2.016 4.32 ;
  LAYER M3 ;
        RECT 1.984 1.832 2.016 1.864 ;
  LAYER M1 ;
        RECT 1.92 1.812 1.952 4.32 ;
  LAYER M3 ;
        RECT 1.92 4.268 1.952 4.3 ;
  LAYER M1 ;
        RECT 1.856 1.812 1.888 4.32 ;
  LAYER M3 ;
        RECT 1.856 1.832 1.888 1.864 ;
  LAYER M1 ;
        RECT 1.792 1.812 1.824 4.32 ;
  LAYER M3 ;
        RECT 1.792 4.268 1.824 4.3 ;
  LAYER M1 ;
        RECT 1.728 1.812 1.76 4.32 ;
  LAYER M3 ;
        RECT 1.728 1.832 1.76 1.864 ;
  LAYER M1 ;
        RECT 1.664 1.812 1.696 4.32 ;
  LAYER M3 ;
        RECT 1.664 4.268 1.696 4.3 ;
  LAYER M1 ;
        RECT 1.6 1.812 1.632 4.32 ;
  LAYER M3 ;
        RECT 1.6 1.832 1.632 1.864 ;
  LAYER M1 ;
        RECT 1.536 1.812 1.568 4.32 ;
  LAYER M3 ;
        RECT 1.536 4.268 1.568 4.3 ;
  LAYER M1 ;
        RECT 1.472 1.812 1.504 4.32 ;
  LAYER M3 ;
        RECT 1.472 1.832 1.504 1.864 ;
  LAYER M1 ;
        RECT 1.408 1.812 1.44 4.32 ;
  LAYER M3 ;
        RECT 1.408 4.268 1.44 4.3 ;
  LAYER M1 ;
        RECT 1.344 1.812 1.376 4.32 ;
  LAYER M3 ;
        RECT 1.344 1.832 1.376 1.864 ;
  LAYER M1 ;
        RECT 1.28 1.812 1.312 4.32 ;
  LAYER M3 ;
        RECT 1.28 4.268 1.312 4.3 ;
  LAYER M1 ;
        RECT 1.216 1.812 1.248 4.32 ;
  LAYER M3 ;
        RECT 1.216 1.832 1.248 1.864 ;
  LAYER M1 ;
        RECT 1.152 1.812 1.184 4.32 ;
  LAYER M3 ;
        RECT 1.152 4.268 1.184 4.3 ;
  LAYER M1 ;
        RECT 1.088 1.812 1.12 4.32 ;
  LAYER M3 ;
        RECT 3.456 1.896 3.488 1.928 ;
  LAYER M2 ;
        RECT 1.088 1.96 1.12 1.992 ;
  LAYER M2 ;
        RECT 3.456 2.024 3.488 2.056 ;
  LAYER M2 ;
        RECT 1.088 2.088 1.12 2.12 ;
  LAYER M2 ;
        RECT 3.456 2.152 3.488 2.184 ;
  LAYER M2 ;
        RECT 1.088 2.216 1.12 2.248 ;
  LAYER M2 ;
        RECT 3.456 2.28 3.488 2.312 ;
  LAYER M2 ;
        RECT 1.088 2.344 1.12 2.376 ;
  LAYER M2 ;
        RECT 3.456 2.408 3.488 2.44 ;
  LAYER M2 ;
        RECT 1.088 2.472 1.12 2.504 ;
  LAYER M2 ;
        RECT 3.456 2.536 3.488 2.568 ;
  LAYER M2 ;
        RECT 1.088 2.6 1.12 2.632 ;
  LAYER M2 ;
        RECT 3.456 2.664 3.488 2.696 ;
  LAYER M2 ;
        RECT 1.088 2.728 1.12 2.76 ;
  LAYER M2 ;
        RECT 3.456 2.792 3.488 2.824 ;
  LAYER M2 ;
        RECT 1.088 2.856 1.12 2.888 ;
  LAYER M2 ;
        RECT 3.456 2.92 3.488 2.952 ;
  LAYER M2 ;
        RECT 1.088 2.984 1.12 3.016 ;
  LAYER M2 ;
        RECT 3.456 3.048 3.488 3.08 ;
  LAYER M2 ;
        RECT 1.088 3.112 1.12 3.144 ;
  LAYER M2 ;
        RECT 3.456 3.176 3.488 3.208 ;
  LAYER M2 ;
        RECT 1.088 3.24 1.12 3.272 ;
  LAYER M2 ;
        RECT 3.456 3.304 3.488 3.336 ;
  LAYER M2 ;
        RECT 1.088 3.368 1.12 3.4 ;
  LAYER M2 ;
        RECT 3.456 3.432 3.488 3.464 ;
  LAYER M2 ;
        RECT 1.088 3.496 1.12 3.528 ;
  LAYER M2 ;
        RECT 3.456 3.56 3.488 3.592 ;
  LAYER M2 ;
        RECT 1.088 3.624 1.12 3.656 ;
  LAYER M2 ;
        RECT 3.456 3.688 3.488 3.72 ;
  LAYER M2 ;
        RECT 1.088 3.752 1.12 3.784 ;
  LAYER M2 ;
        RECT 3.456 3.816 3.488 3.848 ;
  LAYER M2 ;
        RECT 1.088 3.88 1.12 3.912 ;
  LAYER M2 ;
        RECT 3.456 3.944 3.488 3.976 ;
  LAYER M2 ;
        RECT 1.088 4.008 1.12 4.04 ;
  LAYER M2 ;
        RECT 3.456 4.072 3.488 4.104 ;
  LAYER M2 ;
        RECT 1.088 4.136 1.12 4.168 ;
  LAYER M2 ;
        RECT 1.04 1.764 3.536 4.368 ;
  LAYER M1 ;
        RECT 3.456 4.92 3.488 7.428 ;
  LAYER M3 ;
        RECT 3.456 7.376 3.488 7.408 ;
  LAYER M1 ;
        RECT 3.392 4.92 3.424 7.428 ;
  LAYER M3 ;
        RECT 3.392 4.94 3.424 4.972 ;
  LAYER M1 ;
        RECT 3.328 4.92 3.36 7.428 ;
  LAYER M3 ;
        RECT 3.328 7.376 3.36 7.408 ;
  LAYER M1 ;
        RECT 3.264 4.92 3.296 7.428 ;
  LAYER M3 ;
        RECT 3.264 4.94 3.296 4.972 ;
  LAYER M1 ;
        RECT 3.2 4.92 3.232 7.428 ;
  LAYER M3 ;
        RECT 3.2 7.376 3.232 7.408 ;
  LAYER M1 ;
        RECT 3.136 4.92 3.168 7.428 ;
  LAYER M3 ;
        RECT 3.136 4.94 3.168 4.972 ;
  LAYER M1 ;
        RECT 3.072 4.92 3.104 7.428 ;
  LAYER M3 ;
        RECT 3.072 7.376 3.104 7.408 ;
  LAYER M1 ;
        RECT 3.008 4.92 3.04 7.428 ;
  LAYER M3 ;
        RECT 3.008 4.94 3.04 4.972 ;
  LAYER M1 ;
        RECT 2.944 4.92 2.976 7.428 ;
  LAYER M3 ;
        RECT 2.944 7.376 2.976 7.408 ;
  LAYER M1 ;
        RECT 2.88 4.92 2.912 7.428 ;
  LAYER M3 ;
        RECT 2.88 4.94 2.912 4.972 ;
  LAYER M1 ;
        RECT 2.816 4.92 2.848 7.428 ;
  LAYER M3 ;
        RECT 2.816 7.376 2.848 7.408 ;
  LAYER M1 ;
        RECT 2.752 4.92 2.784 7.428 ;
  LAYER M3 ;
        RECT 2.752 4.94 2.784 4.972 ;
  LAYER M1 ;
        RECT 2.688 4.92 2.72 7.428 ;
  LAYER M3 ;
        RECT 2.688 7.376 2.72 7.408 ;
  LAYER M1 ;
        RECT 2.624 4.92 2.656 7.428 ;
  LAYER M3 ;
        RECT 2.624 4.94 2.656 4.972 ;
  LAYER M1 ;
        RECT 2.56 4.92 2.592 7.428 ;
  LAYER M3 ;
        RECT 2.56 7.376 2.592 7.408 ;
  LAYER M1 ;
        RECT 2.496 4.92 2.528 7.428 ;
  LAYER M3 ;
        RECT 2.496 4.94 2.528 4.972 ;
  LAYER M1 ;
        RECT 2.432 4.92 2.464 7.428 ;
  LAYER M3 ;
        RECT 2.432 7.376 2.464 7.408 ;
  LAYER M1 ;
        RECT 2.368 4.92 2.4 7.428 ;
  LAYER M3 ;
        RECT 2.368 4.94 2.4 4.972 ;
  LAYER M1 ;
        RECT 2.304 4.92 2.336 7.428 ;
  LAYER M3 ;
        RECT 2.304 7.376 2.336 7.408 ;
  LAYER M1 ;
        RECT 2.24 4.92 2.272 7.428 ;
  LAYER M3 ;
        RECT 2.24 4.94 2.272 4.972 ;
  LAYER M1 ;
        RECT 2.176 4.92 2.208 7.428 ;
  LAYER M3 ;
        RECT 2.176 7.376 2.208 7.408 ;
  LAYER M1 ;
        RECT 2.112 4.92 2.144 7.428 ;
  LAYER M3 ;
        RECT 2.112 4.94 2.144 4.972 ;
  LAYER M1 ;
        RECT 2.048 4.92 2.08 7.428 ;
  LAYER M3 ;
        RECT 2.048 7.376 2.08 7.408 ;
  LAYER M1 ;
        RECT 1.984 4.92 2.016 7.428 ;
  LAYER M3 ;
        RECT 1.984 4.94 2.016 4.972 ;
  LAYER M1 ;
        RECT 1.92 4.92 1.952 7.428 ;
  LAYER M3 ;
        RECT 1.92 7.376 1.952 7.408 ;
  LAYER M1 ;
        RECT 1.856 4.92 1.888 7.428 ;
  LAYER M3 ;
        RECT 1.856 4.94 1.888 4.972 ;
  LAYER M1 ;
        RECT 1.792 4.92 1.824 7.428 ;
  LAYER M3 ;
        RECT 1.792 7.376 1.824 7.408 ;
  LAYER M1 ;
        RECT 1.728 4.92 1.76 7.428 ;
  LAYER M3 ;
        RECT 1.728 4.94 1.76 4.972 ;
  LAYER M1 ;
        RECT 1.664 4.92 1.696 7.428 ;
  LAYER M3 ;
        RECT 1.664 7.376 1.696 7.408 ;
  LAYER M1 ;
        RECT 1.6 4.92 1.632 7.428 ;
  LAYER M3 ;
        RECT 1.6 4.94 1.632 4.972 ;
  LAYER M1 ;
        RECT 1.536 4.92 1.568 7.428 ;
  LAYER M3 ;
        RECT 1.536 7.376 1.568 7.408 ;
  LAYER M1 ;
        RECT 1.472 4.92 1.504 7.428 ;
  LAYER M3 ;
        RECT 1.472 4.94 1.504 4.972 ;
  LAYER M1 ;
        RECT 1.408 4.92 1.44 7.428 ;
  LAYER M3 ;
        RECT 1.408 7.376 1.44 7.408 ;
  LAYER M1 ;
        RECT 1.344 4.92 1.376 7.428 ;
  LAYER M3 ;
        RECT 1.344 4.94 1.376 4.972 ;
  LAYER M1 ;
        RECT 1.28 4.92 1.312 7.428 ;
  LAYER M3 ;
        RECT 1.28 7.376 1.312 7.408 ;
  LAYER M1 ;
        RECT 1.216 4.92 1.248 7.428 ;
  LAYER M3 ;
        RECT 1.216 4.94 1.248 4.972 ;
  LAYER M1 ;
        RECT 1.152 4.92 1.184 7.428 ;
  LAYER M3 ;
        RECT 1.152 7.376 1.184 7.408 ;
  LAYER M1 ;
        RECT 1.088 4.92 1.12 7.428 ;
  LAYER M3 ;
        RECT 3.456 5.004 3.488 5.036 ;
  LAYER M2 ;
        RECT 1.088 5.068 1.12 5.1 ;
  LAYER M2 ;
        RECT 3.456 5.132 3.488 5.164 ;
  LAYER M2 ;
        RECT 1.088 5.196 1.12 5.228 ;
  LAYER M2 ;
        RECT 3.456 5.26 3.488 5.292 ;
  LAYER M2 ;
        RECT 1.088 5.324 1.12 5.356 ;
  LAYER M2 ;
        RECT 3.456 5.388 3.488 5.42 ;
  LAYER M2 ;
        RECT 1.088 5.452 1.12 5.484 ;
  LAYER M2 ;
        RECT 3.456 5.516 3.488 5.548 ;
  LAYER M2 ;
        RECT 1.088 5.58 1.12 5.612 ;
  LAYER M2 ;
        RECT 3.456 5.644 3.488 5.676 ;
  LAYER M2 ;
        RECT 1.088 5.708 1.12 5.74 ;
  LAYER M2 ;
        RECT 3.456 5.772 3.488 5.804 ;
  LAYER M2 ;
        RECT 1.088 5.836 1.12 5.868 ;
  LAYER M2 ;
        RECT 3.456 5.9 3.488 5.932 ;
  LAYER M2 ;
        RECT 1.088 5.964 1.12 5.996 ;
  LAYER M2 ;
        RECT 3.456 6.028 3.488 6.06 ;
  LAYER M2 ;
        RECT 1.088 6.092 1.12 6.124 ;
  LAYER M2 ;
        RECT 3.456 6.156 3.488 6.188 ;
  LAYER M2 ;
        RECT 1.088 6.22 1.12 6.252 ;
  LAYER M2 ;
        RECT 3.456 6.284 3.488 6.316 ;
  LAYER M2 ;
        RECT 1.088 6.348 1.12 6.38 ;
  LAYER M2 ;
        RECT 3.456 6.412 3.488 6.444 ;
  LAYER M2 ;
        RECT 1.088 6.476 1.12 6.508 ;
  LAYER M2 ;
        RECT 3.456 6.54 3.488 6.572 ;
  LAYER M2 ;
        RECT 1.088 6.604 1.12 6.636 ;
  LAYER M2 ;
        RECT 3.456 6.668 3.488 6.7 ;
  LAYER M2 ;
        RECT 1.088 6.732 1.12 6.764 ;
  LAYER M2 ;
        RECT 3.456 6.796 3.488 6.828 ;
  LAYER M2 ;
        RECT 1.088 6.86 1.12 6.892 ;
  LAYER M2 ;
        RECT 3.456 6.924 3.488 6.956 ;
  LAYER M2 ;
        RECT 1.088 6.988 1.12 7.02 ;
  LAYER M2 ;
        RECT 3.456 7.052 3.488 7.084 ;
  LAYER M2 ;
        RECT 1.088 7.116 1.12 7.148 ;
  LAYER M2 ;
        RECT 3.456 7.18 3.488 7.212 ;
  LAYER M2 ;
        RECT 1.088 7.244 1.12 7.276 ;
  LAYER M2 ;
        RECT 1.04 4.872 3.536 7.476 ;
  LAYER M1 ;
        RECT 3.456 8.028 3.488 10.536 ;
  LAYER M3 ;
        RECT 3.456 10.484 3.488 10.516 ;
  LAYER M1 ;
        RECT 3.392 8.028 3.424 10.536 ;
  LAYER M3 ;
        RECT 3.392 8.048 3.424 8.08 ;
  LAYER M1 ;
        RECT 3.328 8.028 3.36 10.536 ;
  LAYER M3 ;
        RECT 3.328 10.484 3.36 10.516 ;
  LAYER M1 ;
        RECT 3.264 8.028 3.296 10.536 ;
  LAYER M3 ;
        RECT 3.264 8.048 3.296 8.08 ;
  LAYER M1 ;
        RECT 3.2 8.028 3.232 10.536 ;
  LAYER M3 ;
        RECT 3.2 10.484 3.232 10.516 ;
  LAYER M1 ;
        RECT 3.136 8.028 3.168 10.536 ;
  LAYER M3 ;
        RECT 3.136 8.048 3.168 8.08 ;
  LAYER M1 ;
        RECT 3.072 8.028 3.104 10.536 ;
  LAYER M3 ;
        RECT 3.072 10.484 3.104 10.516 ;
  LAYER M1 ;
        RECT 3.008 8.028 3.04 10.536 ;
  LAYER M3 ;
        RECT 3.008 8.048 3.04 8.08 ;
  LAYER M1 ;
        RECT 2.944 8.028 2.976 10.536 ;
  LAYER M3 ;
        RECT 2.944 10.484 2.976 10.516 ;
  LAYER M1 ;
        RECT 2.88 8.028 2.912 10.536 ;
  LAYER M3 ;
        RECT 2.88 8.048 2.912 8.08 ;
  LAYER M1 ;
        RECT 2.816 8.028 2.848 10.536 ;
  LAYER M3 ;
        RECT 2.816 10.484 2.848 10.516 ;
  LAYER M1 ;
        RECT 2.752 8.028 2.784 10.536 ;
  LAYER M3 ;
        RECT 2.752 8.048 2.784 8.08 ;
  LAYER M1 ;
        RECT 2.688 8.028 2.72 10.536 ;
  LAYER M3 ;
        RECT 2.688 10.484 2.72 10.516 ;
  LAYER M1 ;
        RECT 2.624 8.028 2.656 10.536 ;
  LAYER M3 ;
        RECT 2.624 8.048 2.656 8.08 ;
  LAYER M1 ;
        RECT 2.56 8.028 2.592 10.536 ;
  LAYER M3 ;
        RECT 2.56 10.484 2.592 10.516 ;
  LAYER M1 ;
        RECT 2.496 8.028 2.528 10.536 ;
  LAYER M3 ;
        RECT 2.496 8.048 2.528 8.08 ;
  LAYER M1 ;
        RECT 2.432 8.028 2.464 10.536 ;
  LAYER M3 ;
        RECT 2.432 10.484 2.464 10.516 ;
  LAYER M1 ;
        RECT 2.368 8.028 2.4 10.536 ;
  LAYER M3 ;
        RECT 2.368 8.048 2.4 8.08 ;
  LAYER M1 ;
        RECT 2.304 8.028 2.336 10.536 ;
  LAYER M3 ;
        RECT 2.304 10.484 2.336 10.516 ;
  LAYER M1 ;
        RECT 2.24 8.028 2.272 10.536 ;
  LAYER M3 ;
        RECT 2.24 8.048 2.272 8.08 ;
  LAYER M1 ;
        RECT 2.176 8.028 2.208 10.536 ;
  LAYER M3 ;
        RECT 2.176 10.484 2.208 10.516 ;
  LAYER M1 ;
        RECT 2.112 8.028 2.144 10.536 ;
  LAYER M3 ;
        RECT 2.112 8.048 2.144 8.08 ;
  LAYER M1 ;
        RECT 2.048 8.028 2.08 10.536 ;
  LAYER M3 ;
        RECT 2.048 10.484 2.08 10.516 ;
  LAYER M1 ;
        RECT 1.984 8.028 2.016 10.536 ;
  LAYER M3 ;
        RECT 1.984 8.048 2.016 8.08 ;
  LAYER M1 ;
        RECT 1.92 8.028 1.952 10.536 ;
  LAYER M3 ;
        RECT 1.92 10.484 1.952 10.516 ;
  LAYER M1 ;
        RECT 1.856 8.028 1.888 10.536 ;
  LAYER M3 ;
        RECT 1.856 8.048 1.888 8.08 ;
  LAYER M1 ;
        RECT 1.792 8.028 1.824 10.536 ;
  LAYER M3 ;
        RECT 1.792 10.484 1.824 10.516 ;
  LAYER M1 ;
        RECT 1.728 8.028 1.76 10.536 ;
  LAYER M3 ;
        RECT 1.728 8.048 1.76 8.08 ;
  LAYER M1 ;
        RECT 1.664 8.028 1.696 10.536 ;
  LAYER M3 ;
        RECT 1.664 10.484 1.696 10.516 ;
  LAYER M1 ;
        RECT 1.6 8.028 1.632 10.536 ;
  LAYER M3 ;
        RECT 1.6 8.048 1.632 8.08 ;
  LAYER M1 ;
        RECT 1.536 8.028 1.568 10.536 ;
  LAYER M3 ;
        RECT 1.536 10.484 1.568 10.516 ;
  LAYER M1 ;
        RECT 1.472 8.028 1.504 10.536 ;
  LAYER M3 ;
        RECT 1.472 8.048 1.504 8.08 ;
  LAYER M1 ;
        RECT 1.408 8.028 1.44 10.536 ;
  LAYER M3 ;
        RECT 1.408 10.484 1.44 10.516 ;
  LAYER M1 ;
        RECT 1.344 8.028 1.376 10.536 ;
  LAYER M3 ;
        RECT 1.344 8.048 1.376 8.08 ;
  LAYER M1 ;
        RECT 1.28 8.028 1.312 10.536 ;
  LAYER M3 ;
        RECT 1.28 10.484 1.312 10.516 ;
  LAYER M1 ;
        RECT 1.216 8.028 1.248 10.536 ;
  LAYER M3 ;
        RECT 1.216 8.048 1.248 8.08 ;
  LAYER M1 ;
        RECT 1.152 8.028 1.184 10.536 ;
  LAYER M3 ;
        RECT 1.152 10.484 1.184 10.516 ;
  LAYER M1 ;
        RECT 1.088 8.028 1.12 10.536 ;
  LAYER M3 ;
        RECT 3.456 8.112 3.488 8.144 ;
  LAYER M2 ;
        RECT 1.088 8.176 1.12 8.208 ;
  LAYER M2 ;
        RECT 3.456 8.24 3.488 8.272 ;
  LAYER M2 ;
        RECT 1.088 8.304 1.12 8.336 ;
  LAYER M2 ;
        RECT 3.456 8.368 3.488 8.4 ;
  LAYER M2 ;
        RECT 1.088 8.432 1.12 8.464 ;
  LAYER M2 ;
        RECT 3.456 8.496 3.488 8.528 ;
  LAYER M2 ;
        RECT 1.088 8.56 1.12 8.592 ;
  LAYER M2 ;
        RECT 3.456 8.624 3.488 8.656 ;
  LAYER M2 ;
        RECT 1.088 8.688 1.12 8.72 ;
  LAYER M2 ;
        RECT 3.456 8.752 3.488 8.784 ;
  LAYER M2 ;
        RECT 1.088 8.816 1.12 8.848 ;
  LAYER M2 ;
        RECT 3.456 8.88 3.488 8.912 ;
  LAYER M2 ;
        RECT 1.088 8.944 1.12 8.976 ;
  LAYER M2 ;
        RECT 3.456 9.008 3.488 9.04 ;
  LAYER M2 ;
        RECT 1.088 9.072 1.12 9.104 ;
  LAYER M2 ;
        RECT 3.456 9.136 3.488 9.168 ;
  LAYER M2 ;
        RECT 1.088 9.2 1.12 9.232 ;
  LAYER M2 ;
        RECT 3.456 9.264 3.488 9.296 ;
  LAYER M2 ;
        RECT 1.088 9.328 1.12 9.36 ;
  LAYER M2 ;
        RECT 3.456 9.392 3.488 9.424 ;
  LAYER M2 ;
        RECT 1.088 9.456 1.12 9.488 ;
  LAYER M2 ;
        RECT 3.456 9.52 3.488 9.552 ;
  LAYER M2 ;
        RECT 1.088 9.584 1.12 9.616 ;
  LAYER M2 ;
        RECT 3.456 9.648 3.488 9.68 ;
  LAYER M2 ;
        RECT 1.088 9.712 1.12 9.744 ;
  LAYER M2 ;
        RECT 3.456 9.776 3.488 9.808 ;
  LAYER M2 ;
        RECT 1.088 9.84 1.12 9.872 ;
  LAYER M2 ;
        RECT 3.456 9.904 3.488 9.936 ;
  LAYER M2 ;
        RECT 1.088 9.968 1.12 10 ;
  LAYER M2 ;
        RECT 3.456 10.032 3.488 10.064 ;
  LAYER M2 ;
        RECT 1.088 10.096 1.12 10.128 ;
  LAYER M2 ;
        RECT 3.456 10.16 3.488 10.192 ;
  LAYER M2 ;
        RECT 1.088 10.224 1.12 10.256 ;
  LAYER M2 ;
        RECT 3.456 10.288 3.488 10.32 ;
  LAYER M2 ;
        RECT 1.088 10.352 1.12 10.384 ;
  LAYER M2 ;
        RECT 1.04 7.98 3.536 10.584 ;
  LAYER M1 ;
        RECT 3.456 11.136 3.488 13.644 ;
  LAYER M3 ;
        RECT 3.456 13.592 3.488 13.624 ;
  LAYER M1 ;
        RECT 3.392 11.136 3.424 13.644 ;
  LAYER M3 ;
        RECT 3.392 11.156 3.424 11.188 ;
  LAYER M1 ;
        RECT 3.328 11.136 3.36 13.644 ;
  LAYER M3 ;
        RECT 3.328 13.592 3.36 13.624 ;
  LAYER M1 ;
        RECT 3.264 11.136 3.296 13.644 ;
  LAYER M3 ;
        RECT 3.264 11.156 3.296 11.188 ;
  LAYER M1 ;
        RECT 3.2 11.136 3.232 13.644 ;
  LAYER M3 ;
        RECT 3.2 13.592 3.232 13.624 ;
  LAYER M1 ;
        RECT 3.136 11.136 3.168 13.644 ;
  LAYER M3 ;
        RECT 3.136 11.156 3.168 11.188 ;
  LAYER M1 ;
        RECT 3.072 11.136 3.104 13.644 ;
  LAYER M3 ;
        RECT 3.072 13.592 3.104 13.624 ;
  LAYER M1 ;
        RECT 3.008 11.136 3.04 13.644 ;
  LAYER M3 ;
        RECT 3.008 11.156 3.04 11.188 ;
  LAYER M1 ;
        RECT 2.944 11.136 2.976 13.644 ;
  LAYER M3 ;
        RECT 2.944 13.592 2.976 13.624 ;
  LAYER M1 ;
        RECT 2.88 11.136 2.912 13.644 ;
  LAYER M3 ;
        RECT 2.88 11.156 2.912 11.188 ;
  LAYER M1 ;
        RECT 2.816 11.136 2.848 13.644 ;
  LAYER M3 ;
        RECT 2.816 13.592 2.848 13.624 ;
  LAYER M1 ;
        RECT 2.752 11.136 2.784 13.644 ;
  LAYER M3 ;
        RECT 2.752 11.156 2.784 11.188 ;
  LAYER M1 ;
        RECT 2.688 11.136 2.72 13.644 ;
  LAYER M3 ;
        RECT 2.688 13.592 2.72 13.624 ;
  LAYER M1 ;
        RECT 2.624 11.136 2.656 13.644 ;
  LAYER M3 ;
        RECT 2.624 11.156 2.656 11.188 ;
  LAYER M1 ;
        RECT 2.56 11.136 2.592 13.644 ;
  LAYER M3 ;
        RECT 2.56 13.592 2.592 13.624 ;
  LAYER M1 ;
        RECT 2.496 11.136 2.528 13.644 ;
  LAYER M3 ;
        RECT 2.496 11.156 2.528 11.188 ;
  LAYER M1 ;
        RECT 2.432 11.136 2.464 13.644 ;
  LAYER M3 ;
        RECT 2.432 13.592 2.464 13.624 ;
  LAYER M1 ;
        RECT 2.368 11.136 2.4 13.644 ;
  LAYER M3 ;
        RECT 2.368 11.156 2.4 11.188 ;
  LAYER M1 ;
        RECT 2.304 11.136 2.336 13.644 ;
  LAYER M3 ;
        RECT 2.304 13.592 2.336 13.624 ;
  LAYER M1 ;
        RECT 2.24 11.136 2.272 13.644 ;
  LAYER M3 ;
        RECT 2.24 11.156 2.272 11.188 ;
  LAYER M1 ;
        RECT 2.176 11.136 2.208 13.644 ;
  LAYER M3 ;
        RECT 2.176 13.592 2.208 13.624 ;
  LAYER M1 ;
        RECT 2.112 11.136 2.144 13.644 ;
  LAYER M3 ;
        RECT 2.112 11.156 2.144 11.188 ;
  LAYER M1 ;
        RECT 2.048 11.136 2.08 13.644 ;
  LAYER M3 ;
        RECT 2.048 13.592 2.08 13.624 ;
  LAYER M1 ;
        RECT 1.984 11.136 2.016 13.644 ;
  LAYER M3 ;
        RECT 1.984 11.156 2.016 11.188 ;
  LAYER M1 ;
        RECT 1.92 11.136 1.952 13.644 ;
  LAYER M3 ;
        RECT 1.92 13.592 1.952 13.624 ;
  LAYER M1 ;
        RECT 1.856 11.136 1.888 13.644 ;
  LAYER M3 ;
        RECT 1.856 11.156 1.888 11.188 ;
  LAYER M1 ;
        RECT 1.792 11.136 1.824 13.644 ;
  LAYER M3 ;
        RECT 1.792 13.592 1.824 13.624 ;
  LAYER M1 ;
        RECT 1.728 11.136 1.76 13.644 ;
  LAYER M3 ;
        RECT 1.728 11.156 1.76 11.188 ;
  LAYER M1 ;
        RECT 1.664 11.136 1.696 13.644 ;
  LAYER M3 ;
        RECT 1.664 13.592 1.696 13.624 ;
  LAYER M1 ;
        RECT 1.6 11.136 1.632 13.644 ;
  LAYER M3 ;
        RECT 1.6 11.156 1.632 11.188 ;
  LAYER M1 ;
        RECT 1.536 11.136 1.568 13.644 ;
  LAYER M3 ;
        RECT 1.536 13.592 1.568 13.624 ;
  LAYER M1 ;
        RECT 1.472 11.136 1.504 13.644 ;
  LAYER M3 ;
        RECT 1.472 11.156 1.504 11.188 ;
  LAYER M1 ;
        RECT 1.408 11.136 1.44 13.644 ;
  LAYER M3 ;
        RECT 1.408 13.592 1.44 13.624 ;
  LAYER M1 ;
        RECT 1.344 11.136 1.376 13.644 ;
  LAYER M3 ;
        RECT 1.344 11.156 1.376 11.188 ;
  LAYER M1 ;
        RECT 1.28 11.136 1.312 13.644 ;
  LAYER M3 ;
        RECT 1.28 13.592 1.312 13.624 ;
  LAYER M1 ;
        RECT 1.216 11.136 1.248 13.644 ;
  LAYER M3 ;
        RECT 1.216 11.156 1.248 11.188 ;
  LAYER M1 ;
        RECT 1.152 11.136 1.184 13.644 ;
  LAYER M3 ;
        RECT 1.152 13.592 1.184 13.624 ;
  LAYER M1 ;
        RECT 1.088 11.136 1.12 13.644 ;
  LAYER M3 ;
        RECT 3.456 11.22 3.488 11.252 ;
  LAYER M2 ;
        RECT 1.088 11.284 1.12 11.316 ;
  LAYER M2 ;
        RECT 3.456 11.348 3.488 11.38 ;
  LAYER M2 ;
        RECT 1.088 11.412 1.12 11.444 ;
  LAYER M2 ;
        RECT 3.456 11.476 3.488 11.508 ;
  LAYER M2 ;
        RECT 1.088 11.54 1.12 11.572 ;
  LAYER M2 ;
        RECT 3.456 11.604 3.488 11.636 ;
  LAYER M2 ;
        RECT 1.088 11.668 1.12 11.7 ;
  LAYER M2 ;
        RECT 3.456 11.732 3.488 11.764 ;
  LAYER M2 ;
        RECT 1.088 11.796 1.12 11.828 ;
  LAYER M2 ;
        RECT 3.456 11.86 3.488 11.892 ;
  LAYER M2 ;
        RECT 1.088 11.924 1.12 11.956 ;
  LAYER M2 ;
        RECT 3.456 11.988 3.488 12.02 ;
  LAYER M2 ;
        RECT 1.088 12.052 1.12 12.084 ;
  LAYER M2 ;
        RECT 3.456 12.116 3.488 12.148 ;
  LAYER M2 ;
        RECT 1.088 12.18 1.12 12.212 ;
  LAYER M2 ;
        RECT 3.456 12.244 3.488 12.276 ;
  LAYER M2 ;
        RECT 1.088 12.308 1.12 12.34 ;
  LAYER M2 ;
        RECT 3.456 12.372 3.488 12.404 ;
  LAYER M2 ;
        RECT 1.088 12.436 1.12 12.468 ;
  LAYER M2 ;
        RECT 3.456 12.5 3.488 12.532 ;
  LAYER M2 ;
        RECT 1.088 12.564 1.12 12.596 ;
  LAYER M2 ;
        RECT 3.456 12.628 3.488 12.66 ;
  LAYER M2 ;
        RECT 1.088 12.692 1.12 12.724 ;
  LAYER M2 ;
        RECT 3.456 12.756 3.488 12.788 ;
  LAYER M2 ;
        RECT 1.088 12.82 1.12 12.852 ;
  LAYER M2 ;
        RECT 3.456 12.884 3.488 12.916 ;
  LAYER M2 ;
        RECT 1.088 12.948 1.12 12.98 ;
  LAYER M2 ;
        RECT 3.456 13.012 3.488 13.044 ;
  LAYER M2 ;
        RECT 1.088 13.076 1.12 13.108 ;
  LAYER M2 ;
        RECT 3.456 13.14 3.488 13.172 ;
  LAYER M2 ;
        RECT 1.088 13.204 1.12 13.236 ;
  LAYER M2 ;
        RECT 3.456 13.268 3.488 13.3 ;
  LAYER M2 ;
        RECT 1.088 13.332 1.12 13.364 ;
  LAYER M2 ;
        RECT 3.456 13.396 3.488 13.428 ;
  LAYER M2 ;
        RECT 1.088 13.46 1.12 13.492 ;
  LAYER M2 ;
        RECT 1.04 11.088 3.536 13.692 ;
  LAYER M1 ;
        RECT 10.704 0.132 10.736 0.792 ;
  LAYER M1 ;
        RECT 10.784 0.132 10.816 0.792 ;
  LAYER M1 ;
        RECT 10.624 0.572 10.656 0.604 ;
  LAYER M1 ;
        RECT 0.384 0.132 0.416 0.792 ;
  LAYER M1 ;
        RECT 0.304 0.132 0.336 0.792 ;
  LAYER M1 ;
        RECT 0.464 0.572 0.496 0.604 ;
  LAYER M1 ;
        RECT 9.344 0.216 9.376 0.876 ;
  LAYER M1 ;
        RECT 9.984 0.216 10.016 0.876 ;
  LAYER M1 ;
        RECT 9.264 0.216 9.296 0.876 ;
  LAYER M1 ;
        RECT 9.904 0.216 9.936 0.876 ;
  LAYER M1 ;
        RECT 9.424 0.216 9.456 0.876 ;
  LAYER M1 ;
        RECT 10.064 0.404 10.096 0.436 ;
  LAYER M1 ;
        RECT 7.984 0.216 8.016 0.876 ;
  LAYER M1 ;
        RECT 8.624 0.216 8.656 0.876 ;
  LAYER M1 ;
        RECT 7.904 0.216 7.936 0.876 ;
  LAYER M1 ;
        RECT 8.544 0.216 8.576 0.876 ;
  LAYER M1 ;
        RECT 8.064 0.216 8.096 0.876 ;
  LAYER M1 ;
        RECT 8.704 0.404 8.736 0.436 ;
  LAYER M1 ;
        RECT 9.488 24.156 9.52 24.228 ;
  LAYER M2 ;
        RECT 9.468 24.176 9.54 24.208 ;
  LAYER M2 ;
        RECT 6.752 24.176 9.504 24.208 ;
  LAYER M1 ;
        RECT 6.736 24.156 6.768 24.228 ;
  LAYER M2 ;
        RECT 6.716 24.176 6.788 24.208 ;
  LAYER M1 ;
        RECT 6.512 21.048 6.544 21.12 ;
  LAYER M2 ;
        RECT 6.492 21.068 6.564 21.1 ;
  LAYER M1 ;
        RECT 6.512 21.084 6.544 21.252 ;
  LAYER M1 ;
        RECT 6.512 21.216 6.544 21.288 ;
  LAYER M2 ;
        RECT 6.492 21.236 6.564 21.268 ;
  LAYER M2 ;
        RECT 6.528 21.236 6.752 21.268 ;
  LAYER M1 ;
        RECT 6.736 21.216 6.768 21.288 ;
  LAYER M2 ;
        RECT 6.716 21.236 6.788 21.268 ;
  LAYER M1 ;
        RECT 6.736 30.96 6.768 31.032 ;
  LAYER M2 ;
        RECT 6.716 30.98 6.788 31.012 ;
  LAYER M1 ;
        RECT 6.736 30.744 6.768 30.996 ;
  LAYER M1 ;
        RECT 6.736 21.252 6.768 30.744 ;
  LAYER M1 ;
        RECT 12.464 27.264 12.496 27.336 ;
  LAYER M2 ;
        RECT 12.444 27.284 12.516 27.316 ;
  LAYER M2 ;
        RECT 9.728 27.284 12.48 27.316 ;
  LAYER M1 ;
        RECT 9.712 27.264 9.744 27.336 ;
  LAYER M2 ;
        RECT 9.692 27.284 9.764 27.316 ;
  LAYER M1 ;
        RECT 9.712 30.96 9.744 31.032 ;
  LAYER M2 ;
        RECT 9.692 30.98 9.764 31.012 ;
  LAYER M1 ;
        RECT 9.712 30.744 9.744 30.996 ;
  LAYER M1 ;
        RECT 9.712 27.3 9.744 30.744 ;
  LAYER M2 ;
        RECT 6.752 30.98 9.728 31.012 ;
  LAYER M1 ;
        RECT 6.512 24.156 6.544 24.228 ;
  LAYER M2 ;
        RECT 6.492 24.176 6.564 24.208 ;
  LAYER M2 ;
        RECT 3.776 24.176 6.528 24.208 ;
  LAYER M1 ;
        RECT 3.76 24.156 3.792 24.228 ;
  LAYER M2 ;
        RECT 3.74 24.176 3.812 24.208 ;
  LAYER M1 ;
        RECT 6.512 27.264 6.544 27.336 ;
  LAYER M2 ;
        RECT 6.492 27.284 6.564 27.316 ;
  LAYER M2 ;
        RECT 3.776 27.284 6.528 27.316 ;
  LAYER M1 ;
        RECT 3.76 27.264 3.792 27.336 ;
  LAYER M2 ;
        RECT 3.74 27.284 3.812 27.316 ;
  LAYER M1 ;
        RECT 3.76 31.128 3.792 31.2 ;
  LAYER M2 ;
        RECT 3.74 31.148 3.812 31.18 ;
  LAYER M1 ;
        RECT 3.76 30.744 3.792 31.164 ;
  LAYER M1 ;
        RECT 3.76 24.192 3.792 30.744 ;
  LAYER M1 ;
        RECT 12.464 24.156 12.496 24.228 ;
  LAYER M2 ;
        RECT 12.444 24.176 12.516 24.208 ;
  LAYER M1 ;
        RECT 12.464 24.192 12.496 24.36 ;
  LAYER M1 ;
        RECT 12.464 24.324 12.496 24.396 ;
  LAYER M2 ;
        RECT 12.444 24.344 12.516 24.376 ;
  LAYER M2 ;
        RECT 12.48 24.344 12.704 24.376 ;
  LAYER M1 ;
        RECT 12.688 24.324 12.72 24.396 ;
  LAYER M2 ;
        RECT 12.668 24.344 12.74 24.376 ;
  LAYER M1 ;
        RECT 12.464 21.048 12.496 21.12 ;
  LAYER M2 ;
        RECT 12.444 21.068 12.516 21.1 ;
  LAYER M1 ;
        RECT 12.464 21.084 12.496 21.252 ;
  LAYER M1 ;
        RECT 12.464 21.216 12.496 21.288 ;
  LAYER M2 ;
        RECT 12.444 21.236 12.516 21.268 ;
  LAYER M2 ;
        RECT 12.48 21.236 12.704 21.268 ;
  LAYER M1 ;
        RECT 12.688 21.216 12.72 21.288 ;
  LAYER M2 ;
        RECT 12.668 21.236 12.74 21.268 ;
  LAYER M1 ;
        RECT 12.688 31.128 12.72 31.2 ;
  LAYER M2 ;
        RECT 12.668 31.148 12.74 31.18 ;
  LAYER M1 ;
        RECT 12.688 30.744 12.72 31.164 ;
  LAYER M1 ;
        RECT 12.688 21.252 12.72 30.744 ;
  LAYER M2 ;
        RECT 3.776 31.148 12.704 31.18 ;
  LAYER M1 ;
        RECT 9.488 27.264 9.52 27.336 ;
  LAYER M2 ;
        RECT 9.468 27.284 9.54 27.316 ;
  LAYER M2 ;
        RECT 6.528 27.284 9.504 27.316 ;
  LAYER M1 ;
        RECT 6.512 27.264 6.544 27.336 ;
  LAYER M2 ;
        RECT 6.492 27.284 6.564 27.316 ;
  LAYER M1 ;
        RECT 9.488 21.048 9.52 21.12 ;
  LAYER M2 ;
        RECT 9.468 21.068 9.54 21.1 ;
  LAYER M2 ;
        RECT 9.504 21.068 12.48 21.1 ;
  LAYER M1 ;
        RECT 12.464 21.048 12.496 21.12 ;
  LAYER M2 ;
        RECT 12.444 21.068 12.516 21.1 ;
  LAYER M1 ;
        RECT 3.536 30.372 3.568 30.444 ;
  LAYER M2 ;
        RECT 3.516 30.392 3.588 30.424 ;
  LAYER M2 ;
        RECT 0.8 30.392 3.552 30.424 ;
  LAYER M1 ;
        RECT 0.784 30.372 0.816 30.444 ;
  LAYER M2 ;
        RECT 0.764 30.392 0.836 30.424 ;
  LAYER M1 ;
        RECT 3.536 27.264 3.568 27.336 ;
  LAYER M2 ;
        RECT 3.516 27.284 3.588 27.316 ;
  LAYER M2 ;
        RECT 0.8 27.284 3.552 27.316 ;
  LAYER M1 ;
        RECT 0.784 27.264 0.816 27.336 ;
  LAYER M2 ;
        RECT 0.764 27.284 0.836 27.316 ;
  LAYER M1 ;
        RECT 3.536 24.156 3.568 24.228 ;
  LAYER M2 ;
        RECT 3.516 24.176 3.588 24.208 ;
  LAYER M2 ;
        RECT 0.8 24.176 3.552 24.208 ;
  LAYER M1 ;
        RECT 0.784 24.156 0.816 24.228 ;
  LAYER M2 ;
        RECT 0.764 24.176 0.836 24.208 ;
  LAYER M1 ;
        RECT 3.536 21.048 3.568 21.12 ;
  LAYER M2 ;
        RECT 3.516 21.068 3.588 21.1 ;
  LAYER M2 ;
        RECT 0.8 21.068 3.552 21.1 ;
  LAYER M1 ;
        RECT 0.784 21.048 0.816 21.12 ;
  LAYER M2 ;
        RECT 0.764 21.068 0.836 21.1 ;
  LAYER M1 ;
        RECT 3.536 17.94 3.568 18.012 ;
  LAYER M2 ;
        RECT 3.516 17.96 3.588 17.992 ;
  LAYER M2 ;
        RECT 0.8 17.96 3.552 17.992 ;
  LAYER M1 ;
        RECT 0.784 17.94 0.816 18.012 ;
  LAYER M2 ;
        RECT 0.764 17.96 0.836 17.992 ;
  LAYER M1 ;
        RECT 0.784 31.296 0.816 31.368 ;
  LAYER M2 ;
        RECT 0.764 31.316 0.836 31.348 ;
  LAYER M1 ;
        RECT 0.784 30.744 0.816 31.332 ;
  LAYER M1 ;
        RECT 0.784 17.976 0.816 30.744 ;
  LAYER M1 ;
        RECT 15.44 30.372 15.472 30.444 ;
  LAYER M2 ;
        RECT 15.42 30.392 15.492 30.424 ;
  LAYER M1 ;
        RECT 15.44 30.408 15.472 30.576 ;
  LAYER M1 ;
        RECT 15.44 30.54 15.472 30.612 ;
  LAYER M2 ;
        RECT 15.42 30.56 15.492 30.592 ;
  LAYER M2 ;
        RECT 15.456 30.56 15.68 30.592 ;
  LAYER M1 ;
        RECT 15.664 30.54 15.696 30.612 ;
  LAYER M2 ;
        RECT 15.644 30.56 15.716 30.592 ;
  LAYER M1 ;
        RECT 15.44 27.264 15.472 27.336 ;
  LAYER M2 ;
        RECT 15.42 27.284 15.492 27.316 ;
  LAYER M1 ;
        RECT 15.44 27.3 15.472 27.468 ;
  LAYER M1 ;
        RECT 15.44 27.432 15.472 27.504 ;
  LAYER M2 ;
        RECT 15.42 27.452 15.492 27.484 ;
  LAYER M2 ;
        RECT 15.456 27.452 15.68 27.484 ;
  LAYER M1 ;
        RECT 15.664 27.432 15.696 27.504 ;
  LAYER M2 ;
        RECT 15.644 27.452 15.716 27.484 ;
  LAYER M1 ;
        RECT 15.44 24.156 15.472 24.228 ;
  LAYER M2 ;
        RECT 15.42 24.176 15.492 24.208 ;
  LAYER M1 ;
        RECT 15.44 24.192 15.472 24.36 ;
  LAYER M1 ;
        RECT 15.44 24.324 15.472 24.396 ;
  LAYER M2 ;
        RECT 15.42 24.344 15.492 24.376 ;
  LAYER M2 ;
        RECT 15.456 24.344 15.68 24.376 ;
  LAYER M1 ;
        RECT 15.664 24.324 15.696 24.396 ;
  LAYER M2 ;
        RECT 15.644 24.344 15.716 24.376 ;
  LAYER M1 ;
        RECT 15.44 21.048 15.472 21.12 ;
  LAYER M2 ;
        RECT 15.42 21.068 15.492 21.1 ;
  LAYER M1 ;
        RECT 15.44 21.084 15.472 21.252 ;
  LAYER M1 ;
        RECT 15.44 21.216 15.472 21.288 ;
  LAYER M2 ;
        RECT 15.42 21.236 15.492 21.268 ;
  LAYER M2 ;
        RECT 15.456 21.236 15.68 21.268 ;
  LAYER M1 ;
        RECT 15.664 21.216 15.696 21.288 ;
  LAYER M2 ;
        RECT 15.644 21.236 15.716 21.268 ;
  LAYER M1 ;
        RECT 15.44 17.94 15.472 18.012 ;
  LAYER M2 ;
        RECT 15.42 17.96 15.492 17.992 ;
  LAYER M1 ;
        RECT 15.44 17.976 15.472 18.144 ;
  LAYER M1 ;
        RECT 15.44 18.108 15.472 18.18 ;
  LAYER M2 ;
        RECT 15.42 18.128 15.492 18.16 ;
  LAYER M2 ;
        RECT 15.456 18.128 15.68 18.16 ;
  LAYER M1 ;
        RECT 15.664 18.108 15.696 18.18 ;
  LAYER M2 ;
        RECT 15.644 18.128 15.716 18.16 ;
  LAYER M1 ;
        RECT 15.664 31.296 15.696 31.368 ;
  LAYER M2 ;
        RECT 15.644 31.316 15.716 31.348 ;
  LAYER M1 ;
        RECT 15.664 30.744 15.696 31.332 ;
  LAYER M1 ;
        RECT 15.664 18.144 15.696 30.744 ;
  LAYER M2 ;
        RECT 0.8 31.316 15.68 31.348 ;
  LAYER M1 ;
        RECT 6.512 30.372 6.544 30.444 ;
  LAYER M2 ;
        RECT 6.492 30.392 6.564 30.424 ;
  LAYER M2 ;
        RECT 3.552 30.392 6.528 30.424 ;
  LAYER M1 ;
        RECT 3.536 30.372 3.568 30.444 ;
  LAYER M2 ;
        RECT 3.516 30.392 3.588 30.424 ;
  LAYER M1 ;
        RECT 6.512 17.94 6.544 18.012 ;
  LAYER M2 ;
        RECT 6.492 17.96 6.564 17.992 ;
  LAYER M2 ;
        RECT 3.552 17.96 6.528 17.992 ;
  LAYER M1 ;
        RECT 3.536 17.94 3.568 18.012 ;
  LAYER M2 ;
        RECT 3.516 17.96 3.588 17.992 ;
  LAYER M1 ;
        RECT 9.488 17.94 9.52 18.012 ;
  LAYER M2 ;
        RECT 9.468 17.96 9.54 17.992 ;
  LAYER M2 ;
        RECT 6.528 17.96 9.504 17.992 ;
  LAYER M1 ;
        RECT 6.512 17.94 6.544 18.012 ;
  LAYER M2 ;
        RECT 6.492 17.96 6.564 17.992 ;
  LAYER M1 ;
        RECT 12.464 17.94 12.496 18.012 ;
  LAYER M2 ;
        RECT 12.444 17.96 12.516 17.992 ;
  LAYER M2 ;
        RECT 9.504 17.96 12.48 17.992 ;
  LAYER M1 ;
        RECT 9.488 17.94 9.52 18.012 ;
  LAYER M2 ;
        RECT 9.468 17.96 9.54 17.992 ;
  LAYER M1 ;
        RECT 12.464 30.372 12.496 30.444 ;
  LAYER M2 ;
        RECT 12.444 30.392 12.516 30.424 ;
  LAYER M2 ;
        RECT 12.48 30.392 15.456 30.424 ;
  LAYER M1 ;
        RECT 15.44 30.372 15.472 30.444 ;
  LAYER M2 ;
        RECT 15.42 30.392 15.492 30.424 ;
  LAYER M1 ;
        RECT 9.488 30.372 9.52 30.444 ;
  LAYER M2 ;
        RECT 9.468 30.392 9.54 30.424 ;
  LAYER M2 ;
        RECT 9.504 30.392 12.48 30.424 ;
  LAYER M1 ;
        RECT 12.464 30.372 12.496 30.444 ;
  LAYER M2 ;
        RECT 12.444 30.392 12.516 30.424 ;
  LAYER M1 ;
        RECT 7.12 21.72 7.152 21.792 ;
  LAYER M2 ;
        RECT 7.1 21.74 7.172 21.772 ;
  LAYER M2 ;
        RECT 6.912 21.74 7.136 21.772 ;
  LAYER M1 ;
        RECT 6.896 21.72 6.928 21.792 ;
  LAYER M2 ;
        RECT 6.876 21.74 6.948 21.772 ;
  LAYER M1 ;
        RECT 4.144 18.612 4.176 18.684 ;
  LAYER M2 ;
        RECT 4.124 18.632 4.196 18.664 ;
  LAYER M1 ;
        RECT 4.144 18.48 4.176 18.648 ;
  LAYER M1 ;
        RECT 4.144 18.444 4.176 18.516 ;
  LAYER M2 ;
        RECT 4.124 18.464 4.196 18.496 ;
  LAYER M2 ;
        RECT 4.16 18.464 6.912 18.496 ;
  LAYER M1 ;
        RECT 6.896 18.444 6.928 18.516 ;
  LAYER M2 ;
        RECT 6.876 18.464 6.948 18.496 ;
  LAYER M1 ;
        RECT 6.896 14.916 6.928 14.988 ;
  LAYER M2 ;
        RECT 6.876 14.936 6.948 14.968 ;
  LAYER M1 ;
        RECT 6.896 14.952 6.928 15.204 ;
  LAYER M1 ;
        RECT 6.896 15.204 6.928 21.756 ;
  LAYER M1 ;
        RECT 10.096 24.828 10.128 24.9 ;
  LAYER M2 ;
        RECT 10.076 24.848 10.148 24.88 ;
  LAYER M2 ;
        RECT 9.888 24.848 10.112 24.88 ;
  LAYER M1 ;
        RECT 9.872 24.828 9.904 24.9 ;
  LAYER M2 ;
        RECT 9.852 24.848 9.924 24.88 ;
  LAYER M1 ;
        RECT 9.872 14.916 9.904 14.988 ;
  LAYER M2 ;
        RECT 9.852 14.936 9.924 14.968 ;
  LAYER M1 ;
        RECT 9.872 14.952 9.904 15.204 ;
  LAYER M1 ;
        RECT 9.872 15.204 9.904 24.864 ;
  LAYER M2 ;
        RECT 6.912 14.936 9.888 14.968 ;
  LAYER M1 ;
        RECT 4.144 21.72 4.176 21.792 ;
  LAYER M2 ;
        RECT 4.124 21.74 4.196 21.772 ;
  LAYER M2 ;
        RECT 3.936 21.74 4.16 21.772 ;
  LAYER M1 ;
        RECT 3.92 21.72 3.952 21.792 ;
  LAYER M2 ;
        RECT 3.9 21.74 3.972 21.772 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 24.9 ;
  LAYER M2 ;
        RECT 4.124 24.848 4.196 24.88 ;
  LAYER M2 ;
        RECT 3.936 24.848 4.16 24.88 ;
  LAYER M1 ;
        RECT 3.92 24.828 3.952 24.9 ;
  LAYER M2 ;
        RECT 3.9 24.848 3.972 24.88 ;
  LAYER M1 ;
        RECT 3.92 14.748 3.952 14.82 ;
  LAYER M2 ;
        RECT 3.9 14.768 3.972 14.8 ;
  LAYER M1 ;
        RECT 3.92 14.784 3.952 15.204 ;
  LAYER M1 ;
        RECT 3.92 15.204 3.952 24.864 ;
  LAYER M1 ;
        RECT 10.096 21.72 10.128 21.792 ;
  LAYER M2 ;
        RECT 10.076 21.74 10.148 21.772 ;
  LAYER M1 ;
        RECT 10.096 21.588 10.128 21.756 ;
  LAYER M1 ;
        RECT 10.096 21.552 10.128 21.624 ;
  LAYER M2 ;
        RECT 10.076 21.572 10.148 21.604 ;
  LAYER M2 ;
        RECT 10.112 21.572 12.864 21.604 ;
  LAYER M1 ;
        RECT 12.848 21.552 12.88 21.624 ;
  LAYER M2 ;
        RECT 12.828 21.572 12.9 21.604 ;
  LAYER M1 ;
        RECT 10.096 18.612 10.128 18.684 ;
  LAYER M2 ;
        RECT 10.076 18.632 10.148 18.664 ;
  LAYER M1 ;
        RECT 10.096 18.48 10.128 18.648 ;
  LAYER M1 ;
        RECT 10.096 18.444 10.128 18.516 ;
  LAYER M2 ;
        RECT 10.076 18.464 10.148 18.496 ;
  LAYER M2 ;
        RECT 10.112 18.464 12.864 18.496 ;
  LAYER M1 ;
        RECT 12.848 18.444 12.88 18.516 ;
  LAYER M2 ;
        RECT 12.828 18.464 12.9 18.496 ;
  LAYER M1 ;
        RECT 12.848 14.748 12.88 14.82 ;
  LAYER M2 ;
        RECT 12.828 14.768 12.9 14.8 ;
  LAYER M1 ;
        RECT 12.848 14.784 12.88 15.204 ;
  LAYER M1 ;
        RECT 12.848 15.204 12.88 21.588 ;
  LAYER M2 ;
        RECT 3.936 14.768 12.864 14.8 ;
  LAYER M1 ;
        RECT 7.12 24.828 7.152 24.9 ;
  LAYER M2 ;
        RECT 7.1 24.848 7.172 24.88 ;
  LAYER M2 ;
        RECT 4.16 24.848 7.136 24.88 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 24.9 ;
  LAYER M2 ;
        RECT 4.124 24.848 4.196 24.88 ;
  LAYER M1 ;
        RECT 7.12 18.612 7.152 18.684 ;
  LAYER M2 ;
        RECT 7.1 18.632 7.172 18.664 ;
  LAYER M2 ;
        RECT 7.136 18.632 10.112 18.664 ;
  LAYER M1 ;
        RECT 10.096 18.612 10.128 18.684 ;
  LAYER M2 ;
        RECT 10.076 18.632 10.148 18.664 ;
  LAYER M1 ;
        RECT 1.168 27.936 1.2 28.008 ;
  LAYER M2 ;
        RECT 1.148 27.956 1.22 27.988 ;
  LAYER M2 ;
        RECT 0.96 27.956 1.184 27.988 ;
  LAYER M1 ;
        RECT 0.944 27.936 0.976 28.008 ;
  LAYER M2 ;
        RECT 0.924 27.956 0.996 27.988 ;
  LAYER M1 ;
        RECT 1.168 24.828 1.2 24.9 ;
  LAYER M2 ;
        RECT 1.148 24.848 1.22 24.88 ;
  LAYER M2 ;
        RECT 0.96 24.848 1.184 24.88 ;
  LAYER M1 ;
        RECT 0.944 24.828 0.976 24.9 ;
  LAYER M2 ;
        RECT 0.924 24.848 0.996 24.88 ;
  LAYER M1 ;
        RECT 1.168 21.72 1.2 21.792 ;
  LAYER M2 ;
        RECT 1.148 21.74 1.22 21.772 ;
  LAYER M2 ;
        RECT 0.96 21.74 1.184 21.772 ;
  LAYER M1 ;
        RECT 0.944 21.72 0.976 21.792 ;
  LAYER M2 ;
        RECT 0.924 21.74 0.996 21.772 ;
  LAYER M1 ;
        RECT 1.168 18.612 1.2 18.684 ;
  LAYER M2 ;
        RECT 1.148 18.632 1.22 18.664 ;
  LAYER M2 ;
        RECT 0.96 18.632 1.184 18.664 ;
  LAYER M1 ;
        RECT 0.944 18.612 0.976 18.684 ;
  LAYER M2 ;
        RECT 0.924 18.632 0.996 18.664 ;
  LAYER M1 ;
        RECT 1.168 15.504 1.2 15.576 ;
  LAYER M2 ;
        RECT 1.148 15.524 1.22 15.556 ;
  LAYER M2 ;
        RECT 0.96 15.524 1.184 15.556 ;
  LAYER M1 ;
        RECT 0.944 15.504 0.976 15.576 ;
  LAYER M2 ;
        RECT 0.924 15.524 0.996 15.556 ;
  LAYER M1 ;
        RECT 0.944 14.58 0.976 14.652 ;
  LAYER M2 ;
        RECT 0.924 14.6 0.996 14.632 ;
  LAYER M1 ;
        RECT 0.944 14.616 0.976 15.204 ;
  LAYER M1 ;
        RECT 0.944 15.204 0.976 27.972 ;
  LAYER M1 ;
        RECT 13.072 27.936 13.104 28.008 ;
  LAYER M2 ;
        RECT 13.052 27.956 13.124 27.988 ;
  LAYER M1 ;
        RECT 13.072 27.804 13.104 27.972 ;
  LAYER M1 ;
        RECT 13.072 27.768 13.104 27.84 ;
  LAYER M2 ;
        RECT 13.052 27.788 13.124 27.82 ;
  LAYER M2 ;
        RECT 13.088 27.788 15.84 27.82 ;
  LAYER M1 ;
        RECT 15.824 27.768 15.856 27.84 ;
  LAYER M2 ;
        RECT 15.804 27.788 15.876 27.82 ;
  LAYER M1 ;
        RECT 13.072 24.828 13.104 24.9 ;
  LAYER M2 ;
        RECT 13.052 24.848 13.124 24.88 ;
  LAYER M1 ;
        RECT 13.072 24.696 13.104 24.864 ;
  LAYER M1 ;
        RECT 13.072 24.66 13.104 24.732 ;
  LAYER M2 ;
        RECT 13.052 24.68 13.124 24.712 ;
  LAYER M2 ;
        RECT 13.088 24.68 15.84 24.712 ;
  LAYER M1 ;
        RECT 15.824 24.66 15.856 24.732 ;
  LAYER M2 ;
        RECT 15.804 24.68 15.876 24.712 ;
  LAYER M1 ;
        RECT 13.072 21.72 13.104 21.792 ;
  LAYER M2 ;
        RECT 13.052 21.74 13.124 21.772 ;
  LAYER M1 ;
        RECT 13.072 21.588 13.104 21.756 ;
  LAYER M1 ;
        RECT 13.072 21.552 13.104 21.624 ;
  LAYER M2 ;
        RECT 13.052 21.572 13.124 21.604 ;
  LAYER M2 ;
        RECT 13.088 21.572 15.84 21.604 ;
  LAYER M1 ;
        RECT 15.824 21.552 15.856 21.624 ;
  LAYER M2 ;
        RECT 15.804 21.572 15.876 21.604 ;
  LAYER M1 ;
        RECT 13.072 18.612 13.104 18.684 ;
  LAYER M2 ;
        RECT 13.052 18.632 13.124 18.664 ;
  LAYER M1 ;
        RECT 13.072 18.48 13.104 18.648 ;
  LAYER M1 ;
        RECT 13.072 18.444 13.104 18.516 ;
  LAYER M2 ;
        RECT 13.052 18.464 13.124 18.496 ;
  LAYER M2 ;
        RECT 13.088 18.464 15.84 18.496 ;
  LAYER M1 ;
        RECT 15.824 18.444 15.856 18.516 ;
  LAYER M2 ;
        RECT 15.804 18.464 15.876 18.496 ;
  LAYER M1 ;
        RECT 13.072 15.504 13.104 15.576 ;
  LAYER M2 ;
        RECT 13.052 15.524 13.124 15.556 ;
  LAYER M1 ;
        RECT 13.072 15.372 13.104 15.54 ;
  LAYER M1 ;
        RECT 13.072 15.336 13.104 15.408 ;
  LAYER M2 ;
        RECT 13.052 15.356 13.124 15.388 ;
  LAYER M2 ;
        RECT 13.088 15.356 15.84 15.388 ;
  LAYER M1 ;
        RECT 15.824 15.336 15.856 15.408 ;
  LAYER M2 ;
        RECT 15.804 15.356 15.876 15.388 ;
  LAYER M1 ;
        RECT 15.824 14.58 15.856 14.652 ;
  LAYER M2 ;
        RECT 15.804 14.6 15.876 14.632 ;
  LAYER M1 ;
        RECT 15.824 14.616 15.856 15.204 ;
  LAYER M1 ;
        RECT 15.824 15.204 15.856 27.804 ;
  LAYER M2 ;
        RECT 0.96 14.6 15.84 14.632 ;
  LAYER M1 ;
        RECT 4.144 27.936 4.176 28.008 ;
  LAYER M2 ;
        RECT 4.124 27.956 4.196 27.988 ;
  LAYER M2 ;
        RECT 1.184 27.956 4.16 27.988 ;
  LAYER M1 ;
        RECT 1.168 27.936 1.2 28.008 ;
  LAYER M2 ;
        RECT 1.148 27.956 1.22 27.988 ;
  LAYER M1 ;
        RECT 4.144 15.504 4.176 15.576 ;
  LAYER M2 ;
        RECT 4.124 15.524 4.196 15.556 ;
  LAYER M2 ;
        RECT 1.184 15.524 4.16 15.556 ;
  LAYER M1 ;
        RECT 1.168 15.504 1.2 15.576 ;
  LAYER M2 ;
        RECT 1.148 15.524 1.22 15.556 ;
  LAYER M1 ;
        RECT 7.12 15.504 7.152 15.576 ;
  LAYER M2 ;
        RECT 7.1 15.524 7.172 15.556 ;
  LAYER M2 ;
        RECT 4.16 15.524 7.136 15.556 ;
  LAYER M1 ;
        RECT 4.144 15.504 4.176 15.576 ;
  LAYER M2 ;
        RECT 4.124 15.524 4.196 15.556 ;
  LAYER M1 ;
        RECT 10.096 15.504 10.128 15.576 ;
  LAYER M2 ;
        RECT 10.076 15.524 10.148 15.556 ;
  LAYER M2 ;
        RECT 7.136 15.524 10.112 15.556 ;
  LAYER M1 ;
        RECT 7.12 15.504 7.152 15.576 ;
  LAYER M2 ;
        RECT 7.1 15.524 7.172 15.556 ;
  LAYER M1 ;
        RECT 10.096 27.936 10.128 28.008 ;
  LAYER M2 ;
        RECT 10.076 27.956 10.148 27.988 ;
  LAYER M2 ;
        RECT 10.112 27.956 13.088 27.988 ;
  LAYER M1 ;
        RECT 13.072 27.936 13.104 28.008 ;
  LAYER M2 ;
        RECT 13.052 27.956 13.124 27.988 ;
  LAYER M1 ;
        RECT 7.12 27.936 7.152 28.008 ;
  LAYER M2 ;
        RECT 7.1 27.956 7.172 27.988 ;
  LAYER M2 ;
        RECT 7.136 27.956 10.112 27.988 ;
  LAYER M1 ;
        RECT 10.096 27.936 10.128 28.008 ;
  LAYER M2 ;
        RECT 10.076 27.956 10.148 27.988 ;
  LAYER M1 ;
        RECT 1.168 27.936 1.2 30.444 ;
  LAYER M3 ;
        RECT 1.168 27.956 1.2 27.988 ;
  LAYER M1 ;
        RECT 1.232 27.936 1.264 30.444 ;
  LAYER M3 ;
        RECT 1.232 30.392 1.264 30.424 ;
  LAYER M1 ;
        RECT 1.296 27.936 1.328 30.444 ;
  LAYER M3 ;
        RECT 1.296 27.956 1.328 27.988 ;
  LAYER M1 ;
        RECT 1.36 27.936 1.392 30.444 ;
  LAYER M3 ;
        RECT 1.36 30.392 1.392 30.424 ;
  LAYER M1 ;
        RECT 1.424 27.936 1.456 30.444 ;
  LAYER M3 ;
        RECT 1.424 27.956 1.456 27.988 ;
  LAYER M1 ;
        RECT 1.488 27.936 1.52 30.444 ;
  LAYER M3 ;
        RECT 1.488 30.392 1.52 30.424 ;
  LAYER M1 ;
        RECT 1.552 27.936 1.584 30.444 ;
  LAYER M3 ;
        RECT 1.552 27.956 1.584 27.988 ;
  LAYER M1 ;
        RECT 1.616 27.936 1.648 30.444 ;
  LAYER M3 ;
        RECT 1.616 30.392 1.648 30.424 ;
  LAYER M1 ;
        RECT 1.68 27.936 1.712 30.444 ;
  LAYER M3 ;
        RECT 1.68 27.956 1.712 27.988 ;
  LAYER M1 ;
        RECT 1.744 27.936 1.776 30.444 ;
  LAYER M3 ;
        RECT 1.744 30.392 1.776 30.424 ;
  LAYER M1 ;
        RECT 1.808 27.936 1.84 30.444 ;
  LAYER M3 ;
        RECT 1.808 27.956 1.84 27.988 ;
  LAYER M1 ;
        RECT 1.872 27.936 1.904 30.444 ;
  LAYER M3 ;
        RECT 1.872 30.392 1.904 30.424 ;
  LAYER M1 ;
        RECT 1.936 27.936 1.968 30.444 ;
  LAYER M3 ;
        RECT 1.936 27.956 1.968 27.988 ;
  LAYER M1 ;
        RECT 2 27.936 2.032 30.444 ;
  LAYER M3 ;
        RECT 2 30.392 2.032 30.424 ;
  LAYER M1 ;
        RECT 2.064 27.936 2.096 30.444 ;
  LAYER M3 ;
        RECT 2.064 27.956 2.096 27.988 ;
  LAYER M1 ;
        RECT 2.128 27.936 2.16 30.444 ;
  LAYER M3 ;
        RECT 2.128 30.392 2.16 30.424 ;
  LAYER M1 ;
        RECT 2.192 27.936 2.224 30.444 ;
  LAYER M3 ;
        RECT 2.192 27.956 2.224 27.988 ;
  LAYER M1 ;
        RECT 2.256 27.936 2.288 30.444 ;
  LAYER M3 ;
        RECT 2.256 30.392 2.288 30.424 ;
  LAYER M1 ;
        RECT 2.32 27.936 2.352 30.444 ;
  LAYER M3 ;
        RECT 2.32 27.956 2.352 27.988 ;
  LAYER M1 ;
        RECT 2.384 27.936 2.416 30.444 ;
  LAYER M3 ;
        RECT 2.384 30.392 2.416 30.424 ;
  LAYER M1 ;
        RECT 2.448 27.936 2.48 30.444 ;
  LAYER M3 ;
        RECT 2.448 27.956 2.48 27.988 ;
  LAYER M1 ;
        RECT 2.512 27.936 2.544 30.444 ;
  LAYER M3 ;
        RECT 2.512 30.392 2.544 30.424 ;
  LAYER M1 ;
        RECT 2.576 27.936 2.608 30.444 ;
  LAYER M3 ;
        RECT 2.576 27.956 2.608 27.988 ;
  LAYER M1 ;
        RECT 2.64 27.936 2.672 30.444 ;
  LAYER M3 ;
        RECT 2.64 30.392 2.672 30.424 ;
  LAYER M1 ;
        RECT 2.704 27.936 2.736 30.444 ;
  LAYER M3 ;
        RECT 2.704 27.956 2.736 27.988 ;
  LAYER M1 ;
        RECT 2.768 27.936 2.8 30.444 ;
  LAYER M3 ;
        RECT 2.768 30.392 2.8 30.424 ;
  LAYER M1 ;
        RECT 2.832 27.936 2.864 30.444 ;
  LAYER M3 ;
        RECT 2.832 27.956 2.864 27.988 ;
  LAYER M1 ;
        RECT 2.896 27.936 2.928 30.444 ;
  LAYER M3 ;
        RECT 2.896 30.392 2.928 30.424 ;
  LAYER M1 ;
        RECT 2.96 27.936 2.992 30.444 ;
  LAYER M3 ;
        RECT 2.96 27.956 2.992 27.988 ;
  LAYER M1 ;
        RECT 3.024 27.936 3.056 30.444 ;
  LAYER M3 ;
        RECT 3.024 30.392 3.056 30.424 ;
  LAYER M1 ;
        RECT 3.088 27.936 3.12 30.444 ;
  LAYER M3 ;
        RECT 3.088 27.956 3.12 27.988 ;
  LAYER M1 ;
        RECT 3.152 27.936 3.184 30.444 ;
  LAYER M3 ;
        RECT 3.152 30.392 3.184 30.424 ;
  LAYER M1 ;
        RECT 3.216 27.936 3.248 30.444 ;
  LAYER M3 ;
        RECT 3.216 27.956 3.248 27.988 ;
  LAYER M1 ;
        RECT 3.28 27.936 3.312 30.444 ;
  LAYER M3 ;
        RECT 3.28 30.392 3.312 30.424 ;
  LAYER M1 ;
        RECT 3.344 27.936 3.376 30.444 ;
  LAYER M3 ;
        RECT 3.344 27.956 3.376 27.988 ;
  LAYER M1 ;
        RECT 3.408 27.936 3.44 30.444 ;
  LAYER M3 ;
        RECT 3.408 30.392 3.44 30.424 ;
  LAYER M1 ;
        RECT 3.472 27.936 3.504 30.444 ;
  LAYER M3 ;
        RECT 3.472 27.956 3.504 27.988 ;
  LAYER M1 ;
        RECT 3.536 27.936 3.568 30.444 ;
  LAYER M3 ;
        RECT 1.168 30.328 1.2 30.36 ;
  LAYER M2 ;
        RECT 3.536 30.264 3.568 30.296 ;
  LAYER M2 ;
        RECT 1.168 30.2 1.2 30.232 ;
  LAYER M2 ;
        RECT 3.536 30.136 3.568 30.168 ;
  LAYER M2 ;
        RECT 1.168 30.072 1.2 30.104 ;
  LAYER M2 ;
        RECT 3.536 30.008 3.568 30.04 ;
  LAYER M2 ;
        RECT 1.168 29.944 1.2 29.976 ;
  LAYER M2 ;
        RECT 3.536 29.88 3.568 29.912 ;
  LAYER M2 ;
        RECT 1.168 29.816 1.2 29.848 ;
  LAYER M2 ;
        RECT 3.536 29.752 3.568 29.784 ;
  LAYER M2 ;
        RECT 1.168 29.688 1.2 29.72 ;
  LAYER M2 ;
        RECT 3.536 29.624 3.568 29.656 ;
  LAYER M2 ;
        RECT 1.168 29.56 1.2 29.592 ;
  LAYER M2 ;
        RECT 3.536 29.496 3.568 29.528 ;
  LAYER M2 ;
        RECT 1.168 29.432 1.2 29.464 ;
  LAYER M2 ;
        RECT 3.536 29.368 3.568 29.4 ;
  LAYER M2 ;
        RECT 1.168 29.304 1.2 29.336 ;
  LAYER M2 ;
        RECT 3.536 29.24 3.568 29.272 ;
  LAYER M2 ;
        RECT 1.168 29.176 1.2 29.208 ;
  LAYER M2 ;
        RECT 3.536 29.112 3.568 29.144 ;
  LAYER M2 ;
        RECT 1.168 29.048 1.2 29.08 ;
  LAYER M2 ;
        RECT 3.536 28.984 3.568 29.016 ;
  LAYER M2 ;
        RECT 1.168 28.92 1.2 28.952 ;
  LAYER M2 ;
        RECT 3.536 28.856 3.568 28.888 ;
  LAYER M2 ;
        RECT 1.168 28.792 1.2 28.824 ;
  LAYER M2 ;
        RECT 3.536 28.728 3.568 28.76 ;
  LAYER M2 ;
        RECT 1.168 28.664 1.2 28.696 ;
  LAYER M2 ;
        RECT 3.536 28.6 3.568 28.632 ;
  LAYER M2 ;
        RECT 1.168 28.536 1.2 28.568 ;
  LAYER M2 ;
        RECT 3.536 28.472 3.568 28.504 ;
  LAYER M2 ;
        RECT 1.168 28.408 1.2 28.44 ;
  LAYER M2 ;
        RECT 3.536 28.344 3.568 28.376 ;
  LAYER M2 ;
        RECT 1.168 28.28 1.2 28.312 ;
  LAYER M2 ;
        RECT 3.536 28.216 3.568 28.248 ;
  LAYER M2 ;
        RECT 1.168 28.152 1.2 28.184 ;
  LAYER M2 ;
        RECT 3.536 28.088 3.568 28.12 ;
  LAYER M2 ;
        RECT 1.12 27.888 3.616 30.492 ;
  LAYER M1 ;
        RECT 1.168 24.828 1.2 27.336 ;
  LAYER M3 ;
        RECT 1.168 24.848 1.2 24.88 ;
  LAYER M1 ;
        RECT 1.232 24.828 1.264 27.336 ;
  LAYER M3 ;
        RECT 1.232 27.284 1.264 27.316 ;
  LAYER M1 ;
        RECT 1.296 24.828 1.328 27.336 ;
  LAYER M3 ;
        RECT 1.296 24.848 1.328 24.88 ;
  LAYER M1 ;
        RECT 1.36 24.828 1.392 27.336 ;
  LAYER M3 ;
        RECT 1.36 27.284 1.392 27.316 ;
  LAYER M1 ;
        RECT 1.424 24.828 1.456 27.336 ;
  LAYER M3 ;
        RECT 1.424 24.848 1.456 24.88 ;
  LAYER M1 ;
        RECT 1.488 24.828 1.52 27.336 ;
  LAYER M3 ;
        RECT 1.488 27.284 1.52 27.316 ;
  LAYER M1 ;
        RECT 1.552 24.828 1.584 27.336 ;
  LAYER M3 ;
        RECT 1.552 24.848 1.584 24.88 ;
  LAYER M1 ;
        RECT 1.616 24.828 1.648 27.336 ;
  LAYER M3 ;
        RECT 1.616 27.284 1.648 27.316 ;
  LAYER M1 ;
        RECT 1.68 24.828 1.712 27.336 ;
  LAYER M3 ;
        RECT 1.68 24.848 1.712 24.88 ;
  LAYER M1 ;
        RECT 1.744 24.828 1.776 27.336 ;
  LAYER M3 ;
        RECT 1.744 27.284 1.776 27.316 ;
  LAYER M1 ;
        RECT 1.808 24.828 1.84 27.336 ;
  LAYER M3 ;
        RECT 1.808 24.848 1.84 24.88 ;
  LAYER M1 ;
        RECT 1.872 24.828 1.904 27.336 ;
  LAYER M3 ;
        RECT 1.872 27.284 1.904 27.316 ;
  LAYER M1 ;
        RECT 1.936 24.828 1.968 27.336 ;
  LAYER M3 ;
        RECT 1.936 24.848 1.968 24.88 ;
  LAYER M1 ;
        RECT 2 24.828 2.032 27.336 ;
  LAYER M3 ;
        RECT 2 27.284 2.032 27.316 ;
  LAYER M1 ;
        RECT 2.064 24.828 2.096 27.336 ;
  LAYER M3 ;
        RECT 2.064 24.848 2.096 24.88 ;
  LAYER M1 ;
        RECT 2.128 24.828 2.16 27.336 ;
  LAYER M3 ;
        RECT 2.128 27.284 2.16 27.316 ;
  LAYER M1 ;
        RECT 2.192 24.828 2.224 27.336 ;
  LAYER M3 ;
        RECT 2.192 24.848 2.224 24.88 ;
  LAYER M1 ;
        RECT 2.256 24.828 2.288 27.336 ;
  LAYER M3 ;
        RECT 2.256 27.284 2.288 27.316 ;
  LAYER M1 ;
        RECT 2.32 24.828 2.352 27.336 ;
  LAYER M3 ;
        RECT 2.32 24.848 2.352 24.88 ;
  LAYER M1 ;
        RECT 2.384 24.828 2.416 27.336 ;
  LAYER M3 ;
        RECT 2.384 27.284 2.416 27.316 ;
  LAYER M1 ;
        RECT 2.448 24.828 2.48 27.336 ;
  LAYER M3 ;
        RECT 2.448 24.848 2.48 24.88 ;
  LAYER M1 ;
        RECT 2.512 24.828 2.544 27.336 ;
  LAYER M3 ;
        RECT 2.512 27.284 2.544 27.316 ;
  LAYER M1 ;
        RECT 2.576 24.828 2.608 27.336 ;
  LAYER M3 ;
        RECT 2.576 24.848 2.608 24.88 ;
  LAYER M1 ;
        RECT 2.64 24.828 2.672 27.336 ;
  LAYER M3 ;
        RECT 2.64 27.284 2.672 27.316 ;
  LAYER M1 ;
        RECT 2.704 24.828 2.736 27.336 ;
  LAYER M3 ;
        RECT 2.704 24.848 2.736 24.88 ;
  LAYER M1 ;
        RECT 2.768 24.828 2.8 27.336 ;
  LAYER M3 ;
        RECT 2.768 27.284 2.8 27.316 ;
  LAYER M1 ;
        RECT 2.832 24.828 2.864 27.336 ;
  LAYER M3 ;
        RECT 2.832 24.848 2.864 24.88 ;
  LAYER M1 ;
        RECT 2.896 24.828 2.928 27.336 ;
  LAYER M3 ;
        RECT 2.896 27.284 2.928 27.316 ;
  LAYER M1 ;
        RECT 2.96 24.828 2.992 27.336 ;
  LAYER M3 ;
        RECT 2.96 24.848 2.992 24.88 ;
  LAYER M1 ;
        RECT 3.024 24.828 3.056 27.336 ;
  LAYER M3 ;
        RECT 3.024 27.284 3.056 27.316 ;
  LAYER M1 ;
        RECT 3.088 24.828 3.12 27.336 ;
  LAYER M3 ;
        RECT 3.088 24.848 3.12 24.88 ;
  LAYER M1 ;
        RECT 3.152 24.828 3.184 27.336 ;
  LAYER M3 ;
        RECT 3.152 27.284 3.184 27.316 ;
  LAYER M1 ;
        RECT 3.216 24.828 3.248 27.336 ;
  LAYER M3 ;
        RECT 3.216 24.848 3.248 24.88 ;
  LAYER M1 ;
        RECT 3.28 24.828 3.312 27.336 ;
  LAYER M3 ;
        RECT 3.28 27.284 3.312 27.316 ;
  LAYER M1 ;
        RECT 3.344 24.828 3.376 27.336 ;
  LAYER M3 ;
        RECT 3.344 24.848 3.376 24.88 ;
  LAYER M1 ;
        RECT 3.408 24.828 3.44 27.336 ;
  LAYER M3 ;
        RECT 3.408 27.284 3.44 27.316 ;
  LAYER M1 ;
        RECT 3.472 24.828 3.504 27.336 ;
  LAYER M3 ;
        RECT 3.472 24.848 3.504 24.88 ;
  LAYER M1 ;
        RECT 3.536 24.828 3.568 27.336 ;
  LAYER M3 ;
        RECT 1.168 27.22 1.2 27.252 ;
  LAYER M2 ;
        RECT 3.536 27.156 3.568 27.188 ;
  LAYER M2 ;
        RECT 1.168 27.092 1.2 27.124 ;
  LAYER M2 ;
        RECT 3.536 27.028 3.568 27.06 ;
  LAYER M2 ;
        RECT 1.168 26.964 1.2 26.996 ;
  LAYER M2 ;
        RECT 3.536 26.9 3.568 26.932 ;
  LAYER M2 ;
        RECT 1.168 26.836 1.2 26.868 ;
  LAYER M2 ;
        RECT 3.536 26.772 3.568 26.804 ;
  LAYER M2 ;
        RECT 1.168 26.708 1.2 26.74 ;
  LAYER M2 ;
        RECT 3.536 26.644 3.568 26.676 ;
  LAYER M2 ;
        RECT 1.168 26.58 1.2 26.612 ;
  LAYER M2 ;
        RECT 3.536 26.516 3.568 26.548 ;
  LAYER M2 ;
        RECT 1.168 26.452 1.2 26.484 ;
  LAYER M2 ;
        RECT 3.536 26.388 3.568 26.42 ;
  LAYER M2 ;
        RECT 1.168 26.324 1.2 26.356 ;
  LAYER M2 ;
        RECT 3.536 26.26 3.568 26.292 ;
  LAYER M2 ;
        RECT 1.168 26.196 1.2 26.228 ;
  LAYER M2 ;
        RECT 3.536 26.132 3.568 26.164 ;
  LAYER M2 ;
        RECT 1.168 26.068 1.2 26.1 ;
  LAYER M2 ;
        RECT 3.536 26.004 3.568 26.036 ;
  LAYER M2 ;
        RECT 1.168 25.94 1.2 25.972 ;
  LAYER M2 ;
        RECT 3.536 25.876 3.568 25.908 ;
  LAYER M2 ;
        RECT 1.168 25.812 1.2 25.844 ;
  LAYER M2 ;
        RECT 3.536 25.748 3.568 25.78 ;
  LAYER M2 ;
        RECT 1.168 25.684 1.2 25.716 ;
  LAYER M2 ;
        RECT 3.536 25.62 3.568 25.652 ;
  LAYER M2 ;
        RECT 1.168 25.556 1.2 25.588 ;
  LAYER M2 ;
        RECT 3.536 25.492 3.568 25.524 ;
  LAYER M2 ;
        RECT 1.168 25.428 1.2 25.46 ;
  LAYER M2 ;
        RECT 3.536 25.364 3.568 25.396 ;
  LAYER M2 ;
        RECT 1.168 25.3 1.2 25.332 ;
  LAYER M2 ;
        RECT 3.536 25.236 3.568 25.268 ;
  LAYER M2 ;
        RECT 1.168 25.172 1.2 25.204 ;
  LAYER M2 ;
        RECT 3.536 25.108 3.568 25.14 ;
  LAYER M2 ;
        RECT 1.168 25.044 1.2 25.076 ;
  LAYER M2 ;
        RECT 3.536 24.98 3.568 25.012 ;
  LAYER M2 ;
        RECT 1.12 24.78 3.616 27.384 ;
  LAYER M1 ;
        RECT 1.168 21.72 1.2 24.228 ;
  LAYER M3 ;
        RECT 1.168 21.74 1.2 21.772 ;
  LAYER M1 ;
        RECT 1.232 21.72 1.264 24.228 ;
  LAYER M3 ;
        RECT 1.232 24.176 1.264 24.208 ;
  LAYER M1 ;
        RECT 1.296 21.72 1.328 24.228 ;
  LAYER M3 ;
        RECT 1.296 21.74 1.328 21.772 ;
  LAYER M1 ;
        RECT 1.36 21.72 1.392 24.228 ;
  LAYER M3 ;
        RECT 1.36 24.176 1.392 24.208 ;
  LAYER M1 ;
        RECT 1.424 21.72 1.456 24.228 ;
  LAYER M3 ;
        RECT 1.424 21.74 1.456 21.772 ;
  LAYER M1 ;
        RECT 1.488 21.72 1.52 24.228 ;
  LAYER M3 ;
        RECT 1.488 24.176 1.52 24.208 ;
  LAYER M1 ;
        RECT 1.552 21.72 1.584 24.228 ;
  LAYER M3 ;
        RECT 1.552 21.74 1.584 21.772 ;
  LAYER M1 ;
        RECT 1.616 21.72 1.648 24.228 ;
  LAYER M3 ;
        RECT 1.616 24.176 1.648 24.208 ;
  LAYER M1 ;
        RECT 1.68 21.72 1.712 24.228 ;
  LAYER M3 ;
        RECT 1.68 21.74 1.712 21.772 ;
  LAYER M1 ;
        RECT 1.744 21.72 1.776 24.228 ;
  LAYER M3 ;
        RECT 1.744 24.176 1.776 24.208 ;
  LAYER M1 ;
        RECT 1.808 21.72 1.84 24.228 ;
  LAYER M3 ;
        RECT 1.808 21.74 1.84 21.772 ;
  LAYER M1 ;
        RECT 1.872 21.72 1.904 24.228 ;
  LAYER M3 ;
        RECT 1.872 24.176 1.904 24.208 ;
  LAYER M1 ;
        RECT 1.936 21.72 1.968 24.228 ;
  LAYER M3 ;
        RECT 1.936 21.74 1.968 21.772 ;
  LAYER M1 ;
        RECT 2 21.72 2.032 24.228 ;
  LAYER M3 ;
        RECT 2 24.176 2.032 24.208 ;
  LAYER M1 ;
        RECT 2.064 21.72 2.096 24.228 ;
  LAYER M3 ;
        RECT 2.064 21.74 2.096 21.772 ;
  LAYER M1 ;
        RECT 2.128 21.72 2.16 24.228 ;
  LAYER M3 ;
        RECT 2.128 24.176 2.16 24.208 ;
  LAYER M1 ;
        RECT 2.192 21.72 2.224 24.228 ;
  LAYER M3 ;
        RECT 2.192 21.74 2.224 21.772 ;
  LAYER M1 ;
        RECT 2.256 21.72 2.288 24.228 ;
  LAYER M3 ;
        RECT 2.256 24.176 2.288 24.208 ;
  LAYER M1 ;
        RECT 2.32 21.72 2.352 24.228 ;
  LAYER M3 ;
        RECT 2.32 21.74 2.352 21.772 ;
  LAYER M1 ;
        RECT 2.384 21.72 2.416 24.228 ;
  LAYER M3 ;
        RECT 2.384 24.176 2.416 24.208 ;
  LAYER M1 ;
        RECT 2.448 21.72 2.48 24.228 ;
  LAYER M3 ;
        RECT 2.448 21.74 2.48 21.772 ;
  LAYER M1 ;
        RECT 2.512 21.72 2.544 24.228 ;
  LAYER M3 ;
        RECT 2.512 24.176 2.544 24.208 ;
  LAYER M1 ;
        RECT 2.576 21.72 2.608 24.228 ;
  LAYER M3 ;
        RECT 2.576 21.74 2.608 21.772 ;
  LAYER M1 ;
        RECT 2.64 21.72 2.672 24.228 ;
  LAYER M3 ;
        RECT 2.64 24.176 2.672 24.208 ;
  LAYER M1 ;
        RECT 2.704 21.72 2.736 24.228 ;
  LAYER M3 ;
        RECT 2.704 21.74 2.736 21.772 ;
  LAYER M1 ;
        RECT 2.768 21.72 2.8 24.228 ;
  LAYER M3 ;
        RECT 2.768 24.176 2.8 24.208 ;
  LAYER M1 ;
        RECT 2.832 21.72 2.864 24.228 ;
  LAYER M3 ;
        RECT 2.832 21.74 2.864 21.772 ;
  LAYER M1 ;
        RECT 2.896 21.72 2.928 24.228 ;
  LAYER M3 ;
        RECT 2.896 24.176 2.928 24.208 ;
  LAYER M1 ;
        RECT 2.96 21.72 2.992 24.228 ;
  LAYER M3 ;
        RECT 2.96 21.74 2.992 21.772 ;
  LAYER M1 ;
        RECT 3.024 21.72 3.056 24.228 ;
  LAYER M3 ;
        RECT 3.024 24.176 3.056 24.208 ;
  LAYER M1 ;
        RECT 3.088 21.72 3.12 24.228 ;
  LAYER M3 ;
        RECT 3.088 21.74 3.12 21.772 ;
  LAYER M1 ;
        RECT 3.152 21.72 3.184 24.228 ;
  LAYER M3 ;
        RECT 3.152 24.176 3.184 24.208 ;
  LAYER M1 ;
        RECT 3.216 21.72 3.248 24.228 ;
  LAYER M3 ;
        RECT 3.216 21.74 3.248 21.772 ;
  LAYER M1 ;
        RECT 3.28 21.72 3.312 24.228 ;
  LAYER M3 ;
        RECT 3.28 24.176 3.312 24.208 ;
  LAYER M1 ;
        RECT 3.344 21.72 3.376 24.228 ;
  LAYER M3 ;
        RECT 3.344 21.74 3.376 21.772 ;
  LAYER M1 ;
        RECT 3.408 21.72 3.44 24.228 ;
  LAYER M3 ;
        RECT 3.408 24.176 3.44 24.208 ;
  LAYER M1 ;
        RECT 3.472 21.72 3.504 24.228 ;
  LAYER M3 ;
        RECT 3.472 21.74 3.504 21.772 ;
  LAYER M1 ;
        RECT 3.536 21.72 3.568 24.228 ;
  LAYER M3 ;
        RECT 1.168 24.112 1.2 24.144 ;
  LAYER M2 ;
        RECT 3.536 24.048 3.568 24.08 ;
  LAYER M2 ;
        RECT 1.168 23.984 1.2 24.016 ;
  LAYER M2 ;
        RECT 3.536 23.92 3.568 23.952 ;
  LAYER M2 ;
        RECT 1.168 23.856 1.2 23.888 ;
  LAYER M2 ;
        RECT 3.536 23.792 3.568 23.824 ;
  LAYER M2 ;
        RECT 1.168 23.728 1.2 23.76 ;
  LAYER M2 ;
        RECT 3.536 23.664 3.568 23.696 ;
  LAYER M2 ;
        RECT 1.168 23.6 1.2 23.632 ;
  LAYER M2 ;
        RECT 3.536 23.536 3.568 23.568 ;
  LAYER M2 ;
        RECT 1.168 23.472 1.2 23.504 ;
  LAYER M2 ;
        RECT 3.536 23.408 3.568 23.44 ;
  LAYER M2 ;
        RECT 1.168 23.344 1.2 23.376 ;
  LAYER M2 ;
        RECT 3.536 23.28 3.568 23.312 ;
  LAYER M2 ;
        RECT 1.168 23.216 1.2 23.248 ;
  LAYER M2 ;
        RECT 3.536 23.152 3.568 23.184 ;
  LAYER M2 ;
        RECT 1.168 23.088 1.2 23.12 ;
  LAYER M2 ;
        RECT 3.536 23.024 3.568 23.056 ;
  LAYER M2 ;
        RECT 1.168 22.96 1.2 22.992 ;
  LAYER M2 ;
        RECT 3.536 22.896 3.568 22.928 ;
  LAYER M2 ;
        RECT 1.168 22.832 1.2 22.864 ;
  LAYER M2 ;
        RECT 3.536 22.768 3.568 22.8 ;
  LAYER M2 ;
        RECT 1.168 22.704 1.2 22.736 ;
  LAYER M2 ;
        RECT 3.536 22.64 3.568 22.672 ;
  LAYER M2 ;
        RECT 1.168 22.576 1.2 22.608 ;
  LAYER M2 ;
        RECT 3.536 22.512 3.568 22.544 ;
  LAYER M2 ;
        RECT 1.168 22.448 1.2 22.48 ;
  LAYER M2 ;
        RECT 3.536 22.384 3.568 22.416 ;
  LAYER M2 ;
        RECT 1.168 22.32 1.2 22.352 ;
  LAYER M2 ;
        RECT 3.536 22.256 3.568 22.288 ;
  LAYER M2 ;
        RECT 1.168 22.192 1.2 22.224 ;
  LAYER M2 ;
        RECT 3.536 22.128 3.568 22.16 ;
  LAYER M2 ;
        RECT 1.168 22.064 1.2 22.096 ;
  LAYER M2 ;
        RECT 3.536 22 3.568 22.032 ;
  LAYER M2 ;
        RECT 1.168 21.936 1.2 21.968 ;
  LAYER M2 ;
        RECT 3.536 21.872 3.568 21.904 ;
  LAYER M2 ;
        RECT 1.12 21.672 3.616 24.276 ;
  LAYER M1 ;
        RECT 1.168 18.612 1.2 21.12 ;
  LAYER M3 ;
        RECT 1.168 18.632 1.2 18.664 ;
  LAYER M1 ;
        RECT 1.232 18.612 1.264 21.12 ;
  LAYER M3 ;
        RECT 1.232 21.068 1.264 21.1 ;
  LAYER M1 ;
        RECT 1.296 18.612 1.328 21.12 ;
  LAYER M3 ;
        RECT 1.296 18.632 1.328 18.664 ;
  LAYER M1 ;
        RECT 1.36 18.612 1.392 21.12 ;
  LAYER M3 ;
        RECT 1.36 21.068 1.392 21.1 ;
  LAYER M1 ;
        RECT 1.424 18.612 1.456 21.12 ;
  LAYER M3 ;
        RECT 1.424 18.632 1.456 18.664 ;
  LAYER M1 ;
        RECT 1.488 18.612 1.52 21.12 ;
  LAYER M3 ;
        RECT 1.488 21.068 1.52 21.1 ;
  LAYER M1 ;
        RECT 1.552 18.612 1.584 21.12 ;
  LAYER M3 ;
        RECT 1.552 18.632 1.584 18.664 ;
  LAYER M1 ;
        RECT 1.616 18.612 1.648 21.12 ;
  LAYER M3 ;
        RECT 1.616 21.068 1.648 21.1 ;
  LAYER M1 ;
        RECT 1.68 18.612 1.712 21.12 ;
  LAYER M3 ;
        RECT 1.68 18.632 1.712 18.664 ;
  LAYER M1 ;
        RECT 1.744 18.612 1.776 21.12 ;
  LAYER M3 ;
        RECT 1.744 21.068 1.776 21.1 ;
  LAYER M1 ;
        RECT 1.808 18.612 1.84 21.12 ;
  LAYER M3 ;
        RECT 1.808 18.632 1.84 18.664 ;
  LAYER M1 ;
        RECT 1.872 18.612 1.904 21.12 ;
  LAYER M3 ;
        RECT 1.872 21.068 1.904 21.1 ;
  LAYER M1 ;
        RECT 1.936 18.612 1.968 21.12 ;
  LAYER M3 ;
        RECT 1.936 18.632 1.968 18.664 ;
  LAYER M1 ;
        RECT 2 18.612 2.032 21.12 ;
  LAYER M3 ;
        RECT 2 21.068 2.032 21.1 ;
  LAYER M1 ;
        RECT 2.064 18.612 2.096 21.12 ;
  LAYER M3 ;
        RECT 2.064 18.632 2.096 18.664 ;
  LAYER M1 ;
        RECT 2.128 18.612 2.16 21.12 ;
  LAYER M3 ;
        RECT 2.128 21.068 2.16 21.1 ;
  LAYER M1 ;
        RECT 2.192 18.612 2.224 21.12 ;
  LAYER M3 ;
        RECT 2.192 18.632 2.224 18.664 ;
  LAYER M1 ;
        RECT 2.256 18.612 2.288 21.12 ;
  LAYER M3 ;
        RECT 2.256 21.068 2.288 21.1 ;
  LAYER M1 ;
        RECT 2.32 18.612 2.352 21.12 ;
  LAYER M3 ;
        RECT 2.32 18.632 2.352 18.664 ;
  LAYER M1 ;
        RECT 2.384 18.612 2.416 21.12 ;
  LAYER M3 ;
        RECT 2.384 21.068 2.416 21.1 ;
  LAYER M1 ;
        RECT 2.448 18.612 2.48 21.12 ;
  LAYER M3 ;
        RECT 2.448 18.632 2.48 18.664 ;
  LAYER M1 ;
        RECT 2.512 18.612 2.544 21.12 ;
  LAYER M3 ;
        RECT 2.512 21.068 2.544 21.1 ;
  LAYER M1 ;
        RECT 2.576 18.612 2.608 21.12 ;
  LAYER M3 ;
        RECT 2.576 18.632 2.608 18.664 ;
  LAYER M1 ;
        RECT 2.64 18.612 2.672 21.12 ;
  LAYER M3 ;
        RECT 2.64 21.068 2.672 21.1 ;
  LAYER M1 ;
        RECT 2.704 18.612 2.736 21.12 ;
  LAYER M3 ;
        RECT 2.704 18.632 2.736 18.664 ;
  LAYER M1 ;
        RECT 2.768 18.612 2.8 21.12 ;
  LAYER M3 ;
        RECT 2.768 21.068 2.8 21.1 ;
  LAYER M1 ;
        RECT 2.832 18.612 2.864 21.12 ;
  LAYER M3 ;
        RECT 2.832 18.632 2.864 18.664 ;
  LAYER M1 ;
        RECT 2.896 18.612 2.928 21.12 ;
  LAYER M3 ;
        RECT 2.896 21.068 2.928 21.1 ;
  LAYER M1 ;
        RECT 2.96 18.612 2.992 21.12 ;
  LAYER M3 ;
        RECT 2.96 18.632 2.992 18.664 ;
  LAYER M1 ;
        RECT 3.024 18.612 3.056 21.12 ;
  LAYER M3 ;
        RECT 3.024 21.068 3.056 21.1 ;
  LAYER M1 ;
        RECT 3.088 18.612 3.12 21.12 ;
  LAYER M3 ;
        RECT 3.088 18.632 3.12 18.664 ;
  LAYER M1 ;
        RECT 3.152 18.612 3.184 21.12 ;
  LAYER M3 ;
        RECT 3.152 21.068 3.184 21.1 ;
  LAYER M1 ;
        RECT 3.216 18.612 3.248 21.12 ;
  LAYER M3 ;
        RECT 3.216 18.632 3.248 18.664 ;
  LAYER M1 ;
        RECT 3.28 18.612 3.312 21.12 ;
  LAYER M3 ;
        RECT 3.28 21.068 3.312 21.1 ;
  LAYER M1 ;
        RECT 3.344 18.612 3.376 21.12 ;
  LAYER M3 ;
        RECT 3.344 18.632 3.376 18.664 ;
  LAYER M1 ;
        RECT 3.408 18.612 3.44 21.12 ;
  LAYER M3 ;
        RECT 3.408 21.068 3.44 21.1 ;
  LAYER M1 ;
        RECT 3.472 18.612 3.504 21.12 ;
  LAYER M3 ;
        RECT 3.472 18.632 3.504 18.664 ;
  LAYER M1 ;
        RECT 3.536 18.612 3.568 21.12 ;
  LAYER M3 ;
        RECT 1.168 21.004 1.2 21.036 ;
  LAYER M2 ;
        RECT 3.536 20.94 3.568 20.972 ;
  LAYER M2 ;
        RECT 1.168 20.876 1.2 20.908 ;
  LAYER M2 ;
        RECT 3.536 20.812 3.568 20.844 ;
  LAYER M2 ;
        RECT 1.168 20.748 1.2 20.78 ;
  LAYER M2 ;
        RECT 3.536 20.684 3.568 20.716 ;
  LAYER M2 ;
        RECT 1.168 20.62 1.2 20.652 ;
  LAYER M2 ;
        RECT 3.536 20.556 3.568 20.588 ;
  LAYER M2 ;
        RECT 1.168 20.492 1.2 20.524 ;
  LAYER M2 ;
        RECT 3.536 20.428 3.568 20.46 ;
  LAYER M2 ;
        RECT 1.168 20.364 1.2 20.396 ;
  LAYER M2 ;
        RECT 3.536 20.3 3.568 20.332 ;
  LAYER M2 ;
        RECT 1.168 20.236 1.2 20.268 ;
  LAYER M2 ;
        RECT 3.536 20.172 3.568 20.204 ;
  LAYER M2 ;
        RECT 1.168 20.108 1.2 20.14 ;
  LAYER M2 ;
        RECT 3.536 20.044 3.568 20.076 ;
  LAYER M2 ;
        RECT 1.168 19.98 1.2 20.012 ;
  LAYER M2 ;
        RECT 3.536 19.916 3.568 19.948 ;
  LAYER M2 ;
        RECT 1.168 19.852 1.2 19.884 ;
  LAYER M2 ;
        RECT 3.536 19.788 3.568 19.82 ;
  LAYER M2 ;
        RECT 1.168 19.724 1.2 19.756 ;
  LAYER M2 ;
        RECT 3.536 19.66 3.568 19.692 ;
  LAYER M2 ;
        RECT 1.168 19.596 1.2 19.628 ;
  LAYER M2 ;
        RECT 3.536 19.532 3.568 19.564 ;
  LAYER M2 ;
        RECT 1.168 19.468 1.2 19.5 ;
  LAYER M2 ;
        RECT 3.536 19.404 3.568 19.436 ;
  LAYER M2 ;
        RECT 1.168 19.34 1.2 19.372 ;
  LAYER M2 ;
        RECT 3.536 19.276 3.568 19.308 ;
  LAYER M2 ;
        RECT 1.168 19.212 1.2 19.244 ;
  LAYER M2 ;
        RECT 3.536 19.148 3.568 19.18 ;
  LAYER M2 ;
        RECT 1.168 19.084 1.2 19.116 ;
  LAYER M2 ;
        RECT 3.536 19.02 3.568 19.052 ;
  LAYER M2 ;
        RECT 1.168 18.956 1.2 18.988 ;
  LAYER M2 ;
        RECT 3.536 18.892 3.568 18.924 ;
  LAYER M2 ;
        RECT 1.168 18.828 1.2 18.86 ;
  LAYER M2 ;
        RECT 3.536 18.764 3.568 18.796 ;
  LAYER M2 ;
        RECT 1.12 18.564 3.616 21.168 ;
  LAYER M1 ;
        RECT 1.168 15.504 1.2 18.012 ;
  LAYER M3 ;
        RECT 1.168 15.524 1.2 15.556 ;
  LAYER M1 ;
        RECT 1.232 15.504 1.264 18.012 ;
  LAYER M3 ;
        RECT 1.232 17.96 1.264 17.992 ;
  LAYER M1 ;
        RECT 1.296 15.504 1.328 18.012 ;
  LAYER M3 ;
        RECT 1.296 15.524 1.328 15.556 ;
  LAYER M1 ;
        RECT 1.36 15.504 1.392 18.012 ;
  LAYER M3 ;
        RECT 1.36 17.96 1.392 17.992 ;
  LAYER M1 ;
        RECT 1.424 15.504 1.456 18.012 ;
  LAYER M3 ;
        RECT 1.424 15.524 1.456 15.556 ;
  LAYER M1 ;
        RECT 1.488 15.504 1.52 18.012 ;
  LAYER M3 ;
        RECT 1.488 17.96 1.52 17.992 ;
  LAYER M1 ;
        RECT 1.552 15.504 1.584 18.012 ;
  LAYER M3 ;
        RECT 1.552 15.524 1.584 15.556 ;
  LAYER M1 ;
        RECT 1.616 15.504 1.648 18.012 ;
  LAYER M3 ;
        RECT 1.616 17.96 1.648 17.992 ;
  LAYER M1 ;
        RECT 1.68 15.504 1.712 18.012 ;
  LAYER M3 ;
        RECT 1.68 15.524 1.712 15.556 ;
  LAYER M1 ;
        RECT 1.744 15.504 1.776 18.012 ;
  LAYER M3 ;
        RECT 1.744 17.96 1.776 17.992 ;
  LAYER M1 ;
        RECT 1.808 15.504 1.84 18.012 ;
  LAYER M3 ;
        RECT 1.808 15.524 1.84 15.556 ;
  LAYER M1 ;
        RECT 1.872 15.504 1.904 18.012 ;
  LAYER M3 ;
        RECT 1.872 17.96 1.904 17.992 ;
  LAYER M1 ;
        RECT 1.936 15.504 1.968 18.012 ;
  LAYER M3 ;
        RECT 1.936 15.524 1.968 15.556 ;
  LAYER M1 ;
        RECT 2 15.504 2.032 18.012 ;
  LAYER M3 ;
        RECT 2 17.96 2.032 17.992 ;
  LAYER M1 ;
        RECT 2.064 15.504 2.096 18.012 ;
  LAYER M3 ;
        RECT 2.064 15.524 2.096 15.556 ;
  LAYER M1 ;
        RECT 2.128 15.504 2.16 18.012 ;
  LAYER M3 ;
        RECT 2.128 17.96 2.16 17.992 ;
  LAYER M1 ;
        RECT 2.192 15.504 2.224 18.012 ;
  LAYER M3 ;
        RECT 2.192 15.524 2.224 15.556 ;
  LAYER M1 ;
        RECT 2.256 15.504 2.288 18.012 ;
  LAYER M3 ;
        RECT 2.256 17.96 2.288 17.992 ;
  LAYER M1 ;
        RECT 2.32 15.504 2.352 18.012 ;
  LAYER M3 ;
        RECT 2.32 15.524 2.352 15.556 ;
  LAYER M1 ;
        RECT 2.384 15.504 2.416 18.012 ;
  LAYER M3 ;
        RECT 2.384 17.96 2.416 17.992 ;
  LAYER M1 ;
        RECT 2.448 15.504 2.48 18.012 ;
  LAYER M3 ;
        RECT 2.448 15.524 2.48 15.556 ;
  LAYER M1 ;
        RECT 2.512 15.504 2.544 18.012 ;
  LAYER M3 ;
        RECT 2.512 17.96 2.544 17.992 ;
  LAYER M1 ;
        RECT 2.576 15.504 2.608 18.012 ;
  LAYER M3 ;
        RECT 2.576 15.524 2.608 15.556 ;
  LAYER M1 ;
        RECT 2.64 15.504 2.672 18.012 ;
  LAYER M3 ;
        RECT 2.64 17.96 2.672 17.992 ;
  LAYER M1 ;
        RECT 2.704 15.504 2.736 18.012 ;
  LAYER M3 ;
        RECT 2.704 15.524 2.736 15.556 ;
  LAYER M1 ;
        RECT 2.768 15.504 2.8 18.012 ;
  LAYER M3 ;
        RECT 2.768 17.96 2.8 17.992 ;
  LAYER M1 ;
        RECT 2.832 15.504 2.864 18.012 ;
  LAYER M3 ;
        RECT 2.832 15.524 2.864 15.556 ;
  LAYER M1 ;
        RECT 2.896 15.504 2.928 18.012 ;
  LAYER M3 ;
        RECT 2.896 17.96 2.928 17.992 ;
  LAYER M1 ;
        RECT 2.96 15.504 2.992 18.012 ;
  LAYER M3 ;
        RECT 2.96 15.524 2.992 15.556 ;
  LAYER M1 ;
        RECT 3.024 15.504 3.056 18.012 ;
  LAYER M3 ;
        RECT 3.024 17.96 3.056 17.992 ;
  LAYER M1 ;
        RECT 3.088 15.504 3.12 18.012 ;
  LAYER M3 ;
        RECT 3.088 15.524 3.12 15.556 ;
  LAYER M1 ;
        RECT 3.152 15.504 3.184 18.012 ;
  LAYER M3 ;
        RECT 3.152 17.96 3.184 17.992 ;
  LAYER M1 ;
        RECT 3.216 15.504 3.248 18.012 ;
  LAYER M3 ;
        RECT 3.216 15.524 3.248 15.556 ;
  LAYER M1 ;
        RECT 3.28 15.504 3.312 18.012 ;
  LAYER M3 ;
        RECT 3.28 17.96 3.312 17.992 ;
  LAYER M1 ;
        RECT 3.344 15.504 3.376 18.012 ;
  LAYER M3 ;
        RECT 3.344 15.524 3.376 15.556 ;
  LAYER M1 ;
        RECT 3.408 15.504 3.44 18.012 ;
  LAYER M3 ;
        RECT 3.408 17.96 3.44 17.992 ;
  LAYER M1 ;
        RECT 3.472 15.504 3.504 18.012 ;
  LAYER M3 ;
        RECT 3.472 15.524 3.504 15.556 ;
  LAYER M1 ;
        RECT 3.536 15.504 3.568 18.012 ;
  LAYER M3 ;
        RECT 1.168 17.896 1.2 17.928 ;
  LAYER M2 ;
        RECT 3.536 17.832 3.568 17.864 ;
  LAYER M2 ;
        RECT 1.168 17.768 1.2 17.8 ;
  LAYER M2 ;
        RECT 3.536 17.704 3.568 17.736 ;
  LAYER M2 ;
        RECT 1.168 17.64 1.2 17.672 ;
  LAYER M2 ;
        RECT 3.536 17.576 3.568 17.608 ;
  LAYER M2 ;
        RECT 1.168 17.512 1.2 17.544 ;
  LAYER M2 ;
        RECT 3.536 17.448 3.568 17.48 ;
  LAYER M2 ;
        RECT 1.168 17.384 1.2 17.416 ;
  LAYER M2 ;
        RECT 3.536 17.32 3.568 17.352 ;
  LAYER M2 ;
        RECT 1.168 17.256 1.2 17.288 ;
  LAYER M2 ;
        RECT 3.536 17.192 3.568 17.224 ;
  LAYER M2 ;
        RECT 1.168 17.128 1.2 17.16 ;
  LAYER M2 ;
        RECT 3.536 17.064 3.568 17.096 ;
  LAYER M2 ;
        RECT 1.168 17 1.2 17.032 ;
  LAYER M2 ;
        RECT 3.536 16.936 3.568 16.968 ;
  LAYER M2 ;
        RECT 1.168 16.872 1.2 16.904 ;
  LAYER M2 ;
        RECT 3.536 16.808 3.568 16.84 ;
  LAYER M2 ;
        RECT 1.168 16.744 1.2 16.776 ;
  LAYER M2 ;
        RECT 3.536 16.68 3.568 16.712 ;
  LAYER M2 ;
        RECT 1.168 16.616 1.2 16.648 ;
  LAYER M2 ;
        RECT 3.536 16.552 3.568 16.584 ;
  LAYER M2 ;
        RECT 1.168 16.488 1.2 16.52 ;
  LAYER M2 ;
        RECT 3.536 16.424 3.568 16.456 ;
  LAYER M2 ;
        RECT 1.168 16.36 1.2 16.392 ;
  LAYER M2 ;
        RECT 3.536 16.296 3.568 16.328 ;
  LAYER M2 ;
        RECT 1.168 16.232 1.2 16.264 ;
  LAYER M2 ;
        RECT 3.536 16.168 3.568 16.2 ;
  LAYER M2 ;
        RECT 1.168 16.104 1.2 16.136 ;
  LAYER M2 ;
        RECT 3.536 16.04 3.568 16.072 ;
  LAYER M2 ;
        RECT 1.168 15.976 1.2 16.008 ;
  LAYER M2 ;
        RECT 3.536 15.912 3.568 15.944 ;
  LAYER M2 ;
        RECT 1.168 15.848 1.2 15.88 ;
  LAYER M2 ;
        RECT 3.536 15.784 3.568 15.816 ;
  LAYER M2 ;
        RECT 1.168 15.72 1.2 15.752 ;
  LAYER M2 ;
        RECT 3.536 15.656 3.568 15.688 ;
  LAYER M2 ;
        RECT 1.12 15.456 3.616 18.06 ;
  LAYER M1 ;
        RECT 4.144 27.936 4.176 30.444 ;
  LAYER M3 ;
        RECT 4.144 27.956 4.176 27.988 ;
  LAYER M1 ;
        RECT 4.208 27.936 4.24 30.444 ;
  LAYER M3 ;
        RECT 4.208 30.392 4.24 30.424 ;
  LAYER M1 ;
        RECT 4.272 27.936 4.304 30.444 ;
  LAYER M3 ;
        RECT 4.272 27.956 4.304 27.988 ;
  LAYER M1 ;
        RECT 4.336 27.936 4.368 30.444 ;
  LAYER M3 ;
        RECT 4.336 30.392 4.368 30.424 ;
  LAYER M1 ;
        RECT 4.4 27.936 4.432 30.444 ;
  LAYER M3 ;
        RECT 4.4 27.956 4.432 27.988 ;
  LAYER M1 ;
        RECT 4.464 27.936 4.496 30.444 ;
  LAYER M3 ;
        RECT 4.464 30.392 4.496 30.424 ;
  LAYER M1 ;
        RECT 4.528 27.936 4.56 30.444 ;
  LAYER M3 ;
        RECT 4.528 27.956 4.56 27.988 ;
  LAYER M1 ;
        RECT 4.592 27.936 4.624 30.444 ;
  LAYER M3 ;
        RECT 4.592 30.392 4.624 30.424 ;
  LAYER M1 ;
        RECT 4.656 27.936 4.688 30.444 ;
  LAYER M3 ;
        RECT 4.656 27.956 4.688 27.988 ;
  LAYER M1 ;
        RECT 4.72 27.936 4.752 30.444 ;
  LAYER M3 ;
        RECT 4.72 30.392 4.752 30.424 ;
  LAYER M1 ;
        RECT 4.784 27.936 4.816 30.444 ;
  LAYER M3 ;
        RECT 4.784 27.956 4.816 27.988 ;
  LAYER M1 ;
        RECT 4.848 27.936 4.88 30.444 ;
  LAYER M3 ;
        RECT 4.848 30.392 4.88 30.424 ;
  LAYER M1 ;
        RECT 4.912 27.936 4.944 30.444 ;
  LAYER M3 ;
        RECT 4.912 27.956 4.944 27.988 ;
  LAYER M1 ;
        RECT 4.976 27.936 5.008 30.444 ;
  LAYER M3 ;
        RECT 4.976 30.392 5.008 30.424 ;
  LAYER M1 ;
        RECT 5.04 27.936 5.072 30.444 ;
  LAYER M3 ;
        RECT 5.04 27.956 5.072 27.988 ;
  LAYER M1 ;
        RECT 5.104 27.936 5.136 30.444 ;
  LAYER M3 ;
        RECT 5.104 30.392 5.136 30.424 ;
  LAYER M1 ;
        RECT 5.168 27.936 5.2 30.444 ;
  LAYER M3 ;
        RECT 5.168 27.956 5.2 27.988 ;
  LAYER M1 ;
        RECT 5.232 27.936 5.264 30.444 ;
  LAYER M3 ;
        RECT 5.232 30.392 5.264 30.424 ;
  LAYER M1 ;
        RECT 5.296 27.936 5.328 30.444 ;
  LAYER M3 ;
        RECT 5.296 27.956 5.328 27.988 ;
  LAYER M1 ;
        RECT 5.36 27.936 5.392 30.444 ;
  LAYER M3 ;
        RECT 5.36 30.392 5.392 30.424 ;
  LAYER M1 ;
        RECT 5.424 27.936 5.456 30.444 ;
  LAYER M3 ;
        RECT 5.424 27.956 5.456 27.988 ;
  LAYER M1 ;
        RECT 5.488 27.936 5.52 30.444 ;
  LAYER M3 ;
        RECT 5.488 30.392 5.52 30.424 ;
  LAYER M1 ;
        RECT 5.552 27.936 5.584 30.444 ;
  LAYER M3 ;
        RECT 5.552 27.956 5.584 27.988 ;
  LAYER M1 ;
        RECT 5.616 27.936 5.648 30.444 ;
  LAYER M3 ;
        RECT 5.616 30.392 5.648 30.424 ;
  LAYER M1 ;
        RECT 5.68 27.936 5.712 30.444 ;
  LAYER M3 ;
        RECT 5.68 27.956 5.712 27.988 ;
  LAYER M1 ;
        RECT 5.744 27.936 5.776 30.444 ;
  LAYER M3 ;
        RECT 5.744 30.392 5.776 30.424 ;
  LAYER M1 ;
        RECT 5.808 27.936 5.84 30.444 ;
  LAYER M3 ;
        RECT 5.808 27.956 5.84 27.988 ;
  LAYER M1 ;
        RECT 5.872 27.936 5.904 30.444 ;
  LAYER M3 ;
        RECT 5.872 30.392 5.904 30.424 ;
  LAYER M1 ;
        RECT 5.936 27.936 5.968 30.444 ;
  LAYER M3 ;
        RECT 5.936 27.956 5.968 27.988 ;
  LAYER M1 ;
        RECT 6 27.936 6.032 30.444 ;
  LAYER M3 ;
        RECT 6 30.392 6.032 30.424 ;
  LAYER M1 ;
        RECT 6.064 27.936 6.096 30.444 ;
  LAYER M3 ;
        RECT 6.064 27.956 6.096 27.988 ;
  LAYER M1 ;
        RECT 6.128 27.936 6.16 30.444 ;
  LAYER M3 ;
        RECT 6.128 30.392 6.16 30.424 ;
  LAYER M1 ;
        RECT 6.192 27.936 6.224 30.444 ;
  LAYER M3 ;
        RECT 6.192 27.956 6.224 27.988 ;
  LAYER M1 ;
        RECT 6.256 27.936 6.288 30.444 ;
  LAYER M3 ;
        RECT 6.256 30.392 6.288 30.424 ;
  LAYER M1 ;
        RECT 6.32 27.936 6.352 30.444 ;
  LAYER M3 ;
        RECT 6.32 27.956 6.352 27.988 ;
  LAYER M1 ;
        RECT 6.384 27.936 6.416 30.444 ;
  LAYER M3 ;
        RECT 6.384 30.392 6.416 30.424 ;
  LAYER M1 ;
        RECT 6.448 27.936 6.48 30.444 ;
  LAYER M3 ;
        RECT 6.448 27.956 6.48 27.988 ;
  LAYER M1 ;
        RECT 6.512 27.936 6.544 30.444 ;
  LAYER M3 ;
        RECT 4.144 30.328 4.176 30.36 ;
  LAYER M2 ;
        RECT 6.512 30.264 6.544 30.296 ;
  LAYER M2 ;
        RECT 4.144 30.2 4.176 30.232 ;
  LAYER M2 ;
        RECT 6.512 30.136 6.544 30.168 ;
  LAYER M2 ;
        RECT 4.144 30.072 4.176 30.104 ;
  LAYER M2 ;
        RECT 6.512 30.008 6.544 30.04 ;
  LAYER M2 ;
        RECT 4.144 29.944 4.176 29.976 ;
  LAYER M2 ;
        RECT 6.512 29.88 6.544 29.912 ;
  LAYER M2 ;
        RECT 4.144 29.816 4.176 29.848 ;
  LAYER M2 ;
        RECT 6.512 29.752 6.544 29.784 ;
  LAYER M2 ;
        RECT 4.144 29.688 4.176 29.72 ;
  LAYER M2 ;
        RECT 6.512 29.624 6.544 29.656 ;
  LAYER M2 ;
        RECT 4.144 29.56 4.176 29.592 ;
  LAYER M2 ;
        RECT 6.512 29.496 6.544 29.528 ;
  LAYER M2 ;
        RECT 4.144 29.432 4.176 29.464 ;
  LAYER M2 ;
        RECT 6.512 29.368 6.544 29.4 ;
  LAYER M2 ;
        RECT 4.144 29.304 4.176 29.336 ;
  LAYER M2 ;
        RECT 6.512 29.24 6.544 29.272 ;
  LAYER M2 ;
        RECT 4.144 29.176 4.176 29.208 ;
  LAYER M2 ;
        RECT 6.512 29.112 6.544 29.144 ;
  LAYER M2 ;
        RECT 4.144 29.048 4.176 29.08 ;
  LAYER M2 ;
        RECT 6.512 28.984 6.544 29.016 ;
  LAYER M2 ;
        RECT 4.144 28.92 4.176 28.952 ;
  LAYER M2 ;
        RECT 6.512 28.856 6.544 28.888 ;
  LAYER M2 ;
        RECT 4.144 28.792 4.176 28.824 ;
  LAYER M2 ;
        RECT 6.512 28.728 6.544 28.76 ;
  LAYER M2 ;
        RECT 4.144 28.664 4.176 28.696 ;
  LAYER M2 ;
        RECT 6.512 28.6 6.544 28.632 ;
  LAYER M2 ;
        RECT 4.144 28.536 4.176 28.568 ;
  LAYER M2 ;
        RECT 6.512 28.472 6.544 28.504 ;
  LAYER M2 ;
        RECT 4.144 28.408 4.176 28.44 ;
  LAYER M2 ;
        RECT 6.512 28.344 6.544 28.376 ;
  LAYER M2 ;
        RECT 4.144 28.28 4.176 28.312 ;
  LAYER M2 ;
        RECT 6.512 28.216 6.544 28.248 ;
  LAYER M2 ;
        RECT 4.144 28.152 4.176 28.184 ;
  LAYER M2 ;
        RECT 6.512 28.088 6.544 28.12 ;
  LAYER M2 ;
        RECT 4.096 27.888 6.592 30.492 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 27.336 ;
  LAYER M3 ;
        RECT 4.144 24.848 4.176 24.88 ;
  LAYER M1 ;
        RECT 4.208 24.828 4.24 27.336 ;
  LAYER M3 ;
        RECT 4.208 27.284 4.24 27.316 ;
  LAYER M1 ;
        RECT 4.272 24.828 4.304 27.336 ;
  LAYER M3 ;
        RECT 4.272 24.848 4.304 24.88 ;
  LAYER M1 ;
        RECT 4.336 24.828 4.368 27.336 ;
  LAYER M3 ;
        RECT 4.336 27.284 4.368 27.316 ;
  LAYER M1 ;
        RECT 4.4 24.828 4.432 27.336 ;
  LAYER M3 ;
        RECT 4.4 24.848 4.432 24.88 ;
  LAYER M1 ;
        RECT 4.464 24.828 4.496 27.336 ;
  LAYER M3 ;
        RECT 4.464 27.284 4.496 27.316 ;
  LAYER M1 ;
        RECT 4.528 24.828 4.56 27.336 ;
  LAYER M3 ;
        RECT 4.528 24.848 4.56 24.88 ;
  LAYER M1 ;
        RECT 4.592 24.828 4.624 27.336 ;
  LAYER M3 ;
        RECT 4.592 27.284 4.624 27.316 ;
  LAYER M1 ;
        RECT 4.656 24.828 4.688 27.336 ;
  LAYER M3 ;
        RECT 4.656 24.848 4.688 24.88 ;
  LAYER M1 ;
        RECT 4.72 24.828 4.752 27.336 ;
  LAYER M3 ;
        RECT 4.72 27.284 4.752 27.316 ;
  LAYER M1 ;
        RECT 4.784 24.828 4.816 27.336 ;
  LAYER M3 ;
        RECT 4.784 24.848 4.816 24.88 ;
  LAYER M1 ;
        RECT 4.848 24.828 4.88 27.336 ;
  LAYER M3 ;
        RECT 4.848 27.284 4.88 27.316 ;
  LAYER M1 ;
        RECT 4.912 24.828 4.944 27.336 ;
  LAYER M3 ;
        RECT 4.912 24.848 4.944 24.88 ;
  LAYER M1 ;
        RECT 4.976 24.828 5.008 27.336 ;
  LAYER M3 ;
        RECT 4.976 27.284 5.008 27.316 ;
  LAYER M1 ;
        RECT 5.04 24.828 5.072 27.336 ;
  LAYER M3 ;
        RECT 5.04 24.848 5.072 24.88 ;
  LAYER M1 ;
        RECT 5.104 24.828 5.136 27.336 ;
  LAYER M3 ;
        RECT 5.104 27.284 5.136 27.316 ;
  LAYER M1 ;
        RECT 5.168 24.828 5.2 27.336 ;
  LAYER M3 ;
        RECT 5.168 24.848 5.2 24.88 ;
  LAYER M1 ;
        RECT 5.232 24.828 5.264 27.336 ;
  LAYER M3 ;
        RECT 5.232 27.284 5.264 27.316 ;
  LAYER M1 ;
        RECT 5.296 24.828 5.328 27.336 ;
  LAYER M3 ;
        RECT 5.296 24.848 5.328 24.88 ;
  LAYER M1 ;
        RECT 5.36 24.828 5.392 27.336 ;
  LAYER M3 ;
        RECT 5.36 27.284 5.392 27.316 ;
  LAYER M1 ;
        RECT 5.424 24.828 5.456 27.336 ;
  LAYER M3 ;
        RECT 5.424 24.848 5.456 24.88 ;
  LAYER M1 ;
        RECT 5.488 24.828 5.52 27.336 ;
  LAYER M3 ;
        RECT 5.488 27.284 5.52 27.316 ;
  LAYER M1 ;
        RECT 5.552 24.828 5.584 27.336 ;
  LAYER M3 ;
        RECT 5.552 24.848 5.584 24.88 ;
  LAYER M1 ;
        RECT 5.616 24.828 5.648 27.336 ;
  LAYER M3 ;
        RECT 5.616 27.284 5.648 27.316 ;
  LAYER M1 ;
        RECT 5.68 24.828 5.712 27.336 ;
  LAYER M3 ;
        RECT 5.68 24.848 5.712 24.88 ;
  LAYER M1 ;
        RECT 5.744 24.828 5.776 27.336 ;
  LAYER M3 ;
        RECT 5.744 27.284 5.776 27.316 ;
  LAYER M1 ;
        RECT 5.808 24.828 5.84 27.336 ;
  LAYER M3 ;
        RECT 5.808 24.848 5.84 24.88 ;
  LAYER M1 ;
        RECT 5.872 24.828 5.904 27.336 ;
  LAYER M3 ;
        RECT 5.872 27.284 5.904 27.316 ;
  LAYER M1 ;
        RECT 5.936 24.828 5.968 27.336 ;
  LAYER M3 ;
        RECT 5.936 24.848 5.968 24.88 ;
  LAYER M1 ;
        RECT 6 24.828 6.032 27.336 ;
  LAYER M3 ;
        RECT 6 27.284 6.032 27.316 ;
  LAYER M1 ;
        RECT 6.064 24.828 6.096 27.336 ;
  LAYER M3 ;
        RECT 6.064 24.848 6.096 24.88 ;
  LAYER M1 ;
        RECT 6.128 24.828 6.16 27.336 ;
  LAYER M3 ;
        RECT 6.128 27.284 6.16 27.316 ;
  LAYER M1 ;
        RECT 6.192 24.828 6.224 27.336 ;
  LAYER M3 ;
        RECT 6.192 24.848 6.224 24.88 ;
  LAYER M1 ;
        RECT 6.256 24.828 6.288 27.336 ;
  LAYER M3 ;
        RECT 6.256 27.284 6.288 27.316 ;
  LAYER M1 ;
        RECT 6.32 24.828 6.352 27.336 ;
  LAYER M3 ;
        RECT 6.32 24.848 6.352 24.88 ;
  LAYER M1 ;
        RECT 6.384 24.828 6.416 27.336 ;
  LAYER M3 ;
        RECT 6.384 27.284 6.416 27.316 ;
  LAYER M1 ;
        RECT 6.448 24.828 6.48 27.336 ;
  LAYER M3 ;
        RECT 6.448 24.848 6.48 24.88 ;
  LAYER M1 ;
        RECT 6.512 24.828 6.544 27.336 ;
  LAYER M3 ;
        RECT 4.144 27.22 4.176 27.252 ;
  LAYER M2 ;
        RECT 6.512 27.156 6.544 27.188 ;
  LAYER M2 ;
        RECT 4.144 27.092 4.176 27.124 ;
  LAYER M2 ;
        RECT 6.512 27.028 6.544 27.06 ;
  LAYER M2 ;
        RECT 4.144 26.964 4.176 26.996 ;
  LAYER M2 ;
        RECT 6.512 26.9 6.544 26.932 ;
  LAYER M2 ;
        RECT 4.144 26.836 4.176 26.868 ;
  LAYER M2 ;
        RECT 6.512 26.772 6.544 26.804 ;
  LAYER M2 ;
        RECT 4.144 26.708 4.176 26.74 ;
  LAYER M2 ;
        RECT 6.512 26.644 6.544 26.676 ;
  LAYER M2 ;
        RECT 4.144 26.58 4.176 26.612 ;
  LAYER M2 ;
        RECT 6.512 26.516 6.544 26.548 ;
  LAYER M2 ;
        RECT 4.144 26.452 4.176 26.484 ;
  LAYER M2 ;
        RECT 6.512 26.388 6.544 26.42 ;
  LAYER M2 ;
        RECT 4.144 26.324 4.176 26.356 ;
  LAYER M2 ;
        RECT 6.512 26.26 6.544 26.292 ;
  LAYER M2 ;
        RECT 4.144 26.196 4.176 26.228 ;
  LAYER M2 ;
        RECT 6.512 26.132 6.544 26.164 ;
  LAYER M2 ;
        RECT 4.144 26.068 4.176 26.1 ;
  LAYER M2 ;
        RECT 6.512 26.004 6.544 26.036 ;
  LAYER M2 ;
        RECT 4.144 25.94 4.176 25.972 ;
  LAYER M2 ;
        RECT 6.512 25.876 6.544 25.908 ;
  LAYER M2 ;
        RECT 4.144 25.812 4.176 25.844 ;
  LAYER M2 ;
        RECT 6.512 25.748 6.544 25.78 ;
  LAYER M2 ;
        RECT 4.144 25.684 4.176 25.716 ;
  LAYER M2 ;
        RECT 6.512 25.62 6.544 25.652 ;
  LAYER M2 ;
        RECT 4.144 25.556 4.176 25.588 ;
  LAYER M2 ;
        RECT 6.512 25.492 6.544 25.524 ;
  LAYER M2 ;
        RECT 4.144 25.428 4.176 25.46 ;
  LAYER M2 ;
        RECT 6.512 25.364 6.544 25.396 ;
  LAYER M2 ;
        RECT 4.144 25.3 4.176 25.332 ;
  LAYER M2 ;
        RECT 6.512 25.236 6.544 25.268 ;
  LAYER M2 ;
        RECT 4.144 25.172 4.176 25.204 ;
  LAYER M2 ;
        RECT 6.512 25.108 6.544 25.14 ;
  LAYER M2 ;
        RECT 4.144 25.044 4.176 25.076 ;
  LAYER M2 ;
        RECT 6.512 24.98 6.544 25.012 ;
  LAYER M2 ;
        RECT 4.096 24.78 6.592 27.384 ;
  LAYER M1 ;
        RECT 4.144 21.72 4.176 24.228 ;
  LAYER M3 ;
        RECT 4.144 21.74 4.176 21.772 ;
  LAYER M1 ;
        RECT 4.208 21.72 4.24 24.228 ;
  LAYER M3 ;
        RECT 4.208 24.176 4.24 24.208 ;
  LAYER M1 ;
        RECT 4.272 21.72 4.304 24.228 ;
  LAYER M3 ;
        RECT 4.272 21.74 4.304 21.772 ;
  LAYER M1 ;
        RECT 4.336 21.72 4.368 24.228 ;
  LAYER M3 ;
        RECT 4.336 24.176 4.368 24.208 ;
  LAYER M1 ;
        RECT 4.4 21.72 4.432 24.228 ;
  LAYER M3 ;
        RECT 4.4 21.74 4.432 21.772 ;
  LAYER M1 ;
        RECT 4.464 21.72 4.496 24.228 ;
  LAYER M3 ;
        RECT 4.464 24.176 4.496 24.208 ;
  LAYER M1 ;
        RECT 4.528 21.72 4.56 24.228 ;
  LAYER M3 ;
        RECT 4.528 21.74 4.56 21.772 ;
  LAYER M1 ;
        RECT 4.592 21.72 4.624 24.228 ;
  LAYER M3 ;
        RECT 4.592 24.176 4.624 24.208 ;
  LAYER M1 ;
        RECT 4.656 21.72 4.688 24.228 ;
  LAYER M3 ;
        RECT 4.656 21.74 4.688 21.772 ;
  LAYER M1 ;
        RECT 4.72 21.72 4.752 24.228 ;
  LAYER M3 ;
        RECT 4.72 24.176 4.752 24.208 ;
  LAYER M1 ;
        RECT 4.784 21.72 4.816 24.228 ;
  LAYER M3 ;
        RECT 4.784 21.74 4.816 21.772 ;
  LAYER M1 ;
        RECT 4.848 21.72 4.88 24.228 ;
  LAYER M3 ;
        RECT 4.848 24.176 4.88 24.208 ;
  LAYER M1 ;
        RECT 4.912 21.72 4.944 24.228 ;
  LAYER M3 ;
        RECT 4.912 21.74 4.944 21.772 ;
  LAYER M1 ;
        RECT 4.976 21.72 5.008 24.228 ;
  LAYER M3 ;
        RECT 4.976 24.176 5.008 24.208 ;
  LAYER M1 ;
        RECT 5.04 21.72 5.072 24.228 ;
  LAYER M3 ;
        RECT 5.04 21.74 5.072 21.772 ;
  LAYER M1 ;
        RECT 5.104 21.72 5.136 24.228 ;
  LAYER M3 ;
        RECT 5.104 24.176 5.136 24.208 ;
  LAYER M1 ;
        RECT 5.168 21.72 5.2 24.228 ;
  LAYER M3 ;
        RECT 5.168 21.74 5.2 21.772 ;
  LAYER M1 ;
        RECT 5.232 21.72 5.264 24.228 ;
  LAYER M3 ;
        RECT 5.232 24.176 5.264 24.208 ;
  LAYER M1 ;
        RECT 5.296 21.72 5.328 24.228 ;
  LAYER M3 ;
        RECT 5.296 21.74 5.328 21.772 ;
  LAYER M1 ;
        RECT 5.36 21.72 5.392 24.228 ;
  LAYER M3 ;
        RECT 5.36 24.176 5.392 24.208 ;
  LAYER M1 ;
        RECT 5.424 21.72 5.456 24.228 ;
  LAYER M3 ;
        RECT 5.424 21.74 5.456 21.772 ;
  LAYER M1 ;
        RECT 5.488 21.72 5.52 24.228 ;
  LAYER M3 ;
        RECT 5.488 24.176 5.52 24.208 ;
  LAYER M1 ;
        RECT 5.552 21.72 5.584 24.228 ;
  LAYER M3 ;
        RECT 5.552 21.74 5.584 21.772 ;
  LAYER M1 ;
        RECT 5.616 21.72 5.648 24.228 ;
  LAYER M3 ;
        RECT 5.616 24.176 5.648 24.208 ;
  LAYER M1 ;
        RECT 5.68 21.72 5.712 24.228 ;
  LAYER M3 ;
        RECT 5.68 21.74 5.712 21.772 ;
  LAYER M1 ;
        RECT 5.744 21.72 5.776 24.228 ;
  LAYER M3 ;
        RECT 5.744 24.176 5.776 24.208 ;
  LAYER M1 ;
        RECT 5.808 21.72 5.84 24.228 ;
  LAYER M3 ;
        RECT 5.808 21.74 5.84 21.772 ;
  LAYER M1 ;
        RECT 5.872 21.72 5.904 24.228 ;
  LAYER M3 ;
        RECT 5.872 24.176 5.904 24.208 ;
  LAYER M1 ;
        RECT 5.936 21.72 5.968 24.228 ;
  LAYER M3 ;
        RECT 5.936 21.74 5.968 21.772 ;
  LAYER M1 ;
        RECT 6 21.72 6.032 24.228 ;
  LAYER M3 ;
        RECT 6 24.176 6.032 24.208 ;
  LAYER M1 ;
        RECT 6.064 21.72 6.096 24.228 ;
  LAYER M3 ;
        RECT 6.064 21.74 6.096 21.772 ;
  LAYER M1 ;
        RECT 6.128 21.72 6.16 24.228 ;
  LAYER M3 ;
        RECT 6.128 24.176 6.16 24.208 ;
  LAYER M1 ;
        RECT 6.192 21.72 6.224 24.228 ;
  LAYER M3 ;
        RECT 6.192 21.74 6.224 21.772 ;
  LAYER M1 ;
        RECT 6.256 21.72 6.288 24.228 ;
  LAYER M3 ;
        RECT 6.256 24.176 6.288 24.208 ;
  LAYER M1 ;
        RECT 6.32 21.72 6.352 24.228 ;
  LAYER M3 ;
        RECT 6.32 21.74 6.352 21.772 ;
  LAYER M1 ;
        RECT 6.384 21.72 6.416 24.228 ;
  LAYER M3 ;
        RECT 6.384 24.176 6.416 24.208 ;
  LAYER M1 ;
        RECT 6.448 21.72 6.48 24.228 ;
  LAYER M3 ;
        RECT 6.448 21.74 6.48 21.772 ;
  LAYER M1 ;
        RECT 6.512 21.72 6.544 24.228 ;
  LAYER M3 ;
        RECT 4.144 24.112 4.176 24.144 ;
  LAYER M2 ;
        RECT 6.512 24.048 6.544 24.08 ;
  LAYER M2 ;
        RECT 4.144 23.984 4.176 24.016 ;
  LAYER M2 ;
        RECT 6.512 23.92 6.544 23.952 ;
  LAYER M2 ;
        RECT 4.144 23.856 4.176 23.888 ;
  LAYER M2 ;
        RECT 6.512 23.792 6.544 23.824 ;
  LAYER M2 ;
        RECT 4.144 23.728 4.176 23.76 ;
  LAYER M2 ;
        RECT 6.512 23.664 6.544 23.696 ;
  LAYER M2 ;
        RECT 4.144 23.6 4.176 23.632 ;
  LAYER M2 ;
        RECT 6.512 23.536 6.544 23.568 ;
  LAYER M2 ;
        RECT 4.144 23.472 4.176 23.504 ;
  LAYER M2 ;
        RECT 6.512 23.408 6.544 23.44 ;
  LAYER M2 ;
        RECT 4.144 23.344 4.176 23.376 ;
  LAYER M2 ;
        RECT 6.512 23.28 6.544 23.312 ;
  LAYER M2 ;
        RECT 4.144 23.216 4.176 23.248 ;
  LAYER M2 ;
        RECT 6.512 23.152 6.544 23.184 ;
  LAYER M2 ;
        RECT 4.144 23.088 4.176 23.12 ;
  LAYER M2 ;
        RECT 6.512 23.024 6.544 23.056 ;
  LAYER M2 ;
        RECT 4.144 22.96 4.176 22.992 ;
  LAYER M2 ;
        RECT 6.512 22.896 6.544 22.928 ;
  LAYER M2 ;
        RECT 4.144 22.832 4.176 22.864 ;
  LAYER M2 ;
        RECT 6.512 22.768 6.544 22.8 ;
  LAYER M2 ;
        RECT 4.144 22.704 4.176 22.736 ;
  LAYER M2 ;
        RECT 6.512 22.64 6.544 22.672 ;
  LAYER M2 ;
        RECT 4.144 22.576 4.176 22.608 ;
  LAYER M2 ;
        RECT 6.512 22.512 6.544 22.544 ;
  LAYER M2 ;
        RECT 4.144 22.448 4.176 22.48 ;
  LAYER M2 ;
        RECT 6.512 22.384 6.544 22.416 ;
  LAYER M2 ;
        RECT 4.144 22.32 4.176 22.352 ;
  LAYER M2 ;
        RECT 6.512 22.256 6.544 22.288 ;
  LAYER M2 ;
        RECT 4.144 22.192 4.176 22.224 ;
  LAYER M2 ;
        RECT 6.512 22.128 6.544 22.16 ;
  LAYER M2 ;
        RECT 4.144 22.064 4.176 22.096 ;
  LAYER M2 ;
        RECT 6.512 22 6.544 22.032 ;
  LAYER M2 ;
        RECT 4.144 21.936 4.176 21.968 ;
  LAYER M2 ;
        RECT 6.512 21.872 6.544 21.904 ;
  LAYER M2 ;
        RECT 4.096 21.672 6.592 24.276 ;
  LAYER M1 ;
        RECT 4.144 18.612 4.176 21.12 ;
  LAYER M3 ;
        RECT 4.144 18.632 4.176 18.664 ;
  LAYER M1 ;
        RECT 4.208 18.612 4.24 21.12 ;
  LAYER M3 ;
        RECT 4.208 21.068 4.24 21.1 ;
  LAYER M1 ;
        RECT 4.272 18.612 4.304 21.12 ;
  LAYER M3 ;
        RECT 4.272 18.632 4.304 18.664 ;
  LAYER M1 ;
        RECT 4.336 18.612 4.368 21.12 ;
  LAYER M3 ;
        RECT 4.336 21.068 4.368 21.1 ;
  LAYER M1 ;
        RECT 4.4 18.612 4.432 21.12 ;
  LAYER M3 ;
        RECT 4.4 18.632 4.432 18.664 ;
  LAYER M1 ;
        RECT 4.464 18.612 4.496 21.12 ;
  LAYER M3 ;
        RECT 4.464 21.068 4.496 21.1 ;
  LAYER M1 ;
        RECT 4.528 18.612 4.56 21.12 ;
  LAYER M3 ;
        RECT 4.528 18.632 4.56 18.664 ;
  LAYER M1 ;
        RECT 4.592 18.612 4.624 21.12 ;
  LAYER M3 ;
        RECT 4.592 21.068 4.624 21.1 ;
  LAYER M1 ;
        RECT 4.656 18.612 4.688 21.12 ;
  LAYER M3 ;
        RECT 4.656 18.632 4.688 18.664 ;
  LAYER M1 ;
        RECT 4.72 18.612 4.752 21.12 ;
  LAYER M3 ;
        RECT 4.72 21.068 4.752 21.1 ;
  LAYER M1 ;
        RECT 4.784 18.612 4.816 21.12 ;
  LAYER M3 ;
        RECT 4.784 18.632 4.816 18.664 ;
  LAYER M1 ;
        RECT 4.848 18.612 4.88 21.12 ;
  LAYER M3 ;
        RECT 4.848 21.068 4.88 21.1 ;
  LAYER M1 ;
        RECT 4.912 18.612 4.944 21.12 ;
  LAYER M3 ;
        RECT 4.912 18.632 4.944 18.664 ;
  LAYER M1 ;
        RECT 4.976 18.612 5.008 21.12 ;
  LAYER M3 ;
        RECT 4.976 21.068 5.008 21.1 ;
  LAYER M1 ;
        RECT 5.04 18.612 5.072 21.12 ;
  LAYER M3 ;
        RECT 5.04 18.632 5.072 18.664 ;
  LAYER M1 ;
        RECT 5.104 18.612 5.136 21.12 ;
  LAYER M3 ;
        RECT 5.104 21.068 5.136 21.1 ;
  LAYER M1 ;
        RECT 5.168 18.612 5.2 21.12 ;
  LAYER M3 ;
        RECT 5.168 18.632 5.2 18.664 ;
  LAYER M1 ;
        RECT 5.232 18.612 5.264 21.12 ;
  LAYER M3 ;
        RECT 5.232 21.068 5.264 21.1 ;
  LAYER M1 ;
        RECT 5.296 18.612 5.328 21.12 ;
  LAYER M3 ;
        RECT 5.296 18.632 5.328 18.664 ;
  LAYER M1 ;
        RECT 5.36 18.612 5.392 21.12 ;
  LAYER M3 ;
        RECT 5.36 21.068 5.392 21.1 ;
  LAYER M1 ;
        RECT 5.424 18.612 5.456 21.12 ;
  LAYER M3 ;
        RECT 5.424 18.632 5.456 18.664 ;
  LAYER M1 ;
        RECT 5.488 18.612 5.52 21.12 ;
  LAYER M3 ;
        RECT 5.488 21.068 5.52 21.1 ;
  LAYER M1 ;
        RECT 5.552 18.612 5.584 21.12 ;
  LAYER M3 ;
        RECT 5.552 18.632 5.584 18.664 ;
  LAYER M1 ;
        RECT 5.616 18.612 5.648 21.12 ;
  LAYER M3 ;
        RECT 5.616 21.068 5.648 21.1 ;
  LAYER M1 ;
        RECT 5.68 18.612 5.712 21.12 ;
  LAYER M3 ;
        RECT 5.68 18.632 5.712 18.664 ;
  LAYER M1 ;
        RECT 5.744 18.612 5.776 21.12 ;
  LAYER M3 ;
        RECT 5.744 21.068 5.776 21.1 ;
  LAYER M1 ;
        RECT 5.808 18.612 5.84 21.12 ;
  LAYER M3 ;
        RECT 5.808 18.632 5.84 18.664 ;
  LAYER M1 ;
        RECT 5.872 18.612 5.904 21.12 ;
  LAYER M3 ;
        RECT 5.872 21.068 5.904 21.1 ;
  LAYER M1 ;
        RECT 5.936 18.612 5.968 21.12 ;
  LAYER M3 ;
        RECT 5.936 18.632 5.968 18.664 ;
  LAYER M1 ;
        RECT 6 18.612 6.032 21.12 ;
  LAYER M3 ;
        RECT 6 21.068 6.032 21.1 ;
  LAYER M1 ;
        RECT 6.064 18.612 6.096 21.12 ;
  LAYER M3 ;
        RECT 6.064 18.632 6.096 18.664 ;
  LAYER M1 ;
        RECT 6.128 18.612 6.16 21.12 ;
  LAYER M3 ;
        RECT 6.128 21.068 6.16 21.1 ;
  LAYER M1 ;
        RECT 6.192 18.612 6.224 21.12 ;
  LAYER M3 ;
        RECT 6.192 18.632 6.224 18.664 ;
  LAYER M1 ;
        RECT 6.256 18.612 6.288 21.12 ;
  LAYER M3 ;
        RECT 6.256 21.068 6.288 21.1 ;
  LAYER M1 ;
        RECT 6.32 18.612 6.352 21.12 ;
  LAYER M3 ;
        RECT 6.32 18.632 6.352 18.664 ;
  LAYER M1 ;
        RECT 6.384 18.612 6.416 21.12 ;
  LAYER M3 ;
        RECT 6.384 21.068 6.416 21.1 ;
  LAYER M1 ;
        RECT 6.448 18.612 6.48 21.12 ;
  LAYER M3 ;
        RECT 6.448 18.632 6.48 18.664 ;
  LAYER M1 ;
        RECT 6.512 18.612 6.544 21.12 ;
  LAYER M3 ;
        RECT 4.144 21.004 4.176 21.036 ;
  LAYER M2 ;
        RECT 6.512 20.94 6.544 20.972 ;
  LAYER M2 ;
        RECT 4.144 20.876 4.176 20.908 ;
  LAYER M2 ;
        RECT 6.512 20.812 6.544 20.844 ;
  LAYER M2 ;
        RECT 4.144 20.748 4.176 20.78 ;
  LAYER M2 ;
        RECT 6.512 20.684 6.544 20.716 ;
  LAYER M2 ;
        RECT 4.144 20.62 4.176 20.652 ;
  LAYER M2 ;
        RECT 6.512 20.556 6.544 20.588 ;
  LAYER M2 ;
        RECT 4.144 20.492 4.176 20.524 ;
  LAYER M2 ;
        RECT 6.512 20.428 6.544 20.46 ;
  LAYER M2 ;
        RECT 4.144 20.364 4.176 20.396 ;
  LAYER M2 ;
        RECT 6.512 20.3 6.544 20.332 ;
  LAYER M2 ;
        RECT 4.144 20.236 4.176 20.268 ;
  LAYER M2 ;
        RECT 6.512 20.172 6.544 20.204 ;
  LAYER M2 ;
        RECT 4.144 20.108 4.176 20.14 ;
  LAYER M2 ;
        RECT 6.512 20.044 6.544 20.076 ;
  LAYER M2 ;
        RECT 4.144 19.98 4.176 20.012 ;
  LAYER M2 ;
        RECT 6.512 19.916 6.544 19.948 ;
  LAYER M2 ;
        RECT 4.144 19.852 4.176 19.884 ;
  LAYER M2 ;
        RECT 6.512 19.788 6.544 19.82 ;
  LAYER M2 ;
        RECT 4.144 19.724 4.176 19.756 ;
  LAYER M2 ;
        RECT 6.512 19.66 6.544 19.692 ;
  LAYER M2 ;
        RECT 4.144 19.596 4.176 19.628 ;
  LAYER M2 ;
        RECT 6.512 19.532 6.544 19.564 ;
  LAYER M2 ;
        RECT 4.144 19.468 4.176 19.5 ;
  LAYER M2 ;
        RECT 6.512 19.404 6.544 19.436 ;
  LAYER M2 ;
        RECT 4.144 19.34 4.176 19.372 ;
  LAYER M2 ;
        RECT 6.512 19.276 6.544 19.308 ;
  LAYER M2 ;
        RECT 4.144 19.212 4.176 19.244 ;
  LAYER M2 ;
        RECT 6.512 19.148 6.544 19.18 ;
  LAYER M2 ;
        RECT 4.144 19.084 4.176 19.116 ;
  LAYER M2 ;
        RECT 6.512 19.02 6.544 19.052 ;
  LAYER M2 ;
        RECT 4.144 18.956 4.176 18.988 ;
  LAYER M2 ;
        RECT 6.512 18.892 6.544 18.924 ;
  LAYER M2 ;
        RECT 4.144 18.828 4.176 18.86 ;
  LAYER M2 ;
        RECT 6.512 18.764 6.544 18.796 ;
  LAYER M2 ;
        RECT 4.096 18.564 6.592 21.168 ;
  LAYER M1 ;
        RECT 4.144 15.504 4.176 18.012 ;
  LAYER M3 ;
        RECT 4.144 15.524 4.176 15.556 ;
  LAYER M1 ;
        RECT 4.208 15.504 4.24 18.012 ;
  LAYER M3 ;
        RECT 4.208 17.96 4.24 17.992 ;
  LAYER M1 ;
        RECT 4.272 15.504 4.304 18.012 ;
  LAYER M3 ;
        RECT 4.272 15.524 4.304 15.556 ;
  LAYER M1 ;
        RECT 4.336 15.504 4.368 18.012 ;
  LAYER M3 ;
        RECT 4.336 17.96 4.368 17.992 ;
  LAYER M1 ;
        RECT 4.4 15.504 4.432 18.012 ;
  LAYER M3 ;
        RECT 4.4 15.524 4.432 15.556 ;
  LAYER M1 ;
        RECT 4.464 15.504 4.496 18.012 ;
  LAYER M3 ;
        RECT 4.464 17.96 4.496 17.992 ;
  LAYER M1 ;
        RECT 4.528 15.504 4.56 18.012 ;
  LAYER M3 ;
        RECT 4.528 15.524 4.56 15.556 ;
  LAYER M1 ;
        RECT 4.592 15.504 4.624 18.012 ;
  LAYER M3 ;
        RECT 4.592 17.96 4.624 17.992 ;
  LAYER M1 ;
        RECT 4.656 15.504 4.688 18.012 ;
  LAYER M3 ;
        RECT 4.656 15.524 4.688 15.556 ;
  LAYER M1 ;
        RECT 4.72 15.504 4.752 18.012 ;
  LAYER M3 ;
        RECT 4.72 17.96 4.752 17.992 ;
  LAYER M1 ;
        RECT 4.784 15.504 4.816 18.012 ;
  LAYER M3 ;
        RECT 4.784 15.524 4.816 15.556 ;
  LAYER M1 ;
        RECT 4.848 15.504 4.88 18.012 ;
  LAYER M3 ;
        RECT 4.848 17.96 4.88 17.992 ;
  LAYER M1 ;
        RECT 4.912 15.504 4.944 18.012 ;
  LAYER M3 ;
        RECT 4.912 15.524 4.944 15.556 ;
  LAYER M1 ;
        RECT 4.976 15.504 5.008 18.012 ;
  LAYER M3 ;
        RECT 4.976 17.96 5.008 17.992 ;
  LAYER M1 ;
        RECT 5.04 15.504 5.072 18.012 ;
  LAYER M3 ;
        RECT 5.04 15.524 5.072 15.556 ;
  LAYER M1 ;
        RECT 5.104 15.504 5.136 18.012 ;
  LAYER M3 ;
        RECT 5.104 17.96 5.136 17.992 ;
  LAYER M1 ;
        RECT 5.168 15.504 5.2 18.012 ;
  LAYER M3 ;
        RECT 5.168 15.524 5.2 15.556 ;
  LAYER M1 ;
        RECT 5.232 15.504 5.264 18.012 ;
  LAYER M3 ;
        RECT 5.232 17.96 5.264 17.992 ;
  LAYER M1 ;
        RECT 5.296 15.504 5.328 18.012 ;
  LAYER M3 ;
        RECT 5.296 15.524 5.328 15.556 ;
  LAYER M1 ;
        RECT 5.36 15.504 5.392 18.012 ;
  LAYER M3 ;
        RECT 5.36 17.96 5.392 17.992 ;
  LAYER M1 ;
        RECT 5.424 15.504 5.456 18.012 ;
  LAYER M3 ;
        RECT 5.424 15.524 5.456 15.556 ;
  LAYER M1 ;
        RECT 5.488 15.504 5.52 18.012 ;
  LAYER M3 ;
        RECT 5.488 17.96 5.52 17.992 ;
  LAYER M1 ;
        RECT 5.552 15.504 5.584 18.012 ;
  LAYER M3 ;
        RECT 5.552 15.524 5.584 15.556 ;
  LAYER M1 ;
        RECT 5.616 15.504 5.648 18.012 ;
  LAYER M3 ;
        RECT 5.616 17.96 5.648 17.992 ;
  LAYER M1 ;
        RECT 5.68 15.504 5.712 18.012 ;
  LAYER M3 ;
        RECT 5.68 15.524 5.712 15.556 ;
  LAYER M1 ;
        RECT 5.744 15.504 5.776 18.012 ;
  LAYER M3 ;
        RECT 5.744 17.96 5.776 17.992 ;
  LAYER M1 ;
        RECT 5.808 15.504 5.84 18.012 ;
  LAYER M3 ;
        RECT 5.808 15.524 5.84 15.556 ;
  LAYER M1 ;
        RECT 5.872 15.504 5.904 18.012 ;
  LAYER M3 ;
        RECT 5.872 17.96 5.904 17.992 ;
  LAYER M1 ;
        RECT 5.936 15.504 5.968 18.012 ;
  LAYER M3 ;
        RECT 5.936 15.524 5.968 15.556 ;
  LAYER M1 ;
        RECT 6 15.504 6.032 18.012 ;
  LAYER M3 ;
        RECT 6 17.96 6.032 17.992 ;
  LAYER M1 ;
        RECT 6.064 15.504 6.096 18.012 ;
  LAYER M3 ;
        RECT 6.064 15.524 6.096 15.556 ;
  LAYER M1 ;
        RECT 6.128 15.504 6.16 18.012 ;
  LAYER M3 ;
        RECT 6.128 17.96 6.16 17.992 ;
  LAYER M1 ;
        RECT 6.192 15.504 6.224 18.012 ;
  LAYER M3 ;
        RECT 6.192 15.524 6.224 15.556 ;
  LAYER M1 ;
        RECT 6.256 15.504 6.288 18.012 ;
  LAYER M3 ;
        RECT 6.256 17.96 6.288 17.992 ;
  LAYER M1 ;
        RECT 6.32 15.504 6.352 18.012 ;
  LAYER M3 ;
        RECT 6.32 15.524 6.352 15.556 ;
  LAYER M1 ;
        RECT 6.384 15.504 6.416 18.012 ;
  LAYER M3 ;
        RECT 6.384 17.96 6.416 17.992 ;
  LAYER M1 ;
        RECT 6.448 15.504 6.48 18.012 ;
  LAYER M3 ;
        RECT 6.448 15.524 6.48 15.556 ;
  LAYER M1 ;
        RECT 6.512 15.504 6.544 18.012 ;
  LAYER M3 ;
        RECT 4.144 17.896 4.176 17.928 ;
  LAYER M2 ;
        RECT 6.512 17.832 6.544 17.864 ;
  LAYER M2 ;
        RECT 4.144 17.768 4.176 17.8 ;
  LAYER M2 ;
        RECT 6.512 17.704 6.544 17.736 ;
  LAYER M2 ;
        RECT 4.144 17.64 4.176 17.672 ;
  LAYER M2 ;
        RECT 6.512 17.576 6.544 17.608 ;
  LAYER M2 ;
        RECT 4.144 17.512 4.176 17.544 ;
  LAYER M2 ;
        RECT 6.512 17.448 6.544 17.48 ;
  LAYER M2 ;
        RECT 4.144 17.384 4.176 17.416 ;
  LAYER M2 ;
        RECT 6.512 17.32 6.544 17.352 ;
  LAYER M2 ;
        RECT 4.144 17.256 4.176 17.288 ;
  LAYER M2 ;
        RECT 6.512 17.192 6.544 17.224 ;
  LAYER M2 ;
        RECT 4.144 17.128 4.176 17.16 ;
  LAYER M2 ;
        RECT 6.512 17.064 6.544 17.096 ;
  LAYER M2 ;
        RECT 4.144 17 4.176 17.032 ;
  LAYER M2 ;
        RECT 6.512 16.936 6.544 16.968 ;
  LAYER M2 ;
        RECT 4.144 16.872 4.176 16.904 ;
  LAYER M2 ;
        RECT 6.512 16.808 6.544 16.84 ;
  LAYER M2 ;
        RECT 4.144 16.744 4.176 16.776 ;
  LAYER M2 ;
        RECT 6.512 16.68 6.544 16.712 ;
  LAYER M2 ;
        RECT 4.144 16.616 4.176 16.648 ;
  LAYER M2 ;
        RECT 6.512 16.552 6.544 16.584 ;
  LAYER M2 ;
        RECT 4.144 16.488 4.176 16.52 ;
  LAYER M2 ;
        RECT 6.512 16.424 6.544 16.456 ;
  LAYER M2 ;
        RECT 4.144 16.36 4.176 16.392 ;
  LAYER M2 ;
        RECT 6.512 16.296 6.544 16.328 ;
  LAYER M2 ;
        RECT 4.144 16.232 4.176 16.264 ;
  LAYER M2 ;
        RECT 6.512 16.168 6.544 16.2 ;
  LAYER M2 ;
        RECT 4.144 16.104 4.176 16.136 ;
  LAYER M2 ;
        RECT 6.512 16.04 6.544 16.072 ;
  LAYER M2 ;
        RECT 4.144 15.976 4.176 16.008 ;
  LAYER M2 ;
        RECT 6.512 15.912 6.544 15.944 ;
  LAYER M2 ;
        RECT 4.144 15.848 4.176 15.88 ;
  LAYER M2 ;
        RECT 6.512 15.784 6.544 15.816 ;
  LAYER M2 ;
        RECT 4.144 15.72 4.176 15.752 ;
  LAYER M2 ;
        RECT 6.512 15.656 6.544 15.688 ;
  LAYER M2 ;
        RECT 4.096 15.456 6.592 18.06 ;
  LAYER M1 ;
        RECT 7.12 27.936 7.152 30.444 ;
  LAYER M3 ;
        RECT 7.12 27.956 7.152 27.988 ;
  LAYER M1 ;
        RECT 7.184 27.936 7.216 30.444 ;
  LAYER M3 ;
        RECT 7.184 30.392 7.216 30.424 ;
  LAYER M1 ;
        RECT 7.248 27.936 7.28 30.444 ;
  LAYER M3 ;
        RECT 7.248 27.956 7.28 27.988 ;
  LAYER M1 ;
        RECT 7.312 27.936 7.344 30.444 ;
  LAYER M3 ;
        RECT 7.312 30.392 7.344 30.424 ;
  LAYER M1 ;
        RECT 7.376 27.936 7.408 30.444 ;
  LAYER M3 ;
        RECT 7.376 27.956 7.408 27.988 ;
  LAYER M1 ;
        RECT 7.44 27.936 7.472 30.444 ;
  LAYER M3 ;
        RECT 7.44 30.392 7.472 30.424 ;
  LAYER M1 ;
        RECT 7.504 27.936 7.536 30.444 ;
  LAYER M3 ;
        RECT 7.504 27.956 7.536 27.988 ;
  LAYER M1 ;
        RECT 7.568 27.936 7.6 30.444 ;
  LAYER M3 ;
        RECT 7.568 30.392 7.6 30.424 ;
  LAYER M1 ;
        RECT 7.632 27.936 7.664 30.444 ;
  LAYER M3 ;
        RECT 7.632 27.956 7.664 27.988 ;
  LAYER M1 ;
        RECT 7.696 27.936 7.728 30.444 ;
  LAYER M3 ;
        RECT 7.696 30.392 7.728 30.424 ;
  LAYER M1 ;
        RECT 7.76 27.936 7.792 30.444 ;
  LAYER M3 ;
        RECT 7.76 27.956 7.792 27.988 ;
  LAYER M1 ;
        RECT 7.824 27.936 7.856 30.444 ;
  LAYER M3 ;
        RECT 7.824 30.392 7.856 30.424 ;
  LAYER M1 ;
        RECT 7.888 27.936 7.92 30.444 ;
  LAYER M3 ;
        RECT 7.888 27.956 7.92 27.988 ;
  LAYER M1 ;
        RECT 7.952 27.936 7.984 30.444 ;
  LAYER M3 ;
        RECT 7.952 30.392 7.984 30.424 ;
  LAYER M1 ;
        RECT 8.016 27.936 8.048 30.444 ;
  LAYER M3 ;
        RECT 8.016 27.956 8.048 27.988 ;
  LAYER M1 ;
        RECT 8.08 27.936 8.112 30.444 ;
  LAYER M3 ;
        RECT 8.08 30.392 8.112 30.424 ;
  LAYER M1 ;
        RECT 8.144 27.936 8.176 30.444 ;
  LAYER M3 ;
        RECT 8.144 27.956 8.176 27.988 ;
  LAYER M1 ;
        RECT 8.208 27.936 8.24 30.444 ;
  LAYER M3 ;
        RECT 8.208 30.392 8.24 30.424 ;
  LAYER M1 ;
        RECT 8.272 27.936 8.304 30.444 ;
  LAYER M3 ;
        RECT 8.272 27.956 8.304 27.988 ;
  LAYER M1 ;
        RECT 8.336 27.936 8.368 30.444 ;
  LAYER M3 ;
        RECT 8.336 30.392 8.368 30.424 ;
  LAYER M1 ;
        RECT 8.4 27.936 8.432 30.444 ;
  LAYER M3 ;
        RECT 8.4 27.956 8.432 27.988 ;
  LAYER M1 ;
        RECT 8.464 27.936 8.496 30.444 ;
  LAYER M3 ;
        RECT 8.464 30.392 8.496 30.424 ;
  LAYER M1 ;
        RECT 8.528 27.936 8.56 30.444 ;
  LAYER M3 ;
        RECT 8.528 27.956 8.56 27.988 ;
  LAYER M1 ;
        RECT 8.592 27.936 8.624 30.444 ;
  LAYER M3 ;
        RECT 8.592 30.392 8.624 30.424 ;
  LAYER M1 ;
        RECT 8.656 27.936 8.688 30.444 ;
  LAYER M3 ;
        RECT 8.656 27.956 8.688 27.988 ;
  LAYER M1 ;
        RECT 8.72 27.936 8.752 30.444 ;
  LAYER M3 ;
        RECT 8.72 30.392 8.752 30.424 ;
  LAYER M1 ;
        RECT 8.784 27.936 8.816 30.444 ;
  LAYER M3 ;
        RECT 8.784 27.956 8.816 27.988 ;
  LAYER M1 ;
        RECT 8.848 27.936 8.88 30.444 ;
  LAYER M3 ;
        RECT 8.848 30.392 8.88 30.424 ;
  LAYER M1 ;
        RECT 8.912 27.936 8.944 30.444 ;
  LAYER M3 ;
        RECT 8.912 27.956 8.944 27.988 ;
  LAYER M1 ;
        RECT 8.976 27.936 9.008 30.444 ;
  LAYER M3 ;
        RECT 8.976 30.392 9.008 30.424 ;
  LAYER M1 ;
        RECT 9.04 27.936 9.072 30.444 ;
  LAYER M3 ;
        RECT 9.04 27.956 9.072 27.988 ;
  LAYER M1 ;
        RECT 9.104 27.936 9.136 30.444 ;
  LAYER M3 ;
        RECT 9.104 30.392 9.136 30.424 ;
  LAYER M1 ;
        RECT 9.168 27.936 9.2 30.444 ;
  LAYER M3 ;
        RECT 9.168 27.956 9.2 27.988 ;
  LAYER M1 ;
        RECT 9.232 27.936 9.264 30.444 ;
  LAYER M3 ;
        RECT 9.232 30.392 9.264 30.424 ;
  LAYER M1 ;
        RECT 9.296 27.936 9.328 30.444 ;
  LAYER M3 ;
        RECT 9.296 27.956 9.328 27.988 ;
  LAYER M1 ;
        RECT 9.36 27.936 9.392 30.444 ;
  LAYER M3 ;
        RECT 9.36 30.392 9.392 30.424 ;
  LAYER M1 ;
        RECT 9.424 27.936 9.456 30.444 ;
  LAYER M3 ;
        RECT 9.424 27.956 9.456 27.988 ;
  LAYER M1 ;
        RECT 9.488 27.936 9.52 30.444 ;
  LAYER M3 ;
        RECT 7.12 30.328 7.152 30.36 ;
  LAYER M2 ;
        RECT 9.488 30.264 9.52 30.296 ;
  LAYER M2 ;
        RECT 7.12 30.2 7.152 30.232 ;
  LAYER M2 ;
        RECT 9.488 30.136 9.52 30.168 ;
  LAYER M2 ;
        RECT 7.12 30.072 7.152 30.104 ;
  LAYER M2 ;
        RECT 9.488 30.008 9.52 30.04 ;
  LAYER M2 ;
        RECT 7.12 29.944 7.152 29.976 ;
  LAYER M2 ;
        RECT 9.488 29.88 9.52 29.912 ;
  LAYER M2 ;
        RECT 7.12 29.816 7.152 29.848 ;
  LAYER M2 ;
        RECT 9.488 29.752 9.52 29.784 ;
  LAYER M2 ;
        RECT 7.12 29.688 7.152 29.72 ;
  LAYER M2 ;
        RECT 9.488 29.624 9.52 29.656 ;
  LAYER M2 ;
        RECT 7.12 29.56 7.152 29.592 ;
  LAYER M2 ;
        RECT 9.488 29.496 9.52 29.528 ;
  LAYER M2 ;
        RECT 7.12 29.432 7.152 29.464 ;
  LAYER M2 ;
        RECT 9.488 29.368 9.52 29.4 ;
  LAYER M2 ;
        RECT 7.12 29.304 7.152 29.336 ;
  LAYER M2 ;
        RECT 9.488 29.24 9.52 29.272 ;
  LAYER M2 ;
        RECT 7.12 29.176 7.152 29.208 ;
  LAYER M2 ;
        RECT 9.488 29.112 9.52 29.144 ;
  LAYER M2 ;
        RECT 7.12 29.048 7.152 29.08 ;
  LAYER M2 ;
        RECT 9.488 28.984 9.52 29.016 ;
  LAYER M2 ;
        RECT 7.12 28.92 7.152 28.952 ;
  LAYER M2 ;
        RECT 9.488 28.856 9.52 28.888 ;
  LAYER M2 ;
        RECT 7.12 28.792 7.152 28.824 ;
  LAYER M2 ;
        RECT 9.488 28.728 9.52 28.76 ;
  LAYER M2 ;
        RECT 7.12 28.664 7.152 28.696 ;
  LAYER M2 ;
        RECT 9.488 28.6 9.52 28.632 ;
  LAYER M2 ;
        RECT 7.12 28.536 7.152 28.568 ;
  LAYER M2 ;
        RECT 9.488 28.472 9.52 28.504 ;
  LAYER M2 ;
        RECT 7.12 28.408 7.152 28.44 ;
  LAYER M2 ;
        RECT 9.488 28.344 9.52 28.376 ;
  LAYER M2 ;
        RECT 7.12 28.28 7.152 28.312 ;
  LAYER M2 ;
        RECT 9.488 28.216 9.52 28.248 ;
  LAYER M2 ;
        RECT 7.12 28.152 7.152 28.184 ;
  LAYER M2 ;
        RECT 9.488 28.088 9.52 28.12 ;
  LAYER M2 ;
        RECT 7.072 27.888 9.568 30.492 ;
  LAYER M1 ;
        RECT 7.12 24.828 7.152 27.336 ;
  LAYER M3 ;
        RECT 7.12 24.848 7.152 24.88 ;
  LAYER M1 ;
        RECT 7.184 24.828 7.216 27.336 ;
  LAYER M3 ;
        RECT 7.184 27.284 7.216 27.316 ;
  LAYER M1 ;
        RECT 7.248 24.828 7.28 27.336 ;
  LAYER M3 ;
        RECT 7.248 24.848 7.28 24.88 ;
  LAYER M1 ;
        RECT 7.312 24.828 7.344 27.336 ;
  LAYER M3 ;
        RECT 7.312 27.284 7.344 27.316 ;
  LAYER M1 ;
        RECT 7.376 24.828 7.408 27.336 ;
  LAYER M3 ;
        RECT 7.376 24.848 7.408 24.88 ;
  LAYER M1 ;
        RECT 7.44 24.828 7.472 27.336 ;
  LAYER M3 ;
        RECT 7.44 27.284 7.472 27.316 ;
  LAYER M1 ;
        RECT 7.504 24.828 7.536 27.336 ;
  LAYER M3 ;
        RECT 7.504 24.848 7.536 24.88 ;
  LAYER M1 ;
        RECT 7.568 24.828 7.6 27.336 ;
  LAYER M3 ;
        RECT 7.568 27.284 7.6 27.316 ;
  LAYER M1 ;
        RECT 7.632 24.828 7.664 27.336 ;
  LAYER M3 ;
        RECT 7.632 24.848 7.664 24.88 ;
  LAYER M1 ;
        RECT 7.696 24.828 7.728 27.336 ;
  LAYER M3 ;
        RECT 7.696 27.284 7.728 27.316 ;
  LAYER M1 ;
        RECT 7.76 24.828 7.792 27.336 ;
  LAYER M3 ;
        RECT 7.76 24.848 7.792 24.88 ;
  LAYER M1 ;
        RECT 7.824 24.828 7.856 27.336 ;
  LAYER M3 ;
        RECT 7.824 27.284 7.856 27.316 ;
  LAYER M1 ;
        RECT 7.888 24.828 7.92 27.336 ;
  LAYER M3 ;
        RECT 7.888 24.848 7.92 24.88 ;
  LAYER M1 ;
        RECT 7.952 24.828 7.984 27.336 ;
  LAYER M3 ;
        RECT 7.952 27.284 7.984 27.316 ;
  LAYER M1 ;
        RECT 8.016 24.828 8.048 27.336 ;
  LAYER M3 ;
        RECT 8.016 24.848 8.048 24.88 ;
  LAYER M1 ;
        RECT 8.08 24.828 8.112 27.336 ;
  LAYER M3 ;
        RECT 8.08 27.284 8.112 27.316 ;
  LAYER M1 ;
        RECT 8.144 24.828 8.176 27.336 ;
  LAYER M3 ;
        RECT 8.144 24.848 8.176 24.88 ;
  LAYER M1 ;
        RECT 8.208 24.828 8.24 27.336 ;
  LAYER M3 ;
        RECT 8.208 27.284 8.24 27.316 ;
  LAYER M1 ;
        RECT 8.272 24.828 8.304 27.336 ;
  LAYER M3 ;
        RECT 8.272 24.848 8.304 24.88 ;
  LAYER M1 ;
        RECT 8.336 24.828 8.368 27.336 ;
  LAYER M3 ;
        RECT 8.336 27.284 8.368 27.316 ;
  LAYER M1 ;
        RECT 8.4 24.828 8.432 27.336 ;
  LAYER M3 ;
        RECT 8.4 24.848 8.432 24.88 ;
  LAYER M1 ;
        RECT 8.464 24.828 8.496 27.336 ;
  LAYER M3 ;
        RECT 8.464 27.284 8.496 27.316 ;
  LAYER M1 ;
        RECT 8.528 24.828 8.56 27.336 ;
  LAYER M3 ;
        RECT 8.528 24.848 8.56 24.88 ;
  LAYER M1 ;
        RECT 8.592 24.828 8.624 27.336 ;
  LAYER M3 ;
        RECT 8.592 27.284 8.624 27.316 ;
  LAYER M1 ;
        RECT 8.656 24.828 8.688 27.336 ;
  LAYER M3 ;
        RECT 8.656 24.848 8.688 24.88 ;
  LAYER M1 ;
        RECT 8.72 24.828 8.752 27.336 ;
  LAYER M3 ;
        RECT 8.72 27.284 8.752 27.316 ;
  LAYER M1 ;
        RECT 8.784 24.828 8.816 27.336 ;
  LAYER M3 ;
        RECT 8.784 24.848 8.816 24.88 ;
  LAYER M1 ;
        RECT 8.848 24.828 8.88 27.336 ;
  LAYER M3 ;
        RECT 8.848 27.284 8.88 27.316 ;
  LAYER M1 ;
        RECT 8.912 24.828 8.944 27.336 ;
  LAYER M3 ;
        RECT 8.912 24.848 8.944 24.88 ;
  LAYER M1 ;
        RECT 8.976 24.828 9.008 27.336 ;
  LAYER M3 ;
        RECT 8.976 27.284 9.008 27.316 ;
  LAYER M1 ;
        RECT 9.04 24.828 9.072 27.336 ;
  LAYER M3 ;
        RECT 9.04 24.848 9.072 24.88 ;
  LAYER M1 ;
        RECT 9.104 24.828 9.136 27.336 ;
  LAYER M3 ;
        RECT 9.104 27.284 9.136 27.316 ;
  LAYER M1 ;
        RECT 9.168 24.828 9.2 27.336 ;
  LAYER M3 ;
        RECT 9.168 24.848 9.2 24.88 ;
  LAYER M1 ;
        RECT 9.232 24.828 9.264 27.336 ;
  LAYER M3 ;
        RECT 9.232 27.284 9.264 27.316 ;
  LAYER M1 ;
        RECT 9.296 24.828 9.328 27.336 ;
  LAYER M3 ;
        RECT 9.296 24.848 9.328 24.88 ;
  LAYER M1 ;
        RECT 9.36 24.828 9.392 27.336 ;
  LAYER M3 ;
        RECT 9.36 27.284 9.392 27.316 ;
  LAYER M1 ;
        RECT 9.424 24.828 9.456 27.336 ;
  LAYER M3 ;
        RECT 9.424 24.848 9.456 24.88 ;
  LAYER M1 ;
        RECT 9.488 24.828 9.52 27.336 ;
  LAYER M3 ;
        RECT 7.12 27.22 7.152 27.252 ;
  LAYER M2 ;
        RECT 9.488 27.156 9.52 27.188 ;
  LAYER M2 ;
        RECT 7.12 27.092 7.152 27.124 ;
  LAYER M2 ;
        RECT 9.488 27.028 9.52 27.06 ;
  LAYER M2 ;
        RECT 7.12 26.964 7.152 26.996 ;
  LAYER M2 ;
        RECT 9.488 26.9 9.52 26.932 ;
  LAYER M2 ;
        RECT 7.12 26.836 7.152 26.868 ;
  LAYER M2 ;
        RECT 9.488 26.772 9.52 26.804 ;
  LAYER M2 ;
        RECT 7.12 26.708 7.152 26.74 ;
  LAYER M2 ;
        RECT 9.488 26.644 9.52 26.676 ;
  LAYER M2 ;
        RECT 7.12 26.58 7.152 26.612 ;
  LAYER M2 ;
        RECT 9.488 26.516 9.52 26.548 ;
  LAYER M2 ;
        RECT 7.12 26.452 7.152 26.484 ;
  LAYER M2 ;
        RECT 9.488 26.388 9.52 26.42 ;
  LAYER M2 ;
        RECT 7.12 26.324 7.152 26.356 ;
  LAYER M2 ;
        RECT 9.488 26.26 9.52 26.292 ;
  LAYER M2 ;
        RECT 7.12 26.196 7.152 26.228 ;
  LAYER M2 ;
        RECT 9.488 26.132 9.52 26.164 ;
  LAYER M2 ;
        RECT 7.12 26.068 7.152 26.1 ;
  LAYER M2 ;
        RECT 9.488 26.004 9.52 26.036 ;
  LAYER M2 ;
        RECT 7.12 25.94 7.152 25.972 ;
  LAYER M2 ;
        RECT 9.488 25.876 9.52 25.908 ;
  LAYER M2 ;
        RECT 7.12 25.812 7.152 25.844 ;
  LAYER M2 ;
        RECT 9.488 25.748 9.52 25.78 ;
  LAYER M2 ;
        RECT 7.12 25.684 7.152 25.716 ;
  LAYER M2 ;
        RECT 9.488 25.62 9.52 25.652 ;
  LAYER M2 ;
        RECT 7.12 25.556 7.152 25.588 ;
  LAYER M2 ;
        RECT 9.488 25.492 9.52 25.524 ;
  LAYER M2 ;
        RECT 7.12 25.428 7.152 25.46 ;
  LAYER M2 ;
        RECT 9.488 25.364 9.52 25.396 ;
  LAYER M2 ;
        RECT 7.12 25.3 7.152 25.332 ;
  LAYER M2 ;
        RECT 9.488 25.236 9.52 25.268 ;
  LAYER M2 ;
        RECT 7.12 25.172 7.152 25.204 ;
  LAYER M2 ;
        RECT 9.488 25.108 9.52 25.14 ;
  LAYER M2 ;
        RECT 7.12 25.044 7.152 25.076 ;
  LAYER M2 ;
        RECT 9.488 24.98 9.52 25.012 ;
  LAYER M2 ;
        RECT 7.072 24.78 9.568 27.384 ;
  LAYER M1 ;
        RECT 7.12 21.72 7.152 24.228 ;
  LAYER M3 ;
        RECT 7.12 21.74 7.152 21.772 ;
  LAYER M1 ;
        RECT 7.184 21.72 7.216 24.228 ;
  LAYER M3 ;
        RECT 7.184 24.176 7.216 24.208 ;
  LAYER M1 ;
        RECT 7.248 21.72 7.28 24.228 ;
  LAYER M3 ;
        RECT 7.248 21.74 7.28 21.772 ;
  LAYER M1 ;
        RECT 7.312 21.72 7.344 24.228 ;
  LAYER M3 ;
        RECT 7.312 24.176 7.344 24.208 ;
  LAYER M1 ;
        RECT 7.376 21.72 7.408 24.228 ;
  LAYER M3 ;
        RECT 7.376 21.74 7.408 21.772 ;
  LAYER M1 ;
        RECT 7.44 21.72 7.472 24.228 ;
  LAYER M3 ;
        RECT 7.44 24.176 7.472 24.208 ;
  LAYER M1 ;
        RECT 7.504 21.72 7.536 24.228 ;
  LAYER M3 ;
        RECT 7.504 21.74 7.536 21.772 ;
  LAYER M1 ;
        RECT 7.568 21.72 7.6 24.228 ;
  LAYER M3 ;
        RECT 7.568 24.176 7.6 24.208 ;
  LAYER M1 ;
        RECT 7.632 21.72 7.664 24.228 ;
  LAYER M3 ;
        RECT 7.632 21.74 7.664 21.772 ;
  LAYER M1 ;
        RECT 7.696 21.72 7.728 24.228 ;
  LAYER M3 ;
        RECT 7.696 24.176 7.728 24.208 ;
  LAYER M1 ;
        RECT 7.76 21.72 7.792 24.228 ;
  LAYER M3 ;
        RECT 7.76 21.74 7.792 21.772 ;
  LAYER M1 ;
        RECT 7.824 21.72 7.856 24.228 ;
  LAYER M3 ;
        RECT 7.824 24.176 7.856 24.208 ;
  LAYER M1 ;
        RECT 7.888 21.72 7.92 24.228 ;
  LAYER M3 ;
        RECT 7.888 21.74 7.92 21.772 ;
  LAYER M1 ;
        RECT 7.952 21.72 7.984 24.228 ;
  LAYER M3 ;
        RECT 7.952 24.176 7.984 24.208 ;
  LAYER M1 ;
        RECT 8.016 21.72 8.048 24.228 ;
  LAYER M3 ;
        RECT 8.016 21.74 8.048 21.772 ;
  LAYER M1 ;
        RECT 8.08 21.72 8.112 24.228 ;
  LAYER M3 ;
        RECT 8.08 24.176 8.112 24.208 ;
  LAYER M1 ;
        RECT 8.144 21.72 8.176 24.228 ;
  LAYER M3 ;
        RECT 8.144 21.74 8.176 21.772 ;
  LAYER M1 ;
        RECT 8.208 21.72 8.24 24.228 ;
  LAYER M3 ;
        RECT 8.208 24.176 8.24 24.208 ;
  LAYER M1 ;
        RECT 8.272 21.72 8.304 24.228 ;
  LAYER M3 ;
        RECT 8.272 21.74 8.304 21.772 ;
  LAYER M1 ;
        RECT 8.336 21.72 8.368 24.228 ;
  LAYER M3 ;
        RECT 8.336 24.176 8.368 24.208 ;
  LAYER M1 ;
        RECT 8.4 21.72 8.432 24.228 ;
  LAYER M3 ;
        RECT 8.4 21.74 8.432 21.772 ;
  LAYER M1 ;
        RECT 8.464 21.72 8.496 24.228 ;
  LAYER M3 ;
        RECT 8.464 24.176 8.496 24.208 ;
  LAYER M1 ;
        RECT 8.528 21.72 8.56 24.228 ;
  LAYER M3 ;
        RECT 8.528 21.74 8.56 21.772 ;
  LAYER M1 ;
        RECT 8.592 21.72 8.624 24.228 ;
  LAYER M3 ;
        RECT 8.592 24.176 8.624 24.208 ;
  LAYER M1 ;
        RECT 8.656 21.72 8.688 24.228 ;
  LAYER M3 ;
        RECT 8.656 21.74 8.688 21.772 ;
  LAYER M1 ;
        RECT 8.72 21.72 8.752 24.228 ;
  LAYER M3 ;
        RECT 8.72 24.176 8.752 24.208 ;
  LAYER M1 ;
        RECT 8.784 21.72 8.816 24.228 ;
  LAYER M3 ;
        RECT 8.784 21.74 8.816 21.772 ;
  LAYER M1 ;
        RECT 8.848 21.72 8.88 24.228 ;
  LAYER M3 ;
        RECT 8.848 24.176 8.88 24.208 ;
  LAYER M1 ;
        RECT 8.912 21.72 8.944 24.228 ;
  LAYER M3 ;
        RECT 8.912 21.74 8.944 21.772 ;
  LAYER M1 ;
        RECT 8.976 21.72 9.008 24.228 ;
  LAYER M3 ;
        RECT 8.976 24.176 9.008 24.208 ;
  LAYER M1 ;
        RECT 9.04 21.72 9.072 24.228 ;
  LAYER M3 ;
        RECT 9.04 21.74 9.072 21.772 ;
  LAYER M1 ;
        RECT 9.104 21.72 9.136 24.228 ;
  LAYER M3 ;
        RECT 9.104 24.176 9.136 24.208 ;
  LAYER M1 ;
        RECT 9.168 21.72 9.2 24.228 ;
  LAYER M3 ;
        RECT 9.168 21.74 9.2 21.772 ;
  LAYER M1 ;
        RECT 9.232 21.72 9.264 24.228 ;
  LAYER M3 ;
        RECT 9.232 24.176 9.264 24.208 ;
  LAYER M1 ;
        RECT 9.296 21.72 9.328 24.228 ;
  LAYER M3 ;
        RECT 9.296 21.74 9.328 21.772 ;
  LAYER M1 ;
        RECT 9.36 21.72 9.392 24.228 ;
  LAYER M3 ;
        RECT 9.36 24.176 9.392 24.208 ;
  LAYER M1 ;
        RECT 9.424 21.72 9.456 24.228 ;
  LAYER M3 ;
        RECT 9.424 21.74 9.456 21.772 ;
  LAYER M1 ;
        RECT 9.488 21.72 9.52 24.228 ;
  LAYER M3 ;
        RECT 7.12 24.112 7.152 24.144 ;
  LAYER M2 ;
        RECT 9.488 24.048 9.52 24.08 ;
  LAYER M2 ;
        RECT 7.12 23.984 7.152 24.016 ;
  LAYER M2 ;
        RECT 9.488 23.92 9.52 23.952 ;
  LAYER M2 ;
        RECT 7.12 23.856 7.152 23.888 ;
  LAYER M2 ;
        RECT 9.488 23.792 9.52 23.824 ;
  LAYER M2 ;
        RECT 7.12 23.728 7.152 23.76 ;
  LAYER M2 ;
        RECT 9.488 23.664 9.52 23.696 ;
  LAYER M2 ;
        RECT 7.12 23.6 7.152 23.632 ;
  LAYER M2 ;
        RECT 9.488 23.536 9.52 23.568 ;
  LAYER M2 ;
        RECT 7.12 23.472 7.152 23.504 ;
  LAYER M2 ;
        RECT 9.488 23.408 9.52 23.44 ;
  LAYER M2 ;
        RECT 7.12 23.344 7.152 23.376 ;
  LAYER M2 ;
        RECT 9.488 23.28 9.52 23.312 ;
  LAYER M2 ;
        RECT 7.12 23.216 7.152 23.248 ;
  LAYER M2 ;
        RECT 9.488 23.152 9.52 23.184 ;
  LAYER M2 ;
        RECT 7.12 23.088 7.152 23.12 ;
  LAYER M2 ;
        RECT 9.488 23.024 9.52 23.056 ;
  LAYER M2 ;
        RECT 7.12 22.96 7.152 22.992 ;
  LAYER M2 ;
        RECT 9.488 22.896 9.52 22.928 ;
  LAYER M2 ;
        RECT 7.12 22.832 7.152 22.864 ;
  LAYER M2 ;
        RECT 9.488 22.768 9.52 22.8 ;
  LAYER M2 ;
        RECT 7.12 22.704 7.152 22.736 ;
  LAYER M2 ;
        RECT 9.488 22.64 9.52 22.672 ;
  LAYER M2 ;
        RECT 7.12 22.576 7.152 22.608 ;
  LAYER M2 ;
        RECT 9.488 22.512 9.52 22.544 ;
  LAYER M2 ;
        RECT 7.12 22.448 7.152 22.48 ;
  LAYER M2 ;
        RECT 9.488 22.384 9.52 22.416 ;
  LAYER M2 ;
        RECT 7.12 22.32 7.152 22.352 ;
  LAYER M2 ;
        RECT 9.488 22.256 9.52 22.288 ;
  LAYER M2 ;
        RECT 7.12 22.192 7.152 22.224 ;
  LAYER M2 ;
        RECT 9.488 22.128 9.52 22.16 ;
  LAYER M2 ;
        RECT 7.12 22.064 7.152 22.096 ;
  LAYER M2 ;
        RECT 9.488 22 9.52 22.032 ;
  LAYER M2 ;
        RECT 7.12 21.936 7.152 21.968 ;
  LAYER M2 ;
        RECT 9.488 21.872 9.52 21.904 ;
  LAYER M2 ;
        RECT 7.072 21.672 9.568 24.276 ;
  LAYER M1 ;
        RECT 7.12 18.612 7.152 21.12 ;
  LAYER M3 ;
        RECT 7.12 18.632 7.152 18.664 ;
  LAYER M1 ;
        RECT 7.184 18.612 7.216 21.12 ;
  LAYER M3 ;
        RECT 7.184 21.068 7.216 21.1 ;
  LAYER M1 ;
        RECT 7.248 18.612 7.28 21.12 ;
  LAYER M3 ;
        RECT 7.248 18.632 7.28 18.664 ;
  LAYER M1 ;
        RECT 7.312 18.612 7.344 21.12 ;
  LAYER M3 ;
        RECT 7.312 21.068 7.344 21.1 ;
  LAYER M1 ;
        RECT 7.376 18.612 7.408 21.12 ;
  LAYER M3 ;
        RECT 7.376 18.632 7.408 18.664 ;
  LAYER M1 ;
        RECT 7.44 18.612 7.472 21.12 ;
  LAYER M3 ;
        RECT 7.44 21.068 7.472 21.1 ;
  LAYER M1 ;
        RECT 7.504 18.612 7.536 21.12 ;
  LAYER M3 ;
        RECT 7.504 18.632 7.536 18.664 ;
  LAYER M1 ;
        RECT 7.568 18.612 7.6 21.12 ;
  LAYER M3 ;
        RECT 7.568 21.068 7.6 21.1 ;
  LAYER M1 ;
        RECT 7.632 18.612 7.664 21.12 ;
  LAYER M3 ;
        RECT 7.632 18.632 7.664 18.664 ;
  LAYER M1 ;
        RECT 7.696 18.612 7.728 21.12 ;
  LAYER M3 ;
        RECT 7.696 21.068 7.728 21.1 ;
  LAYER M1 ;
        RECT 7.76 18.612 7.792 21.12 ;
  LAYER M3 ;
        RECT 7.76 18.632 7.792 18.664 ;
  LAYER M1 ;
        RECT 7.824 18.612 7.856 21.12 ;
  LAYER M3 ;
        RECT 7.824 21.068 7.856 21.1 ;
  LAYER M1 ;
        RECT 7.888 18.612 7.92 21.12 ;
  LAYER M3 ;
        RECT 7.888 18.632 7.92 18.664 ;
  LAYER M1 ;
        RECT 7.952 18.612 7.984 21.12 ;
  LAYER M3 ;
        RECT 7.952 21.068 7.984 21.1 ;
  LAYER M1 ;
        RECT 8.016 18.612 8.048 21.12 ;
  LAYER M3 ;
        RECT 8.016 18.632 8.048 18.664 ;
  LAYER M1 ;
        RECT 8.08 18.612 8.112 21.12 ;
  LAYER M3 ;
        RECT 8.08 21.068 8.112 21.1 ;
  LAYER M1 ;
        RECT 8.144 18.612 8.176 21.12 ;
  LAYER M3 ;
        RECT 8.144 18.632 8.176 18.664 ;
  LAYER M1 ;
        RECT 8.208 18.612 8.24 21.12 ;
  LAYER M3 ;
        RECT 8.208 21.068 8.24 21.1 ;
  LAYER M1 ;
        RECT 8.272 18.612 8.304 21.12 ;
  LAYER M3 ;
        RECT 8.272 18.632 8.304 18.664 ;
  LAYER M1 ;
        RECT 8.336 18.612 8.368 21.12 ;
  LAYER M3 ;
        RECT 8.336 21.068 8.368 21.1 ;
  LAYER M1 ;
        RECT 8.4 18.612 8.432 21.12 ;
  LAYER M3 ;
        RECT 8.4 18.632 8.432 18.664 ;
  LAYER M1 ;
        RECT 8.464 18.612 8.496 21.12 ;
  LAYER M3 ;
        RECT 8.464 21.068 8.496 21.1 ;
  LAYER M1 ;
        RECT 8.528 18.612 8.56 21.12 ;
  LAYER M3 ;
        RECT 8.528 18.632 8.56 18.664 ;
  LAYER M1 ;
        RECT 8.592 18.612 8.624 21.12 ;
  LAYER M3 ;
        RECT 8.592 21.068 8.624 21.1 ;
  LAYER M1 ;
        RECT 8.656 18.612 8.688 21.12 ;
  LAYER M3 ;
        RECT 8.656 18.632 8.688 18.664 ;
  LAYER M1 ;
        RECT 8.72 18.612 8.752 21.12 ;
  LAYER M3 ;
        RECT 8.72 21.068 8.752 21.1 ;
  LAYER M1 ;
        RECT 8.784 18.612 8.816 21.12 ;
  LAYER M3 ;
        RECT 8.784 18.632 8.816 18.664 ;
  LAYER M1 ;
        RECT 8.848 18.612 8.88 21.12 ;
  LAYER M3 ;
        RECT 8.848 21.068 8.88 21.1 ;
  LAYER M1 ;
        RECT 8.912 18.612 8.944 21.12 ;
  LAYER M3 ;
        RECT 8.912 18.632 8.944 18.664 ;
  LAYER M1 ;
        RECT 8.976 18.612 9.008 21.12 ;
  LAYER M3 ;
        RECT 8.976 21.068 9.008 21.1 ;
  LAYER M1 ;
        RECT 9.04 18.612 9.072 21.12 ;
  LAYER M3 ;
        RECT 9.04 18.632 9.072 18.664 ;
  LAYER M1 ;
        RECT 9.104 18.612 9.136 21.12 ;
  LAYER M3 ;
        RECT 9.104 21.068 9.136 21.1 ;
  LAYER M1 ;
        RECT 9.168 18.612 9.2 21.12 ;
  LAYER M3 ;
        RECT 9.168 18.632 9.2 18.664 ;
  LAYER M1 ;
        RECT 9.232 18.612 9.264 21.12 ;
  LAYER M3 ;
        RECT 9.232 21.068 9.264 21.1 ;
  LAYER M1 ;
        RECT 9.296 18.612 9.328 21.12 ;
  LAYER M3 ;
        RECT 9.296 18.632 9.328 18.664 ;
  LAYER M1 ;
        RECT 9.36 18.612 9.392 21.12 ;
  LAYER M3 ;
        RECT 9.36 21.068 9.392 21.1 ;
  LAYER M1 ;
        RECT 9.424 18.612 9.456 21.12 ;
  LAYER M3 ;
        RECT 9.424 18.632 9.456 18.664 ;
  LAYER M1 ;
        RECT 9.488 18.612 9.52 21.12 ;
  LAYER M3 ;
        RECT 7.12 21.004 7.152 21.036 ;
  LAYER M2 ;
        RECT 9.488 20.94 9.52 20.972 ;
  LAYER M2 ;
        RECT 7.12 20.876 7.152 20.908 ;
  LAYER M2 ;
        RECT 9.488 20.812 9.52 20.844 ;
  LAYER M2 ;
        RECT 7.12 20.748 7.152 20.78 ;
  LAYER M2 ;
        RECT 9.488 20.684 9.52 20.716 ;
  LAYER M2 ;
        RECT 7.12 20.62 7.152 20.652 ;
  LAYER M2 ;
        RECT 9.488 20.556 9.52 20.588 ;
  LAYER M2 ;
        RECT 7.12 20.492 7.152 20.524 ;
  LAYER M2 ;
        RECT 9.488 20.428 9.52 20.46 ;
  LAYER M2 ;
        RECT 7.12 20.364 7.152 20.396 ;
  LAYER M2 ;
        RECT 9.488 20.3 9.52 20.332 ;
  LAYER M2 ;
        RECT 7.12 20.236 7.152 20.268 ;
  LAYER M2 ;
        RECT 9.488 20.172 9.52 20.204 ;
  LAYER M2 ;
        RECT 7.12 20.108 7.152 20.14 ;
  LAYER M2 ;
        RECT 9.488 20.044 9.52 20.076 ;
  LAYER M2 ;
        RECT 7.12 19.98 7.152 20.012 ;
  LAYER M2 ;
        RECT 9.488 19.916 9.52 19.948 ;
  LAYER M2 ;
        RECT 7.12 19.852 7.152 19.884 ;
  LAYER M2 ;
        RECT 9.488 19.788 9.52 19.82 ;
  LAYER M2 ;
        RECT 7.12 19.724 7.152 19.756 ;
  LAYER M2 ;
        RECT 9.488 19.66 9.52 19.692 ;
  LAYER M2 ;
        RECT 7.12 19.596 7.152 19.628 ;
  LAYER M2 ;
        RECT 9.488 19.532 9.52 19.564 ;
  LAYER M2 ;
        RECT 7.12 19.468 7.152 19.5 ;
  LAYER M2 ;
        RECT 9.488 19.404 9.52 19.436 ;
  LAYER M2 ;
        RECT 7.12 19.34 7.152 19.372 ;
  LAYER M2 ;
        RECT 9.488 19.276 9.52 19.308 ;
  LAYER M2 ;
        RECT 7.12 19.212 7.152 19.244 ;
  LAYER M2 ;
        RECT 9.488 19.148 9.52 19.18 ;
  LAYER M2 ;
        RECT 7.12 19.084 7.152 19.116 ;
  LAYER M2 ;
        RECT 9.488 19.02 9.52 19.052 ;
  LAYER M2 ;
        RECT 7.12 18.956 7.152 18.988 ;
  LAYER M2 ;
        RECT 9.488 18.892 9.52 18.924 ;
  LAYER M2 ;
        RECT 7.12 18.828 7.152 18.86 ;
  LAYER M2 ;
        RECT 9.488 18.764 9.52 18.796 ;
  LAYER M2 ;
        RECT 7.072 18.564 9.568 21.168 ;
  LAYER M1 ;
        RECT 7.12 15.504 7.152 18.012 ;
  LAYER M3 ;
        RECT 7.12 15.524 7.152 15.556 ;
  LAYER M1 ;
        RECT 7.184 15.504 7.216 18.012 ;
  LAYER M3 ;
        RECT 7.184 17.96 7.216 17.992 ;
  LAYER M1 ;
        RECT 7.248 15.504 7.28 18.012 ;
  LAYER M3 ;
        RECT 7.248 15.524 7.28 15.556 ;
  LAYER M1 ;
        RECT 7.312 15.504 7.344 18.012 ;
  LAYER M3 ;
        RECT 7.312 17.96 7.344 17.992 ;
  LAYER M1 ;
        RECT 7.376 15.504 7.408 18.012 ;
  LAYER M3 ;
        RECT 7.376 15.524 7.408 15.556 ;
  LAYER M1 ;
        RECT 7.44 15.504 7.472 18.012 ;
  LAYER M3 ;
        RECT 7.44 17.96 7.472 17.992 ;
  LAYER M1 ;
        RECT 7.504 15.504 7.536 18.012 ;
  LAYER M3 ;
        RECT 7.504 15.524 7.536 15.556 ;
  LAYER M1 ;
        RECT 7.568 15.504 7.6 18.012 ;
  LAYER M3 ;
        RECT 7.568 17.96 7.6 17.992 ;
  LAYER M1 ;
        RECT 7.632 15.504 7.664 18.012 ;
  LAYER M3 ;
        RECT 7.632 15.524 7.664 15.556 ;
  LAYER M1 ;
        RECT 7.696 15.504 7.728 18.012 ;
  LAYER M3 ;
        RECT 7.696 17.96 7.728 17.992 ;
  LAYER M1 ;
        RECT 7.76 15.504 7.792 18.012 ;
  LAYER M3 ;
        RECT 7.76 15.524 7.792 15.556 ;
  LAYER M1 ;
        RECT 7.824 15.504 7.856 18.012 ;
  LAYER M3 ;
        RECT 7.824 17.96 7.856 17.992 ;
  LAYER M1 ;
        RECT 7.888 15.504 7.92 18.012 ;
  LAYER M3 ;
        RECT 7.888 15.524 7.92 15.556 ;
  LAYER M1 ;
        RECT 7.952 15.504 7.984 18.012 ;
  LAYER M3 ;
        RECT 7.952 17.96 7.984 17.992 ;
  LAYER M1 ;
        RECT 8.016 15.504 8.048 18.012 ;
  LAYER M3 ;
        RECT 8.016 15.524 8.048 15.556 ;
  LAYER M1 ;
        RECT 8.08 15.504 8.112 18.012 ;
  LAYER M3 ;
        RECT 8.08 17.96 8.112 17.992 ;
  LAYER M1 ;
        RECT 8.144 15.504 8.176 18.012 ;
  LAYER M3 ;
        RECT 8.144 15.524 8.176 15.556 ;
  LAYER M1 ;
        RECT 8.208 15.504 8.24 18.012 ;
  LAYER M3 ;
        RECT 8.208 17.96 8.24 17.992 ;
  LAYER M1 ;
        RECT 8.272 15.504 8.304 18.012 ;
  LAYER M3 ;
        RECT 8.272 15.524 8.304 15.556 ;
  LAYER M1 ;
        RECT 8.336 15.504 8.368 18.012 ;
  LAYER M3 ;
        RECT 8.336 17.96 8.368 17.992 ;
  LAYER M1 ;
        RECT 8.4 15.504 8.432 18.012 ;
  LAYER M3 ;
        RECT 8.4 15.524 8.432 15.556 ;
  LAYER M1 ;
        RECT 8.464 15.504 8.496 18.012 ;
  LAYER M3 ;
        RECT 8.464 17.96 8.496 17.992 ;
  LAYER M1 ;
        RECT 8.528 15.504 8.56 18.012 ;
  LAYER M3 ;
        RECT 8.528 15.524 8.56 15.556 ;
  LAYER M1 ;
        RECT 8.592 15.504 8.624 18.012 ;
  LAYER M3 ;
        RECT 8.592 17.96 8.624 17.992 ;
  LAYER M1 ;
        RECT 8.656 15.504 8.688 18.012 ;
  LAYER M3 ;
        RECT 8.656 15.524 8.688 15.556 ;
  LAYER M1 ;
        RECT 8.72 15.504 8.752 18.012 ;
  LAYER M3 ;
        RECT 8.72 17.96 8.752 17.992 ;
  LAYER M1 ;
        RECT 8.784 15.504 8.816 18.012 ;
  LAYER M3 ;
        RECT 8.784 15.524 8.816 15.556 ;
  LAYER M1 ;
        RECT 8.848 15.504 8.88 18.012 ;
  LAYER M3 ;
        RECT 8.848 17.96 8.88 17.992 ;
  LAYER M1 ;
        RECT 8.912 15.504 8.944 18.012 ;
  LAYER M3 ;
        RECT 8.912 15.524 8.944 15.556 ;
  LAYER M1 ;
        RECT 8.976 15.504 9.008 18.012 ;
  LAYER M3 ;
        RECT 8.976 17.96 9.008 17.992 ;
  LAYER M1 ;
        RECT 9.04 15.504 9.072 18.012 ;
  LAYER M3 ;
        RECT 9.04 15.524 9.072 15.556 ;
  LAYER M1 ;
        RECT 9.104 15.504 9.136 18.012 ;
  LAYER M3 ;
        RECT 9.104 17.96 9.136 17.992 ;
  LAYER M1 ;
        RECT 9.168 15.504 9.2 18.012 ;
  LAYER M3 ;
        RECT 9.168 15.524 9.2 15.556 ;
  LAYER M1 ;
        RECT 9.232 15.504 9.264 18.012 ;
  LAYER M3 ;
        RECT 9.232 17.96 9.264 17.992 ;
  LAYER M1 ;
        RECT 9.296 15.504 9.328 18.012 ;
  LAYER M3 ;
        RECT 9.296 15.524 9.328 15.556 ;
  LAYER M1 ;
        RECT 9.36 15.504 9.392 18.012 ;
  LAYER M3 ;
        RECT 9.36 17.96 9.392 17.992 ;
  LAYER M1 ;
        RECT 9.424 15.504 9.456 18.012 ;
  LAYER M3 ;
        RECT 9.424 15.524 9.456 15.556 ;
  LAYER M1 ;
        RECT 9.488 15.504 9.52 18.012 ;
  LAYER M3 ;
        RECT 7.12 17.896 7.152 17.928 ;
  LAYER M2 ;
        RECT 9.488 17.832 9.52 17.864 ;
  LAYER M2 ;
        RECT 7.12 17.768 7.152 17.8 ;
  LAYER M2 ;
        RECT 9.488 17.704 9.52 17.736 ;
  LAYER M2 ;
        RECT 7.12 17.64 7.152 17.672 ;
  LAYER M2 ;
        RECT 9.488 17.576 9.52 17.608 ;
  LAYER M2 ;
        RECT 7.12 17.512 7.152 17.544 ;
  LAYER M2 ;
        RECT 9.488 17.448 9.52 17.48 ;
  LAYER M2 ;
        RECT 7.12 17.384 7.152 17.416 ;
  LAYER M2 ;
        RECT 9.488 17.32 9.52 17.352 ;
  LAYER M2 ;
        RECT 7.12 17.256 7.152 17.288 ;
  LAYER M2 ;
        RECT 9.488 17.192 9.52 17.224 ;
  LAYER M2 ;
        RECT 7.12 17.128 7.152 17.16 ;
  LAYER M2 ;
        RECT 9.488 17.064 9.52 17.096 ;
  LAYER M2 ;
        RECT 7.12 17 7.152 17.032 ;
  LAYER M2 ;
        RECT 9.488 16.936 9.52 16.968 ;
  LAYER M2 ;
        RECT 7.12 16.872 7.152 16.904 ;
  LAYER M2 ;
        RECT 9.488 16.808 9.52 16.84 ;
  LAYER M2 ;
        RECT 7.12 16.744 7.152 16.776 ;
  LAYER M2 ;
        RECT 9.488 16.68 9.52 16.712 ;
  LAYER M2 ;
        RECT 7.12 16.616 7.152 16.648 ;
  LAYER M2 ;
        RECT 9.488 16.552 9.52 16.584 ;
  LAYER M2 ;
        RECT 7.12 16.488 7.152 16.52 ;
  LAYER M2 ;
        RECT 9.488 16.424 9.52 16.456 ;
  LAYER M2 ;
        RECT 7.12 16.36 7.152 16.392 ;
  LAYER M2 ;
        RECT 9.488 16.296 9.52 16.328 ;
  LAYER M2 ;
        RECT 7.12 16.232 7.152 16.264 ;
  LAYER M2 ;
        RECT 9.488 16.168 9.52 16.2 ;
  LAYER M2 ;
        RECT 7.12 16.104 7.152 16.136 ;
  LAYER M2 ;
        RECT 9.488 16.04 9.52 16.072 ;
  LAYER M2 ;
        RECT 7.12 15.976 7.152 16.008 ;
  LAYER M2 ;
        RECT 9.488 15.912 9.52 15.944 ;
  LAYER M2 ;
        RECT 7.12 15.848 7.152 15.88 ;
  LAYER M2 ;
        RECT 9.488 15.784 9.52 15.816 ;
  LAYER M2 ;
        RECT 7.12 15.72 7.152 15.752 ;
  LAYER M2 ;
        RECT 9.488 15.656 9.52 15.688 ;
  LAYER M2 ;
        RECT 7.072 15.456 9.568 18.06 ;
  LAYER M1 ;
        RECT 10.096 27.936 10.128 30.444 ;
  LAYER M3 ;
        RECT 10.096 27.956 10.128 27.988 ;
  LAYER M1 ;
        RECT 10.16 27.936 10.192 30.444 ;
  LAYER M3 ;
        RECT 10.16 30.392 10.192 30.424 ;
  LAYER M1 ;
        RECT 10.224 27.936 10.256 30.444 ;
  LAYER M3 ;
        RECT 10.224 27.956 10.256 27.988 ;
  LAYER M1 ;
        RECT 10.288 27.936 10.32 30.444 ;
  LAYER M3 ;
        RECT 10.288 30.392 10.32 30.424 ;
  LAYER M1 ;
        RECT 10.352 27.936 10.384 30.444 ;
  LAYER M3 ;
        RECT 10.352 27.956 10.384 27.988 ;
  LAYER M1 ;
        RECT 10.416 27.936 10.448 30.444 ;
  LAYER M3 ;
        RECT 10.416 30.392 10.448 30.424 ;
  LAYER M1 ;
        RECT 10.48 27.936 10.512 30.444 ;
  LAYER M3 ;
        RECT 10.48 27.956 10.512 27.988 ;
  LAYER M1 ;
        RECT 10.544 27.936 10.576 30.444 ;
  LAYER M3 ;
        RECT 10.544 30.392 10.576 30.424 ;
  LAYER M1 ;
        RECT 10.608 27.936 10.64 30.444 ;
  LAYER M3 ;
        RECT 10.608 27.956 10.64 27.988 ;
  LAYER M1 ;
        RECT 10.672 27.936 10.704 30.444 ;
  LAYER M3 ;
        RECT 10.672 30.392 10.704 30.424 ;
  LAYER M1 ;
        RECT 10.736 27.936 10.768 30.444 ;
  LAYER M3 ;
        RECT 10.736 27.956 10.768 27.988 ;
  LAYER M1 ;
        RECT 10.8 27.936 10.832 30.444 ;
  LAYER M3 ;
        RECT 10.8 30.392 10.832 30.424 ;
  LAYER M1 ;
        RECT 10.864 27.936 10.896 30.444 ;
  LAYER M3 ;
        RECT 10.864 27.956 10.896 27.988 ;
  LAYER M1 ;
        RECT 10.928 27.936 10.96 30.444 ;
  LAYER M3 ;
        RECT 10.928 30.392 10.96 30.424 ;
  LAYER M1 ;
        RECT 10.992 27.936 11.024 30.444 ;
  LAYER M3 ;
        RECT 10.992 27.956 11.024 27.988 ;
  LAYER M1 ;
        RECT 11.056 27.936 11.088 30.444 ;
  LAYER M3 ;
        RECT 11.056 30.392 11.088 30.424 ;
  LAYER M1 ;
        RECT 11.12 27.936 11.152 30.444 ;
  LAYER M3 ;
        RECT 11.12 27.956 11.152 27.988 ;
  LAYER M1 ;
        RECT 11.184 27.936 11.216 30.444 ;
  LAYER M3 ;
        RECT 11.184 30.392 11.216 30.424 ;
  LAYER M1 ;
        RECT 11.248 27.936 11.28 30.444 ;
  LAYER M3 ;
        RECT 11.248 27.956 11.28 27.988 ;
  LAYER M1 ;
        RECT 11.312 27.936 11.344 30.444 ;
  LAYER M3 ;
        RECT 11.312 30.392 11.344 30.424 ;
  LAYER M1 ;
        RECT 11.376 27.936 11.408 30.444 ;
  LAYER M3 ;
        RECT 11.376 27.956 11.408 27.988 ;
  LAYER M1 ;
        RECT 11.44 27.936 11.472 30.444 ;
  LAYER M3 ;
        RECT 11.44 30.392 11.472 30.424 ;
  LAYER M1 ;
        RECT 11.504 27.936 11.536 30.444 ;
  LAYER M3 ;
        RECT 11.504 27.956 11.536 27.988 ;
  LAYER M1 ;
        RECT 11.568 27.936 11.6 30.444 ;
  LAYER M3 ;
        RECT 11.568 30.392 11.6 30.424 ;
  LAYER M1 ;
        RECT 11.632 27.936 11.664 30.444 ;
  LAYER M3 ;
        RECT 11.632 27.956 11.664 27.988 ;
  LAYER M1 ;
        RECT 11.696 27.936 11.728 30.444 ;
  LAYER M3 ;
        RECT 11.696 30.392 11.728 30.424 ;
  LAYER M1 ;
        RECT 11.76 27.936 11.792 30.444 ;
  LAYER M3 ;
        RECT 11.76 27.956 11.792 27.988 ;
  LAYER M1 ;
        RECT 11.824 27.936 11.856 30.444 ;
  LAYER M3 ;
        RECT 11.824 30.392 11.856 30.424 ;
  LAYER M1 ;
        RECT 11.888 27.936 11.92 30.444 ;
  LAYER M3 ;
        RECT 11.888 27.956 11.92 27.988 ;
  LAYER M1 ;
        RECT 11.952 27.936 11.984 30.444 ;
  LAYER M3 ;
        RECT 11.952 30.392 11.984 30.424 ;
  LAYER M1 ;
        RECT 12.016 27.936 12.048 30.444 ;
  LAYER M3 ;
        RECT 12.016 27.956 12.048 27.988 ;
  LAYER M1 ;
        RECT 12.08 27.936 12.112 30.444 ;
  LAYER M3 ;
        RECT 12.08 30.392 12.112 30.424 ;
  LAYER M1 ;
        RECT 12.144 27.936 12.176 30.444 ;
  LAYER M3 ;
        RECT 12.144 27.956 12.176 27.988 ;
  LAYER M1 ;
        RECT 12.208 27.936 12.24 30.444 ;
  LAYER M3 ;
        RECT 12.208 30.392 12.24 30.424 ;
  LAYER M1 ;
        RECT 12.272 27.936 12.304 30.444 ;
  LAYER M3 ;
        RECT 12.272 27.956 12.304 27.988 ;
  LAYER M1 ;
        RECT 12.336 27.936 12.368 30.444 ;
  LAYER M3 ;
        RECT 12.336 30.392 12.368 30.424 ;
  LAYER M1 ;
        RECT 12.4 27.936 12.432 30.444 ;
  LAYER M3 ;
        RECT 12.4 27.956 12.432 27.988 ;
  LAYER M1 ;
        RECT 12.464 27.936 12.496 30.444 ;
  LAYER M3 ;
        RECT 10.096 30.328 10.128 30.36 ;
  LAYER M2 ;
        RECT 12.464 30.264 12.496 30.296 ;
  LAYER M2 ;
        RECT 10.096 30.2 10.128 30.232 ;
  LAYER M2 ;
        RECT 12.464 30.136 12.496 30.168 ;
  LAYER M2 ;
        RECT 10.096 30.072 10.128 30.104 ;
  LAYER M2 ;
        RECT 12.464 30.008 12.496 30.04 ;
  LAYER M2 ;
        RECT 10.096 29.944 10.128 29.976 ;
  LAYER M2 ;
        RECT 12.464 29.88 12.496 29.912 ;
  LAYER M2 ;
        RECT 10.096 29.816 10.128 29.848 ;
  LAYER M2 ;
        RECT 12.464 29.752 12.496 29.784 ;
  LAYER M2 ;
        RECT 10.096 29.688 10.128 29.72 ;
  LAYER M2 ;
        RECT 12.464 29.624 12.496 29.656 ;
  LAYER M2 ;
        RECT 10.096 29.56 10.128 29.592 ;
  LAYER M2 ;
        RECT 12.464 29.496 12.496 29.528 ;
  LAYER M2 ;
        RECT 10.096 29.432 10.128 29.464 ;
  LAYER M2 ;
        RECT 12.464 29.368 12.496 29.4 ;
  LAYER M2 ;
        RECT 10.096 29.304 10.128 29.336 ;
  LAYER M2 ;
        RECT 12.464 29.24 12.496 29.272 ;
  LAYER M2 ;
        RECT 10.096 29.176 10.128 29.208 ;
  LAYER M2 ;
        RECT 12.464 29.112 12.496 29.144 ;
  LAYER M2 ;
        RECT 10.096 29.048 10.128 29.08 ;
  LAYER M2 ;
        RECT 12.464 28.984 12.496 29.016 ;
  LAYER M2 ;
        RECT 10.096 28.92 10.128 28.952 ;
  LAYER M2 ;
        RECT 12.464 28.856 12.496 28.888 ;
  LAYER M2 ;
        RECT 10.096 28.792 10.128 28.824 ;
  LAYER M2 ;
        RECT 12.464 28.728 12.496 28.76 ;
  LAYER M2 ;
        RECT 10.096 28.664 10.128 28.696 ;
  LAYER M2 ;
        RECT 12.464 28.6 12.496 28.632 ;
  LAYER M2 ;
        RECT 10.096 28.536 10.128 28.568 ;
  LAYER M2 ;
        RECT 12.464 28.472 12.496 28.504 ;
  LAYER M2 ;
        RECT 10.096 28.408 10.128 28.44 ;
  LAYER M2 ;
        RECT 12.464 28.344 12.496 28.376 ;
  LAYER M2 ;
        RECT 10.096 28.28 10.128 28.312 ;
  LAYER M2 ;
        RECT 12.464 28.216 12.496 28.248 ;
  LAYER M2 ;
        RECT 10.096 28.152 10.128 28.184 ;
  LAYER M2 ;
        RECT 12.464 28.088 12.496 28.12 ;
  LAYER M2 ;
        RECT 10.048 27.888 12.544 30.492 ;
  LAYER M1 ;
        RECT 10.096 24.828 10.128 27.336 ;
  LAYER M3 ;
        RECT 10.096 24.848 10.128 24.88 ;
  LAYER M1 ;
        RECT 10.16 24.828 10.192 27.336 ;
  LAYER M3 ;
        RECT 10.16 27.284 10.192 27.316 ;
  LAYER M1 ;
        RECT 10.224 24.828 10.256 27.336 ;
  LAYER M3 ;
        RECT 10.224 24.848 10.256 24.88 ;
  LAYER M1 ;
        RECT 10.288 24.828 10.32 27.336 ;
  LAYER M3 ;
        RECT 10.288 27.284 10.32 27.316 ;
  LAYER M1 ;
        RECT 10.352 24.828 10.384 27.336 ;
  LAYER M3 ;
        RECT 10.352 24.848 10.384 24.88 ;
  LAYER M1 ;
        RECT 10.416 24.828 10.448 27.336 ;
  LAYER M3 ;
        RECT 10.416 27.284 10.448 27.316 ;
  LAYER M1 ;
        RECT 10.48 24.828 10.512 27.336 ;
  LAYER M3 ;
        RECT 10.48 24.848 10.512 24.88 ;
  LAYER M1 ;
        RECT 10.544 24.828 10.576 27.336 ;
  LAYER M3 ;
        RECT 10.544 27.284 10.576 27.316 ;
  LAYER M1 ;
        RECT 10.608 24.828 10.64 27.336 ;
  LAYER M3 ;
        RECT 10.608 24.848 10.64 24.88 ;
  LAYER M1 ;
        RECT 10.672 24.828 10.704 27.336 ;
  LAYER M3 ;
        RECT 10.672 27.284 10.704 27.316 ;
  LAYER M1 ;
        RECT 10.736 24.828 10.768 27.336 ;
  LAYER M3 ;
        RECT 10.736 24.848 10.768 24.88 ;
  LAYER M1 ;
        RECT 10.8 24.828 10.832 27.336 ;
  LAYER M3 ;
        RECT 10.8 27.284 10.832 27.316 ;
  LAYER M1 ;
        RECT 10.864 24.828 10.896 27.336 ;
  LAYER M3 ;
        RECT 10.864 24.848 10.896 24.88 ;
  LAYER M1 ;
        RECT 10.928 24.828 10.96 27.336 ;
  LAYER M3 ;
        RECT 10.928 27.284 10.96 27.316 ;
  LAYER M1 ;
        RECT 10.992 24.828 11.024 27.336 ;
  LAYER M3 ;
        RECT 10.992 24.848 11.024 24.88 ;
  LAYER M1 ;
        RECT 11.056 24.828 11.088 27.336 ;
  LAYER M3 ;
        RECT 11.056 27.284 11.088 27.316 ;
  LAYER M1 ;
        RECT 11.12 24.828 11.152 27.336 ;
  LAYER M3 ;
        RECT 11.12 24.848 11.152 24.88 ;
  LAYER M1 ;
        RECT 11.184 24.828 11.216 27.336 ;
  LAYER M3 ;
        RECT 11.184 27.284 11.216 27.316 ;
  LAYER M1 ;
        RECT 11.248 24.828 11.28 27.336 ;
  LAYER M3 ;
        RECT 11.248 24.848 11.28 24.88 ;
  LAYER M1 ;
        RECT 11.312 24.828 11.344 27.336 ;
  LAYER M3 ;
        RECT 11.312 27.284 11.344 27.316 ;
  LAYER M1 ;
        RECT 11.376 24.828 11.408 27.336 ;
  LAYER M3 ;
        RECT 11.376 24.848 11.408 24.88 ;
  LAYER M1 ;
        RECT 11.44 24.828 11.472 27.336 ;
  LAYER M3 ;
        RECT 11.44 27.284 11.472 27.316 ;
  LAYER M1 ;
        RECT 11.504 24.828 11.536 27.336 ;
  LAYER M3 ;
        RECT 11.504 24.848 11.536 24.88 ;
  LAYER M1 ;
        RECT 11.568 24.828 11.6 27.336 ;
  LAYER M3 ;
        RECT 11.568 27.284 11.6 27.316 ;
  LAYER M1 ;
        RECT 11.632 24.828 11.664 27.336 ;
  LAYER M3 ;
        RECT 11.632 24.848 11.664 24.88 ;
  LAYER M1 ;
        RECT 11.696 24.828 11.728 27.336 ;
  LAYER M3 ;
        RECT 11.696 27.284 11.728 27.316 ;
  LAYER M1 ;
        RECT 11.76 24.828 11.792 27.336 ;
  LAYER M3 ;
        RECT 11.76 24.848 11.792 24.88 ;
  LAYER M1 ;
        RECT 11.824 24.828 11.856 27.336 ;
  LAYER M3 ;
        RECT 11.824 27.284 11.856 27.316 ;
  LAYER M1 ;
        RECT 11.888 24.828 11.92 27.336 ;
  LAYER M3 ;
        RECT 11.888 24.848 11.92 24.88 ;
  LAYER M1 ;
        RECT 11.952 24.828 11.984 27.336 ;
  LAYER M3 ;
        RECT 11.952 27.284 11.984 27.316 ;
  LAYER M1 ;
        RECT 12.016 24.828 12.048 27.336 ;
  LAYER M3 ;
        RECT 12.016 24.848 12.048 24.88 ;
  LAYER M1 ;
        RECT 12.08 24.828 12.112 27.336 ;
  LAYER M3 ;
        RECT 12.08 27.284 12.112 27.316 ;
  LAYER M1 ;
        RECT 12.144 24.828 12.176 27.336 ;
  LAYER M3 ;
        RECT 12.144 24.848 12.176 24.88 ;
  LAYER M1 ;
        RECT 12.208 24.828 12.24 27.336 ;
  LAYER M3 ;
        RECT 12.208 27.284 12.24 27.316 ;
  LAYER M1 ;
        RECT 12.272 24.828 12.304 27.336 ;
  LAYER M3 ;
        RECT 12.272 24.848 12.304 24.88 ;
  LAYER M1 ;
        RECT 12.336 24.828 12.368 27.336 ;
  LAYER M3 ;
        RECT 12.336 27.284 12.368 27.316 ;
  LAYER M1 ;
        RECT 12.4 24.828 12.432 27.336 ;
  LAYER M3 ;
        RECT 12.4 24.848 12.432 24.88 ;
  LAYER M1 ;
        RECT 12.464 24.828 12.496 27.336 ;
  LAYER M3 ;
        RECT 10.096 27.22 10.128 27.252 ;
  LAYER M2 ;
        RECT 12.464 27.156 12.496 27.188 ;
  LAYER M2 ;
        RECT 10.096 27.092 10.128 27.124 ;
  LAYER M2 ;
        RECT 12.464 27.028 12.496 27.06 ;
  LAYER M2 ;
        RECT 10.096 26.964 10.128 26.996 ;
  LAYER M2 ;
        RECT 12.464 26.9 12.496 26.932 ;
  LAYER M2 ;
        RECT 10.096 26.836 10.128 26.868 ;
  LAYER M2 ;
        RECT 12.464 26.772 12.496 26.804 ;
  LAYER M2 ;
        RECT 10.096 26.708 10.128 26.74 ;
  LAYER M2 ;
        RECT 12.464 26.644 12.496 26.676 ;
  LAYER M2 ;
        RECT 10.096 26.58 10.128 26.612 ;
  LAYER M2 ;
        RECT 12.464 26.516 12.496 26.548 ;
  LAYER M2 ;
        RECT 10.096 26.452 10.128 26.484 ;
  LAYER M2 ;
        RECT 12.464 26.388 12.496 26.42 ;
  LAYER M2 ;
        RECT 10.096 26.324 10.128 26.356 ;
  LAYER M2 ;
        RECT 12.464 26.26 12.496 26.292 ;
  LAYER M2 ;
        RECT 10.096 26.196 10.128 26.228 ;
  LAYER M2 ;
        RECT 12.464 26.132 12.496 26.164 ;
  LAYER M2 ;
        RECT 10.096 26.068 10.128 26.1 ;
  LAYER M2 ;
        RECT 12.464 26.004 12.496 26.036 ;
  LAYER M2 ;
        RECT 10.096 25.94 10.128 25.972 ;
  LAYER M2 ;
        RECT 12.464 25.876 12.496 25.908 ;
  LAYER M2 ;
        RECT 10.096 25.812 10.128 25.844 ;
  LAYER M2 ;
        RECT 12.464 25.748 12.496 25.78 ;
  LAYER M2 ;
        RECT 10.096 25.684 10.128 25.716 ;
  LAYER M2 ;
        RECT 12.464 25.62 12.496 25.652 ;
  LAYER M2 ;
        RECT 10.096 25.556 10.128 25.588 ;
  LAYER M2 ;
        RECT 12.464 25.492 12.496 25.524 ;
  LAYER M2 ;
        RECT 10.096 25.428 10.128 25.46 ;
  LAYER M2 ;
        RECT 12.464 25.364 12.496 25.396 ;
  LAYER M2 ;
        RECT 10.096 25.3 10.128 25.332 ;
  LAYER M2 ;
        RECT 12.464 25.236 12.496 25.268 ;
  LAYER M2 ;
        RECT 10.096 25.172 10.128 25.204 ;
  LAYER M2 ;
        RECT 12.464 25.108 12.496 25.14 ;
  LAYER M2 ;
        RECT 10.096 25.044 10.128 25.076 ;
  LAYER M2 ;
        RECT 12.464 24.98 12.496 25.012 ;
  LAYER M2 ;
        RECT 10.048 24.78 12.544 27.384 ;
  LAYER M1 ;
        RECT 10.096 21.72 10.128 24.228 ;
  LAYER M3 ;
        RECT 10.096 21.74 10.128 21.772 ;
  LAYER M1 ;
        RECT 10.16 21.72 10.192 24.228 ;
  LAYER M3 ;
        RECT 10.16 24.176 10.192 24.208 ;
  LAYER M1 ;
        RECT 10.224 21.72 10.256 24.228 ;
  LAYER M3 ;
        RECT 10.224 21.74 10.256 21.772 ;
  LAYER M1 ;
        RECT 10.288 21.72 10.32 24.228 ;
  LAYER M3 ;
        RECT 10.288 24.176 10.32 24.208 ;
  LAYER M1 ;
        RECT 10.352 21.72 10.384 24.228 ;
  LAYER M3 ;
        RECT 10.352 21.74 10.384 21.772 ;
  LAYER M1 ;
        RECT 10.416 21.72 10.448 24.228 ;
  LAYER M3 ;
        RECT 10.416 24.176 10.448 24.208 ;
  LAYER M1 ;
        RECT 10.48 21.72 10.512 24.228 ;
  LAYER M3 ;
        RECT 10.48 21.74 10.512 21.772 ;
  LAYER M1 ;
        RECT 10.544 21.72 10.576 24.228 ;
  LAYER M3 ;
        RECT 10.544 24.176 10.576 24.208 ;
  LAYER M1 ;
        RECT 10.608 21.72 10.64 24.228 ;
  LAYER M3 ;
        RECT 10.608 21.74 10.64 21.772 ;
  LAYER M1 ;
        RECT 10.672 21.72 10.704 24.228 ;
  LAYER M3 ;
        RECT 10.672 24.176 10.704 24.208 ;
  LAYER M1 ;
        RECT 10.736 21.72 10.768 24.228 ;
  LAYER M3 ;
        RECT 10.736 21.74 10.768 21.772 ;
  LAYER M1 ;
        RECT 10.8 21.72 10.832 24.228 ;
  LAYER M3 ;
        RECT 10.8 24.176 10.832 24.208 ;
  LAYER M1 ;
        RECT 10.864 21.72 10.896 24.228 ;
  LAYER M3 ;
        RECT 10.864 21.74 10.896 21.772 ;
  LAYER M1 ;
        RECT 10.928 21.72 10.96 24.228 ;
  LAYER M3 ;
        RECT 10.928 24.176 10.96 24.208 ;
  LAYER M1 ;
        RECT 10.992 21.72 11.024 24.228 ;
  LAYER M3 ;
        RECT 10.992 21.74 11.024 21.772 ;
  LAYER M1 ;
        RECT 11.056 21.72 11.088 24.228 ;
  LAYER M3 ;
        RECT 11.056 24.176 11.088 24.208 ;
  LAYER M1 ;
        RECT 11.12 21.72 11.152 24.228 ;
  LAYER M3 ;
        RECT 11.12 21.74 11.152 21.772 ;
  LAYER M1 ;
        RECT 11.184 21.72 11.216 24.228 ;
  LAYER M3 ;
        RECT 11.184 24.176 11.216 24.208 ;
  LAYER M1 ;
        RECT 11.248 21.72 11.28 24.228 ;
  LAYER M3 ;
        RECT 11.248 21.74 11.28 21.772 ;
  LAYER M1 ;
        RECT 11.312 21.72 11.344 24.228 ;
  LAYER M3 ;
        RECT 11.312 24.176 11.344 24.208 ;
  LAYER M1 ;
        RECT 11.376 21.72 11.408 24.228 ;
  LAYER M3 ;
        RECT 11.376 21.74 11.408 21.772 ;
  LAYER M1 ;
        RECT 11.44 21.72 11.472 24.228 ;
  LAYER M3 ;
        RECT 11.44 24.176 11.472 24.208 ;
  LAYER M1 ;
        RECT 11.504 21.72 11.536 24.228 ;
  LAYER M3 ;
        RECT 11.504 21.74 11.536 21.772 ;
  LAYER M1 ;
        RECT 11.568 21.72 11.6 24.228 ;
  LAYER M3 ;
        RECT 11.568 24.176 11.6 24.208 ;
  LAYER M1 ;
        RECT 11.632 21.72 11.664 24.228 ;
  LAYER M3 ;
        RECT 11.632 21.74 11.664 21.772 ;
  LAYER M1 ;
        RECT 11.696 21.72 11.728 24.228 ;
  LAYER M3 ;
        RECT 11.696 24.176 11.728 24.208 ;
  LAYER M1 ;
        RECT 11.76 21.72 11.792 24.228 ;
  LAYER M3 ;
        RECT 11.76 21.74 11.792 21.772 ;
  LAYER M1 ;
        RECT 11.824 21.72 11.856 24.228 ;
  LAYER M3 ;
        RECT 11.824 24.176 11.856 24.208 ;
  LAYER M1 ;
        RECT 11.888 21.72 11.92 24.228 ;
  LAYER M3 ;
        RECT 11.888 21.74 11.92 21.772 ;
  LAYER M1 ;
        RECT 11.952 21.72 11.984 24.228 ;
  LAYER M3 ;
        RECT 11.952 24.176 11.984 24.208 ;
  LAYER M1 ;
        RECT 12.016 21.72 12.048 24.228 ;
  LAYER M3 ;
        RECT 12.016 21.74 12.048 21.772 ;
  LAYER M1 ;
        RECT 12.08 21.72 12.112 24.228 ;
  LAYER M3 ;
        RECT 12.08 24.176 12.112 24.208 ;
  LAYER M1 ;
        RECT 12.144 21.72 12.176 24.228 ;
  LAYER M3 ;
        RECT 12.144 21.74 12.176 21.772 ;
  LAYER M1 ;
        RECT 12.208 21.72 12.24 24.228 ;
  LAYER M3 ;
        RECT 12.208 24.176 12.24 24.208 ;
  LAYER M1 ;
        RECT 12.272 21.72 12.304 24.228 ;
  LAYER M3 ;
        RECT 12.272 21.74 12.304 21.772 ;
  LAYER M1 ;
        RECT 12.336 21.72 12.368 24.228 ;
  LAYER M3 ;
        RECT 12.336 24.176 12.368 24.208 ;
  LAYER M1 ;
        RECT 12.4 21.72 12.432 24.228 ;
  LAYER M3 ;
        RECT 12.4 21.74 12.432 21.772 ;
  LAYER M1 ;
        RECT 12.464 21.72 12.496 24.228 ;
  LAYER M3 ;
        RECT 10.096 24.112 10.128 24.144 ;
  LAYER M2 ;
        RECT 12.464 24.048 12.496 24.08 ;
  LAYER M2 ;
        RECT 10.096 23.984 10.128 24.016 ;
  LAYER M2 ;
        RECT 12.464 23.92 12.496 23.952 ;
  LAYER M2 ;
        RECT 10.096 23.856 10.128 23.888 ;
  LAYER M2 ;
        RECT 12.464 23.792 12.496 23.824 ;
  LAYER M2 ;
        RECT 10.096 23.728 10.128 23.76 ;
  LAYER M2 ;
        RECT 12.464 23.664 12.496 23.696 ;
  LAYER M2 ;
        RECT 10.096 23.6 10.128 23.632 ;
  LAYER M2 ;
        RECT 12.464 23.536 12.496 23.568 ;
  LAYER M2 ;
        RECT 10.096 23.472 10.128 23.504 ;
  LAYER M2 ;
        RECT 12.464 23.408 12.496 23.44 ;
  LAYER M2 ;
        RECT 10.096 23.344 10.128 23.376 ;
  LAYER M2 ;
        RECT 12.464 23.28 12.496 23.312 ;
  LAYER M2 ;
        RECT 10.096 23.216 10.128 23.248 ;
  LAYER M2 ;
        RECT 12.464 23.152 12.496 23.184 ;
  LAYER M2 ;
        RECT 10.096 23.088 10.128 23.12 ;
  LAYER M2 ;
        RECT 12.464 23.024 12.496 23.056 ;
  LAYER M2 ;
        RECT 10.096 22.96 10.128 22.992 ;
  LAYER M2 ;
        RECT 12.464 22.896 12.496 22.928 ;
  LAYER M2 ;
        RECT 10.096 22.832 10.128 22.864 ;
  LAYER M2 ;
        RECT 12.464 22.768 12.496 22.8 ;
  LAYER M2 ;
        RECT 10.096 22.704 10.128 22.736 ;
  LAYER M2 ;
        RECT 12.464 22.64 12.496 22.672 ;
  LAYER M2 ;
        RECT 10.096 22.576 10.128 22.608 ;
  LAYER M2 ;
        RECT 12.464 22.512 12.496 22.544 ;
  LAYER M2 ;
        RECT 10.096 22.448 10.128 22.48 ;
  LAYER M2 ;
        RECT 12.464 22.384 12.496 22.416 ;
  LAYER M2 ;
        RECT 10.096 22.32 10.128 22.352 ;
  LAYER M2 ;
        RECT 12.464 22.256 12.496 22.288 ;
  LAYER M2 ;
        RECT 10.096 22.192 10.128 22.224 ;
  LAYER M2 ;
        RECT 12.464 22.128 12.496 22.16 ;
  LAYER M2 ;
        RECT 10.096 22.064 10.128 22.096 ;
  LAYER M2 ;
        RECT 12.464 22 12.496 22.032 ;
  LAYER M2 ;
        RECT 10.096 21.936 10.128 21.968 ;
  LAYER M2 ;
        RECT 12.464 21.872 12.496 21.904 ;
  LAYER M2 ;
        RECT 10.048 21.672 12.544 24.276 ;
  LAYER M1 ;
        RECT 10.096 18.612 10.128 21.12 ;
  LAYER M3 ;
        RECT 10.096 18.632 10.128 18.664 ;
  LAYER M1 ;
        RECT 10.16 18.612 10.192 21.12 ;
  LAYER M3 ;
        RECT 10.16 21.068 10.192 21.1 ;
  LAYER M1 ;
        RECT 10.224 18.612 10.256 21.12 ;
  LAYER M3 ;
        RECT 10.224 18.632 10.256 18.664 ;
  LAYER M1 ;
        RECT 10.288 18.612 10.32 21.12 ;
  LAYER M3 ;
        RECT 10.288 21.068 10.32 21.1 ;
  LAYER M1 ;
        RECT 10.352 18.612 10.384 21.12 ;
  LAYER M3 ;
        RECT 10.352 18.632 10.384 18.664 ;
  LAYER M1 ;
        RECT 10.416 18.612 10.448 21.12 ;
  LAYER M3 ;
        RECT 10.416 21.068 10.448 21.1 ;
  LAYER M1 ;
        RECT 10.48 18.612 10.512 21.12 ;
  LAYER M3 ;
        RECT 10.48 18.632 10.512 18.664 ;
  LAYER M1 ;
        RECT 10.544 18.612 10.576 21.12 ;
  LAYER M3 ;
        RECT 10.544 21.068 10.576 21.1 ;
  LAYER M1 ;
        RECT 10.608 18.612 10.64 21.12 ;
  LAYER M3 ;
        RECT 10.608 18.632 10.64 18.664 ;
  LAYER M1 ;
        RECT 10.672 18.612 10.704 21.12 ;
  LAYER M3 ;
        RECT 10.672 21.068 10.704 21.1 ;
  LAYER M1 ;
        RECT 10.736 18.612 10.768 21.12 ;
  LAYER M3 ;
        RECT 10.736 18.632 10.768 18.664 ;
  LAYER M1 ;
        RECT 10.8 18.612 10.832 21.12 ;
  LAYER M3 ;
        RECT 10.8 21.068 10.832 21.1 ;
  LAYER M1 ;
        RECT 10.864 18.612 10.896 21.12 ;
  LAYER M3 ;
        RECT 10.864 18.632 10.896 18.664 ;
  LAYER M1 ;
        RECT 10.928 18.612 10.96 21.12 ;
  LAYER M3 ;
        RECT 10.928 21.068 10.96 21.1 ;
  LAYER M1 ;
        RECT 10.992 18.612 11.024 21.12 ;
  LAYER M3 ;
        RECT 10.992 18.632 11.024 18.664 ;
  LAYER M1 ;
        RECT 11.056 18.612 11.088 21.12 ;
  LAYER M3 ;
        RECT 11.056 21.068 11.088 21.1 ;
  LAYER M1 ;
        RECT 11.12 18.612 11.152 21.12 ;
  LAYER M3 ;
        RECT 11.12 18.632 11.152 18.664 ;
  LAYER M1 ;
        RECT 11.184 18.612 11.216 21.12 ;
  LAYER M3 ;
        RECT 11.184 21.068 11.216 21.1 ;
  LAYER M1 ;
        RECT 11.248 18.612 11.28 21.12 ;
  LAYER M3 ;
        RECT 11.248 18.632 11.28 18.664 ;
  LAYER M1 ;
        RECT 11.312 18.612 11.344 21.12 ;
  LAYER M3 ;
        RECT 11.312 21.068 11.344 21.1 ;
  LAYER M1 ;
        RECT 11.376 18.612 11.408 21.12 ;
  LAYER M3 ;
        RECT 11.376 18.632 11.408 18.664 ;
  LAYER M1 ;
        RECT 11.44 18.612 11.472 21.12 ;
  LAYER M3 ;
        RECT 11.44 21.068 11.472 21.1 ;
  LAYER M1 ;
        RECT 11.504 18.612 11.536 21.12 ;
  LAYER M3 ;
        RECT 11.504 18.632 11.536 18.664 ;
  LAYER M1 ;
        RECT 11.568 18.612 11.6 21.12 ;
  LAYER M3 ;
        RECT 11.568 21.068 11.6 21.1 ;
  LAYER M1 ;
        RECT 11.632 18.612 11.664 21.12 ;
  LAYER M3 ;
        RECT 11.632 18.632 11.664 18.664 ;
  LAYER M1 ;
        RECT 11.696 18.612 11.728 21.12 ;
  LAYER M3 ;
        RECT 11.696 21.068 11.728 21.1 ;
  LAYER M1 ;
        RECT 11.76 18.612 11.792 21.12 ;
  LAYER M3 ;
        RECT 11.76 18.632 11.792 18.664 ;
  LAYER M1 ;
        RECT 11.824 18.612 11.856 21.12 ;
  LAYER M3 ;
        RECT 11.824 21.068 11.856 21.1 ;
  LAYER M1 ;
        RECT 11.888 18.612 11.92 21.12 ;
  LAYER M3 ;
        RECT 11.888 18.632 11.92 18.664 ;
  LAYER M1 ;
        RECT 11.952 18.612 11.984 21.12 ;
  LAYER M3 ;
        RECT 11.952 21.068 11.984 21.1 ;
  LAYER M1 ;
        RECT 12.016 18.612 12.048 21.12 ;
  LAYER M3 ;
        RECT 12.016 18.632 12.048 18.664 ;
  LAYER M1 ;
        RECT 12.08 18.612 12.112 21.12 ;
  LAYER M3 ;
        RECT 12.08 21.068 12.112 21.1 ;
  LAYER M1 ;
        RECT 12.144 18.612 12.176 21.12 ;
  LAYER M3 ;
        RECT 12.144 18.632 12.176 18.664 ;
  LAYER M1 ;
        RECT 12.208 18.612 12.24 21.12 ;
  LAYER M3 ;
        RECT 12.208 21.068 12.24 21.1 ;
  LAYER M1 ;
        RECT 12.272 18.612 12.304 21.12 ;
  LAYER M3 ;
        RECT 12.272 18.632 12.304 18.664 ;
  LAYER M1 ;
        RECT 12.336 18.612 12.368 21.12 ;
  LAYER M3 ;
        RECT 12.336 21.068 12.368 21.1 ;
  LAYER M1 ;
        RECT 12.4 18.612 12.432 21.12 ;
  LAYER M3 ;
        RECT 12.4 18.632 12.432 18.664 ;
  LAYER M1 ;
        RECT 12.464 18.612 12.496 21.12 ;
  LAYER M3 ;
        RECT 10.096 21.004 10.128 21.036 ;
  LAYER M2 ;
        RECT 12.464 20.94 12.496 20.972 ;
  LAYER M2 ;
        RECT 10.096 20.876 10.128 20.908 ;
  LAYER M2 ;
        RECT 12.464 20.812 12.496 20.844 ;
  LAYER M2 ;
        RECT 10.096 20.748 10.128 20.78 ;
  LAYER M2 ;
        RECT 12.464 20.684 12.496 20.716 ;
  LAYER M2 ;
        RECT 10.096 20.62 10.128 20.652 ;
  LAYER M2 ;
        RECT 12.464 20.556 12.496 20.588 ;
  LAYER M2 ;
        RECT 10.096 20.492 10.128 20.524 ;
  LAYER M2 ;
        RECT 12.464 20.428 12.496 20.46 ;
  LAYER M2 ;
        RECT 10.096 20.364 10.128 20.396 ;
  LAYER M2 ;
        RECT 12.464 20.3 12.496 20.332 ;
  LAYER M2 ;
        RECT 10.096 20.236 10.128 20.268 ;
  LAYER M2 ;
        RECT 12.464 20.172 12.496 20.204 ;
  LAYER M2 ;
        RECT 10.096 20.108 10.128 20.14 ;
  LAYER M2 ;
        RECT 12.464 20.044 12.496 20.076 ;
  LAYER M2 ;
        RECT 10.096 19.98 10.128 20.012 ;
  LAYER M2 ;
        RECT 12.464 19.916 12.496 19.948 ;
  LAYER M2 ;
        RECT 10.096 19.852 10.128 19.884 ;
  LAYER M2 ;
        RECT 12.464 19.788 12.496 19.82 ;
  LAYER M2 ;
        RECT 10.096 19.724 10.128 19.756 ;
  LAYER M2 ;
        RECT 12.464 19.66 12.496 19.692 ;
  LAYER M2 ;
        RECT 10.096 19.596 10.128 19.628 ;
  LAYER M2 ;
        RECT 12.464 19.532 12.496 19.564 ;
  LAYER M2 ;
        RECT 10.096 19.468 10.128 19.5 ;
  LAYER M2 ;
        RECT 12.464 19.404 12.496 19.436 ;
  LAYER M2 ;
        RECT 10.096 19.34 10.128 19.372 ;
  LAYER M2 ;
        RECT 12.464 19.276 12.496 19.308 ;
  LAYER M2 ;
        RECT 10.096 19.212 10.128 19.244 ;
  LAYER M2 ;
        RECT 12.464 19.148 12.496 19.18 ;
  LAYER M2 ;
        RECT 10.096 19.084 10.128 19.116 ;
  LAYER M2 ;
        RECT 12.464 19.02 12.496 19.052 ;
  LAYER M2 ;
        RECT 10.096 18.956 10.128 18.988 ;
  LAYER M2 ;
        RECT 12.464 18.892 12.496 18.924 ;
  LAYER M2 ;
        RECT 10.096 18.828 10.128 18.86 ;
  LAYER M2 ;
        RECT 12.464 18.764 12.496 18.796 ;
  LAYER M2 ;
        RECT 10.048 18.564 12.544 21.168 ;
  LAYER M1 ;
        RECT 10.096 15.504 10.128 18.012 ;
  LAYER M3 ;
        RECT 10.096 15.524 10.128 15.556 ;
  LAYER M1 ;
        RECT 10.16 15.504 10.192 18.012 ;
  LAYER M3 ;
        RECT 10.16 17.96 10.192 17.992 ;
  LAYER M1 ;
        RECT 10.224 15.504 10.256 18.012 ;
  LAYER M3 ;
        RECT 10.224 15.524 10.256 15.556 ;
  LAYER M1 ;
        RECT 10.288 15.504 10.32 18.012 ;
  LAYER M3 ;
        RECT 10.288 17.96 10.32 17.992 ;
  LAYER M1 ;
        RECT 10.352 15.504 10.384 18.012 ;
  LAYER M3 ;
        RECT 10.352 15.524 10.384 15.556 ;
  LAYER M1 ;
        RECT 10.416 15.504 10.448 18.012 ;
  LAYER M3 ;
        RECT 10.416 17.96 10.448 17.992 ;
  LAYER M1 ;
        RECT 10.48 15.504 10.512 18.012 ;
  LAYER M3 ;
        RECT 10.48 15.524 10.512 15.556 ;
  LAYER M1 ;
        RECT 10.544 15.504 10.576 18.012 ;
  LAYER M3 ;
        RECT 10.544 17.96 10.576 17.992 ;
  LAYER M1 ;
        RECT 10.608 15.504 10.64 18.012 ;
  LAYER M3 ;
        RECT 10.608 15.524 10.64 15.556 ;
  LAYER M1 ;
        RECT 10.672 15.504 10.704 18.012 ;
  LAYER M3 ;
        RECT 10.672 17.96 10.704 17.992 ;
  LAYER M1 ;
        RECT 10.736 15.504 10.768 18.012 ;
  LAYER M3 ;
        RECT 10.736 15.524 10.768 15.556 ;
  LAYER M1 ;
        RECT 10.8 15.504 10.832 18.012 ;
  LAYER M3 ;
        RECT 10.8 17.96 10.832 17.992 ;
  LAYER M1 ;
        RECT 10.864 15.504 10.896 18.012 ;
  LAYER M3 ;
        RECT 10.864 15.524 10.896 15.556 ;
  LAYER M1 ;
        RECT 10.928 15.504 10.96 18.012 ;
  LAYER M3 ;
        RECT 10.928 17.96 10.96 17.992 ;
  LAYER M1 ;
        RECT 10.992 15.504 11.024 18.012 ;
  LAYER M3 ;
        RECT 10.992 15.524 11.024 15.556 ;
  LAYER M1 ;
        RECT 11.056 15.504 11.088 18.012 ;
  LAYER M3 ;
        RECT 11.056 17.96 11.088 17.992 ;
  LAYER M1 ;
        RECT 11.12 15.504 11.152 18.012 ;
  LAYER M3 ;
        RECT 11.12 15.524 11.152 15.556 ;
  LAYER M1 ;
        RECT 11.184 15.504 11.216 18.012 ;
  LAYER M3 ;
        RECT 11.184 17.96 11.216 17.992 ;
  LAYER M1 ;
        RECT 11.248 15.504 11.28 18.012 ;
  LAYER M3 ;
        RECT 11.248 15.524 11.28 15.556 ;
  LAYER M1 ;
        RECT 11.312 15.504 11.344 18.012 ;
  LAYER M3 ;
        RECT 11.312 17.96 11.344 17.992 ;
  LAYER M1 ;
        RECT 11.376 15.504 11.408 18.012 ;
  LAYER M3 ;
        RECT 11.376 15.524 11.408 15.556 ;
  LAYER M1 ;
        RECT 11.44 15.504 11.472 18.012 ;
  LAYER M3 ;
        RECT 11.44 17.96 11.472 17.992 ;
  LAYER M1 ;
        RECT 11.504 15.504 11.536 18.012 ;
  LAYER M3 ;
        RECT 11.504 15.524 11.536 15.556 ;
  LAYER M1 ;
        RECT 11.568 15.504 11.6 18.012 ;
  LAYER M3 ;
        RECT 11.568 17.96 11.6 17.992 ;
  LAYER M1 ;
        RECT 11.632 15.504 11.664 18.012 ;
  LAYER M3 ;
        RECT 11.632 15.524 11.664 15.556 ;
  LAYER M1 ;
        RECT 11.696 15.504 11.728 18.012 ;
  LAYER M3 ;
        RECT 11.696 17.96 11.728 17.992 ;
  LAYER M1 ;
        RECT 11.76 15.504 11.792 18.012 ;
  LAYER M3 ;
        RECT 11.76 15.524 11.792 15.556 ;
  LAYER M1 ;
        RECT 11.824 15.504 11.856 18.012 ;
  LAYER M3 ;
        RECT 11.824 17.96 11.856 17.992 ;
  LAYER M1 ;
        RECT 11.888 15.504 11.92 18.012 ;
  LAYER M3 ;
        RECT 11.888 15.524 11.92 15.556 ;
  LAYER M1 ;
        RECT 11.952 15.504 11.984 18.012 ;
  LAYER M3 ;
        RECT 11.952 17.96 11.984 17.992 ;
  LAYER M1 ;
        RECT 12.016 15.504 12.048 18.012 ;
  LAYER M3 ;
        RECT 12.016 15.524 12.048 15.556 ;
  LAYER M1 ;
        RECT 12.08 15.504 12.112 18.012 ;
  LAYER M3 ;
        RECT 12.08 17.96 12.112 17.992 ;
  LAYER M1 ;
        RECT 12.144 15.504 12.176 18.012 ;
  LAYER M3 ;
        RECT 12.144 15.524 12.176 15.556 ;
  LAYER M1 ;
        RECT 12.208 15.504 12.24 18.012 ;
  LAYER M3 ;
        RECT 12.208 17.96 12.24 17.992 ;
  LAYER M1 ;
        RECT 12.272 15.504 12.304 18.012 ;
  LAYER M3 ;
        RECT 12.272 15.524 12.304 15.556 ;
  LAYER M1 ;
        RECT 12.336 15.504 12.368 18.012 ;
  LAYER M3 ;
        RECT 12.336 17.96 12.368 17.992 ;
  LAYER M1 ;
        RECT 12.4 15.504 12.432 18.012 ;
  LAYER M3 ;
        RECT 12.4 15.524 12.432 15.556 ;
  LAYER M1 ;
        RECT 12.464 15.504 12.496 18.012 ;
  LAYER M3 ;
        RECT 10.096 17.896 10.128 17.928 ;
  LAYER M2 ;
        RECT 12.464 17.832 12.496 17.864 ;
  LAYER M2 ;
        RECT 10.096 17.768 10.128 17.8 ;
  LAYER M2 ;
        RECT 12.464 17.704 12.496 17.736 ;
  LAYER M2 ;
        RECT 10.096 17.64 10.128 17.672 ;
  LAYER M2 ;
        RECT 12.464 17.576 12.496 17.608 ;
  LAYER M2 ;
        RECT 10.096 17.512 10.128 17.544 ;
  LAYER M2 ;
        RECT 12.464 17.448 12.496 17.48 ;
  LAYER M2 ;
        RECT 10.096 17.384 10.128 17.416 ;
  LAYER M2 ;
        RECT 12.464 17.32 12.496 17.352 ;
  LAYER M2 ;
        RECT 10.096 17.256 10.128 17.288 ;
  LAYER M2 ;
        RECT 12.464 17.192 12.496 17.224 ;
  LAYER M2 ;
        RECT 10.096 17.128 10.128 17.16 ;
  LAYER M2 ;
        RECT 12.464 17.064 12.496 17.096 ;
  LAYER M2 ;
        RECT 10.096 17 10.128 17.032 ;
  LAYER M2 ;
        RECT 12.464 16.936 12.496 16.968 ;
  LAYER M2 ;
        RECT 10.096 16.872 10.128 16.904 ;
  LAYER M2 ;
        RECT 12.464 16.808 12.496 16.84 ;
  LAYER M2 ;
        RECT 10.096 16.744 10.128 16.776 ;
  LAYER M2 ;
        RECT 12.464 16.68 12.496 16.712 ;
  LAYER M2 ;
        RECT 10.096 16.616 10.128 16.648 ;
  LAYER M2 ;
        RECT 12.464 16.552 12.496 16.584 ;
  LAYER M2 ;
        RECT 10.096 16.488 10.128 16.52 ;
  LAYER M2 ;
        RECT 12.464 16.424 12.496 16.456 ;
  LAYER M2 ;
        RECT 10.096 16.36 10.128 16.392 ;
  LAYER M2 ;
        RECT 12.464 16.296 12.496 16.328 ;
  LAYER M2 ;
        RECT 10.096 16.232 10.128 16.264 ;
  LAYER M2 ;
        RECT 12.464 16.168 12.496 16.2 ;
  LAYER M2 ;
        RECT 10.096 16.104 10.128 16.136 ;
  LAYER M2 ;
        RECT 12.464 16.04 12.496 16.072 ;
  LAYER M2 ;
        RECT 10.096 15.976 10.128 16.008 ;
  LAYER M2 ;
        RECT 12.464 15.912 12.496 15.944 ;
  LAYER M2 ;
        RECT 10.096 15.848 10.128 15.88 ;
  LAYER M2 ;
        RECT 12.464 15.784 12.496 15.816 ;
  LAYER M2 ;
        RECT 10.096 15.72 10.128 15.752 ;
  LAYER M2 ;
        RECT 12.464 15.656 12.496 15.688 ;
  LAYER M2 ;
        RECT 10.048 15.456 12.544 18.06 ;
  LAYER M1 ;
        RECT 13.072 27.936 13.104 30.444 ;
  LAYER M3 ;
        RECT 13.072 27.956 13.104 27.988 ;
  LAYER M1 ;
        RECT 13.136 27.936 13.168 30.444 ;
  LAYER M3 ;
        RECT 13.136 30.392 13.168 30.424 ;
  LAYER M1 ;
        RECT 13.2 27.936 13.232 30.444 ;
  LAYER M3 ;
        RECT 13.2 27.956 13.232 27.988 ;
  LAYER M1 ;
        RECT 13.264 27.936 13.296 30.444 ;
  LAYER M3 ;
        RECT 13.264 30.392 13.296 30.424 ;
  LAYER M1 ;
        RECT 13.328 27.936 13.36 30.444 ;
  LAYER M3 ;
        RECT 13.328 27.956 13.36 27.988 ;
  LAYER M1 ;
        RECT 13.392 27.936 13.424 30.444 ;
  LAYER M3 ;
        RECT 13.392 30.392 13.424 30.424 ;
  LAYER M1 ;
        RECT 13.456 27.936 13.488 30.444 ;
  LAYER M3 ;
        RECT 13.456 27.956 13.488 27.988 ;
  LAYER M1 ;
        RECT 13.52 27.936 13.552 30.444 ;
  LAYER M3 ;
        RECT 13.52 30.392 13.552 30.424 ;
  LAYER M1 ;
        RECT 13.584 27.936 13.616 30.444 ;
  LAYER M3 ;
        RECT 13.584 27.956 13.616 27.988 ;
  LAYER M1 ;
        RECT 13.648 27.936 13.68 30.444 ;
  LAYER M3 ;
        RECT 13.648 30.392 13.68 30.424 ;
  LAYER M1 ;
        RECT 13.712 27.936 13.744 30.444 ;
  LAYER M3 ;
        RECT 13.712 27.956 13.744 27.988 ;
  LAYER M1 ;
        RECT 13.776 27.936 13.808 30.444 ;
  LAYER M3 ;
        RECT 13.776 30.392 13.808 30.424 ;
  LAYER M1 ;
        RECT 13.84 27.936 13.872 30.444 ;
  LAYER M3 ;
        RECT 13.84 27.956 13.872 27.988 ;
  LAYER M1 ;
        RECT 13.904 27.936 13.936 30.444 ;
  LAYER M3 ;
        RECT 13.904 30.392 13.936 30.424 ;
  LAYER M1 ;
        RECT 13.968 27.936 14 30.444 ;
  LAYER M3 ;
        RECT 13.968 27.956 14 27.988 ;
  LAYER M1 ;
        RECT 14.032 27.936 14.064 30.444 ;
  LAYER M3 ;
        RECT 14.032 30.392 14.064 30.424 ;
  LAYER M1 ;
        RECT 14.096 27.936 14.128 30.444 ;
  LAYER M3 ;
        RECT 14.096 27.956 14.128 27.988 ;
  LAYER M1 ;
        RECT 14.16 27.936 14.192 30.444 ;
  LAYER M3 ;
        RECT 14.16 30.392 14.192 30.424 ;
  LAYER M1 ;
        RECT 14.224 27.936 14.256 30.444 ;
  LAYER M3 ;
        RECT 14.224 27.956 14.256 27.988 ;
  LAYER M1 ;
        RECT 14.288 27.936 14.32 30.444 ;
  LAYER M3 ;
        RECT 14.288 30.392 14.32 30.424 ;
  LAYER M1 ;
        RECT 14.352 27.936 14.384 30.444 ;
  LAYER M3 ;
        RECT 14.352 27.956 14.384 27.988 ;
  LAYER M1 ;
        RECT 14.416 27.936 14.448 30.444 ;
  LAYER M3 ;
        RECT 14.416 30.392 14.448 30.424 ;
  LAYER M1 ;
        RECT 14.48 27.936 14.512 30.444 ;
  LAYER M3 ;
        RECT 14.48 27.956 14.512 27.988 ;
  LAYER M1 ;
        RECT 14.544 27.936 14.576 30.444 ;
  LAYER M3 ;
        RECT 14.544 30.392 14.576 30.424 ;
  LAYER M1 ;
        RECT 14.608 27.936 14.64 30.444 ;
  LAYER M3 ;
        RECT 14.608 27.956 14.64 27.988 ;
  LAYER M1 ;
        RECT 14.672 27.936 14.704 30.444 ;
  LAYER M3 ;
        RECT 14.672 30.392 14.704 30.424 ;
  LAYER M1 ;
        RECT 14.736 27.936 14.768 30.444 ;
  LAYER M3 ;
        RECT 14.736 27.956 14.768 27.988 ;
  LAYER M1 ;
        RECT 14.8 27.936 14.832 30.444 ;
  LAYER M3 ;
        RECT 14.8 30.392 14.832 30.424 ;
  LAYER M1 ;
        RECT 14.864 27.936 14.896 30.444 ;
  LAYER M3 ;
        RECT 14.864 27.956 14.896 27.988 ;
  LAYER M1 ;
        RECT 14.928 27.936 14.96 30.444 ;
  LAYER M3 ;
        RECT 14.928 30.392 14.96 30.424 ;
  LAYER M1 ;
        RECT 14.992 27.936 15.024 30.444 ;
  LAYER M3 ;
        RECT 14.992 27.956 15.024 27.988 ;
  LAYER M1 ;
        RECT 15.056 27.936 15.088 30.444 ;
  LAYER M3 ;
        RECT 15.056 30.392 15.088 30.424 ;
  LAYER M1 ;
        RECT 15.12 27.936 15.152 30.444 ;
  LAYER M3 ;
        RECT 15.12 27.956 15.152 27.988 ;
  LAYER M1 ;
        RECT 15.184 27.936 15.216 30.444 ;
  LAYER M3 ;
        RECT 15.184 30.392 15.216 30.424 ;
  LAYER M1 ;
        RECT 15.248 27.936 15.28 30.444 ;
  LAYER M3 ;
        RECT 15.248 27.956 15.28 27.988 ;
  LAYER M1 ;
        RECT 15.312 27.936 15.344 30.444 ;
  LAYER M3 ;
        RECT 15.312 30.392 15.344 30.424 ;
  LAYER M1 ;
        RECT 15.376 27.936 15.408 30.444 ;
  LAYER M3 ;
        RECT 15.376 27.956 15.408 27.988 ;
  LAYER M1 ;
        RECT 15.44 27.936 15.472 30.444 ;
  LAYER M3 ;
        RECT 13.072 30.328 13.104 30.36 ;
  LAYER M2 ;
        RECT 15.44 30.264 15.472 30.296 ;
  LAYER M2 ;
        RECT 13.072 30.2 13.104 30.232 ;
  LAYER M2 ;
        RECT 15.44 30.136 15.472 30.168 ;
  LAYER M2 ;
        RECT 13.072 30.072 13.104 30.104 ;
  LAYER M2 ;
        RECT 15.44 30.008 15.472 30.04 ;
  LAYER M2 ;
        RECT 13.072 29.944 13.104 29.976 ;
  LAYER M2 ;
        RECT 15.44 29.88 15.472 29.912 ;
  LAYER M2 ;
        RECT 13.072 29.816 13.104 29.848 ;
  LAYER M2 ;
        RECT 15.44 29.752 15.472 29.784 ;
  LAYER M2 ;
        RECT 13.072 29.688 13.104 29.72 ;
  LAYER M2 ;
        RECT 15.44 29.624 15.472 29.656 ;
  LAYER M2 ;
        RECT 13.072 29.56 13.104 29.592 ;
  LAYER M2 ;
        RECT 15.44 29.496 15.472 29.528 ;
  LAYER M2 ;
        RECT 13.072 29.432 13.104 29.464 ;
  LAYER M2 ;
        RECT 15.44 29.368 15.472 29.4 ;
  LAYER M2 ;
        RECT 13.072 29.304 13.104 29.336 ;
  LAYER M2 ;
        RECT 15.44 29.24 15.472 29.272 ;
  LAYER M2 ;
        RECT 13.072 29.176 13.104 29.208 ;
  LAYER M2 ;
        RECT 15.44 29.112 15.472 29.144 ;
  LAYER M2 ;
        RECT 13.072 29.048 13.104 29.08 ;
  LAYER M2 ;
        RECT 15.44 28.984 15.472 29.016 ;
  LAYER M2 ;
        RECT 13.072 28.92 13.104 28.952 ;
  LAYER M2 ;
        RECT 15.44 28.856 15.472 28.888 ;
  LAYER M2 ;
        RECT 13.072 28.792 13.104 28.824 ;
  LAYER M2 ;
        RECT 15.44 28.728 15.472 28.76 ;
  LAYER M2 ;
        RECT 13.072 28.664 13.104 28.696 ;
  LAYER M2 ;
        RECT 15.44 28.6 15.472 28.632 ;
  LAYER M2 ;
        RECT 13.072 28.536 13.104 28.568 ;
  LAYER M2 ;
        RECT 15.44 28.472 15.472 28.504 ;
  LAYER M2 ;
        RECT 13.072 28.408 13.104 28.44 ;
  LAYER M2 ;
        RECT 15.44 28.344 15.472 28.376 ;
  LAYER M2 ;
        RECT 13.072 28.28 13.104 28.312 ;
  LAYER M2 ;
        RECT 15.44 28.216 15.472 28.248 ;
  LAYER M2 ;
        RECT 13.072 28.152 13.104 28.184 ;
  LAYER M2 ;
        RECT 15.44 28.088 15.472 28.12 ;
  LAYER M2 ;
        RECT 13.024 27.888 15.52 30.492 ;
  LAYER M1 ;
        RECT 13.072 24.828 13.104 27.336 ;
  LAYER M3 ;
        RECT 13.072 24.848 13.104 24.88 ;
  LAYER M1 ;
        RECT 13.136 24.828 13.168 27.336 ;
  LAYER M3 ;
        RECT 13.136 27.284 13.168 27.316 ;
  LAYER M1 ;
        RECT 13.2 24.828 13.232 27.336 ;
  LAYER M3 ;
        RECT 13.2 24.848 13.232 24.88 ;
  LAYER M1 ;
        RECT 13.264 24.828 13.296 27.336 ;
  LAYER M3 ;
        RECT 13.264 27.284 13.296 27.316 ;
  LAYER M1 ;
        RECT 13.328 24.828 13.36 27.336 ;
  LAYER M3 ;
        RECT 13.328 24.848 13.36 24.88 ;
  LAYER M1 ;
        RECT 13.392 24.828 13.424 27.336 ;
  LAYER M3 ;
        RECT 13.392 27.284 13.424 27.316 ;
  LAYER M1 ;
        RECT 13.456 24.828 13.488 27.336 ;
  LAYER M3 ;
        RECT 13.456 24.848 13.488 24.88 ;
  LAYER M1 ;
        RECT 13.52 24.828 13.552 27.336 ;
  LAYER M3 ;
        RECT 13.52 27.284 13.552 27.316 ;
  LAYER M1 ;
        RECT 13.584 24.828 13.616 27.336 ;
  LAYER M3 ;
        RECT 13.584 24.848 13.616 24.88 ;
  LAYER M1 ;
        RECT 13.648 24.828 13.68 27.336 ;
  LAYER M3 ;
        RECT 13.648 27.284 13.68 27.316 ;
  LAYER M1 ;
        RECT 13.712 24.828 13.744 27.336 ;
  LAYER M3 ;
        RECT 13.712 24.848 13.744 24.88 ;
  LAYER M1 ;
        RECT 13.776 24.828 13.808 27.336 ;
  LAYER M3 ;
        RECT 13.776 27.284 13.808 27.316 ;
  LAYER M1 ;
        RECT 13.84 24.828 13.872 27.336 ;
  LAYER M3 ;
        RECT 13.84 24.848 13.872 24.88 ;
  LAYER M1 ;
        RECT 13.904 24.828 13.936 27.336 ;
  LAYER M3 ;
        RECT 13.904 27.284 13.936 27.316 ;
  LAYER M1 ;
        RECT 13.968 24.828 14 27.336 ;
  LAYER M3 ;
        RECT 13.968 24.848 14 24.88 ;
  LAYER M1 ;
        RECT 14.032 24.828 14.064 27.336 ;
  LAYER M3 ;
        RECT 14.032 27.284 14.064 27.316 ;
  LAYER M1 ;
        RECT 14.096 24.828 14.128 27.336 ;
  LAYER M3 ;
        RECT 14.096 24.848 14.128 24.88 ;
  LAYER M1 ;
        RECT 14.16 24.828 14.192 27.336 ;
  LAYER M3 ;
        RECT 14.16 27.284 14.192 27.316 ;
  LAYER M1 ;
        RECT 14.224 24.828 14.256 27.336 ;
  LAYER M3 ;
        RECT 14.224 24.848 14.256 24.88 ;
  LAYER M1 ;
        RECT 14.288 24.828 14.32 27.336 ;
  LAYER M3 ;
        RECT 14.288 27.284 14.32 27.316 ;
  LAYER M1 ;
        RECT 14.352 24.828 14.384 27.336 ;
  LAYER M3 ;
        RECT 14.352 24.848 14.384 24.88 ;
  LAYER M1 ;
        RECT 14.416 24.828 14.448 27.336 ;
  LAYER M3 ;
        RECT 14.416 27.284 14.448 27.316 ;
  LAYER M1 ;
        RECT 14.48 24.828 14.512 27.336 ;
  LAYER M3 ;
        RECT 14.48 24.848 14.512 24.88 ;
  LAYER M1 ;
        RECT 14.544 24.828 14.576 27.336 ;
  LAYER M3 ;
        RECT 14.544 27.284 14.576 27.316 ;
  LAYER M1 ;
        RECT 14.608 24.828 14.64 27.336 ;
  LAYER M3 ;
        RECT 14.608 24.848 14.64 24.88 ;
  LAYER M1 ;
        RECT 14.672 24.828 14.704 27.336 ;
  LAYER M3 ;
        RECT 14.672 27.284 14.704 27.316 ;
  LAYER M1 ;
        RECT 14.736 24.828 14.768 27.336 ;
  LAYER M3 ;
        RECT 14.736 24.848 14.768 24.88 ;
  LAYER M1 ;
        RECT 14.8 24.828 14.832 27.336 ;
  LAYER M3 ;
        RECT 14.8 27.284 14.832 27.316 ;
  LAYER M1 ;
        RECT 14.864 24.828 14.896 27.336 ;
  LAYER M3 ;
        RECT 14.864 24.848 14.896 24.88 ;
  LAYER M1 ;
        RECT 14.928 24.828 14.96 27.336 ;
  LAYER M3 ;
        RECT 14.928 27.284 14.96 27.316 ;
  LAYER M1 ;
        RECT 14.992 24.828 15.024 27.336 ;
  LAYER M3 ;
        RECT 14.992 24.848 15.024 24.88 ;
  LAYER M1 ;
        RECT 15.056 24.828 15.088 27.336 ;
  LAYER M3 ;
        RECT 15.056 27.284 15.088 27.316 ;
  LAYER M1 ;
        RECT 15.12 24.828 15.152 27.336 ;
  LAYER M3 ;
        RECT 15.12 24.848 15.152 24.88 ;
  LAYER M1 ;
        RECT 15.184 24.828 15.216 27.336 ;
  LAYER M3 ;
        RECT 15.184 27.284 15.216 27.316 ;
  LAYER M1 ;
        RECT 15.248 24.828 15.28 27.336 ;
  LAYER M3 ;
        RECT 15.248 24.848 15.28 24.88 ;
  LAYER M1 ;
        RECT 15.312 24.828 15.344 27.336 ;
  LAYER M3 ;
        RECT 15.312 27.284 15.344 27.316 ;
  LAYER M1 ;
        RECT 15.376 24.828 15.408 27.336 ;
  LAYER M3 ;
        RECT 15.376 24.848 15.408 24.88 ;
  LAYER M1 ;
        RECT 15.44 24.828 15.472 27.336 ;
  LAYER M3 ;
        RECT 13.072 27.22 13.104 27.252 ;
  LAYER M2 ;
        RECT 15.44 27.156 15.472 27.188 ;
  LAYER M2 ;
        RECT 13.072 27.092 13.104 27.124 ;
  LAYER M2 ;
        RECT 15.44 27.028 15.472 27.06 ;
  LAYER M2 ;
        RECT 13.072 26.964 13.104 26.996 ;
  LAYER M2 ;
        RECT 15.44 26.9 15.472 26.932 ;
  LAYER M2 ;
        RECT 13.072 26.836 13.104 26.868 ;
  LAYER M2 ;
        RECT 15.44 26.772 15.472 26.804 ;
  LAYER M2 ;
        RECT 13.072 26.708 13.104 26.74 ;
  LAYER M2 ;
        RECT 15.44 26.644 15.472 26.676 ;
  LAYER M2 ;
        RECT 13.072 26.58 13.104 26.612 ;
  LAYER M2 ;
        RECT 15.44 26.516 15.472 26.548 ;
  LAYER M2 ;
        RECT 13.072 26.452 13.104 26.484 ;
  LAYER M2 ;
        RECT 15.44 26.388 15.472 26.42 ;
  LAYER M2 ;
        RECT 13.072 26.324 13.104 26.356 ;
  LAYER M2 ;
        RECT 15.44 26.26 15.472 26.292 ;
  LAYER M2 ;
        RECT 13.072 26.196 13.104 26.228 ;
  LAYER M2 ;
        RECT 15.44 26.132 15.472 26.164 ;
  LAYER M2 ;
        RECT 13.072 26.068 13.104 26.1 ;
  LAYER M2 ;
        RECT 15.44 26.004 15.472 26.036 ;
  LAYER M2 ;
        RECT 13.072 25.94 13.104 25.972 ;
  LAYER M2 ;
        RECT 15.44 25.876 15.472 25.908 ;
  LAYER M2 ;
        RECT 13.072 25.812 13.104 25.844 ;
  LAYER M2 ;
        RECT 15.44 25.748 15.472 25.78 ;
  LAYER M2 ;
        RECT 13.072 25.684 13.104 25.716 ;
  LAYER M2 ;
        RECT 15.44 25.62 15.472 25.652 ;
  LAYER M2 ;
        RECT 13.072 25.556 13.104 25.588 ;
  LAYER M2 ;
        RECT 15.44 25.492 15.472 25.524 ;
  LAYER M2 ;
        RECT 13.072 25.428 13.104 25.46 ;
  LAYER M2 ;
        RECT 15.44 25.364 15.472 25.396 ;
  LAYER M2 ;
        RECT 13.072 25.3 13.104 25.332 ;
  LAYER M2 ;
        RECT 15.44 25.236 15.472 25.268 ;
  LAYER M2 ;
        RECT 13.072 25.172 13.104 25.204 ;
  LAYER M2 ;
        RECT 15.44 25.108 15.472 25.14 ;
  LAYER M2 ;
        RECT 13.072 25.044 13.104 25.076 ;
  LAYER M2 ;
        RECT 15.44 24.98 15.472 25.012 ;
  LAYER M2 ;
        RECT 13.024 24.78 15.52 27.384 ;
  LAYER M1 ;
        RECT 13.072 21.72 13.104 24.228 ;
  LAYER M3 ;
        RECT 13.072 21.74 13.104 21.772 ;
  LAYER M1 ;
        RECT 13.136 21.72 13.168 24.228 ;
  LAYER M3 ;
        RECT 13.136 24.176 13.168 24.208 ;
  LAYER M1 ;
        RECT 13.2 21.72 13.232 24.228 ;
  LAYER M3 ;
        RECT 13.2 21.74 13.232 21.772 ;
  LAYER M1 ;
        RECT 13.264 21.72 13.296 24.228 ;
  LAYER M3 ;
        RECT 13.264 24.176 13.296 24.208 ;
  LAYER M1 ;
        RECT 13.328 21.72 13.36 24.228 ;
  LAYER M3 ;
        RECT 13.328 21.74 13.36 21.772 ;
  LAYER M1 ;
        RECT 13.392 21.72 13.424 24.228 ;
  LAYER M3 ;
        RECT 13.392 24.176 13.424 24.208 ;
  LAYER M1 ;
        RECT 13.456 21.72 13.488 24.228 ;
  LAYER M3 ;
        RECT 13.456 21.74 13.488 21.772 ;
  LAYER M1 ;
        RECT 13.52 21.72 13.552 24.228 ;
  LAYER M3 ;
        RECT 13.52 24.176 13.552 24.208 ;
  LAYER M1 ;
        RECT 13.584 21.72 13.616 24.228 ;
  LAYER M3 ;
        RECT 13.584 21.74 13.616 21.772 ;
  LAYER M1 ;
        RECT 13.648 21.72 13.68 24.228 ;
  LAYER M3 ;
        RECT 13.648 24.176 13.68 24.208 ;
  LAYER M1 ;
        RECT 13.712 21.72 13.744 24.228 ;
  LAYER M3 ;
        RECT 13.712 21.74 13.744 21.772 ;
  LAYER M1 ;
        RECT 13.776 21.72 13.808 24.228 ;
  LAYER M3 ;
        RECT 13.776 24.176 13.808 24.208 ;
  LAYER M1 ;
        RECT 13.84 21.72 13.872 24.228 ;
  LAYER M3 ;
        RECT 13.84 21.74 13.872 21.772 ;
  LAYER M1 ;
        RECT 13.904 21.72 13.936 24.228 ;
  LAYER M3 ;
        RECT 13.904 24.176 13.936 24.208 ;
  LAYER M1 ;
        RECT 13.968 21.72 14 24.228 ;
  LAYER M3 ;
        RECT 13.968 21.74 14 21.772 ;
  LAYER M1 ;
        RECT 14.032 21.72 14.064 24.228 ;
  LAYER M3 ;
        RECT 14.032 24.176 14.064 24.208 ;
  LAYER M1 ;
        RECT 14.096 21.72 14.128 24.228 ;
  LAYER M3 ;
        RECT 14.096 21.74 14.128 21.772 ;
  LAYER M1 ;
        RECT 14.16 21.72 14.192 24.228 ;
  LAYER M3 ;
        RECT 14.16 24.176 14.192 24.208 ;
  LAYER M1 ;
        RECT 14.224 21.72 14.256 24.228 ;
  LAYER M3 ;
        RECT 14.224 21.74 14.256 21.772 ;
  LAYER M1 ;
        RECT 14.288 21.72 14.32 24.228 ;
  LAYER M3 ;
        RECT 14.288 24.176 14.32 24.208 ;
  LAYER M1 ;
        RECT 14.352 21.72 14.384 24.228 ;
  LAYER M3 ;
        RECT 14.352 21.74 14.384 21.772 ;
  LAYER M1 ;
        RECT 14.416 21.72 14.448 24.228 ;
  LAYER M3 ;
        RECT 14.416 24.176 14.448 24.208 ;
  LAYER M1 ;
        RECT 14.48 21.72 14.512 24.228 ;
  LAYER M3 ;
        RECT 14.48 21.74 14.512 21.772 ;
  LAYER M1 ;
        RECT 14.544 21.72 14.576 24.228 ;
  LAYER M3 ;
        RECT 14.544 24.176 14.576 24.208 ;
  LAYER M1 ;
        RECT 14.608 21.72 14.64 24.228 ;
  LAYER M3 ;
        RECT 14.608 21.74 14.64 21.772 ;
  LAYER M1 ;
        RECT 14.672 21.72 14.704 24.228 ;
  LAYER M3 ;
        RECT 14.672 24.176 14.704 24.208 ;
  LAYER M1 ;
        RECT 14.736 21.72 14.768 24.228 ;
  LAYER M3 ;
        RECT 14.736 21.74 14.768 21.772 ;
  LAYER M1 ;
        RECT 14.8 21.72 14.832 24.228 ;
  LAYER M3 ;
        RECT 14.8 24.176 14.832 24.208 ;
  LAYER M1 ;
        RECT 14.864 21.72 14.896 24.228 ;
  LAYER M3 ;
        RECT 14.864 21.74 14.896 21.772 ;
  LAYER M1 ;
        RECT 14.928 21.72 14.96 24.228 ;
  LAYER M3 ;
        RECT 14.928 24.176 14.96 24.208 ;
  LAYER M1 ;
        RECT 14.992 21.72 15.024 24.228 ;
  LAYER M3 ;
        RECT 14.992 21.74 15.024 21.772 ;
  LAYER M1 ;
        RECT 15.056 21.72 15.088 24.228 ;
  LAYER M3 ;
        RECT 15.056 24.176 15.088 24.208 ;
  LAYER M1 ;
        RECT 15.12 21.72 15.152 24.228 ;
  LAYER M3 ;
        RECT 15.12 21.74 15.152 21.772 ;
  LAYER M1 ;
        RECT 15.184 21.72 15.216 24.228 ;
  LAYER M3 ;
        RECT 15.184 24.176 15.216 24.208 ;
  LAYER M1 ;
        RECT 15.248 21.72 15.28 24.228 ;
  LAYER M3 ;
        RECT 15.248 21.74 15.28 21.772 ;
  LAYER M1 ;
        RECT 15.312 21.72 15.344 24.228 ;
  LAYER M3 ;
        RECT 15.312 24.176 15.344 24.208 ;
  LAYER M1 ;
        RECT 15.376 21.72 15.408 24.228 ;
  LAYER M3 ;
        RECT 15.376 21.74 15.408 21.772 ;
  LAYER M1 ;
        RECT 15.44 21.72 15.472 24.228 ;
  LAYER M3 ;
        RECT 13.072 24.112 13.104 24.144 ;
  LAYER M2 ;
        RECT 15.44 24.048 15.472 24.08 ;
  LAYER M2 ;
        RECT 13.072 23.984 13.104 24.016 ;
  LAYER M2 ;
        RECT 15.44 23.92 15.472 23.952 ;
  LAYER M2 ;
        RECT 13.072 23.856 13.104 23.888 ;
  LAYER M2 ;
        RECT 15.44 23.792 15.472 23.824 ;
  LAYER M2 ;
        RECT 13.072 23.728 13.104 23.76 ;
  LAYER M2 ;
        RECT 15.44 23.664 15.472 23.696 ;
  LAYER M2 ;
        RECT 13.072 23.6 13.104 23.632 ;
  LAYER M2 ;
        RECT 15.44 23.536 15.472 23.568 ;
  LAYER M2 ;
        RECT 13.072 23.472 13.104 23.504 ;
  LAYER M2 ;
        RECT 15.44 23.408 15.472 23.44 ;
  LAYER M2 ;
        RECT 13.072 23.344 13.104 23.376 ;
  LAYER M2 ;
        RECT 15.44 23.28 15.472 23.312 ;
  LAYER M2 ;
        RECT 13.072 23.216 13.104 23.248 ;
  LAYER M2 ;
        RECT 15.44 23.152 15.472 23.184 ;
  LAYER M2 ;
        RECT 13.072 23.088 13.104 23.12 ;
  LAYER M2 ;
        RECT 15.44 23.024 15.472 23.056 ;
  LAYER M2 ;
        RECT 13.072 22.96 13.104 22.992 ;
  LAYER M2 ;
        RECT 15.44 22.896 15.472 22.928 ;
  LAYER M2 ;
        RECT 13.072 22.832 13.104 22.864 ;
  LAYER M2 ;
        RECT 15.44 22.768 15.472 22.8 ;
  LAYER M2 ;
        RECT 13.072 22.704 13.104 22.736 ;
  LAYER M2 ;
        RECT 15.44 22.64 15.472 22.672 ;
  LAYER M2 ;
        RECT 13.072 22.576 13.104 22.608 ;
  LAYER M2 ;
        RECT 15.44 22.512 15.472 22.544 ;
  LAYER M2 ;
        RECT 13.072 22.448 13.104 22.48 ;
  LAYER M2 ;
        RECT 15.44 22.384 15.472 22.416 ;
  LAYER M2 ;
        RECT 13.072 22.32 13.104 22.352 ;
  LAYER M2 ;
        RECT 15.44 22.256 15.472 22.288 ;
  LAYER M2 ;
        RECT 13.072 22.192 13.104 22.224 ;
  LAYER M2 ;
        RECT 15.44 22.128 15.472 22.16 ;
  LAYER M2 ;
        RECT 13.072 22.064 13.104 22.096 ;
  LAYER M2 ;
        RECT 15.44 22 15.472 22.032 ;
  LAYER M2 ;
        RECT 13.072 21.936 13.104 21.968 ;
  LAYER M2 ;
        RECT 15.44 21.872 15.472 21.904 ;
  LAYER M2 ;
        RECT 13.024 21.672 15.52 24.276 ;
  LAYER M1 ;
        RECT 13.072 18.612 13.104 21.12 ;
  LAYER M3 ;
        RECT 13.072 18.632 13.104 18.664 ;
  LAYER M1 ;
        RECT 13.136 18.612 13.168 21.12 ;
  LAYER M3 ;
        RECT 13.136 21.068 13.168 21.1 ;
  LAYER M1 ;
        RECT 13.2 18.612 13.232 21.12 ;
  LAYER M3 ;
        RECT 13.2 18.632 13.232 18.664 ;
  LAYER M1 ;
        RECT 13.264 18.612 13.296 21.12 ;
  LAYER M3 ;
        RECT 13.264 21.068 13.296 21.1 ;
  LAYER M1 ;
        RECT 13.328 18.612 13.36 21.12 ;
  LAYER M3 ;
        RECT 13.328 18.632 13.36 18.664 ;
  LAYER M1 ;
        RECT 13.392 18.612 13.424 21.12 ;
  LAYER M3 ;
        RECT 13.392 21.068 13.424 21.1 ;
  LAYER M1 ;
        RECT 13.456 18.612 13.488 21.12 ;
  LAYER M3 ;
        RECT 13.456 18.632 13.488 18.664 ;
  LAYER M1 ;
        RECT 13.52 18.612 13.552 21.12 ;
  LAYER M3 ;
        RECT 13.52 21.068 13.552 21.1 ;
  LAYER M1 ;
        RECT 13.584 18.612 13.616 21.12 ;
  LAYER M3 ;
        RECT 13.584 18.632 13.616 18.664 ;
  LAYER M1 ;
        RECT 13.648 18.612 13.68 21.12 ;
  LAYER M3 ;
        RECT 13.648 21.068 13.68 21.1 ;
  LAYER M1 ;
        RECT 13.712 18.612 13.744 21.12 ;
  LAYER M3 ;
        RECT 13.712 18.632 13.744 18.664 ;
  LAYER M1 ;
        RECT 13.776 18.612 13.808 21.12 ;
  LAYER M3 ;
        RECT 13.776 21.068 13.808 21.1 ;
  LAYER M1 ;
        RECT 13.84 18.612 13.872 21.12 ;
  LAYER M3 ;
        RECT 13.84 18.632 13.872 18.664 ;
  LAYER M1 ;
        RECT 13.904 18.612 13.936 21.12 ;
  LAYER M3 ;
        RECT 13.904 21.068 13.936 21.1 ;
  LAYER M1 ;
        RECT 13.968 18.612 14 21.12 ;
  LAYER M3 ;
        RECT 13.968 18.632 14 18.664 ;
  LAYER M1 ;
        RECT 14.032 18.612 14.064 21.12 ;
  LAYER M3 ;
        RECT 14.032 21.068 14.064 21.1 ;
  LAYER M1 ;
        RECT 14.096 18.612 14.128 21.12 ;
  LAYER M3 ;
        RECT 14.096 18.632 14.128 18.664 ;
  LAYER M1 ;
        RECT 14.16 18.612 14.192 21.12 ;
  LAYER M3 ;
        RECT 14.16 21.068 14.192 21.1 ;
  LAYER M1 ;
        RECT 14.224 18.612 14.256 21.12 ;
  LAYER M3 ;
        RECT 14.224 18.632 14.256 18.664 ;
  LAYER M1 ;
        RECT 14.288 18.612 14.32 21.12 ;
  LAYER M3 ;
        RECT 14.288 21.068 14.32 21.1 ;
  LAYER M1 ;
        RECT 14.352 18.612 14.384 21.12 ;
  LAYER M3 ;
        RECT 14.352 18.632 14.384 18.664 ;
  LAYER M1 ;
        RECT 14.416 18.612 14.448 21.12 ;
  LAYER M3 ;
        RECT 14.416 21.068 14.448 21.1 ;
  LAYER M1 ;
        RECT 14.48 18.612 14.512 21.12 ;
  LAYER M3 ;
        RECT 14.48 18.632 14.512 18.664 ;
  LAYER M1 ;
        RECT 14.544 18.612 14.576 21.12 ;
  LAYER M3 ;
        RECT 14.544 21.068 14.576 21.1 ;
  LAYER M1 ;
        RECT 14.608 18.612 14.64 21.12 ;
  LAYER M3 ;
        RECT 14.608 18.632 14.64 18.664 ;
  LAYER M1 ;
        RECT 14.672 18.612 14.704 21.12 ;
  LAYER M3 ;
        RECT 14.672 21.068 14.704 21.1 ;
  LAYER M1 ;
        RECT 14.736 18.612 14.768 21.12 ;
  LAYER M3 ;
        RECT 14.736 18.632 14.768 18.664 ;
  LAYER M1 ;
        RECT 14.8 18.612 14.832 21.12 ;
  LAYER M3 ;
        RECT 14.8 21.068 14.832 21.1 ;
  LAYER M1 ;
        RECT 14.864 18.612 14.896 21.12 ;
  LAYER M3 ;
        RECT 14.864 18.632 14.896 18.664 ;
  LAYER M1 ;
        RECT 14.928 18.612 14.96 21.12 ;
  LAYER M3 ;
        RECT 14.928 21.068 14.96 21.1 ;
  LAYER M1 ;
        RECT 14.992 18.612 15.024 21.12 ;
  LAYER M3 ;
        RECT 14.992 18.632 15.024 18.664 ;
  LAYER M1 ;
        RECT 15.056 18.612 15.088 21.12 ;
  LAYER M3 ;
        RECT 15.056 21.068 15.088 21.1 ;
  LAYER M1 ;
        RECT 15.12 18.612 15.152 21.12 ;
  LAYER M3 ;
        RECT 15.12 18.632 15.152 18.664 ;
  LAYER M1 ;
        RECT 15.184 18.612 15.216 21.12 ;
  LAYER M3 ;
        RECT 15.184 21.068 15.216 21.1 ;
  LAYER M1 ;
        RECT 15.248 18.612 15.28 21.12 ;
  LAYER M3 ;
        RECT 15.248 18.632 15.28 18.664 ;
  LAYER M1 ;
        RECT 15.312 18.612 15.344 21.12 ;
  LAYER M3 ;
        RECT 15.312 21.068 15.344 21.1 ;
  LAYER M1 ;
        RECT 15.376 18.612 15.408 21.12 ;
  LAYER M3 ;
        RECT 15.376 18.632 15.408 18.664 ;
  LAYER M1 ;
        RECT 15.44 18.612 15.472 21.12 ;
  LAYER M3 ;
        RECT 13.072 21.004 13.104 21.036 ;
  LAYER M2 ;
        RECT 15.44 20.94 15.472 20.972 ;
  LAYER M2 ;
        RECT 13.072 20.876 13.104 20.908 ;
  LAYER M2 ;
        RECT 15.44 20.812 15.472 20.844 ;
  LAYER M2 ;
        RECT 13.072 20.748 13.104 20.78 ;
  LAYER M2 ;
        RECT 15.44 20.684 15.472 20.716 ;
  LAYER M2 ;
        RECT 13.072 20.62 13.104 20.652 ;
  LAYER M2 ;
        RECT 15.44 20.556 15.472 20.588 ;
  LAYER M2 ;
        RECT 13.072 20.492 13.104 20.524 ;
  LAYER M2 ;
        RECT 15.44 20.428 15.472 20.46 ;
  LAYER M2 ;
        RECT 13.072 20.364 13.104 20.396 ;
  LAYER M2 ;
        RECT 15.44 20.3 15.472 20.332 ;
  LAYER M2 ;
        RECT 13.072 20.236 13.104 20.268 ;
  LAYER M2 ;
        RECT 15.44 20.172 15.472 20.204 ;
  LAYER M2 ;
        RECT 13.072 20.108 13.104 20.14 ;
  LAYER M2 ;
        RECT 15.44 20.044 15.472 20.076 ;
  LAYER M2 ;
        RECT 13.072 19.98 13.104 20.012 ;
  LAYER M2 ;
        RECT 15.44 19.916 15.472 19.948 ;
  LAYER M2 ;
        RECT 13.072 19.852 13.104 19.884 ;
  LAYER M2 ;
        RECT 15.44 19.788 15.472 19.82 ;
  LAYER M2 ;
        RECT 13.072 19.724 13.104 19.756 ;
  LAYER M2 ;
        RECT 15.44 19.66 15.472 19.692 ;
  LAYER M2 ;
        RECT 13.072 19.596 13.104 19.628 ;
  LAYER M2 ;
        RECT 15.44 19.532 15.472 19.564 ;
  LAYER M2 ;
        RECT 13.072 19.468 13.104 19.5 ;
  LAYER M2 ;
        RECT 15.44 19.404 15.472 19.436 ;
  LAYER M2 ;
        RECT 13.072 19.34 13.104 19.372 ;
  LAYER M2 ;
        RECT 15.44 19.276 15.472 19.308 ;
  LAYER M2 ;
        RECT 13.072 19.212 13.104 19.244 ;
  LAYER M2 ;
        RECT 15.44 19.148 15.472 19.18 ;
  LAYER M2 ;
        RECT 13.072 19.084 13.104 19.116 ;
  LAYER M2 ;
        RECT 15.44 19.02 15.472 19.052 ;
  LAYER M2 ;
        RECT 13.072 18.956 13.104 18.988 ;
  LAYER M2 ;
        RECT 15.44 18.892 15.472 18.924 ;
  LAYER M2 ;
        RECT 13.072 18.828 13.104 18.86 ;
  LAYER M2 ;
        RECT 15.44 18.764 15.472 18.796 ;
  LAYER M2 ;
        RECT 13.024 18.564 15.52 21.168 ;
  LAYER M1 ;
        RECT 13.072 15.504 13.104 18.012 ;
  LAYER M3 ;
        RECT 13.072 15.524 13.104 15.556 ;
  LAYER M1 ;
        RECT 13.136 15.504 13.168 18.012 ;
  LAYER M3 ;
        RECT 13.136 17.96 13.168 17.992 ;
  LAYER M1 ;
        RECT 13.2 15.504 13.232 18.012 ;
  LAYER M3 ;
        RECT 13.2 15.524 13.232 15.556 ;
  LAYER M1 ;
        RECT 13.264 15.504 13.296 18.012 ;
  LAYER M3 ;
        RECT 13.264 17.96 13.296 17.992 ;
  LAYER M1 ;
        RECT 13.328 15.504 13.36 18.012 ;
  LAYER M3 ;
        RECT 13.328 15.524 13.36 15.556 ;
  LAYER M1 ;
        RECT 13.392 15.504 13.424 18.012 ;
  LAYER M3 ;
        RECT 13.392 17.96 13.424 17.992 ;
  LAYER M1 ;
        RECT 13.456 15.504 13.488 18.012 ;
  LAYER M3 ;
        RECT 13.456 15.524 13.488 15.556 ;
  LAYER M1 ;
        RECT 13.52 15.504 13.552 18.012 ;
  LAYER M3 ;
        RECT 13.52 17.96 13.552 17.992 ;
  LAYER M1 ;
        RECT 13.584 15.504 13.616 18.012 ;
  LAYER M3 ;
        RECT 13.584 15.524 13.616 15.556 ;
  LAYER M1 ;
        RECT 13.648 15.504 13.68 18.012 ;
  LAYER M3 ;
        RECT 13.648 17.96 13.68 17.992 ;
  LAYER M1 ;
        RECT 13.712 15.504 13.744 18.012 ;
  LAYER M3 ;
        RECT 13.712 15.524 13.744 15.556 ;
  LAYER M1 ;
        RECT 13.776 15.504 13.808 18.012 ;
  LAYER M3 ;
        RECT 13.776 17.96 13.808 17.992 ;
  LAYER M1 ;
        RECT 13.84 15.504 13.872 18.012 ;
  LAYER M3 ;
        RECT 13.84 15.524 13.872 15.556 ;
  LAYER M1 ;
        RECT 13.904 15.504 13.936 18.012 ;
  LAYER M3 ;
        RECT 13.904 17.96 13.936 17.992 ;
  LAYER M1 ;
        RECT 13.968 15.504 14 18.012 ;
  LAYER M3 ;
        RECT 13.968 15.524 14 15.556 ;
  LAYER M1 ;
        RECT 14.032 15.504 14.064 18.012 ;
  LAYER M3 ;
        RECT 14.032 17.96 14.064 17.992 ;
  LAYER M1 ;
        RECT 14.096 15.504 14.128 18.012 ;
  LAYER M3 ;
        RECT 14.096 15.524 14.128 15.556 ;
  LAYER M1 ;
        RECT 14.16 15.504 14.192 18.012 ;
  LAYER M3 ;
        RECT 14.16 17.96 14.192 17.992 ;
  LAYER M1 ;
        RECT 14.224 15.504 14.256 18.012 ;
  LAYER M3 ;
        RECT 14.224 15.524 14.256 15.556 ;
  LAYER M1 ;
        RECT 14.288 15.504 14.32 18.012 ;
  LAYER M3 ;
        RECT 14.288 17.96 14.32 17.992 ;
  LAYER M1 ;
        RECT 14.352 15.504 14.384 18.012 ;
  LAYER M3 ;
        RECT 14.352 15.524 14.384 15.556 ;
  LAYER M1 ;
        RECT 14.416 15.504 14.448 18.012 ;
  LAYER M3 ;
        RECT 14.416 17.96 14.448 17.992 ;
  LAYER M1 ;
        RECT 14.48 15.504 14.512 18.012 ;
  LAYER M3 ;
        RECT 14.48 15.524 14.512 15.556 ;
  LAYER M1 ;
        RECT 14.544 15.504 14.576 18.012 ;
  LAYER M3 ;
        RECT 14.544 17.96 14.576 17.992 ;
  LAYER M1 ;
        RECT 14.608 15.504 14.64 18.012 ;
  LAYER M3 ;
        RECT 14.608 15.524 14.64 15.556 ;
  LAYER M1 ;
        RECT 14.672 15.504 14.704 18.012 ;
  LAYER M3 ;
        RECT 14.672 17.96 14.704 17.992 ;
  LAYER M1 ;
        RECT 14.736 15.504 14.768 18.012 ;
  LAYER M3 ;
        RECT 14.736 15.524 14.768 15.556 ;
  LAYER M1 ;
        RECT 14.8 15.504 14.832 18.012 ;
  LAYER M3 ;
        RECT 14.8 17.96 14.832 17.992 ;
  LAYER M1 ;
        RECT 14.864 15.504 14.896 18.012 ;
  LAYER M3 ;
        RECT 14.864 15.524 14.896 15.556 ;
  LAYER M1 ;
        RECT 14.928 15.504 14.96 18.012 ;
  LAYER M3 ;
        RECT 14.928 17.96 14.96 17.992 ;
  LAYER M1 ;
        RECT 14.992 15.504 15.024 18.012 ;
  LAYER M3 ;
        RECT 14.992 15.524 15.024 15.556 ;
  LAYER M1 ;
        RECT 15.056 15.504 15.088 18.012 ;
  LAYER M3 ;
        RECT 15.056 17.96 15.088 17.992 ;
  LAYER M1 ;
        RECT 15.12 15.504 15.152 18.012 ;
  LAYER M3 ;
        RECT 15.12 15.524 15.152 15.556 ;
  LAYER M1 ;
        RECT 15.184 15.504 15.216 18.012 ;
  LAYER M3 ;
        RECT 15.184 17.96 15.216 17.992 ;
  LAYER M1 ;
        RECT 15.248 15.504 15.28 18.012 ;
  LAYER M3 ;
        RECT 15.248 15.524 15.28 15.556 ;
  LAYER M1 ;
        RECT 15.312 15.504 15.344 18.012 ;
  LAYER M3 ;
        RECT 15.312 17.96 15.344 17.992 ;
  LAYER M1 ;
        RECT 15.376 15.504 15.408 18.012 ;
  LAYER M3 ;
        RECT 15.376 15.524 15.408 15.556 ;
  LAYER M1 ;
        RECT 15.44 15.504 15.472 18.012 ;
  LAYER M3 ;
        RECT 13.072 17.896 13.104 17.928 ;
  LAYER M2 ;
        RECT 15.44 17.832 15.472 17.864 ;
  LAYER M2 ;
        RECT 13.072 17.768 13.104 17.8 ;
  LAYER M2 ;
        RECT 15.44 17.704 15.472 17.736 ;
  LAYER M2 ;
        RECT 13.072 17.64 13.104 17.672 ;
  LAYER M2 ;
        RECT 15.44 17.576 15.472 17.608 ;
  LAYER M2 ;
        RECT 13.072 17.512 13.104 17.544 ;
  LAYER M2 ;
        RECT 15.44 17.448 15.472 17.48 ;
  LAYER M2 ;
        RECT 13.072 17.384 13.104 17.416 ;
  LAYER M2 ;
        RECT 15.44 17.32 15.472 17.352 ;
  LAYER M2 ;
        RECT 13.072 17.256 13.104 17.288 ;
  LAYER M2 ;
        RECT 15.44 17.192 15.472 17.224 ;
  LAYER M2 ;
        RECT 13.072 17.128 13.104 17.16 ;
  LAYER M2 ;
        RECT 15.44 17.064 15.472 17.096 ;
  LAYER M2 ;
        RECT 13.072 17 13.104 17.032 ;
  LAYER M2 ;
        RECT 15.44 16.936 15.472 16.968 ;
  LAYER M2 ;
        RECT 13.072 16.872 13.104 16.904 ;
  LAYER M2 ;
        RECT 15.44 16.808 15.472 16.84 ;
  LAYER M2 ;
        RECT 13.072 16.744 13.104 16.776 ;
  LAYER M2 ;
        RECT 15.44 16.68 15.472 16.712 ;
  LAYER M2 ;
        RECT 13.072 16.616 13.104 16.648 ;
  LAYER M2 ;
        RECT 15.44 16.552 15.472 16.584 ;
  LAYER M2 ;
        RECT 13.072 16.488 13.104 16.52 ;
  LAYER M2 ;
        RECT 15.44 16.424 15.472 16.456 ;
  LAYER M2 ;
        RECT 13.072 16.36 13.104 16.392 ;
  LAYER M2 ;
        RECT 15.44 16.296 15.472 16.328 ;
  LAYER M2 ;
        RECT 13.072 16.232 13.104 16.264 ;
  LAYER M2 ;
        RECT 15.44 16.168 15.472 16.2 ;
  LAYER M2 ;
        RECT 13.072 16.104 13.104 16.136 ;
  LAYER M2 ;
        RECT 15.44 16.04 15.472 16.072 ;
  LAYER M2 ;
        RECT 13.072 15.976 13.104 16.008 ;
  LAYER M2 ;
        RECT 15.44 15.912 15.472 15.944 ;
  LAYER M2 ;
        RECT 13.072 15.848 13.104 15.88 ;
  LAYER M2 ;
        RECT 15.44 15.784 15.472 15.816 ;
  LAYER M2 ;
        RECT 13.072 15.72 13.104 15.752 ;
  LAYER M2 ;
        RECT 15.44 15.656 15.472 15.688 ;
  LAYER M2 ;
        RECT 13.024 15.456 15.52 18.06 ;
  END 
END switched_capacitor_combination
