module testcase_EA_placer ( 0, 1 ); 
input 0, 1;

CMC_PMOS_S_n12_X1_Y1_Pin_3 m1 ( .G1(0), .G2(3), .G3(29) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m2 ( .G1(2), .G2(5) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m3 ( .G1(2), .G2(3), .G3(4), .G4(6) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m4 ( .G1(4), .G2(7) );
CMC_PMOS_S_n12_X1_Y1_Pin_3 m5 ( .G1(5), .G2(8), .G3(10) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m6 ( .G1(6), .G2(8), .G3(11), .G4(9) );
CMC_PMOS_S_n12_X1_Y1_Pin_3 m7 ( .G1(7), .G2(9), .G3(12) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m8 ( .G1(10), .G2(13) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m9 ( .G1(11), .G2(13), .G3(15), .G4(14) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m10 ( .G1(12), .G2(14) );
CMC_PMOS_S_n12_X1_Y1_Pin_3 m11 ( .G1(15), .G2(1), .G3(28) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m12 ( .G1(16), .G2(18) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m13 ( .G1(16), .G2(29), .G3(17), .G4(19) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m14 ( .G1(17), .G2(20) );
CMC_PMOS_S_n12_X1_Y1_Pin_3 m15 ( .G1(18), .G2(23), .G3(21) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m16 ( .G1(19), .G2(21), .G3(22), .G4(24) );
CMC_PMOS_S_n12_X1_Y1_Pin_3 m17 ( .G1(22), .G2(20), .G3(25) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m18 ( .G1(23), .G2(26) );
CMC_PMOS_S_n12_X1_Y1_Pin_4 m19 ( .G1(24), .G2(26), .G3(27), .G4(28) );
CMC_PMOS_S_n12_X1_Y1_Pin_2 m20 ( .G1(25), .G2(27) );

endmodule

