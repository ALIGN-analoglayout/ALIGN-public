MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 15.04 BY 13.44 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 13.152 6.208 13.224 ;
      LAYER M2 ;
        RECT 6.156 13.172 6.228 13.204 ;
      LAYER M1 ;
        RECT 9.152 13.152 9.184 13.224 ;
      LAYER M2 ;
        RECT 9.132 13.172 9.204 13.204 ;
      LAYER M2 ;
        RECT 6.192 13.172 9.168 13.204 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
      LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
      LAYER M2 ;
        RECT 6.032 0.236 9.008 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 6.032 3.932 8.784 3.964 ;
  LAYER M1 ;
        RECT 6.016 3.912 6.048 3.984 ;
  LAYER M2 ;
        RECT 5.996 3.932 6.068 3.964 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M2 ;
        RECT 6.032 7.04 8.784 7.072 ;
  LAYER M1 ;
        RECT 6.016 7.02 6.048 7.092 ;
  LAYER M2 ;
        RECT 5.996 7.04 6.068 7.072 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M1 ;
        RECT 5.792 3.78 5.824 3.948 ;
  LAYER M1 ;
        RECT 5.792 3.744 5.824 3.816 ;
  LAYER M2 ;
        RECT 5.772 3.764 5.844 3.796 ;
  LAYER M2 ;
        RECT 5.808 3.764 6.032 3.796 ;
  LAYER M1 ;
        RECT 6.016 3.744 6.048 3.816 ;
  LAYER M2 ;
        RECT 5.996 3.764 6.068 3.796 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M1 ;
        RECT 5.792 6.888 5.824 7.056 ;
  LAYER M1 ;
        RECT 5.792 6.852 5.824 6.924 ;
  LAYER M2 ;
        RECT 5.772 6.872 5.844 6.904 ;
  LAYER M2 ;
        RECT 5.808 6.872 6.032 6.904 ;
  LAYER M1 ;
        RECT 6.016 6.852 6.048 6.924 ;
  LAYER M2 ;
        RECT 5.996 6.872 6.068 6.904 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.504 ;
  LAYER M1 ;
        RECT 6.016 0.504 6.048 7.056 ;
  LAYER M1 ;
        RECT 11.744 7.02 11.776 7.092 ;
  LAYER M2 ;
        RECT 11.724 7.04 11.796 7.072 ;
  LAYER M2 ;
        RECT 9.008 7.04 11.76 7.072 ;
  LAYER M1 ;
        RECT 8.992 7.02 9.024 7.092 ;
  LAYER M2 ;
        RECT 8.972 7.04 9.044 7.072 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 9.008 3.932 11.76 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
  LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
  LAYER M1 ;
        RECT 8.992 0.252 9.024 0.504 ;
  LAYER M1 ;
        RECT 8.992 0.504 9.024 7.056 ;
  LAYER M2 ;
        RECT 6.032 0.236 9.008 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M1 ;
        RECT 2.816 0.672 2.848 0.84 ;
  LAYER M1 ;
        RECT 2.816 0.636 2.848 0.708 ;
  LAYER M2 ;
        RECT 2.796 0.656 2.868 0.688 ;
  LAYER M2 ;
        RECT 2.832 0.656 3.056 0.688 ;
  LAYER M1 ;
        RECT 3.04 0.636 3.072 0.708 ;
  LAYER M2 ;
        RECT 3.02 0.656 3.092 0.688 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M1 ;
        RECT 2.816 3.78 2.848 3.948 ;
  LAYER M1 ;
        RECT 2.816 3.744 2.848 3.816 ;
  LAYER M2 ;
        RECT 2.796 3.764 2.868 3.796 ;
  LAYER M2 ;
        RECT 2.832 3.764 3.056 3.796 ;
  LAYER M1 ;
        RECT 3.04 3.744 3.072 3.816 ;
  LAYER M2 ;
        RECT 3.02 3.764 3.092 3.796 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M1 ;
        RECT 2.816 6.888 2.848 7.056 ;
  LAYER M1 ;
        RECT 2.816 6.852 2.848 6.924 ;
  LAYER M2 ;
        RECT 2.796 6.872 2.868 6.904 ;
  LAYER M2 ;
        RECT 2.832 6.872 3.056 6.904 ;
  LAYER M1 ;
        RECT 3.04 6.852 3.072 6.924 ;
  LAYER M2 ;
        RECT 3.02 6.872 3.092 6.904 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M1 ;
        RECT 2.816 9.996 2.848 10.164 ;
  LAYER M1 ;
        RECT 2.816 9.96 2.848 10.032 ;
  LAYER M2 ;
        RECT 2.796 9.98 2.868 10.012 ;
  LAYER M2 ;
        RECT 2.832 9.98 3.056 10.012 ;
  LAYER M1 ;
        RECT 3.04 9.96 3.072 10.032 ;
  LAYER M2 ;
        RECT 3.02 9.98 3.092 10.012 ;
  LAYER M1 ;
        RECT 5.792 0.804 5.824 0.876 ;
  LAYER M2 ;
        RECT 5.772 0.824 5.844 0.856 ;
  LAYER M2 ;
        RECT 3.056 0.824 5.808 0.856 ;
  LAYER M1 ;
        RECT 3.04 0.804 3.072 0.876 ;
  LAYER M2 ;
        RECT 3.02 0.824 3.092 0.856 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 3.056 10.148 5.808 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 3.04 0.048 3.072 0.12 ;
  LAYER M2 ;
        RECT 3.02 0.068 3.092 0.1 ;
  LAYER M1 ;
        RECT 3.04 0.084 3.072 0.504 ;
  LAYER M1 ;
        RECT 3.04 0.504 3.072 10.164 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M1 ;
        RECT 11.744 0.672 11.776 0.84 ;
  LAYER M1 ;
        RECT 11.744 0.636 11.776 0.708 ;
  LAYER M2 ;
        RECT 11.724 0.656 11.796 0.688 ;
  LAYER M2 ;
        RECT 11.76 0.656 11.984 0.688 ;
  LAYER M1 ;
        RECT 11.968 0.636 12 0.708 ;
  LAYER M2 ;
        RECT 11.948 0.656 12.02 0.688 ;
  LAYER M1 ;
        RECT 11.744 10.128 11.776 10.2 ;
  LAYER M2 ;
        RECT 11.724 10.148 11.796 10.18 ;
  LAYER M1 ;
        RECT 11.744 9.996 11.776 10.164 ;
  LAYER M1 ;
        RECT 11.744 9.96 11.776 10.032 ;
  LAYER M2 ;
        RECT 11.724 9.98 11.796 10.012 ;
  LAYER M2 ;
        RECT 11.76 9.98 11.984 10.012 ;
  LAYER M1 ;
        RECT 11.968 9.96 12 10.032 ;
  LAYER M2 ;
        RECT 11.948 9.98 12.02 10.012 ;
  LAYER M1 ;
        RECT 14.72 0.804 14.752 0.876 ;
  LAYER M2 ;
        RECT 14.7 0.824 14.772 0.856 ;
  LAYER M2 ;
        RECT 11.984 0.824 14.736 0.856 ;
  LAYER M1 ;
        RECT 11.968 0.804 12 0.876 ;
  LAYER M2 ;
        RECT 11.948 0.824 12.02 0.856 ;
  LAYER M1 ;
        RECT 14.72 3.912 14.752 3.984 ;
  LAYER M2 ;
        RECT 14.7 3.932 14.772 3.964 ;
  LAYER M2 ;
        RECT 11.984 3.932 14.736 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 14.72 7.02 14.752 7.092 ;
  LAYER M2 ;
        RECT 14.7 7.04 14.772 7.072 ;
  LAYER M2 ;
        RECT 11.984 7.04 14.736 7.072 ;
  LAYER M1 ;
        RECT 11.968 7.02 12 7.092 ;
  LAYER M2 ;
        RECT 11.948 7.04 12.02 7.072 ;
  LAYER M1 ;
        RECT 14.72 10.128 14.752 10.2 ;
  LAYER M2 ;
        RECT 14.7 10.148 14.772 10.18 ;
  LAYER M2 ;
        RECT 11.984 10.148 14.736 10.18 ;
  LAYER M1 ;
        RECT 11.968 10.128 12 10.2 ;
  LAYER M2 ;
        RECT 11.948 10.148 12.02 10.18 ;
  LAYER M1 ;
        RECT 11.968 0.048 12 0.12 ;
  LAYER M2 ;
        RECT 11.948 0.068 12.02 0.1 ;
  LAYER M1 ;
        RECT 11.968 0.084 12 0.504 ;
  LAYER M1 ;
        RECT 11.968 0.504 12 10.164 ;
  LAYER M2 ;
        RECT 3.056 0.068 11.984 0.1 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 8.784 10.18 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M1 ;
        RECT 8.768 0.804 8.8 0.876 ;
  LAYER M2 ;
        RECT 8.748 0.824 8.82 0.856 ;
  LAYER M2 ;
        RECT 8.784 0.824 11.76 0.856 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M1 ;
        RECT 6.4 6.348 6.432 6.42 ;
  LAYER M2 ;
        RECT 6.38 6.368 6.452 6.4 ;
  LAYER M2 ;
        RECT 6.192 6.368 6.416 6.4 ;
  LAYER M1 ;
        RECT 6.176 6.348 6.208 6.42 ;
  LAYER M2 ;
        RECT 6.156 6.368 6.228 6.4 ;
  LAYER M1 ;
        RECT 6.4 9.456 6.432 9.528 ;
  LAYER M2 ;
        RECT 6.38 9.476 6.452 9.508 ;
  LAYER M2 ;
        RECT 6.192 9.476 6.416 9.508 ;
  LAYER M1 ;
        RECT 6.176 9.456 6.208 9.528 ;
  LAYER M2 ;
        RECT 6.156 9.476 6.228 9.508 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M1 ;
        RECT 3.424 6.384 3.456 6.552 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 3.44 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M1 ;
        RECT 3.424 9.492 3.456 9.66 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.44 9.644 6.192 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 6.176 13.152 6.208 13.224 ;
  LAYER M2 ;
        RECT 6.156 13.172 6.228 13.204 ;
  LAYER M1 ;
        RECT 6.176 12.936 6.208 13.188 ;
  LAYER M1 ;
        RECT 6.176 6.384 6.208 12.936 ;
  LAYER M1 ;
        RECT 9.376 9.456 9.408 9.528 ;
  LAYER M2 ;
        RECT 9.356 9.476 9.428 9.508 ;
  LAYER M2 ;
        RECT 9.168 9.476 9.392 9.508 ;
  LAYER M1 ;
        RECT 9.152 9.456 9.184 9.528 ;
  LAYER M2 ;
        RECT 9.132 9.476 9.204 9.508 ;
  LAYER M1 ;
        RECT 9.376 6.348 9.408 6.42 ;
  LAYER M2 ;
        RECT 9.356 6.368 9.428 6.4 ;
  LAYER M2 ;
        RECT 9.168 6.368 9.392 6.4 ;
  LAYER M1 ;
        RECT 9.152 6.348 9.184 6.42 ;
  LAYER M2 ;
        RECT 9.132 6.368 9.204 6.4 ;
  LAYER M1 ;
        RECT 9.152 13.152 9.184 13.224 ;
  LAYER M2 ;
        RECT 9.132 13.172 9.204 13.204 ;
  LAYER M1 ;
        RECT 9.152 12.936 9.184 13.188 ;
  LAYER M1 ;
        RECT 9.152 6.384 9.184 12.936 ;
  LAYER M2 ;
        RECT 6.192 13.172 9.168 13.204 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M2 ;
        RECT 0.08 3.26 0.464 3.292 ;
  LAYER M1 ;
        RECT 0.064 3.24 0.096 3.312 ;
  LAYER M2 ;
        RECT 0.044 3.26 0.116 3.292 ;
  LAYER M1 ;
        RECT 0.448 6.348 0.48 6.42 ;
  LAYER M2 ;
        RECT 0.428 6.368 0.5 6.4 ;
  LAYER M2 ;
        RECT 0.08 6.368 0.464 6.4 ;
  LAYER M1 ;
        RECT 0.064 6.348 0.096 6.42 ;
  LAYER M2 ;
        RECT 0.044 6.368 0.116 6.4 ;
  LAYER M1 ;
        RECT 0.448 9.456 0.48 9.528 ;
  LAYER M2 ;
        RECT 0.428 9.476 0.5 9.508 ;
  LAYER M2 ;
        RECT 0.08 9.476 0.464 9.508 ;
  LAYER M1 ;
        RECT 0.064 9.456 0.096 9.528 ;
  LAYER M2 ;
        RECT 0.044 9.476 0.116 9.508 ;
  LAYER M1 ;
        RECT 0.448 12.564 0.48 12.636 ;
  LAYER M2 ;
        RECT 0.428 12.584 0.5 12.616 ;
  LAYER M2 ;
        RECT 0.08 12.584 0.464 12.616 ;
  LAYER M1 ;
        RECT 0.064 12.564 0.096 12.636 ;
  LAYER M2 ;
        RECT 0.044 12.584 0.116 12.616 ;
  LAYER M1 ;
        RECT 0.064 13.32 0.096 13.392 ;
  LAYER M2 ;
        RECT 0.044 13.34 0.116 13.372 ;
  LAYER M1 ;
        RECT 0.064 12.936 0.096 13.356 ;
  LAYER M1 ;
        RECT 0.064 3.276 0.096 12.936 ;
  LAYER M1 ;
        RECT 12.352 3.24 12.384 3.312 ;
  LAYER M2 ;
        RECT 12.332 3.26 12.404 3.292 ;
  LAYER M1 ;
        RECT 12.352 3.276 12.384 3.444 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M2 ;
        RECT 12.368 3.428 14.96 3.46 ;
  LAYER M1 ;
        RECT 14.944 3.408 14.976 3.48 ;
  LAYER M2 ;
        RECT 14.924 3.428 14.996 3.46 ;
  LAYER M1 ;
        RECT 12.352 6.348 12.384 6.42 ;
  LAYER M2 ;
        RECT 12.332 6.368 12.404 6.4 ;
  LAYER M1 ;
        RECT 12.352 6.384 12.384 6.552 ;
  LAYER M1 ;
        RECT 12.352 6.516 12.384 6.588 ;
  LAYER M2 ;
        RECT 12.332 6.536 12.404 6.568 ;
  LAYER M2 ;
        RECT 12.368 6.536 14.96 6.568 ;
  LAYER M1 ;
        RECT 14.944 6.516 14.976 6.588 ;
  LAYER M2 ;
        RECT 14.924 6.536 14.996 6.568 ;
  LAYER M1 ;
        RECT 12.352 9.456 12.384 9.528 ;
  LAYER M2 ;
        RECT 12.332 9.476 12.404 9.508 ;
  LAYER M1 ;
        RECT 12.352 9.492 12.384 9.66 ;
  LAYER M1 ;
        RECT 12.352 9.624 12.384 9.696 ;
  LAYER M2 ;
        RECT 12.332 9.644 12.404 9.676 ;
  LAYER M2 ;
        RECT 12.368 9.644 14.96 9.676 ;
  LAYER M1 ;
        RECT 14.944 9.624 14.976 9.696 ;
  LAYER M2 ;
        RECT 14.924 9.644 14.996 9.676 ;
  LAYER M1 ;
        RECT 12.352 12.564 12.384 12.636 ;
  LAYER M2 ;
        RECT 12.332 12.584 12.404 12.616 ;
  LAYER M1 ;
        RECT 12.352 12.6 12.384 12.768 ;
  LAYER M1 ;
        RECT 12.352 12.732 12.384 12.804 ;
  LAYER M2 ;
        RECT 12.332 12.752 12.404 12.784 ;
  LAYER M2 ;
        RECT 12.368 12.752 14.96 12.784 ;
  LAYER M1 ;
        RECT 14.944 12.732 14.976 12.804 ;
  LAYER M2 ;
        RECT 14.924 12.752 14.996 12.784 ;
  LAYER M1 ;
        RECT 14.944 13.32 14.976 13.392 ;
  LAYER M2 ;
        RECT 14.924 13.34 14.996 13.372 ;
  LAYER M1 ;
        RECT 14.944 12.936 14.976 13.356 ;
  LAYER M1 ;
        RECT 14.944 3.444 14.976 12.936 ;
  LAYER M2 ;
        RECT 0.08 13.34 14.96 13.372 ;
  LAYER M1 ;
        RECT 3.424 3.24 3.456 3.312 ;
  LAYER M2 ;
        RECT 3.404 3.26 3.476 3.292 ;
  LAYER M2 ;
        RECT 0.464 3.26 3.44 3.292 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M2 ;
        RECT 0.464 12.584 3.44 12.616 ;
  LAYER M1 ;
        RECT 0.448 12.564 0.48 12.636 ;
  LAYER M2 ;
        RECT 0.428 12.584 0.5 12.616 ;
  LAYER M1 ;
        RECT 6.4 12.564 6.432 12.636 ;
  LAYER M2 ;
        RECT 6.38 12.584 6.452 12.616 ;
  LAYER M2 ;
        RECT 3.44 12.584 6.416 12.616 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M1 ;
        RECT 9.376 12.564 9.408 12.636 ;
  LAYER M2 ;
        RECT 9.356 12.584 9.428 12.616 ;
  LAYER M2 ;
        RECT 6.416 12.584 9.392 12.616 ;
  LAYER M1 ;
        RECT 6.4 12.564 6.432 12.636 ;
  LAYER M2 ;
        RECT 6.38 12.584 6.452 12.616 ;
  LAYER M1 ;
        RECT 9.376 3.24 9.408 3.312 ;
  LAYER M2 ;
        RECT 9.356 3.26 9.428 3.292 ;
  LAYER M2 ;
        RECT 9.392 3.26 12.368 3.292 ;
  LAYER M1 ;
        RECT 12.352 3.24 12.384 3.312 ;
  LAYER M2 ;
        RECT 12.332 3.26 12.404 3.292 ;
  LAYER M1 ;
        RECT 6.4 3.24 6.432 3.312 ;
  LAYER M2 ;
        RECT 6.38 3.26 6.452 3.292 ;
  LAYER M2 ;
        RECT 6.416 3.26 9.392 3.292 ;
  LAYER M1 ;
        RECT 9.376 3.24 9.408 3.312 ;
  LAYER M2 ;
        RECT 9.356 3.26 9.428 3.292 ;
  LAYER M1 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M3 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M1 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M3 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M1 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M3 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M2 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M1 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M3 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M2 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M1 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M3 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M2 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M1 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M3 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M2 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M1 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M3 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M2 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M1 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M3 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M2 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M1 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M3 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M2 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M1 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M3 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M2 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M1 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M3 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M2 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M1 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M3 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M2 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M1 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M3 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M2 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M1 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M3 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M2 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M1 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M3 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M2 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M1 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M3 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M2 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M1 ;
        RECT 12.304 0.756 14.8 3.36 ;
  LAYER M3 ;
        RECT 12.304 0.756 14.8 3.36 ;
  LAYER M2 ;
        RECT 12.304 0.756 14.8 3.36 ;
  LAYER M1 ;
        RECT 12.304 3.864 14.8 6.468 ;
  LAYER M3 ;
        RECT 12.304 3.864 14.8 6.468 ;
  LAYER M2 ;
        RECT 12.304 3.864 14.8 6.468 ;
  LAYER M1 ;
        RECT 12.304 6.972 14.8 9.576 ;
  LAYER M3 ;
        RECT 12.304 6.972 14.8 9.576 ;
  LAYER M2 ;
        RECT 12.304 6.972 14.8 9.576 ;
  LAYER M1 ;
        RECT 12.304 10.08 14.8 12.684 ;
  LAYER M3 ;
        RECT 12.304 10.08 14.8 12.684 ;
  LAYER M2 ;
        RECT 12.304 10.08 14.8 12.684 ;
  END 
END Cap_60fF
