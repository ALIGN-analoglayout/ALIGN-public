MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 0.3200 BY 0.7560 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.1000 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2200 0.0680 0.2920 0.1000 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.0480 0.0480 0.0800 0.7080 ;
    LAYER M1 ;
      RECT 0.0480 0.6560 0.1440 0.6880 ;
    LAYER M1 ;
      RECT 0.1120 0.0480 0.1440 0.7080 ;
    LAYER M1 ;
      RECT 0.1120 0.0680 0.2080 0.1000 ;
    LAYER M1 ;
      RECT 0.1760 0.0480 0.2080 0.7080 ;
    LAYER M1 ;
      RECT 0.1760 0.6560 0.2720 0.6880 ;
    LAYER M1 ;
      RECT 0.2400 0.0480 0.2720 0.7080 ;
    LAYER V1 ;
      RECT 0.0480 0.0680 0.0800 0.1000 ;
    LAYER V1 ;
      RECT 0.2400 0.0680 0.2720 0.1000 ;
    LAYER boundary ;
      RECT 0.0000 0.0000 0.3200 0.7560 ;
  END
END test
