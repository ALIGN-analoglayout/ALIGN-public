MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 9.36 BY 25.872 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.328 25.584 3.36 25.656 ;
      LAYER M2 ;
        RECT 3.308 25.604 3.38 25.636 ;
      LAYER M1 ;
        RECT 6.304 25.584 6.336 25.656 ;
      LAYER M2 ;
        RECT 6.284 25.604 6.356 25.636 ;
      LAYER M2 ;
        RECT 3.344 25.604 6.32 25.636 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.856 10.128 5.888 10.2 ;
  LAYER M2 ;
        RECT 5.836 10.148 5.908 10.18 ;
  LAYER M2 ;
        RECT 3.056 10.148 5.872 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 5.856 13.236 5.888 13.308 ;
  LAYER M2 ;
        RECT 5.836 13.256 5.908 13.288 ;
  LAYER M2 ;
        RECT 3.056 13.256 5.872 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 5.856 7.02 5.888 7.092 ;
  LAYER M2 ;
        RECT 5.836 7.04 5.908 7.072 ;
  LAYER M2 ;
        RECT 3.056 7.04 5.872 7.072 ;
  LAYER M1 ;
        RECT 3.04 7.02 3.072 7.092 ;
  LAYER M2 ;
        RECT 3.02 7.04 3.092 7.072 ;
  LAYER M1 ;
        RECT 5.856 16.344 5.888 16.416 ;
  LAYER M2 ;
        RECT 5.836 16.364 5.908 16.396 ;
  LAYER M2 ;
        RECT 3.056 16.364 5.872 16.396 ;
  LAYER M1 ;
        RECT 3.04 16.344 3.072 16.416 ;
  LAYER M2 ;
        RECT 3.02 16.364 3.092 16.396 ;
  LAYER M1 ;
        RECT 5.856 3.912 5.888 3.984 ;
  LAYER M2 ;
        RECT 5.836 3.932 5.908 3.964 ;
  LAYER M2 ;
        RECT 3.056 3.932 5.872 3.964 ;
  LAYER M1 ;
        RECT 3.04 3.912 3.072 3.984 ;
  LAYER M2 ;
        RECT 3.02 3.932 3.092 3.964 ;
  LAYER M1 ;
        RECT 5.856 19.452 5.888 19.524 ;
  LAYER M2 ;
        RECT 5.836 19.472 5.908 19.504 ;
  LAYER M2 ;
        RECT 3.056 19.472 5.872 19.504 ;
  LAYER M1 ;
        RECT 3.04 19.452 3.072 19.524 ;
  LAYER M2 ;
        RECT 3.02 19.472 3.092 19.504 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.504 ;
  LAYER M1 ;
        RECT 3.04 0.504 3.072 19.488 ;
  LAYER M1 ;
        RECT 5.856 10.128 5.888 10.2 ;
  LAYER M2 ;
        RECT 5.836 10.148 5.908 10.18 ;
  LAYER M1 ;
        RECT 5.856 9.996 5.888 10.164 ;
  LAYER M1 ;
        RECT 5.856 9.96 5.888 10.032 ;
  LAYER M2 ;
        RECT 5.836 9.98 5.908 10.012 ;
  LAYER M2 ;
        RECT 5.872 9.98 6.032 10.012 ;
  LAYER M1 ;
        RECT 6.016 9.96 6.048 10.032 ;
  LAYER M2 ;
        RECT 5.996 9.98 6.068 10.012 ;
  LAYER M1 ;
        RECT 5.856 13.236 5.888 13.308 ;
  LAYER M2 ;
        RECT 5.836 13.256 5.908 13.288 ;
  LAYER M1 ;
        RECT 5.856 13.104 5.888 13.272 ;
  LAYER M1 ;
        RECT 5.856 13.068 5.888 13.14 ;
  LAYER M2 ;
        RECT 5.836 13.088 5.908 13.12 ;
  LAYER M2 ;
        RECT 5.872 13.088 6.032 13.12 ;
  LAYER M1 ;
        RECT 6.016 13.068 6.048 13.14 ;
  LAYER M2 ;
        RECT 5.996 13.088 6.068 13.12 ;
  LAYER M1 ;
        RECT 5.856 7.02 5.888 7.092 ;
  LAYER M2 ;
        RECT 5.836 7.04 5.908 7.072 ;
  LAYER M1 ;
        RECT 5.856 6.888 5.888 7.056 ;
  LAYER M1 ;
        RECT 5.856 6.852 5.888 6.924 ;
  LAYER M2 ;
        RECT 5.836 6.872 5.908 6.904 ;
  LAYER M2 ;
        RECT 5.872 6.872 6.032 6.904 ;
  LAYER M1 ;
        RECT 6.016 6.852 6.048 6.924 ;
  LAYER M2 ;
        RECT 5.996 6.872 6.068 6.904 ;
  LAYER M1 ;
        RECT 5.856 16.344 5.888 16.416 ;
  LAYER M2 ;
        RECT 5.836 16.364 5.908 16.396 ;
  LAYER M1 ;
        RECT 5.856 16.212 5.888 16.38 ;
  LAYER M1 ;
        RECT 5.856 16.176 5.888 16.248 ;
  LAYER M2 ;
        RECT 5.836 16.196 5.908 16.228 ;
  LAYER M2 ;
        RECT 5.872 16.196 6.032 16.228 ;
  LAYER M1 ;
        RECT 6.016 16.176 6.048 16.248 ;
  LAYER M2 ;
        RECT 5.996 16.196 6.068 16.228 ;
  LAYER M1 ;
        RECT 5.856 3.912 5.888 3.984 ;
  LAYER M2 ;
        RECT 5.836 3.932 5.908 3.964 ;
  LAYER M1 ;
        RECT 5.856 3.78 5.888 3.948 ;
  LAYER M1 ;
        RECT 5.856 3.744 5.888 3.816 ;
  LAYER M2 ;
        RECT 5.836 3.764 5.908 3.796 ;
  LAYER M2 ;
        RECT 5.872 3.764 6.032 3.796 ;
  LAYER M1 ;
        RECT 6.016 3.744 6.048 3.816 ;
  LAYER M2 ;
        RECT 5.996 3.764 6.068 3.796 ;
  LAYER M1 ;
        RECT 5.856 19.452 5.888 19.524 ;
  LAYER M2 ;
        RECT 5.836 19.472 5.908 19.504 ;
  LAYER M1 ;
        RECT 5.856 19.32 5.888 19.488 ;
  LAYER M1 ;
        RECT 5.856 19.284 5.888 19.356 ;
  LAYER M2 ;
        RECT 5.836 19.304 5.908 19.336 ;
  LAYER M2 ;
        RECT 5.872 19.304 6.032 19.336 ;
  LAYER M1 ;
        RECT 6.016 19.284 6.048 19.356 ;
  LAYER M2 ;
        RECT 5.996 19.304 6.068 19.336 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.504 ;
  LAYER M1 ;
        RECT 6.016 0.504 6.048 19.32 ;
  LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
  LAYER M1 ;
        RECT 2.88 0.804 2.912 0.876 ;
  LAYER M2 ;
        RECT 2.86 0.824 2.932 0.856 ;
  LAYER M2 ;
        RECT 0.08 0.824 2.896 0.856 ;
  LAYER M1 ;
        RECT 0.064 0.804 0.096 0.876 ;
  LAYER M2 ;
        RECT 0.044 0.824 0.116 0.856 ;
  LAYER M1 ;
        RECT 2.88 3.912 2.912 3.984 ;
  LAYER M2 ;
        RECT 2.86 3.932 2.932 3.964 ;
  LAYER M2 ;
        RECT 0.08 3.932 2.896 3.964 ;
  LAYER M1 ;
        RECT 0.064 3.912 0.096 3.984 ;
  LAYER M2 ;
        RECT 0.044 3.932 0.116 3.964 ;
  LAYER M1 ;
        RECT 2.88 7.02 2.912 7.092 ;
  LAYER M2 ;
        RECT 2.86 7.04 2.932 7.072 ;
  LAYER M2 ;
        RECT 0.08 7.04 2.896 7.072 ;
  LAYER M1 ;
        RECT 0.064 7.02 0.096 7.092 ;
  LAYER M2 ;
        RECT 0.044 7.04 0.116 7.072 ;
  LAYER M1 ;
        RECT 2.88 10.128 2.912 10.2 ;
  LAYER M2 ;
        RECT 2.86 10.148 2.932 10.18 ;
  LAYER M2 ;
        RECT 0.08 10.148 2.896 10.18 ;
  LAYER M1 ;
        RECT 0.064 10.128 0.096 10.2 ;
  LAYER M2 ;
        RECT 0.044 10.148 0.116 10.18 ;
  LAYER M1 ;
        RECT 2.88 13.236 2.912 13.308 ;
  LAYER M2 ;
        RECT 2.86 13.256 2.932 13.288 ;
  LAYER M2 ;
        RECT 0.08 13.256 2.896 13.288 ;
  LAYER M1 ;
        RECT 0.064 13.236 0.096 13.308 ;
  LAYER M2 ;
        RECT 0.044 13.256 0.116 13.288 ;
  LAYER M1 ;
        RECT 2.88 16.344 2.912 16.416 ;
  LAYER M2 ;
        RECT 2.86 16.364 2.932 16.396 ;
  LAYER M2 ;
        RECT 0.08 16.364 2.896 16.396 ;
  LAYER M1 ;
        RECT 0.064 16.344 0.096 16.416 ;
  LAYER M2 ;
        RECT 0.044 16.364 0.116 16.396 ;
  LAYER M1 ;
        RECT 2.88 19.452 2.912 19.524 ;
  LAYER M2 ;
        RECT 2.86 19.472 2.932 19.504 ;
  LAYER M2 ;
        RECT 0.08 19.472 2.896 19.504 ;
  LAYER M1 ;
        RECT 0.064 19.452 0.096 19.524 ;
  LAYER M2 ;
        RECT 0.044 19.472 0.116 19.504 ;
  LAYER M1 ;
        RECT 2.88 22.56 2.912 22.632 ;
  LAYER M2 ;
        RECT 2.86 22.58 2.932 22.612 ;
  LAYER M2 ;
        RECT 0.08 22.58 2.896 22.612 ;
  LAYER M1 ;
        RECT 0.064 22.56 0.096 22.632 ;
  LAYER M2 ;
        RECT 0.044 22.58 0.116 22.612 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.504 ;
  LAYER M1 ;
        RECT 0.064 0.504 0.096 22.596 ;
  LAYER M1 ;
        RECT 8.832 0.804 8.864 0.876 ;
  LAYER M2 ;
        RECT 8.812 0.824 8.884 0.856 ;
  LAYER M1 ;
        RECT 8.832 0.672 8.864 0.84 ;
  LAYER M1 ;
        RECT 8.832 0.636 8.864 0.708 ;
  LAYER M2 ;
        RECT 8.812 0.656 8.884 0.688 ;
  LAYER M2 ;
        RECT 8.848 0.656 9.008 0.688 ;
  LAYER M1 ;
        RECT 8.992 0.636 9.024 0.708 ;
  LAYER M2 ;
        RECT 8.972 0.656 9.044 0.688 ;
  LAYER M1 ;
        RECT 8.832 3.912 8.864 3.984 ;
  LAYER M2 ;
        RECT 8.812 3.932 8.884 3.964 ;
  LAYER M1 ;
        RECT 8.832 3.78 8.864 3.948 ;
  LAYER M1 ;
        RECT 8.832 3.744 8.864 3.816 ;
  LAYER M2 ;
        RECT 8.812 3.764 8.884 3.796 ;
  LAYER M2 ;
        RECT 8.848 3.764 9.008 3.796 ;
  LAYER M1 ;
        RECT 8.992 3.744 9.024 3.816 ;
  LAYER M2 ;
        RECT 8.972 3.764 9.044 3.796 ;
  LAYER M1 ;
        RECT 8.832 7.02 8.864 7.092 ;
  LAYER M2 ;
        RECT 8.812 7.04 8.884 7.072 ;
  LAYER M1 ;
        RECT 8.832 6.888 8.864 7.056 ;
  LAYER M1 ;
        RECT 8.832 6.852 8.864 6.924 ;
  LAYER M2 ;
        RECT 8.812 6.872 8.884 6.904 ;
  LAYER M2 ;
        RECT 8.848 6.872 9.008 6.904 ;
  LAYER M1 ;
        RECT 8.992 6.852 9.024 6.924 ;
  LAYER M2 ;
        RECT 8.972 6.872 9.044 6.904 ;
  LAYER M1 ;
        RECT 8.832 10.128 8.864 10.2 ;
  LAYER M2 ;
        RECT 8.812 10.148 8.884 10.18 ;
  LAYER M1 ;
        RECT 8.832 9.996 8.864 10.164 ;
  LAYER M1 ;
        RECT 8.832 9.96 8.864 10.032 ;
  LAYER M2 ;
        RECT 8.812 9.98 8.884 10.012 ;
  LAYER M2 ;
        RECT 8.848 9.98 9.008 10.012 ;
  LAYER M1 ;
        RECT 8.992 9.96 9.024 10.032 ;
  LAYER M2 ;
        RECT 8.972 9.98 9.044 10.012 ;
  LAYER M1 ;
        RECT 8.832 13.236 8.864 13.308 ;
  LAYER M2 ;
        RECT 8.812 13.256 8.884 13.288 ;
  LAYER M1 ;
        RECT 8.832 13.104 8.864 13.272 ;
  LAYER M1 ;
        RECT 8.832 13.068 8.864 13.14 ;
  LAYER M2 ;
        RECT 8.812 13.088 8.884 13.12 ;
  LAYER M2 ;
        RECT 8.848 13.088 9.008 13.12 ;
  LAYER M1 ;
        RECT 8.992 13.068 9.024 13.14 ;
  LAYER M2 ;
        RECT 8.972 13.088 9.044 13.12 ;
  LAYER M1 ;
        RECT 8.832 16.344 8.864 16.416 ;
  LAYER M2 ;
        RECT 8.812 16.364 8.884 16.396 ;
  LAYER M1 ;
        RECT 8.832 16.212 8.864 16.38 ;
  LAYER M1 ;
        RECT 8.832 16.176 8.864 16.248 ;
  LAYER M2 ;
        RECT 8.812 16.196 8.884 16.228 ;
  LAYER M2 ;
        RECT 8.848 16.196 9.008 16.228 ;
  LAYER M1 ;
        RECT 8.992 16.176 9.024 16.248 ;
  LAYER M2 ;
        RECT 8.972 16.196 9.044 16.228 ;
  LAYER M1 ;
        RECT 8.832 19.452 8.864 19.524 ;
  LAYER M2 ;
        RECT 8.812 19.472 8.884 19.504 ;
  LAYER M1 ;
        RECT 8.832 19.32 8.864 19.488 ;
  LAYER M1 ;
        RECT 8.832 19.284 8.864 19.356 ;
  LAYER M2 ;
        RECT 8.812 19.304 8.884 19.336 ;
  LAYER M2 ;
        RECT 8.848 19.304 9.008 19.336 ;
  LAYER M1 ;
        RECT 8.992 19.284 9.024 19.356 ;
  LAYER M2 ;
        RECT 8.972 19.304 9.044 19.336 ;
  LAYER M1 ;
        RECT 8.832 22.56 8.864 22.632 ;
  LAYER M2 ;
        RECT 8.812 22.58 8.884 22.612 ;
  LAYER M1 ;
        RECT 8.832 22.428 8.864 22.596 ;
  LAYER M1 ;
        RECT 8.832 22.392 8.864 22.464 ;
  LAYER M2 ;
        RECT 8.812 22.412 8.884 22.444 ;
  LAYER M2 ;
        RECT 8.848 22.412 9.008 22.444 ;
  LAYER M1 ;
        RECT 8.992 22.392 9.024 22.464 ;
  LAYER M2 ;
        RECT 8.972 22.412 9.044 22.444 ;
  LAYER M1 ;
        RECT 8.992 0.048 9.024 0.12 ;
  LAYER M2 ;
        RECT 8.972 0.068 9.044 0.1 ;
  LAYER M1 ;
        RECT 8.992 0.084 9.024 0.504 ;
  LAYER M1 ;
        RECT 8.992 0.504 9.024 22.428 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.008 0.1 ;
  LAYER M1 ;
        RECT 5.856 0.804 5.888 0.876 ;
  LAYER M2 ;
        RECT 5.836 0.824 5.908 0.856 ;
  LAYER M2 ;
        RECT 2.896 0.824 5.872 0.856 ;
  LAYER M1 ;
        RECT 2.88 0.804 2.912 0.876 ;
  LAYER M2 ;
        RECT 2.86 0.824 2.932 0.856 ;
  LAYER M1 ;
        RECT 5.856 22.56 5.888 22.632 ;
  LAYER M2 ;
        RECT 5.836 22.58 5.908 22.612 ;
  LAYER M2 ;
        RECT 2.896 22.58 5.872 22.612 ;
  LAYER M1 ;
        RECT 2.88 22.56 2.912 22.632 ;
  LAYER M2 ;
        RECT 2.86 22.58 2.932 22.612 ;
  LAYER M1 ;
        RECT 3.488 12.564 3.52 12.636 ;
  LAYER M2 ;
        RECT 3.468 12.584 3.54 12.616 ;
  LAYER M2 ;
        RECT 3.344 12.584 3.504 12.616 ;
  LAYER M1 ;
        RECT 3.328 12.564 3.36 12.636 ;
  LAYER M2 ;
        RECT 3.308 12.584 3.38 12.616 ;
  LAYER M1 ;
        RECT 3.488 15.672 3.52 15.744 ;
  LAYER M2 ;
        RECT 3.468 15.692 3.54 15.724 ;
  LAYER M2 ;
        RECT 3.344 15.692 3.504 15.724 ;
  LAYER M1 ;
        RECT 3.328 15.672 3.36 15.744 ;
  LAYER M2 ;
        RECT 3.308 15.692 3.38 15.724 ;
  LAYER M1 ;
        RECT 3.488 9.456 3.52 9.528 ;
  LAYER M2 ;
        RECT 3.468 9.476 3.54 9.508 ;
  LAYER M2 ;
        RECT 3.344 9.476 3.504 9.508 ;
  LAYER M1 ;
        RECT 3.328 9.456 3.36 9.528 ;
  LAYER M2 ;
        RECT 3.308 9.476 3.38 9.508 ;
  LAYER M1 ;
        RECT 3.488 18.78 3.52 18.852 ;
  LAYER M2 ;
        RECT 3.468 18.8 3.54 18.832 ;
  LAYER M2 ;
        RECT 3.344 18.8 3.504 18.832 ;
  LAYER M1 ;
        RECT 3.328 18.78 3.36 18.852 ;
  LAYER M2 ;
        RECT 3.308 18.8 3.38 18.832 ;
  LAYER M1 ;
        RECT 3.488 6.348 3.52 6.42 ;
  LAYER M2 ;
        RECT 3.468 6.368 3.54 6.4 ;
  LAYER M2 ;
        RECT 3.344 6.368 3.504 6.4 ;
  LAYER M1 ;
        RECT 3.328 6.348 3.36 6.42 ;
  LAYER M2 ;
        RECT 3.308 6.368 3.38 6.4 ;
  LAYER M1 ;
        RECT 3.488 21.888 3.52 21.96 ;
  LAYER M2 ;
        RECT 3.468 21.908 3.54 21.94 ;
  LAYER M2 ;
        RECT 3.344 21.908 3.504 21.94 ;
  LAYER M1 ;
        RECT 3.328 21.888 3.36 21.96 ;
  LAYER M2 ;
        RECT 3.308 21.908 3.38 21.94 ;
  LAYER M1 ;
        RECT 3.328 25.584 3.36 25.656 ;
  LAYER M2 ;
        RECT 3.308 25.604 3.38 25.636 ;
  LAYER M1 ;
        RECT 3.328 25.368 3.36 25.62 ;
  LAYER M1 ;
        RECT 3.328 6.384 3.36 25.368 ;
  LAYER M1 ;
        RECT 3.488 12.564 3.52 12.636 ;
  LAYER M2 ;
        RECT 3.468 12.584 3.54 12.616 ;
  LAYER M1 ;
        RECT 3.488 12.6 3.52 12.768 ;
  LAYER M1 ;
        RECT 3.488 12.732 3.52 12.804 ;
  LAYER M2 ;
        RECT 3.468 12.752 3.54 12.784 ;
  LAYER M2 ;
        RECT 3.504 12.752 6.32 12.784 ;
  LAYER M1 ;
        RECT 6.304 12.732 6.336 12.804 ;
  LAYER M2 ;
        RECT 6.284 12.752 6.356 12.784 ;
  LAYER M1 ;
        RECT 3.488 15.672 3.52 15.744 ;
  LAYER M2 ;
        RECT 3.468 15.692 3.54 15.724 ;
  LAYER M1 ;
        RECT 3.488 15.708 3.52 15.876 ;
  LAYER M1 ;
        RECT 3.488 15.84 3.52 15.912 ;
  LAYER M2 ;
        RECT 3.468 15.86 3.54 15.892 ;
  LAYER M2 ;
        RECT 3.504 15.86 6.32 15.892 ;
  LAYER M1 ;
        RECT 6.304 15.84 6.336 15.912 ;
  LAYER M2 ;
        RECT 6.284 15.86 6.356 15.892 ;
  LAYER M1 ;
        RECT 3.488 9.456 3.52 9.528 ;
  LAYER M2 ;
        RECT 3.468 9.476 3.54 9.508 ;
  LAYER M1 ;
        RECT 3.488 9.492 3.52 9.66 ;
  LAYER M1 ;
        RECT 3.488 9.624 3.52 9.696 ;
  LAYER M2 ;
        RECT 3.468 9.644 3.54 9.676 ;
  LAYER M2 ;
        RECT 3.504 9.644 6.32 9.676 ;
  LAYER M1 ;
        RECT 6.304 9.624 6.336 9.696 ;
  LAYER M2 ;
        RECT 6.284 9.644 6.356 9.676 ;
  LAYER M1 ;
        RECT 3.488 18.78 3.52 18.852 ;
  LAYER M2 ;
        RECT 3.468 18.8 3.54 18.832 ;
  LAYER M1 ;
        RECT 3.488 18.816 3.52 18.984 ;
  LAYER M1 ;
        RECT 3.488 18.948 3.52 19.02 ;
  LAYER M2 ;
        RECT 3.468 18.968 3.54 19 ;
  LAYER M2 ;
        RECT 3.504 18.968 6.32 19 ;
  LAYER M1 ;
        RECT 6.304 18.948 6.336 19.02 ;
  LAYER M2 ;
        RECT 6.284 18.968 6.356 19 ;
  LAYER M1 ;
        RECT 3.488 6.348 3.52 6.42 ;
  LAYER M2 ;
        RECT 3.468 6.368 3.54 6.4 ;
  LAYER M1 ;
        RECT 3.488 6.384 3.52 6.552 ;
  LAYER M1 ;
        RECT 3.488 6.516 3.52 6.588 ;
  LAYER M2 ;
        RECT 3.468 6.536 3.54 6.568 ;
  LAYER M2 ;
        RECT 3.504 6.536 6.32 6.568 ;
  LAYER M1 ;
        RECT 6.304 6.516 6.336 6.588 ;
  LAYER M2 ;
        RECT 6.284 6.536 6.356 6.568 ;
  LAYER M1 ;
        RECT 3.488 21.888 3.52 21.96 ;
  LAYER M2 ;
        RECT 3.468 21.908 3.54 21.94 ;
  LAYER M1 ;
        RECT 3.488 21.924 3.52 22.092 ;
  LAYER M1 ;
        RECT 3.488 22.056 3.52 22.128 ;
  LAYER M2 ;
        RECT 3.468 22.076 3.54 22.108 ;
  LAYER M2 ;
        RECT 3.504 22.076 6.32 22.108 ;
  LAYER M1 ;
        RECT 6.304 22.056 6.336 22.128 ;
  LAYER M2 ;
        RECT 6.284 22.076 6.356 22.108 ;
  LAYER M1 ;
        RECT 6.304 25.584 6.336 25.656 ;
  LAYER M2 ;
        RECT 6.284 25.604 6.356 25.636 ;
  LAYER M1 ;
        RECT 6.304 25.368 6.336 25.62 ;
  LAYER M1 ;
        RECT 6.304 6.552 6.336 25.368 ;
  LAYER M2 ;
        RECT 3.344 25.604 6.32 25.636 ;
  LAYER M1 ;
        RECT 0.512 3.24 0.544 3.312 ;
  LAYER M2 ;
        RECT 0.492 3.26 0.564 3.292 ;
  LAYER M2 ;
        RECT 0.368 3.26 0.528 3.292 ;
  LAYER M1 ;
        RECT 0.352 3.24 0.384 3.312 ;
  LAYER M2 ;
        RECT 0.332 3.26 0.404 3.292 ;
  LAYER M1 ;
        RECT 0.512 6.348 0.544 6.42 ;
  LAYER M2 ;
        RECT 0.492 6.368 0.564 6.4 ;
  LAYER M2 ;
        RECT 0.368 6.368 0.528 6.4 ;
  LAYER M1 ;
        RECT 0.352 6.348 0.384 6.42 ;
  LAYER M2 ;
        RECT 0.332 6.368 0.404 6.4 ;
  LAYER M1 ;
        RECT 0.512 9.456 0.544 9.528 ;
  LAYER M2 ;
        RECT 0.492 9.476 0.564 9.508 ;
  LAYER M2 ;
        RECT 0.368 9.476 0.528 9.508 ;
  LAYER M1 ;
        RECT 0.352 9.456 0.384 9.528 ;
  LAYER M2 ;
        RECT 0.332 9.476 0.404 9.508 ;
  LAYER M1 ;
        RECT 0.512 12.564 0.544 12.636 ;
  LAYER M2 ;
        RECT 0.492 12.584 0.564 12.616 ;
  LAYER M2 ;
        RECT 0.368 12.584 0.528 12.616 ;
  LAYER M1 ;
        RECT 0.352 12.564 0.384 12.636 ;
  LAYER M2 ;
        RECT 0.332 12.584 0.404 12.616 ;
  LAYER M1 ;
        RECT 0.512 15.672 0.544 15.744 ;
  LAYER M2 ;
        RECT 0.492 15.692 0.564 15.724 ;
  LAYER M2 ;
        RECT 0.368 15.692 0.528 15.724 ;
  LAYER M1 ;
        RECT 0.352 15.672 0.384 15.744 ;
  LAYER M2 ;
        RECT 0.332 15.692 0.404 15.724 ;
  LAYER M1 ;
        RECT 0.512 18.78 0.544 18.852 ;
  LAYER M2 ;
        RECT 0.492 18.8 0.564 18.832 ;
  LAYER M2 ;
        RECT 0.368 18.8 0.528 18.832 ;
  LAYER M1 ;
        RECT 0.352 18.78 0.384 18.852 ;
  LAYER M2 ;
        RECT 0.332 18.8 0.404 18.832 ;
  LAYER M1 ;
        RECT 0.512 21.888 0.544 21.96 ;
  LAYER M2 ;
        RECT 0.492 21.908 0.564 21.94 ;
  LAYER M2 ;
        RECT 0.368 21.908 0.528 21.94 ;
  LAYER M1 ;
        RECT 0.352 21.888 0.384 21.96 ;
  LAYER M2 ;
        RECT 0.332 21.908 0.404 21.94 ;
  LAYER M1 ;
        RECT 0.512 24.996 0.544 25.068 ;
  LAYER M2 ;
        RECT 0.492 25.016 0.564 25.048 ;
  LAYER M2 ;
        RECT 0.368 25.016 0.528 25.048 ;
  LAYER M1 ;
        RECT 0.352 24.996 0.384 25.068 ;
  LAYER M2 ;
        RECT 0.332 25.016 0.404 25.048 ;
  LAYER M1 ;
        RECT 0.352 25.752 0.384 25.824 ;
  LAYER M2 ;
        RECT 0.332 25.772 0.404 25.804 ;
  LAYER M1 ;
        RECT 0.352 25.368 0.384 25.788 ;
  LAYER M1 ;
        RECT 0.352 3.276 0.384 25.368 ;
  LAYER M1 ;
        RECT 6.464 3.24 6.496 3.312 ;
  LAYER M2 ;
        RECT 6.444 3.26 6.516 3.292 ;
  LAYER M1 ;
        RECT 6.464 3.276 6.496 3.444 ;
  LAYER M1 ;
        RECT 6.464 3.408 6.496 3.48 ;
  LAYER M2 ;
        RECT 6.444 3.428 6.516 3.46 ;
  LAYER M2 ;
        RECT 6.48 3.428 9.296 3.46 ;
  LAYER M1 ;
        RECT 9.28 3.408 9.312 3.48 ;
  LAYER M2 ;
        RECT 9.26 3.428 9.332 3.46 ;
  LAYER M1 ;
        RECT 6.464 6.348 6.496 6.42 ;
  LAYER M2 ;
        RECT 6.444 6.368 6.516 6.4 ;
  LAYER M1 ;
        RECT 6.464 6.384 6.496 6.552 ;
  LAYER M1 ;
        RECT 6.464 6.516 6.496 6.588 ;
  LAYER M2 ;
        RECT 6.444 6.536 6.516 6.568 ;
  LAYER M2 ;
        RECT 6.48 6.536 9.296 6.568 ;
  LAYER M1 ;
        RECT 9.28 6.516 9.312 6.588 ;
  LAYER M2 ;
        RECT 9.26 6.536 9.332 6.568 ;
  LAYER M1 ;
        RECT 6.464 9.456 6.496 9.528 ;
  LAYER M2 ;
        RECT 6.444 9.476 6.516 9.508 ;
  LAYER M1 ;
        RECT 6.464 9.492 6.496 9.66 ;
  LAYER M1 ;
        RECT 6.464 9.624 6.496 9.696 ;
  LAYER M2 ;
        RECT 6.444 9.644 6.516 9.676 ;
  LAYER M2 ;
        RECT 6.48 9.644 9.296 9.676 ;
  LAYER M1 ;
        RECT 9.28 9.624 9.312 9.696 ;
  LAYER M2 ;
        RECT 9.26 9.644 9.332 9.676 ;
  LAYER M1 ;
        RECT 6.464 12.564 6.496 12.636 ;
  LAYER M2 ;
        RECT 6.444 12.584 6.516 12.616 ;
  LAYER M1 ;
        RECT 6.464 12.6 6.496 12.768 ;
  LAYER M1 ;
        RECT 6.464 12.732 6.496 12.804 ;
  LAYER M2 ;
        RECT 6.444 12.752 6.516 12.784 ;
  LAYER M2 ;
        RECT 6.48 12.752 9.296 12.784 ;
  LAYER M1 ;
        RECT 9.28 12.732 9.312 12.804 ;
  LAYER M2 ;
        RECT 9.26 12.752 9.332 12.784 ;
  LAYER M1 ;
        RECT 6.464 15.672 6.496 15.744 ;
  LAYER M2 ;
        RECT 6.444 15.692 6.516 15.724 ;
  LAYER M1 ;
        RECT 6.464 15.708 6.496 15.876 ;
  LAYER M1 ;
        RECT 6.464 15.84 6.496 15.912 ;
  LAYER M2 ;
        RECT 6.444 15.86 6.516 15.892 ;
  LAYER M2 ;
        RECT 6.48 15.86 9.296 15.892 ;
  LAYER M1 ;
        RECT 9.28 15.84 9.312 15.912 ;
  LAYER M2 ;
        RECT 9.26 15.86 9.332 15.892 ;
  LAYER M1 ;
        RECT 6.464 18.78 6.496 18.852 ;
  LAYER M2 ;
        RECT 6.444 18.8 6.516 18.832 ;
  LAYER M1 ;
        RECT 6.464 18.816 6.496 18.984 ;
  LAYER M1 ;
        RECT 6.464 18.948 6.496 19.02 ;
  LAYER M2 ;
        RECT 6.444 18.968 6.516 19 ;
  LAYER M2 ;
        RECT 6.48 18.968 9.296 19 ;
  LAYER M1 ;
        RECT 9.28 18.948 9.312 19.02 ;
  LAYER M2 ;
        RECT 9.26 18.968 9.332 19 ;
  LAYER M1 ;
        RECT 6.464 21.888 6.496 21.96 ;
  LAYER M2 ;
        RECT 6.444 21.908 6.516 21.94 ;
  LAYER M1 ;
        RECT 6.464 21.924 6.496 22.092 ;
  LAYER M1 ;
        RECT 6.464 22.056 6.496 22.128 ;
  LAYER M2 ;
        RECT 6.444 22.076 6.516 22.108 ;
  LAYER M2 ;
        RECT 6.48 22.076 9.296 22.108 ;
  LAYER M1 ;
        RECT 9.28 22.056 9.312 22.128 ;
  LAYER M2 ;
        RECT 9.26 22.076 9.332 22.108 ;
  LAYER M1 ;
        RECT 6.464 24.996 6.496 25.068 ;
  LAYER M2 ;
        RECT 6.444 25.016 6.516 25.048 ;
  LAYER M1 ;
        RECT 6.464 25.032 6.496 25.2 ;
  LAYER M1 ;
        RECT 6.464 25.164 6.496 25.236 ;
  LAYER M2 ;
        RECT 6.444 25.184 6.516 25.216 ;
  LAYER M2 ;
        RECT 6.48 25.184 9.296 25.216 ;
  LAYER M1 ;
        RECT 9.28 25.164 9.312 25.236 ;
  LAYER M2 ;
        RECT 9.26 25.184 9.332 25.216 ;
  LAYER M1 ;
        RECT 9.28 25.752 9.312 25.824 ;
  LAYER M2 ;
        RECT 9.26 25.772 9.332 25.804 ;
  LAYER M1 ;
        RECT 9.28 25.368 9.312 25.788 ;
  LAYER M1 ;
        RECT 9.28 3.444 9.312 25.368 ;
  LAYER M2 ;
        RECT 0.368 25.772 9.296 25.804 ;
  LAYER M1 ;
        RECT 3.488 3.24 3.52 3.312 ;
  LAYER M2 ;
        RECT 3.468 3.26 3.54 3.292 ;
  LAYER M2 ;
        RECT 0.528 3.26 3.504 3.292 ;
  LAYER M1 ;
        RECT 0.512 3.24 0.544 3.312 ;
  LAYER M2 ;
        RECT 0.492 3.26 0.564 3.292 ;
  LAYER M1 ;
        RECT 3.488 24.996 3.52 25.068 ;
  LAYER M2 ;
        RECT 3.468 25.016 3.54 25.048 ;
  LAYER M2 ;
        RECT 0.528 25.016 3.504 25.048 ;
  LAYER M1 ;
        RECT 0.512 24.996 0.544 25.068 ;
  LAYER M2 ;
        RECT 0.492 25.016 0.564 25.048 ;
  LAYER M1 ;
        RECT 0.464 0.756 2.96 3.36 ;
  LAYER M3 ;
        RECT 0.464 0.756 2.96 3.36 ;
  LAYER M2 ;
        RECT 0.464 0.756 2.96 3.36 ;
  LAYER M1 ;
        RECT 0.464 3.864 2.96 6.468 ;
  LAYER M3 ;
        RECT 0.464 3.864 2.96 6.468 ;
  LAYER M2 ;
        RECT 0.464 3.864 2.96 6.468 ;
  LAYER M1 ;
        RECT 0.464 6.972 2.96 9.576 ;
  LAYER M3 ;
        RECT 0.464 6.972 2.96 9.576 ;
  LAYER M2 ;
        RECT 0.464 6.972 2.96 9.576 ;
  LAYER M1 ;
        RECT 0.464 10.08 2.96 12.684 ;
  LAYER M3 ;
        RECT 0.464 10.08 2.96 12.684 ;
  LAYER M2 ;
        RECT 0.464 10.08 2.96 12.684 ;
  LAYER M1 ;
        RECT 0.464 13.188 2.96 15.792 ;
  LAYER M3 ;
        RECT 0.464 13.188 2.96 15.792 ;
  LAYER M2 ;
        RECT 0.464 13.188 2.96 15.792 ;
  LAYER M1 ;
        RECT 0.464 16.296 2.96 18.9 ;
  LAYER M3 ;
        RECT 0.464 16.296 2.96 18.9 ;
  LAYER M2 ;
        RECT 0.464 16.296 2.96 18.9 ;
  LAYER M1 ;
        RECT 0.464 19.404 2.96 22.008 ;
  LAYER M3 ;
        RECT 0.464 19.404 2.96 22.008 ;
  LAYER M2 ;
        RECT 0.464 19.404 2.96 22.008 ;
  LAYER M1 ;
        RECT 0.464 22.512 2.96 25.116 ;
  LAYER M3 ;
        RECT 0.464 22.512 2.96 25.116 ;
  LAYER M2 ;
        RECT 0.464 22.512 2.96 25.116 ;
  LAYER M1 ;
        RECT 3.44 0.756 5.936 3.36 ;
  LAYER M3 ;
        RECT 3.44 0.756 5.936 3.36 ;
  LAYER M2 ;
        RECT 3.44 0.756 5.936 3.36 ;
  LAYER M1 ;
        RECT 3.44 3.864 5.936 6.468 ;
  LAYER M3 ;
        RECT 3.44 3.864 5.936 6.468 ;
  LAYER M2 ;
        RECT 3.44 3.864 5.936 6.468 ;
  LAYER M1 ;
        RECT 3.44 6.972 5.936 9.576 ;
  LAYER M3 ;
        RECT 3.44 6.972 5.936 9.576 ;
  LAYER M2 ;
        RECT 3.44 6.972 5.936 9.576 ;
  LAYER M1 ;
        RECT 3.44 10.08 5.936 12.684 ;
  LAYER M3 ;
        RECT 3.44 10.08 5.936 12.684 ;
  LAYER M2 ;
        RECT 3.44 10.08 5.936 12.684 ;
  LAYER M1 ;
        RECT 3.44 13.188 5.936 15.792 ;
  LAYER M3 ;
        RECT 3.44 13.188 5.936 15.792 ;
  LAYER M2 ;
        RECT 3.44 13.188 5.936 15.792 ;
  LAYER M1 ;
        RECT 3.44 16.296 5.936 18.9 ;
  LAYER M3 ;
        RECT 3.44 16.296 5.936 18.9 ;
  LAYER M2 ;
        RECT 3.44 16.296 5.936 18.9 ;
  LAYER M1 ;
        RECT 3.44 19.404 5.936 22.008 ;
  LAYER M3 ;
        RECT 3.44 19.404 5.936 22.008 ;
  LAYER M2 ;
        RECT 3.44 19.404 5.936 22.008 ;
  LAYER M1 ;
        RECT 3.44 22.512 5.936 25.116 ;
  LAYER M3 ;
        RECT 3.44 22.512 5.936 25.116 ;
  LAYER M2 ;
        RECT 3.44 22.512 5.936 25.116 ;
  LAYER M1 ;
        RECT 6.416 0.756 8.912 3.36 ;
  LAYER M3 ;
        RECT 6.416 0.756 8.912 3.36 ;
  LAYER M2 ;
        RECT 6.416 0.756 8.912 3.36 ;
  LAYER M1 ;
        RECT 6.416 3.864 8.912 6.468 ;
  LAYER M3 ;
        RECT 6.416 3.864 8.912 6.468 ;
  LAYER M2 ;
        RECT 6.416 3.864 8.912 6.468 ;
  LAYER M1 ;
        RECT 6.416 6.972 8.912 9.576 ;
  LAYER M3 ;
        RECT 6.416 6.972 8.912 9.576 ;
  LAYER M2 ;
        RECT 6.416 6.972 8.912 9.576 ;
  LAYER M1 ;
        RECT 6.416 10.08 8.912 12.684 ;
  LAYER M3 ;
        RECT 6.416 10.08 8.912 12.684 ;
  LAYER M2 ;
        RECT 6.416 10.08 8.912 12.684 ;
  LAYER M1 ;
        RECT 6.416 13.188 8.912 15.792 ;
  LAYER M3 ;
        RECT 6.416 13.188 8.912 15.792 ;
  LAYER M2 ;
        RECT 6.416 13.188 8.912 15.792 ;
  LAYER M1 ;
        RECT 6.416 16.296 8.912 18.9 ;
  LAYER M3 ;
        RECT 6.416 16.296 8.912 18.9 ;
  LAYER M2 ;
        RECT 6.416 16.296 8.912 18.9 ;
  LAYER M1 ;
        RECT 6.416 19.404 8.912 22.008 ;
  LAYER M3 ;
        RECT 6.416 19.404 8.912 22.008 ;
  LAYER M2 ;
        RECT 6.416 19.404 8.912 22.008 ;
  LAYER M1 ;
        RECT 6.416 22.512 8.912 25.116 ;
  LAYER M3 ;
        RECT 6.416 22.512 8.912 25.116 ;
  LAYER M2 ;
        RECT 6.416 22.512 8.912 25.116 ;
  END 
END Cap_60fF
