MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 16.64 BY 18.984 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.624 18.528 6.656 18.6 ;
      LAYER M2 ;
        RECT 6.604 18.548 6.676 18.58 ;
      LAYER M1 ;
        RECT 10.144 18.528 10.176 18.6 ;
      LAYER M2 ;
        RECT 10.124 18.548 10.196 18.58 ;
      LAYER M2 ;
        RECT 6.64 18.548 10.16 18.58 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.144 0.384 6.176 0.456 ;
      LAYER M2 ;
        RECT 6.124 0.404 6.196 0.436 ;
      LAYER M1 ;
        RECT 9.664 0.384 9.696 0.456 ;
      LAYER M2 ;
        RECT 9.644 0.404 9.716 0.436 ;
      LAYER M2 ;
        RECT 6.16 0.404 9.68 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.784 18.696 6.816 18.768 ;
      LAYER M2 ;
        RECT 6.764 18.716 6.836 18.748 ;
      LAYER M1 ;
        RECT 10.304 18.696 10.336 18.768 ;
      LAYER M2 ;
        RECT 10.284 18.716 10.356 18.748 ;
      LAYER M2 ;
        RECT 6.8 18.716 10.32 18.748 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.304 0.216 6.336 0.288 ;
      LAYER M2 ;
        RECT 6.284 0.236 6.356 0.268 ;
      LAYER M1 ;
        RECT 9.824 0.216 9.856 0.288 ;
      LAYER M2 ;
        RECT 9.804 0.236 9.876 0.268 ;
      LAYER M2 ;
        RECT 6.32 0.236 9.84 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 7.104 6.768 7.136 6.84 ;
  LAYER M2 ;
        RECT 7.084 6.788 7.156 6.82 ;
  LAYER M2 ;
        RECT 6.16 6.788 7.12 6.82 ;
  LAYER M1 ;
        RECT 6.144 6.768 6.176 6.84 ;
  LAYER M2 ;
        RECT 6.124 6.788 6.196 6.82 ;
  LAYER M1 ;
        RECT 3.584 12.648 3.616 12.72 ;
  LAYER M2 ;
        RECT 3.564 12.668 3.636 12.7 ;
  LAYER M1 ;
        RECT 3.584 12.516 3.616 12.684 ;
  LAYER M1 ;
        RECT 3.584 12.48 3.616 12.552 ;
  LAYER M2 ;
        RECT 3.564 12.5 3.636 12.532 ;
  LAYER M2 ;
        RECT 3.6 12.5 6.16 12.532 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 12.552 ;
  LAYER M2 ;
        RECT 6.124 12.5 6.196 12.532 ;
  LAYER M1 ;
        RECT 6.144 0.384 6.176 0.456 ;
  LAYER M2 ;
        RECT 6.124 0.404 6.196 0.436 ;
  LAYER M1 ;
        RECT 6.144 0.42 6.176 0.588 ;
  LAYER M1 ;
        RECT 6.144 0.588 6.176 12.516 ;
  LAYER M1 ;
        RECT 10.624 3.828 10.656 3.9 ;
  LAYER M2 ;
        RECT 10.604 3.848 10.676 3.88 ;
  LAYER M2 ;
        RECT 9.68 3.848 10.64 3.88 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 3.9 ;
  LAYER M2 ;
        RECT 9.644 3.848 9.716 3.88 ;
  LAYER M1 ;
        RECT 9.664 0.384 9.696 0.456 ;
  LAYER M2 ;
        RECT 9.644 0.404 9.716 0.436 ;
  LAYER M1 ;
        RECT 9.664 0.42 9.696 0.588 ;
  LAYER M1 ;
        RECT 9.664 0.588 9.696 3.864 ;
  LAYER M2 ;
        RECT 6.16 0.404 9.68 0.436 ;
  LAYER M1 ;
        RECT 3.584 6.768 3.616 6.84 ;
  LAYER M2 ;
        RECT 3.564 6.788 3.636 6.82 ;
  LAYER M1 ;
        RECT 3.584 6.636 3.616 6.804 ;
  LAYER M1 ;
        RECT 3.584 6.6 3.616 6.672 ;
  LAYER M2 ;
        RECT 3.564 6.62 3.636 6.652 ;
  LAYER M2 ;
        RECT 3.6 6.62 6.32 6.652 ;
  LAYER M1 ;
        RECT 6.304 6.6 6.336 6.672 ;
  LAYER M2 ;
        RECT 6.284 6.62 6.356 6.652 ;
  LAYER M1 ;
        RECT 3.584 9.708 3.616 9.78 ;
  LAYER M2 ;
        RECT 3.564 9.728 3.636 9.76 ;
  LAYER M1 ;
        RECT 3.584 9.576 3.616 9.744 ;
  LAYER M1 ;
        RECT 3.584 9.54 3.616 9.612 ;
  LAYER M2 ;
        RECT 3.564 9.56 3.636 9.592 ;
  LAYER M2 ;
        RECT 3.6 9.56 6.32 9.592 ;
  LAYER M1 ;
        RECT 6.304 9.54 6.336 9.612 ;
  LAYER M2 ;
        RECT 6.284 9.56 6.356 9.592 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 3.9 ;
  LAYER M2 ;
        RECT 7.084 3.848 7.156 3.88 ;
  LAYER M2 ;
        RECT 6.32 3.848 7.12 3.88 ;
  LAYER M1 ;
        RECT 6.304 3.828 6.336 3.9 ;
  LAYER M2 ;
        RECT 6.284 3.848 6.356 3.88 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 12.72 ;
  LAYER M2 ;
        RECT 7.084 12.668 7.156 12.7 ;
  LAYER M2 ;
        RECT 6.32 12.668 7.12 12.7 ;
  LAYER M1 ;
        RECT 6.304 12.648 6.336 12.72 ;
  LAYER M2 ;
        RECT 6.284 12.668 6.356 12.7 ;
  LAYER M1 ;
        RECT 6.304 0.216 6.336 0.288 ;
  LAYER M2 ;
        RECT 6.284 0.236 6.356 0.268 ;
  LAYER M1 ;
        RECT 6.304 0.252 6.336 0.588 ;
  LAYER M1 ;
        RECT 6.304 0.588 6.336 12.684 ;
  LAYER M1 ;
        RECT 10.624 9.708 10.656 9.78 ;
  LAYER M2 ;
        RECT 10.604 9.728 10.676 9.76 ;
  LAYER M2 ;
        RECT 9.84 9.728 10.64 9.76 ;
  LAYER M1 ;
        RECT 9.824 9.708 9.856 9.78 ;
  LAYER M2 ;
        RECT 9.804 9.728 9.876 9.76 ;
  LAYER M1 ;
        RECT 10.624 6.768 10.656 6.84 ;
  LAYER M2 ;
        RECT 10.604 6.788 10.676 6.82 ;
  LAYER M2 ;
        RECT 9.84 6.788 10.64 6.82 ;
  LAYER M1 ;
        RECT 9.824 6.768 9.856 6.84 ;
  LAYER M2 ;
        RECT 9.804 6.788 9.876 6.82 ;
  LAYER M1 ;
        RECT 9.824 0.216 9.856 0.288 ;
  LAYER M2 ;
        RECT 9.804 0.236 9.876 0.268 ;
  LAYER M1 ;
        RECT 9.824 0.252 9.856 0.588 ;
  LAYER M1 ;
        RECT 9.824 0.588 9.856 9.744 ;
  LAYER M2 ;
        RECT 6.32 0.236 9.84 0.268 ;
  LAYER M1 ;
        RECT 3.584 0.888 3.616 0.96 ;
  LAYER M2 ;
        RECT 3.564 0.908 3.636 0.94 ;
  LAYER M1 ;
        RECT 3.584 0.756 3.616 0.924 ;
  LAYER M1 ;
        RECT 3.584 0.72 3.616 0.792 ;
  LAYER M2 ;
        RECT 3.564 0.74 3.636 0.772 ;
  LAYER M2 ;
        RECT 3.6 0.74 6.48 0.772 ;
  LAYER M1 ;
        RECT 6.464 0.72 6.496 0.792 ;
  LAYER M2 ;
        RECT 6.444 0.74 6.516 0.772 ;
  LAYER M1 ;
        RECT 3.584 3.828 3.616 3.9 ;
  LAYER M2 ;
        RECT 3.564 3.848 3.636 3.88 ;
  LAYER M1 ;
        RECT 3.584 3.696 3.616 3.864 ;
  LAYER M1 ;
        RECT 3.584 3.66 3.616 3.732 ;
  LAYER M2 ;
        RECT 3.564 3.68 3.636 3.712 ;
  LAYER M2 ;
        RECT 3.6 3.68 6.48 3.712 ;
  LAYER M1 ;
        RECT 6.464 3.66 6.496 3.732 ;
  LAYER M2 ;
        RECT 6.444 3.68 6.516 3.712 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 15.66 ;
  LAYER M2 ;
        RECT 3.564 15.608 3.636 15.64 ;
  LAYER M1 ;
        RECT 3.584 15.456 3.616 15.624 ;
  LAYER M1 ;
        RECT 3.584 15.42 3.616 15.492 ;
  LAYER M2 ;
        RECT 3.564 15.44 3.636 15.472 ;
  LAYER M2 ;
        RECT 3.6 15.44 6.48 15.472 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 15.492 ;
  LAYER M2 ;
        RECT 6.444 15.44 6.516 15.472 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 0.96 ;
  LAYER M2 ;
        RECT 7.084 0.908 7.156 0.94 ;
  LAYER M2 ;
        RECT 6.48 0.908 7.12 0.94 ;
  LAYER M1 ;
        RECT 6.464 0.888 6.496 0.96 ;
  LAYER M2 ;
        RECT 6.444 0.908 6.516 0.94 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 9.78 ;
  LAYER M2 ;
        RECT 7.084 9.728 7.156 9.76 ;
  LAYER M2 ;
        RECT 6.48 9.728 7.12 9.76 ;
  LAYER M1 ;
        RECT 6.464 9.708 6.496 9.78 ;
  LAYER M2 ;
        RECT 6.444 9.728 6.516 9.76 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 15.66 ;
  LAYER M2 ;
        RECT 7.084 15.608 7.156 15.64 ;
  LAYER M2 ;
        RECT 6.48 15.608 7.12 15.64 ;
  LAYER M1 ;
        RECT 6.464 15.588 6.496 15.66 ;
  LAYER M2 ;
        RECT 6.444 15.608 6.516 15.64 ;
  LAYER M1 ;
        RECT 6.464 0.048 6.496 0.12 ;
  LAYER M2 ;
        RECT 6.444 0.068 6.516 0.1 ;
  LAYER M1 ;
        RECT 6.464 0.084 6.496 0.588 ;
  LAYER M1 ;
        RECT 6.464 0.588 6.496 15.624 ;
  LAYER M1 ;
        RECT 10.624 0.888 10.656 0.96 ;
  LAYER M2 ;
        RECT 10.604 0.908 10.676 0.94 ;
  LAYER M2 ;
        RECT 10 0.908 10.64 0.94 ;
  LAYER M1 ;
        RECT 9.984 0.888 10.016 0.96 ;
  LAYER M2 ;
        RECT 9.964 0.908 10.036 0.94 ;
  LAYER M1 ;
        RECT 10.624 12.648 10.656 12.72 ;
  LAYER M2 ;
        RECT 10.604 12.668 10.676 12.7 ;
  LAYER M2 ;
        RECT 10 12.668 10.64 12.7 ;
  LAYER M1 ;
        RECT 9.984 12.648 10.016 12.72 ;
  LAYER M2 ;
        RECT 9.964 12.668 10.036 12.7 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 15.66 ;
  LAYER M2 ;
        RECT 10.604 15.608 10.676 15.64 ;
  LAYER M2 ;
        RECT 10 15.608 10.64 15.64 ;
  LAYER M1 ;
        RECT 9.984 15.588 10.016 15.66 ;
  LAYER M2 ;
        RECT 9.964 15.608 10.036 15.64 ;
  LAYER M1 ;
        RECT 9.984 0.048 10.016 0.12 ;
  LAYER M2 ;
        RECT 9.964 0.068 10.036 0.1 ;
  LAYER M1 ;
        RECT 9.984 0.084 10.016 0.588 ;
  LAYER M1 ;
        RECT 9.984 0.588 10.016 15.624 ;
  LAYER M2 ;
        RECT 6.48 0.068 10 0.1 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M2 ;
        RECT 0.08 15.608 3.6 15.64 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 15.66 ;
  LAYER M2 ;
        RECT 3.564 15.608 3.636 15.64 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.684 0.096 15.624 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.744 0.096 12.684 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.804 0.096 9.744 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.864 0.096 6.804 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.924 0.096 3.864 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 14.144 15.588 14.176 15.66 ;
  LAYER M2 ;
        RECT 14.124 15.608 14.196 15.64 ;
  LAYER M2 ;
        RECT 10.64 15.608 14.16 15.64 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 15.66 ;
  LAYER M2 ;
        RECT 10.604 15.608 10.676 15.64 ;
  LAYER M1 ;
        RECT 14.144 12.648 14.176 12.72 ;
  LAYER M2 ;
        RECT 14.124 12.668 14.196 12.7 ;
  LAYER M2 ;
        RECT 10.64 12.668 14.16 12.7 ;
  LAYER M1 ;
        RECT 10.624 12.648 10.656 12.72 ;
  LAYER M2 ;
        RECT 10.604 12.668 10.676 12.7 ;
  LAYER M1 ;
        RECT 14.144 9.708 14.176 9.78 ;
  LAYER M2 ;
        RECT 14.124 9.728 14.196 9.76 ;
  LAYER M1 ;
        RECT 14.144 9.744 14.176 12.684 ;
  LAYER M1 ;
        RECT 14.144 12.648 14.176 12.72 ;
  LAYER M2 ;
        RECT 14.124 12.668 14.196 12.7 ;
  LAYER M1 ;
        RECT 14.144 6.768 14.176 6.84 ;
  LAYER M2 ;
        RECT 14.124 6.788 14.196 6.82 ;
  LAYER M1 ;
        RECT 14.144 6.804 14.176 9.744 ;
  LAYER M1 ;
        RECT 14.144 9.708 14.176 9.78 ;
  LAYER M2 ;
        RECT 14.124 9.728 14.196 9.76 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 3.9 ;
  LAYER M2 ;
        RECT 14.124 3.848 14.196 3.88 ;
  LAYER M1 ;
        RECT 14.144 3.864 14.176 6.804 ;
  LAYER M1 ;
        RECT 14.144 6.768 14.176 6.84 ;
  LAYER M2 ;
        RECT 14.124 6.788 14.196 6.82 ;
  LAYER M1 ;
        RECT 14.144 0.888 14.176 0.96 ;
  LAYER M2 ;
        RECT 14.124 0.908 14.196 0.94 ;
  LAYER M1 ;
        RECT 14.144 0.924 14.176 3.864 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 3.9 ;
  LAYER M2 ;
        RECT 14.124 3.848 14.196 3.88 ;
  LAYER M1 ;
        RECT 9.504 9.204 9.536 9.276 ;
  LAYER M2 ;
        RECT 9.484 9.224 9.556 9.256 ;
  LAYER M2 ;
        RECT 6.64 9.224 9.52 9.256 ;
  LAYER M1 ;
        RECT 6.624 9.204 6.656 9.276 ;
  LAYER M2 ;
        RECT 6.604 9.224 6.676 9.256 ;
  LAYER M1 ;
        RECT 5.984 15.084 6.016 15.156 ;
  LAYER M2 ;
        RECT 5.964 15.104 6.036 15.136 ;
  LAYER M1 ;
        RECT 5.984 15.12 6.016 15.288 ;
  LAYER M1 ;
        RECT 5.984 15.252 6.016 15.324 ;
  LAYER M2 ;
        RECT 5.964 15.272 6.036 15.304 ;
  LAYER M2 ;
        RECT 6 15.272 6.64 15.304 ;
  LAYER M1 ;
        RECT 6.624 15.252 6.656 15.324 ;
  LAYER M2 ;
        RECT 6.604 15.272 6.676 15.304 ;
  LAYER M1 ;
        RECT 6.624 18.528 6.656 18.6 ;
  LAYER M2 ;
        RECT 6.604 18.548 6.676 18.58 ;
  LAYER M1 ;
        RECT 6.624 18.396 6.656 18.564 ;
  LAYER M1 ;
        RECT 6.624 9.24 6.656 18.396 ;
  LAYER M1 ;
        RECT 13.024 6.264 13.056 6.336 ;
  LAYER M2 ;
        RECT 13.004 6.284 13.076 6.316 ;
  LAYER M2 ;
        RECT 10.16 6.284 13.04 6.316 ;
  LAYER M1 ;
        RECT 10.144 6.264 10.176 6.336 ;
  LAYER M2 ;
        RECT 10.124 6.284 10.196 6.316 ;
  LAYER M1 ;
        RECT 10.144 18.528 10.176 18.6 ;
  LAYER M2 ;
        RECT 10.124 18.548 10.196 18.58 ;
  LAYER M1 ;
        RECT 10.144 18.396 10.176 18.564 ;
  LAYER M1 ;
        RECT 10.144 6.3 10.176 18.396 ;
  LAYER M2 ;
        RECT 6.64 18.548 10.16 18.58 ;
  LAYER M1 ;
        RECT 5.984 9.204 6.016 9.276 ;
  LAYER M2 ;
        RECT 5.964 9.224 6.036 9.256 ;
  LAYER M1 ;
        RECT 5.984 9.24 6.016 9.408 ;
  LAYER M1 ;
        RECT 5.984 9.372 6.016 9.444 ;
  LAYER M2 ;
        RECT 5.964 9.392 6.036 9.424 ;
  LAYER M2 ;
        RECT 6 9.392 6.8 9.424 ;
  LAYER M1 ;
        RECT 6.784 9.372 6.816 9.444 ;
  LAYER M2 ;
        RECT 6.764 9.392 6.836 9.424 ;
  LAYER M1 ;
        RECT 5.984 12.144 6.016 12.216 ;
  LAYER M2 ;
        RECT 5.964 12.164 6.036 12.196 ;
  LAYER M1 ;
        RECT 5.984 12.18 6.016 12.348 ;
  LAYER M1 ;
        RECT 5.984 12.312 6.016 12.384 ;
  LAYER M2 ;
        RECT 5.964 12.332 6.036 12.364 ;
  LAYER M2 ;
        RECT 6 12.332 6.8 12.364 ;
  LAYER M1 ;
        RECT 6.784 12.312 6.816 12.384 ;
  LAYER M2 ;
        RECT 6.764 12.332 6.836 12.364 ;
  LAYER M1 ;
        RECT 9.504 6.264 9.536 6.336 ;
  LAYER M2 ;
        RECT 9.484 6.284 9.556 6.316 ;
  LAYER M2 ;
        RECT 6.8 6.284 9.52 6.316 ;
  LAYER M1 ;
        RECT 6.784 6.264 6.816 6.336 ;
  LAYER M2 ;
        RECT 6.764 6.284 6.836 6.316 ;
  LAYER M1 ;
        RECT 9.504 15.084 9.536 15.156 ;
  LAYER M2 ;
        RECT 9.484 15.104 9.556 15.136 ;
  LAYER M2 ;
        RECT 6.8 15.104 9.52 15.136 ;
  LAYER M1 ;
        RECT 6.784 15.084 6.816 15.156 ;
  LAYER M2 ;
        RECT 6.764 15.104 6.836 15.136 ;
  LAYER M1 ;
        RECT 6.784 18.696 6.816 18.768 ;
  LAYER M2 ;
        RECT 6.764 18.716 6.836 18.748 ;
  LAYER M1 ;
        RECT 6.784 18.396 6.816 18.732 ;
  LAYER M1 ;
        RECT 6.784 6.3 6.816 18.396 ;
  LAYER M1 ;
        RECT 13.024 12.144 13.056 12.216 ;
  LAYER M2 ;
        RECT 13.004 12.164 13.076 12.196 ;
  LAYER M2 ;
        RECT 10.32 12.164 13.04 12.196 ;
  LAYER M1 ;
        RECT 10.304 12.144 10.336 12.216 ;
  LAYER M2 ;
        RECT 10.284 12.164 10.356 12.196 ;
  LAYER M1 ;
        RECT 13.024 9.204 13.056 9.276 ;
  LAYER M2 ;
        RECT 13.004 9.224 13.076 9.256 ;
  LAYER M2 ;
        RECT 10.32 9.224 13.04 9.256 ;
  LAYER M1 ;
        RECT 10.304 9.204 10.336 9.276 ;
  LAYER M2 ;
        RECT 10.284 9.224 10.356 9.256 ;
  LAYER M1 ;
        RECT 10.304 18.696 10.336 18.768 ;
  LAYER M2 ;
        RECT 10.284 18.716 10.356 18.748 ;
  LAYER M1 ;
        RECT 10.304 18.396 10.336 18.732 ;
  LAYER M1 ;
        RECT 10.304 9.24 10.336 18.396 ;
  LAYER M2 ;
        RECT 6.8 18.716 10.32 18.748 ;
  LAYER M1 ;
        RECT 5.984 3.324 6.016 3.396 ;
  LAYER M2 ;
        RECT 5.964 3.344 6.036 3.376 ;
  LAYER M1 ;
        RECT 5.984 3.36 6.016 3.528 ;
  LAYER M1 ;
        RECT 5.984 3.492 6.016 3.564 ;
  LAYER M2 ;
        RECT 5.964 3.512 6.036 3.544 ;
  LAYER M2 ;
        RECT 6 3.512 6.96 3.544 ;
  LAYER M1 ;
        RECT 6.944 3.492 6.976 3.564 ;
  LAYER M2 ;
        RECT 6.924 3.512 6.996 3.544 ;
  LAYER M1 ;
        RECT 5.984 6.264 6.016 6.336 ;
  LAYER M2 ;
        RECT 5.964 6.284 6.036 6.316 ;
  LAYER M1 ;
        RECT 5.984 6.3 6.016 6.468 ;
  LAYER M1 ;
        RECT 5.984 6.432 6.016 6.504 ;
  LAYER M2 ;
        RECT 5.964 6.452 6.036 6.484 ;
  LAYER M2 ;
        RECT 6 6.452 6.96 6.484 ;
  LAYER M1 ;
        RECT 6.944 6.432 6.976 6.504 ;
  LAYER M2 ;
        RECT 6.924 6.452 6.996 6.484 ;
  LAYER M1 ;
        RECT 5.984 18.024 6.016 18.096 ;
  LAYER M2 ;
        RECT 5.964 18.044 6.036 18.076 ;
  LAYER M1 ;
        RECT 5.984 18.06 6.016 18.228 ;
  LAYER M1 ;
        RECT 5.984 18.192 6.016 18.264 ;
  LAYER M2 ;
        RECT 5.964 18.212 6.036 18.244 ;
  LAYER M2 ;
        RECT 6 18.212 6.96 18.244 ;
  LAYER M1 ;
        RECT 6.944 18.192 6.976 18.264 ;
  LAYER M2 ;
        RECT 6.924 18.212 6.996 18.244 ;
  LAYER M1 ;
        RECT 9.504 3.324 9.536 3.396 ;
  LAYER M2 ;
        RECT 9.484 3.344 9.556 3.376 ;
  LAYER M2 ;
        RECT 6.96 3.344 9.52 3.376 ;
  LAYER M1 ;
        RECT 6.944 3.324 6.976 3.396 ;
  LAYER M2 ;
        RECT 6.924 3.344 6.996 3.376 ;
  LAYER M1 ;
        RECT 9.504 12.144 9.536 12.216 ;
  LAYER M2 ;
        RECT 9.484 12.164 9.556 12.196 ;
  LAYER M2 ;
        RECT 6.96 12.164 9.52 12.196 ;
  LAYER M1 ;
        RECT 6.944 12.144 6.976 12.216 ;
  LAYER M2 ;
        RECT 6.924 12.164 6.996 12.196 ;
  LAYER M1 ;
        RECT 9.504 18.024 9.536 18.096 ;
  LAYER M2 ;
        RECT 9.484 18.044 9.556 18.076 ;
  LAYER M2 ;
        RECT 6.96 18.044 9.52 18.076 ;
  LAYER M1 ;
        RECT 6.944 18.024 6.976 18.096 ;
  LAYER M2 ;
        RECT 6.924 18.044 6.996 18.076 ;
  LAYER M1 ;
        RECT 6.944 18.864 6.976 18.936 ;
  LAYER M2 ;
        RECT 6.924 18.884 6.996 18.916 ;
  LAYER M1 ;
        RECT 6.944 18.396 6.976 18.9 ;
  LAYER M1 ;
        RECT 6.944 3.36 6.976 18.396 ;
  LAYER M1 ;
        RECT 13.024 3.324 13.056 3.396 ;
  LAYER M2 ;
        RECT 13.004 3.344 13.076 3.376 ;
  LAYER M2 ;
        RECT 10.48 3.344 13.04 3.376 ;
  LAYER M1 ;
        RECT 10.464 3.324 10.496 3.396 ;
  LAYER M2 ;
        RECT 10.444 3.344 10.516 3.376 ;
  LAYER M1 ;
        RECT 13.024 15.084 13.056 15.156 ;
  LAYER M2 ;
        RECT 13.004 15.104 13.076 15.136 ;
  LAYER M2 ;
        RECT 10.48 15.104 13.04 15.136 ;
  LAYER M1 ;
        RECT 10.464 15.084 10.496 15.156 ;
  LAYER M2 ;
        RECT 10.444 15.104 10.516 15.136 ;
  LAYER M1 ;
        RECT 13.024 18.024 13.056 18.096 ;
  LAYER M2 ;
        RECT 13.004 18.044 13.076 18.076 ;
  LAYER M2 ;
        RECT 10.48 18.044 13.04 18.076 ;
  LAYER M1 ;
        RECT 10.464 18.024 10.496 18.096 ;
  LAYER M2 ;
        RECT 10.444 18.044 10.516 18.076 ;
  LAYER M1 ;
        RECT 10.464 18.864 10.496 18.936 ;
  LAYER M2 ;
        RECT 10.444 18.884 10.516 18.916 ;
  LAYER M1 ;
        RECT 10.464 18.396 10.496 18.9 ;
  LAYER M1 ;
        RECT 10.464 3.36 10.496 18.396 ;
  LAYER M2 ;
        RECT 6.96 18.884 10.48 18.916 ;
  LAYER M1 ;
        RECT 2.464 18.024 2.496 18.096 ;
  LAYER M2 ;
        RECT 2.444 18.044 2.516 18.076 ;
  LAYER M2 ;
        RECT 2.48 18.044 6 18.076 ;
  LAYER M1 ;
        RECT 5.984 18.024 6.016 18.096 ;
  LAYER M2 ;
        RECT 5.964 18.044 6.036 18.076 ;
  LAYER M1 ;
        RECT 2.464 15.084 2.496 15.156 ;
  LAYER M2 ;
        RECT 2.444 15.104 2.516 15.136 ;
  LAYER M1 ;
        RECT 2.464 15.12 2.496 18.06 ;
  LAYER M1 ;
        RECT 2.464 18.024 2.496 18.096 ;
  LAYER M2 ;
        RECT 2.444 18.044 2.516 18.076 ;
  LAYER M1 ;
        RECT 2.464 12.144 2.496 12.216 ;
  LAYER M2 ;
        RECT 2.444 12.164 2.516 12.196 ;
  LAYER M1 ;
        RECT 2.464 12.18 2.496 15.12 ;
  LAYER M1 ;
        RECT 2.464 15.084 2.496 15.156 ;
  LAYER M2 ;
        RECT 2.444 15.104 2.516 15.136 ;
  LAYER M1 ;
        RECT 2.464 9.204 2.496 9.276 ;
  LAYER M2 ;
        RECT 2.444 9.224 2.516 9.256 ;
  LAYER M1 ;
        RECT 2.464 9.24 2.496 12.18 ;
  LAYER M1 ;
        RECT 2.464 12.144 2.496 12.216 ;
  LAYER M2 ;
        RECT 2.444 12.164 2.516 12.196 ;
  LAYER M1 ;
        RECT 2.464 6.264 2.496 6.336 ;
  LAYER M2 ;
        RECT 2.444 6.284 2.516 6.316 ;
  LAYER M1 ;
        RECT 2.464 6.3 2.496 9.24 ;
  LAYER M1 ;
        RECT 2.464 9.204 2.496 9.276 ;
  LAYER M2 ;
        RECT 2.444 9.224 2.516 9.256 ;
  LAYER M1 ;
        RECT 2.464 3.324 2.496 3.396 ;
  LAYER M2 ;
        RECT 2.444 3.344 2.516 3.376 ;
  LAYER M1 ;
        RECT 2.464 3.36 2.496 6.3 ;
  LAYER M1 ;
        RECT 2.464 6.264 2.496 6.336 ;
  LAYER M2 ;
        RECT 2.444 6.284 2.516 6.316 ;
  LAYER M1 ;
        RECT 16.544 18.024 16.576 18.096 ;
  LAYER M2 ;
        RECT 16.524 18.044 16.596 18.076 ;
  LAYER M2 ;
        RECT 13.04 18.044 16.56 18.076 ;
  LAYER M1 ;
        RECT 13.024 18.024 13.056 18.096 ;
  LAYER M2 ;
        RECT 13.004 18.044 13.076 18.076 ;
  LAYER M1 ;
        RECT 16.544 15.084 16.576 15.156 ;
  LAYER M2 ;
        RECT 16.524 15.104 16.596 15.136 ;
  LAYER M2 ;
        RECT 13.04 15.104 16.56 15.136 ;
  LAYER M1 ;
        RECT 13.024 15.084 13.056 15.156 ;
  LAYER M2 ;
        RECT 13.004 15.104 13.076 15.136 ;
  LAYER M1 ;
        RECT 16.544 12.144 16.576 12.216 ;
  LAYER M2 ;
        RECT 16.524 12.164 16.596 12.196 ;
  LAYER M1 ;
        RECT 16.544 12.18 16.576 15.12 ;
  LAYER M1 ;
        RECT 16.544 15.084 16.576 15.156 ;
  LAYER M2 ;
        RECT 16.524 15.104 16.596 15.136 ;
  LAYER M1 ;
        RECT 16.544 9.204 16.576 9.276 ;
  LAYER M2 ;
        RECT 16.524 9.224 16.596 9.256 ;
  LAYER M1 ;
        RECT 16.544 9.24 16.576 12.18 ;
  LAYER M1 ;
        RECT 16.544 12.144 16.576 12.216 ;
  LAYER M2 ;
        RECT 16.524 12.164 16.596 12.196 ;
  LAYER M1 ;
        RECT 16.544 6.264 16.576 6.336 ;
  LAYER M2 ;
        RECT 16.524 6.284 16.596 6.316 ;
  LAYER M1 ;
        RECT 16.544 6.3 16.576 9.24 ;
  LAYER M1 ;
        RECT 16.544 9.204 16.576 9.276 ;
  LAYER M2 ;
        RECT 16.524 9.224 16.596 9.256 ;
  LAYER M1 ;
        RECT 16.544 3.324 16.576 3.396 ;
  LAYER M2 ;
        RECT 16.524 3.344 16.596 3.376 ;
  LAYER M1 ;
        RECT 16.544 3.36 16.576 6.3 ;
  LAYER M1 ;
        RECT 16.544 6.264 16.576 6.336 ;
  LAYER M2 ;
        RECT 16.524 6.284 16.596 6.316 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 3.396 ;
  LAYER M1 ;
        RECT 0.128 0.888 0.16 3.396 ;
  LAYER M1 ;
        RECT 0.192 0.888 0.224 3.396 ;
  LAYER M1 ;
        RECT 0.256 0.888 0.288 3.396 ;
  LAYER M1 ;
        RECT 0.32 0.888 0.352 3.396 ;
  LAYER M1 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M1 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M1 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M1 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M1 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M1 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M1 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M1 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M1 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M1 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M1 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M1 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M1 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M1 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M1 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M1 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M1 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M1 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M1 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M1 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M1 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M1 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M1 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M1 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M1 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M1 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M1 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M1 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M1 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M1 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M1 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M2 ;
        RECT 0.044 0.972 2.516 1.004 ;
  LAYER M2 ;
        RECT 0.044 1.036 2.516 1.068 ;
  LAYER M2 ;
        RECT 0.044 1.1 2.516 1.132 ;
  LAYER M2 ;
        RECT 0.044 1.164 2.516 1.196 ;
  LAYER M2 ;
        RECT 0.044 1.228 2.516 1.26 ;
  LAYER M2 ;
        RECT 0.044 1.292 2.516 1.324 ;
  LAYER M2 ;
        RECT 0.044 1.356 2.516 1.388 ;
  LAYER M2 ;
        RECT 0.044 1.42 2.516 1.452 ;
  LAYER M2 ;
        RECT 0.044 1.484 2.516 1.516 ;
  LAYER M2 ;
        RECT 0.044 1.548 2.516 1.58 ;
  LAYER M2 ;
        RECT 0.044 1.612 2.516 1.644 ;
  LAYER M2 ;
        RECT 0.044 1.676 2.516 1.708 ;
  LAYER M2 ;
        RECT 0.044 1.74 2.516 1.772 ;
  LAYER M2 ;
        RECT 0.044 1.804 2.516 1.836 ;
  LAYER M2 ;
        RECT 0.044 1.868 2.516 1.9 ;
  LAYER M2 ;
        RECT 0.044 1.932 2.516 1.964 ;
  LAYER M2 ;
        RECT 0.044 1.996 2.516 2.028 ;
  LAYER M2 ;
        RECT 0.044 2.06 2.516 2.092 ;
  LAYER M2 ;
        RECT 0.044 2.124 2.516 2.156 ;
  LAYER M2 ;
        RECT 0.044 2.188 2.516 2.22 ;
  LAYER M2 ;
        RECT 0.044 2.252 2.516 2.284 ;
  LAYER M2 ;
        RECT 0.044 2.316 2.516 2.348 ;
  LAYER M2 ;
        RECT 0.044 2.38 2.516 2.412 ;
  LAYER M2 ;
        RECT 0.044 2.444 2.516 2.476 ;
  LAYER M2 ;
        RECT 0.044 2.508 2.516 2.54 ;
  LAYER M2 ;
        RECT 0.044 2.572 2.516 2.604 ;
  LAYER M2 ;
        RECT 0.044 2.636 2.516 2.668 ;
  LAYER M2 ;
        RECT 0.044 2.7 2.516 2.732 ;
  LAYER M2 ;
        RECT 0.044 2.764 2.516 2.796 ;
  LAYER M2 ;
        RECT 0.044 2.828 2.516 2.86 ;
  LAYER M2 ;
        RECT 0.044 2.892 2.516 2.924 ;
  LAYER M2 ;
        RECT 0.044 2.956 2.516 2.988 ;
  LAYER M2 ;
        RECT 0.044 3.02 2.516 3.052 ;
  LAYER M2 ;
        RECT 0.044 3.084 2.516 3.116 ;
  LAYER M2 ;
        RECT 0.044 3.148 2.516 3.18 ;
  LAYER M2 ;
        RECT 0.044 3.212 2.516 3.244 ;
  LAYER M3 ;
        RECT 0.064 0.888 0.096 3.396 ;
  LAYER M3 ;
        RECT 0.128 0.888 0.16 3.396 ;
  LAYER M3 ;
        RECT 0.192 0.888 0.224 3.396 ;
  LAYER M3 ;
        RECT 0.256 0.888 0.288 3.396 ;
  LAYER M3 ;
        RECT 0.32 0.888 0.352 3.396 ;
  LAYER M3 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M3 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M3 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M3 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M3 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M3 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M3 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M3 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M3 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M3 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M3 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M3 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M3 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M3 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M3 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M3 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M3 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M3 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M3 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M3 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M3 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M3 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M3 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M3 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M3 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M3 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M3 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M3 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M3 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M3 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M3 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M3 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M3 ;
        RECT 2.464 0.888 2.496 3.396 ;
  LAYER M1 ;
        RECT 0.079 0.924 0.081 3.36 ;
  LAYER M1 ;
        RECT 0.159 0.924 0.161 3.36 ;
  LAYER M1 ;
        RECT 0.239 0.924 0.241 3.36 ;
  LAYER M1 ;
        RECT 0.319 0.924 0.321 3.36 ;
  LAYER M1 ;
        RECT 0.399 0.924 0.401 3.36 ;
  LAYER M1 ;
        RECT 0.479 0.924 0.481 3.36 ;
  LAYER M1 ;
        RECT 0.559 0.924 0.561 3.36 ;
  LAYER M1 ;
        RECT 0.639 0.924 0.641 3.36 ;
  LAYER M1 ;
        RECT 0.719 0.924 0.721 3.36 ;
  LAYER M1 ;
        RECT 0.799 0.924 0.801 3.36 ;
  LAYER M1 ;
        RECT 0.879 0.924 0.881 3.36 ;
  LAYER M1 ;
        RECT 0.959 0.924 0.961 3.36 ;
  LAYER M1 ;
        RECT 1.039 0.924 1.041 3.36 ;
  LAYER M1 ;
        RECT 1.119 0.924 1.121 3.36 ;
  LAYER M1 ;
        RECT 1.199 0.924 1.201 3.36 ;
  LAYER M1 ;
        RECT 1.279 0.924 1.281 3.36 ;
  LAYER M1 ;
        RECT 1.359 0.924 1.361 3.36 ;
  LAYER M1 ;
        RECT 1.439 0.924 1.441 3.36 ;
  LAYER M1 ;
        RECT 1.519 0.924 1.521 3.36 ;
  LAYER M1 ;
        RECT 1.599 0.924 1.601 3.36 ;
  LAYER M1 ;
        RECT 1.679 0.924 1.681 3.36 ;
  LAYER M1 ;
        RECT 1.759 0.924 1.761 3.36 ;
  LAYER M1 ;
        RECT 1.839 0.924 1.841 3.36 ;
  LAYER M1 ;
        RECT 1.919 0.924 1.921 3.36 ;
  LAYER M1 ;
        RECT 1.999 0.924 2.001 3.36 ;
  LAYER M1 ;
        RECT 2.079 0.924 2.081 3.36 ;
  LAYER M1 ;
        RECT 2.159 0.924 2.161 3.36 ;
  LAYER M1 ;
        RECT 2.239 0.924 2.241 3.36 ;
  LAYER M1 ;
        RECT 2.319 0.924 2.321 3.36 ;
  LAYER M1 ;
        RECT 2.399 0.924 2.401 3.36 ;
  LAYER M2 ;
        RECT 0.08 0.923 2.48 0.925 ;
  LAYER M2 ;
        RECT 0.08 1.007 2.48 1.009 ;
  LAYER M2 ;
        RECT 0.08 1.091 2.48 1.093 ;
  LAYER M2 ;
        RECT 0.08 1.175 2.48 1.177 ;
  LAYER M2 ;
        RECT 0.08 1.259 2.48 1.261 ;
  LAYER M2 ;
        RECT 0.08 1.343 2.48 1.345 ;
  LAYER M2 ;
        RECT 0.08 1.427 2.48 1.429 ;
  LAYER M2 ;
        RECT 0.08 1.511 2.48 1.513 ;
  LAYER M2 ;
        RECT 0.08 1.595 2.48 1.597 ;
  LAYER M2 ;
        RECT 0.08 1.679 2.48 1.681 ;
  LAYER M2 ;
        RECT 0.08 1.763 2.48 1.765 ;
  LAYER M2 ;
        RECT 0.08 1.847 2.48 1.849 ;
  LAYER M2 ;
        RECT 0.08 1.9305 2.48 1.9325 ;
  LAYER M2 ;
        RECT 0.08 2.015 2.48 2.017 ;
  LAYER M2 ;
        RECT 0.08 2.099 2.48 2.101 ;
  LAYER M2 ;
        RECT 0.08 2.183 2.48 2.185 ;
  LAYER M2 ;
        RECT 0.08 2.267 2.48 2.269 ;
  LAYER M2 ;
        RECT 0.08 2.351 2.48 2.353 ;
  LAYER M2 ;
        RECT 0.08 2.435 2.48 2.437 ;
  LAYER M2 ;
        RECT 0.08 2.519 2.48 2.521 ;
  LAYER M2 ;
        RECT 0.08 2.603 2.48 2.605 ;
  LAYER M2 ;
        RECT 0.08 2.687 2.48 2.689 ;
  LAYER M2 ;
        RECT 0.08 2.771 2.48 2.773 ;
  LAYER M2 ;
        RECT 0.08 2.855 2.48 2.857 ;
  LAYER M2 ;
        RECT 0.08 2.939 2.48 2.941 ;
  LAYER M2 ;
        RECT 0.08 3.023 2.48 3.025 ;
  LAYER M2 ;
        RECT 0.08 3.107 2.48 3.109 ;
  LAYER M2 ;
        RECT 0.08 3.191 2.48 3.193 ;
  LAYER M2 ;
        RECT 0.08 3.275 2.48 3.277 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 6.336 ;
  LAYER M1 ;
        RECT 0.128 3.828 0.16 6.336 ;
  LAYER M1 ;
        RECT 0.192 3.828 0.224 6.336 ;
  LAYER M1 ;
        RECT 0.256 3.828 0.288 6.336 ;
  LAYER M1 ;
        RECT 0.32 3.828 0.352 6.336 ;
  LAYER M1 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M1 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M1 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M1 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M1 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M1 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M1 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M1 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M1 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M1 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M1 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M1 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M1 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M1 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M1 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M1 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M1 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M1 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M1 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M1 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M1 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M1 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M1 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M1 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M1 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M1 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M1 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M1 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M1 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M1 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M1 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M1 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M2 ;
        RECT 0.044 3.912 2.516 3.944 ;
  LAYER M2 ;
        RECT 0.044 3.976 2.516 4.008 ;
  LAYER M2 ;
        RECT 0.044 4.04 2.516 4.072 ;
  LAYER M2 ;
        RECT 0.044 4.104 2.516 4.136 ;
  LAYER M2 ;
        RECT 0.044 4.168 2.516 4.2 ;
  LAYER M2 ;
        RECT 0.044 4.232 2.516 4.264 ;
  LAYER M2 ;
        RECT 0.044 4.296 2.516 4.328 ;
  LAYER M2 ;
        RECT 0.044 4.36 2.516 4.392 ;
  LAYER M2 ;
        RECT 0.044 4.424 2.516 4.456 ;
  LAYER M2 ;
        RECT 0.044 4.488 2.516 4.52 ;
  LAYER M2 ;
        RECT 0.044 4.552 2.516 4.584 ;
  LAYER M2 ;
        RECT 0.044 4.616 2.516 4.648 ;
  LAYER M2 ;
        RECT 0.044 4.68 2.516 4.712 ;
  LAYER M2 ;
        RECT 0.044 4.744 2.516 4.776 ;
  LAYER M2 ;
        RECT 0.044 4.808 2.516 4.84 ;
  LAYER M2 ;
        RECT 0.044 4.872 2.516 4.904 ;
  LAYER M2 ;
        RECT 0.044 4.936 2.516 4.968 ;
  LAYER M2 ;
        RECT 0.044 5 2.516 5.032 ;
  LAYER M2 ;
        RECT 0.044 5.064 2.516 5.096 ;
  LAYER M2 ;
        RECT 0.044 5.128 2.516 5.16 ;
  LAYER M2 ;
        RECT 0.044 5.192 2.516 5.224 ;
  LAYER M2 ;
        RECT 0.044 5.256 2.516 5.288 ;
  LAYER M2 ;
        RECT 0.044 5.32 2.516 5.352 ;
  LAYER M2 ;
        RECT 0.044 5.384 2.516 5.416 ;
  LAYER M2 ;
        RECT 0.044 5.448 2.516 5.48 ;
  LAYER M2 ;
        RECT 0.044 5.512 2.516 5.544 ;
  LAYER M2 ;
        RECT 0.044 5.576 2.516 5.608 ;
  LAYER M2 ;
        RECT 0.044 5.64 2.516 5.672 ;
  LAYER M2 ;
        RECT 0.044 5.704 2.516 5.736 ;
  LAYER M2 ;
        RECT 0.044 5.768 2.516 5.8 ;
  LAYER M2 ;
        RECT 0.044 5.832 2.516 5.864 ;
  LAYER M2 ;
        RECT 0.044 5.896 2.516 5.928 ;
  LAYER M2 ;
        RECT 0.044 5.96 2.516 5.992 ;
  LAYER M2 ;
        RECT 0.044 6.024 2.516 6.056 ;
  LAYER M2 ;
        RECT 0.044 6.088 2.516 6.12 ;
  LAYER M2 ;
        RECT 0.044 6.152 2.516 6.184 ;
  LAYER M3 ;
        RECT 0.064 3.828 0.096 6.336 ;
  LAYER M3 ;
        RECT 0.128 3.828 0.16 6.336 ;
  LAYER M3 ;
        RECT 0.192 3.828 0.224 6.336 ;
  LAYER M3 ;
        RECT 0.256 3.828 0.288 6.336 ;
  LAYER M3 ;
        RECT 0.32 3.828 0.352 6.336 ;
  LAYER M3 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M3 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M3 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M3 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M3 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M3 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M3 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M3 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M3 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M3 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M3 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M3 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M3 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M3 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M3 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M3 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M3 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M3 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M3 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M3 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M3 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M3 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M3 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M3 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M3 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M3 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M3 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M3 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M3 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M3 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M3 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M3 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M3 ;
        RECT 2.464 3.828 2.496 6.336 ;
  LAYER M1 ;
        RECT 0.079 3.864 0.081 6.3 ;
  LAYER M1 ;
        RECT 0.159 3.864 0.161 6.3 ;
  LAYER M1 ;
        RECT 0.239 3.864 0.241 6.3 ;
  LAYER M1 ;
        RECT 0.319 3.864 0.321 6.3 ;
  LAYER M1 ;
        RECT 0.399 3.864 0.401 6.3 ;
  LAYER M1 ;
        RECT 0.479 3.864 0.481 6.3 ;
  LAYER M1 ;
        RECT 0.559 3.864 0.561 6.3 ;
  LAYER M1 ;
        RECT 0.639 3.864 0.641 6.3 ;
  LAYER M1 ;
        RECT 0.719 3.864 0.721 6.3 ;
  LAYER M1 ;
        RECT 0.799 3.864 0.801 6.3 ;
  LAYER M1 ;
        RECT 0.879 3.864 0.881 6.3 ;
  LAYER M1 ;
        RECT 0.959 3.864 0.961 6.3 ;
  LAYER M1 ;
        RECT 1.039 3.864 1.041 6.3 ;
  LAYER M1 ;
        RECT 1.119 3.864 1.121 6.3 ;
  LAYER M1 ;
        RECT 1.199 3.864 1.201 6.3 ;
  LAYER M1 ;
        RECT 1.279 3.864 1.281 6.3 ;
  LAYER M1 ;
        RECT 1.359 3.864 1.361 6.3 ;
  LAYER M1 ;
        RECT 1.439 3.864 1.441 6.3 ;
  LAYER M1 ;
        RECT 1.519 3.864 1.521 6.3 ;
  LAYER M1 ;
        RECT 1.599 3.864 1.601 6.3 ;
  LAYER M1 ;
        RECT 1.679 3.864 1.681 6.3 ;
  LAYER M1 ;
        RECT 1.759 3.864 1.761 6.3 ;
  LAYER M1 ;
        RECT 1.839 3.864 1.841 6.3 ;
  LAYER M1 ;
        RECT 1.919 3.864 1.921 6.3 ;
  LAYER M1 ;
        RECT 1.999 3.864 2.001 6.3 ;
  LAYER M1 ;
        RECT 2.079 3.864 2.081 6.3 ;
  LAYER M1 ;
        RECT 2.159 3.864 2.161 6.3 ;
  LAYER M1 ;
        RECT 2.239 3.864 2.241 6.3 ;
  LAYER M1 ;
        RECT 2.319 3.864 2.321 6.3 ;
  LAYER M1 ;
        RECT 2.399 3.864 2.401 6.3 ;
  LAYER M2 ;
        RECT 0.08 3.863 2.48 3.865 ;
  LAYER M2 ;
        RECT 0.08 3.947 2.48 3.949 ;
  LAYER M2 ;
        RECT 0.08 4.031 2.48 4.033 ;
  LAYER M2 ;
        RECT 0.08 4.115 2.48 4.117 ;
  LAYER M2 ;
        RECT 0.08 4.199 2.48 4.201 ;
  LAYER M2 ;
        RECT 0.08 4.283 2.48 4.285 ;
  LAYER M2 ;
        RECT 0.08 4.367 2.48 4.369 ;
  LAYER M2 ;
        RECT 0.08 4.451 2.48 4.453 ;
  LAYER M2 ;
        RECT 0.08 4.535 2.48 4.537 ;
  LAYER M2 ;
        RECT 0.08 4.619 2.48 4.621 ;
  LAYER M2 ;
        RECT 0.08 4.703 2.48 4.705 ;
  LAYER M2 ;
        RECT 0.08 4.787 2.48 4.789 ;
  LAYER M2 ;
        RECT 0.08 4.8705 2.48 4.8725 ;
  LAYER M2 ;
        RECT 0.08 4.955 2.48 4.957 ;
  LAYER M2 ;
        RECT 0.08 5.039 2.48 5.041 ;
  LAYER M2 ;
        RECT 0.08 5.123 2.48 5.125 ;
  LAYER M2 ;
        RECT 0.08 5.207 2.48 5.209 ;
  LAYER M2 ;
        RECT 0.08 5.291 2.48 5.293 ;
  LAYER M2 ;
        RECT 0.08 5.375 2.48 5.377 ;
  LAYER M2 ;
        RECT 0.08 5.459 2.48 5.461 ;
  LAYER M2 ;
        RECT 0.08 5.543 2.48 5.545 ;
  LAYER M2 ;
        RECT 0.08 5.627 2.48 5.629 ;
  LAYER M2 ;
        RECT 0.08 5.711 2.48 5.713 ;
  LAYER M2 ;
        RECT 0.08 5.795 2.48 5.797 ;
  LAYER M2 ;
        RECT 0.08 5.879 2.48 5.881 ;
  LAYER M2 ;
        RECT 0.08 5.963 2.48 5.965 ;
  LAYER M2 ;
        RECT 0.08 6.047 2.48 6.049 ;
  LAYER M2 ;
        RECT 0.08 6.131 2.48 6.133 ;
  LAYER M2 ;
        RECT 0.08 6.215 2.48 6.217 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 9.276 ;
  LAYER M1 ;
        RECT 0.128 6.768 0.16 9.276 ;
  LAYER M1 ;
        RECT 0.192 6.768 0.224 9.276 ;
  LAYER M1 ;
        RECT 0.256 6.768 0.288 9.276 ;
  LAYER M1 ;
        RECT 0.32 6.768 0.352 9.276 ;
  LAYER M1 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M1 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M1 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M1 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M1 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M1 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M1 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M1 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M1 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M1 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M1 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M1 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M1 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M1 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M1 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M1 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M1 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M1 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M1 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M1 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M1 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M1 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M1 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M1 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M1 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M1 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M1 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M1 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M1 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M1 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M1 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M1 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M2 ;
        RECT 0.044 6.852 2.516 6.884 ;
  LAYER M2 ;
        RECT 0.044 6.916 2.516 6.948 ;
  LAYER M2 ;
        RECT 0.044 6.98 2.516 7.012 ;
  LAYER M2 ;
        RECT 0.044 7.044 2.516 7.076 ;
  LAYER M2 ;
        RECT 0.044 7.108 2.516 7.14 ;
  LAYER M2 ;
        RECT 0.044 7.172 2.516 7.204 ;
  LAYER M2 ;
        RECT 0.044 7.236 2.516 7.268 ;
  LAYER M2 ;
        RECT 0.044 7.3 2.516 7.332 ;
  LAYER M2 ;
        RECT 0.044 7.364 2.516 7.396 ;
  LAYER M2 ;
        RECT 0.044 7.428 2.516 7.46 ;
  LAYER M2 ;
        RECT 0.044 7.492 2.516 7.524 ;
  LAYER M2 ;
        RECT 0.044 7.556 2.516 7.588 ;
  LAYER M2 ;
        RECT 0.044 7.62 2.516 7.652 ;
  LAYER M2 ;
        RECT 0.044 7.684 2.516 7.716 ;
  LAYER M2 ;
        RECT 0.044 7.748 2.516 7.78 ;
  LAYER M2 ;
        RECT 0.044 7.812 2.516 7.844 ;
  LAYER M2 ;
        RECT 0.044 7.876 2.516 7.908 ;
  LAYER M2 ;
        RECT 0.044 7.94 2.516 7.972 ;
  LAYER M2 ;
        RECT 0.044 8.004 2.516 8.036 ;
  LAYER M2 ;
        RECT 0.044 8.068 2.516 8.1 ;
  LAYER M2 ;
        RECT 0.044 8.132 2.516 8.164 ;
  LAYER M2 ;
        RECT 0.044 8.196 2.516 8.228 ;
  LAYER M2 ;
        RECT 0.044 8.26 2.516 8.292 ;
  LAYER M2 ;
        RECT 0.044 8.324 2.516 8.356 ;
  LAYER M2 ;
        RECT 0.044 8.388 2.516 8.42 ;
  LAYER M2 ;
        RECT 0.044 8.452 2.516 8.484 ;
  LAYER M2 ;
        RECT 0.044 8.516 2.516 8.548 ;
  LAYER M2 ;
        RECT 0.044 8.58 2.516 8.612 ;
  LAYER M2 ;
        RECT 0.044 8.644 2.516 8.676 ;
  LAYER M2 ;
        RECT 0.044 8.708 2.516 8.74 ;
  LAYER M2 ;
        RECT 0.044 8.772 2.516 8.804 ;
  LAYER M2 ;
        RECT 0.044 8.836 2.516 8.868 ;
  LAYER M2 ;
        RECT 0.044 8.9 2.516 8.932 ;
  LAYER M2 ;
        RECT 0.044 8.964 2.516 8.996 ;
  LAYER M2 ;
        RECT 0.044 9.028 2.516 9.06 ;
  LAYER M2 ;
        RECT 0.044 9.092 2.516 9.124 ;
  LAYER M3 ;
        RECT 0.064 6.768 0.096 9.276 ;
  LAYER M3 ;
        RECT 0.128 6.768 0.16 9.276 ;
  LAYER M3 ;
        RECT 0.192 6.768 0.224 9.276 ;
  LAYER M3 ;
        RECT 0.256 6.768 0.288 9.276 ;
  LAYER M3 ;
        RECT 0.32 6.768 0.352 9.276 ;
  LAYER M3 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M3 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M3 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M3 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M3 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M3 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M3 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M3 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M3 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M3 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M3 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M3 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M3 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M3 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M3 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M3 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M3 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M3 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M3 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M3 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M3 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M3 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M3 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M3 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M3 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M3 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M3 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M3 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M3 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M3 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M3 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M3 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M3 ;
        RECT 2.464 6.768 2.496 9.276 ;
  LAYER M1 ;
        RECT 0.079 6.804 0.081 9.24 ;
  LAYER M1 ;
        RECT 0.159 6.804 0.161 9.24 ;
  LAYER M1 ;
        RECT 0.239 6.804 0.241 9.24 ;
  LAYER M1 ;
        RECT 0.319 6.804 0.321 9.24 ;
  LAYER M1 ;
        RECT 0.399 6.804 0.401 9.24 ;
  LAYER M1 ;
        RECT 0.479 6.804 0.481 9.24 ;
  LAYER M1 ;
        RECT 0.559 6.804 0.561 9.24 ;
  LAYER M1 ;
        RECT 0.639 6.804 0.641 9.24 ;
  LAYER M1 ;
        RECT 0.719 6.804 0.721 9.24 ;
  LAYER M1 ;
        RECT 0.799 6.804 0.801 9.24 ;
  LAYER M1 ;
        RECT 0.879 6.804 0.881 9.24 ;
  LAYER M1 ;
        RECT 0.959 6.804 0.961 9.24 ;
  LAYER M1 ;
        RECT 1.039 6.804 1.041 9.24 ;
  LAYER M1 ;
        RECT 1.119 6.804 1.121 9.24 ;
  LAYER M1 ;
        RECT 1.199 6.804 1.201 9.24 ;
  LAYER M1 ;
        RECT 1.279 6.804 1.281 9.24 ;
  LAYER M1 ;
        RECT 1.359 6.804 1.361 9.24 ;
  LAYER M1 ;
        RECT 1.439 6.804 1.441 9.24 ;
  LAYER M1 ;
        RECT 1.519 6.804 1.521 9.24 ;
  LAYER M1 ;
        RECT 1.599 6.804 1.601 9.24 ;
  LAYER M1 ;
        RECT 1.679 6.804 1.681 9.24 ;
  LAYER M1 ;
        RECT 1.759 6.804 1.761 9.24 ;
  LAYER M1 ;
        RECT 1.839 6.804 1.841 9.24 ;
  LAYER M1 ;
        RECT 1.919 6.804 1.921 9.24 ;
  LAYER M1 ;
        RECT 1.999 6.804 2.001 9.24 ;
  LAYER M1 ;
        RECT 2.079 6.804 2.081 9.24 ;
  LAYER M1 ;
        RECT 2.159 6.804 2.161 9.24 ;
  LAYER M1 ;
        RECT 2.239 6.804 2.241 9.24 ;
  LAYER M1 ;
        RECT 2.319 6.804 2.321 9.24 ;
  LAYER M1 ;
        RECT 2.399 6.804 2.401 9.24 ;
  LAYER M2 ;
        RECT 0.08 6.803 2.48 6.805 ;
  LAYER M2 ;
        RECT 0.08 6.887 2.48 6.889 ;
  LAYER M2 ;
        RECT 0.08 6.971 2.48 6.973 ;
  LAYER M2 ;
        RECT 0.08 7.055 2.48 7.057 ;
  LAYER M2 ;
        RECT 0.08 7.139 2.48 7.141 ;
  LAYER M2 ;
        RECT 0.08 7.223 2.48 7.225 ;
  LAYER M2 ;
        RECT 0.08 7.307 2.48 7.309 ;
  LAYER M2 ;
        RECT 0.08 7.391 2.48 7.393 ;
  LAYER M2 ;
        RECT 0.08 7.475 2.48 7.477 ;
  LAYER M2 ;
        RECT 0.08 7.559 2.48 7.561 ;
  LAYER M2 ;
        RECT 0.08 7.643 2.48 7.645 ;
  LAYER M2 ;
        RECT 0.08 7.727 2.48 7.729 ;
  LAYER M2 ;
        RECT 0.08 7.8105 2.48 7.8125 ;
  LAYER M2 ;
        RECT 0.08 7.895 2.48 7.897 ;
  LAYER M2 ;
        RECT 0.08 7.979 2.48 7.981 ;
  LAYER M2 ;
        RECT 0.08 8.063 2.48 8.065 ;
  LAYER M2 ;
        RECT 0.08 8.147 2.48 8.149 ;
  LAYER M2 ;
        RECT 0.08 8.231 2.48 8.233 ;
  LAYER M2 ;
        RECT 0.08 8.315 2.48 8.317 ;
  LAYER M2 ;
        RECT 0.08 8.399 2.48 8.401 ;
  LAYER M2 ;
        RECT 0.08 8.483 2.48 8.485 ;
  LAYER M2 ;
        RECT 0.08 8.567 2.48 8.569 ;
  LAYER M2 ;
        RECT 0.08 8.651 2.48 8.653 ;
  LAYER M2 ;
        RECT 0.08 8.735 2.48 8.737 ;
  LAYER M2 ;
        RECT 0.08 8.819 2.48 8.821 ;
  LAYER M2 ;
        RECT 0.08 8.903 2.48 8.905 ;
  LAYER M2 ;
        RECT 0.08 8.987 2.48 8.989 ;
  LAYER M2 ;
        RECT 0.08 9.071 2.48 9.073 ;
  LAYER M2 ;
        RECT 0.08 9.155 2.48 9.157 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 12.216 ;
  LAYER M1 ;
        RECT 0.128 9.708 0.16 12.216 ;
  LAYER M1 ;
        RECT 0.192 9.708 0.224 12.216 ;
  LAYER M1 ;
        RECT 0.256 9.708 0.288 12.216 ;
  LAYER M1 ;
        RECT 0.32 9.708 0.352 12.216 ;
  LAYER M1 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M1 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M1 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M1 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M1 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M1 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M1 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M1 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M1 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M1 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M1 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M1 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M1 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M1 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M1 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M1 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M1 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M1 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M1 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M1 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M1 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M1 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M1 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M1 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M1 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M1 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M1 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M1 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M1 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M1 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M1 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M1 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M2 ;
        RECT 0.044 9.792 2.516 9.824 ;
  LAYER M2 ;
        RECT 0.044 9.856 2.516 9.888 ;
  LAYER M2 ;
        RECT 0.044 9.92 2.516 9.952 ;
  LAYER M2 ;
        RECT 0.044 9.984 2.516 10.016 ;
  LAYER M2 ;
        RECT 0.044 10.048 2.516 10.08 ;
  LAYER M2 ;
        RECT 0.044 10.112 2.516 10.144 ;
  LAYER M2 ;
        RECT 0.044 10.176 2.516 10.208 ;
  LAYER M2 ;
        RECT 0.044 10.24 2.516 10.272 ;
  LAYER M2 ;
        RECT 0.044 10.304 2.516 10.336 ;
  LAYER M2 ;
        RECT 0.044 10.368 2.516 10.4 ;
  LAYER M2 ;
        RECT 0.044 10.432 2.516 10.464 ;
  LAYER M2 ;
        RECT 0.044 10.496 2.516 10.528 ;
  LAYER M2 ;
        RECT 0.044 10.56 2.516 10.592 ;
  LAYER M2 ;
        RECT 0.044 10.624 2.516 10.656 ;
  LAYER M2 ;
        RECT 0.044 10.688 2.516 10.72 ;
  LAYER M2 ;
        RECT 0.044 10.752 2.516 10.784 ;
  LAYER M2 ;
        RECT 0.044 10.816 2.516 10.848 ;
  LAYER M2 ;
        RECT 0.044 10.88 2.516 10.912 ;
  LAYER M2 ;
        RECT 0.044 10.944 2.516 10.976 ;
  LAYER M2 ;
        RECT 0.044 11.008 2.516 11.04 ;
  LAYER M2 ;
        RECT 0.044 11.072 2.516 11.104 ;
  LAYER M2 ;
        RECT 0.044 11.136 2.516 11.168 ;
  LAYER M2 ;
        RECT 0.044 11.2 2.516 11.232 ;
  LAYER M2 ;
        RECT 0.044 11.264 2.516 11.296 ;
  LAYER M2 ;
        RECT 0.044 11.328 2.516 11.36 ;
  LAYER M2 ;
        RECT 0.044 11.392 2.516 11.424 ;
  LAYER M2 ;
        RECT 0.044 11.456 2.516 11.488 ;
  LAYER M2 ;
        RECT 0.044 11.52 2.516 11.552 ;
  LAYER M2 ;
        RECT 0.044 11.584 2.516 11.616 ;
  LAYER M2 ;
        RECT 0.044 11.648 2.516 11.68 ;
  LAYER M2 ;
        RECT 0.044 11.712 2.516 11.744 ;
  LAYER M2 ;
        RECT 0.044 11.776 2.516 11.808 ;
  LAYER M2 ;
        RECT 0.044 11.84 2.516 11.872 ;
  LAYER M2 ;
        RECT 0.044 11.904 2.516 11.936 ;
  LAYER M2 ;
        RECT 0.044 11.968 2.516 12 ;
  LAYER M2 ;
        RECT 0.044 12.032 2.516 12.064 ;
  LAYER M3 ;
        RECT 0.064 9.708 0.096 12.216 ;
  LAYER M3 ;
        RECT 0.128 9.708 0.16 12.216 ;
  LAYER M3 ;
        RECT 0.192 9.708 0.224 12.216 ;
  LAYER M3 ;
        RECT 0.256 9.708 0.288 12.216 ;
  LAYER M3 ;
        RECT 0.32 9.708 0.352 12.216 ;
  LAYER M3 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M3 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M3 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M3 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M3 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M3 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M3 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M3 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M3 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M3 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M3 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M3 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M3 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M3 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M3 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M3 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M3 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M3 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M3 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M3 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M3 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M3 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M3 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M3 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M3 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M3 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M3 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M3 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M3 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M3 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M3 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M3 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M3 ;
        RECT 2.464 9.708 2.496 12.216 ;
  LAYER M1 ;
        RECT 0.079 9.744 0.081 12.18 ;
  LAYER M1 ;
        RECT 0.159 9.744 0.161 12.18 ;
  LAYER M1 ;
        RECT 0.239 9.744 0.241 12.18 ;
  LAYER M1 ;
        RECT 0.319 9.744 0.321 12.18 ;
  LAYER M1 ;
        RECT 0.399 9.744 0.401 12.18 ;
  LAYER M1 ;
        RECT 0.479 9.744 0.481 12.18 ;
  LAYER M1 ;
        RECT 0.559 9.744 0.561 12.18 ;
  LAYER M1 ;
        RECT 0.639 9.744 0.641 12.18 ;
  LAYER M1 ;
        RECT 0.719 9.744 0.721 12.18 ;
  LAYER M1 ;
        RECT 0.799 9.744 0.801 12.18 ;
  LAYER M1 ;
        RECT 0.879 9.744 0.881 12.18 ;
  LAYER M1 ;
        RECT 0.959 9.744 0.961 12.18 ;
  LAYER M1 ;
        RECT 1.039 9.744 1.041 12.18 ;
  LAYER M1 ;
        RECT 1.119 9.744 1.121 12.18 ;
  LAYER M1 ;
        RECT 1.199 9.744 1.201 12.18 ;
  LAYER M1 ;
        RECT 1.279 9.744 1.281 12.18 ;
  LAYER M1 ;
        RECT 1.359 9.744 1.361 12.18 ;
  LAYER M1 ;
        RECT 1.439 9.744 1.441 12.18 ;
  LAYER M1 ;
        RECT 1.519 9.744 1.521 12.18 ;
  LAYER M1 ;
        RECT 1.599 9.744 1.601 12.18 ;
  LAYER M1 ;
        RECT 1.679 9.744 1.681 12.18 ;
  LAYER M1 ;
        RECT 1.759 9.744 1.761 12.18 ;
  LAYER M1 ;
        RECT 1.839 9.744 1.841 12.18 ;
  LAYER M1 ;
        RECT 1.919 9.744 1.921 12.18 ;
  LAYER M1 ;
        RECT 1.999 9.744 2.001 12.18 ;
  LAYER M1 ;
        RECT 2.079 9.744 2.081 12.18 ;
  LAYER M1 ;
        RECT 2.159 9.744 2.161 12.18 ;
  LAYER M1 ;
        RECT 2.239 9.744 2.241 12.18 ;
  LAYER M1 ;
        RECT 2.319 9.744 2.321 12.18 ;
  LAYER M1 ;
        RECT 2.399 9.744 2.401 12.18 ;
  LAYER M2 ;
        RECT 0.08 9.743 2.48 9.745 ;
  LAYER M2 ;
        RECT 0.08 9.827 2.48 9.829 ;
  LAYER M2 ;
        RECT 0.08 9.911 2.48 9.913 ;
  LAYER M2 ;
        RECT 0.08 9.995 2.48 9.997 ;
  LAYER M2 ;
        RECT 0.08 10.079 2.48 10.081 ;
  LAYER M2 ;
        RECT 0.08 10.163 2.48 10.165 ;
  LAYER M2 ;
        RECT 0.08 10.247 2.48 10.249 ;
  LAYER M2 ;
        RECT 0.08 10.331 2.48 10.333 ;
  LAYER M2 ;
        RECT 0.08 10.415 2.48 10.417 ;
  LAYER M2 ;
        RECT 0.08 10.499 2.48 10.501 ;
  LAYER M2 ;
        RECT 0.08 10.583 2.48 10.585 ;
  LAYER M2 ;
        RECT 0.08 10.667 2.48 10.669 ;
  LAYER M2 ;
        RECT 0.08 10.7505 2.48 10.7525 ;
  LAYER M2 ;
        RECT 0.08 10.835 2.48 10.837 ;
  LAYER M2 ;
        RECT 0.08 10.919 2.48 10.921 ;
  LAYER M2 ;
        RECT 0.08 11.003 2.48 11.005 ;
  LAYER M2 ;
        RECT 0.08 11.087 2.48 11.089 ;
  LAYER M2 ;
        RECT 0.08 11.171 2.48 11.173 ;
  LAYER M2 ;
        RECT 0.08 11.255 2.48 11.257 ;
  LAYER M2 ;
        RECT 0.08 11.339 2.48 11.341 ;
  LAYER M2 ;
        RECT 0.08 11.423 2.48 11.425 ;
  LAYER M2 ;
        RECT 0.08 11.507 2.48 11.509 ;
  LAYER M2 ;
        RECT 0.08 11.591 2.48 11.593 ;
  LAYER M2 ;
        RECT 0.08 11.675 2.48 11.677 ;
  LAYER M2 ;
        RECT 0.08 11.759 2.48 11.761 ;
  LAYER M2 ;
        RECT 0.08 11.843 2.48 11.845 ;
  LAYER M2 ;
        RECT 0.08 11.927 2.48 11.929 ;
  LAYER M2 ;
        RECT 0.08 12.011 2.48 12.013 ;
  LAYER M2 ;
        RECT 0.08 12.095 2.48 12.097 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 15.156 ;
  LAYER M1 ;
        RECT 0.128 12.648 0.16 15.156 ;
  LAYER M1 ;
        RECT 0.192 12.648 0.224 15.156 ;
  LAYER M1 ;
        RECT 0.256 12.648 0.288 15.156 ;
  LAYER M1 ;
        RECT 0.32 12.648 0.352 15.156 ;
  LAYER M1 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M1 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M1 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M1 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M1 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M1 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M1 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M1 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M1 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M1 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M1 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M1 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M1 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M1 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M1 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M1 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M1 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M1 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M1 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M1 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M1 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M1 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M1 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M1 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M1 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M1 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M1 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M1 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M1 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M1 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M1 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M1 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M2 ;
        RECT 0.044 12.732 2.516 12.764 ;
  LAYER M2 ;
        RECT 0.044 12.796 2.516 12.828 ;
  LAYER M2 ;
        RECT 0.044 12.86 2.516 12.892 ;
  LAYER M2 ;
        RECT 0.044 12.924 2.516 12.956 ;
  LAYER M2 ;
        RECT 0.044 12.988 2.516 13.02 ;
  LAYER M2 ;
        RECT 0.044 13.052 2.516 13.084 ;
  LAYER M2 ;
        RECT 0.044 13.116 2.516 13.148 ;
  LAYER M2 ;
        RECT 0.044 13.18 2.516 13.212 ;
  LAYER M2 ;
        RECT 0.044 13.244 2.516 13.276 ;
  LAYER M2 ;
        RECT 0.044 13.308 2.516 13.34 ;
  LAYER M2 ;
        RECT 0.044 13.372 2.516 13.404 ;
  LAYER M2 ;
        RECT 0.044 13.436 2.516 13.468 ;
  LAYER M2 ;
        RECT 0.044 13.5 2.516 13.532 ;
  LAYER M2 ;
        RECT 0.044 13.564 2.516 13.596 ;
  LAYER M2 ;
        RECT 0.044 13.628 2.516 13.66 ;
  LAYER M2 ;
        RECT 0.044 13.692 2.516 13.724 ;
  LAYER M2 ;
        RECT 0.044 13.756 2.516 13.788 ;
  LAYER M2 ;
        RECT 0.044 13.82 2.516 13.852 ;
  LAYER M2 ;
        RECT 0.044 13.884 2.516 13.916 ;
  LAYER M2 ;
        RECT 0.044 13.948 2.516 13.98 ;
  LAYER M2 ;
        RECT 0.044 14.012 2.516 14.044 ;
  LAYER M2 ;
        RECT 0.044 14.076 2.516 14.108 ;
  LAYER M2 ;
        RECT 0.044 14.14 2.516 14.172 ;
  LAYER M2 ;
        RECT 0.044 14.204 2.516 14.236 ;
  LAYER M2 ;
        RECT 0.044 14.268 2.516 14.3 ;
  LAYER M2 ;
        RECT 0.044 14.332 2.516 14.364 ;
  LAYER M2 ;
        RECT 0.044 14.396 2.516 14.428 ;
  LAYER M2 ;
        RECT 0.044 14.46 2.516 14.492 ;
  LAYER M2 ;
        RECT 0.044 14.524 2.516 14.556 ;
  LAYER M2 ;
        RECT 0.044 14.588 2.516 14.62 ;
  LAYER M2 ;
        RECT 0.044 14.652 2.516 14.684 ;
  LAYER M2 ;
        RECT 0.044 14.716 2.516 14.748 ;
  LAYER M2 ;
        RECT 0.044 14.78 2.516 14.812 ;
  LAYER M2 ;
        RECT 0.044 14.844 2.516 14.876 ;
  LAYER M2 ;
        RECT 0.044 14.908 2.516 14.94 ;
  LAYER M2 ;
        RECT 0.044 14.972 2.516 15.004 ;
  LAYER M3 ;
        RECT 0.064 12.648 0.096 15.156 ;
  LAYER M3 ;
        RECT 0.128 12.648 0.16 15.156 ;
  LAYER M3 ;
        RECT 0.192 12.648 0.224 15.156 ;
  LAYER M3 ;
        RECT 0.256 12.648 0.288 15.156 ;
  LAYER M3 ;
        RECT 0.32 12.648 0.352 15.156 ;
  LAYER M3 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M3 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M3 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M3 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M3 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M3 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M3 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M3 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M3 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M3 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M3 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M3 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M3 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M3 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M3 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M3 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M3 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M3 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M3 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M3 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M3 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M3 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M3 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M3 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M3 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M3 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M3 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M3 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M3 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M3 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M3 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M3 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M3 ;
        RECT 2.464 12.648 2.496 15.156 ;
  LAYER M1 ;
        RECT 0.079 12.684 0.081 15.12 ;
  LAYER M1 ;
        RECT 0.159 12.684 0.161 15.12 ;
  LAYER M1 ;
        RECT 0.239 12.684 0.241 15.12 ;
  LAYER M1 ;
        RECT 0.319 12.684 0.321 15.12 ;
  LAYER M1 ;
        RECT 0.399 12.684 0.401 15.12 ;
  LAYER M1 ;
        RECT 0.479 12.684 0.481 15.12 ;
  LAYER M1 ;
        RECT 0.559 12.684 0.561 15.12 ;
  LAYER M1 ;
        RECT 0.639 12.684 0.641 15.12 ;
  LAYER M1 ;
        RECT 0.719 12.684 0.721 15.12 ;
  LAYER M1 ;
        RECT 0.799 12.684 0.801 15.12 ;
  LAYER M1 ;
        RECT 0.879 12.684 0.881 15.12 ;
  LAYER M1 ;
        RECT 0.959 12.684 0.961 15.12 ;
  LAYER M1 ;
        RECT 1.039 12.684 1.041 15.12 ;
  LAYER M1 ;
        RECT 1.119 12.684 1.121 15.12 ;
  LAYER M1 ;
        RECT 1.199 12.684 1.201 15.12 ;
  LAYER M1 ;
        RECT 1.279 12.684 1.281 15.12 ;
  LAYER M1 ;
        RECT 1.359 12.684 1.361 15.12 ;
  LAYER M1 ;
        RECT 1.439 12.684 1.441 15.12 ;
  LAYER M1 ;
        RECT 1.519 12.684 1.521 15.12 ;
  LAYER M1 ;
        RECT 1.599 12.684 1.601 15.12 ;
  LAYER M1 ;
        RECT 1.679 12.684 1.681 15.12 ;
  LAYER M1 ;
        RECT 1.759 12.684 1.761 15.12 ;
  LAYER M1 ;
        RECT 1.839 12.684 1.841 15.12 ;
  LAYER M1 ;
        RECT 1.919 12.684 1.921 15.12 ;
  LAYER M1 ;
        RECT 1.999 12.684 2.001 15.12 ;
  LAYER M1 ;
        RECT 2.079 12.684 2.081 15.12 ;
  LAYER M1 ;
        RECT 2.159 12.684 2.161 15.12 ;
  LAYER M1 ;
        RECT 2.239 12.684 2.241 15.12 ;
  LAYER M1 ;
        RECT 2.319 12.684 2.321 15.12 ;
  LAYER M1 ;
        RECT 2.399 12.684 2.401 15.12 ;
  LAYER M2 ;
        RECT 0.08 12.683 2.48 12.685 ;
  LAYER M2 ;
        RECT 0.08 12.767 2.48 12.769 ;
  LAYER M2 ;
        RECT 0.08 12.851 2.48 12.853 ;
  LAYER M2 ;
        RECT 0.08 12.935 2.48 12.937 ;
  LAYER M2 ;
        RECT 0.08 13.019 2.48 13.021 ;
  LAYER M2 ;
        RECT 0.08 13.103 2.48 13.105 ;
  LAYER M2 ;
        RECT 0.08 13.187 2.48 13.189 ;
  LAYER M2 ;
        RECT 0.08 13.271 2.48 13.273 ;
  LAYER M2 ;
        RECT 0.08 13.355 2.48 13.357 ;
  LAYER M2 ;
        RECT 0.08 13.439 2.48 13.441 ;
  LAYER M2 ;
        RECT 0.08 13.523 2.48 13.525 ;
  LAYER M2 ;
        RECT 0.08 13.607 2.48 13.609 ;
  LAYER M2 ;
        RECT 0.08 13.6905 2.48 13.6925 ;
  LAYER M2 ;
        RECT 0.08 13.775 2.48 13.777 ;
  LAYER M2 ;
        RECT 0.08 13.859 2.48 13.861 ;
  LAYER M2 ;
        RECT 0.08 13.943 2.48 13.945 ;
  LAYER M2 ;
        RECT 0.08 14.027 2.48 14.029 ;
  LAYER M2 ;
        RECT 0.08 14.111 2.48 14.113 ;
  LAYER M2 ;
        RECT 0.08 14.195 2.48 14.197 ;
  LAYER M2 ;
        RECT 0.08 14.279 2.48 14.281 ;
  LAYER M2 ;
        RECT 0.08 14.363 2.48 14.365 ;
  LAYER M2 ;
        RECT 0.08 14.447 2.48 14.449 ;
  LAYER M2 ;
        RECT 0.08 14.531 2.48 14.533 ;
  LAYER M2 ;
        RECT 0.08 14.615 2.48 14.617 ;
  LAYER M2 ;
        RECT 0.08 14.699 2.48 14.701 ;
  LAYER M2 ;
        RECT 0.08 14.783 2.48 14.785 ;
  LAYER M2 ;
        RECT 0.08 14.867 2.48 14.869 ;
  LAYER M2 ;
        RECT 0.08 14.951 2.48 14.953 ;
  LAYER M2 ;
        RECT 0.08 15.035 2.48 15.037 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 18.096 ;
  LAYER M1 ;
        RECT 0.128 15.588 0.16 18.096 ;
  LAYER M1 ;
        RECT 0.192 15.588 0.224 18.096 ;
  LAYER M1 ;
        RECT 0.256 15.588 0.288 18.096 ;
  LAYER M1 ;
        RECT 0.32 15.588 0.352 18.096 ;
  LAYER M1 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M1 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M1 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M1 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M1 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M1 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M1 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M1 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M1 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M1 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M1 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M1 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M1 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M1 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M1 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M1 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M1 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M1 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M1 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M1 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M1 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M1 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M1 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M1 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M1 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M1 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M1 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M1 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M1 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M1 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M1 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M1 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M2 ;
        RECT 0.044 15.672 2.516 15.704 ;
  LAYER M2 ;
        RECT 0.044 15.736 2.516 15.768 ;
  LAYER M2 ;
        RECT 0.044 15.8 2.516 15.832 ;
  LAYER M2 ;
        RECT 0.044 15.864 2.516 15.896 ;
  LAYER M2 ;
        RECT 0.044 15.928 2.516 15.96 ;
  LAYER M2 ;
        RECT 0.044 15.992 2.516 16.024 ;
  LAYER M2 ;
        RECT 0.044 16.056 2.516 16.088 ;
  LAYER M2 ;
        RECT 0.044 16.12 2.516 16.152 ;
  LAYER M2 ;
        RECT 0.044 16.184 2.516 16.216 ;
  LAYER M2 ;
        RECT 0.044 16.248 2.516 16.28 ;
  LAYER M2 ;
        RECT 0.044 16.312 2.516 16.344 ;
  LAYER M2 ;
        RECT 0.044 16.376 2.516 16.408 ;
  LAYER M2 ;
        RECT 0.044 16.44 2.516 16.472 ;
  LAYER M2 ;
        RECT 0.044 16.504 2.516 16.536 ;
  LAYER M2 ;
        RECT 0.044 16.568 2.516 16.6 ;
  LAYER M2 ;
        RECT 0.044 16.632 2.516 16.664 ;
  LAYER M2 ;
        RECT 0.044 16.696 2.516 16.728 ;
  LAYER M2 ;
        RECT 0.044 16.76 2.516 16.792 ;
  LAYER M2 ;
        RECT 0.044 16.824 2.516 16.856 ;
  LAYER M2 ;
        RECT 0.044 16.888 2.516 16.92 ;
  LAYER M2 ;
        RECT 0.044 16.952 2.516 16.984 ;
  LAYER M2 ;
        RECT 0.044 17.016 2.516 17.048 ;
  LAYER M2 ;
        RECT 0.044 17.08 2.516 17.112 ;
  LAYER M2 ;
        RECT 0.044 17.144 2.516 17.176 ;
  LAYER M2 ;
        RECT 0.044 17.208 2.516 17.24 ;
  LAYER M2 ;
        RECT 0.044 17.272 2.516 17.304 ;
  LAYER M2 ;
        RECT 0.044 17.336 2.516 17.368 ;
  LAYER M2 ;
        RECT 0.044 17.4 2.516 17.432 ;
  LAYER M2 ;
        RECT 0.044 17.464 2.516 17.496 ;
  LAYER M2 ;
        RECT 0.044 17.528 2.516 17.56 ;
  LAYER M2 ;
        RECT 0.044 17.592 2.516 17.624 ;
  LAYER M2 ;
        RECT 0.044 17.656 2.516 17.688 ;
  LAYER M2 ;
        RECT 0.044 17.72 2.516 17.752 ;
  LAYER M2 ;
        RECT 0.044 17.784 2.516 17.816 ;
  LAYER M2 ;
        RECT 0.044 17.848 2.516 17.88 ;
  LAYER M2 ;
        RECT 0.044 17.912 2.516 17.944 ;
  LAYER M3 ;
        RECT 0.064 15.588 0.096 18.096 ;
  LAYER M3 ;
        RECT 0.128 15.588 0.16 18.096 ;
  LAYER M3 ;
        RECT 0.192 15.588 0.224 18.096 ;
  LAYER M3 ;
        RECT 0.256 15.588 0.288 18.096 ;
  LAYER M3 ;
        RECT 0.32 15.588 0.352 18.096 ;
  LAYER M3 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M3 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M3 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M3 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M3 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M3 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M3 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M3 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M3 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M3 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M3 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M3 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M3 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M3 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M3 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M3 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M3 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M3 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M3 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M3 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M3 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M3 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M3 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M3 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M3 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M3 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M3 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M3 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M3 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M3 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M3 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M3 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M3 ;
        RECT 2.464 15.588 2.496 18.096 ;
  LAYER M1 ;
        RECT 0.079 15.624 0.081 18.06 ;
  LAYER M1 ;
        RECT 0.159 15.624 0.161 18.06 ;
  LAYER M1 ;
        RECT 0.239 15.624 0.241 18.06 ;
  LAYER M1 ;
        RECT 0.319 15.624 0.321 18.06 ;
  LAYER M1 ;
        RECT 0.399 15.624 0.401 18.06 ;
  LAYER M1 ;
        RECT 0.479 15.624 0.481 18.06 ;
  LAYER M1 ;
        RECT 0.559 15.624 0.561 18.06 ;
  LAYER M1 ;
        RECT 0.639 15.624 0.641 18.06 ;
  LAYER M1 ;
        RECT 0.719 15.624 0.721 18.06 ;
  LAYER M1 ;
        RECT 0.799 15.624 0.801 18.06 ;
  LAYER M1 ;
        RECT 0.879 15.624 0.881 18.06 ;
  LAYER M1 ;
        RECT 0.959 15.624 0.961 18.06 ;
  LAYER M1 ;
        RECT 1.039 15.624 1.041 18.06 ;
  LAYER M1 ;
        RECT 1.119 15.624 1.121 18.06 ;
  LAYER M1 ;
        RECT 1.199 15.624 1.201 18.06 ;
  LAYER M1 ;
        RECT 1.279 15.624 1.281 18.06 ;
  LAYER M1 ;
        RECT 1.359 15.624 1.361 18.06 ;
  LAYER M1 ;
        RECT 1.439 15.624 1.441 18.06 ;
  LAYER M1 ;
        RECT 1.519 15.624 1.521 18.06 ;
  LAYER M1 ;
        RECT 1.599 15.624 1.601 18.06 ;
  LAYER M1 ;
        RECT 1.679 15.624 1.681 18.06 ;
  LAYER M1 ;
        RECT 1.759 15.624 1.761 18.06 ;
  LAYER M1 ;
        RECT 1.839 15.624 1.841 18.06 ;
  LAYER M1 ;
        RECT 1.919 15.624 1.921 18.06 ;
  LAYER M1 ;
        RECT 1.999 15.624 2.001 18.06 ;
  LAYER M1 ;
        RECT 2.079 15.624 2.081 18.06 ;
  LAYER M1 ;
        RECT 2.159 15.624 2.161 18.06 ;
  LAYER M1 ;
        RECT 2.239 15.624 2.241 18.06 ;
  LAYER M1 ;
        RECT 2.319 15.624 2.321 18.06 ;
  LAYER M1 ;
        RECT 2.399 15.624 2.401 18.06 ;
  LAYER M2 ;
        RECT 0.08 15.623 2.48 15.625 ;
  LAYER M2 ;
        RECT 0.08 15.707 2.48 15.709 ;
  LAYER M2 ;
        RECT 0.08 15.791 2.48 15.793 ;
  LAYER M2 ;
        RECT 0.08 15.875 2.48 15.877 ;
  LAYER M2 ;
        RECT 0.08 15.959 2.48 15.961 ;
  LAYER M2 ;
        RECT 0.08 16.043 2.48 16.045 ;
  LAYER M2 ;
        RECT 0.08 16.127 2.48 16.129 ;
  LAYER M2 ;
        RECT 0.08 16.211 2.48 16.213 ;
  LAYER M2 ;
        RECT 0.08 16.295 2.48 16.297 ;
  LAYER M2 ;
        RECT 0.08 16.379 2.48 16.381 ;
  LAYER M2 ;
        RECT 0.08 16.463 2.48 16.465 ;
  LAYER M2 ;
        RECT 0.08 16.547 2.48 16.549 ;
  LAYER M2 ;
        RECT 0.08 16.6305 2.48 16.6325 ;
  LAYER M2 ;
        RECT 0.08 16.715 2.48 16.717 ;
  LAYER M2 ;
        RECT 0.08 16.799 2.48 16.801 ;
  LAYER M2 ;
        RECT 0.08 16.883 2.48 16.885 ;
  LAYER M2 ;
        RECT 0.08 16.967 2.48 16.969 ;
  LAYER M2 ;
        RECT 0.08 17.051 2.48 17.053 ;
  LAYER M2 ;
        RECT 0.08 17.135 2.48 17.137 ;
  LAYER M2 ;
        RECT 0.08 17.219 2.48 17.221 ;
  LAYER M2 ;
        RECT 0.08 17.303 2.48 17.305 ;
  LAYER M2 ;
        RECT 0.08 17.387 2.48 17.389 ;
  LAYER M2 ;
        RECT 0.08 17.471 2.48 17.473 ;
  LAYER M2 ;
        RECT 0.08 17.555 2.48 17.557 ;
  LAYER M2 ;
        RECT 0.08 17.639 2.48 17.641 ;
  LAYER M2 ;
        RECT 0.08 17.723 2.48 17.725 ;
  LAYER M2 ;
        RECT 0.08 17.807 2.48 17.809 ;
  LAYER M2 ;
        RECT 0.08 17.891 2.48 17.893 ;
  LAYER M2 ;
        RECT 0.08 17.975 2.48 17.977 ;
  LAYER M1 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M1 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M1 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M1 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M1 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M1 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M1 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M1 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M1 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M1 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M1 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M1 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M1 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M1 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M1 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M1 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M1 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M1 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M1 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M1 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M1 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M1 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M1 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M1 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M1 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M1 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M1 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M1 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M1 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M1 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M1 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M1 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M1 ;
        RECT 5.632 0.888 5.664 3.396 ;
  LAYER M1 ;
        RECT 5.696 0.888 5.728 3.396 ;
  LAYER M1 ;
        RECT 5.76 0.888 5.792 3.396 ;
  LAYER M1 ;
        RECT 5.824 0.888 5.856 3.396 ;
  LAYER M1 ;
        RECT 5.888 0.888 5.92 3.396 ;
  LAYER M2 ;
        RECT 3.564 0.972 6.036 1.004 ;
  LAYER M2 ;
        RECT 3.564 1.036 6.036 1.068 ;
  LAYER M2 ;
        RECT 3.564 1.1 6.036 1.132 ;
  LAYER M2 ;
        RECT 3.564 1.164 6.036 1.196 ;
  LAYER M2 ;
        RECT 3.564 1.228 6.036 1.26 ;
  LAYER M2 ;
        RECT 3.564 1.292 6.036 1.324 ;
  LAYER M2 ;
        RECT 3.564 1.356 6.036 1.388 ;
  LAYER M2 ;
        RECT 3.564 1.42 6.036 1.452 ;
  LAYER M2 ;
        RECT 3.564 1.484 6.036 1.516 ;
  LAYER M2 ;
        RECT 3.564 1.548 6.036 1.58 ;
  LAYER M2 ;
        RECT 3.564 1.612 6.036 1.644 ;
  LAYER M2 ;
        RECT 3.564 1.676 6.036 1.708 ;
  LAYER M2 ;
        RECT 3.564 1.74 6.036 1.772 ;
  LAYER M2 ;
        RECT 3.564 1.804 6.036 1.836 ;
  LAYER M2 ;
        RECT 3.564 1.868 6.036 1.9 ;
  LAYER M2 ;
        RECT 3.564 1.932 6.036 1.964 ;
  LAYER M2 ;
        RECT 3.564 1.996 6.036 2.028 ;
  LAYER M2 ;
        RECT 3.564 2.06 6.036 2.092 ;
  LAYER M2 ;
        RECT 3.564 2.124 6.036 2.156 ;
  LAYER M2 ;
        RECT 3.564 2.188 6.036 2.22 ;
  LAYER M2 ;
        RECT 3.564 2.252 6.036 2.284 ;
  LAYER M2 ;
        RECT 3.564 2.316 6.036 2.348 ;
  LAYER M2 ;
        RECT 3.564 2.38 6.036 2.412 ;
  LAYER M2 ;
        RECT 3.564 2.444 6.036 2.476 ;
  LAYER M2 ;
        RECT 3.564 2.508 6.036 2.54 ;
  LAYER M2 ;
        RECT 3.564 2.572 6.036 2.604 ;
  LAYER M2 ;
        RECT 3.564 2.636 6.036 2.668 ;
  LAYER M2 ;
        RECT 3.564 2.7 6.036 2.732 ;
  LAYER M2 ;
        RECT 3.564 2.764 6.036 2.796 ;
  LAYER M2 ;
        RECT 3.564 2.828 6.036 2.86 ;
  LAYER M2 ;
        RECT 3.564 2.892 6.036 2.924 ;
  LAYER M2 ;
        RECT 3.564 2.956 6.036 2.988 ;
  LAYER M2 ;
        RECT 3.564 3.02 6.036 3.052 ;
  LAYER M2 ;
        RECT 3.564 3.084 6.036 3.116 ;
  LAYER M2 ;
        RECT 3.564 3.148 6.036 3.18 ;
  LAYER M2 ;
        RECT 3.564 3.212 6.036 3.244 ;
  LAYER M3 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M3 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M3 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M3 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M3 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M3 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M3 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M3 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M3 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M3 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M3 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M3 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M3 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M3 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M3 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M3 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M3 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M3 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M3 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M3 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M3 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M3 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M3 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M3 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M3 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M3 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M3 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M3 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M3 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M3 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M3 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M3 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M3 ;
        RECT 5.632 0.888 5.664 3.396 ;
  LAYER M3 ;
        RECT 5.696 0.888 5.728 3.396 ;
  LAYER M3 ;
        RECT 5.76 0.888 5.792 3.396 ;
  LAYER M3 ;
        RECT 5.824 0.888 5.856 3.396 ;
  LAYER M3 ;
        RECT 5.888 0.888 5.92 3.396 ;
  LAYER M3 ;
        RECT 5.984 0.888 6.016 3.396 ;
  LAYER M1 ;
        RECT 3.599 0.924 3.601 3.36 ;
  LAYER M1 ;
        RECT 3.679 0.924 3.681 3.36 ;
  LAYER M1 ;
        RECT 3.759 0.924 3.761 3.36 ;
  LAYER M1 ;
        RECT 3.839 0.924 3.841 3.36 ;
  LAYER M1 ;
        RECT 3.919 0.924 3.921 3.36 ;
  LAYER M1 ;
        RECT 3.999 0.924 4.001 3.36 ;
  LAYER M1 ;
        RECT 4.079 0.924 4.081 3.36 ;
  LAYER M1 ;
        RECT 4.159 0.924 4.161 3.36 ;
  LAYER M1 ;
        RECT 4.239 0.924 4.241 3.36 ;
  LAYER M1 ;
        RECT 4.319 0.924 4.321 3.36 ;
  LAYER M1 ;
        RECT 4.399 0.924 4.401 3.36 ;
  LAYER M1 ;
        RECT 4.479 0.924 4.481 3.36 ;
  LAYER M1 ;
        RECT 4.559 0.924 4.561 3.36 ;
  LAYER M1 ;
        RECT 4.639 0.924 4.641 3.36 ;
  LAYER M1 ;
        RECT 4.719 0.924 4.721 3.36 ;
  LAYER M1 ;
        RECT 4.799 0.924 4.801 3.36 ;
  LAYER M1 ;
        RECT 4.879 0.924 4.881 3.36 ;
  LAYER M1 ;
        RECT 4.959 0.924 4.961 3.36 ;
  LAYER M1 ;
        RECT 5.039 0.924 5.041 3.36 ;
  LAYER M1 ;
        RECT 5.119 0.924 5.121 3.36 ;
  LAYER M1 ;
        RECT 5.199 0.924 5.201 3.36 ;
  LAYER M1 ;
        RECT 5.279 0.924 5.281 3.36 ;
  LAYER M1 ;
        RECT 5.359 0.924 5.361 3.36 ;
  LAYER M1 ;
        RECT 5.439 0.924 5.441 3.36 ;
  LAYER M1 ;
        RECT 5.519 0.924 5.521 3.36 ;
  LAYER M1 ;
        RECT 5.599 0.924 5.601 3.36 ;
  LAYER M1 ;
        RECT 5.679 0.924 5.681 3.36 ;
  LAYER M1 ;
        RECT 5.759 0.924 5.761 3.36 ;
  LAYER M1 ;
        RECT 5.839 0.924 5.841 3.36 ;
  LAYER M1 ;
        RECT 5.919 0.924 5.921 3.36 ;
  LAYER M2 ;
        RECT 3.6 0.923 6 0.925 ;
  LAYER M2 ;
        RECT 3.6 1.007 6 1.009 ;
  LAYER M2 ;
        RECT 3.6 1.091 6 1.093 ;
  LAYER M2 ;
        RECT 3.6 1.175 6 1.177 ;
  LAYER M2 ;
        RECT 3.6 1.259 6 1.261 ;
  LAYER M2 ;
        RECT 3.6 1.343 6 1.345 ;
  LAYER M2 ;
        RECT 3.6 1.427 6 1.429 ;
  LAYER M2 ;
        RECT 3.6 1.511 6 1.513 ;
  LAYER M2 ;
        RECT 3.6 1.595 6 1.597 ;
  LAYER M2 ;
        RECT 3.6 1.679 6 1.681 ;
  LAYER M2 ;
        RECT 3.6 1.763 6 1.765 ;
  LAYER M2 ;
        RECT 3.6 1.847 6 1.849 ;
  LAYER M2 ;
        RECT 3.6 1.9305 6 1.9325 ;
  LAYER M2 ;
        RECT 3.6 2.015 6 2.017 ;
  LAYER M2 ;
        RECT 3.6 2.099 6 2.101 ;
  LAYER M2 ;
        RECT 3.6 2.183 6 2.185 ;
  LAYER M2 ;
        RECT 3.6 2.267 6 2.269 ;
  LAYER M2 ;
        RECT 3.6 2.351 6 2.353 ;
  LAYER M2 ;
        RECT 3.6 2.435 6 2.437 ;
  LAYER M2 ;
        RECT 3.6 2.519 6 2.521 ;
  LAYER M2 ;
        RECT 3.6 2.603 6 2.605 ;
  LAYER M2 ;
        RECT 3.6 2.687 6 2.689 ;
  LAYER M2 ;
        RECT 3.6 2.771 6 2.773 ;
  LAYER M2 ;
        RECT 3.6 2.855 6 2.857 ;
  LAYER M2 ;
        RECT 3.6 2.939 6 2.941 ;
  LAYER M2 ;
        RECT 3.6 3.023 6 3.025 ;
  LAYER M2 ;
        RECT 3.6 3.107 6 3.109 ;
  LAYER M2 ;
        RECT 3.6 3.191 6 3.193 ;
  LAYER M2 ;
        RECT 3.6 3.275 6 3.277 ;
  LAYER M1 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M1 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M1 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M1 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M1 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M1 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M1 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M1 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M1 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M1 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M1 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M1 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M1 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M1 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M1 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M1 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M1 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M1 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M1 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M1 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M1 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M1 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M1 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M1 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M1 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M1 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M1 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M1 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M1 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M1 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M1 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M1 ;
        RECT 5.632 3.828 5.664 6.336 ;
  LAYER M1 ;
        RECT 5.696 3.828 5.728 6.336 ;
  LAYER M1 ;
        RECT 5.76 3.828 5.792 6.336 ;
  LAYER M1 ;
        RECT 5.824 3.828 5.856 6.336 ;
  LAYER M1 ;
        RECT 5.888 3.828 5.92 6.336 ;
  LAYER M2 ;
        RECT 3.564 3.912 6.036 3.944 ;
  LAYER M2 ;
        RECT 3.564 3.976 6.036 4.008 ;
  LAYER M2 ;
        RECT 3.564 4.04 6.036 4.072 ;
  LAYER M2 ;
        RECT 3.564 4.104 6.036 4.136 ;
  LAYER M2 ;
        RECT 3.564 4.168 6.036 4.2 ;
  LAYER M2 ;
        RECT 3.564 4.232 6.036 4.264 ;
  LAYER M2 ;
        RECT 3.564 4.296 6.036 4.328 ;
  LAYER M2 ;
        RECT 3.564 4.36 6.036 4.392 ;
  LAYER M2 ;
        RECT 3.564 4.424 6.036 4.456 ;
  LAYER M2 ;
        RECT 3.564 4.488 6.036 4.52 ;
  LAYER M2 ;
        RECT 3.564 4.552 6.036 4.584 ;
  LAYER M2 ;
        RECT 3.564 4.616 6.036 4.648 ;
  LAYER M2 ;
        RECT 3.564 4.68 6.036 4.712 ;
  LAYER M2 ;
        RECT 3.564 4.744 6.036 4.776 ;
  LAYER M2 ;
        RECT 3.564 4.808 6.036 4.84 ;
  LAYER M2 ;
        RECT 3.564 4.872 6.036 4.904 ;
  LAYER M2 ;
        RECT 3.564 4.936 6.036 4.968 ;
  LAYER M2 ;
        RECT 3.564 5 6.036 5.032 ;
  LAYER M2 ;
        RECT 3.564 5.064 6.036 5.096 ;
  LAYER M2 ;
        RECT 3.564 5.128 6.036 5.16 ;
  LAYER M2 ;
        RECT 3.564 5.192 6.036 5.224 ;
  LAYER M2 ;
        RECT 3.564 5.256 6.036 5.288 ;
  LAYER M2 ;
        RECT 3.564 5.32 6.036 5.352 ;
  LAYER M2 ;
        RECT 3.564 5.384 6.036 5.416 ;
  LAYER M2 ;
        RECT 3.564 5.448 6.036 5.48 ;
  LAYER M2 ;
        RECT 3.564 5.512 6.036 5.544 ;
  LAYER M2 ;
        RECT 3.564 5.576 6.036 5.608 ;
  LAYER M2 ;
        RECT 3.564 5.64 6.036 5.672 ;
  LAYER M2 ;
        RECT 3.564 5.704 6.036 5.736 ;
  LAYER M2 ;
        RECT 3.564 5.768 6.036 5.8 ;
  LAYER M2 ;
        RECT 3.564 5.832 6.036 5.864 ;
  LAYER M2 ;
        RECT 3.564 5.896 6.036 5.928 ;
  LAYER M2 ;
        RECT 3.564 5.96 6.036 5.992 ;
  LAYER M2 ;
        RECT 3.564 6.024 6.036 6.056 ;
  LAYER M2 ;
        RECT 3.564 6.088 6.036 6.12 ;
  LAYER M2 ;
        RECT 3.564 6.152 6.036 6.184 ;
  LAYER M3 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M3 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M3 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M3 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M3 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M3 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M3 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M3 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M3 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M3 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M3 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M3 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M3 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M3 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M3 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M3 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M3 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M3 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M3 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M3 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M3 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M3 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M3 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M3 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M3 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M3 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M3 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M3 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M3 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M3 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M3 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M3 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M3 ;
        RECT 5.632 3.828 5.664 6.336 ;
  LAYER M3 ;
        RECT 5.696 3.828 5.728 6.336 ;
  LAYER M3 ;
        RECT 5.76 3.828 5.792 6.336 ;
  LAYER M3 ;
        RECT 5.824 3.828 5.856 6.336 ;
  LAYER M3 ;
        RECT 5.888 3.828 5.92 6.336 ;
  LAYER M3 ;
        RECT 5.984 3.828 6.016 6.336 ;
  LAYER M1 ;
        RECT 3.599 3.864 3.601 6.3 ;
  LAYER M1 ;
        RECT 3.679 3.864 3.681 6.3 ;
  LAYER M1 ;
        RECT 3.759 3.864 3.761 6.3 ;
  LAYER M1 ;
        RECT 3.839 3.864 3.841 6.3 ;
  LAYER M1 ;
        RECT 3.919 3.864 3.921 6.3 ;
  LAYER M1 ;
        RECT 3.999 3.864 4.001 6.3 ;
  LAYER M1 ;
        RECT 4.079 3.864 4.081 6.3 ;
  LAYER M1 ;
        RECT 4.159 3.864 4.161 6.3 ;
  LAYER M1 ;
        RECT 4.239 3.864 4.241 6.3 ;
  LAYER M1 ;
        RECT 4.319 3.864 4.321 6.3 ;
  LAYER M1 ;
        RECT 4.399 3.864 4.401 6.3 ;
  LAYER M1 ;
        RECT 4.479 3.864 4.481 6.3 ;
  LAYER M1 ;
        RECT 4.559 3.864 4.561 6.3 ;
  LAYER M1 ;
        RECT 4.639 3.864 4.641 6.3 ;
  LAYER M1 ;
        RECT 4.719 3.864 4.721 6.3 ;
  LAYER M1 ;
        RECT 4.799 3.864 4.801 6.3 ;
  LAYER M1 ;
        RECT 4.879 3.864 4.881 6.3 ;
  LAYER M1 ;
        RECT 4.959 3.864 4.961 6.3 ;
  LAYER M1 ;
        RECT 5.039 3.864 5.041 6.3 ;
  LAYER M1 ;
        RECT 5.119 3.864 5.121 6.3 ;
  LAYER M1 ;
        RECT 5.199 3.864 5.201 6.3 ;
  LAYER M1 ;
        RECT 5.279 3.864 5.281 6.3 ;
  LAYER M1 ;
        RECT 5.359 3.864 5.361 6.3 ;
  LAYER M1 ;
        RECT 5.439 3.864 5.441 6.3 ;
  LAYER M1 ;
        RECT 5.519 3.864 5.521 6.3 ;
  LAYER M1 ;
        RECT 5.599 3.864 5.601 6.3 ;
  LAYER M1 ;
        RECT 5.679 3.864 5.681 6.3 ;
  LAYER M1 ;
        RECT 5.759 3.864 5.761 6.3 ;
  LAYER M1 ;
        RECT 5.839 3.864 5.841 6.3 ;
  LAYER M1 ;
        RECT 5.919 3.864 5.921 6.3 ;
  LAYER M2 ;
        RECT 3.6 3.863 6 3.865 ;
  LAYER M2 ;
        RECT 3.6 3.947 6 3.949 ;
  LAYER M2 ;
        RECT 3.6 4.031 6 4.033 ;
  LAYER M2 ;
        RECT 3.6 4.115 6 4.117 ;
  LAYER M2 ;
        RECT 3.6 4.199 6 4.201 ;
  LAYER M2 ;
        RECT 3.6 4.283 6 4.285 ;
  LAYER M2 ;
        RECT 3.6 4.367 6 4.369 ;
  LAYER M2 ;
        RECT 3.6 4.451 6 4.453 ;
  LAYER M2 ;
        RECT 3.6 4.535 6 4.537 ;
  LAYER M2 ;
        RECT 3.6 4.619 6 4.621 ;
  LAYER M2 ;
        RECT 3.6 4.703 6 4.705 ;
  LAYER M2 ;
        RECT 3.6 4.787 6 4.789 ;
  LAYER M2 ;
        RECT 3.6 4.8705 6 4.8725 ;
  LAYER M2 ;
        RECT 3.6 4.955 6 4.957 ;
  LAYER M2 ;
        RECT 3.6 5.039 6 5.041 ;
  LAYER M2 ;
        RECT 3.6 5.123 6 5.125 ;
  LAYER M2 ;
        RECT 3.6 5.207 6 5.209 ;
  LAYER M2 ;
        RECT 3.6 5.291 6 5.293 ;
  LAYER M2 ;
        RECT 3.6 5.375 6 5.377 ;
  LAYER M2 ;
        RECT 3.6 5.459 6 5.461 ;
  LAYER M2 ;
        RECT 3.6 5.543 6 5.545 ;
  LAYER M2 ;
        RECT 3.6 5.627 6 5.629 ;
  LAYER M2 ;
        RECT 3.6 5.711 6 5.713 ;
  LAYER M2 ;
        RECT 3.6 5.795 6 5.797 ;
  LAYER M2 ;
        RECT 3.6 5.879 6 5.881 ;
  LAYER M2 ;
        RECT 3.6 5.963 6 5.965 ;
  LAYER M2 ;
        RECT 3.6 6.047 6 6.049 ;
  LAYER M2 ;
        RECT 3.6 6.131 6 6.133 ;
  LAYER M2 ;
        RECT 3.6 6.215 6 6.217 ;
  LAYER M1 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M1 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M1 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M1 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M1 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M1 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M1 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M1 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M1 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M1 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M1 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M1 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M1 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M1 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M1 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M1 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M1 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M1 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M1 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M1 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M1 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M1 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M1 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M1 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M1 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M1 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M1 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M1 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M1 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M1 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M1 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M1 ;
        RECT 5.632 6.768 5.664 9.276 ;
  LAYER M1 ;
        RECT 5.696 6.768 5.728 9.276 ;
  LAYER M1 ;
        RECT 5.76 6.768 5.792 9.276 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 9.276 ;
  LAYER M1 ;
        RECT 5.888 6.768 5.92 9.276 ;
  LAYER M2 ;
        RECT 3.564 6.852 6.036 6.884 ;
  LAYER M2 ;
        RECT 3.564 6.916 6.036 6.948 ;
  LAYER M2 ;
        RECT 3.564 6.98 6.036 7.012 ;
  LAYER M2 ;
        RECT 3.564 7.044 6.036 7.076 ;
  LAYER M2 ;
        RECT 3.564 7.108 6.036 7.14 ;
  LAYER M2 ;
        RECT 3.564 7.172 6.036 7.204 ;
  LAYER M2 ;
        RECT 3.564 7.236 6.036 7.268 ;
  LAYER M2 ;
        RECT 3.564 7.3 6.036 7.332 ;
  LAYER M2 ;
        RECT 3.564 7.364 6.036 7.396 ;
  LAYER M2 ;
        RECT 3.564 7.428 6.036 7.46 ;
  LAYER M2 ;
        RECT 3.564 7.492 6.036 7.524 ;
  LAYER M2 ;
        RECT 3.564 7.556 6.036 7.588 ;
  LAYER M2 ;
        RECT 3.564 7.62 6.036 7.652 ;
  LAYER M2 ;
        RECT 3.564 7.684 6.036 7.716 ;
  LAYER M2 ;
        RECT 3.564 7.748 6.036 7.78 ;
  LAYER M2 ;
        RECT 3.564 7.812 6.036 7.844 ;
  LAYER M2 ;
        RECT 3.564 7.876 6.036 7.908 ;
  LAYER M2 ;
        RECT 3.564 7.94 6.036 7.972 ;
  LAYER M2 ;
        RECT 3.564 8.004 6.036 8.036 ;
  LAYER M2 ;
        RECT 3.564 8.068 6.036 8.1 ;
  LAYER M2 ;
        RECT 3.564 8.132 6.036 8.164 ;
  LAYER M2 ;
        RECT 3.564 8.196 6.036 8.228 ;
  LAYER M2 ;
        RECT 3.564 8.26 6.036 8.292 ;
  LAYER M2 ;
        RECT 3.564 8.324 6.036 8.356 ;
  LAYER M2 ;
        RECT 3.564 8.388 6.036 8.42 ;
  LAYER M2 ;
        RECT 3.564 8.452 6.036 8.484 ;
  LAYER M2 ;
        RECT 3.564 8.516 6.036 8.548 ;
  LAYER M2 ;
        RECT 3.564 8.58 6.036 8.612 ;
  LAYER M2 ;
        RECT 3.564 8.644 6.036 8.676 ;
  LAYER M2 ;
        RECT 3.564 8.708 6.036 8.74 ;
  LAYER M2 ;
        RECT 3.564 8.772 6.036 8.804 ;
  LAYER M2 ;
        RECT 3.564 8.836 6.036 8.868 ;
  LAYER M2 ;
        RECT 3.564 8.9 6.036 8.932 ;
  LAYER M2 ;
        RECT 3.564 8.964 6.036 8.996 ;
  LAYER M2 ;
        RECT 3.564 9.028 6.036 9.06 ;
  LAYER M2 ;
        RECT 3.564 9.092 6.036 9.124 ;
  LAYER M3 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M3 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M3 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M3 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M3 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M3 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M3 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M3 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M3 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M3 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M3 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M3 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M3 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M3 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M3 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M3 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M3 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M3 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M3 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M3 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M3 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M3 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M3 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M3 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M3 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M3 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M3 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M3 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M3 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M3 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M3 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M3 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M3 ;
        RECT 5.632 6.768 5.664 9.276 ;
  LAYER M3 ;
        RECT 5.696 6.768 5.728 9.276 ;
  LAYER M3 ;
        RECT 5.76 6.768 5.792 9.276 ;
  LAYER M3 ;
        RECT 5.824 6.768 5.856 9.276 ;
  LAYER M3 ;
        RECT 5.888 6.768 5.92 9.276 ;
  LAYER M3 ;
        RECT 5.984 6.768 6.016 9.276 ;
  LAYER M1 ;
        RECT 3.599 6.804 3.601 9.24 ;
  LAYER M1 ;
        RECT 3.679 6.804 3.681 9.24 ;
  LAYER M1 ;
        RECT 3.759 6.804 3.761 9.24 ;
  LAYER M1 ;
        RECT 3.839 6.804 3.841 9.24 ;
  LAYER M1 ;
        RECT 3.919 6.804 3.921 9.24 ;
  LAYER M1 ;
        RECT 3.999 6.804 4.001 9.24 ;
  LAYER M1 ;
        RECT 4.079 6.804 4.081 9.24 ;
  LAYER M1 ;
        RECT 4.159 6.804 4.161 9.24 ;
  LAYER M1 ;
        RECT 4.239 6.804 4.241 9.24 ;
  LAYER M1 ;
        RECT 4.319 6.804 4.321 9.24 ;
  LAYER M1 ;
        RECT 4.399 6.804 4.401 9.24 ;
  LAYER M1 ;
        RECT 4.479 6.804 4.481 9.24 ;
  LAYER M1 ;
        RECT 4.559 6.804 4.561 9.24 ;
  LAYER M1 ;
        RECT 4.639 6.804 4.641 9.24 ;
  LAYER M1 ;
        RECT 4.719 6.804 4.721 9.24 ;
  LAYER M1 ;
        RECT 4.799 6.804 4.801 9.24 ;
  LAYER M1 ;
        RECT 4.879 6.804 4.881 9.24 ;
  LAYER M1 ;
        RECT 4.959 6.804 4.961 9.24 ;
  LAYER M1 ;
        RECT 5.039 6.804 5.041 9.24 ;
  LAYER M1 ;
        RECT 5.119 6.804 5.121 9.24 ;
  LAYER M1 ;
        RECT 5.199 6.804 5.201 9.24 ;
  LAYER M1 ;
        RECT 5.279 6.804 5.281 9.24 ;
  LAYER M1 ;
        RECT 5.359 6.804 5.361 9.24 ;
  LAYER M1 ;
        RECT 5.439 6.804 5.441 9.24 ;
  LAYER M1 ;
        RECT 5.519 6.804 5.521 9.24 ;
  LAYER M1 ;
        RECT 5.599 6.804 5.601 9.24 ;
  LAYER M1 ;
        RECT 5.679 6.804 5.681 9.24 ;
  LAYER M1 ;
        RECT 5.759 6.804 5.761 9.24 ;
  LAYER M1 ;
        RECT 5.839 6.804 5.841 9.24 ;
  LAYER M1 ;
        RECT 5.919 6.804 5.921 9.24 ;
  LAYER M2 ;
        RECT 3.6 6.803 6 6.805 ;
  LAYER M2 ;
        RECT 3.6 6.887 6 6.889 ;
  LAYER M2 ;
        RECT 3.6 6.971 6 6.973 ;
  LAYER M2 ;
        RECT 3.6 7.055 6 7.057 ;
  LAYER M2 ;
        RECT 3.6 7.139 6 7.141 ;
  LAYER M2 ;
        RECT 3.6 7.223 6 7.225 ;
  LAYER M2 ;
        RECT 3.6 7.307 6 7.309 ;
  LAYER M2 ;
        RECT 3.6 7.391 6 7.393 ;
  LAYER M2 ;
        RECT 3.6 7.475 6 7.477 ;
  LAYER M2 ;
        RECT 3.6 7.559 6 7.561 ;
  LAYER M2 ;
        RECT 3.6 7.643 6 7.645 ;
  LAYER M2 ;
        RECT 3.6 7.727 6 7.729 ;
  LAYER M2 ;
        RECT 3.6 7.8105 6 7.8125 ;
  LAYER M2 ;
        RECT 3.6 7.895 6 7.897 ;
  LAYER M2 ;
        RECT 3.6 7.979 6 7.981 ;
  LAYER M2 ;
        RECT 3.6 8.063 6 8.065 ;
  LAYER M2 ;
        RECT 3.6 8.147 6 8.149 ;
  LAYER M2 ;
        RECT 3.6 8.231 6 8.233 ;
  LAYER M2 ;
        RECT 3.6 8.315 6 8.317 ;
  LAYER M2 ;
        RECT 3.6 8.399 6 8.401 ;
  LAYER M2 ;
        RECT 3.6 8.483 6 8.485 ;
  LAYER M2 ;
        RECT 3.6 8.567 6 8.569 ;
  LAYER M2 ;
        RECT 3.6 8.651 6 8.653 ;
  LAYER M2 ;
        RECT 3.6 8.735 6 8.737 ;
  LAYER M2 ;
        RECT 3.6 8.819 6 8.821 ;
  LAYER M2 ;
        RECT 3.6 8.903 6 8.905 ;
  LAYER M2 ;
        RECT 3.6 8.987 6 8.989 ;
  LAYER M2 ;
        RECT 3.6 9.071 6 9.073 ;
  LAYER M2 ;
        RECT 3.6 9.155 6 9.157 ;
  LAYER M1 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M1 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M1 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M1 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M1 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M1 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M1 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M1 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M1 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M1 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M1 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M1 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M1 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M1 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M1 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M1 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M1 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M1 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M1 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M1 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M1 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M1 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M1 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M1 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M1 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M1 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M1 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M1 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M1 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M1 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M1 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M1 ;
        RECT 5.632 9.708 5.664 12.216 ;
  LAYER M1 ;
        RECT 5.696 9.708 5.728 12.216 ;
  LAYER M1 ;
        RECT 5.76 9.708 5.792 12.216 ;
  LAYER M1 ;
        RECT 5.824 9.708 5.856 12.216 ;
  LAYER M1 ;
        RECT 5.888 9.708 5.92 12.216 ;
  LAYER M2 ;
        RECT 3.564 9.792 6.036 9.824 ;
  LAYER M2 ;
        RECT 3.564 9.856 6.036 9.888 ;
  LAYER M2 ;
        RECT 3.564 9.92 6.036 9.952 ;
  LAYER M2 ;
        RECT 3.564 9.984 6.036 10.016 ;
  LAYER M2 ;
        RECT 3.564 10.048 6.036 10.08 ;
  LAYER M2 ;
        RECT 3.564 10.112 6.036 10.144 ;
  LAYER M2 ;
        RECT 3.564 10.176 6.036 10.208 ;
  LAYER M2 ;
        RECT 3.564 10.24 6.036 10.272 ;
  LAYER M2 ;
        RECT 3.564 10.304 6.036 10.336 ;
  LAYER M2 ;
        RECT 3.564 10.368 6.036 10.4 ;
  LAYER M2 ;
        RECT 3.564 10.432 6.036 10.464 ;
  LAYER M2 ;
        RECT 3.564 10.496 6.036 10.528 ;
  LAYER M2 ;
        RECT 3.564 10.56 6.036 10.592 ;
  LAYER M2 ;
        RECT 3.564 10.624 6.036 10.656 ;
  LAYER M2 ;
        RECT 3.564 10.688 6.036 10.72 ;
  LAYER M2 ;
        RECT 3.564 10.752 6.036 10.784 ;
  LAYER M2 ;
        RECT 3.564 10.816 6.036 10.848 ;
  LAYER M2 ;
        RECT 3.564 10.88 6.036 10.912 ;
  LAYER M2 ;
        RECT 3.564 10.944 6.036 10.976 ;
  LAYER M2 ;
        RECT 3.564 11.008 6.036 11.04 ;
  LAYER M2 ;
        RECT 3.564 11.072 6.036 11.104 ;
  LAYER M2 ;
        RECT 3.564 11.136 6.036 11.168 ;
  LAYER M2 ;
        RECT 3.564 11.2 6.036 11.232 ;
  LAYER M2 ;
        RECT 3.564 11.264 6.036 11.296 ;
  LAYER M2 ;
        RECT 3.564 11.328 6.036 11.36 ;
  LAYER M2 ;
        RECT 3.564 11.392 6.036 11.424 ;
  LAYER M2 ;
        RECT 3.564 11.456 6.036 11.488 ;
  LAYER M2 ;
        RECT 3.564 11.52 6.036 11.552 ;
  LAYER M2 ;
        RECT 3.564 11.584 6.036 11.616 ;
  LAYER M2 ;
        RECT 3.564 11.648 6.036 11.68 ;
  LAYER M2 ;
        RECT 3.564 11.712 6.036 11.744 ;
  LAYER M2 ;
        RECT 3.564 11.776 6.036 11.808 ;
  LAYER M2 ;
        RECT 3.564 11.84 6.036 11.872 ;
  LAYER M2 ;
        RECT 3.564 11.904 6.036 11.936 ;
  LAYER M2 ;
        RECT 3.564 11.968 6.036 12 ;
  LAYER M2 ;
        RECT 3.564 12.032 6.036 12.064 ;
  LAYER M3 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M3 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M3 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M3 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M3 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M3 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M3 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M3 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M3 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M3 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M3 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M3 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M3 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M3 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M3 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M3 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M3 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M3 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M3 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M3 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M3 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M3 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M3 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M3 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M3 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M3 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M3 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M3 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M3 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M3 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M3 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M3 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M3 ;
        RECT 5.632 9.708 5.664 12.216 ;
  LAYER M3 ;
        RECT 5.696 9.708 5.728 12.216 ;
  LAYER M3 ;
        RECT 5.76 9.708 5.792 12.216 ;
  LAYER M3 ;
        RECT 5.824 9.708 5.856 12.216 ;
  LAYER M3 ;
        RECT 5.888 9.708 5.92 12.216 ;
  LAYER M3 ;
        RECT 5.984 9.708 6.016 12.216 ;
  LAYER M1 ;
        RECT 3.599 9.744 3.601 12.18 ;
  LAYER M1 ;
        RECT 3.679 9.744 3.681 12.18 ;
  LAYER M1 ;
        RECT 3.759 9.744 3.761 12.18 ;
  LAYER M1 ;
        RECT 3.839 9.744 3.841 12.18 ;
  LAYER M1 ;
        RECT 3.919 9.744 3.921 12.18 ;
  LAYER M1 ;
        RECT 3.999 9.744 4.001 12.18 ;
  LAYER M1 ;
        RECT 4.079 9.744 4.081 12.18 ;
  LAYER M1 ;
        RECT 4.159 9.744 4.161 12.18 ;
  LAYER M1 ;
        RECT 4.239 9.744 4.241 12.18 ;
  LAYER M1 ;
        RECT 4.319 9.744 4.321 12.18 ;
  LAYER M1 ;
        RECT 4.399 9.744 4.401 12.18 ;
  LAYER M1 ;
        RECT 4.479 9.744 4.481 12.18 ;
  LAYER M1 ;
        RECT 4.559 9.744 4.561 12.18 ;
  LAYER M1 ;
        RECT 4.639 9.744 4.641 12.18 ;
  LAYER M1 ;
        RECT 4.719 9.744 4.721 12.18 ;
  LAYER M1 ;
        RECT 4.799 9.744 4.801 12.18 ;
  LAYER M1 ;
        RECT 4.879 9.744 4.881 12.18 ;
  LAYER M1 ;
        RECT 4.959 9.744 4.961 12.18 ;
  LAYER M1 ;
        RECT 5.039 9.744 5.041 12.18 ;
  LAYER M1 ;
        RECT 5.119 9.744 5.121 12.18 ;
  LAYER M1 ;
        RECT 5.199 9.744 5.201 12.18 ;
  LAYER M1 ;
        RECT 5.279 9.744 5.281 12.18 ;
  LAYER M1 ;
        RECT 5.359 9.744 5.361 12.18 ;
  LAYER M1 ;
        RECT 5.439 9.744 5.441 12.18 ;
  LAYER M1 ;
        RECT 5.519 9.744 5.521 12.18 ;
  LAYER M1 ;
        RECT 5.599 9.744 5.601 12.18 ;
  LAYER M1 ;
        RECT 5.679 9.744 5.681 12.18 ;
  LAYER M1 ;
        RECT 5.759 9.744 5.761 12.18 ;
  LAYER M1 ;
        RECT 5.839 9.744 5.841 12.18 ;
  LAYER M1 ;
        RECT 5.919 9.744 5.921 12.18 ;
  LAYER M2 ;
        RECT 3.6 9.743 6 9.745 ;
  LAYER M2 ;
        RECT 3.6 9.827 6 9.829 ;
  LAYER M2 ;
        RECT 3.6 9.911 6 9.913 ;
  LAYER M2 ;
        RECT 3.6 9.995 6 9.997 ;
  LAYER M2 ;
        RECT 3.6 10.079 6 10.081 ;
  LAYER M2 ;
        RECT 3.6 10.163 6 10.165 ;
  LAYER M2 ;
        RECT 3.6 10.247 6 10.249 ;
  LAYER M2 ;
        RECT 3.6 10.331 6 10.333 ;
  LAYER M2 ;
        RECT 3.6 10.415 6 10.417 ;
  LAYER M2 ;
        RECT 3.6 10.499 6 10.501 ;
  LAYER M2 ;
        RECT 3.6 10.583 6 10.585 ;
  LAYER M2 ;
        RECT 3.6 10.667 6 10.669 ;
  LAYER M2 ;
        RECT 3.6 10.7505 6 10.7525 ;
  LAYER M2 ;
        RECT 3.6 10.835 6 10.837 ;
  LAYER M2 ;
        RECT 3.6 10.919 6 10.921 ;
  LAYER M2 ;
        RECT 3.6 11.003 6 11.005 ;
  LAYER M2 ;
        RECT 3.6 11.087 6 11.089 ;
  LAYER M2 ;
        RECT 3.6 11.171 6 11.173 ;
  LAYER M2 ;
        RECT 3.6 11.255 6 11.257 ;
  LAYER M2 ;
        RECT 3.6 11.339 6 11.341 ;
  LAYER M2 ;
        RECT 3.6 11.423 6 11.425 ;
  LAYER M2 ;
        RECT 3.6 11.507 6 11.509 ;
  LAYER M2 ;
        RECT 3.6 11.591 6 11.593 ;
  LAYER M2 ;
        RECT 3.6 11.675 6 11.677 ;
  LAYER M2 ;
        RECT 3.6 11.759 6 11.761 ;
  LAYER M2 ;
        RECT 3.6 11.843 6 11.845 ;
  LAYER M2 ;
        RECT 3.6 11.927 6 11.929 ;
  LAYER M2 ;
        RECT 3.6 12.011 6 12.013 ;
  LAYER M2 ;
        RECT 3.6 12.095 6 12.097 ;
  LAYER M1 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M1 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M1 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M1 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M1 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M1 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M1 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M1 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M1 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M1 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M1 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M1 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M1 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M1 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M1 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M1 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M1 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M1 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M1 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M1 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M1 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M1 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M1 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M1 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M1 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M1 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M1 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M1 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M1 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M1 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M1 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M1 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M1 ;
        RECT 5.632 12.648 5.664 15.156 ;
  LAYER M1 ;
        RECT 5.696 12.648 5.728 15.156 ;
  LAYER M1 ;
        RECT 5.76 12.648 5.792 15.156 ;
  LAYER M1 ;
        RECT 5.824 12.648 5.856 15.156 ;
  LAYER M1 ;
        RECT 5.888 12.648 5.92 15.156 ;
  LAYER M2 ;
        RECT 3.564 12.732 6.036 12.764 ;
  LAYER M2 ;
        RECT 3.564 12.796 6.036 12.828 ;
  LAYER M2 ;
        RECT 3.564 12.86 6.036 12.892 ;
  LAYER M2 ;
        RECT 3.564 12.924 6.036 12.956 ;
  LAYER M2 ;
        RECT 3.564 12.988 6.036 13.02 ;
  LAYER M2 ;
        RECT 3.564 13.052 6.036 13.084 ;
  LAYER M2 ;
        RECT 3.564 13.116 6.036 13.148 ;
  LAYER M2 ;
        RECT 3.564 13.18 6.036 13.212 ;
  LAYER M2 ;
        RECT 3.564 13.244 6.036 13.276 ;
  LAYER M2 ;
        RECT 3.564 13.308 6.036 13.34 ;
  LAYER M2 ;
        RECT 3.564 13.372 6.036 13.404 ;
  LAYER M2 ;
        RECT 3.564 13.436 6.036 13.468 ;
  LAYER M2 ;
        RECT 3.564 13.5 6.036 13.532 ;
  LAYER M2 ;
        RECT 3.564 13.564 6.036 13.596 ;
  LAYER M2 ;
        RECT 3.564 13.628 6.036 13.66 ;
  LAYER M2 ;
        RECT 3.564 13.692 6.036 13.724 ;
  LAYER M2 ;
        RECT 3.564 13.756 6.036 13.788 ;
  LAYER M2 ;
        RECT 3.564 13.82 6.036 13.852 ;
  LAYER M2 ;
        RECT 3.564 13.884 6.036 13.916 ;
  LAYER M2 ;
        RECT 3.564 13.948 6.036 13.98 ;
  LAYER M2 ;
        RECT 3.564 14.012 6.036 14.044 ;
  LAYER M2 ;
        RECT 3.564 14.076 6.036 14.108 ;
  LAYER M2 ;
        RECT 3.564 14.14 6.036 14.172 ;
  LAYER M2 ;
        RECT 3.564 14.204 6.036 14.236 ;
  LAYER M2 ;
        RECT 3.564 14.268 6.036 14.3 ;
  LAYER M2 ;
        RECT 3.564 14.332 6.036 14.364 ;
  LAYER M2 ;
        RECT 3.564 14.396 6.036 14.428 ;
  LAYER M2 ;
        RECT 3.564 14.46 6.036 14.492 ;
  LAYER M2 ;
        RECT 3.564 14.524 6.036 14.556 ;
  LAYER M2 ;
        RECT 3.564 14.588 6.036 14.62 ;
  LAYER M2 ;
        RECT 3.564 14.652 6.036 14.684 ;
  LAYER M2 ;
        RECT 3.564 14.716 6.036 14.748 ;
  LAYER M2 ;
        RECT 3.564 14.78 6.036 14.812 ;
  LAYER M2 ;
        RECT 3.564 14.844 6.036 14.876 ;
  LAYER M2 ;
        RECT 3.564 14.908 6.036 14.94 ;
  LAYER M2 ;
        RECT 3.564 14.972 6.036 15.004 ;
  LAYER M3 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M3 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M3 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M3 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M3 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M3 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M3 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M3 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M3 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M3 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M3 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M3 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M3 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M3 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M3 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M3 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M3 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M3 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M3 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M3 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M3 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M3 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M3 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M3 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M3 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M3 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M3 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M3 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M3 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M3 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M3 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M3 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M3 ;
        RECT 5.632 12.648 5.664 15.156 ;
  LAYER M3 ;
        RECT 5.696 12.648 5.728 15.156 ;
  LAYER M3 ;
        RECT 5.76 12.648 5.792 15.156 ;
  LAYER M3 ;
        RECT 5.824 12.648 5.856 15.156 ;
  LAYER M3 ;
        RECT 5.888 12.648 5.92 15.156 ;
  LAYER M3 ;
        RECT 5.984 12.648 6.016 15.156 ;
  LAYER M1 ;
        RECT 3.599 12.684 3.601 15.12 ;
  LAYER M1 ;
        RECT 3.679 12.684 3.681 15.12 ;
  LAYER M1 ;
        RECT 3.759 12.684 3.761 15.12 ;
  LAYER M1 ;
        RECT 3.839 12.684 3.841 15.12 ;
  LAYER M1 ;
        RECT 3.919 12.684 3.921 15.12 ;
  LAYER M1 ;
        RECT 3.999 12.684 4.001 15.12 ;
  LAYER M1 ;
        RECT 4.079 12.684 4.081 15.12 ;
  LAYER M1 ;
        RECT 4.159 12.684 4.161 15.12 ;
  LAYER M1 ;
        RECT 4.239 12.684 4.241 15.12 ;
  LAYER M1 ;
        RECT 4.319 12.684 4.321 15.12 ;
  LAYER M1 ;
        RECT 4.399 12.684 4.401 15.12 ;
  LAYER M1 ;
        RECT 4.479 12.684 4.481 15.12 ;
  LAYER M1 ;
        RECT 4.559 12.684 4.561 15.12 ;
  LAYER M1 ;
        RECT 4.639 12.684 4.641 15.12 ;
  LAYER M1 ;
        RECT 4.719 12.684 4.721 15.12 ;
  LAYER M1 ;
        RECT 4.799 12.684 4.801 15.12 ;
  LAYER M1 ;
        RECT 4.879 12.684 4.881 15.12 ;
  LAYER M1 ;
        RECT 4.959 12.684 4.961 15.12 ;
  LAYER M1 ;
        RECT 5.039 12.684 5.041 15.12 ;
  LAYER M1 ;
        RECT 5.119 12.684 5.121 15.12 ;
  LAYER M1 ;
        RECT 5.199 12.684 5.201 15.12 ;
  LAYER M1 ;
        RECT 5.279 12.684 5.281 15.12 ;
  LAYER M1 ;
        RECT 5.359 12.684 5.361 15.12 ;
  LAYER M1 ;
        RECT 5.439 12.684 5.441 15.12 ;
  LAYER M1 ;
        RECT 5.519 12.684 5.521 15.12 ;
  LAYER M1 ;
        RECT 5.599 12.684 5.601 15.12 ;
  LAYER M1 ;
        RECT 5.679 12.684 5.681 15.12 ;
  LAYER M1 ;
        RECT 5.759 12.684 5.761 15.12 ;
  LAYER M1 ;
        RECT 5.839 12.684 5.841 15.12 ;
  LAYER M1 ;
        RECT 5.919 12.684 5.921 15.12 ;
  LAYER M2 ;
        RECT 3.6 12.683 6 12.685 ;
  LAYER M2 ;
        RECT 3.6 12.767 6 12.769 ;
  LAYER M2 ;
        RECT 3.6 12.851 6 12.853 ;
  LAYER M2 ;
        RECT 3.6 12.935 6 12.937 ;
  LAYER M2 ;
        RECT 3.6 13.019 6 13.021 ;
  LAYER M2 ;
        RECT 3.6 13.103 6 13.105 ;
  LAYER M2 ;
        RECT 3.6 13.187 6 13.189 ;
  LAYER M2 ;
        RECT 3.6 13.271 6 13.273 ;
  LAYER M2 ;
        RECT 3.6 13.355 6 13.357 ;
  LAYER M2 ;
        RECT 3.6 13.439 6 13.441 ;
  LAYER M2 ;
        RECT 3.6 13.523 6 13.525 ;
  LAYER M2 ;
        RECT 3.6 13.607 6 13.609 ;
  LAYER M2 ;
        RECT 3.6 13.6905 6 13.6925 ;
  LAYER M2 ;
        RECT 3.6 13.775 6 13.777 ;
  LAYER M2 ;
        RECT 3.6 13.859 6 13.861 ;
  LAYER M2 ;
        RECT 3.6 13.943 6 13.945 ;
  LAYER M2 ;
        RECT 3.6 14.027 6 14.029 ;
  LAYER M2 ;
        RECT 3.6 14.111 6 14.113 ;
  LAYER M2 ;
        RECT 3.6 14.195 6 14.197 ;
  LAYER M2 ;
        RECT 3.6 14.279 6 14.281 ;
  LAYER M2 ;
        RECT 3.6 14.363 6 14.365 ;
  LAYER M2 ;
        RECT 3.6 14.447 6 14.449 ;
  LAYER M2 ;
        RECT 3.6 14.531 6 14.533 ;
  LAYER M2 ;
        RECT 3.6 14.615 6 14.617 ;
  LAYER M2 ;
        RECT 3.6 14.699 6 14.701 ;
  LAYER M2 ;
        RECT 3.6 14.783 6 14.785 ;
  LAYER M2 ;
        RECT 3.6 14.867 6 14.869 ;
  LAYER M2 ;
        RECT 3.6 14.951 6 14.953 ;
  LAYER M2 ;
        RECT 3.6 15.035 6 15.037 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M1 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M1 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M1 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M1 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M1 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M1 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M1 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M1 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M1 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M1 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M1 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M1 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M1 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M1 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M1 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M1 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M1 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M1 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M1 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M1 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M1 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M1 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M1 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M1 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M1 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M1 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M1 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M1 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M1 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M1 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M1 ;
        RECT 5.632 15.588 5.664 18.096 ;
  LAYER M1 ;
        RECT 5.696 15.588 5.728 18.096 ;
  LAYER M1 ;
        RECT 5.76 15.588 5.792 18.096 ;
  LAYER M1 ;
        RECT 5.824 15.588 5.856 18.096 ;
  LAYER M1 ;
        RECT 5.888 15.588 5.92 18.096 ;
  LAYER M2 ;
        RECT 3.564 15.672 6.036 15.704 ;
  LAYER M2 ;
        RECT 3.564 15.736 6.036 15.768 ;
  LAYER M2 ;
        RECT 3.564 15.8 6.036 15.832 ;
  LAYER M2 ;
        RECT 3.564 15.864 6.036 15.896 ;
  LAYER M2 ;
        RECT 3.564 15.928 6.036 15.96 ;
  LAYER M2 ;
        RECT 3.564 15.992 6.036 16.024 ;
  LAYER M2 ;
        RECT 3.564 16.056 6.036 16.088 ;
  LAYER M2 ;
        RECT 3.564 16.12 6.036 16.152 ;
  LAYER M2 ;
        RECT 3.564 16.184 6.036 16.216 ;
  LAYER M2 ;
        RECT 3.564 16.248 6.036 16.28 ;
  LAYER M2 ;
        RECT 3.564 16.312 6.036 16.344 ;
  LAYER M2 ;
        RECT 3.564 16.376 6.036 16.408 ;
  LAYER M2 ;
        RECT 3.564 16.44 6.036 16.472 ;
  LAYER M2 ;
        RECT 3.564 16.504 6.036 16.536 ;
  LAYER M2 ;
        RECT 3.564 16.568 6.036 16.6 ;
  LAYER M2 ;
        RECT 3.564 16.632 6.036 16.664 ;
  LAYER M2 ;
        RECT 3.564 16.696 6.036 16.728 ;
  LAYER M2 ;
        RECT 3.564 16.76 6.036 16.792 ;
  LAYER M2 ;
        RECT 3.564 16.824 6.036 16.856 ;
  LAYER M2 ;
        RECT 3.564 16.888 6.036 16.92 ;
  LAYER M2 ;
        RECT 3.564 16.952 6.036 16.984 ;
  LAYER M2 ;
        RECT 3.564 17.016 6.036 17.048 ;
  LAYER M2 ;
        RECT 3.564 17.08 6.036 17.112 ;
  LAYER M2 ;
        RECT 3.564 17.144 6.036 17.176 ;
  LAYER M2 ;
        RECT 3.564 17.208 6.036 17.24 ;
  LAYER M2 ;
        RECT 3.564 17.272 6.036 17.304 ;
  LAYER M2 ;
        RECT 3.564 17.336 6.036 17.368 ;
  LAYER M2 ;
        RECT 3.564 17.4 6.036 17.432 ;
  LAYER M2 ;
        RECT 3.564 17.464 6.036 17.496 ;
  LAYER M2 ;
        RECT 3.564 17.528 6.036 17.56 ;
  LAYER M2 ;
        RECT 3.564 17.592 6.036 17.624 ;
  LAYER M2 ;
        RECT 3.564 17.656 6.036 17.688 ;
  LAYER M2 ;
        RECT 3.564 17.72 6.036 17.752 ;
  LAYER M2 ;
        RECT 3.564 17.784 6.036 17.816 ;
  LAYER M2 ;
        RECT 3.564 17.848 6.036 17.88 ;
  LAYER M2 ;
        RECT 3.564 17.912 6.036 17.944 ;
  LAYER M3 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M3 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M3 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M3 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M3 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M3 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M3 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M3 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M3 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M3 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M3 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M3 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M3 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M3 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M3 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M3 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M3 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M3 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M3 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M3 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M3 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M3 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M3 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M3 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M3 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M3 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M3 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M3 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M3 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M3 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M3 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M3 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M3 ;
        RECT 5.632 15.588 5.664 18.096 ;
  LAYER M3 ;
        RECT 5.696 15.588 5.728 18.096 ;
  LAYER M3 ;
        RECT 5.76 15.588 5.792 18.096 ;
  LAYER M3 ;
        RECT 5.824 15.588 5.856 18.096 ;
  LAYER M3 ;
        RECT 5.888 15.588 5.92 18.096 ;
  LAYER M3 ;
        RECT 5.984 15.588 6.016 18.096 ;
  LAYER M1 ;
        RECT 3.599 15.624 3.601 18.06 ;
  LAYER M1 ;
        RECT 3.679 15.624 3.681 18.06 ;
  LAYER M1 ;
        RECT 3.759 15.624 3.761 18.06 ;
  LAYER M1 ;
        RECT 3.839 15.624 3.841 18.06 ;
  LAYER M1 ;
        RECT 3.919 15.624 3.921 18.06 ;
  LAYER M1 ;
        RECT 3.999 15.624 4.001 18.06 ;
  LAYER M1 ;
        RECT 4.079 15.624 4.081 18.06 ;
  LAYER M1 ;
        RECT 4.159 15.624 4.161 18.06 ;
  LAYER M1 ;
        RECT 4.239 15.624 4.241 18.06 ;
  LAYER M1 ;
        RECT 4.319 15.624 4.321 18.06 ;
  LAYER M1 ;
        RECT 4.399 15.624 4.401 18.06 ;
  LAYER M1 ;
        RECT 4.479 15.624 4.481 18.06 ;
  LAYER M1 ;
        RECT 4.559 15.624 4.561 18.06 ;
  LAYER M1 ;
        RECT 4.639 15.624 4.641 18.06 ;
  LAYER M1 ;
        RECT 4.719 15.624 4.721 18.06 ;
  LAYER M1 ;
        RECT 4.799 15.624 4.801 18.06 ;
  LAYER M1 ;
        RECT 4.879 15.624 4.881 18.06 ;
  LAYER M1 ;
        RECT 4.959 15.624 4.961 18.06 ;
  LAYER M1 ;
        RECT 5.039 15.624 5.041 18.06 ;
  LAYER M1 ;
        RECT 5.119 15.624 5.121 18.06 ;
  LAYER M1 ;
        RECT 5.199 15.624 5.201 18.06 ;
  LAYER M1 ;
        RECT 5.279 15.624 5.281 18.06 ;
  LAYER M1 ;
        RECT 5.359 15.624 5.361 18.06 ;
  LAYER M1 ;
        RECT 5.439 15.624 5.441 18.06 ;
  LAYER M1 ;
        RECT 5.519 15.624 5.521 18.06 ;
  LAYER M1 ;
        RECT 5.599 15.624 5.601 18.06 ;
  LAYER M1 ;
        RECT 5.679 15.624 5.681 18.06 ;
  LAYER M1 ;
        RECT 5.759 15.624 5.761 18.06 ;
  LAYER M1 ;
        RECT 5.839 15.624 5.841 18.06 ;
  LAYER M1 ;
        RECT 5.919 15.624 5.921 18.06 ;
  LAYER M2 ;
        RECT 3.6 15.623 6 15.625 ;
  LAYER M2 ;
        RECT 3.6 15.707 6 15.709 ;
  LAYER M2 ;
        RECT 3.6 15.791 6 15.793 ;
  LAYER M2 ;
        RECT 3.6 15.875 6 15.877 ;
  LAYER M2 ;
        RECT 3.6 15.959 6 15.961 ;
  LAYER M2 ;
        RECT 3.6 16.043 6 16.045 ;
  LAYER M2 ;
        RECT 3.6 16.127 6 16.129 ;
  LAYER M2 ;
        RECT 3.6 16.211 6 16.213 ;
  LAYER M2 ;
        RECT 3.6 16.295 6 16.297 ;
  LAYER M2 ;
        RECT 3.6 16.379 6 16.381 ;
  LAYER M2 ;
        RECT 3.6 16.463 6 16.465 ;
  LAYER M2 ;
        RECT 3.6 16.547 6 16.549 ;
  LAYER M2 ;
        RECT 3.6 16.6305 6 16.6325 ;
  LAYER M2 ;
        RECT 3.6 16.715 6 16.717 ;
  LAYER M2 ;
        RECT 3.6 16.799 6 16.801 ;
  LAYER M2 ;
        RECT 3.6 16.883 6 16.885 ;
  LAYER M2 ;
        RECT 3.6 16.967 6 16.969 ;
  LAYER M2 ;
        RECT 3.6 17.051 6 17.053 ;
  LAYER M2 ;
        RECT 3.6 17.135 6 17.137 ;
  LAYER M2 ;
        RECT 3.6 17.219 6 17.221 ;
  LAYER M2 ;
        RECT 3.6 17.303 6 17.305 ;
  LAYER M2 ;
        RECT 3.6 17.387 6 17.389 ;
  LAYER M2 ;
        RECT 3.6 17.471 6 17.473 ;
  LAYER M2 ;
        RECT 3.6 17.555 6 17.557 ;
  LAYER M2 ;
        RECT 3.6 17.639 6 17.641 ;
  LAYER M2 ;
        RECT 3.6 17.723 6 17.725 ;
  LAYER M2 ;
        RECT 3.6 17.807 6 17.809 ;
  LAYER M2 ;
        RECT 3.6 17.891 6 17.893 ;
  LAYER M2 ;
        RECT 3.6 17.975 6 17.977 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M1 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M1 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M1 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M1 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M1 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M1 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M1 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M1 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M1 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M1 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M1 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M1 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M1 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M1 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M1 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M1 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M1 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M1 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M1 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M1 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M1 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M1 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M1 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M1 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M1 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M1 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M1 ;
        RECT 8.832 0.888 8.864 3.396 ;
  LAYER M1 ;
        RECT 8.896 0.888 8.928 3.396 ;
  LAYER M1 ;
        RECT 8.96 0.888 8.992 3.396 ;
  LAYER M1 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M1 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M1 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M1 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M1 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M1 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M1 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M2 ;
        RECT 7.084 0.972 9.556 1.004 ;
  LAYER M2 ;
        RECT 7.084 1.036 9.556 1.068 ;
  LAYER M2 ;
        RECT 7.084 1.1 9.556 1.132 ;
  LAYER M2 ;
        RECT 7.084 1.164 9.556 1.196 ;
  LAYER M2 ;
        RECT 7.084 1.228 9.556 1.26 ;
  LAYER M2 ;
        RECT 7.084 1.292 9.556 1.324 ;
  LAYER M2 ;
        RECT 7.084 1.356 9.556 1.388 ;
  LAYER M2 ;
        RECT 7.084 1.42 9.556 1.452 ;
  LAYER M2 ;
        RECT 7.084 1.484 9.556 1.516 ;
  LAYER M2 ;
        RECT 7.084 1.548 9.556 1.58 ;
  LAYER M2 ;
        RECT 7.084 1.612 9.556 1.644 ;
  LAYER M2 ;
        RECT 7.084 1.676 9.556 1.708 ;
  LAYER M2 ;
        RECT 7.084 1.74 9.556 1.772 ;
  LAYER M2 ;
        RECT 7.084 1.804 9.556 1.836 ;
  LAYER M2 ;
        RECT 7.084 1.868 9.556 1.9 ;
  LAYER M2 ;
        RECT 7.084 1.932 9.556 1.964 ;
  LAYER M2 ;
        RECT 7.084 1.996 9.556 2.028 ;
  LAYER M2 ;
        RECT 7.084 2.06 9.556 2.092 ;
  LAYER M2 ;
        RECT 7.084 2.124 9.556 2.156 ;
  LAYER M2 ;
        RECT 7.084 2.188 9.556 2.22 ;
  LAYER M2 ;
        RECT 7.084 2.252 9.556 2.284 ;
  LAYER M2 ;
        RECT 7.084 2.316 9.556 2.348 ;
  LAYER M2 ;
        RECT 7.084 2.38 9.556 2.412 ;
  LAYER M2 ;
        RECT 7.084 2.444 9.556 2.476 ;
  LAYER M2 ;
        RECT 7.084 2.508 9.556 2.54 ;
  LAYER M2 ;
        RECT 7.084 2.572 9.556 2.604 ;
  LAYER M2 ;
        RECT 7.084 2.636 9.556 2.668 ;
  LAYER M2 ;
        RECT 7.084 2.7 9.556 2.732 ;
  LAYER M2 ;
        RECT 7.084 2.764 9.556 2.796 ;
  LAYER M2 ;
        RECT 7.084 2.828 9.556 2.86 ;
  LAYER M2 ;
        RECT 7.084 2.892 9.556 2.924 ;
  LAYER M2 ;
        RECT 7.084 2.956 9.556 2.988 ;
  LAYER M2 ;
        RECT 7.084 3.02 9.556 3.052 ;
  LAYER M2 ;
        RECT 7.084 3.084 9.556 3.116 ;
  LAYER M2 ;
        RECT 7.084 3.148 9.556 3.18 ;
  LAYER M2 ;
        RECT 7.084 3.212 9.556 3.244 ;
  LAYER M3 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M3 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M3 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M3 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M3 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M3 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M3 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M3 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M3 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M3 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M3 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M3 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M3 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M3 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M3 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M3 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M3 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M3 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M3 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M3 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M3 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M3 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M3 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M3 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M3 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M3 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M3 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M3 ;
        RECT 8.832 0.888 8.864 3.396 ;
  LAYER M3 ;
        RECT 8.896 0.888 8.928 3.396 ;
  LAYER M3 ;
        RECT 8.96 0.888 8.992 3.396 ;
  LAYER M3 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M3 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M3 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M3 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M3 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M3 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M3 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M3 ;
        RECT 9.504 0.888 9.536 3.396 ;
  LAYER M1 ;
        RECT 7.119 0.924 7.121 3.36 ;
  LAYER M1 ;
        RECT 7.199 0.924 7.201 3.36 ;
  LAYER M1 ;
        RECT 7.279 0.924 7.281 3.36 ;
  LAYER M1 ;
        RECT 7.359 0.924 7.361 3.36 ;
  LAYER M1 ;
        RECT 7.439 0.924 7.441 3.36 ;
  LAYER M1 ;
        RECT 7.519 0.924 7.521 3.36 ;
  LAYER M1 ;
        RECT 7.599 0.924 7.601 3.36 ;
  LAYER M1 ;
        RECT 7.679 0.924 7.681 3.36 ;
  LAYER M1 ;
        RECT 7.759 0.924 7.761 3.36 ;
  LAYER M1 ;
        RECT 7.839 0.924 7.841 3.36 ;
  LAYER M1 ;
        RECT 7.919 0.924 7.921 3.36 ;
  LAYER M1 ;
        RECT 7.999 0.924 8.001 3.36 ;
  LAYER M1 ;
        RECT 8.079 0.924 8.081 3.36 ;
  LAYER M1 ;
        RECT 8.159 0.924 8.161 3.36 ;
  LAYER M1 ;
        RECT 8.239 0.924 8.241 3.36 ;
  LAYER M1 ;
        RECT 8.319 0.924 8.321 3.36 ;
  LAYER M1 ;
        RECT 8.399 0.924 8.401 3.36 ;
  LAYER M1 ;
        RECT 8.479 0.924 8.481 3.36 ;
  LAYER M1 ;
        RECT 8.559 0.924 8.561 3.36 ;
  LAYER M1 ;
        RECT 8.639 0.924 8.641 3.36 ;
  LAYER M1 ;
        RECT 8.719 0.924 8.721 3.36 ;
  LAYER M1 ;
        RECT 8.799 0.924 8.801 3.36 ;
  LAYER M1 ;
        RECT 8.879 0.924 8.881 3.36 ;
  LAYER M1 ;
        RECT 8.959 0.924 8.961 3.36 ;
  LAYER M1 ;
        RECT 9.039 0.924 9.041 3.36 ;
  LAYER M1 ;
        RECT 9.119 0.924 9.121 3.36 ;
  LAYER M1 ;
        RECT 9.199 0.924 9.201 3.36 ;
  LAYER M1 ;
        RECT 9.279 0.924 9.281 3.36 ;
  LAYER M1 ;
        RECT 9.359 0.924 9.361 3.36 ;
  LAYER M1 ;
        RECT 9.439 0.924 9.441 3.36 ;
  LAYER M2 ;
        RECT 7.12 0.923 9.52 0.925 ;
  LAYER M2 ;
        RECT 7.12 1.007 9.52 1.009 ;
  LAYER M2 ;
        RECT 7.12 1.091 9.52 1.093 ;
  LAYER M2 ;
        RECT 7.12 1.175 9.52 1.177 ;
  LAYER M2 ;
        RECT 7.12 1.259 9.52 1.261 ;
  LAYER M2 ;
        RECT 7.12 1.343 9.52 1.345 ;
  LAYER M2 ;
        RECT 7.12 1.427 9.52 1.429 ;
  LAYER M2 ;
        RECT 7.12 1.511 9.52 1.513 ;
  LAYER M2 ;
        RECT 7.12 1.595 9.52 1.597 ;
  LAYER M2 ;
        RECT 7.12 1.679 9.52 1.681 ;
  LAYER M2 ;
        RECT 7.12 1.763 9.52 1.765 ;
  LAYER M2 ;
        RECT 7.12 1.847 9.52 1.849 ;
  LAYER M2 ;
        RECT 7.12 1.9305 9.52 1.9325 ;
  LAYER M2 ;
        RECT 7.12 2.015 9.52 2.017 ;
  LAYER M2 ;
        RECT 7.12 2.099 9.52 2.101 ;
  LAYER M2 ;
        RECT 7.12 2.183 9.52 2.185 ;
  LAYER M2 ;
        RECT 7.12 2.267 9.52 2.269 ;
  LAYER M2 ;
        RECT 7.12 2.351 9.52 2.353 ;
  LAYER M2 ;
        RECT 7.12 2.435 9.52 2.437 ;
  LAYER M2 ;
        RECT 7.12 2.519 9.52 2.521 ;
  LAYER M2 ;
        RECT 7.12 2.603 9.52 2.605 ;
  LAYER M2 ;
        RECT 7.12 2.687 9.52 2.689 ;
  LAYER M2 ;
        RECT 7.12 2.771 9.52 2.773 ;
  LAYER M2 ;
        RECT 7.12 2.855 9.52 2.857 ;
  LAYER M2 ;
        RECT 7.12 2.939 9.52 2.941 ;
  LAYER M2 ;
        RECT 7.12 3.023 9.52 3.025 ;
  LAYER M2 ;
        RECT 7.12 3.107 9.52 3.109 ;
  LAYER M2 ;
        RECT 7.12 3.191 9.52 3.193 ;
  LAYER M2 ;
        RECT 7.12 3.275 9.52 3.277 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M1 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M1 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M1 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M1 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M1 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M1 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M1 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M1 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M1 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M1 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M1 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M1 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M1 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M1 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M1 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M1 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M1 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M1 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M1 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M1 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M1 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M1 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M1 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M1 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M1 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M1 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M1 ;
        RECT 8.832 3.828 8.864 6.336 ;
  LAYER M1 ;
        RECT 8.896 3.828 8.928 6.336 ;
  LAYER M1 ;
        RECT 8.96 3.828 8.992 6.336 ;
  LAYER M1 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M1 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M1 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M1 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M1 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M1 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M1 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M2 ;
        RECT 7.084 3.912 9.556 3.944 ;
  LAYER M2 ;
        RECT 7.084 3.976 9.556 4.008 ;
  LAYER M2 ;
        RECT 7.084 4.04 9.556 4.072 ;
  LAYER M2 ;
        RECT 7.084 4.104 9.556 4.136 ;
  LAYER M2 ;
        RECT 7.084 4.168 9.556 4.2 ;
  LAYER M2 ;
        RECT 7.084 4.232 9.556 4.264 ;
  LAYER M2 ;
        RECT 7.084 4.296 9.556 4.328 ;
  LAYER M2 ;
        RECT 7.084 4.36 9.556 4.392 ;
  LAYER M2 ;
        RECT 7.084 4.424 9.556 4.456 ;
  LAYER M2 ;
        RECT 7.084 4.488 9.556 4.52 ;
  LAYER M2 ;
        RECT 7.084 4.552 9.556 4.584 ;
  LAYER M2 ;
        RECT 7.084 4.616 9.556 4.648 ;
  LAYER M2 ;
        RECT 7.084 4.68 9.556 4.712 ;
  LAYER M2 ;
        RECT 7.084 4.744 9.556 4.776 ;
  LAYER M2 ;
        RECT 7.084 4.808 9.556 4.84 ;
  LAYER M2 ;
        RECT 7.084 4.872 9.556 4.904 ;
  LAYER M2 ;
        RECT 7.084 4.936 9.556 4.968 ;
  LAYER M2 ;
        RECT 7.084 5 9.556 5.032 ;
  LAYER M2 ;
        RECT 7.084 5.064 9.556 5.096 ;
  LAYER M2 ;
        RECT 7.084 5.128 9.556 5.16 ;
  LAYER M2 ;
        RECT 7.084 5.192 9.556 5.224 ;
  LAYER M2 ;
        RECT 7.084 5.256 9.556 5.288 ;
  LAYER M2 ;
        RECT 7.084 5.32 9.556 5.352 ;
  LAYER M2 ;
        RECT 7.084 5.384 9.556 5.416 ;
  LAYER M2 ;
        RECT 7.084 5.448 9.556 5.48 ;
  LAYER M2 ;
        RECT 7.084 5.512 9.556 5.544 ;
  LAYER M2 ;
        RECT 7.084 5.576 9.556 5.608 ;
  LAYER M2 ;
        RECT 7.084 5.64 9.556 5.672 ;
  LAYER M2 ;
        RECT 7.084 5.704 9.556 5.736 ;
  LAYER M2 ;
        RECT 7.084 5.768 9.556 5.8 ;
  LAYER M2 ;
        RECT 7.084 5.832 9.556 5.864 ;
  LAYER M2 ;
        RECT 7.084 5.896 9.556 5.928 ;
  LAYER M2 ;
        RECT 7.084 5.96 9.556 5.992 ;
  LAYER M2 ;
        RECT 7.084 6.024 9.556 6.056 ;
  LAYER M2 ;
        RECT 7.084 6.088 9.556 6.12 ;
  LAYER M2 ;
        RECT 7.084 6.152 9.556 6.184 ;
  LAYER M3 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M3 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M3 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M3 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M3 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M3 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M3 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M3 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M3 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M3 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M3 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M3 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M3 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M3 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M3 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M3 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M3 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M3 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M3 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M3 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M3 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M3 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M3 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M3 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M3 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M3 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M3 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M3 ;
        RECT 8.832 3.828 8.864 6.336 ;
  LAYER M3 ;
        RECT 8.896 3.828 8.928 6.336 ;
  LAYER M3 ;
        RECT 8.96 3.828 8.992 6.336 ;
  LAYER M3 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M3 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M3 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M3 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M3 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M3 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M3 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M3 ;
        RECT 9.504 3.828 9.536 6.336 ;
  LAYER M1 ;
        RECT 7.119 3.864 7.121 6.3 ;
  LAYER M1 ;
        RECT 7.199 3.864 7.201 6.3 ;
  LAYER M1 ;
        RECT 7.279 3.864 7.281 6.3 ;
  LAYER M1 ;
        RECT 7.359 3.864 7.361 6.3 ;
  LAYER M1 ;
        RECT 7.439 3.864 7.441 6.3 ;
  LAYER M1 ;
        RECT 7.519 3.864 7.521 6.3 ;
  LAYER M1 ;
        RECT 7.599 3.864 7.601 6.3 ;
  LAYER M1 ;
        RECT 7.679 3.864 7.681 6.3 ;
  LAYER M1 ;
        RECT 7.759 3.864 7.761 6.3 ;
  LAYER M1 ;
        RECT 7.839 3.864 7.841 6.3 ;
  LAYER M1 ;
        RECT 7.919 3.864 7.921 6.3 ;
  LAYER M1 ;
        RECT 7.999 3.864 8.001 6.3 ;
  LAYER M1 ;
        RECT 8.079 3.864 8.081 6.3 ;
  LAYER M1 ;
        RECT 8.159 3.864 8.161 6.3 ;
  LAYER M1 ;
        RECT 8.239 3.864 8.241 6.3 ;
  LAYER M1 ;
        RECT 8.319 3.864 8.321 6.3 ;
  LAYER M1 ;
        RECT 8.399 3.864 8.401 6.3 ;
  LAYER M1 ;
        RECT 8.479 3.864 8.481 6.3 ;
  LAYER M1 ;
        RECT 8.559 3.864 8.561 6.3 ;
  LAYER M1 ;
        RECT 8.639 3.864 8.641 6.3 ;
  LAYER M1 ;
        RECT 8.719 3.864 8.721 6.3 ;
  LAYER M1 ;
        RECT 8.799 3.864 8.801 6.3 ;
  LAYER M1 ;
        RECT 8.879 3.864 8.881 6.3 ;
  LAYER M1 ;
        RECT 8.959 3.864 8.961 6.3 ;
  LAYER M1 ;
        RECT 9.039 3.864 9.041 6.3 ;
  LAYER M1 ;
        RECT 9.119 3.864 9.121 6.3 ;
  LAYER M1 ;
        RECT 9.199 3.864 9.201 6.3 ;
  LAYER M1 ;
        RECT 9.279 3.864 9.281 6.3 ;
  LAYER M1 ;
        RECT 9.359 3.864 9.361 6.3 ;
  LAYER M1 ;
        RECT 9.439 3.864 9.441 6.3 ;
  LAYER M2 ;
        RECT 7.12 3.863 9.52 3.865 ;
  LAYER M2 ;
        RECT 7.12 3.947 9.52 3.949 ;
  LAYER M2 ;
        RECT 7.12 4.031 9.52 4.033 ;
  LAYER M2 ;
        RECT 7.12 4.115 9.52 4.117 ;
  LAYER M2 ;
        RECT 7.12 4.199 9.52 4.201 ;
  LAYER M2 ;
        RECT 7.12 4.283 9.52 4.285 ;
  LAYER M2 ;
        RECT 7.12 4.367 9.52 4.369 ;
  LAYER M2 ;
        RECT 7.12 4.451 9.52 4.453 ;
  LAYER M2 ;
        RECT 7.12 4.535 9.52 4.537 ;
  LAYER M2 ;
        RECT 7.12 4.619 9.52 4.621 ;
  LAYER M2 ;
        RECT 7.12 4.703 9.52 4.705 ;
  LAYER M2 ;
        RECT 7.12 4.787 9.52 4.789 ;
  LAYER M2 ;
        RECT 7.12 4.8705 9.52 4.8725 ;
  LAYER M2 ;
        RECT 7.12 4.955 9.52 4.957 ;
  LAYER M2 ;
        RECT 7.12 5.039 9.52 5.041 ;
  LAYER M2 ;
        RECT 7.12 5.123 9.52 5.125 ;
  LAYER M2 ;
        RECT 7.12 5.207 9.52 5.209 ;
  LAYER M2 ;
        RECT 7.12 5.291 9.52 5.293 ;
  LAYER M2 ;
        RECT 7.12 5.375 9.52 5.377 ;
  LAYER M2 ;
        RECT 7.12 5.459 9.52 5.461 ;
  LAYER M2 ;
        RECT 7.12 5.543 9.52 5.545 ;
  LAYER M2 ;
        RECT 7.12 5.627 9.52 5.629 ;
  LAYER M2 ;
        RECT 7.12 5.711 9.52 5.713 ;
  LAYER M2 ;
        RECT 7.12 5.795 9.52 5.797 ;
  LAYER M2 ;
        RECT 7.12 5.879 9.52 5.881 ;
  LAYER M2 ;
        RECT 7.12 5.963 9.52 5.965 ;
  LAYER M2 ;
        RECT 7.12 6.047 9.52 6.049 ;
  LAYER M2 ;
        RECT 7.12 6.131 9.52 6.133 ;
  LAYER M2 ;
        RECT 7.12 6.215 9.52 6.217 ;
  LAYER M1 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M1 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M1 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M1 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M1 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M1 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M1 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M1 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M1 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M1 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M1 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M1 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M1 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M1 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M1 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M1 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M1 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M1 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M1 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M1 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M1 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M1 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M1 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M1 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M1 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M1 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M1 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M1 ;
        RECT 8.832 6.768 8.864 9.276 ;
  LAYER M1 ;
        RECT 8.896 6.768 8.928 9.276 ;
  LAYER M1 ;
        RECT 8.96 6.768 8.992 9.276 ;
  LAYER M1 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M1 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M1 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M1 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M1 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M1 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M1 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M2 ;
        RECT 7.084 6.852 9.556 6.884 ;
  LAYER M2 ;
        RECT 7.084 6.916 9.556 6.948 ;
  LAYER M2 ;
        RECT 7.084 6.98 9.556 7.012 ;
  LAYER M2 ;
        RECT 7.084 7.044 9.556 7.076 ;
  LAYER M2 ;
        RECT 7.084 7.108 9.556 7.14 ;
  LAYER M2 ;
        RECT 7.084 7.172 9.556 7.204 ;
  LAYER M2 ;
        RECT 7.084 7.236 9.556 7.268 ;
  LAYER M2 ;
        RECT 7.084 7.3 9.556 7.332 ;
  LAYER M2 ;
        RECT 7.084 7.364 9.556 7.396 ;
  LAYER M2 ;
        RECT 7.084 7.428 9.556 7.46 ;
  LAYER M2 ;
        RECT 7.084 7.492 9.556 7.524 ;
  LAYER M2 ;
        RECT 7.084 7.556 9.556 7.588 ;
  LAYER M2 ;
        RECT 7.084 7.62 9.556 7.652 ;
  LAYER M2 ;
        RECT 7.084 7.684 9.556 7.716 ;
  LAYER M2 ;
        RECT 7.084 7.748 9.556 7.78 ;
  LAYER M2 ;
        RECT 7.084 7.812 9.556 7.844 ;
  LAYER M2 ;
        RECT 7.084 7.876 9.556 7.908 ;
  LAYER M2 ;
        RECT 7.084 7.94 9.556 7.972 ;
  LAYER M2 ;
        RECT 7.084 8.004 9.556 8.036 ;
  LAYER M2 ;
        RECT 7.084 8.068 9.556 8.1 ;
  LAYER M2 ;
        RECT 7.084 8.132 9.556 8.164 ;
  LAYER M2 ;
        RECT 7.084 8.196 9.556 8.228 ;
  LAYER M2 ;
        RECT 7.084 8.26 9.556 8.292 ;
  LAYER M2 ;
        RECT 7.084 8.324 9.556 8.356 ;
  LAYER M2 ;
        RECT 7.084 8.388 9.556 8.42 ;
  LAYER M2 ;
        RECT 7.084 8.452 9.556 8.484 ;
  LAYER M2 ;
        RECT 7.084 8.516 9.556 8.548 ;
  LAYER M2 ;
        RECT 7.084 8.58 9.556 8.612 ;
  LAYER M2 ;
        RECT 7.084 8.644 9.556 8.676 ;
  LAYER M2 ;
        RECT 7.084 8.708 9.556 8.74 ;
  LAYER M2 ;
        RECT 7.084 8.772 9.556 8.804 ;
  LAYER M2 ;
        RECT 7.084 8.836 9.556 8.868 ;
  LAYER M2 ;
        RECT 7.084 8.9 9.556 8.932 ;
  LAYER M2 ;
        RECT 7.084 8.964 9.556 8.996 ;
  LAYER M2 ;
        RECT 7.084 9.028 9.556 9.06 ;
  LAYER M2 ;
        RECT 7.084 9.092 9.556 9.124 ;
  LAYER M3 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M3 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M3 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M3 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M3 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M3 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M3 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M3 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M3 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M3 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M3 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M3 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M3 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M3 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M3 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M3 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M3 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M3 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M3 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M3 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M3 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M3 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M3 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M3 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M3 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M3 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M3 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M3 ;
        RECT 8.832 6.768 8.864 9.276 ;
  LAYER M3 ;
        RECT 8.896 6.768 8.928 9.276 ;
  LAYER M3 ;
        RECT 8.96 6.768 8.992 9.276 ;
  LAYER M3 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M3 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M3 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M3 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M3 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M3 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M3 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M3 ;
        RECT 9.504 6.768 9.536 9.276 ;
  LAYER M1 ;
        RECT 7.119 6.804 7.121 9.24 ;
  LAYER M1 ;
        RECT 7.199 6.804 7.201 9.24 ;
  LAYER M1 ;
        RECT 7.279 6.804 7.281 9.24 ;
  LAYER M1 ;
        RECT 7.359 6.804 7.361 9.24 ;
  LAYER M1 ;
        RECT 7.439 6.804 7.441 9.24 ;
  LAYER M1 ;
        RECT 7.519 6.804 7.521 9.24 ;
  LAYER M1 ;
        RECT 7.599 6.804 7.601 9.24 ;
  LAYER M1 ;
        RECT 7.679 6.804 7.681 9.24 ;
  LAYER M1 ;
        RECT 7.759 6.804 7.761 9.24 ;
  LAYER M1 ;
        RECT 7.839 6.804 7.841 9.24 ;
  LAYER M1 ;
        RECT 7.919 6.804 7.921 9.24 ;
  LAYER M1 ;
        RECT 7.999 6.804 8.001 9.24 ;
  LAYER M1 ;
        RECT 8.079 6.804 8.081 9.24 ;
  LAYER M1 ;
        RECT 8.159 6.804 8.161 9.24 ;
  LAYER M1 ;
        RECT 8.239 6.804 8.241 9.24 ;
  LAYER M1 ;
        RECT 8.319 6.804 8.321 9.24 ;
  LAYER M1 ;
        RECT 8.399 6.804 8.401 9.24 ;
  LAYER M1 ;
        RECT 8.479 6.804 8.481 9.24 ;
  LAYER M1 ;
        RECT 8.559 6.804 8.561 9.24 ;
  LAYER M1 ;
        RECT 8.639 6.804 8.641 9.24 ;
  LAYER M1 ;
        RECT 8.719 6.804 8.721 9.24 ;
  LAYER M1 ;
        RECT 8.799 6.804 8.801 9.24 ;
  LAYER M1 ;
        RECT 8.879 6.804 8.881 9.24 ;
  LAYER M1 ;
        RECT 8.959 6.804 8.961 9.24 ;
  LAYER M1 ;
        RECT 9.039 6.804 9.041 9.24 ;
  LAYER M1 ;
        RECT 9.119 6.804 9.121 9.24 ;
  LAYER M1 ;
        RECT 9.199 6.804 9.201 9.24 ;
  LAYER M1 ;
        RECT 9.279 6.804 9.281 9.24 ;
  LAYER M1 ;
        RECT 9.359 6.804 9.361 9.24 ;
  LAYER M1 ;
        RECT 9.439 6.804 9.441 9.24 ;
  LAYER M2 ;
        RECT 7.12 6.803 9.52 6.805 ;
  LAYER M2 ;
        RECT 7.12 6.887 9.52 6.889 ;
  LAYER M2 ;
        RECT 7.12 6.971 9.52 6.973 ;
  LAYER M2 ;
        RECT 7.12 7.055 9.52 7.057 ;
  LAYER M2 ;
        RECT 7.12 7.139 9.52 7.141 ;
  LAYER M2 ;
        RECT 7.12 7.223 9.52 7.225 ;
  LAYER M2 ;
        RECT 7.12 7.307 9.52 7.309 ;
  LAYER M2 ;
        RECT 7.12 7.391 9.52 7.393 ;
  LAYER M2 ;
        RECT 7.12 7.475 9.52 7.477 ;
  LAYER M2 ;
        RECT 7.12 7.559 9.52 7.561 ;
  LAYER M2 ;
        RECT 7.12 7.643 9.52 7.645 ;
  LAYER M2 ;
        RECT 7.12 7.727 9.52 7.729 ;
  LAYER M2 ;
        RECT 7.12 7.8105 9.52 7.8125 ;
  LAYER M2 ;
        RECT 7.12 7.895 9.52 7.897 ;
  LAYER M2 ;
        RECT 7.12 7.979 9.52 7.981 ;
  LAYER M2 ;
        RECT 7.12 8.063 9.52 8.065 ;
  LAYER M2 ;
        RECT 7.12 8.147 9.52 8.149 ;
  LAYER M2 ;
        RECT 7.12 8.231 9.52 8.233 ;
  LAYER M2 ;
        RECT 7.12 8.315 9.52 8.317 ;
  LAYER M2 ;
        RECT 7.12 8.399 9.52 8.401 ;
  LAYER M2 ;
        RECT 7.12 8.483 9.52 8.485 ;
  LAYER M2 ;
        RECT 7.12 8.567 9.52 8.569 ;
  LAYER M2 ;
        RECT 7.12 8.651 9.52 8.653 ;
  LAYER M2 ;
        RECT 7.12 8.735 9.52 8.737 ;
  LAYER M2 ;
        RECT 7.12 8.819 9.52 8.821 ;
  LAYER M2 ;
        RECT 7.12 8.903 9.52 8.905 ;
  LAYER M2 ;
        RECT 7.12 8.987 9.52 8.989 ;
  LAYER M2 ;
        RECT 7.12 9.071 9.52 9.073 ;
  LAYER M2 ;
        RECT 7.12 9.155 9.52 9.157 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M1 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M1 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M1 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M1 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M1 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M1 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M1 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M1 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M1 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M1 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M1 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M1 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M1 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M1 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M1 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M1 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M1 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M1 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M1 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M1 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M1 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M1 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M1 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M1 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M1 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M1 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M1 ;
        RECT 8.832 9.708 8.864 12.216 ;
  LAYER M1 ;
        RECT 8.896 9.708 8.928 12.216 ;
  LAYER M1 ;
        RECT 8.96 9.708 8.992 12.216 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M1 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M1 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M1 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M1 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M1 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M1 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M2 ;
        RECT 7.084 9.792 9.556 9.824 ;
  LAYER M2 ;
        RECT 7.084 9.856 9.556 9.888 ;
  LAYER M2 ;
        RECT 7.084 9.92 9.556 9.952 ;
  LAYER M2 ;
        RECT 7.084 9.984 9.556 10.016 ;
  LAYER M2 ;
        RECT 7.084 10.048 9.556 10.08 ;
  LAYER M2 ;
        RECT 7.084 10.112 9.556 10.144 ;
  LAYER M2 ;
        RECT 7.084 10.176 9.556 10.208 ;
  LAYER M2 ;
        RECT 7.084 10.24 9.556 10.272 ;
  LAYER M2 ;
        RECT 7.084 10.304 9.556 10.336 ;
  LAYER M2 ;
        RECT 7.084 10.368 9.556 10.4 ;
  LAYER M2 ;
        RECT 7.084 10.432 9.556 10.464 ;
  LAYER M2 ;
        RECT 7.084 10.496 9.556 10.528 ;
  LAYER M2 ;
        RECT 7.084 10.56 9.556 10.592 ;
  LAYER M2 ;
        RECT 7.084 10.624 9.556 10.656 ;
  LAYER M2 ;
        RECT 7.084 10.688 9.556 10.72 ;
  LAYER M2 ;
        RECT 7.084 10.752 9.556 10.784 ;
  LAYER M2 ;
        RECT 7.084 10.816 9.556 10.848 ;
  LAYER M2 ;
        RECT 7.084 10.88 9.556 10.912 ;
  LAYER M2 ;
        RECT 7.084 10.944 9.556 10.976 ;
  LAYER M2 ;
        RECT 7.084 11.008 9.556 11.04 ;
  LAYER M2 ;
        RECT 7.084 11.072 9.556 11.104 ;
  LAYER M2 ;
        RECT 7.084 11.136 9.556 11.168 ;
  LAYER M2 ;
        RECT 7.084 11.2 9.556 11.232 ;
  LAYER M2 ;
        RECT 7.084 11.264 9.556 11.296 ;
  LAYER M2 ;
        RECT 7.084 11.328 9.556 11.36 ;
  LAYER M2 ;
        RECT 7.084 11.392 9.556 11.424 ;
  LAYER M2 ;
        RECT 7.084 11.456 9.556 11.488 ;
  LAYER M2 ;
        RECT 7.084 11.52 9.556 11.552 ;
  LAYER M2 ;
        RECT 7.084 11.584 9.556 11.616 ;
  LAYER M2 ;
        RECT 7.084 11.648 9.556 11.68 ;
  LAYER M2 ;
        RECT 7.084 11.712 9.556 11.744 ;
  LAYER M2 ;
        RECT 7.084 11.776 9.556 11.808 ;
  LAYER M2 ;
        RECT 7.084 11.84 9.556 11.872 ;
  LAYER M2 ;
        RECT 7.084 11.904 9.556 11.936 ;
  LAYER M2 ;
        RECT 7.084 11.968 9.556 12 ;
  LAYER M2 ;
        RECT 7.084 12.032 9.556 12.064 ;
  LAYER M3 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M3 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M3 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M3 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M3 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M3 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M3 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M3 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M3 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M3 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M3 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M3 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M3 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M3 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M3 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M3 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M3 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M3 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M3 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M3 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M3 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M3 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M3 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M3 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M3 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M3 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M3 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M3 ;
        RECT 8.832 9.708 8.864 12.216 ;
  LAYER M3 ;
        RECT 8.896 9.708 8.928 12.216 ;
  LAYER M3 ;
        RECT 8.96 9.708 8.992 12.216 ;
  LAYER M3 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M3 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M3 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M3 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M3 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M3 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M3 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M3 ;
        RECT 9.504 9.708 9.536 12.216 ;
  LAYER M1 ;
        RECT 7.119 9.744 7.121 12.18 ;
  LAYER M1 ;
        RECT 7.199 9.744 7.201 12.18 ;
  LAYER M1 ;
        RECT 7.279 9.744 7.281 12.18 ;
  LAYER M1 ;
        RECT 7.359 9.744 7.361 12.18 ;
  LAYER M1 ;
        RECT 7.439 9.744 7.441 12.18 ;
  LAYER M1 ;
        RECT 7.519 9.744 7.521 12.18 ;
  LAYER M1 ;
        RECT 7.599 9.744 7.601 12.18 ;
  LAYER M1 ;
        RECT 7.679 9.744 7.681 12.18 ;
  LAYER M1 ;
        RECT 7.759 9.744 7.761 12.18 ;
  LAYER M1 ;
        RECT 7.839 9.744 7.841 12.18 ;
  LAYER M1 ;
        RECT 7.919 9.744 7.921 12.18 ;
  LAYER M1 ;
        RECT 7.999 9.744 8.001 12.18 ;
  LAYER M1 ;
        RECT 8.079 9.744 8.081 12.18 ;
  LAYER M1 ;
        RECT 8.159 9.744 8.161 12.18 ;
  LAYER M1 ;
        RECT 8.239 9.744 8.241 12.18 ;
  LAYER M1 ;
        RECT 8.319 9.744 8.321 12.18 ;
  LAYER M1 ;
        RECT 8.399 9.744 8.401 12.18 ;
  LAYER M1 ;
        RECT 8.479 9.744 8.481 12.18 ;
  LAYER M1 ;
        RECT 8.559 9.744 8.561 12.18 ;
  LAYER M1 ;
        RECT 8.639 9.744 8.641 12.18 ;
  LAYER M1 ;
        RECT 8.719 9.744 8.721 12.18 ;
  LAYER M1 ;
        RECT 8.799 9.744 8.801 12.18 ;
  LAYER M1 ;
        RECT 8.879 9.744 8.881 12.18 ;
  LAYER M1 ;
        RECT 8.959 9.744 8.961 12.18 ;
  LAYER M1 ;
        RECT 9.039 9.744 9.041 12.18 ;
  LAYER M1 ;
        RECT 9.119 9.744 9.121 12.18 ;
  LAYER M1 ;
        RECT 9.199 9.744 9.201 12.18 ;
  LAYER M1 ;
        RECT 9.279 9.744 9.281 12.18 ;
  LAYER M1 ;
        RECT 9.359 9.744 9.361 12.18 ;
  LAYER M1 ;
        RECT 9.439 9.744 9.441 12.18 ;
  LAYER M2 ;
        RECT 7.12 9.743 9.52 9.745 ;
  LAYER M2 ;
        RECT 7.12 9.827 9.52 9.829 ;
  LAYER M2 ;
        RECT 7.12 9.911 9.52 9.913 ;
  LAYER M2 ;
        RECT 7.12 9.995 9.52 9.997 ;
  LAYER M2 ;
        RECT 7.12 10.079 9.52 10.081 ;
  LAYER M2 ;
        RECT 7.12 10.163 9.52 10.165 ;
  LAYER M2 ;
        RECT 7.12 10.247 9.52 10.249 ;
  LAYER M2 ;
        RECT 7.12 10.331 9.52 10.333 ;
  LAYER M2 ;
        RECT 7.12 10.415 9.52 10.417 ;
  LAYER M2 ;
        RECT 7.12 10.499 9.52 10.501 ;
  LAYER M2 ;
        RECT 7.12 10.583 9.52 10.585 ;
  LAYER M2 ;
        RECT 7.12 10.667 9.52 10.669 ;
  LAYER M2 ;
        RECT 7.12 10.7505 9.52 10.7525 ;
  LAYER M2 ;
        RECT 7.12 10.835 9.52 10.837 ;
  LAYER M2 ;
        RECT 7.12 10.919 9.52 10.921 ;
  LAYER M2 ;
        RECT 7.12 11.003 9.52 11.005 ;
  LAYER M2 ;
        RECT 7.12 11.087 9.52 11.089 ;
  LAYER M2 ;
        RECT 7.12 11.171 9.52 11.173 ;
  LAYER M2 ;
        RECT 7.12 11.255 9.52 11.257 ;
  LAYER M2 ;
        RECT 7.12 11.339 9.52 11.341 ;
  LAYER M2 ;
        RECT 7.12 11.423 9.52 11.425 ;
  LAYER M2 ;
        RECT 7.12 11.507 9.52 11.509 ;
  LAYER M2 ;
        RECT 7.12 11.591 9.52 11.593 ;
  LAYER M2 ;
        RECT 7.12 11.675 9.52 11.677 ;
  LAYER M2 ;
        RECT 7.12 11.759 9.52 11.761 ;
  LAYER M2 ;
        RECT 7.12 11.843 9.52 11.845 ;
  LAYER M2 ;
        RECT 7.12 11.927 9.52 11.929 ;
  LAYER M2 ;
        RECT 7.12 12.011 9.52 12.013 ;
  LAYER M2 ;
        RECT 7.12 12.095 9.52 12.097 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M1 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M1 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M1 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M1 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M1 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M1 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M1 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M1 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M1 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M1 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M1 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M1 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M1 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M1 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M1 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M1 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M1 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M1 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M1 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M1 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M1 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M1 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M1 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M1 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M1 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M1 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M1 ;
        RECT 8.832 12.648 8.864 15.156 ;
  LAYER M1 ;
        RECT 8.896 12.648 8.928 15.156 ;
  LAYER M1 ;
        RECT 8.96 12.648 8.992 15.156 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M1 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M1 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M1 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M1 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M1 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M1 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M2 ;
        RECT 7.084 12.732 9.556 12.764 ;
  LAYER M2 ;
        RECT 7.084 12.796 9.556 12.828 ;
  LAYER M2 ;
        RECT 7.084 12.86 9.556 12.892 ;
  LAYER M2 ;
        RECT 7.084 12.924 9.556 12.956 ;
  LAYER M2 ;
        RECT 7.084 12.988 9.556 13.02 ;
  LAYER M2 ;
        RECT 7.084 13.052 9.556 13.084 ;
  LAYER M2 ;
        RECT 7.084 13.116 9.556 13.148 ;
  LAYER M2 ;
        RECT 7.084 13.18 9.556 13.212 ;
  LAYER M2 ;
        RECT 7.084 13.244 9.556 13.276 ;
  LAYER M2 ;
        RECT 7.084 13.308 9.556 13.34 ;
  LAYER M2 ;
        RECT 7.084 13.372 9.556 13.404 ;
  LAYER M2 ;
        RECT 7.084 13.436 9.556 13.468 ;
  LAYER M2 ;
        RECT 7.084 13.5 9.556 13.532 ;
  LAYER M2 ;
        RECT 7.084 13.564 9.556 13.596 ;
  LAYER M2 ;
        RECT 7.084 13.628 9.556 13.66 ;
  LAYER M2 ;
        RECT 7.084 13.692 9.556 13.724 ;
  LAYER M2 ;
        RECT 7.084 13.756 9.556 13.788 ;
  LAYER M2 ;
        RECT 7.084 13.82 9.556 13.852 ;
  LAYER M2 ;
        RECT 7.084 13.884 9.556 13.916 ;
  LAYER M2 ;
        RECT 7.084 13.948 9.556 13.98 ;
  LAYER M2 ;
        RECT 7.084 14.012 9.556 14.044 ;
  LAYER M2 ;
        RECT 7.084 14.076 9.556 14.108 ;
  LAYER M2 ;
        RECT 7.084 14.14 9.556 14.172 ;
  LAYER M2 ;
        RECT 7.084 14.204 9.556 14.236 ;
  LAYER M2 ;
        RECT 7.084 14.268 9.556 14.3 ;
  LAYER M2 ;
        RECT 7.084 14.332 9.556 14.364 ;
  LAYER M2 ;
        RECT 7.084 14.396 9.556 14.428 ;
  LAYER M2 ;
        RECT 7.084 14.46 9.556 14.492 ;
  LAYER M2 ;
        RECT 7.084 14.524 9.556 14.556 ;
  LAYER M2 ;
        RECT 7.084 14.588 9.556 14.62 ;
  LAYER M2 ;
        RECT 7.084 14.652 9.556 14.684 ;
  LAYER M2 ;
        RECT 7.084 14.716 9.556 14.748 ;
  LAYER M2 ;
        RECT 7.084 14.78 9.556 14.812 ;
  LAYER M2 ;
        RECT 7.084 14.844 9.556 14.876 ;
  LAYER M2 ;
        RECT 7.084 14.908 9.556 14.94 ;
  LAYER M2 ;
        RECT 7.084 14.972 9.556 15.004 ;
  LAYER M3 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M3 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M3 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M3 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M3 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M3 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M3 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M3 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M3 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M3 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M3 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M3 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M3 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M3 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M3 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M3 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M3 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M3 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M3 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M3 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M3 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M3 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M3 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M3 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M3 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M3 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M3 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M3 ;
        RECT 8.832 12.648 8.864 15.156 ;
  LAYER M3 ;
        RECT 8.896 12.648 8.928 15.156 ;
  LAYER M3 ;
        RECT 8.96 12.648 8.992 15.156 ;
  LAYER M3 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M3 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M3 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M3 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M3 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M3 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M3 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M3 ;
        RECT 9.504 12.648 9.536 15.156 ;
  LAYER M1 ;
        RECT 7.119 12.684 7.121 15.12 ;
  LAYER M1 ;
        RECT 7.199 12.684 7.201 15.12 ;
  LAYER M1 ;
        RECT 7.279 12.684 7.281 15.12 ;
  LAYER M1 ;
        RECT 7.359 12.684 7.361 15.12 ;
  LAYER M1 ;
        RECT 7.439 12.684 7.441 15.12 ;
  LAYER M1 ;
        RECT 7.519 12.684 7.521 15.12 ;
  LAYER M1 ;
        RECT 7.599 12.684 7.601 15.12 ;
  LAYER M1 ;
        RECT 7.679 12.684 7.681 15.12 ;
  LAYER M1 ;
        RECT 7.759 12.684 7.761 15.12 ;
  LAYER M1 ;
        RECT 7.839 12.684 7.841 15.12 ;
  LAYER M1 ;
        RECT 7.919 12.684 7.921 15.12 ;
  LAYER M1 ;
        RECT 7.999 12.684 8.001 15.12 ;
  LAYER M1 ;
        RECT 8.079 12.684 8.081 15.12 ;
  LAYER M1 ;
        RECT 8.159 12.684 8.161 15.12 ;
  LAYER M1 ;
        RECT 8.239 12.684 8.241 15.12 ;
  LAYER M1 ;
        RECT 8.319 12.684 8.321 15.12 ;
  LAYER M1 ;
        RECT 8.399 12.684 8.401 15.12 ;
  LAYER M1 ;
        RECT 8.479 12.684 8.481 15.12 ;
  LAYER M1 ;
        RECT 8.559 12.684 8.561 15.12 ;
  LAYER M1 ;
        RECT 8.639 12.684 8.641 15.12 ;
  LAYER M1 ;
        RECT 8.719 12.684 8.721 15.12 ;
  LAYER M1 ;
        RECT 8.799 12.684 8.801 15.12 ;
  LAYER M1 ;
        RECT 8.879 12.684 8.881 15.12 ;
  LAYER M1 ;
        RECT 8.959 12.684 8.961 15.12 ;
  LAYER M1 ;
        RECT 9.039 12.684 9.041 15.12 ;
  LAYER M1 ;
        RECT 9.119 12.684 9.121 15.12 ;
  LAYER M1 ;
        RECT 9.199 12.684 9.201 15.12 ;
  LAYER M1 ;
        RECT 9.279 12.684 9.281 15.12 ;
  LAYER M1 ;
        RECT 9.359 12.684 9.361 15.12 ;
  LAYER M1 ;
        RECT 9.439 12.684 9.441 15.12 ;
  LAYER M2 ;
        RECT 7.12 12.683 9.52 12.685 ;
  LAYER M2 ;
        RECT 7.12 12.767 9.52 12.769 ;
  LAYER M2 ;
        RECT 7.12 12.851 9.52 12.853 ;
  LAYER M2 ;
        RECT 7.12 12.935 9.52 12.937 ;
  LAYER M2 ;
        RECT 7.12 13.019 9.52 13.021 ;
  LAYER M2 ;
        RECT 7.12 13.103 9.52 13.105 ;
  LAYER M2 ;
        RECT 7.12 13.187 9.52 13.189 ;
  LAYER M2 ;
        RECT 7.12 13.271 9.52 13.273 ;
  LAYER M2 ;
        RECT 7.12 13.355 9.52 13.357 ;
  LAYER M2 ;
        RECT 7.12 13.439 9.52 13.441 ;
  LAYER M2 ;
        RECT 7.12 13.523 9.52 13.525 ;
  LAYER M2 ;
        RECT 7.12 13.607 9.52 13.609 ;
  LAYER M2 ;
        RECT 7.12 13.6905 9.52 13.6925 ;
  LAYER M2 ;
        RECT 7.12 13.775 9.52 13.777 ;
  LAYER M2 ;
        RECT 7.12 13.859 9.52 13.861 ;
  LAYER M2 ;
        RECT 7.12 13.943 9.52 13.945 ;
  LAYER M2 ;
        RECT 7.12 14.027 9.52 14.029 ;
  LAYER M2 ;
        RECT 7.12 14.111 9.52 14.113 ;
  LAYER M2 ;
        RECT 7.12 14.195 9.52 14.197 ;
  LAYER M2 ;
        RECT 7.12 14.279 9.52 14.281 ;
  LAYER M2 ;
        RECT 7.12 14.363 9.52 14.365 ;
  LAYER M2 ;
        RECT 7.12 14.447 9.52 14.449 ;
  LAYER M2 ;
        RECT 7.12 14.531 9.52 14.533 ;
  LAYER M2 ;
        RECT 7.12 14.615 9.52 14.617 ;
  LAYER M2 ;
        RECT 7.12 14.699 9.52 14.701 ;
  LAYER M2 ;
        RECT 7.12 14.783 9.52 14.785 ;
  LAYER M2 ;
        RECT 7.12 14.867 9.52 14.869 ;
  LAYER M2 ;
        RECT 7.12 14.951 9.52 14.953 ;
  LAYER M2 ;
        RECT 7.12 15.035 9.52 15.037 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M1 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M1 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M1 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M1 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M1 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M1 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M1 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M1 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M1 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M1 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M1 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M1 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M1 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M1 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M1 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M1 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M1 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M1 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M1 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M1 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M1 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M1 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M1 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M1 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M1 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M1 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M1 ;
        RECT 8.832 15.588 8.864 18.096 ;
  LAYER M1 ;
        RECT 8.896 15.588 8.928 18.096 ;
  LAYER M1 ;
        RECT 8.96 15.588 8.992 18.096 ;
  LAYER M1 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M1 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M1 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M1 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M1 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M1 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M1 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M2 ;
        RECT 7.084 15.672 9.556 15.704 ;
  LAYER M2 ;
        RECT 7.084 15.736 9.556 15.768 ;
  LAYER M2 ;
        RECT 7.084 15.8 9.556 15.832 ;
  LAYER M2 ;
        RECT 7.084 15.864 9.556 15.896 ;
  LAYER M2 ;
        RECT 7.084 15.928 9.556 15.96 ;
  LAYER M2 ;
        RECT 7.084 15.992 9.556 16.024 ;
  LAYER M2 ;
        RECT 7.084 16.056 9.556 16.088 ;
  LAYER M2 ;
        RECT 7.084 16.12 9.556 16.152 ;
  LAYER M2 ;
        RECT 7.084 16.184 9.556 16.216 ;
  LAYER M2 ;
        RECT 7.084 16.248 9.556 16.28 ;
  LAYER M2 ;
        RECT 7.084 16.312 9.556 16.344 ;
  LAYER M2 ;
        RECT 7.084 16.376 9.556 16.408 ;
  LAYER M2 ;
        RECT 7.084 16.44 9.556 16.472 ;
  LAYER M2 ;
        RECT 7.084 16.504 9.556 16.536 ;
  LAYER M2 ;
        RECT 7.084 16.568 9.556 16.6 ;
  LAYER M2 ;
        RECT 7.084 16.632 9.556 16.664 ;
  LAYER M2 ;
        RECT 7.084 16.696 9.556 16.728 ;
  LAYER M2 ;
        RECT 7.084 16.76 9.556 16.792 ;
  LAYER M2 ;
        RECT 7.084 16.824 9.556 16.856 ;
  LAYER M2 ;
        RECT 7.084 16.888 9.556 16.92 ;
  LAYER M2 ;
        RECT 7.084 16.952 9.556 16.984 ;
  LAYER M2 ;
        RECT 7.084 17.016 9.556 17.048 ;
  LAYER M2 ;
        RECT 7.084 17.08 9.556 17.112 ;
  LAYER M2 ;
        RECT 7.084 17.144 9.556 17.176 ;
  LAYER M2 ;
        RECT 7.084 17.208 9.556 17.24 ;
  LAYER M2 ;
        RECT 7.084 17.272 9.556 17.304 ;
  LAYER M2 ;
        RECT 7.084 17.336 9.556 17.368 ;
  LAYER M2 ;
        RECT 7.084 17.4 9.556 17.432 ;
  LAYER M2 ;
        RECT 7.084 17.464 9.556 17.496 ;
  LAYER M2 ;
        RECT 7.084 17.528 9.556 17.56 ;
  LAYER M2 ;
        RECT 7.084 17.592 9.556 17.624 ;
  LAYER M2 ;
        RECT 7.084 17.656 9.556 17.688 ;
  LAYER M2 ;
        RECT 7.084 17.72 9.556 17.752 ;
  LAYER M2 ;
        RECT 7.084 17.784 9.556 17.816 ;
  LAYER M2 ;
        RECT 7.084 17.848 9.556 17.88 ;
  LAYER M2 ;
        RECT 7.084 17.912 9.556 17.944 ;
  LAYER M3 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M3 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M3 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M3 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M3 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M3 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M3 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M3 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M3 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M3 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M3 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M3 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M3 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M3 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M3 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M3 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M3 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M3 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M3 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M3 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M3 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M3 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M3 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M3 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M3 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M3 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M3 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M3 ;
        RECT 8.832 15.588 8.864 18.096 ;
  LAYER M3 ;
        RECT 8.896 15.588 8.928 18.096 ;
  LAYER M3 ;
        RECT 8.96 15.588 8.992 18.096 ;
  LAYER M3 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M3 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M3 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M3 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M3 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M3 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M3 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M3 ;
        RECT 9.504 15.588 9.536 18.096 ;
  LAYER M1 ;
        RECT 7.119 15.624 7.121 18.06 ;
  LAYER M1 ;
        RECT 7.199 15.624 7.201 18.06 ;
  LAYER M1 ;
        RECT 7.279 15.624 7.281 18.06 ;
  LAYER M1 ;
        RECT 7.359 15.624 7.361 18.06 ;
  LAYER M1 ;
        RECT 7.439 15.624 7.441 18.06 ;
  LAYER M1 ;
        RECT 7.519 15.624 7.521 18.06 ;
  LAYER M1 ;
        RECT 7.599 15.624 7.601 18.06 ;
  LAYER M1 ;
        RECT 7.679 15.624 7.681 18.06 ;
  LAYER M1 ;
        RECT 7.759 15.624 7.761 18.06 ;
  LAYER M1 ;
        RECT 7.839 15.624 7.841 18.06 ;
  LAYER M1 ;
        RECT 7.919 15.624 7.921 18.06 ;
  LAYER M1 ;
        RECT 7.999 15.624 8.001 18.06 ;
  LAYER M1 ;
        RECT 8.079 15.624 8.081 18.06 ;
  LAYER M1 ;
        RECT 8.159 15.624 8.161 18.06 ;
  LAYER M1 ;
        RECT 8.239 15.624 8.241 18.06 ;
  LAYER M1 ;
        RECT 8.319 15.624 8.321 18.06 ;
  LAYER M1 ;
        RECT 8.399 15.624 8.401 18.06 ;
  LAYER M1 ;
        RECT 8.479 15.624 8.481 18.06 ;
  LAYER M1 ;
        RECT 8.559 15.624 8.561 18.06 ;
  LAYER M1 ;
        RECT 8.639 15.624 8.641 18.06 ;
  LAYER M1 ;
        RECT 8.719 15.624 8.721 18.06 ;
  LAYER M1 ;
        RECT 8.799 15.624 8.801 18.06 ;
  LAYER M1 ;
        RECT 8.879 15.624 8.881 18.06 ;
  LAYER M1 ;
        RECT 8.959 15.624 8.961 18.06 ;
  LAYER M1 ;
        RECT 9.039 15.624 9.041 18.06 ;
  LAYER M1 ;
        RECT 9.119 15.624 9.121 18.06 ;
  LAYER M1 ;
        RECT 9.199 15.624 9.201 18.06 ;
  LAYER M1 ;
        RECT 9.279 15.624 9.281 18.06 ;
  LAYER M1 ;
        RECT 9.359 15.624 9.361 18.06 ;
  LAYER M1 ;
        RECT 9.439 15.624 9.441 18.06 ;
  LAYER M2 ;
        RECT 7.12 15.623 9.52 15.625 ;
  LAYER M2 ;
        RECT 7.12 15.707 9.52 15.709 ;
  LAYER M2 ;
        RECT 7.12 15.791 9.52 15.793 ;
  LAYER M2 ;
        RECT 7.12 15.875 9.52 15.877 ;
  LAYER M2 ;
        RECT 7.12 15.959 9.52 15.961 ;
  LAYER M2 ;
        RECT 7.12 16.043 9.52 16.045 ;
  LAYER M2 ;
        RECT 7.12 16.127 9.52 16.129 ;
  LAYER M2 ;
        RECT 7.12 16.211 9.52 16.213 ;
  LAYER M2 ;
        RECT 7.12 16.295 9.52 16.297 ;
  LAYER M2 ;
        RECT 7.12 16.379 9.52 16.381 ;
  LAYER M2 ;
        RECT 7.12 16.463 9.52 16.465 ;
  LAYER M2 ;
        RECT 7.12 16.547 9.52 16.549 ;
  LAYER M2 ;
        RECT 7.12 16.6305 9.52 16.6325 ;
  LAYER M2 ;
        RECT 7.12 16.715 9.52 16.717 ;
  LAYER M2 ;
        RECT 7.12 16.799 9.52 16.801 ;
  LAYER M2 ;
        RECT 7.12 16.883 9.52 16.885 ;
  LAYER M2 ;
        RECT 7.12 16.967 9.52 16.969 ;
  LAYER M2 ;
        RECT 7.12 17.051 9.52 17.053 ;
  LAYER M2 ;
        RECT 7.12 17.135 9.52 17.137 ;
  LAYER M2 ;
        RECT 7.12 17.219 9.52 17.221 ;
  LAYER M2 ;
        RECT 7.12 17.303 9.52 17.305 ;
  LAYER M2 ;
        RECT 7.12 17.387 9.52 17.389 ;
  LAYER M2 ;
        RECT 7.12 17.471 9.52 17.473 ;
  LAYER M2 ;
        RECT 7.12 17.555 9.52 17.557 ;
  LAYER M2 ;
        RECT 7.12 17.639 9.52 17.641 ;
  LAYER M2 ;
        RECT 7.12 17.723 9.52 17.725 ;
  LAYER M2 ;
        RECT 7.12 17.807 9.52 17.809 ;
  LAYER M2 ;
        RECT 7.12 17.891 9.52 17.893 ;
  LAYER M2 ;
        RECT 7.12 17.975 9.52 17.977 ;
  LAYER M1 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M1 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M1 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M1 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M1 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M1 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M1 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M1 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M1 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M1 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M1 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M1 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M1 ;
        RECT 11.392 0.888 11.424 3.396 ;
  LAYER M1 ;
        RECT 11.456 0.888 11.488 3.396 ;
  LAYER M1 ;
        RECT 11.52 0.888 11.552 3.396 ;
  LAYER M1 ;
        RECT 11.584 0.888 11.616 3.396 ;
  LAYER M1 ;
        RECT 11.648 0.888 11.68 3.396 ;
  LAYER M1 ;
        RECT 11.712 0.888 11.744 3.396 ;
  LAYER M1 ;
        RECT 11.776 0.888 11.808 3.396 ;
  LAYER M1 ;
        RECT 11.84 0.888 11.872 3.396 ;
  LAYER M1 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M1 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M1 ;
        RECT 12.032 0.888 12.064 3.396 ;
  LAYER M1 ;
        RECT 12.096 0.888 12.128 3.396 ;
  LAYER M1 ;
        RECT 12.16 0.888 12.192 3.396 ;
  LAYER M1 ;
        RECT 12.224 0.888 12.256 3.396 ;
  LAYER M1 ;
        RECT 12.288 0.888 12.32 3.396 ;
  LAYER M1 ;
        RECT 12.352 0.888 12.384 3.396 ;
  LAYER M1 ;
        RECT 12.416 0.888 12.448 3.396 ;
  LAYER M1 ;
        RECT 12.48 0.888 12.512 3.396 ;
  LAYER M1 ;
        RECT 12.544 0.888 12.576 3.396 ;
  LAYER M1 ;
        RECT 12.608 0.888 12.64 3.396 ;
  LAYER M1 ;
        RECT 12.672 0.888 12.704 3.396 ;
  LAYER M1 ;
        RECT 12.736 0.888 12.768 3.396 ;
  LAYER M1 ;
        RECT 12.8 0.888 12.832 3.396 ;
  LAYER M1 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M1 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M2 ;
        RECT 10.604 0.972 13.076 1.004 ;
  LAYER M2 ;
        RECT 10.604 1.036 13.076 1.068 ;
  LAYER M2 ;
        RECT 10.604 1.1 13.076 1.132 ;
  LAYER M2 ;
        RECT 10.604 1.164 13.076 1.196 ;
  LAYER M2 ;
        RECT 10.604 1.228 13.076 1.26 ;
  LAYER M2 ;
        RECT 10.604 1.292 13.076 1.324 ;
  LAYER M2 ;
        RECT 10.604 1.356 13.076 1.388 ;
  LAYER M2 ;
        RECT 10.604 1.42 13.076 1.452 ;
  LAYER M2 ;
        RECT 10.604 1.484 13.076 1.516 ;
  LAYER M2 ;
        RECT 10.604 1.548 13.076 1.58 ;
  LAYER M2 ;
        RECT 10.604 1.612 13.076 1.644 ;
  LAYER M2 ;
        RECT 10.604 1.676 13.076 1.708 ;
  LAYER M2 ;
        RECT 10.604 1.74 13.076 1.772 ;
  LAYER M2 ;
        RECT 10.604 1.804 13.076 1.836 ;
  LAYER M2 ;
        RECT 10.604 1.868 13.076 1.9 ;
  LAYER M2 ;
        RECT 10.604 1.932 13.076 1.964 ;
  LAYER M2 ;
        RECT 10.604 1.996 13.076 2.028 ;
  LAYER M2 ;
        RECT 10.604 2.06 13.076 2.092 ;
  LAYER M2 ;
        RECT 10.604 2.124 13.076 2.156 ;
  LAYER M2 ;
        RECT 10.604 2.188 13.076 2.22 ;
  LAYER M2 ;
        RECT 10.604 2.252 13.076 2.284 ;
  LAYER M2 ;
        RECT 10.604 2.316 13.076 2.348 ;
  LAYER M2 ;
        RECT 10.604 2.38 13.076 2.412 ;
  LAYER M2 ;
        RECT 10.604 2.444 13.076 2.476 ;
  LAYER M2 ;
        RECT 10.604 2.508 13.076 2.54 ;
  LAYER M2 ;
        RECT 10.604 2.572 13.076 2.604 ;
  LAYER M2 ;
        RECT 10.604 2.636 13.076 2.668 ;
  LAYER M2 ;
        RECT 10.604 2.7 13.076 2.732 ;
  LAYER M2 ;
        RECT 10.604 2.764 13.076 2.796 ;
  LAYER M2 ;
        RECT 10.604 2.828 13.076 2.86 ;
  LAYER M2 ;
        RECT 10.604 2.892 13.076 2.924 ;
  LAYER M2 ;
        RECT 10.604 2.956 13.076 2.988 ;
  LAYER M2 ;
        RECT 10.604 3.02 13.076 3.052 ;
  LAYER M2 ;
        RECT 10.604 3.084 13.076 3.116 ;
  LAYER M2 ;
        RECT 10.604 3.148 13.076 3.18 ;
  LAYER M2 ;
        RECT 10.604 3.212 13.076 3.244 ;
  LAYER M3 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M3 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M3 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M3 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M3 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M3 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M3 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M3 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M3 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M3 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M3 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M3 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M3 ;
        RECT 11.392 0.888 11.424 3.396 ;
  LAYER M3 ;
        RECT 11.456 0.888 11.488 3.396 ;
  LAYER M3 ;
        RECT 11.52 0.888 11.552 3.396 ;
  LAYER M3 ;
        RECT 11.584 0.888 11.616 3.396 ;
  LAYER M3 ;
        RECT 11.648 0.888 11.68 3.396 ;
  LAYER M3 ;
        RECT 11.712 0.888 11.744 3.396 ;
  LAYER M3 ;
        RECT 11.776 0.888 11.808 3.396 ;
  LAYER M3 ;
        RECT 11.84 0.888 11.872 3.396 ;
  LAYER M3 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M3 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M3 ;
        RECT 12.032 0.888 12.064 3.396 ;
  LAYER M3 ;
        RECT 12.096 0.888 12.128 3.396 ;
  LAYER M3 ;
        RECT 12.16 0.888 12.192 3.396 ;
  LAYER M3 ;
        RECT 12.224 0.888 12.256 3.396 ;
  LAYER M3 ;
        RECT 12.288 0.888 12.32 3.396 ;
  LAYER M3 ;
        RECT 12.352 0.888 12.384 3.396 ;
  LAYER M3 ;
        RECT 12.416 0.888 12.448 3.396 ;
  LAYER M3 ;
        RECT 12.48 0.888 12.512 3.396 ;
  LAYER M3 ;
        RECT 12.544 0.888 12.576 3.396 ;
  LAYER M3 ;
        RECT 12.608 0.888 12.64 3.396 ;
  LAYER M3 ;
        RECT 12.672 0.888 12.704 3.396 ;
  LAYER M3 ;
        RECT 12.736 0.888 12.768 3.396 ;
  LAYER M3 ;
        RECT 12.8 0.888 12.832 3.396 ;
  LAYER M3 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M3 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M3 ;
        RECT 13.024 0.888 13.056 3.396 ;
  LAYER M1 ;
        RECT 10.639 0.924 10.641 3.36 ;
  LAYER M1 ;
        RECT 10.719 0.924 10.721 3.36 ;
  LAYER M1 ;
        RECT 10.799 0.924 10.801 3.36 ;
  LAYER M1 ;
        RECT 10.879 0.924 10.881 3.36 ;
  LAYER M1 ;
        RECT 10.959 0.924 10.961 3.36 ;
  LAYER M1 ;
        RECT 11.039 0.924 11.041 3.36 ;
  LAYER M1 ;
        RECT 11.119 0.924 11.121 3.36 ;
  LAYER M1 ;
        RECT 11.199 0.924 11.201 3.36 ;
  LAYER M1 ;
        RECT 11.279 0.924 11.281 3.36 ;
  LAYER M1 ;
        RECT 11.359 0.924 11.361 3.36 ;
  LAYER M1 ;
        RECT 11.439 0.924 11.441 3.36 ;
  LAYER M1 ;
        RECT 11.519 0.924 11.521 3.36 ;
  LAYER M1 ;
        RECT 11.599 0.924 11.601 3.36 ;
  LAYER M1 ;
        RECT 11.679 0.924 11.681 3.36 ;
  LAYER M1 ;
        RECT 11.759 0.924 11.761 3.36 ;
  LAYER M1 ;
        RECT 11.839 0.924 11.841 3.36 ;
  LAYER M1 ;
        RECT 11.919 0.924 11.921 3.36 ;
  LAYER M1 ;
        RECT 11.999 0.924 12.001 3.36 ;
  LAYER M1 ;
        RECT 12.079 0.924 12.081 3.36 ;
  LAYER M1 ;
        RECT 12.159 0.924 12.161 3.36 ;
  LAYER M1 ;
        RECT 12.239 0.924 12.241 3.36 ;
  LAYER M1 ;
        RECT 12.319 0.924 12.321 3.36 ;
  LAYER M1 ;
        RECT 12.399 0.924 12.401 3.36 ;
  LAYER M1 ;
        RECT 12.479 0.924 12.481 3.36 ;
  LAYER M1 ;
        RECT 12.559 0.924 12.561 3.36 ;
  LAYER M1 ;
        RECT 12.639 0.924 12.641 3.36 ;
  LAYER M1 ;
        RECT 12.719 0.924 12.721 3.36 ;
  LAYER M1 ;
        RECT 12.799 0.924 12.801 3.36 ;
  LAYER M1 ;
        RECT 12.879 0.924 12.881 3.36 ;
  LAYER M1 ;
        RECT 12.959 0.924 12.961 3.36 ;
  LAYER M2 ;
        RECT 10.64 0.923 13.04 0.925 ;
  LAYER M2 ;
        RECT 10.64 1.007 13.04 1.009 ;
  LAYER M2 ;
        RECT 10.64 1.091 13.04 1.093 ;
  LAYER M2 ;
        RECT 10.64 1.175 13.04 1.177 ;
  LAYER M2 ;
        RECT 10.64 1.259 13.04 1.261 ;
  LAYER M2 ;
        RECT 10.64 1.343 13.04 1.345 ;
  LAYER M2 ;
        RECT 10.64 1.427 13.04 1.429 ;
  LAYER M2 ;
        RECT 10.64 1.511 13.04 1.513 ;
  LAYER M2 ;
        RECT 10.64 1.595 13.04 1.597 ;
  LAYER M2 ;
        RECT 10.64 1.679 13.04 1.681 ;
  LAYER M2 ;
        RECT 10.64 1.763 13.04 1.765 ;
  LAYER M2 ;
        RECT 10.64 1.847 13.04 1.849 ;
  LAYER M2 ;
        RECT 10.64 1.9305 13.04 1.9325 ;
  LAYER M2 ;
        RECT 10.64 2.015 13.04 2.017 ;
  LAYER M2 ;
        RECT 10.64 2.099 13.04 2.101 ;
  LAYER M2 ;
        RECT 10.64 2.183 13.04 2.185 ;
  LAYER M2 ;
        RECT 10.64 2.267 13.04 2.269 ;
  LAYER M2 ;
        RECT 10.64 2.351 13.04 2.353 ;
  LAYER M2 ;
        RECT 10.64 2.435 13.04 2.437 ;
  LAYER M2 ;
        RECT 10.64 2.519 13.04 2.521 ;
  LAYER M2 ;
        RECT 10.64 2.603 13.04 2.605 ;
  LAYER M2 ;
        RECT 10.64 2.687 13.04 2.689 ;
  LAYER M2 ;
        RECT 10.64 2.771 13.04 2.773 ;
  LAYER M2 ;
        RECT 10.64 2.855 13.04 2.857 ;
  LAYER M2 ;
        RECT 10.64 2.939 13.04 2.941 ;
  LAYER M2 ;
        RECT 10.64 3.023 13.04 3.025 ;
  LAYER M2 ;
        RECT 10.64 3.107 13.04 3.109 ;
  LAYER M2 ;
        RECT 10.64 3.191 13.04 3.193 ;
  LAYER M2 ;
        RECT 10.64 3.275 13.04 3.277 ;
  LAYER M1 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M1 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M1 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M1 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M1 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M1 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M1 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M1 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M1 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M1 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M1 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M1 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M1 ;
        RECT 11.392 3.828 11.424 6.336 ;
  LAYER M1 ;
        RECT 11.456 3.828 11.488 6.336 ;
  LAYER M1 ;
        RECT 11.52 3.828 11.552 6.336 ;
  LAYER M1 ;
        RECT 11.584 3.828 11.616 6.336 ;
  LAYER M1 ;
        RECT 11.648 3.828 11.68 6.336 ;
  LAYER M1 ;
        RECT 11.712 3.828 11.744 6.336 ;
  LAYER M1 ;
        RECT 11.776 3.828 11.808 6.336 ;
  LAYER M1 ;
        RECT 11.84 3.828 11.872 6.336 ;
  LAYER M1 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M1 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M1 ;
        RECT 12.032 3.828 12.064 6.336 ;
  LAYER M1 ;
        RECT 12.096 3.828 12.128 6.336 ;
  LAYER M1 ;
        RECT 12.16 3.828 12.192 6.336 ;
  LAYER M1 ;
        RECT 12.224 3.828 12.256 6.336 ;
  LAYER M1 ;
        RECT 12.288 3.828 12.32 6.336 ;
  LAYER M1 ;
        RECT 12.352 3.828 12.384 6.336 ;
  LAYER M1 ;
        RECT 12.416 3.828 12.448 6.336 ;
  LAYER M1 ;
        RECT 12.48 3.828 12.512 6.336 ;
  LAYER M1 ;
        RECT 12.544 3.828 12.576 6.336 ;
  LAYER M1 ;
        RECT 12.608 3.828 12.64 6.336 ;
  LAYER M1 ;
        RECT 12.672 3.828 12.704 6.336 ;
  LAYER M1 ;
        RECT 12.736 3.828 12.768 6.336 ;
  LAYER M1 ;
        RECT 12.8 3.828 12.832 6.336 ;
  LAYER M1 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M1 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M2 ;
        RECT 10.604 3.912 13.076 3.944 ;
  LAYER M2 ;
        RECT 10.604 3.976 13.076 4.008 ;
  LAYER M2 ;
        RECT 10.604 4.04 13.076 4.072 ;
  LAYER M2 ;
        RECT 10.604 4.104 13.076 4.136 ;
  LAYER M2 ;
        RECT 10.604 4.168 13.076 4.2 ;
  LAYER M2 ;
        RECT 10.604 4.232 13.076 4.264 ;
  LAYER M2 ;
        RECT 10.604 4.296 13.076 4.328 ;
  LAYER M2 ;
        RECT 10.604 4.36 13.076 4.392 ;
  LAYER M2 ;
        RECT 10.604 4.424 13.076 4.456 ;
  LAYER M2 ;
        RECT 10.604 4.488 13.076 4.52 ;
  LAYER M2 ;
        RECT 10.604 4.552 13.076 4.584 ;
  LAYER M2 ;
        RECT 10.604 4.616 13.076 4.648 ;
  LAYER M2 ;
        RECT 10.604 4.68 13.076 4.712 ;
  LAYER M2 ;
        RECT 10.604 4.744 13.076 4.776 ;
  LAYER M2 ;
        RECT 10.604 4.808 13.076 4.84 ;
  LAYER M2 ;
        RECT 10.604 4.872 13.076 4.904 ;
  LAYER M2 ;
        RECT 10.604 4.936 13.076 4.968 ;
  LAYER M2 ;
        RECT 10.604 5 13.076 5.032 ;
  LAYER M2 ;
        RECT 10.604 5.064 13.076 5.096 ;
  LAYER M2 ;
        RECT 10.604 5.128 13.076 5.16 ;
  LAYER M2 ;
        RECT 10.604 5.192 13.076 5.224 ;
  LAYER M2 ;
        RECT 10.604 5.256 13.076 5.288 ;
  LAYER M2 ;
        RECT 10.604 5.32 13.076 5.352 ;
  LAYER M2 ;
        RECT 10.604 5.384 13.076 5.416 ;
  LAYER M2 ;
        RECT 10.604 5.448 13.076 5.48 ;
  LAYER M2 ;
        RECT 10.604 5.512 13.076 5.544 ;
  LAYER M2 ;
        RECT 10.604 5.576 13.076 5.608 ;
  LAYER M2 ;
        RECT 10.604 5.64 13.076 5.672 ;
  LAYER M2 ;
        RECT 10.604 5.704 13.076 5.736 ;
  LAYER M2 ;
        RECT 10.604 5.768 13.076 5.8 ;
  LAYER M2 ;
        RECT 10.604 5.832 13.076 5.864 ;
  LAYER M2 ;
        RECT 10.604 5.896 13.076 5.928 ;
  LAYER M2 ;
        RECT 10.604 5.96 13.076 5.992 ;
  LAYER M2 ;
        RECT 10.604 6.024 13.076 6.056 ;
  LAYER M2 ;
        RECT 10.604 6.088 13.076 6.12 ;
  LAYER M2 ;
        RECT 10.604 6.152 13.076 6.184 ;
  LAYER M3 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M3 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M3 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M3 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M3 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M3 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M3 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M3 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M3 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M3 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M3 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M3 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M3 ;
        RECT 11.392 3.828 11.424 6.336 ;
  LAYER M3 ;
        RECT 11.456 3.828 11.488 6.336 ;
  LAYER M3 ;
        RECT 11.52 3.828 11.552 6.336 ;
  LAYER M3 ;
        RECT 11.584 3.828 11.616 6.336 ;
  LAYER M3 ;
        RECT 11.648 3.828 11.68 6.336 ;
  LAYER M3 ;
        RECT 11.712 3.828 11.744 6.336 ;
  LAYER M3 ;
        RECT 11.776 3.828 11.808 6.336 ;
  LAYER M3 ;
        RECT 11.84 3.828 11.872 6.336 ;
  LAYER M3 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M3 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M3 ;
        RECT 12.032 3.828 12.064 6.336 ;
  LAYER M3 ;
        RECT 12.096 3.828 12.128 6.336 ;
  LAYER M3 ;
        RECT 12.16 3.828 12.192 6.336 ;
  LAYER M3 ;
        RECT 12.224 3.828 12.256 6.336 ;
  LAYER M3 ;
        RECT 12.288 3.828 12.32 6.336 ;
  LAYER M3 ;
        RECT 12.352 3.828 12.384 6.336 ;
  LAYER M3 ;
        RECT 12.416 3.828 12.448 6.336 ;
  LAYER M3 ;
        RECT 12.48 3.828 12.512 6.336 ;
  LAYER M3 ;
        RECT 12.544 3.828 12.576 6.336 ;
  LAYER M3 ;
        RECT 12.608 3.828 12.64 6.336 ;
  LAYER M3 ;
        RECT 12.672 3.828 12.704 6.336 ;
  LAYER M3 ;
        RECT 12.736 3.828 12.768 6.336 ;
  LAYER M3 ;
        RECT 12.8 3.828 12.832 6.336 ;
  LAYER M3 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M3 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M3 ;
        RECT 13.024 3.828 13.056 6.336 ;
  LAYER M1 ;
        RECT 10.639 3.864 10.641 6.3 ;
  LAYER M1 ;
        RECT 10.719 3.864 10.721 6.3 ;
  LAYER M1 ;
        RECT 10.799 3.864 10.801 6.3 ;
  LAYER M1 ;
        RECT 10.879 3.864 10.881 6.3 ;
  LAYER M1 ;
        RECT 10.959 3.864 10.961 6.3 ;
  LAYER M1 ;
        RECT 11.039 3.864 11.041 6.3 ;
  LAYER M1 ;
        RECT 11.119 3.864 11.121 6.3 ;
  LAYER M1 ;
        RECT 11.199 3.864 11.201 6.3 ;
  LAYER M1 ;
        RECT 11.279 3.864 11.281 6.3 ;
  LAYER M1 ;
        RECT 11.359 3.864 11.361 6.3 ;
  LAYER M1 ;
        RECT 11.439 3.864 11.441 6.3 ;
  LAYER M1 ;
        RECT 11.519 3.864 11.521 6.3 ;
  LAYER M1 ;
        RECT 11.599 3.864 11.601 6.3 ;
  LAYER M1 ;
        RECT 11.679 3.864 11.681 6.3 ;
  LAYER M1 ;
        RECT 11.759 3.864 11.761 6.3 ;
  LAYER M1 ;
        RECT 11.839 3.864 11.841 6.3 ;
  LAYER M1 ;
        RECT 11.919 3.864 11.921 6.3 ;
  LAYER M1 ;
        RECT 11.999 3.864 12.001 6.3 ;
  LAYER M1 ;
        RECT 12.079 3.864 12.081 6.3 ;
  LAYER M1 ;
        RECT 12.159 3.864 12.161 6.3 ;
  LAYER M1 ;
        RECT 12.239 3.864 12.241 6.3 ;
  LAYER M1 ;
        RECT 12.319 3.864 12.321 6.3 ;
  LAYER M1 ;
        RECT 12.399 3.864 12.401 6.3 ;
  LAYER M1 ;
        RECT 12.479 3.864 12.481 6.3 ;
  LAYER M1 ;
        RECT 12.559 3.864 12.561 6.3 ;
  LAYER M1 ;
        RECT 12.639 3.864 12.641 6.3 ;
  LAYER M1 ;
        RECT 12.719 3.864 12.721 6.3 ;
  LAYER M1 ;
        RECT 12.799 3.864 12.801 6.3 ;
  LAYER M1 ;
        RECT 12.879 3.864 12.881 6.3 ;
  LAYER M1 ;
        RECT 12.959 3.864 12.961 6.3 ;
  LAYER M2 ;
        RECT 10.64 3.863 13.04 3.865 ;
  LAYER M2 ;
        RECT 10.64 3.947 13.04 3.949 ;
  LAYER M2 ;
        RECT 10.64 4.031 13.04 4.033 ;
  LAYER M2 ;
        RECT 10.64 4.115 13.04 4.117 ;
  LAYER M2 ;
        RECT 10.64 4.199 13.04 4.201 ;
  LAYER M2 ;
        RECT 10.64 4.283 13.04 4.285 ;
  LAYER M2 ;
        RECT 10.64 4.367 13.04 4.369 ;
  LAYER M2 ;
        RECT 10.64 4.451 13.04 4.453 ;
  LAYER M2 ;
        RECT 10.64 4.535 13.04 4.537 ;
  LAYER M2 ;
        RECT 10.64 4.619 13.04 4.621 ;
  LAYER M2 ;
        RECT 10.64 4.703 13.04 4.705 ;
  LAYER M2 ;
        RECT 10.64 4.787 13.04 4.789 ;
  LAYER M2 ;
        RECT 10.64 4.8705 13.04 4.8725 ;
  LAYER M2 ;
        RECT 10.64 4.955 13.04 4.957 ;
  LAYER M2 ;
        RECT 10.64 5.039 13.04 5.041 ;
  LAYER M2 ;
        RECT 10.64 5.123 13.04 5.125 ;
  LAYER M2 ;
        RECT 10.64 5.207 13.04 5.209 ;
  LAYER M2 ;
        RECT 10.64 5.291 13.04 5.293 ;
  LAYER M2 ;
        RECT 10.64 5.375 13.04 5.377 ;
  LAYER M2 ;
        RECT 10.64 5.459 13.04 5.461 ;
  LAYER M2 ;
        RECT 10.64 5.543 13.04 5.545 ;
  LAYER M2 ;
        RECT 10.64 5.627 13.04 5.629 ;
  LAYER M2 ;
        RECT 10.64 5.711 13.04 5.713 ;
  LAYER M2 ;
        RECT 10.64 5.795 13.04 5.797 ;
  LAYER M2 ;
        RECT 10.64 5.879 13.04 5.881 ;
  LAYER M2 ;
        RECT 10.64 5.963 13.04 5.965 ;
  LAYER M2 ;
        RECT 10.64 6.047 13.04 6.049 ;
  LAYER M2 ;
        RECT 10.64 6.131 13.04 6.133 ;
  LAYER M2 ;
        RECT 10.64 6.215 13.04 6.217 ;
  LAYER M1 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M1 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M1 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M1 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M1 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M1 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M1 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M1 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M1 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M1 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M1 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M1 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M1 ;
        RECT 11.392 6.768 11.424 9.276 ;
  LAYER M1 ;
        RECT 11.456 6.768 11.488 9.276 ;
  LAYER M1 ;
        RECT 11.52 6.768 11.552 9.276 ;
  LAYER M1 ;
        RECT 11.584 6.768 11.616 9.276 ;
  LAYER M1 ;
        RECT 11.648 6.768 11.68 9.276 ;
  LAYER M1 ;
        RECT 11.712 6.768 11.744 9.276 ;
  LAYER M1 ;
        RECT 11.776 6.768 11.808 9.276 ;
  LAYER M1 ;
        RECT 11.84 6.768 11.872 9.276 ;
  LAYER M1 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M1 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M1 ;
        RECT 12.032 6.768 12.064 9.276 ;
  LAYER M1 ;
        RECT 12.096 6.768 12.128 9.276 ;
  LAYER M1 ;
        RECT 12.16 6.768 12.192 9.276 ;
  LAYER M1 ;
        RECT 12.224 6.768 12.256 9.276 ;
  LAYER M1 ;
        RECT 12.288 6.768 12.32 9.276 ;
  LAYER M1 ;
        RECT 12.352 6.768 12.384 9.276 ;
  LAYER M1 ;
        RECT 12.416 6.768 12.448 9.276 ;
  LAYER M1 ;
        RECT 12.48 6.768 12.512 9.276 ;
  LAYER M1 ;
        RECT 12.544 6.768 12.576 9.276 ;
  LAYER M1 ;
        RECT 12.608 6.768 12.64 9.276 ;
  LAYER M1 ;
        RECT 12.672 6.768 12.704 9.276 ;
  LAYER M1 ;
        RECT 12.736 6.768 12.768 9.276 ;
  LAYER M1 ;
        RECT 12.8 6.768 12.832 9.276 ;
  LAYER M1 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M1 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M2 ;
        RECT 10.604 6.852 13.076 6.884 ;
  LAYER M2 ;
        RECT 10.604 6.916 13.076 6.948 ;
  LAYER M2 ;
        RECT 10.604 6.98 13.076 7.012 ;
  LAYER M2 ;
        RECT 10.604 7.044 13.076 7.076 ;
  LAYER M2 ;
        RECT 10.604 7.108 13.076 7.14 ;
  LAYER M2 ;
        RECT 10.604 7.172 13.076 7.204 ;
  LAYER M2 ;
        RECT 10.604 7.236 13.076 7.268 ;
  LAYER M2 ;
        RECT 10.604 7.3 13.076 7.332 ;
  LAYER M2 ;
        RECT 10.604 7.364 13.076 7.396 ;
  LAYER M2 ;
        RECT 10.604 7.428 13.076 7.46 ;
  LAYER M2 ;
        RECT 10.604 7.492 13.076 7.524 ;
  LAYER M2 ;
        RECT 10.604 7.556 13.076 7.588 ;
  LAYER M2 ;
        RECT 10.604 7.62 13.076 7.652 ;
  LAYER M2 ;
        RECT 10.604 7.684 13.076 7.716 ;
  LAYER M2 ;
        RECT 10.604 7.748 13.076 7.78 ;
  LAYER M2 ;
        RECT 10.604 7.812 13.076 7.844 ;
  LAYER M2 ;
        RECT 10.604 7.876 13.076 7.908 ;
  LAYER M2 ;
        RECT 10.604 7.94 13.076 7.972 ;
  LAYER M2 ;
        RECT 10.604 8.004 13.076 8.036 ;
  LAYER M2 ;
        RECT 10.604 8.068 13.076 8.1 ;
  LAYER M2 ;
        RECT 10.604 8.132 13.076 8.164 ;
  LAYER M2 ;
        RECT 10.604 8.196 13.076 8.228 ;
  LAYER M2 ;
        RECT 10.604 8.26 13.076 8.292 ;
  LAYER M2 ;
        RECT 10.604 8.324 13.076 8.356 ;
  LAYER M2 ;
        RECT 10.604 8.388 13.076 8.42 ;
  LAYER M2 ;
        RECT 10.604 8.452 13.076 8.484 ;
  LAYER M2 ;
        RECT 10.604 8.516 13.076 8.548 ;
  LAYER M2 ;
        RECT 10.604 8.58 13.076 8.612 ;
  LAYER M2 ;
        RECT 10.604 8.644 13.076 8.676 ;
  LAYER M2 ;
        RECT 10.604 8.708 13.076 8.74 ;
  LAYER M2 ;
        RECT 10.604 8.772 13.076 8.804 ;
  LAYER M2 ;
        RECT 10.604 8.836 13.076 8.868 ;
  LAYER M2 ;
        RECT 10.604 8.9 13.076 8.932 ;
  LAYER M2 ;
        RECT 10.604 8.964 13.076 8.996 ;
  LAYER M2 ;
        RECT 10.604 9.028 13.076 9.06 ;
  LAYER M2 ;
        RECT 10.604 9.092 13.076 9.124 ;
  LAYER M3 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M3 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M3 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M3 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M3 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M3 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M3 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M3 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M3 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M3 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M3 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M3 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M3 ;
        RECT 11.392 6.768 11.424 9.276 ;
  LAYER M3 ;
        RECT 11.456 6.768 11.488 9.276 ;
  LAYER M3 ;
        RECT 11.52 6.768 11.552 9.276 ;
  LAYER M3 ;
        RECT 11.584 6.768 11.616 9.276 ;
  LAYER M3 ;
        RECT 11.648 6.768 11.68 9.276 ;
  LAYER M3 ;
        RECT 11.712 6.768 11.744 9.276 ;
  LAYER M3 ;
        RECT 11.776 6.768 11.808 9.276 ;
  LAYER M3 ;
        RECT 11.84 6.768 11.872 9.276 ;
  LAYER M3 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M3 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M3 ;
        RECT 12.032 6.768 12.064 9.276 ;
  LAYER M3 ;
        RECT 12.096 6.768 12.128 9.276 ;
  LAYER M3 ;
        RECT 12.16 6.768 12.192 9.276 ;
  LAYER M3 ;
        RECT 12.224 6.768 12.256 9.276 ;
  LAYER M3 ;
        RECT 12.288 6.768 12.32 9.276 ;
  LAYER M3 ;
        RECT 12.352 6.768 12.384 9.276 ;
  LAYER M3 ;
        RECT 12.416 6.768 12.448 9.276 ;
  LAYER M3 ;
        RECT 12.48 6.768 12.512 9.276 ;
  LAYER M3 ;
        RECT 12.544 6.768 12.576 9.276 ;
  LAYER M3 ;
        RECT 12.608 6.768 12.64 9.276 ;
  LAYER M3 ;
        RECT 12.672 6.768 12.704 9.276 ;
  LAYER M3 ;
        RECT 12.736 6.768 12.768 9.276 ;
  LAYER M3 ;
        RECT 12.8 6.768 12.832 9.276 ;
  LAYER M3 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M3 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M3 ;
        RECT 13.024 6.768 13.056 9.276 ;
  LAYER M1 ;
        RECT 10.639 6.804 10.641 9.24 ;
  LAYER M1 ;
        RECT 10.719 6.804 10.721 9.24 ;
  LAYER M1 ;
        RECT 10.799 6.804 10.801 9.24 ;
  LAYER M1 ;
        RECT 10.879 6.804 10.881 9.24 ;
  LAYER M1 ;
        RECT 10.959 6.804 10.961 9.24 ;
  LAYER M1 ;
        RECT 11.039 6.804 11.041 9.24 ;
  LAYER M1 ;
        RECT 11.119 6.804 11.121 9.24 ;
  LAYER M1 ;
        RECT 11.199 6.804 11.201 9.24 ;
  LAYER M1 ;
        RECT 11.279 6.804 11.281 9.24 ;
  LAYER M1 ;
        RECT 11.359 6.804 11.361 9.24 ;
  LAYER M1 ;
        RECT 11.439 6.804 11.441 9.24 ;
  LAYER M1 ;
        RECT 11.519 6.804 11.521 9.24 ;
  LAYER M1 ;
        RECT 11.599 6.804 11.601 9.24 ;
  LAYER M1 ;
        RECT 11.679 6.804 11.681 9.24 ;
  LAYER M1 ;
        RECT 11.759 6.804 11.761 9.24 ;
  LAYER M1 ;
        RECT 11.839 6.804 11.841 9.24 ;
  LAYER M1 ;
        RECT 11.919 6.804 11.921 9.24 ;
  LAYER M1 ;
        RECT 11.999 6.804 12.001 9.24 ;
  LAYER M1 ;
        RECT 12.079 6.804 12.081 9.24 ;
  LAYER M1 ;
        RECT 12.159 6.804 12.161 9.24 ;
  LAYER M1 ;
        RECT 12.239 6.804 12.241 9.24 ;
  LAYER M1 ;
        RECT 12.319 6.804 12.321 9.24 ;
  LAYER M1 ;
        RECT 12.399 6.804 12.401 9.24 ;
  LAYER M1 ;
        RECT 12.479 6.804 12.481 9.24 ;
  LAYER M1 ;
        RECT 12.559 6.804 12.561 9.24 ;
  LAYER M1 ;
        RECT 12.639 6.804 12.641 9.24 ;
  LAYER M1 ;
        RECT 12.719 6.804 12.721 9.24 ;
  LAYER M1 ;
        RECT 12.799 6.804 12.801 9.24 ;
  LAYER M1 ;
        RECT 12.879 6.804 12.881 9.24 ;
  LAYER M1 ;
        RECT 12.959 6.804 12.961 9.24 ;
  LAYER M2 ;
        RECT 10.64 6.803 13.04 6.805 ;
  LAYER M2 ;
        RECT 10.64 6.887 13.04 6.889 ;
  LAYER M2 ;
        RECT 10.64 6.971 13.04 6.973 ;
  LAYER M2 ;
        RECT 10.64 7.055 13.04 7.057 ;
  LAYER M2 ;
        RECT 10.64 7.139 13.04 7.141 ;
  LAYER M2 ;
        RECT 10.64 7.223 13.04 7.225 ;
  LAYER M2 ;
        RECT 10.64 7.307 13.04 7.309 ;
  LAYER M2 ;
        RECT 10.64 7.391 13.04 7.393 ;
  LAYER M2 ;
        RECT 10.64 7.475 13.04 7.477 ;
  LAYER M2 ;
        RECT 10.64 7.559 13.04 7.561 ;
  LAYER M2 ;
        RECT 10.64 7.643 13.04 7.645 ;
  LAYER M2 ;
        RECT 10.64 7.727 13.04 7.729 ;
  LAYER M2 ;
        RECT 10.64 7.8105 13.04 7.8125 ;
  LAYER M2 ;
        RECT 10.64 7.895 13.04 7.897 ;
  LAYER M2 ;
        RECT 10.64 7.979 13.04 7.981 ;
  LAYER M2 ;
        RECT 10.64 8.063 13.04 8.065 ;
  LAYER M2 ;
        RECT 10.64 8.147 13.04 8.149 ;
  LAYER M2 ;
        RECT 10.64 8.231 13.04 8.233 ;
  LAYER M2 ;
        RECT 10.64 8.315 13.04 8.317 ;
  LAYER M2 ;
        RECT 10.64 8.399 13.04 8.401 ;
  LAYER M2 ;
        RECT 10.64 8.483 13.04 8.485 ;
  LAYER M2 ;
        RECT 10.64 8.567 13.04 8.569 ;
  LAYER M2 ;
        RECT 10.64 8.651 13.04 8.653 ;
  LAYER M2 ;
        RECT 10.64 8.735 13.04 8.737 ;
  LAYER M2 ;
        RECT 10.64 8.819 13.04 8.821 ;
  LAYER M2 ;
        RECT 10.64 8.903 13.04 8.905 ;
  LAYER M2 ;
        RECT 10.64 8.987 13.04 8.989 ;
  LAYER M2 ;
        RECT 10.64 9.071 13.04 9.073 ;
  LAYER M2 ;
        RECT 10.64 9.155 13.04 9.157 ;
  LAYER M1 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M1 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M1 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M1 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M1 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M1 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M1 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M1 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M1 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M1 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M1 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M1 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M1 ;
        RECT 11.392 9.708 11.424 12.216 ;
  LAYER M1 ;
        RECT 11.456 9.708 11.488 12.216 ;
  LAYER M1 ;
        RECT 11.52 9.708 11.552 12.216 ;
  LAYER M1 ;
        RECT 11.584 9.708 11.616 12.216 ;
  LAYER M1 ;
        RECT 11.648 9.708 11.68 12.216 ;
  LAYER M1 ;
        RECT 11.712 9.708 11.744 12.216 ;
  LAYER M1 ;
        RECT 11.776 9.708 11.808 12.216 ;
  LAYER M1 ;
        RECT 11.84 9.708 11.872 12.216 ;
  LAYER M1 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M1 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M1 ;
        RECT 12.032 9.708 12.064 12.216 ;
  LAYER M1 ;
        RECT 12.096 9.708 12.128 12.216 ;
  LAYER M1 ;
        RECT 12.16 9.708 12.192 12.216 ;
  LAYER M1 ;
        RECT 12.224 9.708 12.256 12.216 ;
  LAYER M1 ;
        RECT 12.288 9.708 12.32 12.216 ;
  LAYER M1 ;
        RECT 12.352 9.708 12.384 12.216 ;
  LAYER M1 ;
        RECT 12.416 9.708 12.448 12.216 ;
  LAYER M1 ;
        RECT 12.48 9.708 12.512 12.216 ;
  LAYER M1 ;
        RECT 12.544 9.708 12.576 12.216 ;
  LAYER M1 ;
        RECT 12.608 9.708 12.64 12.216 ;
  LAYER M1 ;
        RECT 12.672 9.708 12.704 12.216 ;
  LAYER M1 ;
        RECT 12.736 9.708 12.768 12.216 ;
  LAYER M1 ;
        RECT 12.8 9.708 12.832 12.216 ;
  LAYER M1 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M1 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M2 ;
        RECT 10.604 9.792 13.076 9.824 ;
  LAYER M2 ;
        RECT 10.604 9.856 13.076 9.888 ;
  LAYER M2 ;
        RECT 10.604 9.92 13.076 9.952 ;
  LAYER M2 ;
        RECT 10.604 9.984 13.076 10.016 ;
  LAYER M2 ;
        RECT 10.604 10.048 13.076 10.08 ;
  LAYER M2 ;
        RECT 10.604 10.112 13.076 10.144 ;
  LAYER M2 ;
        RECT 10.604 10.176 13.076 10.208 ;
  LAYER M2 ;
        RECT 10.604 10.24 13.076 10.272 ;
  LAYER M2 ;
        RECT 10.604 10.304 13.076 10.336 ;
  LAYER M2 ;
        RECT 10.604 10.368 13.076 10.4 ;
  LAYER M2 ;
        RECT 10.604 10.432 13.076 10.464 ;
  LAYER M2 ;
        RECT 10.604 10.496 13.076 10.528 ;
  LAYER M2 ;
        RECT 10.604 10.56 13.076 10.592 ;
  LAYER M2 ;
        RECT 10.604 10.624 13.076 10.656 ;
  LAYER M2 ;
        RECT 10.604 10.688 13.076 10.72 ;
  LAYER M2 ;
        RECT 10.604 10.752 13.076 10.784 ;
  LAYER M2 ;
        RECT 10.604 10.816 13.076 10.848 ;
  LAYER M2 ;
        RECT 10.604 10.88 13.076 10.912 ;
  LAYER M2 ;
        RECT 10.604 10.944 13.076 10.976 ;
  LAYER M2 ;
        RECT 10.604 11.008 13.076 11.04 ;
  LAYER M2 ;
        RECT 10.604 11.072 13.076 11.104 ;
  LAYER M2 ;
        RECT 10.604 11.136 13.076 11.168 ;
  LAYER M2 ;
        RECT 10.604 11.2 13.076 11.232 ;
  LAYER M2 ;
        RECT 10.604 11.264 13.076 11.296 ;
  LAYER M2 ;
        RECT 10.604 11.328 13.076 11.36 ;
  LAYER M2 ;
        RECT 10.604 11.392 13.076 11.424 ;
  LAYER M2 ;
        RECT 10.604 11.456 13.076 11.488 ;
  LAYER M2 ;
        RECT 10.604 11.52 13.076 11.552 ;
  LAYER M2 ;
        RECT 10.604 11.584 13.076 11.616 ;
  LAYER M2 ;
        RECT 10.604 11.648 13.076 11.68 ;
  LAYER M2 ;
        RECT 10.604 11.712 13.076 11.744 ;
  LAYER M2 ;
        RECT 10.604 11.776 13.076 11.808 ;
  LAYER M2 ;
        RECT 10.604 11.84 13.076 11.872 ;
  LAYER M2 ;
        RECT 10.604 11.904 13.076 11.936 ;
  LAYER M2 ;
        RECT 10.604 11.968 13.076 12 ;
  LAYER M2 ;
        RECT 10.604 12.032 13.076 12.064 ;
  LAYER M3 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M3 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M3 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M3 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M3 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M3 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M3 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M3 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M3 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M3 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M3 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M3 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M3 ;
        RECT 11.392 9.708 11.424 12.216 ;
  LAYER M3 ;
        RECT 11.456 9.708 11.488 12.216 ;
  LAYER M3 ;
        RECT 11.52 9.708 11.552 12.216 ;
  LAYER M3 ;
        RECT 11.584 9.708 11.616 12.216 ;
  LAYER M3 ;
        RECT 11.648 9.708 11.68 12.216 ;
  LAYER M3 ;
        RECT 11.712 9.708 11.744 12.216 ;
  LAYER M3 ;
        RECT 11.776 9.708 11.808 12.216 ;
  LAYER M3 ;
        RECT 11.84 9.708 11.872 12.216 ;
  LAYER M3 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M3 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M3 ;
        RECT 12.032 9.708 12.064 12.216 ;
  LAYER M3 ;
        RECT 12.096 9.708 12.128 12.216 ;
  LAYER M3 ;
        RECT 12.16 9.708 12.192 12.216 ;
  LAYER M3 ;
        RECT 12.224 9.708 12.256 12.216 ;
  LAYER M3 ;
        RECT 12.288 9.708 12.32 12.216 ;
  LAYER M3 ;
        RECT 12.352 9.708 12.384 12.216 ;
  LAYER M3 ;
        RECT 12.416 9.708 12.448 12.216 ;
  LAYER M3 ;
        RECT 12.48 9.708 12.512 12.216 ;
  LAYER M3 ;
        RECT 12.544 9.708 12.576 12.216 ;
  LAYER M3 ;
        RECT 12.608 9.708 12.64 12.216 ;
  LAYER M3 ;
        RECT 12.672 9.708 12.704 12.216 ;
  LAYER M3 ;
        RECT 12.736 9.708 12.768 12.216 ;
  LAYER M3 ;
        RECT 12.8 9.708 12.832 12.216 ;
  LAYER M3 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M3 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M3 ;
        RECT 13.024 9.708 13.056 12.216 ;
  LAYER M1 ;
        RECT 10.639 9.744 10.641 12.18 ;
  LAYER M1 ;
        RECT 10.719 9.744 10.721 12.18 ;
  LAYER M1 ;
        RECT 10.799 9.744 10.801 12.18 ;
  LAYER M1 ;
        RECT 10.879 9.744 10.881 12.18 ;
  LAYER M1 ;
        RECT 10.959 9.744 10.961 12.18 ;
  LAYER M1 ;
        RECT 11.039 9.744 11.041 12.18 ;
  LAYER M1 ;
        RECT 11.119 9.744 11.121 12.18 ;
  LAYER M1 ;
        RECT 11.199 9.744 11.201 12.18 ;
  LAYER M1 ;
        RECT 11.279 9.744 11.281 12.18 ;
  LAYER M1 ;
        RECT 11.359 9.744 11.361 12.18 ;
  LAYER M1 ;
        RECT 11.439 9.744 11.441 12.18 ;
  LAYER M1 ;
        RECT 11.519 9.744 11.521 12.18 ;
  LAYER M1 ;
        RECT 11.599 9.744 11.601 12.18 ;
  LAYER M1 ;
        RECT 11.679 9.744 11.681 12.18 ;
  LAYER M1 ;
        RECT 11.759 9.744 11.761 12.18 ;
  LAYER M1 ;
        RECT 11.839 9.744 11.841 12.18 ;
  LAYER M1 ;
        RECT 11.919 9.744 11.921 12.18 ;
  LAYER M1 ;
        RECT 11.999 9.744 12.001 12.18 ;
  LAYER M1 ;
        RECT 12.079 9.744 12.081 12.18 ;
  LAYER M1 ;
        RECT 12.159 9.744 12.161 12.18 ;
  LAYER M1 ;
        RECT 12.239 9.744 12.241 12.18 ;
  LAYER M1 ;
        RECT 12.319 9.744 12.321 12.18 ;
  LAYER M1 ;
        RECT 12.399 9.744 12.401 12.18 ;
  LAYER M1 ;
        RECT 12.479 9.744 12.481 12.18 ;
  LAYER M1 ;
        RECT 12.559 9.744 12.561 12.18 ;
  LAYER M1 ;
        RECT 12.639 9.744 12.641 12.18 ;
  LAYER M1 ;
        RECT 12.719 9.744 12.721 12.18 ;
  LAYER M1 ;
        RECT 12.799 9.744 12.801 12.18 ;
  LAYER M1 ;
        RECT 12.879 9.744 12.881 12.18 ;
  LAYER M1 ;
        RECT 12.959 9.744 12.961 12.18 ;
  LAYER M2 ;
        RECT 10.64 9.743 13.04 9.745 ;
  LAYER M2 ;
        RECT 10.64 9.827 13.04 9.829 ;
  LAYER M2 ;
        RECT 10.64 9.911 13.04 9.913 ;
  LAYER M2 ;
        RECT 10.64 9.995 13.04 9.997 ;
  LAYER M2 ;
        RECT 10.64 10.079 13.04 10.081 ;
  LAYER M2 ;
        RECT 10.64 10.163 13.04 10.165 ;
  LAYER M2 ;
        RECT 10.64 10.247 13.04 10.249 ;
  LAYER M2 ;
        RECT 10.64 10.331 13.04 10.333 ;
  LAYER M2 ;
        RECT 10.64 10.415 13.04 10.417 ;
  LAYER M2 ;
        RECT 10.64 10.499 13.04 10.501 ;
  LAYER M2 ;
        RECT 10.64 10.583 13.04 10.585 ;
  LAYER M2 ;
        RECT 10.64 10.667 13.04 10.669 ;
  LAYER M2 ;
        RECT 10.64 10.7505 13.04 10.7525 ;
  LAYER M2 ;
        RECT 10.64 10.835 13.04 10.837 ;
  LAYER M2 ;
        RECT 10.64 10.919 13.04 10.921 ;
  LAYER M2 ;
        RECT 10.64 11.003 13.04 11.005 ;
  LAYER M2 ;
        RECT 10.64 11.087 13.04 11.089 ;
  LAYER M2 ;
        RECT 10.64 11.171 13.04 11.173 ;
  LAYER M2 ;
        RECT 10.64 11.255 13.04 11.257 ;
  LAYER M2 ;
        RECT 10.64 11.339 13.04 11.341 ;
  LAYER M2 ;
        RECT 10.64 11.423 13.04 11.425 ;
  LAYER M2 ;
        RECT 10.64 11.507 13.04 11.509 ;
  LAYER M2 ;
        RECT 10.64 11.591 13.04 11.593 ;
  LAYER M2 ;
        RECT 10.64 11.675 13.04 11.677 ;
  LAYER M2 ;
        RECT 10.64 11.759 13.04 11.761 ;
  LAYER M2 ;
        RECT 10.64 11.843 13.04 11.845 ;
  LAYER M2 ;
        RECT 10.64 11.927 13.04 11.929 ;
  LAYER M2 ;
        RECT 10.64 12.011 13.04 12.013 ;
  LAYER M2 ;
        RECT 10.64 12.095 13.04 12.097 ;
  LAYER M1 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M1 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M1 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M1 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M1 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M1 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M1 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M1 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M1 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M1 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M1 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M1 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M1 ;
        RECT 11.392 12.648 11.424 15.156 ;
  LAYER M1 ;
        RECT 11.456 12.648 11.488 15.156 ;
  LAYER M1 ;
        RECT 11.52 12.648 11.552 15.156 ;
  LAYER M1 ;
        RECT 11.584 12.648 11.616 15.156 ;
  LAYER M1 ;
        RECT 11.648 12.648 11.68 15.156 ;
  LAYER M1 ;
        RECT 11.712 12.648 11.744 15.156 ;
  LAYER M1 ;
        RECT 11.776 12.648 11.808 15.156 ;
  LAYER M1 ;
        RECT 11.84 12.648 11.872 15.156 ;
  LAYER M1 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M1 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M1 ;
        RECT 12.032 12.648 12.064 15.156 ;
  LAYER M1 ;
        RECT 12.096 12.648 12.128 15.156 ;
  LAYER M1 ;
        RECT 12.16 12.648 12.192 15.156 ;
  LAYER M1 ;
        RECT 12.224 12.648 12.256 15.156 ;
  LAYER M1 ;
        RECT 12.288 12.648 12.32 15.156 ;
  LAYER M1 ;
        RECT 12.352 12.648 12.384 15.156 ;
  LAYER M1 ;
        RECT 12.416 12.648 12.448 15.156 ;
  LAYER M1 ;
        RECT 12.48 12.648 12.512 15.156 ;
  LAYER M1 ;
        RECT 12.544 12.648 12.576 15.156 ;
  LAYER M1 ;
        RECT 12.608 12.648 12.64 15.156 ;
  LAYER M1 ;
        RECT 12.672 12.648 12.704 15.156 ;
  LAYER M1 ;
        RECT 12.736 12.648 12.768 15.156 ;
  LAYER M1 ;
        RECT 12.8 12.648 12.832 15.156 ;
  LAYER M1 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M1 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M2 ;
        RECT 10.604 12.732 13.076 12.764 ;
  LAYER M2 ;
        RECT 10.604 12.796 13.076 12.828 ;
  LAYER M2 ;
        RECT 10.604 12.86 13.076 12.892 ;
  LAYER M2 ;
        RECT 10.604 12.924 13.076 12.956 ;
  LAYER M2 ;
        RECT 10.604 12.988 13.076 13.02 ;
  LAYER M2 ;
        RECT 10.604 13.052 13.076 13.084 ;
  LAYER M2 ;
        RECT 10.604 13.116 13.076 13.148 ;
  LAYER M2 ;
        RECT 10.604 13.18 13.076 13.212 ;
  LAYER M2 ;
        RECT 10.604 13.244 13.076 13.276 ;
  LAYER M2 ;
        RECT 10.604 13.308 13.076 13.34 ;
  LAYER M2 ;
        RECT 10.604 13.372 13.076 13.404 ;
  LAYER M2 ;
        RECT 10.604 13.436 13.076 13.468 ;
  LAYER M2 ;
        RECT 10.604 13.5 13.076 13.532 ;
  LAYER M2 ;
        RECT 10.604 13.564 13.076 13.596 ;
  LAYER M2 ;
        RECT 10.604 13.628 13.076 13.66 ;
  LAYER M2 ;
        RECT 10.604 13.692 13.076 13.724 ;
  LAYER M2 ;
        RECT 10.604 13.756 13.076 13.788 ;
  LAYER M2 ;
        RECT 10.604 13.82 13.076 13.852 ;
  LAYER M2 ;
        RECT 10.604 13.884 13.076 13.916 ;
  LAYER M2 ;
        RECT 10.604 13.948 13.076 13.98 ;
  LAYER M2 ;
        RECT 10.604 14.012 13.076 14.044 ;
  LAYER M2 ;
        RECT 10.604 14.076 13.076 14.108 ;
  LAYER M2 ;
        RECT 10.604 14.14 13.076 14.172 ;
  LAYER M2 ;
        RECT 10.604 14.204 13.076 14.236 ;
  LAYER M2 ;
        RECT 10.604 14.268 13.076 14.3 ;
  LAYER M2 ;
        RECT 10.604 14.332 13.076 14.364 ;
  LAYER M2 ;
        RECT 10.604 14.396 13.076 14.428 ;
  LAYER M2 ;
        RECT 10.604 14.46 13.076 14.492 ;
  LAYER M2 ;
        RECT 10.604 14.524 13.076 14.556 ;
  LAYER M2 ;
        RECT 10.604 14.588 13.076 14.62 ;
  LAYER M2 ;
        RECT 10.604 14.652 13.076 14.684 ;
  LAYER M2 ;
        RECT 10.604 14.716 13.076 14.748 ;
  LAYER M2 ;
        RECT 10.604 14.78 13.076 14.812 ;
  LAYER M2 ;
        RECT 10.604 14.844 13.076 14.876 ;
  LAYER M2 ;
        RECT 10.604 14.908 13.076 14.94 ;
  LAYER M2 ;
        RECT 10.604 14.972 13.076 15.004 ;
  LAYER M3 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M3 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M3 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M3 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M3 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M3 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M3 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M3 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M3 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M3 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M3 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M3 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M3 ;
        RECT 11.392 12.648 11.424 15.156 ;
  LAYER M3 ;
        RECT 11.456 12.648 11.488 15.156 ;
  LAYER M3 ;
        RECT 11.52 12.648 11.552 15.156 ;
  LAYER M3 ;
        RECT 11.584 12.648 11.616 15.156 ;
  LAYER M3 ;
        RECT 11.648 12.648 11.68 15.156 ;
  LAYER M3 ;
        RECT 11.712 12.648 11.744 15.156 ;
  LAYER M3 ;
        RECT 11.776 12.648 11.808 15.156 ;
  LAYER M3 ;
        RECT 11.84 12.648 11.872 15.156 ;
  LAYER M3 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M3 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M3 ;
        RECT 12.032 12.648 12.064 15.156 ;
  LAYER M3 ;
        RECT 12.096 12.648 12.128 15.156 ;
  LAYER M3 ;
        RECT 12.16 12.648 12.192 15.156 ;
  LAYER M3 ;
        RECT 12.224 12.648 12.256 15.156 ;
  LAYER M3 ;
        RECT 12.288 12.648 12.32 15.156 ;
  LAYER M3 ;
        RECT 12.352 12.648 12.384 15.156 ;
  LAYER M3 ;
        RECT 12.416 12.648 12.448 15.156 ;
  LAYER M3 ;
        RECT 12.48 12.648 12.512 15.156 ;
  LAYER M3 ;
        RECT 12.544 12.648 12.576 15.156 ;
  LAYER M3 ;
        RECT 12.608 12.648 12.64 15.156 ;
  LAYER M3 ;
        RECT 12.672 12.648 12.704 15.156 ;
  LAYER M3 ;
        RECT 12.736 12.648 12.768 15.156 ;
  LAYER M3 ;
        RECT 12.8 12.648 12.832 15.156 ;
  LAYER M3 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M3 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M3 ;
        RECT 13.024 12.648 13.056 15.156 ;
  LAYER M1 ;
        RECT 10.639 12.684 10.641 15.12 ;
  LAYER M1 ;
        RECT 10.719 12.684 10.721 15.12 ;
  LAYER M1 ;
        RECT 10.799 12.684 10.801 15.12 ;
  LAYER M1 ;
        RECT 10.879 12.684 10.881 15.12 ;
  LAYER M1 ;
        RECT 10.959 12.684 10.961 15.12 ;
  LAYER M1 ;
        RECT 11.039 12.684 11.041 15.12 ;
  LAYER M1 ;
        RECT 11.119 12.684 11.121 15.12 ;
  LAYER M1 ;
        RECT 11.199 12.684 11.201 15.12 ;
  LAYER M1 ;
        RECT 11.279 12.684 11.281 15.12 ;
  LAYER M1 ;
        RECT 11.359 12.684 11.361 15.12 ;
  LAYER M1 ;
        RECT 11.439 12.684 11.441 15.12 ;
  LAYER M1 ;
        RECT 11.519 12.684 11.521 15.12 ;
  LAYER M1 ;
        RECT 11.599 12.684 11.601 15.12 ;
  LAYER M1 ;
        RECT 11.679 12.684 11.681 15.12 ;
  LAYER M1 ;
        RECT 11.759 12.684 11.761 15.12 ;
  LAYER M1 ;
        RECT 11.839 12.684 11.841 15.12 ;
  LAYER M1 ;
        RECT 11.919 12.684 11.921 15.12 ;
  LAYER M1 ;
        RECT 11.999 12.684 12.001 15.12 ;
  LAYER M1 ;
        RECT 12.079 12.684 12.081 15.12 ;
  LAYER M1 ;
        RECT 12.159 12.684 12.161 15.12 ;
  LAYER M1 ;
        RECT 12.239 12.684 12.241 15.12 ;
  LAYER M1 ;
        RECT 12.319 12.684 12.321 15.12 ;
  LAYER M1 ;
        RECT 12.399 12.684 12.401 15.12 ;
  LAYER M1 ;
        RECT 12.479 12.684 12.481 15.12 ;
  LAYER M1 ;
        RECT 12.559 12.684 12.561 15.12 ;
  LAYER M1 ;
        RECT 12.639 12.684 12.641 15.12 ;
  LAYER M1 ;
        RECT 12.719 12.684 12.721 15.12 ;
  LAYER M1 ;
        RECT 12.799 12.684 12.801 15.12 ;
  LAYER M1 ;
        RECT 12.879 12.684 12.881 15.12 ;
  LAYER M1 ;
        RECT 12.959 12.684 12.961 15.12 ;
  LAYER M2 ;
        RECT 10.64 12.683 13.04 12.685 ;
  LAYER M2 ;
        RECT 10.64 12.767 13.04 12.769 ;
  LAYER M2 ;
        RECT 10.64 12.851 13.04 12.853 ;
  LAYER M2 ;
        RECT 10.64 12.935 13.04 12.937 ;
  LAYER M2 ;
        RECT 10.64 13.019 13.04 13.021 ;
  LAYER M2 ;
        RECT 10.64 13.103 13.04 13.105 ;
  LAYER M2 ;
        RECT 10.64 13.187 13.04 13.189 ;
  LAYER M2 ;
        RECT 10.64 13.271 13.04 13.273 ;
  LAYER M2 ;
        RECT 10.64 13.355 13.04 13.357 ;
  LAYER M2 ;
        RECT 10.64 13.439 13.04 13.441 ;
  LAYER M2 ;
        RECT 10.64 13.523 13.04 13.525 ;
  LAYER M2 ;
        RECT 10.64 13.607 13.04 13.609 ;
  LAYER M2 ;
        RECT 10.64 13.6905 13.04 13.6925 ;
  LAYER M2 ;
        RECT 10.64 13.775 13.04 13.777 ;
  LAYER M2 ;
        RECT 10.64 13.859 13.04 13.861 ;
  LAYER M2 ;
        RECT 10.64 13.943 13.04 13.945 ;
  LAYER M2 ;
        RECT 10.64 14.027 13.04 14.029 ;
  LAYER M2 ;
        RECT 10.64 14.111 13.04 14.113 ;
  LAYER M2 ;
        RECT 10.64 14.195 13.04 14.197 ;
  LAYER M2 ;
        RECT 10.64 14.279 13.04 14.281 ;
  LAYER M2 ;
        RECT 10.64 14.363 13.04 14.365 ;
  LAYER M2 ;
        RECT 10.64 14.447 13.04 14.449 ;
  LAYER M2 ;
        RECT 10.64 14.531 13.04 14.533 ;
  LAYER M2 ;
        RECT 10.64 14.615 13.04 14.617 ;
  LAYER M2 ;
        RECT 10.64 14.699 13.04 14.701 ;
  LAYER M2 ;
        RECT 10.64 14.783 13.04 14.785 ;
  LAYER M2 ;
        RECT 10.64 14.867 13.04 14.869 ;
  LAYER M2 ;
        RECT 10.64 14.951 13.04 14.953 ;
  LAYER M2 ;
        RECT 10.64 15.035 13.04 15.037 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M1 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M1 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M1 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M1 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M1 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M1 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M1 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M1 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M1 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M1 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M1 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M1 ;
        RECT 11.392 15.588 11.424 18.096 ;
  LAYER M1 ;
        RECT 11.456 15.588 11.488 18.096 ;
  LAYER M1 ;
        RECT 11.52 15.588 11.552 18.096 ;
  LAYER M1 ;
        RECT 11.584 15.588 11.616 18.096 ;
  LAYER M1 ;
        RECT 11.648 15.588 11.68 18.096 ;
  LAYER M1 ;
        RECT 11.712 15.588 11.744 18.096 ;
  LAYER M1 ;
        RECT 11.776 15.588 11.808 18.096 ;
  LAYER M1 ;
        RECT 11.84 15.588 11.872 18.096 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M1 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M1 ;
        RECT 12.032 15.588 12.064 18.096 ;
  LAYER M1 ;
        RECT 12.096 15.588 12.128 18.096 ;
  LAYER M1 ;
        RECT 12.16 15.588 12.192 18.096 ;
  LAYER M1 ;
        RECT 12.224 15.588 12.256 18.096 ;
  LAYER M1 ;
        RECT 12.288 15.588 12.32 18.096 ;
  LAYER M1 ;
        RECT 12.352 15.588 12.384 18.096 ;
  LAYER M1 ;
        RECT 12.416 15.588 12.448 18.096 ;
  LAYER M1 ;
        RECT 12.48 15.588 12.512 18.096 ;
  LAYER M1 ;
        RECT 12.544 15.588 12.576 18.096 ;
  LAYER M1 ;
        RECT 12.608 15.588 12.64 18.096 ;
  LAYER M1 ;
        RECT 12.672 15.588 12.704 18.096 ;
  LAYER M1 ;
        RECT 12.736 15.588 12.768 18.096 ;
  LAYER M1 ;
        RECT 12.8 15.588 12.832 18.096 ;
  LAYER M1 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M1 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M2 ;
        RECT 10.604 15.672 13.076 15.704 ;
  LAYER M2 ;
        RECT 10.604 15.736 13.076 15.768 ;
  LAYER M2 ;
        RECT 10.604 15.8 13.076 15.832 ;
  LAYER M2 ;
        RECT 10.604 15.864 13.076 15.896 ;
  LAYER M2 ;
        RECT 10.604 15.928 13.076 15.96 ;
  LAYER M2 ;
        RECT 10.604 15.992 13.076 16.024 ;
  LAYER M2 ;
        RECT 10.604 16.056 13.076 16.088 ;
  LAYER M2 ;
        RECT 10.604 16.12 13.076 16.152 ;
  LAYER M2 ;
        RECT 10.604 16.184 13.076 16.216 ;
  LAYER M2 ;
        RECT 10.604 16.248 13.076 16.28 ;
  LAYER M2 ;
        RECT 10.604 16.312 13.076 16.344 ;
  LAYER M2 ;
        RECT 10.604 16.376 13.076 16.408 ;
  LAYER M2 ;
        RECT 10.604 16.44 13.076 16.472 ;
  LAYER M2 ;
        RECT 10.604 16.504 13.076 16.536 ;
  LAYER M2 ;
        RECT 10.604 16.568 13.076 16.6 ;
  LAYER M2 ;
        RECT 10.604 16.632 13.076 16.664 ;
  LAYER M2 ;
        RECT 10.604 16.696 13.076 16.728 ;
  LAYER M2 ;
        RECT 10.604 16.76 13.076 16.792 ;
  LAYER M2 ;
        RECT 10.604 16.824 13.076 16.856 ;
  LAYER M2 ;
        RECT 10.604 16.888 13.076 16.92 ;
  LAYER M2 ;
        RECT 10.604 16.952 13.076 16.984 ;
  LAYER M2 ;
        RECT 10.604 17.016 13.076 17.048 ;
  LAYER M2 ;
        RECT 10.604 17.08 13.076 17.112 ;
  LAYER M2 ;
        RECT 10.604 17.144 13.076 17.176 ;
  LAYER M2 ;
        RECT 10.604 17.208 13.076 17.24 ;
  LAYER M2 ;
        RECT 10.604 17.272 13.076 17.304 ;
  LAYER M2 ;
        RECT 10.604 17.336 13.076 17.368 ;
  LAYER M2 ;
        RECT 10.604 17.4 13.076 17.432 ;
  LAYER M2 ;
        RECT 10.604 17.464 13.076 17.496 ;
  LAYER M2 ;
        RECT 10.604 17.528 13.076 17.56 ;
  LAYER M2 ;
        RECT 10.604 17.592 13.076 17.624 ;
  LAYER M2 ;
        RECT 10.604 17.656 13.076 17.688 ;
  LAYER M2 ;
        RECT 10.604 17.72 13.076 17.752 ;
  LAYER M2 ;
        RECT 10.604 17.784 13.076 17.816 ;
  LAYER M2 ;
        RECT 10.604 17.848 13.076 17.88 ;
  LAYER M2 ;
        RECT 10.604 17.912 13.076 17.944 ;
  LAYER M3 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M3 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M3 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M3 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M3 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M3 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M3 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M3 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M3 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M3 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M3 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M3 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M3 ;
        RECT 11.392 15.588 11.424 18.096 ;
  LAYER M3 ;
        RECT 11.456 15.588 11.488 18.096 ;
  LAYER M3 ;
        RECT 11.52 15.588 11.552 18.096 ;
  LAYER M3 ;
        RECT 11.584 15.588 11.616 18.096 ;
  LAYER M3 ;
        RECT 11.648 15.588 11.68 18.096 ;
  LAYER M3 ;
        RECT 11.712 15.588 11.744 18.096 ;
  LAYER M3 ;
        RECT 11.776 15.588 11.808 18.096 ;
  LAYER M3 ;
        RECT 11.84 15.588 11.872 18.096 ;
  LAYER M3 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M3 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M3 ;
        RECT 12.032 15.588 12.064 18.096 ;
  LAYER M3 ;
        RECT 12.096 15.588 12.128 18.096 ;
  LAYER M3 ;
        RECT 12.16 15.588 12.192 18.096 ;
  LAYER M3 ;
        RECT 12.224 15.588 12.256 18.096 ;
  LAYER M3 ;
        RECT 12.288 15.588 12.32 18.096 ;
  LAYER M3 ;
        RECT 12.352 15.588 12.384 18.096 ;
  LAYER M3 ;
        RECT 12.416 15.588 12.448 18.096 ;
  LAYER M3 ;
        RECT 12.48 15.588 12.512 18.096 ;
  LAYER M3 ;
        RECT 12.544 15.588 12.576 18.096 ;
  LAYER M3 ;
        RECT 12.608 15.588 12.64 18.096 ;
  LAYER M3 ;
        RECT 12.672 15.588 12.704 18.096 ;
  LAYER M3 ;
        RECT 12.736 15.588 12.768 18.096 ;
  LAYER M3 ;
        RECT 12.8 15.588 12.832 18.096 ;
  LAYER M3 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M3 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M3 ;
        RECT 13.024 15.588 13.056 18.096 ;
  LAYER M1 ;
        RECT 10.639 15.624 10.641 18.06 ;
  LAYER M1 ;
        RECT 10.719 15.624 10.721 18.06 ;
  LAYER M1 ;
        RECT 10.799 15.624 10.801 18.06 ;
  LAYER M1 ;
        RECT 10.879 15.624 10.881 18.06 ;
  LAYER M1 ;
        RECT 10.959 15.624 10.961 18.06 ;
  LAYER M1 ;
        RECT 11.039 15.624 11.041 18.06 ;
  LAYER M1 ;
        RECT 11.119 15.624 11.121 18.06 ;
  LAYER M1 ;
        RECT 11.199 15.624 11.201 18.06 ;
  LAYER M1 ;
        RECT 11.279 15.624 11.281 18.06 ;
  LAYER M1 ;
        RECT 11.359 15.624 11.361 18.06 ;
  LAYER M1 ;
        RECT 11.439 15.624 11.441 18.06 ;
  LAYER M1 ;
        RECT 11.519 15.624 11.521 18.06 ;
  LAYER M1 ;
        RECT 11.599 15.624 11.601 18.06 ;
  LAYER M1 ;
        RECT 11.679 15.624 11.681 18.06 ;
  LAYER M1 ;
        RECT 11.759 15.624 11.761 18.06 ;
  LAYER M1 ;
        RECT 11.839 15.624 11.841 18.06 ;
  LAYER M1 ;
        RECT 11.919 15.624 11.921 18.06 ;
  LAYER M1 ;
        RECT 11.999 15.624 12.001 18.06 ;
  LAYER M1 ;
        RECT 12.079 15.624 12.081 18.06 ;
  LAYER M1 ;
        RECT 12.159 15.624 12.161 18.06 ;
  LAYER M1 ;
        RECT 12.239 15.624 12.241 18.06 ;
  LAYER M1 ;
        RECT 12.319 15.624 12.321 18.06 ;
  LAYER M1 ;
        RECT 12.399 15.624 12.401 18.06 ;
  LAYER M1 ;
        RECT 12.479 15.624 12.481 18.06 ;
  LAYER M1 ;
        RECT 12.559 15.624 12.561 18.06 ;
  LAYER M1 ;
        RECT 12.639 15.624 12.641 18.06 ;
  LAYER M1 ;
        RECT 12.719 15.624 12.721 18.06 ;
  LAYER M1 ;
        RECT 12.799 15.624 12.801 18.06 ;
  LAYER M1 ;
        RECT 12.879 15.624 12.881 18.06 ;
  LAYER M1 ;
        RECT 12.959 15.624 12.961 18.06 ;
  LAYER M2 ;
        RECT 10.64 15.623 13.04 15.625 ;
  LAYER M2 ;
        RECT 10.64 15.707 13.04 15.709 ;
  LAYER M2 ;
        RECT 10.64 15.791 13.04 15.793 ;
  LAYER M2 ;
        RECT 10.64 15.875 13.04 15.877 ;
  LAYER M2 ;
        RECT 10.64 15.959 13.04 15.961 ;
  LAYER M2 ;
        RECT 10.64 16.043 13.04 16.045 ;
  LAYER M2 ;
        RECT 10.64 16.127 13.04 16.129 ;
  LAYER M2 ;
        RECT 10.64 16.211 13.04 16.213 ;
  LAYER M2 ;
        RECT 10.64 16.295 13.04 16.297 ;
  LAYER M2 ;
        RECT 10.64 16.379 13.04 16.381 ;
  LAYER M2 ;
        RECT 10.64 16.463 13.04 16.465 ;
  LAYER M2 ;
        RECT 10.64 16.547 13.04 16.549 ;
  LAYER M2 ;
        RECT 10.64 16.6305 13.04 16.6325 ;
  LAYER M2 ;
        RECT 10.64 16.715 13.04 16.717 ;
  LAYER M2 ;
        RECT 10.64 16.799 13.04 16.801 ;
  LAYER M2 ;
        RECT 10.64 16.883 13.04 16.885 ;
  LAYER M2 ;
        RECT 10.64 16.967 13.04 16.969 ;
  LAYER M2 ;
        RECT 10.64 17.051 13.04 17.053 ;
  LAYER M2 ;
        RECT 10.64 17.135 13.04 17.137 ;
  LAYER M2 ;
        RECT 10.64 17.219 13.04 17.221 ;
  LAYER M2 ;
        RECT 10.64 17.303 13.04 17.305 ;
  LAYER M2 ;
        RECT 10.64 17.387 13.04 17.389 ;
  LAYER M2 ;
        RECT 10.64 17.471 13.04 17.473 ;
  LAYER M2 ;
        RECT 10.64 17.555 13.04 17.557 ;
  LAYER M2 ;
        RECT 10.64 17.639 13.04 17.641 ;
  LAYER M2 ;
        RECT 10.64 17.723 13.04 17.725 ;
  LAYER M2 ;
        RECT 10.64 17.807 13.04 17.809 ;
  LAYER M2 ;
        RECT 10.64 17.891 13.04 17.893 ;
  LAYER M2 ;
        RECT 10.64 17.975 13.04 17.977 ;
  LAYER M1 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M1 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M1 ;
        RECT 14.272 0.888 14.304 3.396 ;
  LAYER M1 ;
        RECT 14.336 0.888 14.368 3.396 ;
  LAYER M1 ;
        RECT 14.4 0.888 14.432 3.396 ;
  LAYER M1 ;
        RECT 14.464 0.888 14.496 3.396 ;
  LAYER M1 ;
        RECT 14.528 0.888 14.56 3.396 ;
  LAYER M1 ;
        RECT 14.592 0.888 14.624 3.396 ;
  LAYER M1 ;
        RECT 14.656 0.888 14.688 3.396 ;
  LAYER M1 ;
        RECT 14.72 0.888 14.752 3.396 ;
  LAYER M1 ;
        RECT 14.784 0.888 14.816 3.396 ;
  LAYER M1 ;
        RECT 14.848 0.888 14.88 3.396 ;
  LAYER M1 ;
        RECT 14.912 0.888 14.944 3.396 ;
  LAYER M1 ;
        RECT 14.976 0.888 15.008 3.396 ;
  LAYER M1 ;
        RECT 15.04 0.888 15.072 3.396 ;
  LAYER M1 ;
        RECT 15.104 0.888 15.136 3.396 ;
  LAYER M1 ;
        RECT 15.168 0.888 15.2 3.396 ;
  LAYER M1 ;
        RECT 15.232 0.888 15.264 3.396 ;
  LAYER M1 ;
        RECT 15.296 0.888 15.328 3.396 ;
  LAYER M1 ;
        RECT 15.36 0.888 15.392 3.396 ;
  LAYER M1 ;
        RECT 15.424 0.888 15.456 3.396 ;
  LAYER M1 ;
        RECT 15.488 0.888 15.52 3.396 ;
  LAYER M1 ;
        RECT 15.552 0.888 15.584 3.396 ;
  LAYER M1 ;
        RECT 15.616 0.888 15.648 3.396 ;
  LAYER M1 ;
        RECT 15.68 0.888 15.712 3.396 ;
  LAYER M1 ;
        RECT 15.744 0.888 15.776 3.396 ;
  LAYER M1 ;
        RECT 15.808 0.888 15.84 3.396 ;
  LAYER M1 ;
        RECT 15.872 0.888 15.904 3.396 ;
  LAYER M1 ;
        RECT 15.936 0.888 15.968 3.396 ;
  LAYER M1 ;
        RECT 16 0.888 16.032 3.396 ;
  LAYER M1 ;
        RECT 16.064 0.888 16.096 3.396 ;
  LAYER M1 ;
        RECT 16.128 0.888 16.16 3.396 ;
  LAYER M1 ;
        RECT 16.192 0.888 16.224 3.396 ;
  LAYER M1 ;
        RECT 16.256 0.888 16.288 3.396 ;
  LAYER M1 ;
        RECT 16.32 0.888 16.352 3.396 ;
  LAYER M1 ;
        RECT 16.384 0.888 16.416 3.396 ;
  LAYER M1 ;
        RECT 16.448 0.888 16.48 3.396 ;
  LAYER M2 ;
        RECT 14.124 0.972 16.596 1.004 ;
  LAYER M2 ;
        RECT 14.124 1.036 16.596 1.068 ;
  LAYER M2 ;
        RECT 14.124 1.1 16.596 1.132 ;
  LAYER M2 ;
        RECT 14.124 1.164 16.596 1.196 ;
  LAYER M2 ;
        RECT 14.124 1.228 16.596 1.26 ;
  LAYER M2 ;
        RECT 14.124 1.292 16.596 1.324 ;
  LAYER M2 ;
        RECT 14.124 1.356 16.596 1.388 ;
  LAYER M2 ;
        RECT 14.124 1.42 16.596 1.452 ;
  LAYER M2 ;
        RECT 14.124 1.484 16.596 1.516 ;
  LAYER M2 ;
        RECT 14.124 1.548 16.596 1.58 ;
  LAYER M2 ;
        RECT 14.124 1.612 16.596 1.644 ;
  LAYER M2 ;
        RECT 14.124 1.676 16.596 1.708 ;
  LAYER M2 ;
        RECT 14.124 1.74 16.596 1.772 ;
  LAYER M2 ;
        RECT 14.124 1.804 16.596 1.836 ;
  LAYER M2 ;
        RECT 14.124 1.868 16.596 1.9 ;
  LAYER M2 ;
        RECT 14.124 1.932 16.596 1.964 ;
  LAYER M2 ;
        RECT 14.124 1.996 16.596 2.028 ;
  LAYER M2 ;
        RECT 14.124 2.06 16.596 2.092 ;
  LAYER M2 ;
        RECT 14.124 2.124 16.596 2.156 ;
  LAYER M2 ;
        RECT 14.124 2.188 16.596 2.22 ;
  LAYER M2 ;
        RECT 14.124 2.252 16.596 2.284 ;
  LAYER M2 ;
        RECT 14.124 2.316 16.596 2.348 ;
  LAYER M2 ;
        RECT 14.124 2.38 16.596 2.412 ;
  LAYER M2 ;
        RECT 14.124 2.444 16.596 2.476 ;
  LAYER M2 ;
        RECT 14.124 2.508 16.596 2.54 ;
  LAYER M2 ;
        RECT 14.124 2.572 16.596 2.604 ;
  LAYER M2 ;
        RECT 14.124 2.636 16.596 2.668 ;
  LAYER M2 ;
        RECT 14.124 2.7 16.596 2.732 ;
  LAYER M2 ;
        RECT 14.124 2.764 16.596 2.796 ;
  LAYER M2 ;
        RECT 14.124 2.828 16.596 2.86 ;
  LAYER M2 ;
        RECT 14.124 2.892 16.596 2.924 ;
  LAYER M2 ;
        RECT 14.124 2.956 16.596 2.988 ;
  LAYER M2 ;
        RECT 14.124 3.02 16.596 3.052 ;
  LAYER M2 ;
        RECT 14.124 3.084 16.596 3.116 ;
  LAYER M2 ;
        RECT 14.124 3.148 16.596 3.18 ;
  LAYER M2 ;
        RECT 14.124 3.212 16.596 3.244 ;
  LAYER M3 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M3 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M3 ;
        RECT 14.272 0.888 14.304 3.396 ;
  LAYER M3 ;
        RECT 14.336 0.888 14.368 3.396 ;
  LAYER M3 ;
        RECT 14.4 0.888 14.432 3.396 ;
  LAYER M3 ;
        RECT 14.464 0.888 14.496 3.396 ;
  LAYER M3 ;
        RECT 14.528 0.888 14.56 3.396 ;
  LAYER M3 ;
        RECT 14.592 0.888 14.624 3.396 ;
  LAYER M3 ;
        RECT 14.656 0.888 14.688 3.396 ;
  LAYER M3 ;
        RECT 14.72 0.888 14.752 3.396 ;
  LAYER M3 ;
        RECT 14.784 0.888 14.816 3.396 ;
  LAYER M3 ;
        RECT 14.848 0.888 14.88 3.396 ;
  LAYER M3 ;
        RECT 14.912 0.888 14.944 3.396 ;
  LAYER M3 ;
        RECT 14.976 0.888 15.008 3.396 ;
  LAYER M3 ;
        RECT 15.04 0.888 15.072 3.396 ;
  LAYER M3 ;
        RECT 15.104 0.888 15.136 3.396 ;
  LAYER M3 ;
        RECT 15.168 0.888 15.2 3.396 ;
  LAYER M3 ;
        RECT 15.232 0.888 15.264 3.396 ;
  LAYER M3 ;
        RECT 15.296 0.888 15.328 3.396 ;
  LAYER M3 ;
        RECT 15.36 0.888 15.392 3.396 ;
  LAYER M3 ;
        RECT 15.424 0.888 15.456 3.396 ;
  LAYER M3 ;
        RECT 15.488 0.888 15.52 3.396 ;
  LAYER M3 ;
        RECT 15.552 0.888 15.584 3.396 ;
  LAYER M3 ;
        RECT 15.616 0.888 15.648 3.396 ;
  LAYER M3 ;
        RECT 15.68 0.888 15.712 3.396 ;
  LAYER M3 ;
        RECT 15.744 0.888 15.776 3.396 ;
  LAYER M3 ;
        RECT 15.808 0.888 15.84 3.396 ;
  LAYER M3 ;
        RECT 15.872 0.888 15.904 3.396 ;
  LAYER M3 ;
        RECT 15.936 0.888 15.968 3.396 ;
  LAYER M3 ;
        RECT 16 0.888 16.032 3.396 ;
  LAYER M3 ;
        RECT 16.064 0.888 16.096 3.396 ;
  LAYER M3 ;
        RECT 16.128 0.888 16.16 3.396 ;
  LAYER M3 ;
        RECT 16.192 0.888 16.224 3.396 ;
  LAYER M3 ;
        RECT 16.256 0.888 16.288 3.396 ;
  LAYER M3 ;
        RECT 16.32 0.888 16.352 3.396 ;
  LAYER M3 ;
        RECT 16.384 0.888 16.416 3.396 ;
  LAYER M3 ;
        RECT 16.448 0.888 16.48 3.396 ;
  LAYER M3 ;
        RECT 16.544 0.888 16.576 3.396 ;
  LAYER M1 ;
        RECT 14.159 0.924 14.161 3.36 ;
  LAYER M1 ;
        RECT 14.239 0.924 14.241 3.36 ;
  LAYER M1 ;
        RECT 14.319 0.924 14.321 3.36 ;
  LAYER M1 ;
        RECT 14.399 0.924 14.401 3.36 ;
  LAYER M1 ;
        RECT 14.479 0.924 14.481 3.36 ;
  LAYER M1 ;
        RECT 14.559 0.924 14.561 3.36 ;
  LAYER M1 ;
        RECT 14.639 0.924 14.641 3.36 ;
  LAYER M1 ;
        RECT 14.719 0.924 14.721 3.36 ;
  LAYER M1 ;
        RECT 14.799 0.924 14.801 3.36 ;
  LAYER M1 ;
        RECT 14.879 0.924 14.881 3.36 ;
  LAYER M1 ;
        RECT 14.959 0.924 14.961 3.36 ;
  LAYER M1 ;
        RECT 15.039 0.924 15.041 3.36 ;
  LAYER M1 ;
        RECT 15.119 0.924 15.121 3.36 ;
  LAYER M1 ;
        RECT 15.199 0.924 15.201 3.36 ;
  LAYER M1 ;
        RECT 15.279 0.924 15.281 3.36 ;
  LAYER M1 ;
        RECT 15.359 0.924 15.361 3.36 ;
  LAYER M1 ;
        RECT 15.439 0.924 15.441 3.36 ;
  LAYER M1 ;
        RECT 15.519 0.924 15.521 3.36 ;
  LAYER M1 ;
        RECT 15.599 0.924 15.601 3.36 ;
  LAYER M1 ;
        RECT 15.679 0.924 15.681 3.36 ;
  LAYER M1 ;
        RECT 15.759 0.924 15.761 3.36 ;
  LAYER M1 ;
        RECT 15.839 0.924 15.841 3.36 ;
  LAYER M1 ;
        RECT 15.919 0.924 15.921 3.36 ;
  LAYER M1 ;
        RECT 15.999 0.924 16.001 3.36 ;
  LAYER M1 ;
        RECT 16.079 0.924 16.081 3.36 ;
  LAYER M1 ;
        RECT 16.159 0.924 16.161 3.36 ;
  LAYER M1 ;
        RECT 16.239 0.924 16.241 3.36 ;
  LAYER M1 ;
        RECT 16.319 0.924 16.321 3.36 ;
  LAYER M1 ;
        RECT 16.399 0.924 16.401 3.36 ;
  LAYER M1 ;
        RECT 16.479 0.924 16.481 3.36 ;
  LAYER M2 ;
        RECT 14.16 0.923 16.56 0.925 ;
  LAYER M2 ;
        RECT 14.16 1.007 16.56 1.009 ;
  LAYER M2 ;
        RECT 14.16 1.091 16.56 1.093 ;
  LAYER M2 ;
        RECT 14.16 1.175 16.56 1.177 ;
  LAYER M2 ;
        RECT 14.16 1.259 16.56 1.261 ;
  LAYER M2 ;
        RECT 14.16 1.343 16.56 1.345 ;
  LAYER M2 ;
        RECT 14.16 1.427 16.56 1.429 ;
  LAYER M2 ;
        RECT 14.16 1.511 16.56 1.513 ;
  LAYER M2 ;
        RECT 14.16 1.595 16.56 1.597 ;
  LAYER M2 ;
        RECT 14.16 1.679 16.56 1.681 ;
  LAYER M2 ;
        RECT 14.16 1.763 16.56 1.765 ;
  LAYER M2 ;
        RECT 14.16 1.847 16.56 1.849 ;
  LAYER M2 ;
        RECT 14.16 1.9305 16.56 1.9325 ;
  LAYER M2 ;
        RECT 14.16 2.015 16.56 2.017 ;
  LAYER M2 ;
        RECT 14.16 2.099 16.56 2.101 ;
  LAYER M2 ;
        RECT 14.16 2.183 16.56 2.185 ;
  LAYER M2 ;
        RECT 14.16 2.267 16.56 2.269 ;
  LAYER M2 ;
        RECT 14.16 2.351 16.56 2.353 ;
  LAYER M2 ;
        RECT 14.16 2.435 16.56 2.437 ;
  LAYER M2 ;
        RECT 14.16 2.519 16.56 2.521 ;
  LAYER M2 ;
        RECT 14.16 2.603 16.56 2.605 ;
  LAYER M2 ;
        RECT 14.16 2.687 16.56 2.689 ;
  LAYER M2 ;
        RECT 14.16 2.771 16.56 2.773 ;
  LAYER M2 ;
        RECT 14.16 2.855 16.56 2.857 ;
  LAYER M2 ;
        RECT 14.16 2.939 16.56 2.941 ;
  LAYER M2 ;
        RECT 14.16 3.023 16.56 3.025 ;
  LAYER M2 ;
        RECT 14.16 3.107 16.56 3.109 ;
  LAYER M2 ;
        RECT 14.16 3.191 16.56 3.193 ;
  LAYER M2 ;
        RECT 14.16 3.275 16.56 3.277 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M1 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M1 ;
        RECT 14.272 3.828 14.304 6.336 ;
  LAYER M1 ;
        RECT 14.336 3.828 14.368 6.336 ;
  LAYER M1 ;
        RECT 14.4 3.828 14.432 6.336 ;
  LAYER M1 ;
        RECT 14.464 3.828 14.496 6.336 ;
  LAYER M1 ;
        RECT 14.528 3.828 14.56 6.336 ;
  LAYER M1 ;
        RECT 14.592 3.828 14.624 6.336 ;
  LAYER M1 ;
        RECT 14.656 3.828 14.688 6.336 ;
  LAYER M1 ;
        RECT 14.72 3.828 14.752 6.336 ;
  LAYER M1 ;
        RECT 14.784 3.828 14.816 6.336 ;
  LAYER M1 ;
        RECT 14.848 3.828 14.88 6.336 ;
  LAYER M1 ;
        RECT 14.912 3.828 14.944 6.336 ;
  LAYER M1 ;
        RECT 14.976 3.828 15.008 6.336 ;
  LAYER M1 ;
        RECT 15.04 3.828 15.072 6.336 ;
  LAYER M1 ;
        RECT 15.104 3.828 15.136 6.336 ;
  LAYER M1 ;
        RECT 15.168 3.828 15.2 6.336 ;
  LAYER M1 ;
        RECT 15.232 3.828 15.264 6.336 ;
  LAYER M1 ;
        RECT 15.296 3.828 15.328 6.336 ;
  LAYER M1 ;
        RECT 15.36 3.828 15.392 6.336 ;
  LAYER M1 ;
        RECT 15.424 3.828 15.456 6.336 ;
  LAYER M1 ;
        RECT 15.488 3.828 15.52 6.336 ;
  LAYER M1 ;
        RECT 15.552 3.828 15.584 6.336 ;
  LAYER M1 ;
        RECT 15.616 3.828 15.648 6.336 ;
  LAYER M1 ;
        RECT 15.68 3.828 15.712 6.336 ;
  LAYER M1 ;
        RECT 15.744 3.828 15.776 6.336 ;
  LAYER M1 ;
        RECT 15.808 3.828 15.84 6.336 ;
  LAYER M1 ;
        RECT 15.872 3.828 15.904 6.336 ;
  LAYER M1 ;
        RECT 15.936 3.828 15.968 6.336 ;
  LAYER M1 ;
        RECT 16 3.828 16.032 6.336 ;
  LAYER M1 ;
        RECT 16.064 3.828 16.096 6.336 ;
  LAYER M1 ;
        RECT 16.128 3.828 16.16 6.336 ;
  LAYER M1 ;
        RECT 16.192 3.828 16.224 6.336 ;
  LAYER M1 ;
        RECT 16.256 3.828 16.288 6.336 ;
  LAYER M1 ;
        RECT 16.32 3.828 16.352 6.336 ;
  LAYER M1 ;
        RECT 16.384 3.828 16.416 6.336 ;
  LAYER M1 ;
        RECT 16.448 3.828 16.48 6.336 ;
  LAYER M2 ;
        RECT 14.124 3.912 16.596 3.944 ;
  LAYER M2 ;
        RECT 14.124 3.976 16.596 4.008 ;
  LAYER M2 ;
        RECT 14.124 4.04 16.596 4.072 ;
  LAYER M2 ;
        RECT 14.124 4.104 16.596 4.136 ;
  LAYER M2 ;
        RECT 14.124 4.168 16.596 4.2 ;
  LAYER M2 ;
        RECT 14.124 4.232 16.596 4.264 ;
  LAYER M2 ;
        RECT 14.124 4.296 16.596 4.328 ;
  LAYER M2 ;
        RECT 14.124 4.36 16.596 4.392 ;
  LAYER M2 ;
        RECT 14.124 4.424 16.596 4.456 ;
  LAYER M2 ;
        RECT 14.124 4.488 16.596 4.52 ;
  LAYER M2 ;
        RECT 14.124 4.552 16.596 4.584 ;
  LAYER M2 ;
        RECT 14.124 4.616 16.596 4.648 ;
  LAYER M2 ;
        RECT 14.124 4.68 16.596 4.712 ;
  LAYER M2 ;
        RECT 14.124 4.744 16.596 4.776 ;
  LAYER M2 ;
        RECT 14.124 4.808 16.596 4.84 ;
  LAYER M2 ;
        RECT 14.124 4.872 16.596 4.904 ;
  LAYER M2 ;
        RECT 14.124 4.936 16.596 4.968 ;
  LAYER M2 ;
        RECT 14.124 5 16.596 5.032 ;
  LAYER M2 ;
        RECT 14.124 5.064 16.596 5.096 ;
  LAYER M2 ;
        RECT 14.124 5.128 16.596 5.16 ;
  LAYER M2 ;
        RECT 14.124 5.192 16.596 5.224 ;
  LAYER M2 ;
        RECT 14.124 5.256 16.596 5.288 ;
  LAYER M2 ;
        RECT 14.124 5.32 16.596 5.352 ;
  LAYER M2 ;
        RECT 14.124 5.384 16.596 5.416 ;
  LAYER M2 ;
        RECT 14.124 5.448 16.596 5.48 ;
  LAYER M2 ;
        RECT 14.124 5.512 16.596 5.544 ;
  LAYER M2 ;
        RECT 14.124 5.576 16.596 5.608 ;
  LAYER M2 ;
        RECT 14.124 5.64 16.596 5.672 ;
  LAYER M2 ;
        RECT 14.124 5.704 16.596 5.736 ;
  LAYER M2 ;
        RECT 14.124 5.768 16.596 5.8 ;
  LAYER M2 ;
        RECT 14.124 5.832 16.596 5.864 ;
  LAYER M2 ;
        RECT 14.124 5.896 16.596 5.928 ;
  LAYER M2 ;
        RECT 14.124 5.96 16.596 5.992 ;
  LAYER M2 ;
        RECT 14.124 6.024 16.596 6.056 ;
  LAYER M2 ;
        RECT 14.124 6.088 16.596 6.12 ;
  LAYER M2 ;
        RECT 14.124 6.152 16.596 6.184 ;
  LAYER M3 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M3 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M3 ;
        RECT 14.272 3.828 14.304 6.336 ;
  LAYER M3 ;
        RECT 14.336 3.828 14.368 6.336 ;
  LAYER M3 ;
        RECT 14.4 3.828 14.432 6.336 ;
  LAYER M3 ;
        RECT 14.464 3.828 14.496 6.336 ;
  LAYER M3 ;
        RECT 14.528 3.828 14.56 6.336 ;
  LAYER M3 ;
        RECT 14.592 3.828 14.624 6.336 ;
  LAYER M3 ;
        RECT 14.656 3.828 14.688 6.336 ;
  LAYER M3 ;
        RECT 14.72 3.828 14.752 6.336 ;
  LAYER M3 ;
        RECT 14.784 3.828 14.816 6.336 ;
  LAYER M3 ;
        RECT 14.848 3.828 14.88 6.336 ;
  LAYER M3 ;
        RECT 14.912 3.828 14.944 6.336 ;
  LAYER M3 ;
        RECT 14.976 3.828 15.008 6.336 ;
  LAYER M3 ;
        RECT 15.04 3.828 15.072 6.336 ;
  LAYER M3 ;
        RECT 15.104 3.828 15.136 6.336 ;
  LAYER M3 ;
        RECT 15.168 3.828 15.2 6.336 ;
  LAYER M3 ;
        RECT 15.232 3.828 15.264 6.336 ;
  LAYER M3 ;
        RECT 15.296 3.828 15.328 6.336 ;
  LAYER M3 ;
        RECT 15.36 3.828 15.392 6.336 ;
  LAYER M3 ;
        RECT 15.424 3.828 15.456 6.336 ;
  LAYER M3 ;
        RECT 15.488 3.828 15.52 6.336 ;
  LAYER M3 ;
        RECT 15.552 3.828 15.584 6.336 ;
  LAYER M3 ;
        RECT 15.616 3.828 15.648 6.336 ;
  LAYER M3 ;
        RECT 15.68 3.828 15.712 6.336 ;
  LAYER M3 ;
        RECT 15.744 3.828 15.776 6.336 ;
  LAYER M3 ;
        RECT 15.808 3.828 15.84 6.336 ;
  LAYER M3 ;
        RECT 15.872 3.828 15.904 6.336 ;
  LAYER M3 ;
        RECT 15.936 3.828 15.968 6.336 ;
  LAYER M3 ;
        RECT 16 3.828 16.032 6.336 ;
  LAYER M3 ;
        RECT 16.064 3.828 16.096 6.336 ;
  LAYER M3 ;
        RECT 16.128 3.828 16.16 6.336 ;
  LAYER M3 ;
        RECT 16.192 3.828 16.224 6.336 ;
  LAYER M3 ;
        RECT 16.256 3.828 16.288 6.336 ;
  LAYER M3 ;
        RECT 16.32 3.828 16.352 6.336 ;
  LAYER M3 ;
        RECT 16.384 3.828 16.416 6.336 ;
  LAYER M3 ;
        RECT 16.448 3.828 16.48 6.336 ;
  LAYER M3 ;
        RECT 16.544 3.828 16.576 6.336 ;
  LAYER M1 ;
        RECT 14.159 3.864 14.161 6.3 ;
  LAYER M1 ;
        RECT 14.239 3.864 14.241 6.3 ;
  LAYER M1 ;
        RECT 14.319 3.864 14.321 6.3 ;
  LAYER M1 ;
        RECT 14.399 3.864 14.401 6.3 ;
  LAYER M1 ;
        RECT 14.479 3.864 14.481 6.3 ;
  LAYER M1 ;
        RECT 14.559 3.864 14.561 6.3 ;
  LAYER M1 ;
        RECT 14.639 3.864 14.641 6.3 ;
  LAYER M1 ;
        RECT 14.719 3.864 14.721 6.3 ;
  LAYER M1 ;
        RECT 14.799 3.864 14.801 6.3 ;
  LAYER M1 ;
        RECT 14.879 3.864 14.881 6.3 ;
  LAYER M1 ;
        RECT 14.959 3.864 14.961 6.3 ;
  LAYER M1 ;
        RECT 15.039 3.864 15.041 6.3 ;
  LAYER M1 ;
        RECT 15.119 3.864 15.121 6.3 ;
  LAYER M1 ;
        RECT 15.199 3.864 15.201 6.3 ;
  LAYER M1 ;
        RECT 15.279 3.864 15.281 6.3 ;
  LAYER M1 ;
        RECT 15.359 3.864 15.361 6.3 ;
  LAYER M1 ;
        RECT 15.439 3.864 15.441 6.3 ;
  LAYER M1 ;
        RECT 15.519 3.864 15.521 6.3 ;
  LAYER M1 ;
        RECT 15.599 3.864 15.601 6.3 ;
  LAYER M1 ;
        RECT 15.679 3.864 15.681 6.3 ;
  LAYER M1 ;
        RECT 15.759 3.864 15.761 6.3 ;
  LAYER M1 ;
        RECT 15.839 3.864 15.841 6.3 ;
  LAYER M1 ;
        RECT 15.919 3.864 15.921 6.3 ;
  LAYER M1 ;
        RECT 15.999 3.864 16.001 6.3 ;
  LAYER M1 ;
        RECT 16.079 3.864 16.081 6.3 ;
  LAYER M1 ;
        RECT 16.159 3.864 16.161 6.3 ;
  LAYER M1 ;
        RECT 16.239 3.864 16.241 6.3 ;
  LAYER M1 ;
        RECT 16.319 3.864 16.321 6.3 ;
  LAYER M1 ;
        RECT 16.399 3.864 16.401 6.3 ;
  LAYER M1 ;
        RECT 16.479 3.864 16.481 6.3 ;
  LAYER M2 ;
        RECT 14.16 3.863 16.56 3.865 ;
  LAYER M2 ;
        RECT 14.16 3.947 16.56 3.949 ;
  LAYER M2 ;
        RECT 14.16 4.031 16.56 4.033 ;
  LAYER M2 ;
        RECT 14.16 4.115 16.56 4.117 ;
  LAYER M2 ;
        RECT 14.16 4.199 16.56 4.201 ;
  LAYER M2 ;
        RECT 14.16 4.283 16.56 4.285 ;
  LAYER M2 ;
        RECT 14.16 4.367 16.56 4.369 ;
  LAYER M2 ;
        RECT 14.16 4.451 16.56 4.453 ;
  LAYER M2 ;
        RECT 14.16 4.535 16.56 4.537 ;
  LAYER M2 ;
        RECT 14.16 4.619 16.56 4.621 ;
  LAYER M2 ;
        RECT 14.16 4.703 16.56 4.705 ;
  LAYER M2 ;
        RECT 14.16 4.787 16.56 4.789 ;
  LAYER M2 ;
        RECT 14.16 4.8705 16.56 4.8725 ;
  LAYER M2 ;
        RECT 14.16 4.955 16.56 4.957 ;
  LAYER M2 ;
        RECT 14.16 5.039 16.56 5.041 ;
  LAYER M2 ;
        RECT 14.16 5.123 16.56 5.125 ;
  LAYER M2 ;
        RECT 14.16 5.207 16.56 5.209 ;
  LAYER M2 ;
        RECT 14.16 5.291 16.56 5.293 ;
  LAYER M2 ;
        RECT 14.16 5.375 16.56 5.377 ;
  LAYER M2 ;
        RECT 14.16 5.459 16.56 5.461 ;
  LAYER M2 ;
        RECT 14.16 5.543 16.56 5.545 ;
  LAYER M2 ;
        RECT 14.16 5.627 16.56 5.629 ;
  LAYER M2 ;
        RECT 14.16 5.711 16.56 5.713 ;
  LAYER M2 ;
        RECT 14.16 5.795 16.56 5.797 ;
  LAYER M2 ;
        RECT 14.16 5.879 16.56 5.881 ;
  LAYER M2 ;
        RECT 14.16 5.963 16.56 5.965 ;
  LAYER M2 ;
        RECT 14.16 6.047 16.56 6.049 ;
  LAYER M2 ;
        RECT 14.16 6.131 16.56 6.133 ;
  LAYER M2 ;
        RECT 14.16 6.215 16.56 6.217 ;
  LAYER M1 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M1 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M1 ;
        RECT 14.272 6.768 14.304 9.276 ;
  LAYER M1 ;
        RECT 14.336 6.768 14.368 9.276 ;
  LAYER M1 ;
        RECT 14.4 6.768 14.432 9.276 ;
  LAYER M1 ;
        RECT 14.464 6.768 14.496 9.276 ;
  LAYER M1 ;
        RECT 14.528 6.768 14.56 9.276 ;
  LAYER M1 ;
        RECT 14.592 6.768 14.624 9.276 ;
  LAYER M1 ;
        RECT 14.656 6.768 14.688 9.276 ;
  LAYER M1 ;
        RECT 14.72 6.768 14.752 9.276 ;
  LAYER M1 ;
        RECT 14.784 6.768 14.816 9.276 ;
  LAYER M1 ;
        RECT 14.848 6.768 14.88 9.276 ;
  LAYER M1 ;
        RECT 14.912 6.768 14.944 9.276 ;
  LAYER M1 ;
        RECT 14.976 6.768 15.008 9.276 ;
  LAYER M1 ;
        RECT 15.04 6.768 15.072 9.276 ;
  LAYER M1 ;
        RECT 15.104 6.768 15.136 9.276 ;
  LAYER M1 ;
        RECT 15.168 6.768 15.2 9.276 ;
  LAYER M1 ;
        RECT 15.232 6.768 15.264 9.276 ;
  LAYER M1 ;
        RECT 15.296 6.768 15.328 9.276 ;
  LAYER M1 ;
        RECT 15.36 6.768 15.392 9.276 ;
  LAYER M1 ;
        RECT 15.424 6.768 15.456 9.276 ;
  LAYER M1 ;
        RECT 15.488 6.768 15.52 9.276 ;
  LAYER M1 ;
        RECT 15.552 6.768 15.584 9.276 ;
  LAYER M1 ;
        RECT 15.616 6.768 15.648 9.276 ;
  LAYER M1 ;
        RECT 15.68 6.768 15.712 9.276 ;
  LAYER M1 ;
        RECT 15.744 6.768 15.776 9.276 ;
  LAYER M1 ;
        RECT 15.808 6.768 15.84 9.276 ;
  LAYER M1 ;
        RECT 15.872 6.768 15.904 9.276 ;
  LAYER M1 ;
        RECT 15.936 6.768 15.968 9.276 ;
  LAYER M1 ;
        RECT 16 6.768 16.032 9.276 ;
  LAYER M1 ;
        RECT 16.064 6.768 16.096 9.276 ;
  LAYER M1 ;
        RECT 16.128 6.768 16.16 9.276 ;
  LAYER M1 ;
        RECT 16.192 6.768 16.224 9.276 ;
  LAYER M1 ;
        RECT 16.256 6.768 16.288 9.276 ;
  LAYER M1 ;
        RECT 16.32 6.768 16.352 9.276 ;
  LAYER M1 ;
        RECT 16.384 6.768 16.416 9.276 ;
  LAYER M1 ;
        RECT 16.448 6.768 16.48 9.276 ;
  LAYER M2 ;
        RECT 14.124 6.852 16.596 6.884 ;
  LAYER M2 ;
        RECT 14.124 6.916 16.596 6.948 ;
  LAYER M2 ;
        RECT 14.124 6.98 16.596 7.012 ;
  LAYER M2 ;
        RECT 14.124 7.044 16.596 7.076 ;
  LAYER M2 ;
        RECT 14.124 7.108 16.596 7.14 ;
  LAYER M2 ;
        RECT 14.124 7.172 16.596 7.204 ;
  LAYER M2 ;
        RECT 14.124 7.236 16.596 7.268 ;
  LAYER M2 ;
        RECT 14.124 7.3 16.596 7.332 ;
  LAYER M2 ;
        RECT 14.124 7.364 16.596 7.396 ;
  LAYER M2 ;
        RECT 14.124 7.428 16.596 7.46 ;
  LAYER M2 ;
        RECT 14.124 7.492 16.596 7.524 ;
  LAYER M2 ;
        RECT 14.124 7.556 16.596 7.588 ;
  LAYER M2 ;
        RECT 14.124 7.62 16.596 7.652 ;
  LAYER M2 ;
        RECT 14.124 7.684 16.596 7.716 ;
  LAYER M2 ;
        RECT 14.124 7.748 16.596 7.78 ;
  LAYER M2 ;
        RECT 14.124 7.812 16.596 7.844 ;
  LAYER M2 ;
        RECT 14.124 7.876 16.596 7.908 ;
  LAYER M2 ;
        RECT 14.124 7.94 16.596 7.972 ;
  LAYER M2 ;
        RECT 14.124 8.004 16.596 8.036 ;
  LAYER M2 ;
        RECT 14.124 8.068 16.596 8.1 ;
  LAYER M2 ;
        RECT 14.124 8.132 16.596 8.164 ;
  LAYER M2 ;
        RECT 14.124 8.196 16.596 8.228 ;
  LAYER M2 ;
        RECT 14.124 8.26 16.596 8.292 ;
  LAYER M2 ;
        RECT 14.124 8.324 16.596 8.356 ;
  LAYER M2 ;
        RECT 14.124 8.388 16.596 8.42 ;
  LAYER M2 ;
        RECT 14.124 8.452 16.596 8.484 ;
  LAYER M2 ;
        RECT 14.124 8.516 16.596 8.548 ;
  LAYER M2 ;
        RECT 14.124 8.58 16.596 8.612 ;
  LAYER M2 ;
        RECT 14.124 8.644 16.596 8.676 ;
  LAYER M2 ;
        RECT 14.124 8.708 16.596 8.74 ;
  LAYER M2 ;
        RECT 14.124 8.772 16.596 8.804 ;
  LAYER M2 ;
        RECT 14.124 8.836 16.596 8.868 ;
  LAYER M2 ;
        RECT 14.124 8.9 16.596 8.932 ;
  LAYER M2 ;
        RECT 14.124 8.964 16.596 8.996 ;
  LAYER M2 ;
        RECT 14.124 9.028 16.596 9.06 ;
  LAYER M2 ;
        RECT 14.124 9.092 16.596 9.124 ;
  LAYER M3 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M3 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M3 ;
        RECT 14.272 6.768 14.304 9.276 ;
  LAYER M3 ;
        RECT 14.336 6.768 14.368 9.276 ;
  LAYER M3 ;
        RECT 14.4 6.768 14.432 9.276 ;
  LAYER M3 ;
        RECT 14.464 6.768 14.496 9.276 ;
  LAYER M3 ;
        RECT 14.528 6.768 14.56 9.276 ;
  LAYER M3 ;
        RECT 14.592 6.768 14.624 9.276 ;
  LAYER M3 ;
        RECT 14.656 6.768 14.688 9.276 ;
  LAYER M3 ;
        RECT 14.72 6.768 14.752 9.276 ;
  LAYER M3 ;
        RECT 14.784 6.768 14.816 9.276 ;
  LAYER M3 ;
        RECT 14.848 6.768 14.88 9.276 ;
  LAYER M3 ;
        RECT 14.912 6.768 14.944 9.276 ;
  LAYER M3 ;
        RECT 14.976 6.768 15.008 9.276 ;
  LAYER M3 ;
        RECT 15.04 6.768 15.072 9.276 ;
  LAYER M3 ;
        RECT 15.104 6.768 15.136 9.276 ;
  LAYER M3 ;
        RECT 15.168 6.768 15.2 9.276 ;
  LAYER M3 ;
        RECT 15.232 6.768 15.264 9.276 ;
  LAYER M3 ;
        RECT 15.296 6.768 15.328 9.276 ;
  LAYER M3 ;
        RECT 15.36 6.768 15.392 9.276 ;
  LAYER M3 ;
        RECT 15.424 6.768 15.456 9.276 ;
  LAYER M3 ;
        RECT 15.488 6.768 15.52 9.276 ;
  LAYER M3 ;
        RECT 15.552 6.768 15.584 9.276 ;
  LAYER M3 ;
        RECT 15.616 6.768 15.648 9.276 ;
  LAYER M3 ;
        RECT 15.68 6.768 15.712 9.276 ;
  LAYER M3 ;
        RECT 15.744 6.768 15.776 9.276 ;
  LAYER M3 ;
        RECT 15.808 6.768 15.84 9.276 ;
  LAYER M3 ;
        RECT 15.872 6.768 15.904 9.276 ;
  LAYER M3 ;
        RECT 15.936 6.768 15.968 9.276 ;
  LAYER M3 ;
        RECT 16 6.768 16.032 9.276 ;
  LAYER M3 ;
        RECT 16.064 6.768 16.096 9.276 ;
  LAYER M3 ;
        RECT 16.128 6.768 16.16 9.276 ;
  LAYER M3 ;
        RECT 16.192 6.768 16.224 9.276 ;
  LAYER M3 ;
        RECT 16.256 6.768 16.288 9.276 ;
  LAYER M3 ;
        RECT 16.32 6.768 16.352 9.276 ;
  LAYER M3 ;
        RECT 16.384 6.768 16.416 9.276 ;
  LAYER M3 ;
        RECT 16.448 6.768 16.48 9.276 ;
  LAYER M3 ;
        RECT 16.544 6.768 16.576 9.276 ;
  LAYER M1 ;
        RECT 14.159 6.804 14.161 9.24 ;
  LAYER M1 ;
        RECT 14.239 6.804 14.241 9.24 ;
  LAYER M1 ;
        RECT 14.319 6.804 14.321 9.24 ;
  LAYER M1 ;
        RECT 14.399 6.804 14.401 9.24 ;
  LAYER M1 ;
        RECT 14.479 6.804 14.481 9.24 ;
  LAYER M1 ;
        RECT 14.559 6.804 14.561 9.24 ;
  LAYER M1 ;
        RECT 14.639 6.804 14.641 9.24 ;
  LAYER M1 ;
        RECT 14.719 6.804 14.721 9.24 ;
  LAYER M1 ;
        RECT 14.799 6.804 14.801 9.24 ;
  LAYER M1 ;
        RECT 14.879 6.804 14.881 9.24 ;
  LAYER M1 ;
        RECT 14.959 6.804 14.961 9.24 ;
  LAYER M1 ;
        RECT 15.039 6.804 15.041 9.24 ;
  LAYER M1 ;
        RECT 15.119 6.804 15.121 9.24 ;
  LAYER M1 ;
        RECT 15.199 6.804 15.201 9.24 ;
  LAYER M1 ;
        RECT 15.279 6.804 15.281 9.24 ;
  LAYER M1 ;
        RECT 15.359 6.804 15.361 9.24 ;
  LAYER M1 ;
        RECT 15.439 6.804 15.441 9.24 ;
  LAYER M1 ;
        RECT 15.519 6.804 15.521 9.24 ;
  LAYER M1 ;
        RECT 15.599 6.804 15.601 9.24 ;
  LAYER M1 ;
        RECT 15.679 6.804 15.681 9.24 ;
  LAYER M1 ;
        RECT 15.759 6.804 15.761 9.24 ;
  LAYER M1 ;
        RECT 15.839 6.804 15.841 9.24 ;
  LAYER M1 ;
        RECT 15.919 6.804 15.921 9.24 ;
  LAYER M1 ;
        RECT 15.999 6.804 16.001 9.24 ;
  LAYER M1 ;
        RECT 16.079 6.804 16.081 9.24 ;
  LAYER M1 ;
        RECT 16.159 6.804 16.161 9.24 ;
  LAYER M1 ;
        RECT 16.239 6.804 16.241 9.24 ;
  LAYER M1 ;
        RECT 16.319 6.804 16.321 9.24 ;
  LAYER M1 ;
        RECT 16.399 6.804 16.401 9.24 ;
  LAYER M1 ;
        RECT 16.479 6.804 16.481 9.24 ;
  LAYER M2 ;
        RECT 14.16 6.803 16.56 6.805 ;
  LAYER M2 ;
        RECT 14.16 6.887 16.56 6.889 ;
  LAYER M2 ;
        RECT 14.16 6.971 16.56 6.973 ;
  LAYER M2 ;
        RECT 14.16 7.055 16.56 7.057 ;
  LAYER M2 ;
        RECT 14.16 7.139 16.56 7.141 ;
  LAYER M2 ;
        RECT 14.16 7.223 16.56 7.225 ;
  LAYER M2 ;
        RECT 14.16 7.307 16.56 7.309 ;
  LAYER M2 ;
        RECT 14.16 7.391 16.56 7.393 ;
  LAYER M2 ;
        RECT 14.16 7.475 16.56 7.477 ;
  LAYER M2 ;
        RECT 14.16 7.559 16.56 7.561 ;
  LAYER M2 ;
        RECT 14.16 7.643 16.56 7.645 ;
  LAYER M2 ;
        RECT 14.16 7.727 16.56 7.729 ;
  LAYER M2 ;
        RECT 14.16 7.8105 16.56 7.8125 ;
  LAYER M2 ;
        RECT 14.16 7.895 16.56 7.897 ;
  LAYER M2 ;
        RECT 14.16 7.979 16.56 7.981 ;
  LAYER M2 ;
        RECT 14.16 8.063 16.56 8.065 ;
  LAYER M2 ;
        RECT 14.16 8.147 16.56 8.149 ;
  LAYER M2 ;
        RECT 14.16 8.231 16.56 8.233 ;
  LAYER M2 ;
        RECT 14.16 8.315 16.56 8.317 ;
  LAYER M2 ;
        RECT 14.16 8.399 16.56 8.401 ;
  LAYER M2 ;
        RECT 14.16 8.483 16.56 8.485 ;
  LAYER M2 ;
        RECT 14.16 8.567 16.56 8.569 ;
  LAYER M2 ;
        RECT 14.16 8.651 16.56 8.653 ;
  LAYER M2 ;
        RECT 14.16 8.735 16.56 8.737 ;
  LAYER M2 ;
        RECT 14.16 8.819 16.56 8.821 ;
  LAYER M2 ;
        RECT 14.16 8.903 16.56 8.905 ;
  LAYER M2 ;
        RECT 14.16 8.987 16.56 8.989 ;
  LAYER M2 ;
        RECT 14.16 9.071 16.56 9.073 ;
  LAYER M2 ;
        RECT 14.16 9.155 16.56 9.157 ;
  LAYER M1 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M1 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M1 ;
        RECT 14.272 9.708 14.304 12.216 ;
  LAYER M1 ;
        RECT 14.336 9.708 14.368 12.216 ;
  LAYER M1 ;
        RECT 14.4 9.708 14.432 12.216 ;
  LAYER M1 ;
        RECT 14.464 9.708 14.496 12.216 ;
  LAYER M1 ;
        RECT 14.528 9.708 14.56 12.216 ;
  LAYER M1 ;
        RECT 14.592 9.708 14.624 12.216 ;
  LAYER M1 ;
        RECT 14.656 9.708 14.688 12.216 ;
  LAYER M1 ;
        RECT 14.72 9.708 14.752 12.216 ;
  LAYER M1 ;
        RECT 14.784 9.708 14.816 12.216 ;
  LAYER M1 ;
        RECT 14.848 9.708 14.88 12.216 ;
  LAYER M1 ;
        RECT 14.912 9.708 14.944 12.216 ;
  LAYER M1 ;
        RECT 14.976 9.708 15.008 12.216 ;
  LAYER M1 ;
        RECT 15.04 9.708 15.072 12.216 ;
  LAYER M1 ;
        RECT 15.104 9.708 15.136 12.216 ;
  LAYER M1 ;
        RECT 15.168 9.708 15.2 12.216 ;
  LAYER M1 ;
        RECT 15.232 9.708 15.264 12.216 ;
  LAYER M1 ;
        RECT 15.296 9.708 15.328 12.216 ;
  LAYER M1 ;
        RECT 15.36 9.708 15.392 12.216 ;
  LAYER M1 ;
        RECT 15.424 9.708 15.456 12.216 ;
  LAYER M1 ;
        RECT 15.488 9.708 15.52 12.216 ;
  LAYER M1 ;
        RECT 15.552 9.708 15.584 12.216 ;
  LAYER M1 ;
        RECT 15.616 9.708 15.648 12.216 ;
  LAYER M1 ;
        RECT 15.68 9.708 15.712 12.216 ;
  LAYER M1 ;
        RECT 15.744 9.708 15.776 12.216 ;
  LAYER M1 ;
        RECT 15.808 9.708 15.84 12.216 ;
  LAYER M1 ;
        RECT 15.872 9.708 15.904 12.216 ;
  LAYER M1 ;
        RECT 15.936 9.708 15.968 12.216 ;
  LAYER M1 ;
        RECT 16 9.708 16.032 12.216 ;
  LAYER M1 ;
        RECT 16.064 9.708 16.096 12.216 ;
  LAYER M1 ;
        RECT 16.128 9.708 16.16 12.216 ;
  LAYER M1 ;
        RECT 16.192 9.708 16.224 12.216 ;
  LAYER M1 ;
        RECT 16.256 9.708 16.288 12.216 ;
  LAYER M1 ;
        RECT 16.32 9.708 16.352 12.216 ;
  LAYER M1 ;
        RECT 16.384 9.708 16.416 12.216 ;
  LAYER M1 ;
        RECT 16.448 9.708 16.48 12.216 ;
  LAYER M2 ;
        RECT 14.124 9.792 16.596 9.824 ;
  LAYER M2 ;
        RECT 14.124 9.856 16.596 9.888 ;
  LAYER M2 ;
        RECT 14.124 9.92 16.596 9.952 ;
  LAYER M2 ;
        RECT 14.124 9.984 16.596 10.016 ;
  LAYER M2 ;
        RECT 14.124 10.048 16.596 10.08 ;
  LAYER M2 ;
        RECT 14.124 10.112 16.596 10.144 ;
  LAYER M2 ;
        RECT 14.124 10.176 16.596 10.208 ;
  LAYER M2 ;
        RECT 14.124 10.24 16.596 10.272 ;
  LAYER M2 ;
        RECT 14.124 10.304 16.596 10.336 ;
  LAYER M2 ;
        RECT 14.124 10.368 16.596 10.4 ;
  LAYER M2 ;
        RECT 14.124 10.432 16.596 10.464 ;
  LAYER M2 ;
        RECT 14.124 10.496 16.596 10.528 ;
  LAYER M2 ;
        RECT 14.124 10.56 16.596 10.592 ;
  LAYER M2 ;
        RECT 14.124 10.624 16.596 10.656 ;
  LAYER M2 ;
        RECT 14.124 10.688 16.596 10.72 ;
  LAYER M2 ;
        RECT 14.124 10.752 16.596 10.784 ;
  LAYER M2 ;
        RECT 14.124 10.816 16.596 10.848 ;
  LAYER M2 ;
        RECT 14.124 10.88 16.596 10.912 ;
  LAYER M2 ;
        RECT 14.124 10.944 16.596 10.976 ;
  LAYER M2 ;
        RECT 14.124 11.008 16.596 11.04 ;
  LAYER M2 ;
        RECT 14.124 11.072 16.596 11.104 ;
  LAYER M2 ;
        RECT 14.124 11.136 16.596 11.168 ;
  LAYER M2 ;
        RECT 14.124 11.2 16.596 11.232 ;
  LAYER M2 ;
        RECT 14.124 11.264 16.596 11.296 ;
  LAYER M2 ;
        RECT 14.124 11.328 16.596 11.36 ;
  LAYER M2 ;
        RECT 14.124 11.392 16.596 11.424 ;
  LAYER M2 ;
        RECT 14.124 11.456 16.596 11.488 ;
  LAYER M2 ;
        RECT 14.124 11.52 16.596 11.552 ;
  LAYER M2 ;
        RECT 14.124 11.584 16.596 11.616 ;
  LAYER M2 ;
        RECT 14.124 11.648 16.596 11.68 ;
  LAYER M2 ;
        RECT 14.124 11.712 16.596 11.744 ;
  LAYER M2 ;
        RECT 14.124 11.776 16.596 11.808 ;
  LAYER M2 ;
        RECT 14.124 11.84 16.596 11.872 ;
  LAYER M2 ;
        RECT 14.124 11.904 16.596 11.936 ;
  LAYER M2 ;
        RECT 14.124 11.968 16.596 12 ;
  LAYER M2 ;
        RECT 14.124 12.032 16.596 12.064 ;
  LAYER M3 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M3 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M3 ;
        RECT 14.272 9.708 14.304 12.216 ;
  LAYER M3 ;
        RECT 14.336 9.708 14.368 12.216 ;
  LAYER M3 ;
        RECT 14.4 9.708 14.432 12.216 ;
  LAYER M3 ;
        RECT 14.464 9.708 14.496 12.216 ;
  LAYER M3 ;
        RECT 14.528 9.708 14.56 12.216 ;
  LAYER M3 ;
        RECT 14.592 9.708 14.624 12.216 ;
  LAYER M3 ;
        RECT 14.656 9.708 14.688 12.216 ;
  LAYER M3 ;
        RECT 14.72 9.708 14.752 12.216 ;
  LAYER M3 ;
        RECT 14.784 9.708 14.816 12.216 ;
  LAYER M3 ;
        RECT 14.848 9.708 14.88 12.216 ;
  LAYER M3 ;
        RECT 14.912 9.708 14.944 12.216 ;
  LAYER M3 ;
        RECT 14.976 9.708 15.008 12.216 ;
  LAYER M3 ;
        RECT 15.04 9.708 15.072 12.216 ;
  LAYER M3 ;
        RECT 15.104 9.708 15.136 12.216 ;
  LAYER M3 ;
        RECT 15.168 9.708 15.2 12.216 ;
  LAYER M3 ;
        RECT 15.232 9.708 15.264 12.216 ;
  LAYER M3 ;
        RECT 15.296 9.708 15.328 12.216 ;
  LAYER M3 ;
        RECT 15.36 9.708 15.392 12.216 ;
  LAYER M3 ;
        RECT 15.424 9.708 15.456 12.216 ;
  LAYER M3 ;
        RECT 15.488 9.708 15.52 12.216 ;
  LAYER M3 ;
        RECT 15.552 9.708 15.584 12.216 ;
  LAYER M3 ;
        RECT 15.616 9.708 15.648 12.216 ;
  LAYER M3 ;
        RECT 15.68 9.708 15.712 12.216 ;
  LAYER M3 ;
        RECT 15.744 9.708 15.776 12.216 ;
  LAYER M3 ;
        RECT 15.808 9.708 15.84 12.216 ;
  LAYER M3 ;
        RECT 15.872 9.708 15.904 12.216 ;
  LAYER M3 ;
        RECT 15.936 9.708 15.968 12.216 ;
  LAYER M3 ;
        RECT 16 9.708 16.032 12.216 ;
  LAYER M3 ;
        RECT 16.064 9.708 16.096 12.216 ;
  LAYER M3 ;
        RECT 16.128 9.708 16.16 12.216 ;
  LAYER M3 ;
        RECT 16.192 9.708 16.224 12.216 ;
  LAYER M3 ;
        RECT 16.256 9.708 16.288 12.216 ;
  LAYER M3 ;
        RECT 16.32 9.708 16.352 12.216 ;
  LAYER M3 ;
        RECT 16.384 9.708 16.416 12.216 ;
  LAYER M3 ;
        RECT 16.448 9.708 16.48 12.216 ;
  LAYER M3 ;
        RECT 16.544 9.708 16.576 12.216 ;
  LAYER M1 ;
        RECT 14.159 9.744 14.161 12.18 ;
  LAYER M1 ;
        RECT 14.239 9.744 14.241 12.18 ;
  LAYER M1 ;
        RECT 14.319 9.744 14.321 12.18 ;
  LAYER M1 ;
        RECT 14.399 9.744 14.401 12.18 ;
  LAYER M1 ;
        RECT 14.479 9.744 14.481 12.18 ;
  LAYER M1 ;
        RECT 14.559 9.744 14.561 12.18 ;
  LAYER M1 ;
        RECT 14.639 9.744 14.641 12.18 ;
  LAYER M1 ;
        RECT 14.719 9.744 14.721 12.18 ;
  LAYER M1 ;
        RECT 14.799 9.744 14.801 12.18 ;
  LAYER M1 ;
        RECT 14.879 9.744 14.881 12.18 ;
  LAYER M1 ;
        RECT 14.959 9.744 14.961 12.18 ;
  LAYER M1 ;
        RECT 15.039 9.744 15.041 12.18 ;
  LAYER M1 ;
        RECT 15.119 9.744 15.121 12.18 ;
  LAYER M1 ;
        RECT 15.199 9.744 15.201 12.18 ;
  LAYER M1 ;
        RECT 15.279 9.744 15.281 12.18 ;
  LAYER M1 ;
        RECT 15.359 9.744 15.361 12.18 ;
  LAYER M1 ;
        RECT 15.439 9.744 15.441 12.18 ;
  LAYER M1 ;
        RECT 15.519 9.744 15.521 12.18 ;
  LAYER M1 ;
        RECT 15.599 9.744 15.601 12.18 ;
  LAYER M1 ;
        RECT 15.679 9.744 15.681 12.18 ;
  LAYER M1 ;
        RECT 15.759 9.744 15.761 12.18 ;
  LAYER M1 ;
        RECT 15.839 9.744 15.841 12.18 ;
  LAYER M1 ;
        RECT 15.919 9.744 15.921 12.18 ;
  LAYER M1 ;
        RECT 15.999 9.744 16.001 12.18 ;
  LAYER M1 ;
        RECT 16.079 9.744 16.081 12.18 ;
  LAYER M1 ;
        RECT 16.159 9.744 16.161 12.18 ;
  LAYER M1 ;
        RECT 16.239 9.744 16.241 12.18 ;
  LAYER M1 ;
        RECT 16.319 9.744 16.321 12.18 ;
  LAYER M1 ;
        RECT 16.399 9.744 16.401 12.18 ;
  LAYER M1 ;
        RECT 16.479 9.744 16.481 12.18 ;
  LAYER M2 ;
        RECT 14.16 9.743 16.56 9.745 ;
  LAYER M2 ;
        RECT 14.16 9.827 16.56 9.829 ;
  LAYER M2 ;
        RECT 14.16 9.911 16.56 9.913 ;
  LAYER M2 ;
        RECT 14.16 9.995 16.56 9.997 ;
  LAYER M2 ;
        RECT 14.16 10.079 16.56 10.081 ;
  LAYER M2 ;
        RECT 14.16 10.163 16.56 10.165 ;
  LAYER M2 ;
        RECT 14.16 10.247 16.56 10.249 ;
  LAYER M2 ;
        RECT 14.16 10.331 16.56 10.333 ;
  LAYER M2 ;
        RECT 14.16 10.415 16.56 10.417 ;
  LAYER M2 ;
        RECT 14.16 10.499 16.56 10.501 ;
  LAYER M2 ;
        RECT 14.16 10.583 16.56 10.585 ;
  LAYER M2 ;
        RECT 14.16 10.667 16.56 10.669 ;
  LAYER M2 ;
        RECT 14.16 10.7505 16.56 10.7525 ;
  LAYER M2 ;
        RECT 14.16 10.835 16.56 10.837 ;
  LAYER M2 ;
        RECT 14.16 10.919 16.56 10.921 ;
  LAYER M2 ;
        RECT 14.16 11.003 16.56 11.005 ;
  LAYER M2 ;
        RECT 14.16 11.087 16.56 11.089 ;
  LAYER M2 ;
        RECT 14.16 11.171 16.56 11.173 ;
  LAYER M2 ;
        RECT 14.16 11.255 16.56 11.257 ;
  LAYER M2 ;
        RECT 14.16 11.339 16.56 11.341 ;
  LAYER M2 ;
        RECT 14.16 11.423 16.56 11.425 ;
  LAYER M2 ;
        RECT 14.16 11.507 16.56 11.509 ;
  LAYER M2 ;
        RECT 14.16 11.591 16.56 11.593 ;
  LAYER M2 ;
        RECT 14.16 11.675 16.56 11.677 ;
  LAYER M2 ;
        RECT 14.16 11.759 16.56 11.761 ;
  LAYER M2 ;
        RECT 14.16 11.843 16.56 11.845 ;
  LAYER M2 ;
        RECT 14.16 11.927 16.56 11.929 ;
  LAYER M2 ;
        RECT 14.16 12.011 16.56 12.013 ;
  LAYER M2 ;
        RECT 14.16 12.095 16.56 12.097 ;
  LAYER M1 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M1 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M1 ;
        RECT 14.272 12.648 14.304 15.156 ;
  LAYER M1 ;
        RECT 14.336 12.648 14.368 15.156 ;
  LAYER M1 ;
        RECT 14.4 12.648 14.432 15.156 ;
  LAYER M1 ;
        RECT 14.464 12.648 14.496 15.156 ;
  LAYER M1 ;
        RECT 14.528 12.648 14.56 15.156 ;
  LAYER M1 ;
        RECT 14.592 12.648 14.624 15.156 ;
  LAYER M1 ;
        RECT 14.656 12.648 14.688 15.156 ;
  LAYER M1 ;
        RECT 14.72 12.648 14.752 15.156 ;
  LAYER M1 ;
        RECT 14.784 12.648 14.816 15.156 ;
  LAYER M1 ;
        RECT 14.848 12.648 14.88 15.156 ;
  LAYER M1 ;
        RECT 14.912 12.648 14.944 15.156 ;
  LAYER M1 ;
        RECT 14.976 12.648 15.008 15.156 ;
  LAYER M1 ;
        RECT 15.04 12.648 15.072 15.156 ;
  LAYER M1 ;
        RECT 15.104 12.648 15.136 15.156 ;
  LAYER M1 ;
        RECT 15.168 12.648 15.2 15.156 ;
  LAYER M1 ;
        RECT 15.232 12.648 15.264 15.156 ;
  LAYER M1 ;
        RECT 15.296 12.648 15.328 15.156 ;
  LAYER M1 ;
        RECT 15.36 12.648 15.392 15.156 ;
  LAYER M1 ;
        RECT 15.424 12.648 15.456 15.156 ;
  LAYER M1 ;
        RECT 15.488 12.648 15.52 15.156 ;
  LAYER M1 ;
        RECT 15.552 12.648 15.584 15.156 ;
  LAYER M1 ;
        RECT 15.616 12.648 15.648 15.156 ;
  LAYER M1 ;
        RECT 15.68 12.648 15.712 15.156 ;
  LAYER M1 ;
        RECT 15.744 12.648 15.776 15.156 ;
  LAYER M1 ;
        RECT 15.808 12.648 15.84 15.156 ;
  LAYER M1 ;
        RECT 15.872 12.648 15.904 15.156 ;
  LAYER M1 ;
        RECT 15.936 12.648 15.968 15.156 ;
  LAYER M1 ;
        RECT 16 12.648 16.032 15.156 ;
  LAYER M1 ;
        RECT 16.064 12.648 16.096 15.156 ;
  LAYER M1 ;
        RECT 16.128 12.648 16.16 15.156 ;
  LAYER M1 ;
        RECT 16.192 12.648 16.224 15.156 ;
  LAYER M1 ;
        RECT 16.256 12.648 16.288 15.156 ;
  LAYER M1 ;
        RECT 16.32 12.648 16.352 15.156 ;
  LAYER M1 ;
        RECT 16.384 12.648 16.416 15.156 ;
  LAYER M1 ;
        RECT 16.448 12.648 16.48 15.156 ;
  LAYER M2 ;
        RECT 14.124 12.732 16.596 12.764 ;
  LAYER M2 ;
        RECT 14.124 12.796 16.596 12.828 ;
  LAYER M2 ;
        RECT 14.124 12.86 16.596 12.892 ;
  LAYER M2 ;
        RECT 14.124 12.924 16.596 12.956 ;
  LAYER M2 ;
        RECT 14.124 12.988 16.596 13.02 ;
  LAYER M2 ;
        RECT 14.124 13.052 16.596 13.084 ;
  LAYER M2 ;
        RECT 14.124 13.116 16.596 13.148 ;
  LAYER M2 ;
        RECT 14.124 13.18 16.596 13.212 ;
  LAYER M2 ;
        RECT 14.124 13.244 16.596 13.276 ;
  LAYER M2 ;
        RECT 14.124 13.308 16.596 13.34 ;
  LAYER M2 ;
        RECT 14.124 13.372 16.596 13.404 ;
  LAYER M2 ;
        RECT 14.124 13.436 16.596 13.468 ;
  LAYER M2 ;
        RECT 14.124 13.5 16.596 13.532 ;
  LAYER M2 ;
        RECT 14.124 13.564 16.596 13.596 ;
  LAYER M2 ;
        RECT 14.124 13.628 16.596 13.66 ;
  LAYER M2 ;
        RECT 14.124 13.692 16.596 13.724 ;
  LAYER M2 ;
        RECT 14.124 13.756 16.596 13.788 ;
  LAYER M2 ;
        RECT 14.124 13.82 16.596 13.852 ;
  LAYER M2 ;
        RECT 14.124 13.884 16.596 13.916 ;
  LAYER M2 ;
        RECT 14.124 13.948 16.596 13.98 ;
  LAYER M2 ;
        RECT 14.124 14.012 16.596 14.044 ;
  LAYER M2 ;
        RECT 14.124 14.076 16.596 14.108 ;
  LAYER M2 ;
        RECT 14.124 14.14 16.596 14.172 ;
  LAYER M2 ;
        RECT 14.124 14.204 16.596 14.236 ;
  LAYER M2 ;
        RECT 14.124 14.268 16.596 14.3 ;
  LAYER M2 ;
        RECT 14.124 14.332 16.596 14.364 ;
  LAYER M2 ;
        RECT 14.124 14.396 16.596 14.428 ;
  LAYER M2 ;
        RECT 14.124 14.46 16.596 14.492 ;
  LAYER M2 ;
        RECT 14.124 14.524 16.596 14.556 ;
  LAYER M2 ;
        RECT 14.124 14.588 16.596 14.62 ;
  LAYER M2 ;
        RECT 14.124 14.652 16.596 14.684 ;
  LAYER M2 ;
        RECT 14.124 14.716 16.596 14.748 ;
  LAYER M2 ;
        RECT 14.124 14.78 16.596 14.812 ;
  LAYER M2 ;
        RECT 14.124 14.844 16.596 14.876 ;
  LAYER M2 ;
        RECT 14.124 14.908 16.596 14.94 ;
  LAYER M2 ;
        RECT 14.124 14.972 16.596 15.004 ;
  LAYER M3 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M3 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M3 ;
        RECT 14.272 12.648 14.304 15.156 ;
  LAYER M3 ;
        RECT 14.336 12.648 14.368 15.156 ;
  LAYER M3 ;
        RECT 14.4 12.648 14.432 15.156 ;
  LAYER M3 ;
        RECT 14.464 12.648 14.496 15.156 ;
  LAYER M3 ;
        RECT 14.528 12.648 14.56 15.156 ;
  LAYER M3 ;
        RECT 14.592 12.648 14.624 15.156 ;
  LAYER M3 ;
        RECT 14.656 12.648 14.688 15.156 ;
  LAYER M3 ;
        RECT 14.72 12.648 14.752 15.156 ;
  LAYER M3 ;
        RECT 14.784 12.648 14.816 15.156 ;
  LAYER M3 ;
        RECT 14.848 12.648 14.88 15.156 ;
  LAYER M3 ;
        RECT 14.912 12.648 14.944 15.156 ;
  LAYER M3 ;
        RECT 14.976 12.648 15.008 15.156 ;
  LAYER M3 ;
        RECT 15.04 12.648 15.072 15.156 ;
  LAYER M3 ;
        RECT 15.104 12.648 15.136 15.156 ;
  LAYER M3 ;
        RECT 15.168 12.648 15.2 15.156 ;
  LAYER M3 ;
        RECT 15.232 12.648 15.264 15.156 ;
  LAYER M3 ;
        RECT 15.296 12.648 15.328 15.156 ;
  LAYER M3 ;
        RECT 15.36 12.648 15.392 15.156 ;
  LAYER M3 ;
        RECT 15.424 12.648 15.456 15.156 ;
  LAYER M3 ;
        RECT 15.488 12.648 15.52 15.156 ;
  LAYER M3 ;
        RECT 15.552 12.648 15.584 15.156 ;
  LAYER M3 ;
        RECT 15.616 12.648 15.648 15.156 ;
  LAYER M3 ;
        RECT 15.68 12.648 15.712 15.156 ;
  LAYER M3 ;
        RECT 15.744 12.648 15.776 15.156 ;
  LAYER M3 ;
        RECT 15.808 12.648 15.84 15.156 ;
  LAYER M3 ;
        RECT 15.872 12.648 15.904 15.156 ;
  LAYER M3 ;
        RECT 15.936 12.648 15.968 15.156 ;
  LAYER M3 ;
        RECT 16 12.648 16.032 15.156 ;
  LAYER M3 ;
        RECT 16.064 12.648 16.096 15.156 ;
  LAYER M3 ;
        RECT 16.128 12.648 16.16 15.156 ;
  LAYER M3 ;
        RECT 16.192 12.648 16.224 15.156 ;
  LAYER M3 ;
        RECT 16.256 12.648 16.288 15.156 ;
  LAYER M3 ;
        RECT 16.32 12.648 16.352 15.156 ;
  LAYER M3 ;
        RECT 16.384 12.648 16.416 15.156 ;
  LAYER M3 ;
        RECT 16.448 12.648 16.48 15.156 ;
  LAYER M3 ;
        RECT 16.544 12.648 16.576 15.156 ;
  LAYER M1 ;
        RECT 14.159 12.684 14.161 15.12 ;
  LAYER M1 ;
        RECT 14.239 12.684 14.241 15.12 ;
  LAYER M1 ;
        RECT 14.319 12.684 14.321 15.12 ;
  LAYER M1 ;
        RECT 14.399 12.684 14.401 15.12 ;
  LAYER M1 ;
        RECT 14.479 12.684 14.481 15.12 ;
  LAYER M1 ;
        RECT 14.559 12.684 14.561 15.12 ;
  LAYER M1 ;
        RECT 14.639 12.684 14.641 15.12 ;
  LAYER M1 ;
        RECT 14.719 12.684 14.721 15.12 ;
  LAYER M1 ;
        RECT 14.799 12.684 14.801 15.12 ;
  LAYER M1 ;
        RECT 14.879 12.684 14.881 15.12 ;
  LAYER M1 ;
        RECT 14.959 12.684 14.961 15.12 ;
  LAYER M1 ;
        RECT 15.039 12.684 15.041 15.12 ;
  LAYER M1 ;
        RECT 15.119 12.684 15.121 15.12 ;
  LAYER M1 ;
        RECT 15.199 12.684 15.201 15.12 ;
  LAYER M1 ;
        RECT 15.279 12.684 15.281 15.12 ;
  LAYER M1 ;
        RECT 15.359 12.684 15.361 15.12 ;
  LAYER M1 ;
        RECT 15.439 12.684 15.441 15.12 ;
  LAYER M1 ;
        RECT 15.519 12.684 15.521 15.12 ;
  LAYER M1 ;
        RECT 15.599 12.684 15.601 15.12 ;
  LAYER M1 ;
        RECT 15.679 12.684 15.681 15.12 ;
  LAYER M1 ;
        RECT 15.759 12.684 15.761 15.12 ;
  LAYER M1 ;
        RECT 15.839 12.684 15.841 15.12 ;
  LAYER M1 ;
        RECT 15.919 12.684 15.921 15.12 ;
  LAYER M1 ;
        RECT 15.999 12.684 16.001 15.12 ;
  LAYER M1 ;
        RECT 16.079 12.684 16.081 15.12 ;
  LAYER M1 ;
        RECT 16.159 12.684 16.161 15.12 ;
  LAYER M1 ;
        RECT 16.239 12.684 16.241 15.12 ;
  LAYER M1 ;
        RECT 16.319 12.684 16.321 15.12 ;
  LAYER M1 ;
        RECT 16.399 12.684 16.401 15.12 ;
  LAYER M1 ;
        RECT 16.479 12.684 16.481 15.12 ;
  LAYER M2 ;
        RECT 14.16 12.683 16.56 12.685 ;
  LAYER M2 ;
        RECT 14.16 12.767 16.56 12.769 ;
  LAYER M2 ;
        RECT 14.16 12.851 16.56 12.853 ;
  LAYER M2 ;
        RECT 14.16 12.935 16.56 12.937 ;
  LAYER M2 ;
        RECT 14.16 13.019 16.56 13.021 ;
  LAYER M2 ;
        RECT 14.16 13.103 16.56 13.105 ;
  LAYER M2 ;
        RECT 14.16 13.187 16.56 13.189 ;
  LAYER M2 ;
        RECT 14.16 13.271 16.56 13.273 ;
  LAYER M2 ;
        RECT 14.16 13.355 16.56 13.357 ;
  LAYER M2 ;
        RECT 14.16 13.439 16.56 13.441 ;
  LAYER M2 ;
        RECT 14.16 13.523 16.56 13.525 ;
  LAYER M2 ;
        RECT 14.16 13.607 16.56 13.609 ;
  LAYER M2 ;
        RECT 14.16 13.6905 16.56 13.6925 ;
  LAYER M2 ;
        RECT 14.16 13.775 16.56 13.777 ;
  LAYER M2 ;
        RECT 14.16 13.859 16.56 13.861 ;
  LAYER M2 ;
        RECT 14.16 13.943 16.56 13.945 ;
  LAYER M2 ;
        RECT 14.16 14.027 16.56 14.029 ;
  LAYER M2 ;
        RECT 14.16 14.111 16.56 14.113 ;
  LAYER M2 ;
        RECT 14.16 14.195 16.56 14.197 ;
  LAYER M2 ;
        RECT 14.16 14.279 16.56 14.281 ;
  LAYER M2 ;
        RECT 14.16 14.363 16.56 14.365 ;
  LAYER M2 ;
        RECT 14.16 14.447 16.56 14.449 ;
  LAYER M2 ;
        RECT 14.16 14.531 16.56 14.533 ;
  LAYER M2 ;
        RECT 14.16 14.615 16.56 14.617 ;
  LAYER M2 ;
        RECT 14.16 14.699 16.56 14.701 ;
  LAYER M2 ;
        RECT 14.16 14.783 16.56 14.785 ;
  LAYER M2 ;
        RECT 14.16 14.867 16.56 14.869 ;
  LAYER M2 ;
        RECT 14.16 14.951 16.56 14.953 ;
  LAYER M2 ;
        RECT 14.16 15.035 16.56 15.037 ;
  LAYER M1 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M1 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M1 ;
        RECT 14.272 15.588 14.304 18.096 ;
  LAYER M1 ;
        RECT 14.336 15.588 14.368 18.096 ;
  LAYER M1 ;
        RECT 14.4 15.588 14.432 18.096 ;
  LAYER M1 ;
        RECT 14.464 15.588 14.496 18.096 ;
  LAYER M1 ;
        RECT 14.528 15.588 14.56 18.096 ;
  LAYER M1 ;
        RECT 14.592 15.588 14.624 18.096 ;
  LAYER M1 ;
        RECT 14.656 15.588 14.688 18.096 ;
  LAYER M1 ;
        RECT 14.72 15.588 14.752 18.096 ;
  LAYER M1 ;
        RECT 14.784 15.588 14.816 18.096 ;
  LAYER M1 ;
        RECT 14.848 15.588 14.88 18.096 ;
  LAYER M1 ;
        RECT 14.912 15.588 14.944 18.096 ;
  LAYER M1 ;
        RECT 14.976 15.588 15.008 18.096 ;
  LAYER M1 ;
        RECT 15.04 15.588 15.072 18.096 ;
  LAYER M1 ;
        RECT 15.104 15.588 15.136 18.096 ;
  LAYER M1 ;
        RECT 15.168 15.588 15.2 18.096 ;
  LAYER M1 ;
        RECT 15.232 15.588 15.264 18.096 ;
  LAYER M1 ;
        RECT 15.296 15.588 15.328 18.096 ;
  LAYER M1 ;
        RECT 15.36 15.588 15.392 18.096 ;
  LAYER M1 ;
        RECT 15.424 15.588 15.456 18.096 ;
  LAYER M1 ;
        RECT 15.488 15.588 15.52 18.096 ;
  LAYER M1 ;
        RECT 15.552 15.588 15.584 18.096 ;
  LAYER M1 ;
        RECT 15.616 15.588 15.648 18.096 ;
  LAYER M1 ;
        RECT 15.68 15.588 15.712 18.096 ;
  LAYER M1 ;
        RECT 15.744 15.588 15.776 18.096 ;
  LAYER M1 ;
        RECT 15.808 15.588 15.84 18.096 ;
  LAYER M1 ;
        RECT 15.872 15.588 15.904 18.096 ;
  LAYER M1 ;
        RECT 15.936 15.588 15.968 18.096 ;
  LAYER M1 ;
        RECT 16 15.588 16.032 18.096 ;
  LAYER M1 ;
        RECT 16.064 15.588 16.096 18.096 ;
  LAYER M1 ;
        RECT 16.128 15.588 16.16 18.096 ;
  LAYER M1 ;
        RECT 16.192 15.588 16.224 18.096 ;
  LAYER M1 ;
        RECT 16.256 15.588 16.288 18.096 ;
  LAYER M1 ;
        RECT 16.32 15.588 16.352 18.096 ;
  LAYER M1 ;
        RECT 16.384 15.588 16.416 18.096 ;
  LAYER M1 ;
        RECT 16.448 15.588 16.48 18.096 ;
  LAYER M2 ;
        RECT 14.124 15.672 16.596 15.704 ;
  LAYER M2 ;
        RECT 14.124 15.736 16.596 15.768 ;
  LAYER M2 ;
        RECT 14.124 15.8 16.596 15.832 ;
  LAYER M2 ;
        RECT 14.124 15.864 16.596 15.896 ;
  LAYER M2 ;
        RECT 14.124 15.928 16.596 15.96 ;
  LAYER M2 ;
        RECT 14.124 15.992 16.596 16.024 ;
  LAYER M2 ;
        RECT 14.124 16.056 16.596 16.088 ;
  LAYER M2 ;
        RECT 14.124 16.12 16.596 16.152 ;
  LAYER M2 ;
        RECT 14.124 16.184 16.596 16.216 ;
  LAYER M2 ;
        RECT 14.124 16.248 16.596 16.28 ;
  LAYER M2 ;
        RECT 14.124 16.312 16.596 16.344 ;
  LAYER M2 ;
        RECT 14.124 16.376 16.596 16.408 ;
  LAYER M2 ;
        RECT 14.124 16.44 16.596 16.472 ;
  LAYER M2 ;
        RECT 14.124 16.504 16.596 16.536 ;
  LAYER M2 ;
        RECT 14.124 16.568 16.596 16.6 ;
  LAYER M2 ;
        RECT 14.124 16.632 16.596 16.664 ;
  LAYER M2 ;
        RECT 14.124 16.696 16.596 16.728 ;
  LAYER M2 ;
        RECT 14.124 16.76 16.596 16.792 ;
  LAYER M2 ;
        RECT 14.124 16.824 16.596 16.856 ;
  LAYER M2 ;
        RECT 14.124 16.888 16.596 16.92 ;
  LAYER M2 ;
        RECT 14.124 16.952 16.596 16.984 ;
  LAYER M2 ;
        RECT 14.124 17.016 16.596 17.048 ;
  LAYER M2 ;
        RECT 14.124 17.08 16.596 17.112 ;
  LAYER M2 ;
        RECT 14.124 17.144 16.596 17.176 ;
  LAYER M2 ;
        RECT 14.124 17.208 16.596 17.24 ;
  LAYER M2 ;
        RECT 14.124 17.272 16.596 17.304 ;
  LAYER M2 ;
        RECT 14.124 17.336 16.596 17.368 ;
  LAYER M2 ;
        RECT 14.124 17.4 16.596 17.432 ;
  LAYER M2 ;
        RECT 14.124 17.464 16.596 17.496 ;
  LAYER M2 ;
        RECT 14.124 17.528 16.596 17.56 ;
  LAYER M2 ;
        RECT 14.124 17.592 16.596 17.624 ;
  LAYER M2 ;
        RECT 14.124 17.656 16.596 17.688 ;
  LAYER M2 ;
        RECT 14.124 17.72 16.596 17.752 ;
  LAYER M2 ;
        RECT 14.124 17.784 16.596 17.816 ;
  LAYER M2 ;
        RECT 14.124 17.848 16.596 17.88 ;
  LAYER M2 ;
        RECT 14.124 17.912 16.596 17.944 ;
  LAYER M3 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M3 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M3 ;
        RECT 14.272 15.588 14.304 18.096 ;
  LAYER M3 ;
        RECT 14.336 15.588 14.368 18.096 ;
  LAYER M3 ;
        RECT 14.4 15.588 14.432 18.096 ;
  LAYER M3 ;
        RECT 14.464 15.588 14.496 18.096 ;
  LAYER M3 ;
        RECT 14.528 15.588 14.56 18.096 ;
  LAYER M3 ;
        RECT 14.592 15.588 14.624 18.096 ;
  LAYER M3 ;
        RECT 14.656 15.588 14.688 18.096 ;
  LAYER M3 ;
        RECT 14.72 15.588 14.752 18.096 ;
  LAYER M3 ;
        RECT 14.784 15.588 14.816 18.096 ;
  LAYER M3 ;
        RECT 14.848 15.588 14.88 18.096 ;
  LAYER M3 ;
        RECT 14.912 15.588 14.944 18.096 ;
  LAYER M3 ;
        RECT 14.976 15.588 15.008 18.096 ;
  LAYER M3 ;
        RECT 15.04 15.588 15.072 18.096 ;
  LAYER M3 ;
        RECT 15.104 15.588 15.136 18.096 ;
  LAYER M3 ;
        RECT 15.168 15.588 15.2 18.096 ;
  LAYER M3 ;
        RECT 15.232 15.588 15.264 18.096 ;
  LAYER M3 ;
        RECT 15.296 15.588 15.328 18.096 ;
  LAYER M3 ;
        RECT 15.36 15.588 15.392 18.096 ;
  LAYER M3 ;
        RECT 15.424 15.588 15.456 18.096 ;
  LAYER M3 ;
        RECT 15.488 15.588 15.52 18.096 ;
  LAYER M3 ;
        RECT 15.552 15.588 15.584 18.096 ;
  LAYER M3 ;
        RECT 15.616 15.588 15.648 18.096 ;
  LAYER M3 ;
        RECT 15.68 15.588 15.712 18.096 ;
  LAYER M3 ;
        RECT 15.744 15.588 15.776 18.096 ;
  LAYER M3 ;
        RECT 15.808 15.588 15.84 18.096 ;
  LAYER M3 ;
        RECT 15.872 15.588 15.904 18.096 ;
  LAYER M3 ;
        RECT 15.936 15.588 15.968 18.096 ;
  LAYER M3 ;
        RECT 16 15.588 16.032 18.096 ;
  LAYER M3 ;
        RECT 16.064 15.588 16.096 18.096 ;
  LAYER M3 ;
        RECT 16.128 15.588 16.16 18.096 ;
  LAYER M3 ;
        RECT 16.192 15.588 16.224 18.096 ;
  LAYER M3 ;
        RECT 16.256 15.588 16.288 18.096 ;
  LAYER M3 ;
        RECT 16.32 15.588 16.352 18.096 ;
  LAYER M3 ;
        RECT 16.384 15.588 16.416 18.096 ;
  LAYER M3 ;
        RECT 16.448 15.588 16.48 18.096 ;
  LAYER M3 ;
        RECT 16.544 15.588 16.576 18.096 ;
  LAYER M1 ;
        RECT 14.159 15.624 14.161 18.06 ;
  LAYER M1 ;
        RECT 14.239 15.624 14.241 18.06 ;
  LAYER M1 ;
        RECT 14.319 15.624 14.321 18.06 ;
  LAYER M1 ;
        RECT 14.399 15.624 14.401 18.06 ;
  LAYER M1 ;
        RECT 14.479 15.624 14.481 18.06 ;
  LAYER M1 ;
        RECT 14.559 15.624 14.561 18.06 ;
  LAYER M1 ;
        RECT 14.639 15.624 14.641 18.06 ;
  LAYER M1 ;
        RECT 14.719 15.624 14.721 18.06 ;
  LAYER M1 ;
        RECT 14.799 15.624 14.801 18.06 ;
  LAYER M1 ;
        RECT 14.879 15.624 14.881 18.06 ;
  LAYER M1 ;
        RECT 14.959 15.624 14.961 18.06 ;
  LAYER M1 ;
        RECT 15.039 15.624 15.041 18.06 ;
  LAYER M1 ;
        RECT 15.119 15.624 15.121 18.06 ;
  LAYER M1 ;
        RECT 15.199 15.624 15.201 18.06 ;
  LAYER M1 ;
        RECT 15.279 15.624 15.281 18.06 ;
  LAYER M1 ;
        RECT 15.359 15.624 15.361 18.06 ;
  LAYER M1 ;
        RECT 15.439 15.624 15.441 18.06 ;
  LAYER M1 ;
        RECT 15.519 15.624 15.521 18.06 ;
  LAYER M1 ;
        RECT 15.599 15.624 15.601 18.06 ;
  LAYER M1 ;
        RECT 15.679 15.624 15.681 18.06 ;
  LAYER M1 ;
        RECT 15.759 15.624 15.761 18.06 ;
  LAYER M1 ;
        RECT 15.839 15.624 15.841 18.06 ;
  LAYER M1 ;
        RECT 15.919 15.624 15.921 18.06 ;
  LAYER M1 ;
        RECT 15.999 15.624 16.001 18.06 ;
  LAYER M1 ;
        RECT 16.079 15.624 16.081 18.06 ;
  LAYER M1 ;
        RECT 16.159 15.624 16.161 18.06 ;
  LAYER M1 ;
        RECT 16.239 15.624 16.241 18.06 ;
  LAYER M1 ;
        RECT 16.319 15.624 16.321 18.06 ;
  LAYER M1 ;
        RECT 16.399 15.624 16.401 18.06 ;
  LAYER M1 ;
        RECT 16.479 15.624 16.481 18.06 ;
  LAYER M2 ;
        RECT 14.16 15.623 16.56 15.625 ;
  LAYER M2 ;
        RECT 14.16 15.707 16.56 15.709 ;
  LAYER M2 ;
        RECT 14.16 15.791 16.56 15.793 ;
  LAYER M2 ;
        RECT 14.16 15.875 16.56 15.877 ;
  LAYER M2 ;
        RECT 14.16 15.959 16.56 15.961 ;
  LAYER M2 ;
        RECT 14.16 16.043 16.56 16.045 ;
  LAYER M2 ;
        RECT 14.16 16.127 16.56 16.129 ;
  LAYER M2 ;
        RECT 14.16 16.211 16.56 16.213 ;
  LAYER M2 ;
        RECT 14.16 16.295 16.56 16.297 ;
  LAYER M2 ;
        RECT 14.16 16.379 16.56 16.381 ;
  LAYER M2 ;
        RECT 14.16 16.463 16.56 16.465 ;
  LAYER M2 ;
        RECT 14.16 16.547 16.56 16.549 ;
  LAYER M2 ;
        RECT 14.16 16.6305 16.56 16.6325 ;
  LAYER M2 ;
        RECT 14.16 16.715 16.56 16.717 ;
  LAYER M2 ;
        RECT 14.16 16.799 16.56 16.801 ;
  LAYER M2 ;
        RECT 14.16 16.883 16.56 16.885 ;
  LAYER M2 ;
        RECT 14.16 16.967 16.56 16.969 ;
  LAYER M2 ;
        RECT 14.16 17.051 16.56 17.053 ;
  LAYER M2 ;
        RECT 14.16 17.135 16.56 17.137 ;
  LAYER M2 ;
        RECT 14.16 17.219 16.56 17.221 ;
  LAYER M2 ;
        RECT 14.16 17.303 16.56 17.305 ;
  LAYER M2 ;
        RECT 14.16 17.387 16.56 17.389 ;
  LAYER M2 ;
        RECT 14.16 17.471 16.56 17.473 ;
  LAYER M2 ;
        RECT 14.16 17.555 16.56 17.557 ;
  LAYER M2 ;
        RECT 14.16 17.639 16.56 17.641 ;
  LAYER M2 ;
        RECT 14.16 17.723 16.56 17.725 ;
  LAYER M2 ;
        RECT 14.16 17.807 16.56 17.809 ;
  LAYER M2 ;
        RECT 14.16 17.891 16.56 17.893 ;
  LAYER M2 ;
        RECT 14.16 17.975 16.56 17.977 ;
  END 
END Cap_30fF_Cap_60fF
