MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 12.16 BY 19.992 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 19.536 3.232 19.608 ;
      LAYER M2 ;
        RECT 3.18 19.556 3.252 19.588 ;
      LAYER M1 ;
        RECT 9.152 19.536 9.184 19.608 ;
      LAYER M2 ;
        RECT 9.132 19.556 9.204 19.588 ;
      LAYER M2 ;
        RECT 3.216 19.556 9.168 19.588 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
      LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 19.704 6.208 19.776 ;
      LAYER M2 ;
        RECT 6.156 19.724 6.228 19.756 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
      LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M2 ;
        RECT 6.032 10.316 8.784 10.348 ;
  LAYER M1 ;
        RECT 6.016 10.296 6.048 10.368 ;
  LAYER M2 ;
        RECT 5.996 10.316 6.068 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.164 5.824 10.332 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M2 ;
        RECT 6.032 7.208 8.784 7.24 ;
  LAYER M1 ;
        RECT 6.016 7.188 6.048 7.26 ;
  LAYER M2 ;
        RECT 5.996 7.208 6.068 7.24 ;
  LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
  LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
  LAYER M1 ;
        RECT 6.016 0.42 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 10.332 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M2 ;
        RECT 3.056 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 3.04 7.188 3.072 7.26 ;
  LAYER M2 ;
        RECT 3.02 7.208 3.092 7.24 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M2 ;
        RECT 3.056 13.424 5.808 13.456 ;
  LAYER M1 ;
        RECT 3.04 13.404 3.072 13.476 ;
  LAYER M2 ;
        RECT 3.02 13.424 3.092 13.456 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 13.44 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M1 ;
        RECT 8.768 3.948 8.8 4.116 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 8.784 3.932 9.008 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
  LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
  LAYER M1 ;
        RECT 8.992 0.252 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 3.948 ;
  LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 2.832 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 2.832 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 2.832 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 2.832 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 2.832 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 2.816 16.512 2.848 16.584 ;
  LAYER M2 ;
        RECT 2.796 16.532 2.868 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 2.832 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 16.548 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.84 11.776 1.008 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M2 ;
        RECT 11.76 0.824 11.984 0.856 ;
  LAYER M1 ;
        RECT 11.968 0.804 12 0.876 ;
  LAYER M2 ;
        RECT 11.948 0.824 12.02 0.856 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M1 ;
        RECT 11.744 3.948 11.776 4.116 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 11.76 3.932 11.984 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M1 ;
        RECT 11.744 7.056 11.776 7.224 ;
  LAYER M1 ;
        RECT 11.744 7.02 11.776 7.092 ;
  LAYER M2 ;
        RECT 11.724 7.04 11.796 7.072 ;
  LAYER M2 ;
        RECT 11.76 7.04 11.984 7.072 ;
  LAYER M1 ;
        RECT 11.968 7.02 12 7.092 ;
  LAYER M2 ;
        RECT 11.948 7.04 12.02 7.072 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M1 ;
        RECT 11.744 10.164 11.776 10.332 ;
  LAYER M1 ;
        RECT 11.744 10.128 11.776 10.2 ;
  LAYER M2 ;
        RECT 11.724 10.148 11.796 10.18 ;
  LAYER M2 ;
        RECT 11.76 10.148 11.984 10.18 ;
  LAYER M1 ;
        RECT 11.968 10.128 12 10.2 ;
  LAYER M2 ;
        RECT 11.948 10.148 12.02 10.18 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 13.476 ;
  LAYER M2 ;
        RECT 11.724 13.424 11.796 13.456 ;
  LAYER M1 ;
        RECT 11.744 13.272 11.776 13.44 ;
  LAYER M1 ;
        RECT 11.744 13.236 11.776 13.308 ;
  LAYER M2 ;
        RECT 11.724 13.256 11.796 13.288 ;
  LAYER M2 ;
        RECT 11.76 13.256 11.984 13.288 ;
  LAYER M1 ;
        RECT 11.968 13.236 12 13.308 ;
  LAYER M2 ;
        RECT 11.948 13.256 12.02 13.288 ;
  LAYER M1 ;
        RECT 11.744 16.512 11.776 16.584 ;
  LAYER M2 ;
        RECT 11.724 16.532 11.796 16.564 ;
  LAYER M1 ;
        RECT 11.744 16.38 11.776 16.548 ;
  LAYER M1 ;
        RECT 11.744 16.344 11.776 16.416 ;
  LAYER M2 ;
        RECT 11.724 16.364 11.796 16.396 ;
  LAYER M2 ;
        RECT 11.76 16.364 11.984 16.396 ;
  LAYER M1 ;
        RECT 11.968 16.344 12 16.416 ;
  LAYER M2 ;
        RECT 11.948 16.364 12.02 16.396 ;
  LAYER M1 ;
        RECT 11.968 0.048 12 0.12 ;
  LAYER M2 ;
        RECT 11.948 0.068 12.02 0.1 ;
  LAYER M1 ;
        RECT 11.968 0.084 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 16.38 ;
  LAYER M2 ;
        RECT 0.08 0.068 11.984 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 2.832 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M2 ;
        RECT 2.832 4.1 5.808 4.132 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M1 ;
        RECT 5.792 16.512 5.824 16.584 ;
  LAYER M2 ;
        RECT 5.772 16.532 5.844 16.564 ;
  LAYER M2 ;
        RECT 2.832 16.532 5.808 16.564 ;
  LAYER M1 ;
        RECT 2.816 16.512 2.848 16.584 ;
  LAYER M2 ;
        RECT 2.796 16.532 2.868 16.564 ;
  LAYER M1 ;
        RECT 8.768 16.512 8.8 16.584 ;
  LAYER M2 ;
        RECT 8.748 16.532 8.82 16.564 ;
  LAYER M2 ;
        RECT 5.808 16.532 8.784 16.564 ;
  LAYER M1 ;
        RECT 5.792 16.512 5.824 16.584 ;
  LAYER M2 ;
        RECT 5.772 16.532 5.844 16.564 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M1 ;
        RECT 8.768 13.44 8.8 16.548 ;
  LAYER M1 ;
        RECT 8.768 16.512 8.8 16.584 ;
  LAYER M2 ;
        RECT 8.748 16.532 8.82 16.564 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.2 19.536 3.232 19.608 ;
  LAYER M2 ;
        RECT 3.18 19.556 3.252 19.588 ;
  LAYER M1 ;
        RECT 3.2 19.32 3.232 19.572 ;
  LAYER M1 ;
        RECT 3.2 12.768 3.232 19.32 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M1 ;
        RECT 6.4 12.768 6.432 12.936 ;
  LAYER M1 ;
        RECT 6.4 12.9 6.432 12.972 ;
  LAYER M2 ;
        RECT 6.38 12.92 6.452 12.952 ;
  LAYER M2 ;
        RECT 6.416 12.92 9.168 12.952 ;
  LAYER M1 ;
        RECT 9.152 12.9 9.184 12.972 ;
  LAYER M2 ;
        RECT 9.132 12.92 9.204 12.952 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M1 ;
        RECT 6.4 9.66 6.432 9.828 ;
  LAYER M1 ;
        RECT 6.4 9.792 6.432 9.864 ;
  LAYER M2 ;
        RECT 6.38 9.812 6.452 9.844 ;
  LAYER M2 ;
        RECT 6.416 9.812 9.168 9.844 ;
  LAYER M1 ;
        RECT 9.152 9.792 9.184 9.864 ;
  LAYER M2 ;
        RECT 9.132 9.812 9.204 9.844 ;
  LAYER M1 ;
        RECT 9.152 19.536 9.184 19.608 ;
  LAYER M2 ;
        RECT 9.132 19.556 9.204 19.588 ;
  LAYER M1 ;
        RECT 9.152 19.32 9.184 19.572 ;
  LAYER M1 ;
        RECT 9.152 9.828 9.184 19.32 ;
  LAYER M2 ;
        RECT 3.216 19.556 9.168 19.588 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M1 ;
        RECT 3.424 9.66 3.456 9.828 ;
  LAYER M1 ;
        RECT 3.424 9.792 3.456 9.864 ;
  LAYER M2 ;
        RECT 3.404 9.812 3.476 9.844 ;
  LAYER M2 ;
        RECT 3.44 9.812 6.192 9.844 ;
  LAYER M1 ;
        RECT 6.176 9.792 6.208 9.864 ;
  LAYER M2 ;
        RECT 6.156 9.812 6.228 9.844 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M1 ;
        RECT 3.424 15.876 3.456 16.044 ;
  LAYER M1 ;
        RECT 3.424 16.008 3.456 16.08 ;
  LAYER M2 ;
        RECT 3.404 16.028 3.476 16.06 ;
  LAYER M2 ;
        RECT 3.44 16.028 6.192 16.06 ;
  LAYER M1 ;
        RECT 6.176 16.008 6.208 16.08 ;
  LAYER M2 ;
        RECT 6.156 16.028 6.228 16.06 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.416 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 6.176 19.704 6.208 19.776 ;
  LAYER M2 ;
        RECT 6.156 19.724 6.228 19.756 ;
  LAYER M1 ;
        RECT 6.176 19.32 6.208 19.74 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 19.32 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.464 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.448 18.948 0.48 19.02 ;
  LAYER M2 ;
        RECT 0.428 18.968 0.5 19 ;
  LAYER M2 ;
        RECT 0.24 18.968 0.464 19 ;
  LAYER M1 ;
        RECT 0.224 18.948 0.256 19.02 ;
  LAYER M2 ;
        RECT 0.204 18.968 0.276 19 ;
  LAYER M1 ;
        RECT 0.224 19.872 0.256 19.944 ;
  LAYER M2 ;
        RECT 0.204 19.892 0.276 19.924 ;
  LAYER M1 ;
        RECT 0.224 19.32 0.256 19.908 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 19.32 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.444 9.408 3.612 ;
  LAYER M1 ;
        RECT 9.376 3.576 9.408 3.648 ;
  LAYER M2 ;
        RECT 9.356 3.596 9.428 3.628 ;
  LAYER M2 ;
        RECT 9.392 3.596 12.144 3.628 ;
  LAYER M1 ;
        RECT 12.128 3.576 12.16 3.648 ;
  LAYER M2 ;
        RECT 12.108 3.596 12.18 3.628 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.376 6.552 9.408 6.72 ;
  LAYER M1 ;
        RECT 9.376 6.684 9.408 6.756 ;
  LAYER M2 ;
        RECT 9.356 6.704 9.428 6.736 ;
  LAYER M2 ;
        RECT 9.392 6.704 12.144 6.736 ;
  LAYER M1 ;
        RECT 12.128 6.684 12.16 6.756 ;
  LAYER M2 ;
        RECT 12.108 6.704 12.18 6.736 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M1 ;
        RECT 9.376 9.66 9.408 9.828 ;
  LAYER M1 ;
        RECT 9.376 9.792 9.408 9.864 ;
  LAYER M2 ;
        RECT 9.356 9.812 9.428 9.844 ;
  LAYER M2 ;
        RECT 9.392 9.812 12.144 9.844 ;
  LAYER M1 ;
        RECT 12.128 9.792 12.16 9.864 ;
  LAYER M2 ;
        RECT 12.108 9.812 12.18 9.844 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M1 ;
        RECT 9.376 12.768 9.408 12.936 ;
  LAYER M1 ;
        RECT 9.376 12.9 9.408 12.972 ;
  LAYER M2 ;
        RECT 9.356 12.92 9.428 12.952 ;
  LAYER M2 ;
        RECT 9.392 12.92 12.144 12.952 ;
  LAYER M1 ;
        RECT 12.128 12.9 12.16 12.972 ;
  LAYER M2 ;
        RECT 12.108 12.92 12.18 12.952 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.876 9.408 16.044 ;
  LAYER M1 ;
        RECT 9.376 16.008 9.408 16.08 ;
  LAYER M2 ;
        RECT 9.356 16.028 9.428 16.06 ;
  LAYER M2 ;
        RECT 9.392 16.028 12.144 16.06 ;
  LAYER M1 ;
        RECT 12.128 16.008 12.16 16.08 ;
  LAYER M2 ;
        RECT 12.108 16.028 12.18 16.06 ;
  LAYER M1 ;
        RECT 9.376 18.948 9.408 19.02 ;
  LAYER M2 ;
        RECT 9.356 18.968 9.428 19 ;
  LAYER M1 ;
        RECT 9.376 18.984 9.408 19.152 ;
  LAYER M1 ;
        RECT 9.376 19.116 9.408 19.188 ;
  LAYER M2 ;
        RECT 9.356 19.136 9.428 19.168 ;
  LAYER M2 ;
        RECT 9.392 19.136 12.144 19.168 ;
  LAYER M1 ;
        RECT 12.128 19.116 12.16 19.188 ;
  LAYER M2 ;
        RECT 12.108 19.136 12.18 19.168 ;
  LAYER M1 ;
        RECT 12.128 19.872 12.16 19.944 ;
  LAYER M2 ;
        RECT 12.108 19.892 12.18 19.924 ;
  LAYER M1 ;
        RECT 12.128 19.32 12.16 19.908 ;
  LAYER M1 ;
        RECT 12.128 3.612 12.16 19.32 ;
  LAYER M2 ;
        RECT 0.24 19.892 12.144 19.924 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 0.464 6.536 3.44 6.568 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M1 ;
        RECT 3.424 18.948 3.456 19.02 ;
  LAYER M2 ;
        RECT 3.404 18.968 3.476 19 ;
  LAYER M2 ;
        RECT 0.464 18.968 3.44 19 ;
  LAYER M1 ;
        RECT 0.448 18.948 0.48 19.02 ;
  LAYER M2 ;
        RECT 0.428 18.968 0.5 19 ;
  LAYER M1 ;
        RECT 6.4 18.948 6.432 19.02 ;
  LAYER M2 ;
        RECT 6.38 18.968 6.452 19 ;
  LAYER M2 ;
        RECT 3.44 18.968 6.416 19 ;
  LAYER M1 ;
        RECT 3.424 18.948 3.456 19.02 ;
  LAYER M2 ;
        RECT 3.404 18.968 3.476 19 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.876 6.432 18.984 ;
  LAYER M1 ;
        RECT 6.4 18.948 6.432 19.02 ;
  LAYER M2 ;
        RECT 6.38 18.968 6.452 19 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M3 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M3 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M3 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M3 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M2 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M1 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M3 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M2 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M1 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M3 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M3 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M3 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M3 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M3 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M2 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M1 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M3 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M2 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M1 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M3 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M3 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M3 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M3 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M3 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M2 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M1 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M3 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M2 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M1 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M3 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M3 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M3 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M3 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M3 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M2 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M1 ;
        RECT 9.328 16.464 11.824 19.068 ;
  LAYER M3 ;
        RECT 9.328 16.464 11.824 19.068 ;
  LAYER M2 ;
        RECT 9.328 16.464 11.824 19.068 ;
  END 
END Cap_30fF_Cap_30fF
