
.subckt Sanitized_ResTune_Configure VDD VSS INPH RESEN<7> INPHASE<7> RESEN<6> INPHASE<6> RESEN<5> INPHASE<5> RESEN<4> INPHASE<4> RESEN<3> INPHASE<3> RESEN<2> INPHASE<2> RESEN<1> INPHASE<1> RESEN<0> INPHASE<0> OUTPH OUTPHASE<7> OUTPHASE<6> OUTPHASE<5> OUTPHASE<4> OUTPHASE<3> OUTPHASE<2> OUTPHASE<1> OUTPHASE<0>
XI3<1> VDD VSS DCAP8LVT
XI3<0> VDD VSS DCAP8LVT
XI2<7> VDD VSS DCAP16LVT
XI2<6> VDD VSS DCAP16LVT
XI2<5> VDD VSS DCAP16LVT
XI2<4> VDD VSS DCAP16LVT
XI2<3> VDD VSS DCAP16LVT
XI2<2> VDD VSS DCAP16LVT
XI2<1> VDD VSS DCAP16LVT
XI2<0> VDD VSS DCAP16LVT
XI4<3> VDD VSS DCAP32LVT
XI4<2> VDD VSS DCAP32LVT
XI4<1> VDD VSS DCAP32LVT
XI4<0> VDD VSS DCAP32LVT
XI1<7> INPH RESEN<7> VDD VSS INPHASE<7> BUFTD16LVT
XI1<6> INPH RESEN<6> VDD VSS INPHASE<6> BUFTD16LVT
XI1<5> INPH RESEN<5> VDD VSS INPHASE<5> BUFTD16LVT
XI1<4> INPH RESEN<4> VDD VSS INPHASE<4> BUFTD16LVT
XI1<3> INPH RESEN<3> VDD VSS INPHASE<3> BUFTD16LVT
XI1<2> INPH RESEN<2> VDD VSS INPHASE<2> BUFTD16LVT
XI1<1> INPH RESEN<1> VDD VSS INPHASE<1> BUFTD16LVT
XI1<0> INPH RESEN<0> VDD VSS INPHASE<0> BUFTD16LVT
XI0<7> OUTPH RESEN<7> VDD VSS OUTPHASE<7> BUFTD16LVT
XI0<6> OUTPH RESEN<6> VDD VSS OUTPHASE<6> BUFTD16LVT
XI0<5> OUTPH RESEN<5> VDD VSS OUTPHASE<5> BUFTD16LVT
XI0<4> OUTPH RESEN<4> VDD VSS OUTPHASE<4> BUFTD16LVT
XI0<3> OUTPH RESEN<3> VDD VSS OUTPHASE<3> BUFTD16LVT
XI0<2> OUTPH RESEN<2> VDD VSS OUTPHASE<2> BUFTD16LVT
XI0<1> OUTPH RESEN<1> VDD VSS OUTPHASE<1> BUFTD16LVT
XI0<0> OUTPH RESEN<0> VDD VSS OUTPHASE<0> BUFTD16LVT
.ends Sanitized_ResTune_Configure

.subckt DCAP8LVT 
xMMI4 VSS net9 VSS Dcap_NMOS_n12_X1_Y1
xMM_u2 net11 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI3 VDD net11 VDD Dcap_PMOS_n12_X1_Y1
xMM_u1 net9 net11 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DCAP8LVT

.subckt Dcap_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_NMOS_n12_X1_Y1

.subckt Switch_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_NMOS_n12_X1_Y1

.subckt Dcap_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_PMOS_n12_X1_Y1

.subckt Switch_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_PMOS_n12_X1_Y1

.subckt DCAP16LVT 
xMMI4 VSS net11 VSS Dcap_NMOS_n12_X1_Y1
xMM_u2 net5 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI7 VSS net11 VSS Dcap_NMOS_n12_X1_Y1
xMMI3 VDD net5 VDD Dcap_PMOS_n12_X1_Y1
xMM_u1 net11 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 VDD net5 VDD Dcap_PMOS_n12_X1_Y1
.ends DCAP16LVT

.subckt DCAP32LVT 
xMMI39 VSS net11 VSS Dcap_NMOS_n12_X1_Y1
xMM_u2 net5 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI36 VSS net11 VSS Dcap_NMOS_n12_X1_Y1
xMM_u1 net11 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI35 VDD net5 VDD Dcap_PMOS_n12_X1_Y1
xMMI26 VDD net5 VDD Dcap_PMOS_n12_X1_Y1
.ends DCAP32LVT

.subckt CMC_NMOS_S_n12_X1_Y1 B DA G S DB
xM0 DA G S B Switch_NMOS_n12_X1_Y1
xM1 DB G S B Switch_NMOS_n12_X1_Y1
.ends CMC_NMOS_S_n12_X1_Y1

.subckt CMC_PMOS_S_n12_X1_Y1 B DA G S DB
xM0 DA G S B Switch_PMOS_n12_X1_Y1
xM1 DB G S B Switch_PMOS_n12_X1_Y1
.ends CMC_PMOS_S_n12_X1_Y1

.subckt INV_LVT zn i SN SP
xxm0 zn i SN SN Switch_NMOS_n12_X1_Y1
xxm1 zn i SP SP Switch_PMOS_n12_X1_Y1
.ends INV_LVT

.subckt BUFTD16LVT I OE Z
xMMI5_1_M_u4 net25 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5_0_M_u3 net25 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMI7_M_u3 net13 OE net9 VSS Switch_NMOS_n12_X1_Y1
xMM_u7 Z net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI6_M_u3 net13 OE net37 VSS Switch_NMOS_n12_X1_Y1
xMMI5_0_M_u2 net25 net5 net72 VDD Switch_PMOS_n12_X1_Y1
xMMI6_M_u2 net13 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMI7_M_u1 net13 OE VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u6 Z net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5_1_M_u2 net25 net5 net53 VDD Switch_PMOS_n12_X1_Y1
xMMI7_M_u4_MMI6_M_u4 net9 I VSS net37 VSS CMC_NMOS_S_n12_X1_Y1
xMMI5_1_M_u1_MMI5_0_M_u1 net53 I VDD net72 VDD CMC_PMOS_S_n12_X1_Y1
MM_u17_M_u2_MM_u17_M_u3 OE VSS VDD net5 INV_LVT
.ends BUFTD16LVT

.subckt CMC_NMOS_S_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends CMC_NMOS_S_n12_X1_Y1

.subckt CMC_PMOS_S_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends CMC_PMOS_S_n12_X1_Y1
