MACRO CKT_OBS_LEF
  ORIGIN 0 0 ;
  FOREIGN CKT_OBS_LEF 0 0 ;
  SIZE 1.542 BY 3.84 ;
  PIN VOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.294 1.15 1.218 1.19 ;
      LAYER M2 ;
        RECT 0.186 0.79 1.326 0.83 ;
      LAYER M2 ;
        RECT 0.294 1.78 1.218 1.82 ;
      LAYER M2 ;
        RECT 0.186 1.42 1.326 1.46 ;
      LAYER M2 ;
        RECT 0.186 2.95 1.326 2.99 ;
      LAYER M2 ;
        RECT 0.186 2.32 1.326 2.36 ;
      LAYER M3 ;
        RECT 0.618 2.32 0.678 2.99 ;
      LAYER M2 ;
        RECT 0.618 1.78 0.678 1.82 ;
      LAYER M3 ;
        RECT 0.618 1.8 0.678 2.34 ;
    END
  END VOP
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.294 2.59 1.218 2.63 ;
      LAYER M2 ;
        RECT 0.294 1.96 1.218 2 ;
      LAYER M3 ;
        RECT 0.726 1.96 0.786 2.63 ;
    END
  END VIN
  OBS 
  LAYER M1 ;
        RECT 0.186 0.07 0.246 1.64 ;
  LAYER M1 ;
        RECT 0.402 0.07 0.462 1.64 ;
  LAYER M1 ;
        RECT 0.618 0.07 0.678 1.64 ;
  LAYER M1 ;
        RECT 0.834 0.07 0.894 1.64 ;
  LAYER M1 ;
        RECT 1.05 0.07 1.11 1.64 ;
  LAYER M1 ;
        RECT 1.266 0.07 1.326 1.64 ;
  LAYER M1 ;
        RECT 0.294 0.7 0.354 1.82 ;
  LAYER M1 ;
        RECT 0.51 0.7 0.57 1.82 ;
  LAYER M1 ;
        RECT 0.942 0.7 1.002 1.82 ;
  LAYER M1 ;
        RECT 1.158 0.7 1.218 1.82 ;
  LAYER M2 ;
        RECT 0.294 1.15 1.218 1.19 ;
  LAYER M2 ;
        RECT 0.186 0.79 1.326 0.83 ;
  LAYER M2 ;
        RECT 0.294 1.78 1.218 1.82 ;
  LAYER M2 ;
        RECT 0.186 1.42 1.326 1.46 ;
  LAYER M2 ;
        RECT 0.186 0.34 1.326 0.38 ;
  LAYER M2 ;
        RECT 0.186 0.97 1.326 1.01 ;
  LAYER M2 ;
        RECT 0.186 1.6 1.326 1.64 ;
  LAYER M1 ;
        RECT 0.186 2.14 0.246 3.71 ;
  LAYER M1 ;
        RECT 0.402 2.14 0.462 3.71 ;
  LAYER M1 ;
        RECT 0.618 2.14 0.678 3.71 ;
  LAYER M1 ;
        RECT 0.834 2.14 0.894 3.71 ;
  LAYER M1 ;
        RECT 1.05 2.14 1.11 3.71 ;
  LAYER M1 ;
        RECT 1.266 2.14 1.326 3.71 ;
  LAYER M1 ;
        RECT 0.294 2.77 0.354 3.08 ;
  LAYER M1 ;
        RECT 0.294 2.59 0.354 2.72 ;
  LAYER M1 ;
        RECT 0.294 2.14 0.354 2.45 ;
  LAYER M1 ;
        RECT 0.294 1.96 0.354 2.09 ;
  LAYER M1 ;
        RECT 0.51 2.77 0.57 3.08 ;
  LAYER M1 ;
        RECT 0.51 2.59 0.57 2.72 ;
  LAYER M1 ;
        RECT 0.51 2.14 0.57 2.45 ;
  LAYER M1 ;
        RECT 0.51 1.96 0.57 2.09 ;
  LAYER M1 ;
        RECT 0.942 2.77 1.002 3.08 ;
  LAYER M1 ;
        RECT 0.942 2.59 1.002 2.72 ;
  LAYER M1 ;
        RECT 0.942 2.14 1.002 2.45 ;
  LAYER M1 ;
        RECT 0.942 1.96 1.002 2.09 ;
  LAYER M1 ;
        RECT 1.158 2.77 1.218 3.08 ;
  LAYER M1 ;
        RECT 1.158 2.59 1.218 2.72 ;
  LAYER M1 ;
        RECT 1.158 2.14 1.218 2.45 ;
  LAYER M1 ;
        RECT 1.158 1.96 1.218 2.09 ;
  LAYER M2 ;
        RECT 0.186 2.95 1.326 2.99 ;
  LAYER M2 ;
        RECT 0.186 2.32 1.326 2.36 ;
  LAYER M3 ;
        RECT 0.618 2.32 0.678 2.99 ;
  LAYER M2 ;
        RECT 0.294 2.59 1.218 2.63 ;
  LAYER M2 ;
        RECT 0.294 1.96 1.218 2 ;
  LAYER M3 ;
        RECT 0.726 1.96 0.786 2.63 ;
  LAYER M2 ;
        RECT 0.186 3.58 1.326 3.62 ;
  LAYER M2 ;
        RECT 0.186 2.77 1.326 2.81 ;
  LAYER M2 ;
        RECT 0.186 2.14 1.326 2.18 ;
  END 
END CKT_OBS_LEF
