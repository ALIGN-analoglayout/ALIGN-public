MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 12.32 BY 16.884 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.328 16.428 3.36 16.5 ;
      LAYER M2 ;
        RECT 3.308 16.448 3.38 16.48 ;
      LAYER M1 ;
        RECT 9.28 16.428 9.312 16.5 ;
      LAYER M2 ;
        RECT 9.26 16.448 9.332 16.48 ;
      LAYER M2 ;
        RECT 3.344 16.448 9.296 16.48 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
      LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.304 16.596 6.336 16.668 ;
      LAYER M2 ;
        RECT 6.284 16.616 6.356 16.648 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
      LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.832 7.188 8.864 7.26 ;
  LAYER M2 ;
        RECT 8.812 7.208 8.884 7.24 ;
  LAYER M2 ;
        RECT 6.032 7.208 8.848 7.24 ;
  LAYER M1 ;
        RECT 6.016 7.188 6.048 7.26 ;
  LAYER M2 ;
        RECT 5.996 7.208 6.068 7.24 ;
  LAYER M1 ;
        RECT 5.856 10.296 5.888 10.368 ;
  LAYER M2 ;
        RECT 5.836 10.316 5.908 10.348 ;
  LAYER M1 ;
        RECT 5.856 10.164 5.888 10.332 ;
  LAYER M1 ;
        RECT 5.856 10.128 5.888 10.2 ;
  LAYER M2 ;
        RECT 5.836 10.148 5.908 10.18 ;
  LAYER M2 ;
        RECT 5.872 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 8.832 4.08 8.864 4.152 ;
  LAYER M2 ;
        RECT 8.812 4.1 8.884 4.132 ;
  LAYER M2 ;
        RECT 6.032 4.1 8.848 4.132 ;
  LAYER M1 ;
        RECT 6.016 4.08 6.048 4.152 ;
  LAYER M2 ;
        RECT 5.996 4.1 6.068 4.132 ;
  LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
  LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
  LAYER M1 ;
        RECT 6.016 0.42 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 10.164 ;
  LAYER M1 ;
        RECT 5.856 7.188 5.888 7.26 ;
  LAYER M2 ;
        RECT 5.836 7.208 5.908 7.24 ;
  LAYER M2 ;
        RECT 3.056 7.208 5.872 7.24 ;
  LAYER M1 ;
        RECT 3.04 7.188 3.072 7.26 ;
  LAYER M2 ;
        RECT 3.02 7.208 3.092 7.24 ;
  LAYER M1 ;
        RECT 5.856 4.08 5.888 4.152 ;
  LAYER M2 ;
        RECT 5.836 4.1 5.908 4.132 ;
  LAYER M2 ;
        RECT 3.056 4.1 5.872 4.132 ;
  LAYER M1 ;
        RECT 3.04 4.08 3.072 4.152 ;
  LAYER M2 ;
        RECT 3.02 4.1 3.092 4.132 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 7.224 ;
  LAYER M1 ;
        RECT 8.832 10.296 8.864 10.368 ;
  LAYER M2 ;
        RECT 8.812 10.316 8.884 10.348 ;
  LAYER M1 ;
        RECT 8.832 10.164 8.864 10.332 ;
  LAYER M1 ;
        RECT 8.832 10.128 8.864 10.2 ;
  LAYER M2 ;
        RECT 8.812 10.148 8.884 10.18 ;
  LAYER M2 ;
        RECT 8.848 10.148 9.008 10.18 ;
  LAYER M1 ;
        RECT 8.992 10.128 9.024 10.2 ;
  LAYER M2 ;
        RECT 8.972 10.148 9.044 10.18 ;
  LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
  LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
  LAYER M1 ;
        RECT 8.992 0.252 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 10.164 ;
  LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
  LAYER M1 ;
        RECT 2.88 0.972 2.912 1.044 ;
  LAYER M2 ;
        RECT 2.86 0.992 2.932 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 2.896 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 2.88 4.08 2.912 4.152 ;
  LAYER M2 ;
        RECT 2.86 4.1 2.932 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 2.896 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 2.88 7.188 2.912 7.26 ;
  LAYER M2 ;
        RECT 2.86 7.208 2.932 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 2.896 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 2.88 10.296 2.912 10.368 ;
  LAYER M2 ;
        RECT 2.86 10.316 2.932 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 2.896 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 2.88 13.404 2.912 13.476 ;
  LAYER M2 ;
        RECT 2.86 13.424 2.932 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 2.896 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 13.44 ;
  LAYER M1 ;
        RECT 11.808 0.972 11.84 1.044 ;
  LAYER M2 ;
        RECT 11.788 0.992 11.86 1.024 ;
  LAYER M1 ;
        RECT 11.808 0.84 11.84 1.008 ;
  LAYER M1 ;
        RECT 11.808 0.804 11.84 0.876 ;
  LAYER M2 ;
        RECT 11.788 0.824 11.86 0.856 ;
  LAYER M2 ;
        RECT 11.824 0.824 11.984 0.856 ;
  LAYER M1 ;
        RECT 11.968 0.804 12 0.876 ;
  LAYER M2 ;
        RECT 11.948 0.824 12.02 0.856 ;
  LAYER M1 ;
        RECT 11.808 4.08 11.84 4.152 ;
  LAYER M2 ;
        RECT 11.788 4.1 11.86 4.132 ;
  LAYER M1 ;
        RECT 11.808 3.948 11.84 4.116 ;
  LAYER M1 ;
        RECT 11.808 3.912 11.84 3.984 ;
  LAYER M2 ;
        RECT 11.788 3.932 11.86 3.964 ;
  LAYER M2 ;
        RECT 11.824 3.932 11.984 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 11.808 7.188 11.84 7.26 ;
  LAYER M2 ;
        RECT 11.788 7.208 11.86 7.24 ;
  LAYER M1 ;
        RECT 11.808 7.056 11.84 7.224 ;
  LAYER M1 ;
        RECT 11.808 7.02 11.84 7.092 ;
  LAYER M2 ;
        RECT 11.788 7.04 11.86 7.072 ;
  LAYER M2 ;
        RECT 11.824 7.04 11.984 7.072 ;
  LAYER M1 ;
        RECT 11.968 7.02 12 7.092 ;
  LAYER M2 ;
        RECT 11.948 7.04 12.02 7.072 ;
  LAYER M1 ;
        RECT 11.808 10.296 11.84 10.368 ;
  LAYER M2 ;
        RECT 11.788 10.316 11.86 10.348 ;
  LAYER M1 ;
        RECT 11.808 10.164 11.84 10.332 ;
  LAYER M1 ;
        RECT 11.808 10.128 11.84 10.2 ;
  LAYER M2 ;
        RECT 11.788 10.148 11.86 10.18 ;
  LAYER M2 ;
        RECT 11.824 10.148 11.984 10.18 ;
  LAYER M1 ;
        RECT 11.968 10.128 12 10.2 ;
  LAYER M2 ;
        RECT 11.948 10.148 12.02 10.18 ;
  LAYER M1 ;
        RECT 11.808 13.404 11.84 13.476 ;
  LAYER M2 ;
        RECT 11.788 13.424 11.86 13.456 ;
  LAYER M1 ;
        RECT 11.808 13.272 11.84 13.44 ;
  LAYER M1 ;
        RECT 11.808 13.236 11.84 13.308 ;
  LAYER M2 ;
        RECT 11.788 13.256 11.86 13.288 ;
  LAYER M2 ;
        RECT 11.824 13.256 11.984 13.288 ;
  LAYER M1 ;
        RECT 11.968 13.236 12 13.308 ;
  LAYER M2 ;
        RECT 11.948 13.256 12.02 13.288 ;
  LAYER M1 ;
        RECT 11.968 0.048 12 0.12 ;
  LAYER M2 ;
        RECT 11.948 0.068 12.02 0.1 ;
  LAYER M1 ;
        RECT 11.968 0.084 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 13.272 ;
  LAYER M2 ;
        RECT 0.08 0.068 11.984 0.1 ;
  LAYER M1 ;
        RECT 5.856 0.972 5.888 1.044 ;
  LAYER M2 ;
        RECT 5.836 0.992 5.908 1.024 ;
  LAYER M2 ;
        RECT 2.896 0.992 5.872 1.024 ;
  LAYER M1 ;
        RECT 2.88 0.972 2.912 1.044 ;
  LAYER M2 ;
        RECT 2.86 0.992 2.932 1.024 ;
  LAYER M1 ;
        RECT 5.856 13.404 5.888 13.476 ;
  LAYER M2 ;
        RECT 5.836 13.424 5.908 13.456 ;
  LAYER M2 ;
        RECT 2.896 13.424 5.872 13.456 ;
  LAYER M1 ;
        RECT 2.88 13.404 2.912 13.476 ;
  LAYER M2 ;
        RECT 2.86 13.424 2.932 13.456 ;
  LAYER M1 ;
        RECT 8.832 13.404 8.864 13.476 ;
  LAYER M2 ;
        RECT 8.812 13.424 8.884 13.456 ;
  LAYER M2 ;
        RECT 5.872 13.424 8.848 13.456 ;
  LAYER M1 ;
        RECT 5.856 13.404 5.888 13.476 ;
  LAYER M2 ;
        RECT 5.836 13.424 5.908 13.456 ;
  LAYER M1 ;
        RECT 8.832 0.972 8.864 1.044 ;
  LAYER M2 ;
        RECT 8.812 0.992 8.884 1.024 ;
  LAYER M2 ;
        RECT 8.848 0.992 11.824 1.024 ;
  LAYER M1 ;
        RECT 11.808 0.972 11.84 1.044 ;
  LAYER M2 ;
        RECT 11.788 0.992 11.86 1.024 ;
  LAYER M1 ;
        RECT 3.488 12.732 3.52 12.804 ;
  LAYER M2 ;
        RECT 3.468 12.752 3.54 12.784 ;
  LAYER M2 ;
        RECT 3.344 12.752 3.504 12.784 ;
  LAYER M1 ;
        RECT 3.328 12.732 3.36 12.804 ;
  LAYER M2 ;
        RECT 3.308 12.752 3.38 12.784 ;
  LAYER M1 ;
        RECT 3.328 16.428 3.36 16.5 ;
  LAYER M2 ;
        RECT 3.308 16.448 3.38 16.48 ;
  LAYER M1 ;
        RECT 3.328 16.212 3.36 16.464 ;
  LAYER M1 ;
        RECT 3.328 12.768 3.36 16.212 ;
  LAYER M1 ;
        RECT 6.464 9.624 6.496 9.696 ;
  LAYER M2 ;
        RECT 6.444 9.644 6.516 9.676 ;
  LAYER M1 ;
        RECT 6.464 9.66 6.496 9.828 ;
  LAYER M1 ;
        RECT 6.464 9.792 6.496 9.864 ;
  LAYER M2 ;
        RECT 6.444 9.812 6.516 9.844 ;
  LAYER M2 ;
        RECT 6.48 9.812 9.296 9.844 ;
  LAYER M1 ;
        RECT 9.28 9.792 9.312 9.864 ;
  LAYER M2 ;
        RECT 9.26 9.812 9.332 9.844 ;
  LAYER M1 ;
        RECT 6.464 6.516 6.496 6.588 ;
  LAYER M2 ;
        RECT 6.444 6.536 6.516 6.568 ;
  LAYER M1 ;
        RECT 6.464 6.552 6.496 6.72 ;
  LAYER M1 ;
        RECT 6.464 6.684 6.496 6.756 ;
  LAYER M2 ;
        RECT 6.444 6.704 6.516 6.736 ;
  LAYER M2 ;
        RECT 6.48 6.704 9.296 6.736 ;
  LAYER M1 ;
        RECT 9.28 6.684 9.312 6.756 ;
  LAYER M2 ;
        RECT 9.26 6.704 9.332 6.736 ;
  LAYER M1 ;
        RECT 9.28 16.428 9.312 16.5 ;
  LAYER M2 ;
        RECT 9.26 16.448 9.332 16.48 ;
  LAYER M1 ;
        RECT 9.28 16.212 9.312 16.464 ;
  LAYER M1 ;
        RECT 9.28 6.72 9.312 16.212 ;
  LAYER M2 ;
        RECT 3.344 16.448 9.296 16.48 ;
  LAYER M1 ;
        RECT 3.488 9.624 3.52 9.696 ;
  LAYER M2 ;
        RECT 3.468 9.644 3.54 9.676 ;
  LAYER M1 ;
        RECT 3.488 9.66 3.52 9.828 ;
  LAYER M1 ;
        RECT 3.488 9.792 3.52 9.864 ;
  LAYER M2 ;
        RECT 3.468 9.812 3.54 9.844 ;
  LAYER M2 ;
        RECT 3.504 9.812 6.32 9.844 ;
  LAYER M1 ;
        RECT 6.304 9.792 6.336 9.864 ;
  LAYER M2 ;
        RECT 6.284 9.812 6.356 9.844 ;
  LAYER M1 ;
        RECT 3.488 6.516 3.52 6.588 ;
  LAYER M2 ;
        RECT 3.468 6.536 3.54 6.568 ;
  LAYER M1 ;
        RECT 3.488 6.552 3.52 6.72 ;
  LAYER M1 ;
        RECT 3.488 6.684 3.52 6.756 ;
  LAYER M2 ;
        RECT 3.468 6.704 3.54 6.736 ;
  LAYER M2 ;
        RECT 3.504 6.704 6.32 6.736 ;
  LAYER M1 ;
        RECT 6.304 6.684 6.336 6.756 ;
  LAYER M2 ;
        RECT 6.284 6.704 6.356 6.736 ;
  LAYER M1 ;
        RECT 6.464 12.732 6.496 12.804 ;
  LAYER M2 ;
        RECT 6.444 12.752 6.516 12.784 ;
  LAYER M2 ;
        RECT 6.32 12.752 6.48 12.784 ;
  LAYER M1 ;
        RECT 6.304 12.732 6.336 12.804 ;
  LAYER M2 ;
        RECT 6.284 12.752 6.356 12.784 ;
  LAYER M1 ;
        RECT 6.304 16.596 6.336 16.668 ;
  LAYER M2 ;
        RECT 6.284 16.616 6.356 16.648 ;
  LAYER M1 ;
        RECT 6.304 16.212 6.336 16.632 ;
  LAYER M1 ;
        RECT 6.304 6.72 6.336 16.212 ;
  LAYER M1 ;
        RECT 0.512 3.408 0.544 3.48 ;
  LAYER M2 ;
        RECT 0.492 3.428 0.564 3.46 ;
  LAYER M2 ;
        RECT 0.368 3.428 0.528 3.46 ;
  LAYER M1 ;
        RECT 0.352 3.408 0.384 3.48 ;
  LAYER M2 ;
        RECT 0.332 3.428 0.404 3.46 ;
  LAYER M1 ;
        RECT 0.512 6.516 0.544 6.588 ;
  LAYER M2 ;
        RECT 0.492 6.536 0.564 6.568 ;
  LAYER M2 ;
        RECT 0.368 6.536 0.528 6.568 ;
  LAYER M1 ;
        RECT 0.352 6.516 0.384 6.588 ;
  LAYER M2 ;
        RECT 0.332 6.536 0.404 6.568 ;
  LAYER M1 ;
        RECT 0.512 9.624 0.544 9.696 ;
  LAYER M2 ;
        RECT 0.492 9.644 0.564 9.676 ;
  LAYER M2 ;
        RECT 0.368 9.644 0.528 9.676 ;
  LAYER M1 ;
        RECT 0.352 9.624 0.384 9.696 ;
  LAYER M2 ;
        RECT 0.332 9.644 0.404 9.676 ;
  LAYER M1 ;
        RECT 0.512 12.732 0.544 12.804 ;
  LAYER M2 ;
        RECT 0.492 12.752 0.564 12.784 ;
  LAYER M2 ;
        RECT 0.368 12.752 0.528 12.784 ;
  LAYER M1 ;
        RECT 0.352 12.732 0.384 12.804 ;
  LAYER M2 ;
        RECT 0.332 12.752 0.404 12.784 ;
  LAYER M1 ;
        RECT 0.512 15.84 0.544 15.912 ;
  LAYER M2 ;
        RECT 0.492 15.86 0.564 15.892 ;
  LAYER M2 ;
        RECT 0.368 15.86 0.528 15.892 ;
  LAYER M1 ;
        RECT 0.352 15.84 0.384 15.912 ;
  LAYER M2 ;
        RECT 0.332 15.86 0.404 15.892 ;
  LAYER M1 ;
        RECT 0.352 16.764 0.384 16.836 ;
  LAYER M2 ;
        RECT 0.332 16.784 0.404 16.816 ;
  LAYER M1 ;
        RECT 0.352 16.212 0.384 16.8 ;
  LAYER M1 ;
        RECT 0.352 3.444 0.384 16.212 ;
  LAYER M1 ;
        RECT 9.44 3.408 9.472 3.48 ;
  LAYER M2 ;
        RECT 9.42 3.428 9.492 3.46 ;
  LAYER M1 ;
        RECT 9.44 3.444 9.472 3.612 ;
  LAYER M1 ;
        RECT 9.44 3.576 9.472 3.648 ;
  LAYER M2 ;
        RECT 9.42 3.596 9.492 3.628 ;
  LAYER M2 ;
        RECT 9.456 3.596 12.272 3.628 ;
  LAYER M1 ;
        RECT 12.256 3.576 12.288 3.648 ;
  LAYER M2 ;
        RECT 12.236 3.596 12.308 3.628 ;
  LAYER M1 ;
        RECT 9.44 6.516 9.472 6.588 ;
  LAYER M2 ;
        RECT 9.42 6.536 9.492 6.568 ;
  LAYER M1 ;
        RECT 9.44 6.552 9.472 6.72 ;
  LAYER M1 ;
        RECT 9.44 6.684 9.472 6.756 ;
  LAYER M2 ;
        RECT 9.42 6.704 9.492 6.736 ;
  LAYER M2 ;
        RECT 9.456 6.704 12.272 6.736 ;
  LAYER M1 ;
        RECT 12.256 6.684 12.288 6.756 ;
  LAYER M2 ;
        RECT 12.236 6.704 12.308 6.736 ;
  LAYER M1 ;
        RECT 9.44 9.624 9.472 9.696 ;
  LAYER M2 ;
        RECT 9.42 9.644 9.492 9.676 ;
  LAYER M1 ;
        RECT 9.44 9.66 9.472 9.828 ;
  LAYER M1 ;
        RECT 9.44 9.792 9.472 9.864 ;
  LAYER M2 ;
        RECT 9.42 9.812 9.492 9.844 ;
  LAYER M2 ;
        RECT 9.456 9.812 12.272 9.844 ;
  LAYER M1 ;
        RECT 12.256 9.792 12.288 9.864 ;
  LAYER M2 ;
        RECT 12.236 9.812 12.308 9.844 ;
  LAYER M1 ;
        RECT 9.44 12.732 9.472 12.804 ;
  LAYER M2 ;
        RECT 9.42 12.752 9.492 12.784 ;
  LAYER M1 ;
        RECT 9.44 12.768 9.472 12.936 ;
  LAYER M1 ;
        RECT 9.44 12.9 9.472 12.972 ;
  LAYER M2 ;
        RECT 9.42 12.92 9.492 12.952 ;
  LAYER M2 ;
        RECT 9.456 12.92 12.272 12.952 ;
  LAYER M1 ;
        RECT 12.256 12.9 12.288 12.972 ;
  LAYER M2 ;
        RECT 12.236 12.92 12.308 12.952 ;
  LAYER M1 ;
        RECT 9.44 15.84 9.472 15.912 ;
  LAYER M2 ;
        RECT 9.42 15.86 9.492 15.892 ;
  LAYER M1 ;
        RECT 9.44 15.876 9.472 16.044 ;
  LAYER M1 ;
        RECT 9.44 16.008 9.472 16.08 ;
  LAYER M2 ;
        RECT 9.42 16.028 9.492 16.06 ;
  LAYER M2 ;
        RECT 9.456 16.028 12.272 16.06 ;
  LAYER M1 ;
        RECT 12.256 16.008 12.288 16.08 ;
  LAYER M2 ;
        RECT 12.236 16.028 12.308 16.06 ;
  LAYER M1 ;
        RECT 12.256 16.764 12.288 16.836 ;
  LAYER M2 ;
        RECT 12.236 16.784 12.308 16.816 ;
  LAYER M1 ;
        RECT 12.256 16.212 12.288 16.8 ;
  LAYER M1 ;
        RECT 12.256 3.612 12.288 16.212 ;
  LAYER M2 ;
        RECT 0.368 16.784 12.272 16.816 ;
  LAYER M1 ;
        RECT 3.488 3.408 3.52 3.48 ;
  LAYER M2 ;
        RECT 3.468 3.428 3.54 3.46 ;
  LAYER M2 ;
        RECT 0.528 3.428 3.504 3.46 ;
  LAYER M1 ;
        RECT 0.512 3.408 0.544 3.48 ;
  LAYER M2 ;
        RECT 0.492 3.428 0.564 3.46 ;
  LAYER M1 ;
        RECT 3.488 15.84 3.52 15.912 ;
  LAYER M2 ;
        RECT 3.468 15.86 3.54 15.892 ;
  LAYER M2 ;
        RECT 0.528 15.86 3.504 15.892 ;
  LAYER M1 ;
        RECT 0.512 15.84 0.544 15.912 ;
  LAYER M2 ;
        RECT 0.492 15.86 0.564 15.892 ;
  LAYER M1 ;
        RECT 6.464 15.84 6.496 15.912 ;
  LAYER M2 ;
        RECT 6.444 15.86 6.516 15.892 ;
  LAYER M2 ;
        RECT 3.504 15.86 6.48 15.892 ;
  LAYER M1 ;
        RECT 3.488 15.84 3.52 15.912 ;
  LAYER M2 ;
        RECT 3.468 15.86 3.54 15.892 ;
  LAYER M1 ;
        RECT 6.464 3.408 6.496 3.48 ;
  LAYER M2 ;
        RECT 6.444 3.428 6.516 3.46 ;
  LAYER M2 ;
        RECT 6.48 3.428 9.456 3.46 ;
  LAYER M1 ;
        RECT 9.44 3.408 9.472 3.48 ;
  LAYER M2 ;
        RECT 9.42 3.428 9.492 3.46 ;
  LAYER M1 ;
        RECT 0.464 0.924 2.96 3.528 ;
  LAYER M3 ;
        RECT 0.464 0.924 2.96 3.528 ;
  LAYER M2 ;
        RECT 0.464 0.924 2.96 3.528 ;
  LAYER M1 ;
        RECT 0.464 4.032 2.96 6.636 ;
  LAYER M3 ;
        RECT 0.464 4.032 2.96 6.636 ;
  LAYER M2 ;
        RECT 0.464 4.032 2.96 6.636 ;
  LAYER M1 ;
        RECT 0.464 7.14 2.96 9.744 ;
  LAYER M3 ;
        RECT 0.464 7.14 2.96 9.744 ;
  LAYER M2 ;
        RECT 0.464 7.14 2.96 9.744 ;
  LAYER M1 ;
        RECT 0.464 10.248 2.96 12.852 ;
  LAYER M3 ;
        RECT 0.464 10.248 2.96 12.852 ;
  LAYER M2 ;
        RECT 0.464 10.248 2.96 12.852 ;
  LAYER M1 ;
        RECT 0.464 13.356 2.96 15.96 ;
  LAYER M3 ;
        RECT 0.464 13.356 2.96 15.96 ;
  LAYER M2 ;
        RECT 0.464 13.356 2.96 15.96 ;
  LAYER M1 ;
        RECT 3.44 0.924 5.936 3.528 ;
  LAYER M3 ;
        RECT 3.44 0.924 5.936 3.528 ;
  LAYER M2 ;
        RECT 3.44 0.924 5.936 3.528 ;
  LAYER M1 ;
        RECT 3.44 4.032 5.936 6.636 ;
  LAYER M3 ;
        RECT 3.44 4.032 5.936 6.636 ;
  LAYER M2 ;
        RECT 3.44 4.032 5.936 6.636 ;
  LAYER M1 ;
        RECT 3.44 7.14 5.936 9.744 ;
  LAYER M3 ;
        RECT 3.44 7.14 5.936 9.744 ;
  LAYER M2 ;
        RECT 3.44 7.14 5.936 9.744 ;
  LAYER M1 ;
        RECT 3.44 10.248 5.936 12.852 ;
  LAYER M3 ;
        RECT 3.44 10.248 5.936 12.852 ;
  LAYER M2 ;
        RECT 3.44 10.248 5.936 12.852 ;
  LAYER M1 ;
        RECT 3.44 13.356 5.936 15.96 ;
  LAYER M3 ;
        RECT 3.44 13.356 5.936 15.96 ;
  LAYER M2 ;
        RECT 3.44 13.356 5.936 15.96 ;
  LAYER M1 ;
        RECT 6.416 0.924 8.912 3.528 ;
  LAYER M3 ;
        RECT 6.416 0.924 8.912 3.528 ;
  LAYER M2 ;
        RECT 6.416 0.924 8.912 3.528 ;
  LAYER M1 ;
        RECT 6.416 4.032 8.912 6.636 ;
  LAYER M3 ;
        RECT 6.416 4.032 8.912 6.636 ;
  LAYER M2 ;
        RECT 6.416 4.032 8.912 6.636 ;
  LAYER M1 ;
        RECT 6.416 7.14 8.912 9.744 ;
  LAYER M3 ;
        RECT 6.416 7.14 8.912 9.744 ;
  LAYER M2 ;
        RECT 6.416 7.14 8.912 9.744 ;
  LAYER M1 ;
        RECT 6.416 10.248 8.912 12.852 ;
  LAYER M3 ;
        RECT 6.416 10.248 8.912 12.852 ;
  LAYER M2 ;
        RECT 6.416 10.248 8.912 12.852 ;
  LAYER M1 ;
        RECT 6.416 13.356 8.912 15.96 ;
  LAYER M3 ;
        RECT 6.416 13.356 8.912 15.96 ;
  LAYER M2 ;
        RECT 6.416 13.356 8.912 15.96 ;
  LAYER M1 ;
        RECT 9.392 0.924 11.888 3.528 ;
  LAYER M3 ;
        RECT 9.392 0.924 11.888 3.528 ;
  LAYER M2 ;
        RECT 9.392 0.924 11.888 3.528 ;
  LAYER M1 ;
        RECT 9.392 4.032 11.888 6.636 ;
  LAYER M3 ;
        RECT 9.392 4.032 11.888 6.636 ;
  LAYER M2 ;
        RECT 9.392 4.032 11.888 6.636 ;
  LAYER M1 ;
        RECT 9.392 7.14 11.888 9.744 ;
  LAYER M3 ;
        RECT 9.392 7.14 11.888 9.744 ;
  LAYER M2 ;
        RECT 9.392 7.14 11.888 9.744 ;
  LAYER M1 ;
        RECT 9.392 10.248 11.888 12.852 ;
  LAYER M3 ;
        RECT 9.392 10.248 11.888 12.852 ;
  LAYER M2 ;
        RECT 9.392 10.248 11.888 12.852 ;
  LAYER M1 ;
        RECT 9.392 13.356 11.888 15.96 ;
  LAYER M3 ;
        RECT 9.392 13.356 11.888 15.96 ;
  LAYER M2 ;
        RECT 9.392 13.356 11.888 15.96 ;
  END 
END Cap_30fF_Cap_30fF
