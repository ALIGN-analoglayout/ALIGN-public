MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 11.68 BY 18.648 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 18.36 3.136 18.432 ;
      LAYER M2 ;
        RECT 3.084 18.38 3.156 18.412 ;
      LAYER M1 ;
        RECT 8.864 18.36 8.896 18.432 ;
      LAYER M2 ;
        RECT 8.844 18.38 8.916 18.412 ;
      LAYER M2 ;
        RECT 3.12 18.38 8.88 18.412 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
      LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 3.264 6.6 3.296 6.672 ;
  LAYER M2 ;
        RECT 3.244 6.62 3.316 6.652 ;
  LAYER M1 ;
        RECT 3.264 6.468 3.296 6.636 ;
  LAYER M1 ;
        RECT 3.264 6.432 3.296 6.504 ;
  LAYER M2 ;
        RECT 3.244 6.452 3.316 6.484 ;
  LAYER M2 ;
        RECT 3.28 6.452 5.84 6.484 ;
  LAYER M1 ;
        RECT 5.824 6.432 5.856 6.504 ;
  LAYER M2 ;
        RECT 5.804 6.452 5.876 6.484 ;
  LAYER M1 ;
        RECT 6.144 9.54 6.176 9.612 ;
  LAYER M2 ;
        RECT 6.124 9.56 6.196 9.592 ;
  LAYER M2 ;
        RECT 5.84 9.56 6.16 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 9.612 ;
  LAYER M2 ;
        RECT 3.244 9.56 3.316 9.592 ;
  LAYER M1 ;
        RECT 3.264 9.408 3.296 9.576 ;
  LAYER M1 ;
        RECT 3.264 9.372 3.296 9.444 ;
  LAYER M2 ;
        RECT 3.244 9.392 3.316 9.424 ;
  LAYER M2 ;
        RECT 3.28 9.392 5.84 9.424 ;
  LAYER M1 ;
        RECT 5.824 9.372 5.856 9.444 ;
  LAYER M2 ;
        RECT 5.804 9.392 5.876 9.424 ;
  LAYER M1 ;
        RECT 6.144 6.6 6.176 6.672 ;
  LAYER M2 ;
        RECT 6.124 6.62 6.196 6.652 ;
  LAYER M2 ;
        RECT 5.84 6.62 6.16 6.652 ;
  LAYER M1 ;
        RECT 5.824 6.6 5.856 6.672 ;
  LAYER M2 ;
        RECT 5.804 6.62 5.876 6.652 ;
  LAYER M1 ;
        RECT 3.264 12.48 3.296 12.552 ;
  LAYER M2 ;
        RECT 3.244 12.5 3.316 12.532 ;
  LAYER M1 ;
        RECT 3.264 12.348 3.296 12.516 ;
  LAYER M1 ;
        RECT 3.264 12.312 3.296 12.384 ;
  LAYER M2 ;
        RECT 3.244 12.332 3.316 12.364 ;
  LAYER M2 ;
        RECT 3.28 12.332 5.84 12.364 ;
  LAYER M1 ;
        RECT 5.824 12.312 5.856 12.384 ;
  LAYER M2 ;
        RECT 5.804 12.332 5.876 12.364 ;
  LAYER M1 ;
        RECT 6.144 3.66 6.176 3.732 ;
  LAYER M2 ;
        RECT 6.124 3.68 6.196 3.712 ;
  LAYER M2 ;
        RECT 5.84 3.68 6.16 3.712 ;
  LAYER M1 ;
        RECT 5.824 3.66 5.856 3.732 ;
  LAYER M2 ;
        RECT 5.804 3.68 5.876 3.712 ;
  LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
  LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
  LAYER M1 ;
        RECT 5.824 0.252 5.856 0.42 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 12.348 ;
  LAYER M1 ;
        RECT 0.384 0.72 0.416 0.792 ;
  LAYER M2 ;
        RECT 0.364 0.74 0.436 0.772 ;
  LAYER M1 ;
        RECT 0.384 0.588 0.416 0.756 ;
  LAYER M1 ;
        RECT 0.384 0.552 0.416 0.624 ;
  LAYER M2 ;
        RECT 0.364 0.572 0.436 0.604 ;
  LAYER M2 ;
        RECT 0.4 0.572 2.96 0.604 ;
  LAYER M1 ;
        RECT 2.944 0.552 2.976 0.624 ;
  LAYER M2 ;
        RECT 2.924 0.572 2.996 0.604 ;
  LAYER M1 ;
        RECT 0.384 3.66 0.416 3.732 ;
  LAYER M2 ;
        RECT 0.364 3.68 0.436 3.712 ;
  LAYER M1 ;
        RECT 0.384 3.528 0.416 3.696 ;
  LAYER M1 ;
        RECT 0.384 3.492 0.416 3.564 ;
  LAYER M2 ;
        RECT 0.364 3.512 0.436 3.544 ;
  LAYER M2 ;
        RECT 0.4 3.512 2.96 3.544 ;
  LAYER M1 ;
        RECT 2.944 3.492 2.976 3.564 ;
  LAYER M2 ;
        RECT 2.924 3.512 2.996 3.544 ;
  LAYER M1 ;
        RECT 0.384 6.6 0.416 6.672 ;
  LAYER M2 ;
        RECT 0.364 6.62 0.436 6.652 ;
  LAYER M1 ;
        RECT 0.384 6.468 0.416 6.636 ;
  LAYER M1 ;
        RECT 0.384 6.432 0.416 6.504 ;
  LAYER M2 ;
        RECT 0.364 6.452 0.436 6.484 ;
  LAYER M2 ;
        RECT 0.4 6.452 2.96 6.484 ;
  LAYER M1 ;
        RECT 2.944 6.432 2.976 6.504 ;
  LAYER M2 ;
        RECT 2.924 6.452 2.996 6.484 ;
  LAYER M1 ;
        RECT 0.384 9.54 0.416 9.612 ;
  LAYER M2 ;
        RECT 0.364 9.56 0.436 9.592 ;
  LAYER M1 ;
        RECT 0.384 9.408 0.416 9.576 ;
  LAYER M1 ;
        RECT 0.384 9.372 0.416 9.444 ;
  LAYER M2 ;
        RECT 0.364 9.392 0.436 9.424 ;
  LAYER M2 ;
        RECT 0.4 9.392 2.96 9.424 ;
  LAYER M1 ;
        RECT 2.944 9.372 2.976 9.444 ;
  LAYER M2 ;
        RECT 2.924 9.392 2.996 9.424 ;
  LAYER M1 ;
        RECT 0.384 12.48 0.416 12.552 ;
  LAYER M2 ;
        RECT 0.364 12.5 0.436 12.532 ;
  LAYER M1 ;
        RECT 0.384 12.348 0.416 12.516 ;
  LAYER M1 ;
        RECT 0.384 12.312 0.416 12.384 ;
  LAYER M2 ;
        RECT 0.364 12.332 0.436 12.364 ;
  LAYER M2 ;
        RECT 0.4 12.332 2.96 12.364 ;
  LAYER M1 ;
        RECT 2.944 12.312 2.976 12.384 ;
  LAYER M2 ;
        RECT 2.924 12.332 2.996 12.364 ;
  LAYER M1 ;
        RECT 0.384 15.42 0.416 15.492 ;
  LAYER M2 ;
        RECT 0.364 15.44 0.436 15.472 ;
  LAYER M1 ;
        RECT 0.384 15.288 0.416 15.456 ;
  LAYER M1 ;
        RECT 0.384 15.252 0.416 15.324 ;
  LAYER M2 ;
        RECT 0.364 15.272 0.436 15.304 ;
  LAYER M2 ;
        RECT 0.4 15.272 2.96 15.304 ;
  LAYER M1 ;
        RECT 2.944 15.252 2.976 15.324 ;
  LAYER M2 ;
        RECT 2.924 15.272 2.996 15.304 ;
  LAYER M1 ;
        RECT 3.264 0.72 3.296 0.792 ;
  LAYER M2 ;
        RECT 3.244 0.74 3.316 0.772 ;
  LAYER M2 ;
        RECT 2.96 0.74 3.28 0.772 ;
  LAYER M1 ;
        RECT 2.944 0.72 2.976 0.792 ;
  LAYER M2 ;
        RECT 2.924 0.74 2.996 0.772 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 3.732 ;
  LAYER M2 ;
        RECT 3.244 3.68 3.316 3.712 ;
  LAYER M2 ;
        RECT 2.96 3.68 3.28 3.712 ;
  LAYER M1 ;
        RECT 2.944 3.66 2.976 3.732 ;
  LAYER M2 ;
        RECT 2.924 3.68 2.996 3.712 ;
  LAYER M1 ;
        RECT 3.264 15.42 3.296 15.492 ;
  LAYER M2 ;
        RECT 3.244 15.44 3.316 15.472 ;
  LAYER M2 ;
        RECT 2.96 15.44 3.28 15.472 ;
  LAYER M1 ;
        RECT 2.944 15.42 2.976 15.492 ;
  LAYER M2 ;
        RECT 2.924 15.44 2.996 15.472 ;
  LAYER M1 ;
        RECT 2.944 0.048 2.976 0.12 ;
  LAYER M2 ;
        RECT 2.924 0.068 2.996 0.1 ;
  LAYER M1 ;
        RECT 2.944 0.084 2.976 0.42 ;
  LAYER M1 ;
        RECT 2.944 0.42 2.976 15.456 ;
  LAYER M1 ;
        RECT 6.144 0.72 6.176 0.792 ;
  LAYER M2 ;
        RECT 6.124 0.74 6.196 0.772 ;
  LAYER M1 ;
        RECT 6.144 0.588 6.176 0.756 ;
  LAYER M1 ;
        RECT 6.144 0.552 6.176 0.624 ;
  LAYER M2 ;
        RECT 6.124 0.572 6.196 0.604 ;
  LAYER M2 ;
        RECT 6.16 0.572 8.72 0.604 ;
  LAYER M1 ;
        RECT 8.704 0.552 8.736 0.624 ;
  LAYER M2 ;
        RECT 8.684 0.572 8.756 0.604 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 12.552 ;
  LAYER M2 ;
        RECT 6.124 12.5 6.196 12.532 ;
  LAYER M1 ;
        RECT 6.144 12.348 6.176 12.516 ;
  LAYER M1 ;
        RECT 6.144 12.312 6.176 12.384 ;
  LAYER M2 ;
        RECT 6.124 12.332 6.196 12.364 ;
  LAYER M2 ;
        RECT 6.16 12.332 8.72 12.364 ;
  LAYER M1 ;
        RECT 8.704 12.312 8.736 12.384 ;
  LAYER M2 ;
        RECT 8.684 12.332 8.756 12.364 ;
  LAYER M1 ;
        RECT 6.144 15.42 6.176 15.492 ;
  LAYER M2 ;
        RECT 6.124 15.44 6.196 15.472 ;
  LAYER M1 ;
        RECT 6.144 15.288 6.176 15.456 ;
  LAYER M1 ;
        RECT 6.144 15.252 6.176 15.324 ;
  LAYER M2 ;
        RECT 6.124 15.272 6.196 15.304 ;
  LAYER M2 ;
        RECT 6.16 15.272 8.72 15.304 ;
  LAYER M1 ;
        RECT 8.704 15.252 8.736 15.324 ;
  LAYER M2 ;
        RECT 8.684 15.272 8.756 15.304 ;
  LAYER M1 ;
        RECT 9.024 0.72 9.056 0.792 ;
  LAYER M2 ;
        RECT 9.004 0.74 9.076 0.772 ;
  LAYER M2 ;
        RECT 8.72 0.74 9.04 0.772 ;
  LAYER M1 ;
        RECT 8.704 0.72 8.736 0.792 ;
  LAYER M2 ;
        RECT 8.684 0.74 8.756 0.772 ;
  LAYER M1 ;
        RECT 9.024 3.66 9.056 3.732 ;
  LAYER M2 ;
        RECT 9.004 3.68 9.076 3.712 ;
  LAYER M2 ;
        RECT 8.72 3.68 9.04 3.712 ;
  LAYER M1 ;
        RECT 8.704 3.66 8.736 3.732 ;
  LAYER M2 ;
        RECT 8.684 3.68 8.756 3.712 ;
  LAYER M1 ;
        RECT 9.024 6.6 9.056 6.672 ;
  LAYER M2 ;
        RECT 9.004 6.62 9.076 6.652 ;
  LAYER M2 ;
        RECT 8.72 6.62 9.04 6.652 ;
  LAYER M1 ;
        RECT 8.704 6.6 8.736 6.672 ;
  LAYER M2 ;
        RECT 8.684 6.62 8.756 6.652 ;
  LAYER M1 ;
        RECT 9.024 9.54 9.056 9.612 ;
  LAYER M2 ;
        RECT 9.004 9.56 9.076 9.592 ;
  LAYER M2 ;
        RECT 8.72 9.56 9.04 9.592 ;
  LAYER M1 ;
        RECT 8.704 9.54 8.736 9.612 ;
  LAYER M2 ;
        RECT 8.684 9.56 8.756 9.592 ;
  LAYER M1 ;
        RECT 9.024 12.48 9.056 12.552 ;
  LAYER M2 ;
        RECT 9.004 12.5 9.076 12.532 ;
  LAYER M2 ;
        RECT 8.72 12.5 9.04 12.532 ;
  LAYER M1 ;
        RECT 8.704 12.48 8.736 12.552 ;
  LAYER M2 ;
        RECT 8.684 12.5 8.756 12.532 ;
  LAYER M1 ;
        RECT 9.024 15.42 9.056 15.492 ;
  LAYER M2 ;
        RECT 9.004 15.44 9.076 15.472 ;
  LAYER M2 ;
        RECT 8.72 15.44 9.04 15.472 ;
  LAYER M1 ;
        RECT 8.704 15.42 8.736 15.492 ;
  LAYER M2 ;
        RECT 8.684 15.44 8.756 15.472 ;
  LAYER M1 ;
        RECT 8.704 0.048 8.736 0.12 ;
  LAYER M2 ;
        RECT 8.684 0.068 8.756 0.1 ;
  LAYER M1 ;
        RECT 8.704 0.084 8.736 0.42 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 15.456 ;
  LAYER M2 ;
        RECT 2.96 0.068 8.72 0.1 ;
  LAYER M1 ;
        RECT 5.664 9.036 5.696 9.108 ;
  LAYER M2 ;
        RECT 5.644 9.056 5.716 9.088 ;
  LAYER M2 ;
        RECT 3.12 9.056 5.68 9.088 ;
  LAYER M1 ;
        RECT 3.104 9.036 3.136 9.108 ;
  LAYER M2 ;
        RECT 3.084 9.056 3.156 9.088 ;
  LAYER M1 ;
        RECT 5.664 11.976 5.696 12.048 ;
  LAYER M2 ;
        RECT 5.644 11.996 5.716 12.028 ;
  LAYER M2 ;
        RECT 3.12 11.996 5.68 12.028 ;
  LAYER M1 ;
        RECT 3.104 11.976 3.136 12.048 ;
  LAYER M2 ;
        RECT 3.084 11.996 3.156 12.028 ;
  LAYER M1 ;
        RECT 5.664 14.916 5.696 14.988 ;
  LAYER M2 ;
        RECT 5.644 14.936 5.716 14.968 ;
  LAYER M2 ;
        RECT 3.12 14.936 5.68 14.968 ;
  LAYER M1 ;
        RECT 3.104 14.916 3.136 14.988 ;
  LAYER M2 ;
        RECT 3.084 14.936 3.156 14.968 ;
  LAYER M1 ;
        RECT 3.104 18.36 3.136 18.432 ;
  LAYER M2 ;
        RECT 3.084 18.38 3.156 18.412 ;
  LAYER M1 ;
        RECT 3.104 18.228 3.136 18.396 ;
  LAYER M1 ;
        RECT 3.104 9.072 3.136 18.228 ;
  LAYER M1 ;
        RECT 8.544 11.976 8.576 12.048 ;
  LAYER M2 ;
        RECT 8.524 11.996 8.596 12.028 ;
  LAYER M1 ;
        RECT 8.544 12.012 8.576 12.18 ;
  LAYER M1 ;
        RECT 8.544 12.144 8.576 12.216 ;
  LAYER M2 ;
        RECT 8.524 12.164 8.596 12.196 ;
  LAYER M2 ;
        RECT 8.56 12.164 8.88 12.196 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M1 ;
        RECT 8.544 9.036 8.576 9.108 ;
  LAYER M2 ;
        RECT 8.524 9.056 8.596 9.088 ;
  LAYER M1 ;
        RECT 8.544 9.072 8.576 9.24 ;
  LAYER M1 ;
        RECT 8.544 9.204 8.576 9.276 ;
  LAYER M2 ;
        RECT 8.524 9.224 8.596 9.256 ;
  LAYER M2 ;
        RECT 8.56 9.224 8.88 9.256 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M1 ;
        RECT 8.544 6.096 8.576 6.168 ;
  LAYER M2 ;
        RECT 8.524 6.116 8.596 6.148 ;
  LAYER M1 ;
        RECT 8.544 6.132 8.576 6.3 ;
  LAYER M1 ;
        RECT 8.544 6.264 8.576 6.336 ;
  LAYER M2 ;
        RECT 8.524 6.284 8.596 6.316 ;
  LAYER M2 ;
        RECT 8.56 6.284 8.88 6.316 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M1 ;
        RECT 8.864 18.36 8.896 18.432 ;
  LAYER M2 ;
        RECT 8.844 18.38 8.916 18.412 ;
  LAYER M1 ;
        RECT 8.864 18.228 8.896 18.396 ;
  LAYER M1 ;
        RECT 8.864 6.3 8.896 18.228 ;
  LAYER M2 ;
        RECT 3.12 18.38 8.88 18.412 ;
  LAYER M1 ;
        RECT 2.784 3.156 2.816 3.228 ;
  LAYER M2 ;
        RECT 2.764 3.176 2.836 3.208 ;
  LAYER M2 ;
        RECT 0.08 3.176 2.8 3.208 ;
  LAYER M1 ;
        RECT 0.064 3.156 0.096 3.228 ;
  LAYER M2 ;
        RECT 0.044 3.176 0.116 3.208 ;
  LAYER M1 ;
        RECT 2.784 6.096 2.816 6.168 ;
  LAYER M2 ;
        RECT 2.764 6.116 2.836 6.148 ;
  LAYER M2 ;
        RECT 0.08 6.116 2.8 6.148 ;
  LAYER M1 ;
        RECT 0.064 6.096 0.096 6.168 ;
  LAYER M2 ;
        RECT 0.044 6.116 0.116 6.148 ;
  LAYER M1 ;
        RECT 2.784 9.036 2.816 9.108 ;
  LAYER M2 ;
        RECT 2.764 9.056 2.836 9.088 ;
  LAYER M2 ;
        RECT 0.08 9.056 2.8 9.088 ;
  LAYER M1 ;
        RECT 0.064 9.036 0.096 9.108 ;
  LAYER M2 ;
        RECT 0.044 9.056 0.116 9.088 ;
  LAYER M1 ;
        RECT 2.784 11.976 2.816 12.048 ;
  LAYER M2 ;
        RECT 2.764 11.996 2.836 12.028 ;
  LAYER M2 ;
        RECT 0.08 11.996 2.8 12.028 ;
  LAYER M1 ;
        RECT 0.064 11.976 0.096 12.048 ;
  LAYER M2 ;
        RECT 0.044 11.996 0.116 12.028 ;
  LAYER M1 ;
        RECT 2.784 14.916 2.816 14.988 ;
  LAYER M2 ;
        RECT 2.764 14.936 2.836 14.968 ;
  LAYER M2 ;
        RECT 0.08 14.936 2.8 14.968 ;
  LAYER M1 ;
        RECT 0.064 14.916 0.096 14.988 ;
  LAYER M2 ;
        RECT 0.044 14.936 0.116 14.968 ;
  LAYER M1 ;
        RECT 2.784 17.856 2.816 17.928 ;
  LAYER M2 ;
        RECT 2.764 17.876 2.836 17.908 ;
  LAYER M2 ;
        RECT 0.08 17.876 2.8 17.908 ;
  LAYER M1 ;
        RECT 0.064 17.856 0.096 17.928 ;
  LAYER M2 ;
        RECT 0.044 17.876 0.116 17.908 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M1 ;
        RECT 0.064 18.228 0.096 18.564 ;
  LAYER M1 ;
        RECT 0.064 3.192 0.096 18.228 ;
  LAYER M1 ;
        RECT 11.424 3.156 11.456 3.228 ;
  LAYER M2 ;
        RECT 11.404 3.176 11.476 3.208 ;
  LAYER M1 ;
        RECT 11.424 3.192 11.456 3.36 ;
  LAYER M1 ;
        RECT 11.424 3.324 11.456 3.396 ;
  LAYER M2 ;
        RECT 11.404 3.344 11.476 3.376 ;
  LAYER M2 ;
        RECT 11.44 3.344 11.6 3.376 ;
  LAYER M1 ;
        RECT 11.584 3.324 11.616 3.396 ;
  LAYER M2 ;
        RECT 11.564 3.344 11.636 3.376 ;
  LAYER M1 ;
        RECT 11.424 6.096 11.456 6.168 ;
  LAYER M2 ;
        RECT 11.404 6.116 11.476 6.148 ;
  LAYER M1 ;
        RECT 11.424 6.132 11.456 6.3 ;
  LAYER M1 ;
        RECT 11.424 6.264 11.456 6.336 ;
  LAYER M2 ;
        RECT 11.404 6.284 11.476 6.316 ;
  LAYER M2 ;
        RECT 11.44 6.284 11.6 6.316 ;
  LAYER M1 ;
        RECT 11.584 6.264 11.616 6.336 ;
  LAYER M2 ;
        RECT 11.564 6.284 11.636 6.316 ;
  LAYER M1 ;
        RECT 11.424 9.036 11.456 9.108 ;
  LAYER M2 ;
        RECT 11.404 9.056 11.476 9.088 ;
  LAYER M1 ;
        RECT 11.424 9.072 11.456 9.24 ;
  LAYER M1 ;
        RECT 11.424 9.204 11.456 9.276 ;
  LAYER M2 ;
        RECT 11.404 9.224 11.476 9.256 ;
  LAYER M2 ;
        RECT 11.44 9.224 11.6 9.256 ;
  LAYER M1 ;
        RECT 11.584 9.204 11.616 9.276 ;
  LAYER M2 ;
        RECT 11.564 9.224 11.636 9.256 ;
  LAYER M1 ;
        RECT 11.424 11.976 11.456 12.048 ;
  LAYER M2 ;
        RECT 11.404 11.996 11.476 12.028 ;
  LAYER M1 ;
        RECT 11.424 12.012 11.456 12.18 ;
  LAYER M1 ;
        RECT 11.424 12.144 11.456 12.216 ;
  LAYER M2 ;
        RECT 11.404 12.164 11.476 12.196 ;
  LAYER M2 ;
        RECT 11.44 12.164 11.6 12.196 ;
  LAYER M1 ;
        RECT 11.584 12.144 11.616 12.216 ;
  LAYER M2 ;
        RECT 11.564 12.164 11.636 12.196 ;
  LAYER M1 ;
        RECT 11.424 14.916 11.456 14.988 ;
  LAYER M2 ;
        RECT 11.404 14.936 11.476 14.968 ;
  LAYER M1 ;
        RECT 11.424 14.952 11.456 15.12 ;
  LAYER M1 ;
        RECT 11.424 15.084 11.456 15.156 ;
  LAYER M2 ;
        RECT 11.404 15.104 11.476 15.136 ;
  LAYER M2 ;
        RECT 11.44 15.104 11.6 15.136 ;
  LAYER M1 ;
        RECT 11.584 15.084 11.616 15.156 ;
  LAYER M2 ;
        RECT 11.564 15.104 11.636 15.136 ;
  LAYER M1 ;
        RECT 11.424 17.856 11.456 17.928 ;
  LAYER M2 ;
        RECT 11.404 17.876 11.476 17.908 ;
  LAYER M1 ;
        RECT 11.424 17.892 11.456 18.06 ;
  LAYER M1 ;
        RECT 11.424 18.024 11.456 18.096 ;
  LAYER M2 ;
        RECT 11.404 18.044 11.476 18.076 ;
  LAYER M2 ;
        RECT 11.44 18.044 11.6 18.076 ;
  LAYER M1 ;
        RECT 11.584 18.024 11.616 18.096 ;
  LAYER M2 ;
        RECT 11.564 18.044 11.636 18.076 ;
  LAYER M1 ;
        RECT 11.584 18.528 11.616 18.6 ;
  LAYER M2 ;
        RECT 11.564 18.548 11.636 18.58 ;
  LAYER M1 ;
        RECT 11.584 18.228 11.616 18.564 ;
  LAYER M1 ;
        RECT 11.584 3.36 11.616 18.228 ;
  LAYER M2 ;
        RECT 0.08 18.548 11.6 18.58 ;
  LAYER M1 ;
        RECT 5.664 3.156 5.696 3.228 ;
  LAYER M2 ;
        RECT 5.644 3.176 5.716 3.208 ;
  LAYER M2 ;
        RECT 2.8 3.176 5.68 3.208 ;
  LAYER M1 ;
        RECT 2.784 3.156 2.816 3.228 ;
  LAYER M2 ;
        RECT 2.764 3.176 2.836 3.208 ;
  LAYER M1 ;
        RECT 5.664 6.096 5.696 6.168 ;
  LAYER M2 ;
        RECT 5.644 6.116 5.716 6.148 ;
  LAYER M2 ;
        RECT 2.8 6.116 5.68 6.148 ;
  LAYER M1 ;
        RECT 2.784 6.096 2.816 6.168 ;
  LAYER M2 ;
        RECT 2.764 6.116 2.836 6.148 ;
  LAYER M1 ;
        RECT 5.664 17.856 5.696 17.928 ;
  LAYER M2 ;
        RECT 5.644 17.876 5.716 17.908 ;
  LAYER M2 ;
        RECT 2.8 17.876 5.68 17.908 ;
  LAYER M1 ;
        RECT 2.784 17.856 2.816 17.928 ;
  LAYER M2 ;
        RECT 2.764 17.876 2.836 17.908 ;
  LAYER M1 ;
        RECT 8.544 17.856 8.576 17.928 ;
  LAYER M2 ;
        RECT 8.524 17.876 8.596 17.908 ;
  LAYER M2 ;
        RECT 5.68 17.876 8.56 17.908 ;
  LAYER M1 ;
        RECT 5.664 17.856 5.696 17.928 ;
  LAYER M2 ;
        RECT 5.644 17.876 5.716 17.908 ;
  LAYER M1 ;
        RECT 8.544 14.916 8.576 14.988 ;
  LAYER M2 ;
        RECT 8.524 14.936 8.596 14.968 ;
  LAYER M1 ;
        RECT 8.544 14.952 8.576 17.892 ;
  LAYER M1 ;
        RECT 8.544 17.856 8.576 17.928 ;
  LAYER M2 ;
        RECT 8.524 17.876 8.596 17.908 ;
  LAYER M1 ;
        RECT 8.544 3.156 8.576 3.228 ;
  LAYER M2 ;
        RECT 8.524 3.176 8.596 3.208 ;
  LAYER M2 ;
        RECT 8.56 3.176 11.44 3.208 ;
  LAYER M1 ;
        RECT 11.424 3.156 11.456 3.228 ;
  LAYER M2 ;
        RECT 11.404 3.176 11.476 3.208 ;
  LAYER M1 ;
        RECT 0.384 0.72 0.416 3.228 ;
  LAYER M1 ;
        RECT 0.448 0.72 0.48 3.228 ;
  LAYER M1 ;
        RECT 0.512 0.72 0.544 3.228 ;
  LAYER M1 ;
        RECT 0.576 0.72 0.608 3.228 ;
  LAYER M1 ;
        RECT 0.64 0.72 0.672 3.228 ;
  LAYER M1 ;
        RECT 0.704 0.72 0.736 3.228 ;
  LAYER M1 ;
        RECT 0.768 0.72 0.8 3.228 ;
  LAYER M1 ;
        RECT 0.832 0.72 0.864 3.228 ;
  LAYER M1 ;
        RECT 0.896 0.72 0.928 3.228 ;
  LAYER M1 ;
        RECT 0.96 0.72 0.992 3.228 ;
  LAYER M1 ;
        RECT 1.024 0.72 1.056 3.228 ;
  LAYER M1 ;
        RECT 1.088 0.72 1.12 3.228 ;
  LAYER M1 ;
        RECT 1.152 0.72 1.184 3.228 ;
  LAYER M1 ;
        RECT 1.216 0.72 1.248 3.228 ;
  LAYER M1 ;
        RECT 1.28 0.72 1.312 3.228 ;
  LAYER M1 ;
        RECT 1.344 0.72 1.376 3.228 ;
  LAYER M1 ;
        RECT 1.408 0.72 1.44 3.228 ;
  LAYER M1 ;
        RECT 1.472 0.72 1.504 3.228 ;
  LAYER M1 ;
        RECT 1.536 0.72 1.568 3.228 ;
  LAYER M1 ;
        RECT 1.6 0.72 1.632 3.228 ;
  LAYER M1 ;
        RECT 1.664 0.72 1.696 3.228 ;
  LAYER M1 ;
        RECT 1.728 0.72 1.76 3.228 ;
  LAYER M1 ;
        RECT 1.792 0.72 1.824 3.228 ;
  LAYER M1 ;
        RECT 1.856 0.72 1.888 3.228 ;
  LAYER M1 ;
        RECT 1.92 0.72 1.952 3.228 ;
  LAYER M1 ;
        RECT 1.984 0.72 2.016 3.228 ;
  LAYER M1 ;
        RECT 2.048 0.72 2.08 3.228 ;
  LAYER M1 ;
        RECT 2.112 0.72 2.144 3.228 ;
  LAYER M1 ;
        RECT 2.176 0.72 2.208 3.228 ;
  LAYER M1 ;
        RECT 2.24 0.72 2.272 3.228 ;
  LAYER M1 ;
        RECT 2.304 0.72 2.336 3.228 ;
  LAYER M1 ;
        RECT 2.368 0.72 2.4 3.228 ;
  LAYER M1 ;
        RECT 2.432 0.72 2.464 3.228 ;
  LAYER M1 ;
        RECT 2.496 0.72 2.528 3.228 ;
  LAYER M1 ;
        RECT 2.56 0.72 2.592 3.228 ;
  LAYER M1 ;
        RECT 2.624 0.72 2.656 3.228 ;
  LAYER M1 ;
        RECT 2.688 0.72 2.72 3.228 ;
  LAYER M2 ;
        RECT 0.364 0.804 2.836 0.836 ;
  LAYER M2 ;
        RECT 0.364 0.868 2.836 0.9 ;
  LAYER M2 ;
        RECT 0.364 0.932 2.836 0.964 ;
  LAYER M2 ;
        RECT 0.364 0.996 2.836 1.028 ;
  LAYER M2 ;
        RECT 0.364 1.06 2.836 1.092 ;
  LAYER M2 ;
        RECT 0.364 1.124 2.836 1.156 ;
  LAYER M2 ;
        RECT 0.364 1.188 2.836 1.22 ;
  LAYER M2 ;
        RECT 0.364 1.252 2.836 1.284 ;
  LAYER M2 ;
        RECT 0.364 1.316 2.836 1.348 ;
  LAYER M2 ;
        RECT 0.364 1.38 2.836 1.412 ;
  LAYER M2 ;
        RECT 0.364 1.444 2.836 1.476 ;
  LAYER M2 ;
        RECT 0.364 1.508 2.836 1.54 ;
  LAYER M2 ;
        RECT 0.364 1.572 2.836 1.604 ;
  LAYER M2 ;
        RECT 0.364 1.636 2.836 1.668 ;
  LAYER M2 ;
        RECT 0.364 1.7 2.836 1.732 ;
  LAYER M2 ;
        RECT 0.364 1.764 2.836 1.796 ;
  LAYER M2 ;
        RECT 0.364 1.828 2.836 1.86 ;
  LAYER M2 ;
        RECT 0.364 1.892 2.836 1.924 ;
  LAYER M2 ;
        RECT 0.364 1.956 2.836 1.988 ;
  LAYER M2 ;
        RECT 0.364 2.02 2.836 2.052 ;
  LAYER M2 ;
        RECT 0.364 2.084 2.836 2.116 ;
  LAYER M2 ;
        RECT 0.364 2.148 2.836 2.18 ;
  LAYER M2 ;
        RECT 0.364 2.212 2.836 2.244 ;
  LAYER M2 ;
        RECT 0.364 2.276 2.836 2.308 ;
  LAYER M2 ;
        RECT 0.364 2.34 2.836 2.372 ;
  LAYER M2 ;
        RECT 0.364 2.404 2.836 2.436 ;
  LAYER M2 ;
        RECT 0.364 2.468 2.836 2.5 ;
  LAYER M2 ;
        RECT 0.364 2.532 2.836 2.564 ;
  LAYER M2 ;
        RECT 0.364 2.596 2.836 2.628 ;
  LAYER M2 ;
        RECT 0.364 2.66 2.836 2.692 ;
  LAYER M2 ;
        RECT 0.364 2.724 2.836 2.756 ;
  LAYER M2 ;
        RECT 0.364 2.788 2.836 2.82 ;
  LAYER M2 ;
        RECT 0.364 2.852 2.836 2.884 ;
  LAYER M2 ;
        RECT 0.364 2.916 2.836 2.948 ;
  LAYER M2 ;
        RECT 0.364 2.98 2.836 3.012 ;
  LAYER M2 ;
        RECT 0.364 3.044 2.836 3.076 ;
  LAYER M3 ;
        RECT 0.384 0.72 0.416 3.228 ;
  LAYER M3 ;
        RECT 0.448 0.72 0.48 3.228 ;
  LAYER M3 ;
        RECT 0.512 0.72 0.544 3.228 ;
  LAYER M3 ;
        RECT 0.576 0.72 0.608 3.228 ;
  LAYER M3 ;
        RECT 0.64 0.72 0.672 3.228 ;
  LAYER M3 ;
        RECT 0.704 0.72 0.736 3.228 ;
  LAYER M3 ;
        RECT 0.768 0.72 0.8 3.228 ;
  LAYER M3 ;
        RECT 0.832 0.72 0.864 3.228 ;
  LAYER M3 ;
        RECT 0.896 0.72 0.928 3.228 ;
  LAYER M3 ;
        RECT 0.96 0.72 0.992 3.228 ;
  LAYER M3 ;
        RECT 1.024 0.72 1.056 3.228 ;
  LAYER M3 ;
        RECT 1.088 0.72 1.12 3.228 ;
  LAYER M3 ;
        RECT 1.152 0.72 1.184 3.228 ;
  LAYER M3 ;
        RECT 1.216 0.72 1.248 3.228 ;
  LAYER M3 ;
        RECT 1.28 0.72 1.312 3.228 ;
  LAYER M3 ;
        RECT 1.344 0.72 1.376 3.228 ;
  LAYER M3 ;
        RECT 1.408 0.72 1.44 3.228 ;
  LAYER M3 ;
        RECT 1.472 0.72 1.504 3.228 ;
  LAYER M3 ;
        RECT 1.536 0.72 1.568 3.228 ;
  LAYER M3 ;
        RECT 1.6 0.72 1.632 3.228 ;
  LAYER M3 ;
        RECT 1.664 0.72 1.696 3.228 ;
  LAYER M3 ;
        RECT 1.728 0.72 1.76 3.228 ;
  LAYER M3 ;
        RECT 1.792 0.72 1.824 3.228 ;
  LAYER M3 ;
        RECT 1.856 0.72 1.888 3.228 ;
  LAYER M3 ;
        RECT 1.92 0.72 1.952 3.228 ;
  LAYER M3 ;
        RECT 1.984 0.72 2.016 3.228 ;
  LAYER M3 ;
        RECT 2.048 0.72 2.08 3.228 ;
  LAYER M3 ;
        RECT 2.112 0.72 2.144 3.228 ;
  LAYER M3 ;
        RECT 2.176 0.72 2.208 3.228 ;
  LAYER M3 ;
        RECT 2.24 0.72 2.272 3.228 ;
  LAYER M3 ;
        RECT 2.304 0.72 2.336 3.228 ;
  LAYER M3 ;
        RECT 2.368 0.72 2.4 3.228 ;
  LAYER M3 ;
        RECT 2.432 0.72 2.464 3.228 ;
  LAYER M3 ;
        RECT 2.496 0.72 2.528 3.228 ;
  LAYER M3 ;
        RECT 2.56 0.72 2.592 3.228 ;
  LAYER M3 ;
        RECT 2.624 0.72 2.656 3.228 ;
  LAYER M3 ;
        RECT 2.688 0.72 2.72 3.228 ;
  LAYER M3 ;
        RECT 2.784 0.72 2.816 3.228 ;
  LAYER M1 ;
        RECT 0.399 0.756 0.401 3.192 ;
  LAYER M1 ;
        RECT 0.479 0.756 0.481 3.192 ;
  LAYER M1 ;
        RECT 0.559 0.756 0.561 3.192 ;
  LAYER M1 ;
        RECT 0.639 0.756 0.641 3.192 ;
  LAYER M1 ;
        RECT 0.719 0.756 0.721 3.192 ;
  LAYER M1 ;
        RECT 0.799 0.756 0.801 3.192 ;
  LAYER M1 ;
        RECT 0.879 0.756 0.881 3.192 ;
  LAYER M1 ;
        RECT 0.959 0.756 0.961 3.192 ;
  LAYER M1 ;
        RECT 1.039 0.756 1.041 3.192 ;
  LAYER M1 ;
        RECT 1.119 0.756 1.121 3.192 ;
  LAYER M1 ;
        RECT 1.199 0.756 1.201 3.192 ;
  LAYER M1 ;
        RECT 1.279 0.756 1.281 3.192 ;
  LAYER M1 ;
        RECT 1.359 0.756 1.361 3.192 ;
  LAYER M1 ;
        RECT 1.439 0.756 1.441 3.192 ;
  LAYER M1 ;
        RECT 1.519 0.756 1.521 3.192 ;
  LAYER M1 ;
        RECT 1.599 0.756 1.601 3.192 ;
  LAYER M1 ;
        RECT 1.679 0.756 1.681 3.192 ;
  LAYER M1 ;
        RECT 1.759 0.756 1.761 3.192 ;
  LAYER M1 ;
        RECT 1.839 0.756 1.841 3.192 ;
  LAYER M1 ;
        RECT 1.919 0.756 1.921 3.192 ;
  LAYER M1 ;
        RECT 1.999 0.756 2.001 3.192 ;
  LAYER M1 ;
        RECT 2.079 0.756 2.081 3.192 ;
  LAYER M1 ;
        RECT 2.159 0.756 2.161 3.192 ;
  LAYER M1 ;
        RECT 2.239 0.756 2.241 3.192 ;
  LAYER M1 ;
        RECT 2.319 0.756 2.321 3.192 ;
  LAYER M1 ;
        RECT 2.399 0.756 2.401 3.192 ;
  LAYER M1 ;
        RECT 2.479 0.756 2.481 3.192 ;
  LAYER M1 ;
        RECT 2.559 0.756 2.561 3.192 ;
  LAYER M1 ;
        RECT 2.639 0.756 2.641 3.192 ;
  LAYER M1 ;
        RECT 2.719 0.756 2.721 3.192 ;
  LAYER M2 ;
        RECT 0.4 0.755 2.8 0.757 ;
  LAYER M2 ;
        RECT 0.4 0.839 2.8 0.841 ;
  LAYER M2 ;
        RECT 0.4 0.923 2.8 0.925 ;
  LAYER M2 ;
        RECT 0.4 1.007 2.8 1.009 ;
  LAYER M2 ;
        RECT 0.4 1.091 2.8 1.093 ;
  LAYER M2 ;
        RECT 0.4 1.175 2.8 1.177 ;
  LAYER M2 ;
        RECT 0.4 1.259 2.8 1.261 ;
  LAYER M2 ;
        RECT 0.4 1.343 2.8 1.345 ;
  LAYER M2 ;
        RECT 0.4 1.427 2.8 1.429 ;
  LAYER M2 ;
        RECT 0.4 1.511 2.8 1.513 ;
  LAYER M2 ;
        RECT 0.4 1.595 2.8 1.597 ;
  LAYER M2 ;
        RECT 0.4 1.679 2.8 1.681 ;
  LAYER M2 ;
        RECT 0.4 1.7625 2.8 1.7645 ;
  LAYER M2 ;
        RECT 0.4 1.847 2.8 1.849 ;
  LAYER M2 ;
        RECT 0.4 1.931 2.8 1.933 ;
  LAYER M2 ;
        RECT 0.4 2.015 2.8 2.017 ;
  LAYER M2 ;
        RECT 0.4 2.099 2.8 2.101 ;
  LAYER M2 ;
        RECT 0.4 2.183 2.8 2.185 ;
  LAYER M2 ;
        RECT 0.4 2.267 2.8 2.269 ;
  LAYER M2 ;
        RECT 0.4 2.351 2.8 2.353 ;
  LAYER M2 ;
        RECT 0.4 2.435 2.8 2.437 ;
  LAYER M2 ;
        RECT 0.4 2.519 2.8 2.521 ;
  LAYER M2 ;
        RECT 0.4 2.603 2.8 2.605 ;
  LAYER M2 ;
        RECT 0.4 2.687 2.8 2.689 ;
  LAYER M2 ;
        RECT 0.4 2.771 2.8 2.773 ;
  LAYER M2 ;
        RECT 0.4 2.855 2.8 2.857 ;
  LAYER M2 ;
        RECT 0.4 2.939 2.8 2.941 ;
  LAYER M2 ;
        RECT 0.4 3.023 2.8 3.025 ;
  LAYER M2 ;
        RECT 0.4 3.107 2.8 3.109 ;
  LAYER M1 ;
        RECT 0.384 3.66 0.416 6.168 ;
  LAYER M1 ;
        RECT 0.448 3.66 0.48 6.168 ;
  LAYER M1 ;
        RECT 0.512 3.66 0.544 6.168 ;
  LAYER M1 ;
        RECT 0.576 3.66 0.608 6.168 ;
  LAYER M1 ;
        RECT 0.64 3.66 0.672 6.168 ;
  LAYER M1 ;
        RECT 0.704 3.66 0.736 6.168 ;
  LAYER M1 ;
        RECT 0.768 3.66 0.8 6.168 ;
  LAYER M1 ;
        RECT 0.832 3.66 0.864 6.168 ;
  LAYER M1 ;
        RECT 0.896 3.66 0.928 6.168 ;
  LAYER M1 ;
        RECT 0.96 3.66 0.992 6.168 ;
  LAYER M1 ;
        RECT 1.024 3.66 1.056 6.168 ;
  LAYER M1 ;
        RECT 1.088 3.66 1.12 6.168 ;
  LAYER M1 ;
        RECT 1.152 3.66 1.184 6.168 ;
  LAYER M1 ;
        RECT 1.216 3.66 1.248 6.168 ;
  LAYER M1 ;
        RECT 1.28 3.66 1.312 6.168 ;
  LAYER M1 ;
        RECT 1.344 3.66 1.376 6.168 ;
  LAYER M1 ;
        RECT 1.408 3.66 1.44 6.168 ;
  LAYER M1 ;
        RECT 1.472 3.66 1.504 6.168 ;
  LAYER M1 ;
        RECT 1.536 3.66 1.568 6.168 ;
  LAYER M1 ;
        RECT 1.6 3.66 1.632 6.168 ;
  LAYER M1 ;
        RECT 1.664 3.66 1.696 6.168 ;
  LAYER M1 ;
        RECT 1.728 3.66 1.76 6.168 ;
  LAYER M1 ;
        RECT 1.792 3.66 1.824 6.168 ;
  LAYER M1 ;
        RECT 1.856 3.66 1.888 6.168 ;
  LAYER M1 ;
        RECT 1.92 3.66 1.952 6.168 ;
  LAYER M1 ;
        RECT 1.984 3.66 2.016 6.168 ;
  LAYER M1 ;
        RECT 2.048 3.66 2.08 6.168 ;
  LAYER M1 ;
        RECT 2.112 3.66 2.144 6.168 ;
  LAYER M1 ;
        RECT 2.176 3.66 2.208 6.168 ;
  LAYER M1 ;
        RECT 2.24 3.66 2.272 6.168 ;
  LAYER M1 ;
        RECT 2.304 3.66 2.336 6.168 ;
  LAYER M1 ;
        RECT 2.368 3.66 2.4 6.168 ;
  LAYER M1 ;
        RECT 2.432 3.66 2.464 6.168 ;
  LAYER M1 ;
        RECT 2.496 3.66 2.528 6.168 ;
  LAYER M1 ;
        RECT 2.56 3.66 2.592 6.168 ;
  LAYER M1 ;
        RECT 2.624 3.66 2.656 6.168 ;
  LAYER M1 ;
        RECT 2.688 3.66 2.72 6.168 ;
  LAYER M2 ;
        RECT 0.364 3.744 2.836 3.776 ;
  LAYER M2 ;
        RECT 0.364 3.808 2.836 3.84 ;
  LAYER M2 ;
        RECT 0.364 3.872 2.836 3.904 ;
  LAYER M2 ;
        RECT 0.364 3.936 2.836 3.968 ;
  LAYER M2 ;
        RECT 0.364 4 2.836 4.032 ;
  LAYER M2 ;
        RECT 0.364 4.064 2.836 4.096 ;
  LAYER M2 ;
        RECT 0.364 4.128 2.836 4.16 ;
  LAYER M2 ;
        RECT 0.364 4.192 2.836 4.224 ;
  LAYER M2 ;
        RECT 0.364 4.256 2.836 4.288 ;
  LAYER M2 ;
        RECT 0.364 4.32 2.836 4.352 ;
  LAYER M2 ;
        RECT 0.364 4.384 2.836 4.416 ;
  LAYER M2 ;
        RECT 0.364 4.448 2.836 4.48 ;
  LAYER M2 ;
        RECT 0.364 4.512 2.836 4.544 ;
  LAYER M2 ;
        RECT 0.364 4.576 2.836 4.608 ;
  LAYER M2 ;
        RECT 0.364 4.64 2.836 4.672 ;
  LAYER M2 ;
        RECT 0.364 4.704 2.836 4.736 ;
  LAYER M2 ;
        RECT 0.364 4.768 2.836 4.8 ;
  LAYER M2 ;
        RECT 0.364 4.832 2.836 4.864 ;
  LAYER M2 ;
        RECT 0.364 4.896 2.836 4.928 ;
  LAYER M2 ;
        RECT 0.364 4.96 2.836 4.992 ;
  LAYER M2 ;
        RECT 0.364 5.024 2.836 5.056 ;
  LAYER M2 ;
        RECT 0.364 5.088 2.836 5.12 ;
  LAYER M2 ;
        RECT 0.364 5.152 2.836 5.184 ;
  LAYER M2 ;
        RECT 0.364 5.216 2.836 5.248 ;
  LAYER M2 ;
        RECT 0.364 5.28 2.836 5.312 ;
  LAYER M2 ;
        RECT 0.364 5.344 2.836 5.376 ;
  LAYER M2 ;
        RECT 0.364 5.408 2.836 5.44 ;
  LAYER M2 ;
        RECT 0.364 5.472 2.836 5.504 ;
  LAYER M2 ;
        RECT 0.364 5.536 2.836 5.568 ;
  LAYER M2 ;
        RECT 0.364 5.6 2.836 5.632 ;
  LAYER M2 ;
        RECT 0.364 5.664 2.836 5.696 ;
  LAYER M2 ;
        RECT 0.364 5.728 2.836 5.76 ;
  LAYER M2 ;
        RECT 0.364 5.792 2.836 5.824 ;
  LAYER M2 ;
        RECT 0.364 5.856 2.836 5.888 ;
  LAYER M2 ;
        RECT 0.364 5.92 2.836 5.952 ;
  LAYER M2 ;
        RECT 0.364 5.984 2.836 6.016 ;
  LAYER M3 ;
        RECT 0.384 3.66 0.416 6.168 ;
  LAYER M3 ;
        RECT 0.448 3.66 0.48 6.168 ;
  LAYER M3 ;
        RECT 0.512 3.66 0.544 6.168 ;
  LAYER M3 ;
        RECT 0.576 3.66 0.608 6.168 ;
  LAYER M3 ;
        RECT 0.64 3.66 0.672 6.168 ;
  LAYER M3 ;
        RECT 0.704 3.66 0.736 6.168 ;
  LAYER M3 ;
        RECT 0.768 3.66 0.8 6.168 ;
  LAYER M3 ;
        RECT 0.832 3.66 0.864 6.168 ;
  LAYER M3 ;
        RECT 0.896 3.66 0.928 6.168 ;
  LAYER M3 ;
        RECT 0.96 3.66 0.992 6.168 ;
  LAYER M3 ;
        RECT 1.024 3.66 1.056 6.168 ;
  LAYER M3 ;
        RECT 1.088 3.66 1.12 6.168 ;
  LAYER M3 ;
        RECT 1.152 3.66 1.184 6.168 ;
  LAYER M3 ;
        RECT 1.216 3.66 1.248 6.168 ;
  LAYER M3 ;
        RECT 1.28 3.66 1.312 6.168 ;
  LAYER M3 ;
        RECT 1.344 3.66 1.376 6.168 ;
  LAYER M3 ;
        RECT 1.408 3.66 1.44 6.168 ;
  LAYER M3 ;
        RECT 1.472 3.66 1.504 6.168 ;
  LAYER M3 ;
        RECT 1.536 3.66 1.568 6.168 ;
  LAYER M3 ;
        RECT 1.6 3.66 1.632 6.168 ;
  LAYER M3 ;
        RECT 1.664 3.66 1.696 6.168 ;
  LAYER M3 ;
        RECT 1.728 3.66 1.76 6.168 ;
  LAYER M3 ;
        RECT 1.792 3.66 1.824 6.168 ;
  LAYER M3 ;
        RECT 1.856 3.66 1.888 6.168 ;
  LAYER M3 ;
        RECT 1.92 3.66 1.952 6.168 ;
  LAYER M3 ;
        RECT 1.984 3.66 2.016 6.168 ;
  LAYER M3 ;
        RECT 2.048 3.66 2.08 6.168 ;
  LAYER M3 ;
        RECT 2.112 3.66 2.144 6.168 ;
  LAYER M3 ;
        RECT 2.176 3.66 2.208 6.168 ;
  LAYER M3 ;
        RECT 2.24 3.66 2.272 6.168 ;
  LAYER M3 ;
        RECT 2.304 3.66 2.336 6.168 ;
  LAYER M3 ;
        RECT 2.368 3.66 2.4 6.168 ;
  LAYER M3 ;
        RECT 2.432 3.66 2.464 6.168 ;
  LAYER M3 ;
        RECT 2.496 3.66 2.528 6.168 ;
  LAYER M3 ;
        RECT 2.56 3.66 2.592 6.168 ;
  LAYER M3 ;
        RECT 2.624 3.66 2.656 6.168 ;
  LAYER M3 ;
        RECT 2.688 3.66 2.72 6.168 ;
  LAYER M3 ;
        RECT 2.784 3.66 2.816 6.168 ;
  LAYER M1 ;
        RECT 0.399 3.696 0.401 6.132 ;
  LAYER M1 ;
        RECT 0.479 3.696 0.481 6.132 ;
  LAYER M1 ;
        RECT 0.559 3.696 0.561 6.132 ;
  LAYER M1 ;
        RECT 0.639 3.696 0.641 6.132 ;
  LAYER M1 ;
        RECT 0.719 3.696 0.721 6.132 ;
  LAYER M1 ;
        RECT 0.799 3.696 0.801 6.132 ;
  LAYER M1 ;
        RECT 0.879 3.696 0.881 6.132 ;
  LAYER M1 ;
        RECT 0.959 3.696 0.961 6.132 ;
  LAYER M1 ;
        RECT 1.039 3.696 1.041 6.132 ;
  LAYER M1 ;
        RECT 1.119 3.696 1.121 6.132 ;
  LAYER M1 ;
        RECT 1.199 3.696 1.201 6.132 ;
  LAYER M1 ;
        RECT 1.279 3.696 1.281 6.132 ;
  LAYER M1 ;
        RECT 1.359 3.696 1.361 6.132 ;
  LAYER M1 ;
        RECT 1.439 3.696 1.441 6.132 ;
  LAYER M1 ;
        RECT 1.519 3.696 1.521 6.132 ;
  LAYER M1 ;
        RECT 1.599 3.696 1.601 6.132 ;
  LAYER M1 ;
        RECT 1.679 3.696 1.681 6.132 ;
  LAYER M1 ;
        RECT 1.759 3.696 1.761 6.132 ;
  LAYER M1 ;
        RECT 1.839 3.696 1.841 6.132 ;
  LAYER M1 ;
        RECT 1.919 3.696 1.921 6.132 ;
  LAYER M1 ;
        RECT 1.999 3.696 2.001 6.132 ;
  LAYER M1 ;
        RECT 2.079 3.696 2.081 6.132 ;
  LAYER M1 ;
        RECT 2.159 3.696 2.161 6.132 ;
  LAYER M1 ;
        RECT 2.239 3.696 2.241 6.132 ;
  LAYER M1 ;
        RECT 2.319 3.696 2.321 6.132 ;
  LAYER M1 ;
        RECT 2.399 3.696 2.401 6.132 ;
  LAYER M1 ;
        RECT 2.479 3.696 2.481 6.132 ;
  LAYER M1 ;
        RECT 2.559 3.696 2.561 6.132 ;
  LAYER M1 ;
        RECT 2.639 3.696 2.641 6.132 ;
  LAYER M1 ;
        RECT 2.719 3.696 2.721 6.132 ;
  LAYER M2 ;
        RECT 0.4 3.695 2.8 3.697 ;
  LAYER M2 ;
        RECT 0.4 3.779 2.8 3.781 ;
  LAYER M2 ;
        RECT 0.4 3.863 2.8 3.865 ;
  LAYER M2 ;
        RECT 0.4 3.947 2.8 3.949 ;
  LAYER M2 ;
        RECT 0.4 4.031 2.8 4.033 ;
  LAYER M2 ;
        RECT 0.4 4.115 2.8 4.117 ;
  LAYER M2 ;
        RECT 0.4 4.199 2.8 4.201 ;
  LAYER M2 ;
        RECT 0.4 4.283 2.8 4.285 ;
  LAYER M2 ;
        RECT 0.4 4.367 2.8 4.369 ;
  LAYER M2 ;
        RECT 0.4 4.451 2.8 4.453 ;
  LAYER M2 ;
        RECT 0.4 4.535 2.8 4.537 ;
  LAYER M2 ;
        RECT 0.4 4.619 2.8 4.621 ;
  LAYER M2 ;
        RECT 0.4 4.7025 2.8 4.7045 ;
  LAYER M2 ;
        RECT 0.4 4.787 2.8 4.789 ;
  LAYER M2 ;
        RECT 0.4 4.871 2.8 4.873 ;
  LAYER M2 ;
        RECT 0.4 4.955 2.8 4.957 ;
  LAYER M2 ;
        RECT 0.4 5.039 2.8 5.041 ;
  LAYER M2 ;
        RECT 0.4 5.123 2.8 5.125 ;
  LAYER M2 ;
        RECT 0.4 5.207 2.8 5.209 ;
  LAYER M2 ;
        RECT 0.4 5.291 2.8 5.293 ;
  LAYER M2 ;
        RECT 0.4 5.375 2.8 5.377 ;
  LAYER M2 ;
        RECT 0.4 5.459 2.8 5.461 ;
  LAYER M2 ;
        RECT 0.4 5.543 2.8 5.545 ;
  LAYER M2 ;
        RECT 0.4 5.627 2.8 5.629 ;
  LAYER M2 ;
        RECT 0.4 5.711 2.8 5.713 ;
  LAYER M2 ;
        RECT 0.4 5.795 2.8 5.797 ;
  LAYER M2 ;
        RECT 0.4 5.879 2.8 5.881 ;
  LAYER M2 ;
        RECT 0.4 5.963 2.8 5.965 ;
  LAYER M2 ;
        RECT 0.4 6.047 2.8 6.049 ;
  LAYER M1 ;
        RECT 0.384 6.6 0.416 9.108 ;
  LAYER M1 ;
        RECT 0.448 6.6 0.48 9.108 ;
  LAYER M1 ;
        RECT 0.512 6.6 0.544 9.108 ;
  LAYER M1 ;
        RECT 0.576 6.6 0.608 9.108 ;
  LAYER M1 ;
        RECT 0.64 6.6 0.672 9.108 ;
  LAYER M1 ;
        RECT 0.704 6.6 0.736 9.108 ;
  LAYER M1 ;
        RECT 0.768 6.6 0.8 9.108 ;
  LAYER M1 ;
        RECT 0.832 6.6 0.864 9.108 ;
  LAYER M1 ;
        RECT 0.896 6.6 0.928 9.108 ;
  LAYER M1 ;
        RECT 0.96 6.6 0.992 9.108 ;
  LAYER M1 ;
        RECT 1.024 6.6 1.056 9.108 ;
  LAYER M1 ;
        RECT 1.088 6.6 1.12 9.108 ;
  LAYER M1 ;
        RECT 1.152 6.6 1.184 9.108 ;
  LAYER M1 ;
        RECT 1.216 6.6 1.248 9.108 ;
  LAYER M1 ;
        RECT 1.28 6.6 1.312 9.108 ;
  LAYER M1 ;
        RECT 1.344 6.6 1.376 9.108 ;
  LAYER M1 ;
        RECT 1.408 6.6 1.44 9.108 ;
  LAYER M1 ;
        RECT 1.472 6.6 1.504 9.108 ;
  LAYER M1 ;
        RECT 1.536 6.6 1.568 9.108 ;
  LAYER M1 ;
        RECT 1.6 6.6 1.632 9.108 ;
  LAYER M1 ;
        RECT 1.664 6.6 1.696 9.108 ;
  LAYER M1 ;
        RECT 1.728 6.6 1.76 9.108 ;
  LAYER M1 ;
        RECT 1.792 6.6 1.824 9.108 ;
  LAYER M1 ;
        RECT 1.856 6.6 1.888 9.108 ;
  LAYER M1 ;
        RECT 1.92 6.6 1.952 9.108 ;
  LAYER M1 ;
        RECT 1.984 6.6 2.016 9.108 ;
  LAYER M1 ;
        RECT 2.048 6.6 2.08 9.108 ;
  LAYER M1 ;
        RECT 2.112 6.6 2.144 9.108 ;
  LAYER M1 ;
        RECT 2.176 6.6 2.208 9.108 ;
  LAYER M1 ;
        RECT 2.24 6.6 2.272 9.108 ;
  LAYER M1 ;
        RECT 2.304 6.6 2.336 9.108 ;
  LAYER M1 ;
        RECT 2.368 6.6 2.4 9.108 ;
  LAYER M1 ;
        RECT 2.432 6.6 2.464 9.108 ;
  LAYER M1 ;
        RECT 2.496 6.6 2.528 9.108 ;
  LAYER M1 ;
        RECT 2.56 6.6 2.592 9.108 ;
  LAYER M1 ;
        RECT 2.624 6.6 2.656 9.108 ;
  LAYER M1 ;
        RECT 2.688 6.6 2.72 9.108 ;
  LAYER M2 ;
        RECT 0.364 6.684 2.836 6.716 ;
  LAYER M2 ;
        RECT 0.364 6.748 2.836 6.78 ;
  LAYER M2 ;
        RECT 0.364 6.812 2.836 6.844 ;
  LAYER M2 ;
        RECT 0.364 6.876 2.836 6.908 ;
  LAYER M2 ;
        RECT 0.364 6.94 2.836 6.972 ;
  LAYER M2 ;
        RECT 0.364 7.004 2.836 7.036 ;
  LAYER M2 ;
        RECT 0.364 7.068 2.836 7.1 ;
  LAYER M2 ;
        RECT 0.364 7.132 2.836 7.164 ;
  LAYER M2 ;
        RECT 0.364 7.196 2.836 7.228 ;
  LAYER M2 ;
        RECT 0.364 7.26 2.836 7.292 ;
  LAYER M2 ;
        RECT 0.364 7.324 2.836 7.356 ;
  LAYER M2 ;
        RECT 0.364 7.388 2.836 7.42 ;
  LAYER M2 ;
        RECT 0.364 7.452 2.836 7.484 ;
  LAYER M2 ;
        RECT 0.364 7.516 2.836 7.548 ;
  LAYER M2 ;
        RECT 0.364 7.58 2.836 7.612 ;
  LAYER M2 ;
        RECT 0.364 7.644 2.836 7.676 ;
  LAYER M2 ;
        RECT 0.364 7.708 2.836 7.74 ;
  LAYER M2 ;
        RECT 0.364 7.772 2.836 7.804 ;
  LAYER M2 ;
        RECT 0.364 7.836 2.836 7.868 ;
  LAYER M2 ;
        RECT 0.364 7.9 2.836 7.932 ;
  LAYER M2 ;
        RECT 0.364 7.964 2.836 7.996 ;
  LAYER M2 ;
        RECT 0.364 8.028 2.836 8.06 ;
  LAYER M2 ;
        RECT 0.364 8.092 2.836 8.124 ;
  LAYER M2 ;
        RECT 0.364 8.156 2.836 8.188 ;
  LAYER M2 ;
        RECT 0.364 8.22 2.836 8.252 ;
  LAYER M2 ;
        RECT 0.364 8.284 2.836 8.316 ;
  LAYER M2 ;
        RECT 0.364 8.348 2.836 8.38 ;
  LAYER M2 ;
        RECT 0.364 8.412 2.836 8.444 ;
  LAYER M2 ;
        RECT 0.364 8.476 2.836 8.508 ;
  LAYER M2 ;
        RECT 0.364 8.54 2.836 8.572 ;
  LAYER M2 ;
        RECT 0.364 8.604 2.836 8.636 ;
  LAYER M2 ;
        RECT 0.364 8.668 2.836 8.7 ;
  LAYER M2 ;
        RECT 0.364 8.732 2.836 8.764 ;
  LAYER M2 ;
        RECT 0.364 8.796 2.836 8.828 ;
  LAYER M2 ;
        RECT 0.364 8.86 2.836 8.892 ;
  LAYER M2 ;
        RECT 0.364 8.924 2.836 8.956 ;
  LAYER M3 ;
        RECT 0.384 6.6 0.416 9.108 ;
  LAYER M3 ;
        RECT 0.448 6.6 0.48 9.108 ;
  LAYER M3 ;
        RECT 0.512 6.6 0.544 9.108 ;
  LAYER M3 ;
        RECT 0.576 6.6 0.608 9.108 ;
  LAYER M3 ;
        RECT 0.64 6.6 0.672 9.108 ;
  LAYER M3 ;
        RECT 0.704 6.6 0.736 9.108 ;
  LAYER M3 ;
        RECT 0.768 6.6 0.8 9.108 ;
  LAYER M3 ;
        RECT 0.832 6.6 0.864 9.108 ;
  LAYER M3 ;
        RECT 0.896 6.6 0.928 9.108 ;
  LAYER M3 ;
        RECT 0.96 6.6 0.992 9.108 ;
  LAYER M3 ;
        RECT 1.024 6.6 1.056 9.108 ;
  LAYER M3 ;
        RECT 1.088 6.6 1.12 9.108 ;
  LAYER M3 ;
        RECT 1.152 6.6 1.184 9.108 ;
  LAYER M3 ;
        RECT 1.216 6.6 1.248 9.108 ;
  LAYER M3 ;
        RECT 1.28 6.6 1.312 9.108 ;
  LAYER M3 ;
        RECT 1.344 6.6 1.376 9.108 ;
  LAYER M3 ;
        RECT 1.408 6.6 1.44 9.108 ;
  LAYER M3 ;
        RECT 1.472 6.6 1.504 9.108 ;
  LAYER M3 ;
        RECT 1.536 6.6 1.568 9.108 ;
  LAYER M3 ;
        RECT 1.6 6.6 1.632 9.108 ;
  LAYER M3 ;
        RECT 1.664 6.6 1.696 9.108 ;
  LAYER M3 ;
        RECT 1.728 6.6 1.76 9.108 ;
  LAYER M3 ;
        RECT 1.792 6.6 1.824 9.108 ;
  LAYER M3 ;
        RECT 1.856 6.6 1.888 9.108 ;
  LAYER M3 ;
        RECT 1.92 6.6 1.952 9.108 ;
  LAYER M3 ;
        RECT 1.984 6.6 2.016 9.108 ;
  LAYER M3 ;
        RECT 2.048 6.6 2.08 9.108 ;
  LAYER M3 ;
        RECT 2.112 6.6 2.144 9.108 ;
  LAYER M3 ;
        RECT 2.176 6.6 2.208 9.108 ;
  LAYER M3 ;
        RECT 2.24 6.6 2.272 9.108 ;
  LAYER M3 ;
        RECT 2.304 6.6 2.336 9.108 ;
  LAYER M3 ;
        RECT 2.368 6.6 2.4 9.108 ;
  LAYER M3 ;
        RECT 2.432 6.6 2.464 9.108 ;
  LAYER M3 ;
        RECT 2.496 6.6 2.528 9.108 ;
  LAYER M3 ;
        RECT 2.56 6.6 2.592 9.108 ;
  LAYER M3 ;
        RECT 2.624 6.6 2.656 9.108 ;
  LAYER M3 ;
        RECT 2.688 6.6 2.72 9.108 ;
  LAYER M3 ;
        RECT 2.784 6.6 2.816 9.108 ;
  LAYER M1 ;
        RECT 0.399 6.636 0.401 9.072 ;
  LAYER M1 ;
        RECT 0.479 6.636 0.481 9.072 ;
  LAYER M1 ;
        RECT 0.559 6.636 0.561 9.072 ;
  LAYER M1 ;
        RECT 0.639 6.636 0.641 9.072 ;
  LAYER M1 ;
        RECT 0.719 6.636 0.721 9.072 ;
  LAYER M1 ;
        RECT 0.799 6.636 0.801 9.072 ;
  LAYER M1 ;
        RECT 0.879 6.636 0.881 9.072 ;
  LAYER M1 ;
        RECT 0.959 6.636 0.961 9.072 ;
  LAYER M1 ;
        RECT 1.039 6.636 1.041 9.072 ;
  LAYER M1 ;
        RECT 1.119 6.636 1.121 9.072 ;
  LAYER M1 ;
        RECT 1.199 6.636 1.201 9.072 ;
  LAYER M1 ;
        RECT 1.279 6.636 1.281 9.072 ;
  LAYER M1 ;
        RECT 1.359 6.636 1.361 9.072 ;
  LAYER M1 ;
        RECT 1.439 6.636 1.441 9.072 ;
  LAYER M1 ;
        RECT 1.519 6.636 1.521 9.072 ;
  LAYER M1 ;
        RECT 1.599 6.636 1.601 9.072 ;
  LAYER M1 ;
        RECT 1.679 6.636 1.681 9.072 ;
  LAYER M1 ;
        RECT 1.759 6.636 1.761 9.072 ;
  LAYER M1 ;
        RECT 1.839 6.636 1.841 9.072 ;
  LAYER M1 ;
        RECT 1.919 6.636 1.921 9.072 ;
  LAYER M1 ;
        RECT 1.999 6.636 2.001 9.072 ;
  LAYER M1 ;
        RECT 2.079 6.636 2.081 9.072 ;
  LAYER M1 ;
        RECT 2.159 6.636 2.161 9.072 ;
  LAYER M1 ;
        RECT 2.239 6.636 2.241 9.072 ;
  LAYER M1 ;
        RECT 2.319 6.636 2.321 9.072 ;
  LAYER M1 ;
        RECT 2.399 6.636 2.401 9.072 ;
  LAYER M1 ;
        RECT 2.479 6.636 2.481 9.072 ;
  LAYER M1 ;
        RECT 2.559 6.636 2.561 9.072 ;
  LAYER M1 ;
        RECT 2.639 6.636 2.641 9.072 ;
  LAYER M1 ;
        RECT 2.719 6.636 2.721 9.072 ;
  LAYER M2 ;
        RECT 0.4 6.635 2.8 6.637 ;
  LAYER M2 ;
        RECT 0.4 6.719 2.8 6.721 ;
  LAYER M2 ;
        RECT 0.4 6.803 2.8 6.805 ;
  LAYER M2 ;
        RECT 0.4 6.887 2.8 6.889 ;
  LAYER M2 ;
        RECT 0.4 6.971 2.8 6.973 ;
  LAYER M2 ;
        RECT 0.4 7.055 2.8 7.057 ;
  LAYER M2 ;
        RECT 0.4 7.139 2.8 7.141 ;
  LAYER M2 ;
        RECT 0.4 7.223 2.8 7.225 ;
  LAYER M2 ;
        RECT 0.4 7.307 2.8 7.309 ;
  LAYER M2 ;
        RECT 0.4 7.391 2.8 7.393 ;
  LAYER M2 ;
        RECT 0.4 7.475 2.8 7.477 ;
  LAYER M2 ;
        RECT 0.4 7.559 2.8 7.561 ;
  LAYER M2 ;
        RECT 0.4 7.6425 2.8 7.6445 ;
  LAYER M2 ;
        RECT 0.4 7.727 2.8 7.729 ;
  LAYER M2 ;
        RECT 0.4 7.811 2.8 7.813 ;
  LAYER M2 ;
        RECT 0.4 7.895 2.8 7.897 ;
  LAYER M2 ;
        RECT 0.4 7.979 2.8 7.981 ;
  LAYER M2 ;
        RECT 0.4 8.063 2.8 8.065 ;
  LAYER M2 ;
        RECT 0.4 8.147 2.8 8.149 ;
  LAYER M2 ;
        RECT 0.4 8.231 2.8 8.233 ;
  LAYER M2 ;
        RECT 0.4 8.315 2.8 8.317 ;
  LAYER M2 ;
        RECT 0.4 8.399 2.8 8.401 ;
  LAYER M2 ;
        RECT 0.4 8.483 2.8 8.485 ;
  LAYER M2 ;
        RECT 0.4 8.567 2.8 8.569 ;
  LAYER M2 ;
        RECT 0.4 8.651 2.8 8.653 ;
  LAYER M2 ;
        RECT 0.4 8.735 2.8 8.737 ;
  LAYER M2 ;
        RECT 0.4 8.819 2.8 8.821 ;
  LAYER M2 ;
        RECT 0.4 8.903 2.8 8.905 ;
  LAYER M2 ;
        RECT 0.4 8.987 2.8 8.989 ;
  LAYER M1 ;
        RECT 0.384 9.54 0.416 12.048 ;
  LAYER M1 ;
        RECT 0.448 9.54 0.48 12.048 ;
  LAYER M1 ;
        RECT 0.512 9.54 0.544 12.048 ;
  LAYER M1 ;
        RECT 0.576 9.54 0.608 12.048 ;
  LAYER M1 ;
        RECT 0.64 9.54 0.672 12.048 ;
  LAYER M1 ;
        RECT 0.704 9.54 0.736 12.048 ;
  LAYER M1 ;
        RECT 0.768 9.54 0.8 12.048 ;
  LAYER M1 ;
        RECT 0.832 9.54 0.864 12.048 ;
  LAYER M1 ;
        RECT 0.896 9.54 0.928 12.048 ;
  LAYER M1 ;
        RECT 0.96 9.54 0.992 12.048 ;
  LAYER M1 ;
        RECT 1.024 9.54 1.056 12.048 ;
  LAYER M1 ;
        RECT 1.088 9.54 1.12 12.048 ;
  LAYER M1 ;
        RECT 1.152 9.54 1.184 12.048 ;
  LAYER M1 ;
        RECT 1.216 9.54 1.248 12.048 ;
  LAYER M1 ;
        RECT 1.28 9.54 1.312 12.048 ;
  LAYER M1 ;
        RECT 1.344 9.54 1.376 12.048 ;
  LAYER M1 ;
        RECT 1.408 9.54 1.44 12.048 ;
  LAYER M1 ;
        RECT 1.472 9.54 1.504 12.048 ;
  LAYER M1 ;
        RECT 1.536 9.54 1.568 12.048 ;
  LAYER M1 ;
        RECT 1.6 9.54 1.632 12.048 ;
  LAYER M1 ;
        RECT 1.664 9.54 1.696 12.048 ;
  LAYER M1 ;
        RECT 1.728 9.54 1.76 12.048 ;
  LAYER M1 ;
        RECT 1.792 9.54 1.824 12.048 ;
  LAYER M1 ;
        RECT 1.856 9.54 1.888 12.048 ;
  LAYER M1 ;
        RECT 1.92 9.54 1.952 12.048 ;
  LAYER M1 ;
        RECT 1.984 9.54 2.016 12.048 ;
  LAYER M1 ;
        RECT 2.048 9.54 2.08 12.048 ;
  LAYER M1 ;
        RECT 2.112 9.54 2.144 12.048 ;
  LAYER M1 ;
        RECT 2.176 9.54 2.208 12.048 ;
  LAYER M1 ;
        RECT 2.24 9.54 2.272 12.048 ;
  LAYER M1 ;
        RECT 2.304 9.54 2.336 12.048 ;
  LAYER M1 ;
        RECT 2.368 9.54 2.4 12.048 ;
  LAYER M1 ;
        RECT 2.432 9.54 2.464 12.048 ;
  LAYER M1 ;
        RECT 2.496 9.54 2.528 12.048 ;
  LAYER M1 ;
        RECT 2.56 9.54 2.592 12.048 ;
  LAYER M1 ;
        RECT 2.624 9.54 2.656 12.048 ;
  LAYER M1 ;
        RECT 2.688 9.54 2.72 12.048 ;
  LAYER M2 ;
        RECT 0.364 9.624 2.836 9.656 ;
  LAYER M2 ;
        RECT 0.364 9.688 2.836 9.72 ;
  LAYER M2 ;
        RECT 0.364 9.752 2.836 9.784 ;
  LAYER M2 ;
        RECT 0.364 9.816 2.836 9.848 ;
  LAYER M2 ;
        RECT 0.364 9.88 2.836 9.912 ;
  LAYER M2 ;
        RECT 0.364 9.944 2.836 9.976 ;
  LAYER M2 ;
        RECT 0.364 10.008 2.836 10.04 ;
  LAYER M2 ;
        RECT 0.364 10.072 2.836 10.104 ;
  LAYER M2 ;
        RECT 0.364 10.136 2.836 10.168 ;
  LAYER M2 ;
        RECT 0.364 10.2 2.836 10.232 ;
  LAYER M2 ;
        RECT 0.364 10.264 2.836 10.296 ;
  LAYER M2 ;
        RECT 0.364 10.328 2.836 10.36 ;
  LAYER M2 ;
        RECT 0.364 10.392 2.836 10.424 ;
  LAYER M2 ;
        RECT 0.364 10.456 2.836 10.488 ;
  LAYER M2 ;
        RECT 0.364 10.52 2.836 10.552 ;
  LAYER M2 ;
        RECT 0.364 10.584 2.836 10.616 ;
  LAYER M2 ;
        RECT 0.364 10.648 2.836 10.68 ;
  LAYER M2 ;
        RECT 0.364 10.712 2.836 10.744 ;
  LAYER M2 ;
        RECT 0.364 10.776 2.836 10.808 ;
  LAYER M2 ;
        RECT 0.364 10.84 2.836 10.872 ;
  LAYER M2 ;
        RECT 0.364 10.904 2.836 10.936 ;
  LAYER M2 ;
        RECT 0.364 10.968 2.836 11 ;
  LAYER M2 ;
        RECT 0.364 11.032 2.836 11.064 ;
  LAYER M2 ;
        RECT 0.364 11.096 2.836 11.128 ;
  LAYER M2 ;
        RECT 0.364 11.16 2.836 11.192 ;
  LAYER M2 ;
        RECT 0.364 11.224 2.836 11.256 ;
  LAYER M2 ;
        RECT 0.364 11.288 2.836 11.32 ;
  LAYER M2 ;
        RECT 0.364 11.352 2.836 11.384 ;
  LAYER M2 ;
        RECT 0.364 11.416 2.836 11.448 ;
  LAYER M2 ;
        RECT 0.364 11.48 2.836 11.512 ;
  LAYER M2 ;
        RECT 0.364 11.544 2.836 11.576 ;
  LAYER M2 ;
        RECT 0.364 11.608 2.836 11.64 ;
  LAYER M2 ;
        RECT 0.364 11.672 2.836 11.704 ;
  LAYER M2 ;
        RECT 0.364 11.736 2.836 11.768 ;
  LAYER M2 ;
        RECT 0.364 11.8 2.836 11.832 ;
  LAYER M2 ;
        RECT 0.364 11.864 2.836 11.896 ;
  LAYER M3 ;
        RECT 0.384 9.54 0.416 12.048 ;
  LAYER M3 ;
        RECT 0.448 9.54 0.48 12.048 ;
  LAYER M3 ;
        RECT 0.512 9.54 0.544 12.048 ;
  LAYER M3 ;
        RECT 0.576 9.54 0.608 12.048 ;
  LAYER M3 ;
        RECT 0.64 9.54 0.672 12.048 ;
  LAYER M3 ;
        RECT 0.704 9.54 0.736 12.048 ;
  LAYER M3 ;
        RECT 0.768 9.54 0.8 12.048 ;
  LAYER M3 ;
        RECT 0.832 9.54 0.864 12.048 ;
  LAYER M3 ;
        RECT 0.896 9.54 0.928 12.048 ;
  LAYER M3 ;
        RECT 0.96 9.54 0.992 12.048 ;
  LAYER M3 ;
        RECT 1.024 9.54 1.056 12.048 ;
  LAYER M3 ;
        RECT 1.088 9.54 1.12 12.048 ;
  LAYER M3 ;
        RECT 1.152 9.54 1.184 12.048 ;
  LAYER M3 ;
        RECT 1.216 9.54 1.248 12.048 ;
  LAYER M3 ;
        RECT 1.28 9.54 1.312 12.048 ;
  LAYER M3 ;
        RECT 1.344 9.54 1.376 12.048 ;
  LAYER M3 ;
        RECT 1.408 9.54 1.44 12.048 ;
  LAYER M3 ;
        RECT 1.472 9.54 1.504 12.048 ;
  LAYER M3 ;
        RECT 1.536 9.54 1.568 12.048 ;
  LAYER M3 ;
        RECT 1.6 9.54 1.632 12.048 ;
  LAYER M3 ;
        RECT 1.664 9.54 1.696 12.048 ;
  LAYER M3 ;
        RECT 1.728 9.54 1.76 12.048 ;
  LAYER M3 ;
        RECT 1.792 9.54 1.824 12.048 ;
  LAYER M3 ;
        RECT 1.856 9.54 1.888 12.048 ;
  LAYER M3 ;
        RECT 1.92 9.54 1.952 12.048 ;
  LAYER M3 ;
        RECT 1.984 9.54 2.016 12.048 ;
  LAYER M3 ;
        RECT 2.048 9.54 2.08 12.048 ;
  LAYER M3 ;
        RECT 2.112 9.54 2.144 12.048 ;
  LAYER M3 ;
        RECT 2.176 9.54 2.208 12.048 ;
  LAYER M3 ;
        RECT 2.24 9.54 2.272 12.048 ;
  LAYER M3 ;
        RECT 2.304 9.54 2.336 12.048 ;
  LAYER M3 ;
        RECT 2.368 9.54 2.4 12.048 ;
  LAYER M3 ;
        RECT 2.432 9.54 2.464 12.048 ;
  LAYER M3 ;
        RECT 2.496 9.54 2.528 12.048 ;
  LAYER M3 ;
        RECT 2.56 9.54 2.592 12.048 ;
  LAYER M3 ;
        RECT 2.624 9.54 2.656 12.048 ;
  LAYER M3 ;
        RECT 2.688 9.54 2.72 12.048 ;
  LAYER M3 ;
        RECT 2.784 9.54 2.816 12.048 ;
  LAYER M1 ;
        RECT 0.399 9.576 0.401 12.012 ;
  LAYER M1 ;
        RECT 0.479 9.576 0.481 12.012 ;
  LAYER M1 ;
        RECT 0.559 9.576 0.561 12.012 ;
  LAYER M1 ;
        RECT 0.639 9.576 0.641 12.012 ;
  LAYER M1 ;
        RECT 0.719 9.576 0.721 12.012 ;
  LAYER M1 ;
        RECT 0.799 9.576 0.801 12.012 ;
  LAYER M1 ;
        RECT 0.879 9.576 0.881 12.012 ;
  LAYER M1 ;
        RECT 0.959 9.576 0.961 12.012 ;
  LAYER M1 ;
        RECT 1.039 9.576 1.041 12.012 ;
  LAYER M1 ;
        RECT 1.119 9.576 1.121 12.012 ;
  LAYER M1 ;
        RECT 1.199 9.576 1.201 12.012 ;
  LAYER M1 ;
        RECT 1.279 9.576 1.281 12.012 ;
  LAYER M1 ;
        RECT 1.359 9.576 1.361 12.012 ;
  LAYER M1 ;
        RECT 1.439 9.576 1.441 12.012 ;
  LAYER M1 ;
        RECT 1.519 9.576 1.521 12.012 ;
  LAYER M1 ;
        RECT 1.599 9.576 1.601 12.012 ;
  LAYER M1 ;
        RECT 1.679 9.576 1.681 12.012 ;
  LAYER M1 ;
        RECT 1.759 9.576 1.761 12.012 ;
  LAYER M1 ;
        RECT 1.839 9.576 1.841 12.012 ;
  LAYER M1 ;
        RECT 1.919 9.576 1.921 12.012 ;
  LAYER M1 ;
        RECT 1.999 9.576 2.001 12.012 ;
  LAYER M1 ;
        RECT 2.079 9.576 2.081 12.012 ;
  LAYER M1 ;
        RECT 2.159 9.576 2.161 12.012 ;
  LAYER M1 ;
        RECT 2.239 9.576 2.241 12.012 ;
  LAYER M1 ;
        RECT 2.319 9.576 2.321 12.012 ;
  LAYER M1 ;
        RECT 2.399 9.576 2.401 12.012 ;
  LAYER M1 ;
        RECT 2.479 9.576 2.481 12.012 ;
  LAYER M1 ;
        RECT 2.559 9.576 2.561 12.012 ;
  LAYER M1 ;
        RECT 2.639 9.576 2.641 12.012 ;
  LAYER M1 ;
        RECT 2.719 9.576 2.721 12.012 ;
  LAYER M2 ;
        RECT 0.4 9.575 2.8 9.577 ;
  LAYER M2 ;
        RECT 0.4 9.659 2.8 9.661 ;
  LAYER M2 ;
        RECT 0.4 9.743 2.8 9.745 ;
  LAYER M2 ;
        RECT 0.4 9.827 2.8 9.829 ;
  LAYER M2 ;
        RECT 0.4 9.911 2.8 9.913 ;
  LAYER M2 ;
        RECT 0.4 9.995 2.8 9.997 ;
  LAYER M2 ;
        RECT 0.4 10.079 2.8 10.081 ;
  LAYER M2 ;
        RECT 0.4 10.163 2.8 10.165 ;
  LAYER M2 ;
        RECT 0.4 10.247 2.8 10.249 ;
  LAYER M2 ;
        RECT 0.4 10.331 2.8 10.333 ;
  LAYER M2 ;
        RECT 0.4 10.415 2.8 10.417 ;
  LAYER M2 ;
        RECT 0.4 10.499 2.8 10.501 ;
  LAYER M2 ;
        RECT 0.4 10.5825 2.8 10.5845 ;
  LAYER M2 ;
        RECT 0.4 10.667 2.8 10.669 ;
  LAYER M2 ;
        RECT 0.4 10.751 2.8 10.753 ;
  LAYER M2 ;
        RECT 0.4 10.835 2.8 10.837 ;
  LAYER M2 ;
        RECT 0.4 10.919 2.8 10.921 ;
  LAYER M2 ;
        RECT 0.4 11.003 2.8 11.005 ;
  LAYER M2 ;
        RECT 0.4 11.087 2.8 11.089 ;
  LAYER M2 ;
        RECT 0.4 11.171 2.8 11.173 ;
  LAYER M2 ;
        RECT 0.4 11.255 2.8 11.257 ;
  LAYER M2 ;
        RECT 0.4 11.339 2.8 11.341 ;
  LAYER M2 ;
        RECT 0.4 11.423 2.8 11.425 ;
  LAYER M2 ;
        RECT 0.4 11.507 2.8 11.509 ;
  LAYER M2 ;
        RECT 0.4 11.591 2.8 11.593 ;
  LAYER M2 ;
        RECT 0.4 11.675 2.8 11.677 ;
  LAYER M2 ;
        RECT 0.4 11.759 2.8 11.761 ;
  LAYER M2 ;
        RECT 0.4 11.843 2.8 11.845 ;
  LAYER M2 ;
        RECT 0.4 11.927 2.8 11.929 ;
  LAYER M1 ;
        RECT 0.384 12.48 0.416 14.988 ;
  LAYER M1 ;
        RECT 0.448 12.48 0.48 14.988 ;
  LAYER M1 ;
        RECT 0.512 12.48 0.544 14.988 ;
  LAYER M1 ;
        RECT 0.576 12.48 0.608 14.988 ;
  LAYER M1 ;
        RECT 0.64 12.48 0.672 14.988 ;
  LAYER M1 ;
        RECT 0.704 12.48 0.736 14.988 ;
  LAYER M1 ;
        RECT 0.768 12.48 0.8 14.988 ;
  LAYER M1 ;
        RECT 0.832 12.48 0.864 14.988 ;
  LAYER M1 ;
        RECT 0.896 12.48 0.928 14.988 ;
  LAYER M1 ;
        RECT 0.96 12.48 0.992 14.988 ;
  LAYER M1 ;
        RECT 1.024 12.48 1.056 14.988 ;
  LAYER M1 ;
        RECT 1.088 12.48 1.12 14.988 ;
  LAYER M1 ;
        RECT 1.152 12.48 1.184 14.988 ;
  LAYER M1 ;
        RECT 1.216 12.48 1.248 14.988 ;
  LAYER M1 ;
        RECT 1.28 12.48 1.312 14.988 ;
  LAYER M1 ;
        RECT 1.344 12.48 1.376 14.988 ;
  LAYER M1 ;
        RECT 1.408 12.48 1.44 14.988 ;
  LAYER M1 ;
        RECT 1.472 12.48 1.504 14.988 ;
  LAYER M1 ;
        RECT 1.536 12.48 1.568 14.988 ;
  LAYER M1 ;
        RECT 1.6 12.48 1.632 14.988 ;
  LAYER M1 ;
        RECT 1.664 12.48 1.696 14.988 ;
  LAYER M1 ;
        RECT 1.728 12.48 1.76 14.988 ;
  LAYER M1 ;
        RECT 1.792 12.48 1.824 14.988 ;
  LAYER M1 ;
        RECT 1.856 12.48 1.888 14.988 ;
  LAYER M1 ;
        RECT 1.92 12.48 1.952 14.988 ;
  LAYER M1 ;
        RECT 1.984 12.48 2.016 14.988 ;
  LAYER M1 ;
        RECT 2.048 12.48 2.08 14.988 ;
  LAYER M1 ;
        RECT 2.112 12.48 2.144 14.988 ;
  LAYER M1 ;
        RECT 2.176 12.48 2.208 14.988 ;
  LAYER M1 ;
        RECT 2.24 12.48 2.272 14.988 ;
  LAYER M1 ;
        RECT 2.304 12.48 2.336 14.988 ;
  LAYER M1 ;
        RECT 2.368 12.48 2.4 14.988 ;
  LAYER M1 ;
        RECT 2.432 12.48 2.464 14.988 ;
  LAYER M1 ;
        RECT 2.496 12.48 2.528 14.988 ;
  LAYER M1 ;
        RECT 2.56 12.48 2.592 14.988 ;
  LAYER M1 ;
        RECT 2.624 12.48 2.656 14.988 ;
  LAYER M1 ;
        RECT 2.688 12.48 2.72 14.988 ;
  LAYER M2 ;
        RECT 0.364 12.564 2.836 12.596 ;
  LAYER M2 ;
        RECT 0.364 12.628 2.836 12.66 ;
  LAYER M2 ;
        RECT 0.364 12.692 2.836 12.724 ;
  LAYER M2 ;
        RECT 0.364 12.756 2.836 12.788 ;
  LAYER M2 ;
        RECT 0.364 12.82 2.836 12.852 ;
  LAYER M2 ;
        RECT 0.364 12.884 2.836 12.916 ;
  LAYER M2 ;
        RECT 0.364 12.948 2.836 12.98 ;
  LAYER M2 ;
        RECT 0.364 13.012 2.836 13.044 ;
  LAYER M2 ;
        RECT 0.364 13.076 2.836 13.108 ;
  LAYER M2 ;
        RECT 0.364 13.14 2.836 13.172 ;
  LAYER M2 ;
        RECT 0.364 13.204 2.836 13.236 ;
  LAYER M2 ;
        RECT 0.364 13.268 2.836 13.3 ;
  LAYER M2 ;
        RECT 0.364 13.332 2.836 13.364 ;
  LAYER M2 ;
        RECT 0.364 13.396 2.836 13.428 ;
  LAYER M2 ;
        RECT 0.364 13.46 2.836 13.492 ;
  LAYER M2 ;
        RECT 0.364 13.524 2.836 13.556 ;
  LAYER M2 ;
        RECT 0.364 13.588 2.836 13.62 ;
  LAYER M2 ;
        RECT 0.364 13.652 2.836 13.684 ;
  LAYER M2 ;
        RECT 0.364 13.716 2.836 13.748 ;
  LAYER M2 ;
        RECT 0.364 13.78 2.836 13.812 ;
  LAYER M2 ;
        RECT 0.364 13.844 2.836 13.876 ;
  LAYER M2 ;
        RECT 0.364 13.908 2.836 13.94 ;
  LAYER M2 ;
        RECT 0.364 13.972 2.836 14.004 ;
  LAYER M2 ;
        RECT 0.364 14.036 2.836 14.068 ;
  LAYER M2 ;
        RECT 0.364 14.1 2.836 14.132 ;
  LAYER M2 ;
        RECT 0.364 14.164 2.836 14.196 ;
  LAYER M2 ;
        RECT 0.364 14.228 2.836 14.26 ;
  LAYER M2 ;
        RECT 0.364 14.292 2.836 14.324 ;
  LAYER M2 ;
        RECT 0.364 14.356 2.836 14.388 ;
  LAYER M2 ;
        RECT 0.364 14.42 2.836 14.452 ;
  LAYER M2 ;
        RECT 0.364 14.484 2.836 14.516 ;
  LAYER M2 ;
        RECT 0.364 14.548 2.836 14.58 ;
  LAYER M2 ;
        RECT 0.364 14.612 2.836 14.644 ;
  LAYER M2 ;
        RECT 0.364 14.676 2.836 14.708 ;
  LAYER M2 ;
        RECT 0.364 14.74 2.836 14.772 ;
  LAYER M2 ;
        RECT 0.364 14.804 2.836 14.836 ;
  LAYER M3 ;
        RECT 0.384 12.48 0.416 14.988 ;
  LAYER M3 ;
        RECT 0.448 12.48 0.48 14.988 ;
  LAYER M3 ;
        RECT 0.512 12.48 0.544 14.988 ;
  LAYER M3 ;
        RECT 0.576 12.48 0.608 14.988 ;
  LAYER M3 ;
        RECT 0.64 12.48 0.672 14.988 ;
  LAYER M3 ;
        RECT 0.704 12.48 0.736 14.988 ;
  LAYER M3 ;
        RECT 0.768 12.48 0.8 14.988 ;
  LAYER M3 ;
        RECT 0.832 12.48 0.864 14.988 ;
  LAYER M3 ;
        RECT 0.896 12.48 0.928 14.988 ;
  LAYER M3 ;
        RECT 0.96 12.48 0.992 14.988 ;
  LAYER M3 ;
        RECT 1.024 12.48 1.056 14.988 ;
  LAYER M3 ;
        RECT 1.088 12.48 1.12 14.988 ;
  LAYER M3 ;
        RECT 1.152 12.48 1.184 14.988 ;
  LAYER M3 ;
        RECT 1.216 12.48 1.248 14.988 ;
  LAYER M3 ;
        RECT 1.28 12.48 1.312 14.988 ;
  LAYER M3 ;
        RECT 1.344 12.48 1.376 14.988 ;
  LAYER M3 ;
        RECT 1.408 12.48 1.44 14.988 ;
  LAYER M3 ;
        RECT 1.472 12.48 1.504 14.988 ;
  LAYER M3 ;
        RECT 1.536 12.48 1.568 14.988 ;
  LAYER M3 ;
        RECT 1.6 12.48 1.632 14.988 ;
  LAYER M3 ;
        RECT 1.664 12.48 1.696 14.988 ;
  LAYER M3 ;
        RECT 1.728 12.48 1.76 14.988 ;
  LAYER M3 ;
        RECT 1.792 12.48 1.824 14.988 ;
  LAYER M3 ;
        RECT 1.856 12.48 1.888 14.988 ;
  LAYER M3 ;
        RECT 1.92 12.48 1.952 14.988 ;
  LAYER M3 ;
        RECT 1.984 12.48 2.016 14.988 ;
  LAYER M3 ;
        RECT 2.048 12.48 2.08 14.988 ;
  LAYER M3 ;
        RECT 2.112 12.48 2.144 14.988 ;
  LAYER M3 ;
        RECT 2.176 12.48 2.208 14.988 ;
  LAYER M3 ;
        RECT 2.24 12.48 2.272 14.988 ;
  LAYER M3 ;
        RECT 2.304 12.48 2.336 14.988 ;
  LAYER M3 ;
        RECT 2.368 12.48 2.4 14.988 ;
  LAYER M3 ;
        RECT 2.432 12.48 2.464 14.988 ;
  LAYER M3 ;
        RECT 2.496 12.48 2.528 14.988 ;
  LAYER M3 ;
        RECT 2.56 12.48 2.592 14.988 ;
  LAYER M3 ;
        RECT 2.624 12.48 2.656 14.988 ;
  LAYER M3 ;
        RECT 2.688 12.48 2.72 14.988 ;
  LAYER M3 ;
        RECT 2.784 12.48 2.816 14.988 ;
  LAYER M1 ;
        RECT 0.399 12.516 0.401 14.952 ;
  LAYER M1 ;
        RECT 0.479 12.516 0.481 14.952 ;
  LAYER M1 ;
        RECT 0.559 12.516 0.561 14.952 ;
  LAYER M1 ;
        RECT 0.639 12.516 0.641 14.952 ;
  LAYER M1 ;
        RECT 0.719 12.516 0.721 14.952 ;
  LAYER M1 ;
        RECT 0.799 12.516 0.801 14.952 ;
  LAYER M1 ;
        RECT 0.879 12.516 0.881 14.952 ;
  LAYER M1 ;
        RECT 0.959 12.516 0.961 14.952 ;
  LAYER M1 ;
        RECT 1.039 12.516 1.041 14.952 ;
  LAYER M1 ;
        RECT 1.119 12.516 1.121 14.952 ;
  LAYER M1 ;
        RECT 1.199 12.516 1.201 14.952 ;
  LAYER M1 ;
        RECT 1.279 12.516 1.281 14.952 ;
  LAYER M1 ;
        RECT 1.359 12.516 1.361 14.952 ;
  LAYER M1 ;
        RECT 1.439 12.516 1.441 14.952 ;
  LAYER M1 ;
        RECT 1.519 12.516 1.521 14.952 ;
  LAYER M1 ;
        RECT 1.599 12.516 1.601 14.952 ;
  LAYER M1 ;
        RECT 1.679 12.516 1.681 14.952 ;
  LAYER M1 ;
        RECT 1.759 12.516 1.761 14.952 ;
  LAYER M1 ;
        RECT 1.839 12.516 1.841 14.952 ;
  LAYER M1 ;
        RECT 1.919 12.516 1.921 14.952 ;
  LAYER M1 ;
        RECT 1.999 12.516 2.001 14.952 ;
  LAYER M1 ;
        RECT 2.079 12.516 2.081 14.952 ;
  LAYER M1 ;
        RECT 2.159 12.516 2.161 14.952 ;
  LAYER M1 ;
        RECT 2.239 12.516 2.241 14.952 ;
  LAYER M1 ;
        RECT 2.319 12.516 2.321 14.952 ;
  LAYER M1 ;
        RECT 2.399 12.516 2.401 14.952 ;
  LAYER M1 ;
        RECT 2.479 12.516 2.481 14.952 ;
  LAYER M1 ;
        RECT 2.559 12.516 2.561 14.952 ;
  LAYER M1 ;
        RECT 2.639 12.516 2.641 14.952 ;
  LAYER M1 ;
        RECT 2.719 12.516 2.721 14.952 ;
  LAYER M2 ;
        RECT 0.4 12.515 2.8 12.517 ;
  LAYER M2 ;
        RECT 0.4 12.599 2.8 12.601 ;
  LAYER M2 ;
        RECT 0.4 12.683 2.8 12.685 ;
  LAYER M2 ;
        RECT 0.4 12.767 2.8 12.769 ;
  LAYER M2 ;
        RECT 0.4 12.851 2.8 12.853 ;
  LAYER M2 ;
        RECT 0.4 12.935 2.8 12.937 ;
  LAYER M2 ;
        RECT 0.4 13.019 2.8 13.021 ;
  LAYER M2 ;
        RECT 0.4 13.103 2.8 13.105 ;
  LAYER M2 ;
        RECT 0.4 13.187 2.8 13.189 ;
  LAYER M2 ;
        RECT 0.4 13.271 2.8 13.273 ;
  LAYER M2 ;
        RECT 0.4 13.355 2.8 13.357 ;
  LAYER M2 ;
        RECT 0.4 13.439 2.8 13.441 ;
  LAYER M2 ;
        RECT 0.4 13.5225 2.8 13.5245 ;
  LAYER M2 ;
        RECT 0.4 13.607 2.8 13.609 ;
  LAYER M2 ;
        RECT 0.4 13.691 2.8 13.693 ;
  LAYER M2 ;
        RECT 0.4 13.775 2.8 13.777 ;
  LAYER M2 ;
        RECT 0.4 13.859 2.8 13.861 ;
  LAYER M2 ;
        RECT 0.4 13.943 2.8 13.945 ;
  LAYER M2 ;
        RECT 0.4 14.027 2.8 14.029 ;
  LAYER M2 ;
        RECT 0.4 14.111 2.8 14.113 ;
  LAYER M2 ;
        RECT 0.4 14.195 2.8 14.197 ;
  LAYER M2 ;
        RECT 0.4 14.279 2.8 14.281 ;
  LAYER M2 ;
        RECT 0.4 14.363 2.8 14.365 ;
  LAYER M2 ;
        RECT 0.4 14.447 2.8 14.449 ;
  LAYER M2 ;
        RECT 0.4 14.531 2.8 14.533 ;
  LAYER M2 ;
        RECT 0.4 14.615 2.8 14.617 ;
  LAYER M2 ;
        RECT 0.4 14.699 2.8 14.701 ;
  LAYER M2 ;
        RECT 0.4 14.783 2.8 14.785 ;
  LAYER M2 ;
        RECT 0.4 14.867 2.8 14.869 ;
  LAYER M1 ;
        RECT 0.384 15.42 0.416 17.928 ;
  LAYER M1 ;
        RECT 0.448 15.42 0.48 17.928 ;
  LAYER M1 ;
        RECT 0.512 15.42 0.544 17.928 ;
  LAYER M1 ;
        RECT 0.576 15.42 0.608 17.928 ;
  LAYER M1 ;
        RECT 0.64 15.42 0.672 17.928 ;
  LAYER M1 ;
        RECT 0.704 15.42 0.736 17.928 ;
  LAYER M1 ;
        RECT 0.768 15.42 0.8 17.928 ;
  LAYER M1 ;
        RECT 0.832 15.42 0.864 17.928 ;
  LAYER M1 ;
        RECT 0.896 15.42 0.928 17.928 ;
  LAYER M1 ;
        RECT 0.96 15.42 0.992 17.928 ;
  LAYER M1 ;
        RECT 1.024 15.42 1.056 17.928 ;
  LAYER M1 ;
        RECT 1.088 15.42 1.12 17.928 ;
  LAYER M1 ;
        RECT 1.152 15.42 1.184 17.928 ;
  LAYER M1 ;
        RECT 1.216 15.42 1.248 17.928 ;
  LAYER M1 ;
        RECT 1.28 15.42 1.312 17.928 ;
  LAYER M1 ;
        RECT 1.344 15.42 1.376 17.928 ;
  LAYER M1 ;
        RECT 1.408 15.42 1.44 17.928 ;
  LAYER M1 ;
        RECT 1.472 15.42 1.504 17.928 ;
  LAYER M1 ;
        RECT 1.536 15.42 1.568 17.928 ;
  LAYER M1 ;
        RECT 1.6 15.42 1.632 17.928 ;
  LAYER M1 ;
        RECT 1.664 15.42 1.696 17.928 ;
  LAYER M1 ;
        RECT 1.728 15.42 1.76 17.928 ;
  LAYER M1 ;
        RECT 1.792 15.42 1.824 17.928 ;
  LAYER M1 ;
        RECT 1.856 15.42 1.888 17.928 ;
  LAYER M1 ;
        RECT 1.92 15.42 1.952 17.928 ;
  LAYER M1 ;
        RECT 1.984 15.42 2.016 17.928 ;
  LAYER M1 ;
        RECT 2.048 15.42 2.08 17.928 ;
  LAYER M1 ;
        RECT 2.112 15.42 2.144 17.928 ;
  LAYER M1 ;
        RECT 2.176 15.42 2.208 17.928 ;
  LAYER M1 ;
        RECT 2.24 15.42 2.272 17.928 ;
  LAYER M1 ;
        RECT 2.304 15.42 2.336 17.928 ;
  LAYER M1 ;
        RECT 2.368 15.42 2.4 17.928 ;
  LAYER M1 ;
        RECT 2.432 15.42 2.464 17.928 ;
  LAYER M1 ;
        RECT 2.496 15.42 2.528 17.928 ;
  LAYER M1 ;
        RECT 2.56 15.42 2.592 17.928 ;
  LAYER M1 ;
        RECT 2.624 15.42 2.656 17.928 ;
  LAYER M1 ;
        RECT 2.688 15.42 2.72 17.928 ;
  LAYER M2 ;
        RECT 0.364 15.504 2.836 15.536 ;
  LAYER M2 ;
        RECT 0.364 15.568 2.836 15.6 ;
  LAYER M2 ;
        RECT 0.364 15.632 2.836 15.664 ;
  LAYER M2 ;
        RECT 0.364 15.696 2.836 15.728 ;
  LAYER M2 ;
        RECT 0.364 15.76 2.836 15.792 ;
  LAYER M2 ;
        RECT 0.364 15.824 2.836 15.856 ;
  LAYER M2 ;
        RECT 0.364 15.888 2.836 15.92 ;
  LAYER M2 ;
        RECT 0.364 15.952 2.836 15.984 ;
  LAYER M2 ;
        RECT 0.364 16.016 2.836 16.048 ;
  LAYER M2 ;
        RECT 0.364 16.08 2.836 16.112 ;
  LAYER M2 ;
        RECT 0.364 16.144 2.836 16.176 ;
  LAYER M2 ;
        RECT 0.364 16.208 2.836 16.24 ;
  LAYER M2 ;
        RECT 0.364 16.272 2.836 16.304 ;
  LAYER M2 ;
        RECT 0.364 16.336 2.836 16.368 ;
  LAYER M2 ;
        RECT 0.364 16.4 2.836 16.432 ;
  LAYER M2 ;
        RECT 0.364 16.464 2.836 16.496 ;
  LAYER M2 ;
        RECT 0.364 16.528 2.836 16.56 ;
  LAYER M2 ;
        RECT 0.364 16.592 2.836 16.624 ;
  LAYER M2 ;
        RECT 0.364 16.656 2.836 16.688 ;
  LAYER M2 ;
        RECT 0.364 16.72 2.836 16.752 ;
  LAYER M2 ;
        RECT 0.364 16.784 2.836 16.816 ;
  LAYER M2 ;
        RECT 0.364 16.848 2.836 16.88 ;
  LAYER M2 ;
        RECT 0.364 16.912 2.836 16.944 ;
  LAYER M2 ;
        RECT 0.364 16.976 2.836 17.008 ;
  LAYER M2 ;
        RECT 0.364 17.04 2.836 17.072 ;
  LAYER M2 ;
        RECT 0.364 17.104 2.836 17.136 ;
  LAYER M2 ;
        RECT 0.364 17.168 2.836 17.2 ;
  LAYER M2 ;
        RECT 0.364 17.232 2.836 17.264 ;
  LAYER M2 ;
        RECT 0.364 17.296 2.836 17.328 ;
  LAYER M2 ;
        RECT 0.364 17.36 2.836 17.392 ;
  LAYER M2 ;
        RECT 0.364 17.424 2.836 17.456 ;
  LAYER M2 ;
        RECT 0.364 17.488 2.836 17.52 ;
  LAYER M2 ;
        RECT 0.364 17.552 2.836 17.584 ;
  LAYER M2 ;
        RECT 0.364 17.616 2.836 17.648 ;
  LAYER M2 ;
        RECT 0.364 17.68 2.836 17.712 ;
  LAYER M2 ;
        RECT 0.364 17.744 2.836 17.776 ;
  LAYER M3 ;
        RECT 0.384 15.42 0.416 17.928 ;
  LAYER M3 ;
        RECT 0.448 15.42 0.48 17.928 ;
  LAYER M3 ;
        RECT 0.512 15.42 0.544 17.928 ;
  LAYER M3 ;
        RECT 0.576 15.42 0.608 17.928 ;
  LAYER M3 ;
        RECT 0.64 15.42 0.672 17.928 ;
  LAYER M3 ;
        RECT 0.704 15.42 0.736 17.928 ;
  LAYER M3 ;
        RECT 0.768 15.42 0.8 17.928 ;
  LAYER M3 ;
        RECT 0.832 15.42 0.864 17.928 ;
  LAYER M3 ;
        RECT 0.896 15.42 0.928 17.928 ;
  LAYER M3 ;
        RECT 0.96 15.42 0.992 17.928 ;
  LAYER M3 ;
        RECT 1.024 15.42 1.056 17.928 ;
  LAYER M3 ;
        RECT 1.088 15.42 1.12 17.928 ;
  LAYER M3 ;
        RECT 1.152 15.42 1.184 17.928 ;
  LAYER M3 ;
        RECT 1.216 15.42 1.248 17.928 ;
  LAYER M3 ;
        RECT 1.28 15.42 1.312 17.928 ;
  LAYER M3 ;
        RECT 1.344 15.42 1.376 17.928 ;
  LAYER M3 ;
        RECT 1.408 15.42 1.44 17.928 ;
  LAYER M3 ;
        RECT 1.472 15.42 1.504 17.928 ;
  LAYER M3 ;
        RECT 1.536 15.42 1.568 17.928 ;
  LAYER M3 ;
        RECT 1.6 15.42 1.632 17.928 ;
  LAYER M3 ;
        RECT 1.664 15.42 1.696 17.928 ;
  LAYER M3 ;
        RECT 1.728 15.42 1.76 17.928 ;
  LAYER M3 ;
        RECT 1.792 15.42 1.824 17.928 ;
  LAYER M3 ;
        RECT 1.856 15.42 1.888 17.928 ;
  LAYER M3 ;
        RECT 1.92 15.42 1.952 17.928 ;
  LAYER M3 ;
        RECT 1.984 15.42 2.016 17.928 ;
  LAYER M3 ;
        RECT 2.048 15.42 2.08 17.928 ;
  LAYER M3 ;
        RECT 2.112 15.42 2.144 17.928 ;
  LAYER M3 ;
        RECT 2.176 15.42 2.208 17.928 ;
  LAYER M3 ;
        RECT 2.24 15.42 2.272 17.928 ;
  LAYER M3 ;
        RECT 2.304 15.42 2.336 17.928 ;
  LAYER M3 ;
        RECT 2.368 15.42 2.4 17.928 ;
  LAYER M3 ;
        RECT 2.432 15.42 2.464 17.928 ;
  LAYER M3 ;
        RECT 2.496 15.42 2.528 17.928 ;
  LAYER M3 ;
        RECT 2.56 15.42 2.592 17.928 ;
  LAYER M3 ;
        RECT 2.624 15.42 2.656 17.928 ;
  LAYER M3 ;
        RECT 2.688 15.42 2.72 17.928 ;
  LAYER M3 ;
        RECT 2.784 15.42 2.816 17.928 ;
  LAYER M1 ;
        RECT 0.399 15.456 0.401 17.892 ;
  LAYER M1 ;
        RECT 0.479 15.456 0.481 17.892 ;
  LAYER M1 ;
        RECT 0.559 15.456 0.561 17.892 ;
  LAYER M1 ;
        RECT 0.639 15.456 0.641 17.892 ;
  LAYER M1 ;
        RECT 0.719 15.456 0.721 17.892 ;
  LAYER M1 ;
        RECT 0.799 15.456 0.801 17.892 ;
  LAYER M1 ;
        RECT 0.879 15.456 0.881 17.892 ;
  LAYER M1 ;
        RECT 0.959 15.456 0.961 17.892 ;
  LAYER M1 ;
        RECT 1.039 15.456 1.041 17.892 ;
  LAYER M1 ;
        RECT 1.119 15.456 1.121 17.892 ;
  LAYER M1 ;
        RECT 1.199 15.456 1.201 17.892 ;
  LAYER M1 ;
        RECT 1.279 15.456 1.281 17.892 ;
  LAYER M1 ;
        RECT 1.359 15.456 1.361 17.892 ;
  LAYER M1 ;
        RECT 1.439 15.456 1.441 17.892 ;
  LAYER M1 ;
        RECT 1.519 15.456 1.521 17.892 ;
  LAYER M1 ;
        RECT 1.599 15.456 1.601 17.892 ;
  LAYER M1 ;
        RECT 1.679 15.456 1.681 17.892 ;
  LAYER M1 ;
        RECT 1.759 15.456 1.761 17.892 ;
  LAYER M1 ;
        RECT 1.839 15.456 1.841 17.892 ;
  LAYER M1 ;
        RECT 1.919 15.456 1.921 17.892 ;
  LAYER M1 ;
        RECT 1.999 15.456 2.001 17.892 ;
  LAYER M1 ;
        RECT 2.079 15.456 2.081 17.892 ;
  LAYER M1 ;
        RECT 2.159 15.456 2.161 17.892 ;
  LAYER M1 ;
        RECT 2.239 15.456 2.241 17.892 ;
  LAYER M1 ;
        RECT 2.319 15.456 2.321 17.892 ;
  LAYER M1 ;
        RECT 2.399 15.456 2.401 17.892 ;
  LAYER M1 ;
        RECT 2.479 15.456 2.481 17.892 ;
  LAYER M1 ;
        RECT 2.559 15.456 2.561 17.892 ;
  LAYER M1 ;
        RECT 2.639 15.456 2.641 17.892 ;
  LAYER M1 ;
        RECT 2.719 15.456 2.721 17.892 ;
  LAYER M2 ;
        RECT 0.4 15.455 2.8 15.457 ;
  LAYER M2 ;
        RECT 0.4 15.539 2.8 15.541 ;
  LAYER M2 ;
        RECT 0.4 15.623 2.8 15.625 ;
  LAYER M2 ;
        RECT 0.4 15.707 2.8 15.709 ;
  LAYER M2 ;
        RECT 0.4 15.791 2.8 15.793 ;
  LAYER M2 ;
        RECT 0.4 15.875 2.8 15.877 ;
  LAYER M2 ;
        RECT 0.4 15.959 2.8 15.961 ;
  LAYER M2 ;
        RECT 0.4 16.043 2.8 16.045 ;
  LAYER M2 ;
        RECT 0.4 16.127 2.8 16.129 ;
  LAYER M2 ;
        RECT 0.4 16.211 2.8 16.213 ;
  LAYER M2 ;
        RECT 0.4 16.295 2.8 16.297 ;
  LAYER M2 ;
        RECT 0.4 16.379 2.8 16.381 ;
  LAYER M2 ;
        RECT 0.4 16.4625 2.8 16.4645 ;
  LAYER M2 ;
        RECT 0.4 16.547 2.8 16.549 ;
  LAYER M2 ;
        RECT 0.4 16.631 2.8 16.633 ;
  LAYER M2 ;
        RECT 0.4 16.715 2.8 16.717 ;
  LAYER M2 ;
        RECT 0.4 16.799 2.8 16.801 ;
  LAYER M2 ;
        RECT 0.4 16.883 2.8 16.885 ;
  LAYER M2 ;
        RECT 0.4 16.967 2.8 16.969 ;
  LAYER M2 ;
        RECT 0.4 17.051 2.8 17.053 ;
  LAYER M2 ;
        RECT 0.4 17.135 2.8 17.137 ;
  LAYER M2 ;
        RECT 0.4 17.219 2.8 17.221 ;
  LAYER M2 ;
        RECT 0.4 17.303 2.8 17.305 ;
  LAYER M2 ;
        RECT 0.4 17.387 2.8 17.389 ;
  LAYER M2 ;
        RECT 0.4 17.471 2.8 17.473 ;
  LAYER M2 ;
        RECT 0.4 17.555 2.8 17.557 ;
  LAYER M2 ;
        RECT 0.4 17.639 2.8 17.641 ;
  LAYER M2 ;
        RECT 0.4 17.723 2.8 17.725 ;
  LAYER M2 ;
        RECT 0.4 17.807 2.8 17.809 ;
  LAYER M1 ;
        RECT 3.264 0.72 3.296 3.228 ;
  LAYER M1 ;
        RECT 3.328 0.72 3.36 3.228 ;
  LAYER M1 ;
        RECT 3.392 0.72 3.424 3.228 ;
  LAYER M1 ;
        RECT 3.456 0.72 3.488 3.228 ;
  LAYER M1 ;
        RECT 3.52 0.72 3.552 3.228 ;
  LAYER M1 ;
        RECT 3.584 0.72 3.616 3.228 ;
  LAYER M1 ;
        RECT 3.648 0.72 3.68 3.228 ;
  LAYER M1 ;
        RECT 3.712 0.72 3.744 3.228 ;
  LAYER M1 ;
        RECT 3.776 0.72 3.808 3.228 ;
  LAYER M1 ;
        RECT 3.84 0.72 3.872 3.228 ;
  LAYER M1 ;
        RECT 3.904 0.72 3.936 3.228 ;
  LAYER M1 ;
        RECT 3.968 0.72 4 3.228 ;
  LAYER M1 ;
        RECT 4.032 0.72 4.064 3.228 ;
  LAYER M1 ;
        RECT 4.096 0.72 4.128 3.228 ;
  LAYER M1 ;
        RECT 4.16 0.72 4.192 3.228 ;
  LAYER M1 ;
        RECT 4.224 0.72 4.256 3.228 ;
  LAYER M1 ;
        RECT 4.288 0.72 4.32 3.228 ;
  LAYER M1 ;
        RECT 4.352 0.72 4.384 3.228 ;
  LAYER M1 ;
        RECT 4.416 0.72 4.448 3.228 ;
  LAYER M1 ;
        RECT 4.48 0.72 4.512 3.228 ;
  LAYER M1 ;
        RECT 4.544 0.72 4.576 3.228 ;
  LAYER M1 ;
        RECT 4.608 0.72 4.64 3.228 ;
  LAYER M1 ;
        RECT 4.672 0.72 4.704 3.228 ;
  LAYER M1 ;
        RECT 4.736 0.72 4.768 3.228 ;
  LAYER M1 ;
        RECT 4.8 0.72 4.832 3.228 ;
  LAYER M1 ;
        RECT 4.864 0.72 4.896 3.228 ;
  LAYER M1 ;
        RECT 4.928 0.72 4.96 3.228 ;
  LAYER M1 ;
        RECT 4.992 0.72 5.024 3.228 ;
  LAYER M1 ;
        RECT 5.056 0.72 5.088 3.228 ;
  LAYER M1 ;
        RECT 5.12 0.72 5.152 3.228 ;
  LAYER M1 ;
        RECT 5.184 0.72 5.216 3.228 ;
  LAYER M1 ;
        RECT 5.248 0.72 5.28 3.228 ;
  LAYER M1 ;
        RECT 5.312 0.72 5.344 3.228 ;
  LAYER M1 ;
        RECT 5.376 0.72 5.408 3.228 ;
  LAYER M1 ;
        RECT 5.44 0.72 5.472 3.228 ;
  LAYER M1 ;
        RECT 5.504 0.72 5.536 3.228 ;
  LAYER M1 ;
        RECT 5.568 0.72 5.6 3.228 ;
  LAYER M2 ;
        RECT 3.244 0.804 5.716 0.836 ;
  LAYER M2 ;
        RECT 3.244 0.868 5.716 0.9 ;
  LAYER M2 ;
        RECT 3.244 0.932 5.716 0.964 ;
  LAYER M2 ;
        RECT 3.244 0.996 5.716 1.028 ;
  LAYER M2 ;
        RECT 3.244 1.06 5.716 1.092 ;
  LAYER M2 ;
        RECT 3.244 1.124 5.716 1.156 ;
  LAYER M2 ;
        RECT 3.244 1.188 5.716 1.22 ;
  LAYER M2 ;
        RECT 3.244 1.252 5.716 1.284 ;
  LAYER M2 ;
        RECT 3.244 1.316 5.716 1.348 ;
  LAYER M2 ;
        RECT 3.244 1.38 5.716 1.412 ;
  LAYER M2 ;
        RECT 3.244 1.444 5.716 1.476 ;
  LAYER M2 ;
        RECT 3.244 1.508 5.716 1.54 ;
  LAYER M2 ;
        RECT 3.244 1.572 5.716 1.604 ;
  LAYER M2 ;
        RECT 3.244 1.636 5.716 1.668 ;
  LAYER M2 ;
        RECT 3.244 1.7 5.716 1.732 ;
  LAYER M2 ;
        RECT 3.244 1.764 5.716 1.796 ;
  LAYER M2 ;
        RECT 3.244 1.828 5.716 1.86 ;
  LAYER M2 ;
        RECT 3.244 1.892 5.716 1.924 ;
  LAYER M2 ;
        RECT 3.244 1.956 5.716 1.988 ;
  LAYER M2 ;
        RECT 3.244 2.02 5.716 2.052 ;
  LAYER M2 ;
        RECT 3.244 2.084 5.716 2.116 ;
  LAYER M2 ;
        RECT 3.244 2.148 5.716 2.18 ;
  LAYER M2 ;
        RECT 3.244 2.212 5.716 2.244 ;
  LAYER M2 ;
        RECT 3.244 2.276 5.716 2.308 ;
  LAYER M2 ;
        RECT 3.244 2.34 5.716 2.372 ;
  LAYER M2 ;
        RECT 3.244 2.404 5.716 2.436 ;
  LAYER M2 ;
        RECT 3.244 2.468 5.716 2.5 ;
  LAYER M2 ;
        RECT 3.244 2.532 5.716 2.564 ;
  LAYER M2 ;
        RECT 3.244 2.596 5.716 2.628 ;
  LAYER M2 ;
        RECT 3.244 2.66 5.716 2.692 ;
  LAYER M2 ;
        RECT 3.244 2.724 5.716 2.756 ;
  LAYER M2 ;
        RECT 3.244 2.788 5.716 2.82 ;
  LAYER M2 ;
        RECT 3.244 2.852 5.716 2.884 ;
  LAYER M2 ;
        RECT 3.244 2.916 5.716 2.948 ;
  LAYER M2 ;
        RECT 3.244 2.98 5.716 3.012 ;
  LAYER M2 ;
        RECT 3.244 3.044 5.716 3.076 ;
  LAYER M3 ;
        RECT 3.264 0.72 3.296 3.228 ;
  LAYER M3 ;
        RECT 3.328 0.72 3.36 3.228 ;
  LAYER M3 ;
        RECT 3.392 0.72 3.424 3.228 ;
  LAYER M3 ;
        RECT 3.456 0.72 3.488 3.228 ;
  LAYER M3 ;
        RECT 3.52 0.72 3.552 3.228 ;
  LAYER M3 ;
        RECT 3.584 0.72 3.616 3.228 ;
  LAYER M3 ;
        RECT 3.648 0.72 3.68 3.228 ;
  LAYER M3 ;
        RECT 3.712 0.72 3.744 3.228 ;
  LAYER M3 ;
        RECT 3.776 0.72 3.808 3.228 ;
  LAYER M3 ;
        RECT 3.84 0.72 3.872 3.228 ;
  LAYER M3 ;
        RECT 3.904 0.72 3.936 3.228 ;
  LAYER M3 ;
        RECT 3.968 0.72 4 3.228 ;
  LAYER M3 ;
        RECT 4.032 0.72 4.064 3.228 ;
  LAYER M3 ;
        RECT 4.096 0.72 4.128 3.228 ;
  LAYER M3 ;
        RECT 4.16 0.72 4.192 3.228 ;
  LAYER M3 ;
        RECT 4.224 0.72 4.256 3.228 ;
  LAYER M3 ;
        RECT 4.288 0.72 4.32 3.228 ;
  LAYER M3 ;
        RECT 4.352 0.72 4.384 3.228 ;
  LAYER M3 ;
        RECT 4.416 0.72 4.448 3.228 ;
  LAYER M3 ;
        RECT 4.48 0.72 4.512 3.228 ;
  LAYER M3 ;
        RECT 4.544 0.72 4.576 3.228 ;
  LAYER M3 ;
        RECT 4.608 0.72 4.64 3.228 ;
  LAYER M3 ;
        RECT 4.672 0.72 4.704 3.228 ;
  LAYER M3 ;
        RECT 4.736 0.72 4.768 3.228 ;
  LAYER M3 ;
        RECT 4.8 0.72 4.832 3.228 ;
  LAYER M3 ;
        RECT 4.864 0.72 4.896 3.228 ;
  LAYER M3 ;
        RECT 4.928 0.72 4.96 3.228 ;
  LAYER M3 ;
        RECT 4.992 0.72 5.024 3.228 ;
  LAYER M3 ;
        RECT 5.056 0.72 5.088 3.228 ;
  LAYER M3 ;
        RECT 5.12 0.72 5.152 3.228 ;
  LAYER M3 ;
        RECT 5.184 0.72 5.216 3.228 ;
  LAYER M3 ;
        RECT 5.248 0.72 5.28 3.228 ;
  LAYER M3 ;
        RECT 5.312 0.72 5.344 3.228 ;
  LAYER M3 ;
        RECT 5.376 0.72 5.408 3.228 ;
  LAYER M3 ;
        RECT 5.44 0.72 5.472 3.228 ;
  LAYER M3 ;
        RECT 5.504 0.72 5.536 3.228 ;
  LAYER M3 ;
        RECT 5.568 0.72 5.6 3.228 ;
  LAYER M3 ;
        RECT 5.664 0.72 5.696 3.228 ;
  LAYER M1 ;
        RECT 3.279 0.756 3.281 3.192 ;
  LAYER M1 ;
        RECT 3.359 0.756 3.361 3.192 ;
  LAYER M1 ;
        RECT 3.439 0.756 3.441 3.192 ;
  LAYER M1 ;
        RECT 3.519 0.756 3.521 3.192 ;
  LAYER M1 ;
        RECT 3.599 0.756 3.601 3.192 ;
  LAYER M1 ;
        RECT 3.679 0.756 3.681 3.192 ;
  LAYER M1 ;
        RECT 3.759 0.756 3.761 3.192 ;
  LAYER M1 ;
        RECT 3.839 0.756 3.841 3.192 ;
  LAYER M1 ;
        RECT 3.919 0.756 3.921 3.192 ;
  LAYER M1 ;
        RECT 3.999 0.756 4.001 3.192 ;
  LAYER M1 ;
        RECT 4.079 0.756 4.081 3.192 ;
  LAYER M1 ;
        RECT 4.159 0.756 4.161 3.192 ;
  LAYER M1 ;
        RECT 4.239 0.756 4.241 3.192 ;
  LAYER M1 ;
        RECT 4.319 0.756 4.321 3.192 ;
  LAYER M1 ;
        RECT 4.399 0.756 4.401 3.192 ;
  LAYER M1 ;
        RECT 4.479 0.756 4.481 3.192 ;
  LAYER M1 ;
        RECT 4.559 0.756 4.561 3.192 ;
  LAYER M1 ;
        RECT 4.639 0.756 4.641 3.192 ;
  LAYER M1 ;
        RECT 4.719 0.756 4.721 3.192 ;
  LAYER M1 ;
        RECT 4.799 0.756 4.801 3.192 ;
  LAYER M1 ;
        RECT 4.879 0.756 4.881 3.192 ;
  LAYER M1 ;
        RECT 4.959 0.756 4.961 3.192 ;
  LAYER M1 ;
        RECT 5.039 0.756 5.041 3.192 ;
  LAYER M1 ;
        RECT 5.119 0.756 5.121 3.192 ;
  LAYER M1 ;
        RECT 5.199 0.756 5.201 3.192 ;
  LAYER M1 ;
        RECT 5.279 0.756 5.281 3.192 ;
  LAYER M1 ;
        RECT 5.359 0.756 5.361 3.192 ;
  LAYER M1 ;
        RECT 5.439 0.756 5.441 3.192 ;
  LAYER M1 ;
        RECT 5.519 0.756 5.521 3.192 ;
  LAYER M1 ;
        RECT 5.599 0.756 5.601 3.192 ;
  LAYER M2 ;
        RECT 3.28 0.755 5.68 0.757 ;
  LAYER M2 ;
        RECT 3.28 0.839 5.68 0.841 ;
  LAYER M2 ;
        RECT 3.28 0.923 5.68 0.925 ;
  LAYER M2 ;
        RECT 3.28 1.007 5.68 1.009 ;
  LAYER M2 ;
        RECT 3.28 1.091 5.68 1.093 ;
  LAYER M2 ;
        RECT 3.28 1.175 5.68 1.177 ;
  LAYER M2 ;
        RECT 3.28 1.259 5.68 1.261 ;
  LAYER M2 ;
        RECT 3.28 1.343 5.68 1.345 ;
  LAYER M2 ;
        RECT 3.28 1.427 5.68 1.429 ;
  LAYER M2 ;
        RECT 3.28 1.511 5.68 1.513 ;
  LAYER M2 ;
        RECT 3.28 1.595 5.68 1.597 ;
  LAYER M2 ;
        RECT 3.28 1.679 5.68 1.681 ;
  LAYER M2 ;
        RECT 3.28 1.7625 5.68 1.7645 ;
  LAYER M2 ;
        RECT 3.28 1.847 5.68 1.849 ;
  LAYER M2 ;
        RECT 3.28 1.931 5.68 1.933 ;
  LAYER M2 ;
        RECT 3.28 2.015 5.68 2.017 ;
  LAYER M2 ;
        RECT 3.28 2.099 5.68 2.101 ;
  LAYER M2 ;
        RECT 3.28 2.183 5.68 2.185 ;
  LAYER M2 ;
        RECT 3.28 2.267 5.68 2.269 ;
  LAYER M2 ;
        RECT 3.28 2.351 5.68 2.353 ;
  LAYER M2 ;
        RECT 3.28 2.435 5.68 2.437 ;
  LAYER M2 ;
        RECT 3.28 2.519 5.68 2.521 ;
  LAYER M2 ;
        RECT 3.28 2.603 5.68 2.605 ;
  LAYER M2 ;
        RECT 3.28 2.687 5.68 2.689 ;
  LAYER M2 ;
        RECT 3.28 2.771 5.68 2.773 ;
  LAYER M2 ;
        RECT 3.28 2.855 5.68 2.857 ;
  LAYER M2 ;
        RECT 3.28 2.939 5.68 2.941 ;
  LAYER M2 ;
        RECT 3.28 3.023 5.68 3.025 ;
  LAYER M2 ;
        RECT 3.28 3.107 5.68 3.109 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 6.168 ;
  LAYER M1 ;
        RECT 3.328 3.66 3.36 6.168 ;
  LAYER M1 ;
        RECT 3.392 3.66 3.424 6.168 ;
  LAYER M1 ;
        RECT 3.456 3.66 3.488 6.168 ;
  LAYER M1 ;
        RECT 3.52 3.66 3.552 6.168 ;
  LAYER M1 ;
        RECT 3.584 3.66 3.616 6.168 ;
  LAYER M1 ;
        RECT 3.648 3.66 3.68 6.168 ;
  LAYER M1 ;
        RECT 3.712 3.66 3.744 6.168 ;
  LAYER M1 ;
        RECT 3.776 3.66 3.808 6.168 ;
  LAYER M1 ;
        RECT 3.84 3.66 3.872 6.168 ;
  LAYER M1 ;
        RECT 3.904 3.66 3.936 6.168 ;
  LAYER M1 ;
        RECT 3.968 3.66 4 6.168 ;
  LAYER M1 ;
        RECT 4.032 3.66 4.064 6.168 ;
  LAYER M1 ;
        RECT 4.096 3.66 4.128 6.168 ;
  LAYER M1 ;
        RECT 4.16 3.66 4.192 6.168 ;
  LAYER M1 ;
        RECT 4.224 3.66 4.256 6.168 ;
  LAYER M1 ;
        RECT 4.288 3.66 4.32 6.168 ;
  LAYER M1 ;
        RECT 4.352 3.66 4.384 6.168 ;
  LAYER M1 ;
        RECT 4.416 3.66 4.448 6.168 ;
  LAYER M1 ;
        RECT 4.48 3.66 4.512 6.168 ;
  LAYER M1 ;
        RECT 4.544 3.66 4.576 6.168 ;
  LAYER M1 ;
        RECT 4.608 3.66 4.64 6.168 ;
  LAYER M1 ;
        RECT 4.672 3.66 4.704 6.168 ;
  LAYER M1 ;
        RECT 4.736 3.66 4.768 6.168 ;
  LAYER M1 ;
        RECT 4.8 3.66 4.832 6.168 ;
  LAYER M1 ;
        RECT 4.864 3.66 4.896 6.168 ;
  LAYER M1 ;
        RECT 4.928 3.66 4.96 6.168 ;
  LAYER M1 ;
        RECT 4.992 3.66 5.024 6.168 ;
  LAYER M1 ;
        RECT 5.056 3.66 5.088 6.168 ;
  LAYER M1 ;
        RECT 5.12 3.66 5.152 6.168 ;
  LAYER M1 ;
        RECT 5.184 3.66 5.216 6.168 ;
  LAYER M1 ;
        RECT 5.248 3.66 5.28 6.168 ;
  LAYER M1 ;
        RECT 5.312 3.66 5.344 6.168 ;
  LAYER M1 ;
        RECT 5.376 3.66 5.408 6.168 ;
  LAYER M1 ;
        RECT 5.44 3.66 5.472 6.168 ;
  LAYER M1 ;
        RECT 5.504 3.66 5.536 6.168 ;
  LAYER M1 ;
        RECT 5.568 3.66 5.6 6.168 ;
  LAYER M2 ;
        RECT 3.244 3.744 5.716 3.776 ;
  LAYER M2 ;
        RECT 3.244 3.808 5.716 3.84 ;
  LAYER M2 ;
        RECT 3.244 3.872 5.716 3.904 ;
  LAYER M2 ;
        RECT 3.244 3.936 5.716 3.968 ;
  LAYER M2 ;
        RECT 3.244 4 5.716 4.032 ;
  LAYER M2 ;
        RECT 3.244 4.064 5.716 4.096 ;
  LAYER M2 ;
        RECT 3.244 4.128 5.716 4.16 ;
  LAYER M2 ;
        RECT 3.244 4.192 5.716 4.224 ;
  LAYER M2 ;
        RECT 3.244 4.256 5.716 4.288 ;
  LAYER M2 ;
        RECT 3.244 4.32 5.716 4.352 ;
  LAYER M2 ;
        RECT 3.244 4.384 5.716 4.416 ;
  LAYER M2 ;
        RECT 3.244 4.448 5.716 4.48 ;
  LAYER M2 ;
        RECT 3.244 4.512 5.716 4.544 ;
  LAYER M2 ;
        RECT 3.244 4.576 5.716 4.608 ;
  LAYER M2 ;
        RECT 3.244 4.64 5.716 4.672 ;
  LAYER M2 ;
        RECT 3.244 4.704 5.716 4.736 ;
  LAYER M2 ;
        RECT 3.244 4.768 5.716 4.8 ;
  LAYER M2 ;
        RECT 3.244 4.832 5.716 4.864 ;
  LAYER M2 ;
        RECT 3.244 4.896 5.716 4.928 ;
  LAYER M2 ;
        RECT 3.244 4.96 5.716 4.992 ;
  LAYER M2 ;
        RECT 3.244 5.024 5.716 5.056 ;
  LAYER M2 ;
        RECT 3.244 5.088 5.716 5.12 ;
  LAYER M2 ;
        RECT 3.244 5.152 5.716 5.184 ;
  LAYER M2 ;
        RECT 3.244 5.216 5.716 5.248 ;
  LAYER M2 ;
        RECT 3.244 5.28 5.716 5.312 ;
  LAYER M2 ;
        RECT 3.244 5.344 5.716 5.376 ;
  LAYER M2 ;
        RECT 3.244 5.408 5.716 5.44 ;
  LAYER M2 ;
        RECT 3.244 5.472 5.716 5.504 ;
  LAYER M2 ;
        RECT 3.244 5.536 5.716 5.568 ;
  LAYER M2 ;
        RECT 3.244 5.6 5.716 5.632 ;
  LAYER M2 ;
        RECT 3.244 5.664 5.716 5.696 ;
  LAYER M2 ;
        RECT 3.244 5.728 5.716 5.76 ;
  LAYER M2 ;
        RECT 3.244 5.792 5.716 5.824 ;
  LAYER M2 ;
        RECT 3.244 5.856 5.716 5.888 ;
  LAYER M2 ;
        RECT 3.244 5.92 5.716 5.952 ;
  LAYER M2 ;
        RECT 3.244 5.984 5.716 6.016 ;
  LAYER M3 ;
        RECT 3.264 3.66 3.296 6.168 ;
  LAYER M3 ;
        RECT 3.328 3.66 3.36 6.168 ;
  LAYER M3 ;
        RECT 3.392 3.66 3.424 6.168 ;
  LAYER M3 ;
        RECT 3.456 3.66 3.488 6.168 ;
  LAYER M3 ;
        RECT 3.52 3.66 3.552 6.168 ;
  LAYER M3 ;
        RECT 3.584 3.66 3.616 6.168 ;
  LAYER M3 ;
        RECT 3.648 3.66 3.68 6.168 ;
  LAYER M3 ;
        RECT 3.712 3.66 3.744 6.168 ;
  LAYER M3 ;
        RECT 3.776 3.66 3.808 6.168 ;
  LAYER M3 ;
        RECT 3.84 3.66 3.872 6.168 ;
  LAYER M3 ;
        RECT 3.904 3.66 3.936 6.168 ;
  LAYER M3 ;
        RECT 3.968 3.66 4 6.168 ;
  LAYER M3 ;
        RECT 4.032 3.66 4.064 6.168 ;
  LAYER M3 ;
        RECT 4.096 3.66 4.128 6.168 ;
  LAYER M3 ;
        RECT 4.16 3.66 4.192 6.168 ;
  LAYER M3 ;
        RECT 4.224 3.66 4.256 6.168 ;
  LAYER M3 ;
        RECT 4.288 3.66 4.32 6.168 ;
  LAYER M3 ;
        RECT 4.352 3.66 4.384 6.168 ;
  LAYER M3 ;
        RECT 4.416 3.66 4.448 6.168 ;
  LAYER M3 ;
        RECT 4.48 3.66 4.512 6.168 ;
  LAYER M3 ;
        RECT 4.544 3.66 4.576 6.168 ;
  LAYER M3 ;
        RECT 4.608 3.66 4.64 6.168 ;
  LAYER M3 ;
        RECT 4.672 3.66 4.704 6.168 ;
  LAYER M3 ;
        RECT 4.736 3.66 4.768 6.168 ;
  LAYER M3 ;
        RECT 4.8 3.66 4.832 6.168 ;
  LAYER M3 ;
        RECT 4.864 3.66 4.896 6.168 ;
  LAYER M3 ;
        RECT 4.928 3.66 4.96 6.168 ;
  LAYER M3 ;
        RECT 4.992 3.66 5.024 6.168 ;
  LAYER M3 ;
        RECT 5.056 3.66 5.088 6.168 ;
  LAYER M3 ;
        RECT 5.12 3.66 5.152 6.168 ;
  LAYER M3 ;
        RECT 5.184 3.66 5.216 6.168 ;
  LAYER M3 ;
        RECT 5.248 3.66 5.28 6.168 ;
  LAYER M3 ;
        RECT 5.312 3.66 5.344 6.168 ;
  LAYER M3 ;
        RECT 5.376 3.66 5.408 6.168 ;
  LAYER M3 ;
        RECT 5.44 3.66 5.472 6.168 ;
  LAYER M3 ;
        RECT 5.504 3.66 5.536 6.168 ;
  LAYER M3 ;
        RECT 5.568 3.66 5.6 6.168 ;
  LAYER M3 ;
        RECT 5.664 3.66 5.696 6.168 ;
  LAYER M1 ;
        RECT 3.279 3.696 3.281 6.132 ;
  LAYER M1 ;
        RECT 3.359 3.696 3.361 6.132 ;
  LAYER M1 ;
        RECT 3.439 3.696 3.441 6.132 ;
  LAYER M1 ;
        RECT 3.519 3.696 3.521 6.132 ;
  LAYER M1 ;
        RECT 3.599 3.696 3.601 6.132 ;
  LAYER M1 ;
        RECT 3.679 3.696 3.681 6.132 ;
  LAYER M1 ;
        RECT 3.759 3.696 3.761 6.132 ;
  LAYER M1 ;
        RECT 3.839 3.696 3.841 6.132 ;
  LAYER M1 ;
        RECT 3.919 3.696 3.921 6.132 ;
  LAYER M1 ;
        RECT 3.999 3.696 4.001 6.132 ;
  LAYER M1 ;
        RECT 4.079 3.696 4.081 6.132 ;
  LAYER M1 ;
        RECT 4.159 3.696 4.161 6.132 ;
  LAYER M1 ;
        RECT 4.239 3.696 4.241 6.132 ;
  LAYER M1 ;
        RECT 4.319 3.696 4.321 6.132 ;
  LAYER M1 ;
        RECT 4.399 3.696 4.401 6.132 ;
  LAYER M1 ;
        RECT 4.479 3.696 4.481 6.132 ;
  LAYER M1 ;
        RECT 4.559 3.696 4.561 6.132 ;
  LAYER M1 ;
        RECT 4.639 3.696 4.641 6.132 ;
  LAYER M1 ;
        RECT 4.719 3.696 4.721 6.132 ;
  LAYER M1 ;
        RECT 4.799 3.696 4.801 6.132 ;
  LAYER M1 ;
        RECT 4.879 3.696 4.881 6.132 ;
  LAYER M1 ;
        RECT 4.959 3.696 4.961 6.132 ;
  LAYER M1 ;
        RECT 5.039 3.696 5.041 6.132 ;
  LAYER M1 ;
        RECT 5.119 3.696 5.121 6.132 ;
  LAYER M1 ;
        RECT 5.199 3.696 5.201 6.132 ;
  LAYER M1 ;
        RECT 5.279 3.696 5.281 6.132 ;
  LAYER M1 ;
        RECT 5.359 3.696 5.361 6.132 ;
  LAYER M1 ;
        RECT 5.439 3.696 5.441 6.132 ;
  LAYER M1 ;
        RECT 5.519 3.696 5.521 6.132 ;
  LAYER M1 ;
        RECT 5.599 3.696 5.601 6.132 ;
  LAYER M2 ;
        RECT 3.28 3.695 5.68 3.697 ;
  LAYER M2 ;
        RECT 3.28 3.779 5.68 3.781 ;
  LAYER M2 ;
        RECT 3.28 3.863 5.68 3.865 ;
  LAYER M2 ;
        RECT 3.28 3.947 5.68 3.949 ;
  LAYER M2 ;
        RECT 3.28 4.031 5.68 4.033 ;
  LAYER M2 ;
        RECT 3.28 4.115 5.68 4.117 ;
  LAYER M2 ;
        RECT 3.28 4.199 5.68 4.201 ;
  LAYER M2 ;
        RECT 3.28 4.283 5.68 4.285 ;
  LAYER M2 ;
        RECT 3.28 4.367 5.68 4.369 ;
  LAYER M2 ;
        RECT 3.28 4.451 5.68 4.453 ;
  LAYER M2 ;
        RECT 3.28 4.535 5.68 4.537 ;
  LAYER M2 ;
        RECT 3.28 4.619 5.68 4.621 ;
  LAYER M2 ;
        RECT 3.28 4.7025 5.68 4.7045 ;
  LAYER M2 ;
        RECT 3.28 4.787 5.68 4.789 ;
  LAYER M2 ;
        RECT 3.28 4.871 5.68 4.873 ;
  LAYER M2 ;
        RECT 3.28 4.955 5.68 4.957 ;
  LAYER M2 ;
        RECT 3.28 5.039 5.68 5.041 ;
  LAYER M2 ;
        RECT 3.28 5.123 5.68 5.125 ;
  LAYER M2 ;
        RECT 3.28 5.207 5.68 5.209 ;
  LAYER M2 ;
        RECT 3.28 5.291 5.68 5.293 ;
  LAYER M2 ;
        RECT 3.28 5.375 5.68 5.377 ;
  LAYER M2 ;
        RECT 3.28 5.459 5.68 5.461 ;
  LAYER M2 ;
        RECT 3.28 5.543 5.68 5.545 ;
  LAYER M2 ;
        RECT 3.28 5.627 5.68 5.629 ;
  LAYER M2 ;
        RECT 3.28 5.711 5.68 5.713 ;
  LAYER M2 ;
        RECT 3.28 5.795 5.68 5.797 ;
  LAYER M2 ;
        RECT 3.28 5.879 5.68 5.881 ;
  LAYER M2 ;
        RECT 3.28 5.963 5.68 5.965 ;
  LAYER M2 ;
        RECT 3.28 6.047 5.68 6.049 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 9.108 ;
  LAYER M1 ;
        RECT 3.328 6.6 3.36 9.108 ;
  LAYER M1 ;
        RECT 3.392 6.6 3.424 9.108 ;
  LAYER M1 ;
        RECT 3.456 6.6 3.488 9.108 ;
  LAYER M1 ;
        RECT 3.52 6.6 3.552 9.108 ;
  LAYER M1 ;
        RECT 3.584 6.6 3.616 9.108 ;
  LAYER M1 ;
        RECT 3.648 6.6 3.68 9.108 ;
  LAYER M1 ;
        RECT 3.712 6.6 3.744 9.108 ;
  LAYER M1 ;
        RECT 3.776 6.6 3.808 9.108 ;
  LAYER M1 ;
        RECT 3.84 6.6 3.872 9.108 ;
  LAYER M1 ;
        RECT 3.904 6.6 3.936 9.108 ;
  LAYER M1 ;
        RECT 3.968 6.6 4 9.108 ;
  LAYER M1 ;
        RECT 4.032 6.6 4.064 9.108 ;
  LAYER M1 ;
        RECT 4.096 6.6 4.128 9.108 ;
  LAYER M1 ;
        RECT 4.16 6.6 4.192 9.108 ;
  LAYER M1 ;
        RECT 4.224 6.6 4.256 9.108 ;
  LAYER M1 ;
        RECT 4.288 6.6 4.32 9.108 ;
  LAYER M1 ;
        RECT 4.352 6.6 4.384 9.108 ;
  LAYER M1 ;
        RECT 4.416 6.6 4.448 9.108 ;
  LAYER M1 ;
        RECT 4.48 6.6 4.512 9.108 ;
  LAYER M1 ;
        RECT 4.544 6.6 4.576 9.108 ;
  LAYER M1 ;
        RECT 4.608 6.6 4.64 9.108 ;
  LAYER M1 ;
        RECT 4.672 6.6 4.704 9.108 ;
  LAYER M1 ;
        RECT 4.736 6.6 4.768 9.108 ;
  LAYER M1 ;
        RECT 4.8 6.6 4.832 9.108 ;
  LAYER M1 ;
        RECT 4.864 6.6 4.896 9.108 ;
  LAYER M1 ;
        RECT 4.928 6.6 4.96 9.108 ;
  LAYER M1 ;
        RECT 4.992 6.6 5.024 9.108 ;
  LAYER M1 ;
        RECT 5.056 6.6 5.088 9.108 ;
  LAYER M1 ;
        RECT 5.12 6.6 5.152 9.108 ;
  LAYER M1 ;
        RECT 5.184 6.6 5.216 9.108 ;
  LAYER M1 ;
        RECT 5.248 6.6 5.28 9.108 ;
  LAYER M1 ;
        RECT 5.312 6.6 5.344 9.108 ;
  LAYER M1 ;
        RECT 5.376 6.6 5.408 9.108 ;
  LAYER M1 ;
        RECT 5.44 6.6 5.472 9.108 ;
  LAYER M1 ;
        RECT 5.504 6.6 5.536 9.108 ;
  LAYER M1 ;
        RECT 5.568 6.6 5.6 9.108 ;
  LAYER M2 ;
        RECT 3.244 6.684 5.716 6.716 ;
  LAYER M2 ;
        RECT 3.244 6.748 5.716 6.78 ;
  LAYER M2 ;
        RECT 3.244 6.812 5.716 6.844 ;
  LAYER M2 ;
        RECT 3.244 6.876 5.716 6.908 ;
  LAYER M2 ;
        RECT 3.244 6.94 5.716 6.972 ;
  LAYER M2 ;
        RECT 3.244 7.004 5.716 7.036 ;
  LAYER M2 ;
        RECT 3.244 7.068 5.716 7.1 ;
  LAYER M2 ;
        RECT 3.244 7.132 5.716 7.164 ;
  LAYER M2 ;
        RECT 3.244 7.196 5.716 7.228 ;
  LAYER M2 ;
        RECT 3.244 7.26 5.716 7.292 ;
  LAYER M2 ;
        RECT 3.244 7.324 5.716 7.356 ;
  LAYER M2 ;
        RECT 3.244 7.388 5.716 7.42 ;
  LAYER M2 ;
        RECT 3.244 7.452 5.716 7.484 ;
  LAYER M2 ;
        RECT 3.244 7.516 5.716 7.548 ;
  LAYER M2 ;
        RECT 3.244 7.58 5.716 7.612 ;
  LAYER M2 ;
        RECT 3.244 7.644 5.716 7.676 ;
  LAYER M2 ;
        RECT 3.244 7.708 5.716 7.74 ;
  LAYER M2 ;
        RECT 3.244 7.772 5.716 7.804 ;
  LAYER M2 ;
        RECT 3.244 7.836 5.716 7.868 ;
  LAYER M2 ;
        RECT 3.244 7.9 5.716 7.932 ;
  LAYER M2 ;
        RECT 3.244 7.964 5.716 7.996 ;
  LAYER M2 ;
        RECT 3.244 8.028 5.716 8.06 ;
  LAYER M2 ;
        RECT 3.244 8.092 5.716 8.124 ;
  LAYER M2 ;
        RECT 3.244 8.156 5.716 8.188 ;
  LAYER M2 ;
        RECT 3.244 8.22 5.716 8.252 ;
  LAYER M2 ;
        RECT 3.244 8.284 5.716 8.316 ;
  LAYER M2 ;
        RECT 3.244 8.348 5.716 8.38 ;
  LAYER M2 ;
        RECT 3.244 8.412 5.716 8.444 ;
  LAYER M2 ;
        RECT 3.244 8.476 5.716 8.508 ;
  LAYER M2 ;
        RECT 3.244 8.54 5.716 8.572 ;
  LAYER M2 ;
        RECT 3.244 8.604 5.716 8.636 ;
  LAYER M2 ;
        RECT 3.244 8.668 5.716 8.7 ;
  LAYER M2 ;
        RECT 3.244 8.732 5.716 8.764 ;
  LAYER M2 ;
        RECT 3.244 8.796 5.716 8.828 ;
  LAYER M2 ;
        RECT 3.244 8.86 5.716 8.892 ;
  LAYER M2 ;
        RECT 3.244 8.924 5.716 8.956 ;
  LAYER M3 ;
        RECT 3.264 6.6 3.296 9.108 ;
  LAYER M3 ;
        RECT 3.328 6.6 3.36 9.108 ;
  LAYER M3 ;
        RECT 3.392 6.6 3.424 9.108 ;
  LAYER M3 ;
        RECT 3.456 6.6 3.488 9.108 ;
  LAYER M3 ;
        RECT 3.52 6.6 3.552 9.108 ;
  LAYER M3 ;
        RECT 3.584 6.6 3.616 9.108 ;
  LAYER M3 ;
        RECT 3.648 6.6 3.68 9.108 ;
  LAYER M3 ;
        RECT 3.712 6.6 3.744 9.108 ;
  LAYER M3 ;
        RECT 3.776 6.6 3.808 9.108 ;
  LAYER M3 ;
        RECT 3.84 6.6 3.872 9.108 ;
  LAYER M3 ;
        RECT 3.904 6.6 3.936 9.108 ;
  LAYER M3 ;
        RECT 3.968 6.6 4 9.108 ;
  LAYER M3 ;
        RECT 4.032 6.6 4.064 9.108 ;
  LAYER M3 ;
        RECT 4.096 6.6 4.128 9.108 ;
  LAYER M3 ;
        RECT 4.16 6.6 4.192 9.108 ;
  LAYER M3 ;
        RECT 4.224 6.6 4.256 9.108 ;
  LAYER M3 ;
        RECT 4.288 6.6 4.32 9.108 ;
  LAYER M3 ;
        RECT 4.352 6.6 4.384 9.108 ;
  LAYER M3 ;
        RECT 4.416 6.6 4.448 9.108 ;
  LAYER M3 ;
        RECT 4.48 6.6 4.512 9.108 ;
  LAYER M3 ;
        RECT 4.544 6.6 4.576 9.108 ;
  LAYER M3 ;
        RECT 4.608 6.6 4.64 9.108 ;
  LAYER M3 ;
        RECT 4.672 6.6 4.704 9.108 ;
  LAYER M3 ;
        RECT 4.736 6.6 4.768 9.108 ;
  LAYER M3 ;
        RECT 4.8 6.6 4.832 9.108 ;
  LAYER M3 ;
        RECT 4.864 6.6 4.896 9.108 ;
  LAYER M3 ;
        RECT 4.928 6.6 4.96 9.108 ;
  LAYER M3 ;
        RECT 4.992 6.6 5.024 9.108 ;
  LAYER M3 ;
        RECT 5.056 6.6 5.088 9.108 ;
  LAYER M3 ;
        RECT 5.12 6.6 5.152 9.108 ;
  LAYER M3 ;
        RECT 5.184 6.6 5.216 9.108 ;
  LAYER M3 ;
        RECT 5.248 6.6 5.28 9.108 ;
  LAYER M3 ;
        RECT 5.312 6.6 5.344 9.108 ;
  LAYER M3 ;
        RECT 5.376 6.6 5.408 9.108 ;
  LAYER M3 ;
        RECT 5.44 6.6 5.472 9.108 ;
  LAYER M3 ;
        RECT 5.504 6.6 5.536 9.108 ;
  LAYER M3 ;
        RECT 5.568 6.6 5.6 9.108 ;
  LAYER M3 ;
        RECT 5.664 6.6 5.696 9.108 ;
  LAYER M1 ;
        RECT 3.279 6.636 3.281 9.072 ;
  LAYER M1 ;
        RECT 3.359 6.636 3.361 9.072 ;
  LAYER M1 ;
        RECT 3.439 6.636 3.441 9.072 ;
  LAYER M1 ;
        RECT 3.519 6.636 3.521 9.072 ;
  LAYER M1 ;
        RECT 3.599 6.636 3.601 9.072 ;
  LAYER M1 ;
        RECT 3.679 6.636 3.681 9.072 ;
  LAYER M1 ;
        RECT 3.759 6.636 3.761 9.072 ;
  LAYER M1 ;
        RECT 3.839 6.636 3.841 9.072 ;
  LAYER M1 ;
        RECT 3.919 6.636 3.921 9.072 ;
  LAYER M1 ;
        RECT 3.999 6.636 4.001 9.072 ;
  LAYER M1 ;
        RECT 4.079 6.636 4.081 9.072 ;
  LAYER M1 ;
        RECT 4.159 6.636 4.161 9.072 ;
  LAYER M1 ;
        RECT 4.239 6.636 4.241 9.072 ;
  LAYER M1 ;
        RECT 4.319 6.636 4.321 9.072 ;
  LAYER M1 ;
        RECT 4.399 6.636 4.401 9.072 ;
  LAYER M1 ;
        RECT 4.479 6.636 4.481 9.072 ;
  LAYER M1 ;
        RECT 4.559 6.636 4.561 9.072 ;
  LAYER M1 ;
        RECT 4.639 6.636 4.641 9.072 ;
  LAYER M1 ;
        RECT 4.719 6.636 4.721 9.072 ;
  LAYER M1 ;
        RECT 4.799 6.636 4.801 9.072 ;
  LAYER M1 ;
        RECT 4.879 6.636 4.881 9.072 ;
  LAYER M1 ;
        RECT 4.959 6.636 4.961 9.072 ;
  LAYER M1 ;
        RECT 5.039 6.636 5.041 9.072 ;
  LAYER M1 ;
        RECT 5.119 6.636 5.121 9.072 ;
  LAYER M1 ;
        RECT 5.199 6.636 5.201 9.072 ;
  LAYER M1 ;
        RECT 5.279 6.636 5.281 9.072 ;
  LAYER M1 ;
        RECT 5.359 6.636 5.361 9.072 ;
  LAYER M1 ;
        RECT 5.439 6.636 5.441 9.072 ;
  LAYER M1 ;
        RECT 5.519 6.636 5.521 9.072 ;
  LAYER M1 ;
        RECT 5.599 6.636 5.601 9.072 ;
  LAYER M2 ;
        RECT 3.28 6.635 5.68 6.637 ;
  LAYER M2 ;
        RECT 3.28 6.719 5.68 6.721 ;
  LAYER M2 ;
        RECT 3.28 6.803 5.68 6.805 ;
  LAYER M2 ;
        RECT 3.28 6.887 5.68 6.889 ;
  LAYER M2 ;
        RECT 3.28 6.971 5.68 6.973 ;
  LAYER M2 ;
        RECT 3.28 7.055 5.68 7.057 ;
  LAYER M2 ;
        RECT 3.28 7.139 5.68 7.141 ;
  LAYER M2 ;
        RECT 3.28 7.223 5.68 7.225 ;
  LAYER M2 ;
        RECT 3.28 7.307 5.68 7.309 ;
  LAYER M2 ;
        RECT 3.28 7.391 5.68 7.393 ;
  LAYER M2 ;
        RECT 3.28 7.475 5.68 7.477 ;
  LAYER M2 ;
        RECT 3.28 7.559 5.68 7.561 ;
  LAYER M2 ;
        RECT 3.28 7.6425 5.68 7.6445 ;
  LAYER M2 ;
        RECT 3.28 7.727 5.68 7.729 ;
  LAYER M2 ;
        RECT 3.28 7.811 5.68 7.813 ;
  LAYER M2 ;
        RECT 3.28 7.895 5.68 7.897 ;
  LAYER M2 ;
        RECT 3.28 7.979 5.68 7.981 ;
  LAYER M2 ;
        RECT 3.28 8.063 5.68 8.065 ;
  LAYER M2 ;
        RECT 3.28 8.147 5.68 8.149 ;
  LAYER M2 ;
        RECT 3.28 8.231 5.68 8.233 ;
  LAYER M2 ;
        RECT 3.28 8.315 5.68 8.317 ;
  LAYER M2 ;
        RECT 3.28 8.399 5.68 8.401 ;
  LAYER M2 ;
        RECT 3.28 8.483 5.68 8.485 ;
  LAYER M2 ;
        RECT 3.28 8.567 5.68 8.569 ;
  LAYER M2 ;
        RECT 3.28 8.651 5.68 8.653 ;
  LAYER M2 ;
        RECT 3.28 8.735 5.68 8.737 ;
  LAYER M2 ;
        RECT 3.28 8.819 5.68 8.821 ;
  LAYER M2 ;
        RECT 3.28 8.903 5.68 8.905 ;
  LAYER M2 ;
        RECT 3.28 8.987 5.68 8.989 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 12.048 ;
  LAYER M1 ;
        RECT 3.328 9.54 3.36 12.048 ;
  LAYER M1 ;
        RECT 3.392 9.54 3.424 12.048 ;
  LAYER M1 ;
        RECT 3.456 9.54 3.488 12.048 ;
  LAYER M1 ;
        RECT 3.52 9.54 3.552 12.048 ;
  LAYER M1 ;
        RECT 3.584 9.54 3.616 12.048 ;
  LAYER M1 ;
        RECT 3.648 9.54 3.68 12.048 ;
  LAYER M1 ;
        RECT 3.712 9.54 3.744 12.048 ;
  LAYER M1 ;
        RECT 3.776 9.54 3.808 12.048 ;
  LAYER M1 ;
        RECT 3.84 9.54 3.872 12.048 ;
  LAYER M1 ;
        RECT 3.904 9.54 3.936 12.048 ;
  LAYER M1 ;
        RECT 3.968 9.54 4 12.048 ;
  LAYER M1 ;
        RECT 4.032 9.54 4.064 12.048 ;
  LAYER M1 ;
        RECT 4.096 9.54 4.128 12.048 ;
  LAYER M1 ;
        RECT 4.16 9.54 4.192 12.048 ;
  LAYER M1 ;
        RECT 4.224 9.54 4.256 12.048 ;
  LAYER M1 ;
        RECT 4.288 9.54 4.32 12.048 ;
  LAYER M1 ;
        RECT 4.352 9.54 4.384 12.048 ;
  LAYER M1 ;
        RECT 4.416 9.54 4.448 12.048 ;
  LAYER M1 ;
        RECT 4.48 9.54 4.512 12.048 ;
  LAYER M1 ;
        RECT 4.544 9.54 4.576 12.048 ;
  LAYER M1 ;
        RECT 4.608 9.54 4.64 12.048 ;
  LAYER M1 ;
        RECT 4.672 9.54 4.704 12.048 ;
  LAYER M1 ;
        RECT 4.736 9.54 4.768 12.048 ;
  LAYER M1 ;
        RECT 4.8 9.54 4.832 12.048 ;
  LAYER M1 ;
        RECT 4.864 9.54 4.896 12.048 ;
  LAYER M1 ;
        RECT 4.928 9.54 4.96 12.048 ;
  LAYER M1 ;
        RECT 4.992 9.54 5.024 12.048 ;
  LAYER M1 ;
        RECT 5.056 9.54 5.088 12.048 ;
  LAYER M1 ;
        RECT 5.12 9.54 5.152 12.048 ;
  LAYER M1 ;
        RECT 5.184 9.54 5.216 12.048 ;
  LAYER M1 ;
        RECT 5.248 9.54 5.28 12.048 ;
  LAYER M1 ;
        RECT 5.312 9.54 5.344 12.048 ;
  LAYER M1 ;
        RECT 5.376 9.54 5.408 12.048 ;
  LAYER M1 ;
        RECT 5.44 9.54 5.472 12.048 ;
  LAYER M1 ;
        RECT 5.504 9.54 5.536 12.048 ;
  LAYER M1 ;
        RECT 5.568 9.54 5.6 12.048 ;
  LAYER M2 ;
        RECT 3.244 9.624 5.716 9.656 ;
  LAYER M2 ;
        RECT 3.244 9.688 5.716 9.72 ;
  LAYER M2 ;
        RECT 3.244 9.752 5.716 9.784 ;
  LAYER M2 ;
        RECT 3.244 9.816 5.716 9.848 ;
  LAYER M2 ;
        RECT 3.244 9.88 5.716 9.912 ;
  LAYER M2 ;
        RECT 3.244 9.944 5.716 9.976 ;
  LAYER M2 ;
        RECT 3.244 10.008 5.716 10.04 ;
  LAYER M2 ;
        RECT 3.244 10.072 5.716 10.104 ;
  LAYER M2 ;
        RECT 3.244 10.136 5.716 10.168 ;
  LAYER M2 ;
        RECT 3.244 10.2 5.716 10.232 ;
  LAYER M2 ;
        RECT 3.244 10.264 5.716 10.296 ;
  LAYER M2 ;
        RECT 3.244 10.328 5.716 10.36 ;
  LAYER M2 ;
        RECT 3.244 10.392 5.716 10.424 ;
  LAYER M2 ;
        RECT 3.244 10.456 5.716 10.488 ;
  LAYER M2 ;
        RECT 3.244 10.52 5.716 10.552 ;
  LAYER M2 ;
        RECT 3.244 10.584 5.716 10.616 ;
  LAYER M2 ;
        RECT 3.244 10.648 5.716 10.68 ;
  LAYER M2 ;
        RECT 3.244 10.712 5.716 10.744 ;
  LAYER M2 ;
        RECT 3.244 10.776 5.716 10.808 ;
  LAYER M2 ;
        RECT 3.244 10.84 5.716 10.872 ;
  LAYER M2 ;
        RECT 3.244 10.904 5.716 10.936 ;
  LAYER M2 ;
        RECT 3.244 10.968 5.716 11 ;
  LAYER M2 ;
        RECT 3.244 11.032 5.716 11.064 ;
  LAYER M2 ;
        RECT 3.244 11.096 5.716 11.128 ;
  LAYER M2 ;
        RECT 3.244 11.16 5.716 11.192 ;
  LAYER M2 ;
        RECT 3.244 11.224 5.716 11.256 ;
  LAYER M2 ;
        RECT 3.244 11.288 5.716 11.32 ;
  LAYER M2 ;
        RECT 3.244 11.352 5.716 11.384 ;
  LAYER M2 ;
        RECT 3.244 11.416 5.716 11.448 ;
  LAYER M2 ;
        RECT 3.244 11.48 5.716 11.512 ;
  LAYER M2 ;
        RECT 3.244 11.544 5.716 11.576 ;
  LAYER M2 ;
        RECT 3.244 11.608 5.716 11.64 ;
  LAYER M2 ;
        RECT 3.244 11.672 5.716 11.704 ;
  LAYER M2 ;
        RECT 3.244 11.736 5.716 11.768 ;
  LAYER M2 ;
        RECT 3.244 11.8 5.716 11.832 ;
  LAYER M2 ;
        RECT 3.244 11.864 5.716 11.896 ;
  LAYER M3 ;
        RECT 3.264 9.54 3.296 12.048 ;
  LAYER M3 ;
        RECT 3.328 9.54 3.36 12.048 ;
  LAYER M3 ;
        RECT 3.392 9.54 3.424 12.048 ;
  LAYER M3 ;
        RECT 3.456 9.54 3.488 12.048 ;
  LAYER M3 ;
        RECT 3.52 9.54 3.552 12.048 ;
  LAYER M3 ;
        RECT 3.584 9.54 3.616 12.048 ;
  LAYER M3 ;
        RECT 3.648 9.54 3.68 12.048 ;
  LAYER M3 ;
        RECT 3.712 9.54 3.744 12.048 ;
  LAYER M3 ;
        RECT 3.776 9.54 3.808 12.048 ;
  LAYER M3 ;
        RECT 3.84 9.54 3.872 12.048 ;
  LAYER M3 ;
        RECT 3.904 9.54 3.936 12.048 ;
  LAYER M3 ;
        RECT 3.968 9.54 4 12.048 ;
  LAYER M3 ;
        RECT 4.032 9.54 4.064 12.048 ;
  LAYER M3 ;
        RECT 4.096 9.54 4.128 12.048 ;
  LAYER M3 ;
        RECT 4.16 9.54 4.192 12.048 ;
  LAYER M3 ;
        RECT 4.224 9.54 4.256 12.048 ;
  LAYER M3 ;
        RECT 4.288 9.54 4.32 12.048 ;
  LAYER M3 ;
        RECT 4.352 9.54 4.384 12.048 ;
  LAYER M3 ;
        RECT 4.416 9.54 4.448 12.048 ;
  LAYER M3 ;
        RECT 4.48 9.54 4.512 12.048 ;
  LAYER M3 ;
        RECT 4.544 9.54 4.576 12.048 ;
  LAYER M3 ;
        RECT 4.608 9.54 4.64 12.048 ;
  LAYER M3 ;
        RECT 4.672 9.54 4.704 12.048 ;
  LAYER M3 ;
        RECT 4.736 9.54 4.768 12.048 ;
  LAYER M3 ;
        RECT 4.8 9.54 4.832 12.048 ;
  LAYER M3 ;
        RECT 4.864 9.54 4.896 12.048 ;
  LAYER M3 ;
        RECT 4.928 9.54 4.96 12.048 ;
  LAYER M3 ;
        RECT 4.992 9.54 5.024 12.048 ;
  LAYER M3 ;
        RECT 5.056 9.54 5.088 12.048 ;
  LAYER M3 ;
        RECT 5.12 9.54 5.152 12.048 ;
  LAYER M3 ;
        RECT 5.184 9.54 5.216 12.048 ;
  LAYER M3 ;
        RECT 5.248 9.54 5.28 12.048 ;
  LAYER M3 ;
        RECT 5.312 9.54 5.344 12.048 ;
  LAYER M3 ;
        RECT 5.376 9.54 5.408 12.048 ;
  LAYER M3 ;
        RECT 5.44 9.54 5.472 12.048 ;
  LAYER M3 ;
        RECT 5.504 9.54 5.536 12.048 ;
  LAYER M3 ;
        RECT 5.568 9.54 5.6 12.048 ;
  LAYER M3 ;
        RECT 5.664 9.54 5.696 12.048 ;
  LAYER M1 ;
        RECT 3.279 9.576 3.281 12.012 ;
  LAYER M1 ;
        RECT 3.359 9.576 3.361 12.012 ;
  LAYER M1 ;
        RECT 3.439 9.576 3.441 12.012 ;
  LAYER M1 ;
        RECT 3.519 9.576 3.521 12.012 ;
  LAYER M1 ;
        RECT 3.599 9.576 3.601 12.012 ;
  LAYER M1 ;
        RECT 3.679 9.576 3.681 12.012 ;
  LAYER M1 ;
        RECT 3.759 9.576 3.761 12.012 ;
  LAYER M1 ;
        RECT 3.839 9.576 3.841 12.012 ;
  LAYER M1 ;
        RECT 3.919 9.576 3.921 12.012 ;
  LAYER M1 ;
        RECT 3.999 9.576 4.001 12.012 ;
  LAYER M1 ;
        RECT 4.079 9.576 4.081 12.012 ;
  LAYER M1 ;
        RECT 4.159 9.576 4.161 12.012 ;
  LAYER M1 ;
        RECT 4.239 9.576 4.241 12.012 ;
  LAYER M1 ;
        RECT 4.319 9.576 4.321 12.012 ;
  LAYER M1 ;
        RECT 4.399 9.576 4.401 12.012 ;
  LAYER M1 ;
        RECT 4.479 9.576 4.481 12.012 ;
  LAYER M1 ;
        RECT 4.559 9.576 4.561 12.012 ;
  LAYER M1 ;
        RECT 4.639 9.576 4.641 12.012 ;
  LAYER M1 ;
        RECT 4.719 9.576 4.721 12.012 ;
  LAYER M1 ;
        RECT 4.799 9.576 4.801 12.012 ;
  LAYER M1 ;
        RECT 4.879 9.576 4.881 12.012 ;
  LAYER M1 ;
        RECT 4.959 9.576 4.961 12.012 ;
  LAYER M1 ;
        RECT 5.039 9.576 5.041 12.012 ;
  LAYER M1 ;
        RECT 5.119 9.576 5.121 12.012 ;
  LAYER M1 ;
        RECT 5.199 9.576 5.201 12.012 ;
  LAYER M1 ;
        RECT 5.279 9.576 5.281 12.012 ;
  LAYER M1 ;
        RECT 5.359 9.576 5.361 12.012 ;
  LAYER M1 ;
        RECT 5.439 9.576 5.441 12.012 ;
  LAYER M1 ;
        RECT 5.519 9.576 5.521 12.012 ;
  LAYER M1 ;
        RECT 5.599 9.576 5.601 12.012 ;
  LAYER M2 ;
        RECT 3.28 9.575 5.68 9.577 ;
  LAYER M2 ;
        RECT 3.28 9.659 5.68 9.661 ;
  LAYER M2 ;
        RECT 3.28 9.743 5.68 9.745 ;
  LAYER M2 ;
        RECT 3.28 9.827 5.68 9.829 ;
  LAYER M2 ;
        RECT 3.28 9.911 5.68 9.913 ;
  LAYER M2 ;
        RECT 3.28 9.995 5.68 9.997 ;
  LAYER M2 ;
        RECT 3.28 10.079 5.68 10.081 ;
  LAYER M2 ;
        RECT 3.28 10.163 5.68 10.165 ;
  LAYER M2 ;
        RECT 3.28 10.247 5.68 10.249 ;
  LAYER M2 ;
        RECT 3.28 10.331 5.68 10.333 ;
  LAYER M2 ;
        RECT 3.28 10.415 5.68 10.417 ;
  LAYER M2 ;
        RECT 3.28 10.499 5.68 10.501 ;
  LAYER M2 ;
        RECT 3.28 10.5825 5.68 10.5845 ;
  LAYER M2 ;
        RECT 3.28 10.667 5.68 10.669 ;
  LAYER M2 ;
        RECT 3.28 10.751 5.68 10.753 ;
  LAYER M2 ;
        RECT 3.28 10.835 5.68 10.837 ;
  LAYER M2 ;
        RECT 3.28 10.919 5.68 10.921 ;
  LAYER M2 ;
        RECT 3.28 11.003 5.68 11.005 ;
  LAYER M2 ;
        RECT 3.28 11.087 5.68 11.089 ;
  LAYER M2 ;
        RECT 3.28 11.171 5.68 11.173 ;
  LAYER M2 ;
        RECT 3.28 11.255 5.68 11.257 ;
  LAYER M2 ;
        RECT 3.28 11.339 5.68 11.341 ;
  LAYER M2 ;
        RECT 3.28 11.423 5.68 11.425 ;
  LAYER M2 ;
        RECT 3.28 11.507 5.68 11.509 ;
  LAYER M2 ;
        RECT 3.28 11.591 5.68 11.593 ;
  LAYER M2 ;
        RECT 3.28 11.675 5.68 11.677 ;
  LAYER M2 ;
        RECT 3.28 11.759 5.68 11.761 ;
  LAYER M2 ;
        RECT 3.28 11.843 5.68 11.845 ;
  LAYER M2 ;
        RECT 3.28 11.927 5.68 11.929 ;
  LAYER M1 ;
        RECT 3.264 12.48 3.296 14.988 ;
  LAYER M1 ;
        RECT 3.328 12.48 3.36 14.988 ;
  LAYER M1 ;
        RECT 3.392 12.48 3.424 14.988 ;
  LAYER M1 ;
        RECT 3.456 12.48 3.488 14.988 ;
  LAYER M1 ;
        RECT 3.52 12.48 3.552 14.988 ;
  LAYER M1 ;
        RECT 3.584 12.48 3.616 14.988 ;
  LAYER M1 ;
        RECT 3.648 12.48 3.68 14.988 ;
  LAYER M1 ;
        RECT 3.712 12.48 3.744 14.988 ;
  LAYER M1 ;
        RECT 3.776 12.48 3.808 14.988 ;
  LAYER M1 ;
        RECT 3.84 12.48 3.872 14.988 ;
  LAYER M1 ;
        RECT 3.904 12.48 3.936 14.988 ;
  LAYER M1 ;
        RECT 3.968 12.48 4 14.988 ;
  LAYER M1 ;
        RECT 4.032 12.48 4.064 14.988 ;
  LAYER M1 ;
        RECT 4.096 12.48 4.128 14.988 ;
  LAYER M1 ;
        RECT 4.16 12.48 4.192 14.988 ;
  LAYER M1 ;
        RECT 4.224 12.48 4.256 14.988 ;
  LAYER M1 ;
        RECT 4.288 12.48 4.32 14.988 ;
  LAYER M1 ;
        RECT 4.352 12.48 4.384 14.988 ;
  LAYER M1 ;
        RECT 4.416 12.48 4.448 14.988 ;
  LAYER M1 ;
        RECT 4.48 12.48 4.512 14.988 ;
  LAYER M1 ;
        RECT 4.544 12.48 4.576 14.988 ;
  LAYER M1 ;
        RECT 4.608 12.48 4.64 14.988 ;
  LAYER M1 ;
        RECT 4.672 12.48 4.704 14.988 ;
  LAYER M1 ;
        RECT 4.736 12.48 4.768 14.988 ;
  LAYER M1 ;
        RECT 4.8 12.48 4.832 14.988 ;
  LAYER M1 ;
        RECT 4.864 12.48 4.896 14.988 ;
  LAYER M1 ;
        RECT 4.928 12.48 4.96 14.988 ;
  LAYER M1 ;
        RECT 4.992 12.48 5.024 14.988 ;
  LAYER M1 ;
        RECT 5.056 12.48 5.088 14.988 ;
  LAYER M1 ;
        RECT 5.12 12.48 5.152 14.988 ;
  LAYER M1 ;
        RECT 5.184 12.48 5.216 14.988 ;
  LAYER M1 ;
        RECT 5.248 12.48 5.28 14.988 ;
  LAYER M1 ;
        RECT 5.312 12.48 5.344 14.988 ;
  LAYER M1 ;
        RECT 5.376 12.48 5.408 14.988 ;
  LAYER M1 ;
        RECT 5.44 12.48 5.472 14.988 ;
  LAYER M1 ;
        RECT 5.504 12.48 5.536 14.988 ;
  LAYER M1 ;
        RECT 5.568 12.48 5.6 14.988 ;
  LAYER M2 ;
        RECT 3.244 12.564 5.716 12.596 ;
  LAYER M2 ;
        RECT 3.244 12.628 5.716 12.66 ;
  LAYER M2 ;
        RECT 3.244 12.692 5.716 12.724 ;
  LAYER M2 ;
        RECT 3.244 12.756 5.716 12.788 ;
  LAYER M2 ;
        RECT 3.244 12.82 5.716 12.852 ;
  LAYER M2 ;
        RECT 3.244 12.884 5.716 12.916 ;
  LAYER M2 ;
        RECT 3.244 12.948 5.716 12.98 ;
  LAYER M2 ;
        RECT 3.244 13.012 5.716 13.044 ;
  LAYER M2 ;
        RECT 3.244 13.076 5.716 13.108 ;
  LAYER M2 ;
        RECT 3.244 13.14 5.716 13.172 ;
  LAYER M2 ;
        RECT 3.244 13.204 5.716 13.236 ;
  LAYER M2 ;
        RECT 3.244 13.268 5.716 13.3 ;
  LAYER M2 ;
        RECT 3.244 13.332 5.716 13.364 ;
  LAYER M2 ;
        RECT 3.244 13.396 5.716 13.428 ;
  LAYER M2 ;
        RECT 3.244 13.46 5.716 13.492 ;
  LAYER M2 ;
        RECT 3.244 13.524 5.716 13.556 ;
  LAYER M2 ;
        RECT 3.244 13.588 5.716 13.62 ;
  LAYER M2 ;
        RECT 3.244 13.652 5.716 13.684 ;
  LAYER M2 ;
        RECT 3.244 13.716 5.716 13.748 ;
  LAYER M2 ;
        RECT 3.244 13.78 5.716 13.812 ;
  LAYER M2 ;
        RECT 3.244 13.844 5.716 13.876 ;
  LAYER M2 ;
        RECT 3.244 13.908 5.716 13.94 ;
  LAYER M2 ;
        RECT 3.244 13.972 5.716 14.004 ;
  LAYER M2 ;
        RECT 3.244 14.036 5.716 14.068 ;
  LAYER M2 ;
        RECT 3.244 14.1 5.716 14.132 ;
  LAYER M2 ;
        RECT 3.244 14.164 5.716 14.196 ;
  LAYER M2 ;
        RECT 3.244 14.228 5.716 14.26 ;
  LAYER M2 ;
        RECT 3.244 14.292 5.716 14.324 ;
  LAYER M2 ;
        RECT 3.244 14.356 5.716 14.388 ;
  LAYER M2 ;
        RECT 3.244 14.42 5.716 14.452 ;
  LAYER M2 ;
        RECT 3.244 14.484 5.716 14.516 ;
  LAYER M2 ;
        RECT 3.244 14.548 5.716 14.58 ;
  LAYER M2 ;
        RECT 3.244 14.612 5.716 14.644 ;
  LAYER M2 ;
        RECT 3.244 14.676 5.716 14.708 ;
  LAYER M2 ;
        RECT 3.244 14.74 5.716 14.772 ;
  LAYER M2 ;
        RECT 3.244 14.804 5.716 14.836 ;
  LAYER M3 ;
        RECT 3.264 12.48 3.296 14.988 ;
  LAYER M3 ;
        RECT 3.328 12.48 3.36 14.988 ;
  LAYER M3 ;
        RECT 3.392 12.48 3.424 14.988 ;
  LAYER M3 ;
        RECT 3.456 12.48 3.488 14.988 ;
  LAYER M3 ;
        RECT 3.52 12.48 3.552 14.988 ;
  LAYER M3 ;
        RECT 3.584 12.48 3.616 14.988 ;
  LAYER M3 ;
        RECT 3.648 12.48 3.68 14.988 ;
  LAYER M3 ;
        RECT 3.712 12.48 3.744 14.988 ;
  LAYER M3 ;
        RECT 3.776 12.48 3.808 14.988 ;
  LAYER M3 ;
        RECT 3.84 12.48 3.872 14.988 ;
  LAYER M3 ;
        RECT 3.904 12.48 3.936 14.988 ;
  LAYER M3 ;
        RECT 3.968 12.48 4 14.988 ;
  LAYER M3 ;
        RECT 4.032 12.48 4.064 14.988 ;
  LAYER M3 ;
        RECT 4.096 12.48 4.128 14.988 ;
  LAYER M3 ;
        RECT 4.16 12.48 4.192 14.988 ;
  LAYER M3 ;
        RECT 4.224 12.48 4.256 14.988 ;
  LAYER M3 ;
        RECT 4.288 12.48 4.32 14.988 ;
  LAYER M3 ;
        RECT 4.352 12.48 4.384 14.988 ;
  LAYER M3 ;
        RECT 4.416 12.48 4.448 14.988 ;
  LAYER M3 ;
        RECT 4.48 12.48 4.512 14.988 ;
  LAYER M3 ;
        RECT 4.544 12.48 4.576 14.988 ;
  LAYER M3 ;
        RECT 4.608 12.48 4.64 14.988 ;
  LAYER M3 ;
        RECT 4.672 12.48 4.704 14.988 ;
  LAYER M3 ;
        RECT 4.736 12.48 4.768 14.988 ;
  LAYER M3 ;
        RECT 4.8 12.48 4.832 14.988 ;
  LAYER M3 ;
        RECT 4.864 12.48 4.896 14.988 ;
  LAYER M3 ;
        RECT 4.928 12.48 4.96 14.988 ;
  LAYER M3 ;
        RECT 4.992 12.48 5.024 14.988 ;
  LAYER M3 ;
        RECT 5.056 12.48 5.088 14.988 ;
  LAYER M3 ;
        RECT 5.12 12.48 5.152 14.988 ;
  LAYER M3 ;
        RECT 5.184 12.48 5.216 14.988 ;
  LAYER M3 ;
        RECT 5.248 12.48 5.28 14.988 ;
  LAYER M3 ;
        RECT 5.312 12.48 5.344 14.988 ;
  LAYER M3 ;
        RECT 5.376 12.48 5.408 14.988 ;
  LAYER M3 ;
        RECT 5.44 12.48 5.472 14.988 ;
  LAYER M3 ;
        RECT 5.504 12.48 5.536 14.988 ;
  LAYER M3 ;
        RECT 5.568 12.48 5.6 14.988 ;
  LAYER M3 ;
        RECT 5.664 12.48 5.696 14.988 ;
  LAYER M1 ;
        RECT 3.279 12.516 3.281 14.952 ;
  LAYER M1 ;
        RECT 3.359 12.516 3.361 14.952 ;
  LAYER M1 ;
        RECT 3.439 12.516 3.441 14.952 ;
  LAYER M1 ;
        RECT 3.519 12.516 3.521 14.952 ;
  LAYER M1 ;
        RECT 3.599 12.516 3.601 14.952 ;
  LAYER M1 ;
        RECT 3.679 12.516 3.681 14.952 ;
  LAYER M1 ;
        RECT 3.759 12.516 3.761 14.952 ;
  LAYER M1 ;
        RECT 3.839 12.516 3.841 14.952 ;
  LAYER M1 ;
        RECT 3.919 12.516 3.921 14.952 ;
  LAYER M1 ;
        RECT 3.999 12.516 4.001 14.952 ;
  LAYER M1 ;
        RECT 4.079 12.516 4.081 14.952 ;
  LAYER M1 ;
        RECT 4.159 12.516 4.161 14.952 ;
  LAYER M1 ;
        RECT 4.239 12.516 4.241 14.952 ;
  LAYER M1 ;
        RECT 4.319 12.516 4.321 14.952 ;
  LAYER M1 ;
        RECT 4.399 12.516 4.401 14.952 ;
  LAYER M1 ;
        RECT 4.479 12.516 4.481 14.952 ;
  LAYER M1 ;
        RECT 4.559 12.516 4.561 14.952 ;
  LAYER M1 ;
        RECT 4.639 12.516 4.641 14.952 ;
  LAYER M1 ;
        RECT 4.719 12.516 4.721 14.952 ;
  LAYER M1 ;
        RECT 4.799 12.516 4.801 14.952 ;
  LAYER M1 ;
        RECT 4.879 12.516 4.881 14.952 ;
  LAYER M1 ;
        RECT 4.959 12.516 4.961 14.952 ;
  LAYER M1 ;
        RECT 5.039 12.516 5.041 14.952 ;
  LAYER M1 ;
        RECT 5.119 12.516 5.121 14.952 ;
  LAYER M1 ;
        RECT 5.199 12.516 5.201 14.952 ;
  LAYER M1 ;
        RECT 5.279 12.516 5.281 14.952 ;
  LAYER M1 ;
        RECT 5.359 12.516 5.361 14.952 ;
  LAYER M1 ;
        RECT 5.439 12.516 5.441 14.952 ;
  LAYER M1 ;
        RECT 5.519 12.516 5.521 14.952 ;
  LAYER M1 ;
        RECT 5.599 12.516 5.601 14.952 ;
  LAYER M2 ;
        RECT 3.28 12.515 5.68 12.517 ;
  LAYER M2 ;
        RECT 3.28 12.599 5.68 12.601 ;
  LAYER M2 ;
        RECT 3.28 12.683 5.68 12.685 ;
  LAYER M2 ;
        RECT 3.28 12.767 5.68 12.769 ;
  LAYER M2 ;
        RECT 3.28 12.851 5.68 12.853 ;
  LAYER M2 ;
        RECT 3.28 12.935 5.68 12.937 ;
  LAYER M2 ;
        RECT 3.28 13.019 5.68 13.021 ;
  LAYER M2 ;
        RECT 3.28 13.103 5.68 13.105 ;
  LAYER M2 ;
        RECT 3.28 13.187 5.68 13.189 ;
  LAYER M2 ;
        RECT 3.28 13.271 5.68 13.273 ;
  LAYER M2 ;
        RECT 3.28 13.355 5.68 13.357 ;
  LAYER M2 ;
        RECT 3.28 13.439 5.68 13.441 ;
  LAYER M2 ;
        RECT 3.28 13.5225 5.68 13.5245 ;
  LAYER M2 ;
        RECT 3.28 13.607 5.68 13.609 ;
  LAYER M2 ;
        RECT 3.28 13.691 5.68 13.693 ;
  LAYER M2 ;
        RECT 3.28 13.775 5.68 13.777 ;
  LAYER M2 ;
        RECT 3.28 13.859 5.68 13.861 ;
  LAYER M2 ;
        RECT 3.28 13.943 5.68 13.945 ;
  LAYER M2 ;
        RECT 3.28 14.027 5.68 14.029 ;
  LAYER M2 ;
        RECT 3.28 14.111 5.68 14.113 ;
  LAYER M2 ;
        RECT 3.28 14.195 5.68 14.197 ;
  LAYER M2 ;
        RECT 3.28 14.279 5.68 14.281 ;
  LAYER M2 ;
        RECT 3.28 14.363 5.68 14.365 ;
  LAYER M2 ;
        RECT 3.28 14.447 5.68 14.449 ;
  LAYER M2 ;
        RECT 3.28 14.531 5.68 14.533 ;
  LAYER M2 ;
        RECT 3.28 14.615 5.68 14.617 ;
  LAYER M2 ;
        RECT 3.28 14.699 5.68 14.701 ;
  LAYER M2 ;
        RECT 3.28 14.783 5.68 14.785 ;
  LAYER M2 ;
        RECT 3.28 14.867 5.68 14.869 ;
  LAYER M1 ;
        RECT 3.264 15.42 3.296 17.928 ;
  LAYER M1 ;
        RECT 3.328 15.42 3.36 17.928 ;
  LAYER M1 ;
        RECT 3.392 15.42 3.424 17.928 ;
  LAYER M1 ;
        RECT 3.456 15.42 3.488 17.928 ;
  LAYER M1 ;
        RECT 3.52 15.42 3.552 17.928 ;
  LAYER M1 ;
        RECT 3.584 15.42 3.616 17.928 ;
  LAYER M1 ;
        RECT 3.648 15.42 3.68 17.928 ;
  LAYER M1 ;
        RECT 3.712 15.42 3.744 17.928 ;
  LAYER M1 ;
        RECT 3.776 15.42 3.808 17.928 ;
  LAYER M1 ;
        RECT 3.84 15.42 3.872 17.928 ;
  LAYER M1 ;
        RECT 3.904 15.42 3.936 17.928 ;
  LAYER M1 ;
        RECT 3.968 15.42 4 17.928 ;
  LAYER M1 ;
        RECT 4.032 15.42 4.064 17.928 ;
  LAYER M1 ;
        RECT 4.096 15.42 4.128 17.928 ;
  LAYER M1 ;
        RECT 4.16 15.42 4.192 17.928 ;
  LAYER M1 ;
        RECT 4.224 15.42 4.256 17.928 ;
  LAYER M1 ;
        RECT 4.288 15.42 4.32 17.928 ;
  LAYER M1 ;
        RECT 4.352 15.42 4.384 17.928 ;
  LAYER M1 ;
        RECT 4.416 15.42 4.448 17.928 ;
  LAYER M1 ;
        RECT 4.48 15.42 4.512 17.928 ;
  LAYER M1 ;
        RECT 4.544 15.42 4.576 17.928 ;
  LAYER M1 ;
        RECT 4.608 15.42 4.64 17.928 ;
  LAYER M1 ;
        RECT 4.672 15.42 4.704 17.928 ;
  LAYER M1 ;
        RECT 4.736 15.42 4.768 17.928 ;
  LAYER M1 ;
        RECT 4.8 15.42 4.832 17.928 ;
  LAYER M1 ;
        RECT 4.864 15.42 4.896 17.928 ;
  LAYER M1 ;
        RECT 4.928 15.42 4.96 17.928 ;
  LAYER M1 ;
        RECT 4.992 15.42 5.024 17.928 ;
  LAYER M1 ;
        RECT 5.056 15.42 5.088 17.928 ;
  LAYER M1 ;
        RECT 5.12 15.42 5.152 17.928 ;
  LAYER M1 ;
        RECT 5.184 15.42 5.216 17.928 ;
  LAYER M1 ;
        RECT 5.248 15.42 5.28 17.928 ;
  LAYER M1 ;
        RECT 5.312 15.42 5.344 17.928 ;
  LAYER M1 ;
        RECT 5.376 15.42 5.408 17.928 ;
  LAYER M1 ;
        RECT 5.44 15.42 5.472 17.928 ;
  LAYER M1 ;
        RECT 5.504 15.42 5.536 17.928 ;
  LAYER M1 ;
        RECT 5.568 15.42 5.6 17.928 ;
  LAYER M2 ;
        RECT 3.244 15.504 5.716 15.536 ;
  LAYER M2 ;
        RECT 3.244 15.568 5.716 15.6 ;
  LAYER M2 ;
        RECT 3.244 15.632 5.716 15.664 ;
  LAYER M2 ;
        RECT 3.244 15.696 5.716 15.728 ;
  LAYER M2 ;
        RECT 3.244 15.76 5.716 15.792 ;
  LAYER M2 ;
        RECT 3.244 15.824 5.716 15.856 ;
  LAYER M2 ;
        RECT 3.244 15.888 5.716 15.92 ;
  LAYER M2 ;
        RECT 3.244 15.952 5.716 15.984 ;
  LAYER M2 ;
        RECT 3.244 16.016 5.716 16.048 ;
  LAYER M2 ;
        RECT 3.244 16.08 5.716 16.112 ;
  LAYER M2 ;
        RECT 3.244 16.144 5.716 16.176 ;
  LAYER M2 ;
        RECT 3.244 16.208 5.716 16.24 ;
  LAYER M2 ;
        RECT 3.244 16.272 5.716 16.304 ;
  LAYER M2 ;
        RECT 3.244 16.336 5.716 16.368 ;
  LAYER M2 ;
        RECT 3.244 16.4 5.716 16.432 ;
  LAYER M2 ;
        RECT 3.244 16.464 5.716 16.496 ;
  LAYER M2 ;
        RECT 3.244 16.528 5.716 16.56 ;
  LAYER M2 ;
        RECT 3.244 16.592 5.716 16.624 ;
  LAYER M2 ;
        RECT 3.244 16.656 5.716 16.688 ;
  LAYER M2 ;
        RECT 3.244 16.72 5.716 16.752 ;
  LAYER M2 ;
        RECT 3.244 16.784 5.716 16.816 ;
  LAYER M2 ;
        RECT 3.244 16.848 5.716 16.88 ;
  LAYER M2 ;
        RECT 3.244 16.912 5.716 16.944 ;
  LAYER M2 ;
        RECT 3.244 16.976 5.716 17.008 ;
  LAYER M2 ;
        RECT 3.244 17.04 5.716 17.072 ;
  LAYER M2 ;
        RECT 3.244 17.104 5.716 17.136 ;
  LAYER M2 ;
        RECT 3.244 17.168 5.716 17.2 ;
  LAYER M2 ;
        RECT 3.244 17.232 5.716 17.264 ;
  LAYER M2 ;
        RECT 3.244 17.296 5.716 17.328 ;
  LAYER M2 ;
        RECT 3.244 17.36 5.716 17.392 ;
  LAYER M2 ;
        RECT 3.244 17.424 5.716 17.456 ;
  LAYER M2 ;
        RECT 3.244 17.488 5.716 17.52 ;
  LAYER M2 ;
        RECT 3.244 17.552 5.716 17.584 ;
  LAYER M2 ;
        RECT 3.244 17.616 5.716 17.648 ;
  LAYER M2 ;
        RECT 3.244 17.68 5.716 17.712 ;
  LAYER M2 ;
        RECT 3.244 17.744 5.716 17.776 ;
  LAYER M3 ;
        RECT 3.264 15.42 3.296 17.928 ;
  LAYER M3 ;
        RECT 3.328 15.42 3.36 17.928 ;
  LAYER M3 ;
        RECT 3.392 15.42 3.424 17.928 ;
  LAYER M3 ;
        RECT 3.456 15.42 3.488 17.928 ;
  LAYER M3 ;
        RECT 3.52 15.42 3.552 17.928 ;
  LAYER M3 ;
        RECT 3.584 15.42 3.616 17.928 ;
  LAYER M3 ;
        RECT 3.648 15.42 3.68 17.928 ;
  LAYER M3 ;
        RECT 3.712 15.42 3.744 17.928 ;
  LAYER M3 ;
        RECT 3.776 15.42 3.808 17.928 ;
  LAYER M3 ;
        RECT 3.84 15.42 3.872 17.928 ;
  LAYER M3 ;
        RECT 3.904 15.42 3.936 17.928 ;
  LAYER M3 ;
        RECT 3.968 15.42 4 17.928 ;
  LAYER M3 ;
        RECT 4.032 15.42 4.064 17.928 ;
  LAYER M3 ;
        RECT 4.096 15.42 4.128 17.928 ;
  LAYER M3 ;
        RECT 4.16 15.42 4.192 17.928 ;
  LAYER M3 ;
        RECT 4.224 15.42 4.256 17.928 ;
  LAYER M3 ;
        RECT 4.288 15.42 4.32 17.928 ;
  LAYER M3 ;
        RECT 4.352 15.42 4.384 17.928 ;
  LAYER M3 ;
        RECT 4.416 15.42 4.448 17.928 ;
  LAYER M3 ;
        RECT 4.48 15.42 4.512 17.928 ;
  LAYER M3 ;
        RECT 4.544 15.42 4.576 17.928 ;
  LAYER M3 ;
        RECT 4.608 15.42 4.64 17.928 ;
  LAYER M3 ;
        RECT 4.672 15.42 4.704 17.928 ;
  LAYER M3 ;
        RECT 4.736 15.42 4.768 17.928 ;
  LAYER M3 ;
        RECT 4.8 15.42 4.832 17.928 ;
  LAYER M3 ;
        RECT 4.864 15.42 4.896 17.928 ;
  LAYER M3 ;
        RECT 4.928 15.42 4.96 17.928 ;
  LAYER M3 ;
        RECT 4.992 15.42 5.024 17.928 ;
  LAYER M3 ;
        RECT 5.056 15.42 5.088 17.928 ;
  LAYER M3 ;
        RECT 5.12 15.42 5.152 17.928 ;
  LAYER M3 ;
        RECT 5.184 15.42 5.216 17.928 ;
  LAYER M3 ;
        RECT 5.248 15.42 5.28 17.928 ;
  LAYER M3 ;
        RECT 5.312 15.42 5.344 17.928 ;
  LAYER M3 ;
        RECT 5.376 15.42 5.408 17.928 ;
  LAYER M3 ;
        RECT 5.44 15.42 5.472 17.928 ;
  LAYER M3 ;
        RECT 5.504 15.42 5.536 17.928 ;
  LAYER M3 ;
        RECT 5.568 15.42 5.6 17.928 ;
  LAYER M3 ;
        RECT 5.664 15.42 5.696 17.928 ;
  LAYER M1 ;
        RECT 3.279 15.456 3.281 17.892 ;
  LAYER M1 ;
        RECT 3.359 15.456 3.361 17.892 ;
  LAYER M1 ;
        RECT 3.439 15.456 3.441 17.892 ;
  LAYER M1 ;
        RECT 3.519 15.456 3.521 17.892 ;
  LAYER M1 ;
        RECT 3.599 15.456 3.601 17.892 ;
  LAYER M1 ;
        RECT 3.679 15.456 3.681 17.892 ;
  LAYER M1 ;
        RECT 3.759 15.456 3.761 17.892 ;
  LAYER M1 ;
        RECT 3.839 15.456 3.841 17.892 ;
  LAYER M1 ;
        RECT 3.919 15.456 3.921 17.892 ;
  LAYER M1 ;
        RECT 3.999 15.456 4.001 17.892 ;
  LAYER M1 ;
        RECT 4.079 15.456 4.081 17.892 ;
  LAYER M1 ;
        RECT 4.159 15.456 4.161 17.892 ;
  LAYER M1 ;
        RECT 4.239 15.456 4.241 17.892 ;
  LAYER M1 ;
        RECT 4.319 15.456 4.321 17.892 ;
  LAYER M1 ;
        RECT 4.399 15.456 4.401 17.892 ;
  LAYER M1 ;
        RECT 4.479 15.456 4.481 17.892 ;
  LAYER M1 ;
        RECT 4.559 15.456 4.561 17.892 ;
  LAYER M1 ;
        RECT 4.639 15.456 4.641 17.892 ;
  LAYER M1 ;
        RECT 4.719 15.456 4.721 17.892 ;
  LAYER M1 ;
        RECT 4.799 15.456 4.801 17.892 ;
  LAYER M1 ;
        RECT 4.879 15.456 4.881 17.892 ;
  LAYER M1 ;
        RECT 4.959 15.456 4.961 17.892 ;
  LAYER M1 ;
        RECT 5.039 15.456 5.041 17.892 ;
  LAYER M1 ;
        RECT 5.119 15.456 5.121 17.892 ;
  LAYER M1 ;
        RECT 5.199 15.456 5.201 17.892 ;
  LAYER M1 ;
        RECT 5.279 15.456 5.281 17.892 ;
  LAYER M1 ;
        RECT 5.359 15.456 5.361 17.892 ;
  LAYER M1 ;
        RECT 5.439 15.456 5.441 17.892 ;
  LAYER M1 ;
        RECT 5.519 15.456 5.521 17.892 ;
  LAYER M1 ;
        RECT 5.599 15.456 5.601 17.892 ;
  LAYER M2 ;
        RECT 3.28 15.455 5.68 15.457 ;
  LAYER M2 ;
        RECT 3.28 15.539 5.68 15.541 ;
  LAYER M2 ;
        RECT 3.28 15.623 5.68 15.625 ;
  LAYER M2 ;
        RECT 3.28 15.707 5.68 15.709 ;
  LAYER M2 ;
        RECT 3.28 15.791 5.68 15.793 ;
  LAYER M2 ;
        RECT 3.28 15.875 5.68 15.877 ;
  LAYER M2 ;
        RECT 3.28 15.959 5.68 15.961 ;
  LAYER M2 ;
        RECT 3.28 16.043 5.68 16.045 ;
  LAYER M2 ;
        RECT 3.28 16.127 5.68 16.129 ;
  LAYER M2 ;
        RECT 3.28 16.211 5.68 16.213 ;
  LAYER M2 ;
        RECT 3.28 16.295 5.68 16.297 ;
  LAYER M2 ;
        RECT 3.28 16.379 5.68 16.381 ;
  LAYER M2 ;
        RECT 3.28 16.4625 5.68 16.4645 ;
  LAYER M2 ;
        RECT 3.28 16.547 5.68 16.549 ;
  LAYER M2 ;
        RECT 3.28 16.631 5.68 16.633 ;
  LAYER M2 ;
        RECT 3.28 16.715 5.68 16.717 ;
  LAYER M2 ;
        RECT 3.28 16.799 5.68 16.801 ;
  LAYER M2 ;
        RECT 3.28 16.883 5.68 16.885 ;
  LAYER M2 ;
        RECT 3.28 16.967 5.68 16.969 ;
  LAYER M2 ;
        RECT 3.28 17.051 5.68 17.053 ;
  LAYER M2 ;
        RECT 3.28 17.135 5.68 17.137 ;
  LAYER M2 ;
        RECT 3.28 17.219 5.68 17.221 ;
  LAYER M2 ;
        RECT 3.28 17.303 5.68 17.305 ;
  LAYER M2 ;
        RECT 3.28 17.387 5.68 17.389 ;
  LAYER M2 ;
        RECT 3.28 17.471 5.68 17.473 ;
  LAYER M2 ;
        RECT 3.28 17.555 5.68 17.557 ;
  LAYER M2 ;
        RECT 3.28 17.639 5.68 17.641 ;
  LAYER M2 ;
        RECT 3.28 17.723 5.68 17.725 ;
  LAYER M2 ;
        RECT 3.28 17.807 5.68 17.809 ;
  LAYER M1 ;
        RECT 6.144 0.72 6.176 3.228 ;
  LAYER M1 ;
        RECT 6.208 0.72 6.24 3.228 ;
  LAYER M1 ;
        RECT 6.272 0.72 6.304 3.228 ;
  LAYER M1 ;
        RECT 6.336 0.72 6.368 3.228 ;
  LAYER M1 ;
        RECT 6.4 0.72 6.432 3.228 ;
  LAYER M1 ;
        RECT 6.464 0.72 6.496 3.228 ;
  LAYER M1 ;
        RECT 6.528 0.72 6.56 3.228 ;
  LAYER M1 ;
        RECT 6.592 0.72 6.624 3.228 ;
  LAYER M1 ;
        RECT 6.656 0.72 6.688 3.228 ;
  LAYER M1 ;
        RECT 6.72 0.72 6.752 3.228 ;
  LAYER M1 ;
        RECT 6.784 0.72 6.816 3.228 ;
  LAYER M1 ;
        RECT 6.848 0.72 6.88 3.228 ;
  LAYER M1 ;
        RECT 6.912 0.72 6.944 3.228 ;
  LAYER M1 ;
        RECT 6.976 0.72 7.008 3.228 ;
  LAYER M1 ;
        RECT 7.04 0.72 7.072 3.228 ;
  LAYER M1 ;
        RECT 7.104 0.72 7.136 3.228 ;
  LAYER M1 ;
        RECT 7.168 0.72 7.2 3.228 ;
  LAYER M1 ;
        RECT 7.232 0.72 7.264 3.228 ;
  LAYER M1 ;
        RECT 7.296 0.72 7.328 3.228 ;
  LAYER M1 ;
        RECT 7.36 0.72 7.392 3.228 ;
  LAYER M1 ;
        RECT 7.424 0.72 7.456 3.228 ;
  LAYER M1 ;
        RECT 7.488 0.72 7.52 3.228 ;
  LAYER M1 ;
        RECT 7.552 0.72 7.584 3.228 ;
  LAYER M1 ;
        RECT 7.616 0.72 7.648 3.228 ;
  LAYER M1 ;
        RECT 7.68 0.72 7.712 3.228 ;
  LAYER M1 ;
        RECT 7.744 0.72 7.776 3.228 ;
  LAYER M1 ;
        RECT 7.808 0.72 7.84 3.228 ;
  LAYER M1 ;
        RECT 7.872 0.72 7.904 3.228 ;
  LAYER M1 ;
        RECT 7.936 0.72 7.968 3.228 ;
  LAYER M1 ;
        RECT 8 0.72 8.032 3.228 ;
  LAYER M1 ;
        RECT 8.064 0.72 8.096 3.228 ;
  LAYER M1 ;
        RECT 8.128 0.72 8.16 3.228 ;
  LAYER M1 ;
        RECT 8.192 0.72 8.224 3.228 ;
  LAYER M1 ;
        RECT 8.256 0.72 8.288 3.228 ;
  LAYER M1 ;
        RECT 8.32 0.72 8.352 3.228 ;
  LAYER M1 ;
        RECT 8.384 0.72 8.416 3.228 ;
  LAYER M1 ;
        RECT 8.448 0.72 8.48 3.228 ;
  LAYER M2 ;
        RECT 6.124 0.804 8.596 0.836 ;
  LAYER M2 ;
        RECT 6.124 0.868 8.596 0.9 ;
  LAYER M2 ;
        RECT 6.124 0.932 8.596 0.964 ;
  LAYER M2 ;
        RECT 6.124 0.996 8.596 1.028 ;
  LAYER M2 ;
        RECT 6.124 1.06 8.596 1.092 ;
  LAYER M2 ;
        RECT 6.124 1.124 8.596 1.156 ;
  LAYER M2 ;
        RECT 6.124 1.188 8.596 1.22 ;
  LAYER M2 ;
        RECT 6.124 1.252 8.596 1.284 ;
  LAYER M2 ;
        RECT 6.124 1.316 8.596 1.348 ;
  LAYER M2 ;
        RECT 6.124 1.38 8.596 1.412 ;
  LAYER M2 ;
        RECT 6.124 1.444 8.596 1.476 ;
  LAYER M2 ;
        RECT 6.124 1.508 8.596 1.54 ;
  LAYER M2 ;
        RECT 6.124 1.572 8.596 1.604 ;
  LAYER M2 ;
        RECT 6.124 1.636 8.596 1.668 ;
  LAYER M2 ;
        RECT 6.124 1.7 8.596 1.732 ;
  LAYER M2 ;
        RECT 6.124 1.764 8.596 1.796 ;
  LAYER M2 ;
        RECT 6.124 1.828 8.596 1.86 ;
  LAYER M2 ;
        RECT 6.124 1.892 8.596 1.924 ;
  LAYER M2 ;
        RECT 6.124 1.956 8.596 1.988 ;
  LAYER M2 ;
        RECT 6.124 2.02 8.596 2.052 ;
  LAYER M2 ;
        RECT 6.124 2.084 8.596 2.116 ;
  LAYER M2 ;
        RECT 6.124 2.148 8.596 2.18 ;
  LAYER M2 ;
        RECT 6.124 2.212 8.596 2.244 ;
  LAYER M2 ;
        RECT 6.124 2.276 8.596 2.308 ;
  LAYER M2 ;
        RECT 6.124 2.34 8.596 2.372 ;
  LAYER M2 ;
        RECT 6.124 2.404 8.596 2.436 ;
  LAYER M2 ;
        RECT 6.124 2.468 8.596 2.5 ;
  LAYER M2 ;
        RECT 6.124 2.532 8.596 2.564 ;
  LAYER M2 ;
        RECT 6.124 2.596 8.596 2.628 ;
  LAYER M2 ;
        RECT 6.124 2.66 8.596 2.692 ;
  LAYER M2 ;
        RECT 6.124 2.724 8.596 2.756 ;
  LAYER M2 ;
        RECT 6.124 2.788 8.596 2.82 ;
  LAYER M2 ;
        RECT 6.124 2.852 8.596 2.884 ;
  LAYER M2 ;
        RECT 6.124 2.916 8.596 2.948 ;
  LAYER M2 ;
        RECT 6.124 2.98 8.596 3.012 ;
  LAYER M2 ;
        RECT 6.124 3.044 8.596 3.076 ;
  LAYER M3 ;
        RECT 6.144 0.72 6.176 3.228 ;
  LAYER M3 ;
        RECT 6.208 0.72 6.24 3.228 ;
  LAYER M3 ;
        RECT 6.272 0.72 6.304 3.228 ;
  LAYER M3 ;
        RECT 6.336 0.72 6.368 3.228 ;
  LAYER M3 ;
        RECT 6.4 0.72 6.432 3.228 ;
  LAYER M3 ;
        RECT 6.464 0.72 6.496 3.228 ;
  LAYER M3 ;
        RECT 6.528 0.72 6.56 3.228 ;
  LAYER M3 ;
        RECT 6.592 0.72 6.624 3.228 ;
  LAYER M3 ;
        RECT 6.656 0.72 6.688 3.228 ;
  LAYER M3 ;
        RECT 6.72 0.72 6.752 3.228 ;
  LAYER M3 ;
        RECT 6.784 0.72 6.816 3.228 ;
  LAYER M3 ;
        RECT 6.848 0.72 6.88 3.228 ;
  LAYER M3 ;
        RECT 6.912 0.72 6.944 3.228 ;
  LAYER M3 ;
        RECT 6.976 0.72 7.008 3.228 ;
  LAYER M3 ;
        RECT 7.04 0.72 7.072 3.228 ;
  LAYER M3 ;
        RECT 7.104 0.72 7.136 3.228 ;
  LAYER M3 ;
        RECT 7.168 0.72 7.2 3.228 ;
  LAYER M3 ;
        RECT 7.232 0.72 7.264 3.228 ;
  LAYER M3 ;
        RECT 7.296 0.72 7.328 3.228 ;
  LAYER M3 ;
        RECT 7.36 0.72 7.392 3.228 ;
  LAYER M3 ;
        RECT 7.424 0.72 7.456 3.228 ;
  LAYER M3 ;
        RECT 7.488 0.72 7.52 3.228 ;
  LAYER M3 ;
        RECT 7.552 0.72 7.584 3.228 ;
  LAYER M3 ;
        RECT 7.616 0.72 7.648 3.228 ;
  LAYER M3 ;
        RECT 7.68 0.72 7.712 3.228 ;
  LAYER M3 ;
        RECT 7.744 0.72 7.776 3.228 ;
  LAYER M3 ;
        RECT 7.808 0.72 7.84 3.228 ;
  LAYER M3 ;
        RECT 7.872 0.72 7.904 3.228 ;
  LAYER M3 ;
        RECT 7.936 0.72 7.968 3.228 ;
  LAYER M3 ;
        RECT 8 0.72 8.032 3.228 ;
  LAYER M3 ;
        RECT 8.064 0.72 8.096 3.228 ;
  LAYER M3 ;
        RECT 8.128 0.72 8.16 3.228 ;
  LAYER M3 ;
        RECT 8.192 0.72 8.224 3.228 ;
  LAYER M3 ;
        RECT 8.256 0.72 8.288 3.228 ;
  LAYER M3 ;
        RECT 8.32 0.72 8.352 3.228 ;
  LAYER M3 ;
        RECT 8.384 0.72 8.416 3.228 ;
  LAYER M3 ;
        RECT 8.448 0.72 8.48 3.228 ;
  LAYER M3 ;
        RECT 8.544 0.72 8.576 3.228 ;
  LAYER M1 ;
        RECT 6.159 0.756 6.161 3.192 ;
  LAYER M1 ;
        RECT 6.239 0.756 6.241 3.192 ;
  LAYER M1 ;
        RECT 6.319 0.756 6.321 3.192 ;
  LAYER M1 ;
        RECT 6.399 0.756 6.401 3.192 ;
  LAYER M1 ;
        RECT 6.479 0.756 6.481 3.192 ;
  LAYER M1 ;
        RECT 6.559 0.756 6.561 3.192 ;
  LAYER M1 ;
        RECT 6.639 0.756 6.641 3.192 ;
  LAYER M1 ;
        RECT 6.719 0.756 6.721 3.192 ;
  LAYER M1 ;
        RECT 6.799 0.756 6.801 3.192 ;
  LAYER M1 ;
        RECT 6.879 0.756 6.881 3.192 ;
  LAYER M1 ;
        RECT 6.959 0.756 6.961 3.192 ;
  LAYER M1 ;
        RECT 7.039 0.756 7.041 3.192 ;
  LAYER M1 ;
        RECT 7.119 0.756 7.121 3.192 ;
  LAYER M1 ;
        RECT 7.199 0.756 7.201 3.192 ;
  LAYER M1 ;
        RECT 7.279 0.756 7.281 3.192 ;
  LAYER M1 ;
        RECT 7.359 0.756 7.361 3.192 ;
  LAYER M1 ;
        RECT 7.439 0.756 7.441 3.192 ;
  LAYER M1 ;
        RECT 7.519 0.756 7.521 3.192 ;
  LAYER M1 ;
        RECT 7.599 0.756 7.601 3.192 ;
  LAYER M1 ;
        RECT 7.679 0.756 7.681 3.192 ;
  LAYER M1 ;
        RECT 7.759 0.756 7.761 3.192 ;
  LAYER M1 ;
        RECT 7.839 0.756 7.841 3.192 ;
  LAYER M1 ;
        RECT 7.919 0.756 7.921 3.192 ;
  LAYER M1 ;
        RECT 7.999 0.756 8.001 3.192 ;
  LAYER M1 ;
        RECT 8.079 0.756 8.081 3.192 ;
  LAYER M1 ;
        RECT 8.159 0.756 8.161 3.192 ;
  LAYER M1 ;
        RECT 8.239 0.756 8.241 3.192 ;
  LAYER M1 ;
        RECT 8.319 0.756 8.321 3.192 ;
  LAYER M1 ;
        RECT 8.399 0.756 8.401 3.192 ;
  LAYER M1 ;
        RECT 8.479 0.756 8.481 3.192 ;
  LAYER M2 ;
        RECT 6.16 0.755 8.56 0.757 ;
  LAYER M2 ;
        RECT 6.16 0.839 8.56 0.841 ;
  LAYER M2 ;
        RECT 6.16 0.923 8.56 0.925 ;
  LAYER M2 ;
        RECT 6.16 1.007 8.56 1.009 ;
  LAYER M2 ;
        RECT 6.16 1.091 8.56 1.093 ;
  LAYER M2 ;
        RECT 6.16 1.175 8.56 1.177 ;
  LAYER M2 ;
        RECT 6.16 1.259 8.56 1.261 ;
  LAYER M2 ;
        RECT 6.16 1.343 8.56 1.345 ;
  LAYER M2 ;
        RECT 6.16 1.427 8.56 1.429 ;
  LAYER M2 ;
        RECT 6.16 1.511 8.56 1.513 ;
  LAYER M2 ;
        RECT 6.16 1.595 8.56 1.597 ;
  LAYER M2 ;
        RECT 6.16 1.679 8.56 1.681 ;
  LAYER M2 ;
        RECT 6.16 1.7625 8.56 1.7645 ;
  LAYER M2 ;
        RECT 6.16 1.847 8.56 1.849 ;
  LAYER M2 ;
        RECT 6.16 1.931 8.56 1.933 ;
  LAYER M2 ;
        RECT 6.16 2.015 8.56 2.017 ;
  LAYER M2 ;
        RECT 6.16 2.099 8.56 2.101 ;
  LAYER M2 ;
        RECT 6.16 2.183 8.56 2.185 ;
  LAYER M2 ;
        RECT 6.16 2.267 8.56 2.269 ;
  LAYER M2 ;
        RECT 6.16 2.351 8.56 2.353 ;
  LAYER M2 ;
        RECT 6.16 2.435 8.56 2.437 ;
  LAYER M2 ;
        RECT 6.16 2.519 8.56 2.521 ;
  LAYER M2 ;
        RECT 6.16 2.603 8.56 2.605 ;
  LAYER M2 ;
        RECT 6.16 2.687 8.56 2.689 ;
  LAYER M2 ;
        RECT 6.16 2.771 8.56 2.773 ;
  LAYER M2 ;
        RECT 6.16 2.855 8.56 2.857 ;
  LAYER M2 ;
        RECT 6.16 2.939 8.56 2.941 ;
  LAYER M2 ;
        RECT 6.16 3.023 8.56 3.025 ;
  LAYER M2 ;
        RECT 6.16 3.107 8.56 3.109 ;
  LAYER M1 ;
        RECT 6.144 3.66 6.176 6.168 ;
  LAYER M1 ;
        RECT 6.208 3.66 6.24 6.168 ;
  LAYER M1 ;
        RECT 6.272 3.66 6.304 6.168 ;
  LAYER M1 ;
        RECT 6.336 3.66 6.368 6.168 ;
  LAYER M1 ;
        RECT 6.4 3.66 6.432 6.168 ;
  LAYER M1 ;
        RECT 6.464 3.66 6.496 6.168 ;
  LAYER M1 ;
        RECT 6.528 3.66 6.56 6.168 ;
  LAYER M1 ;
        RECT 6.592 3.66 6.624 6.168 ;
  LAYER M1 ;
        RECT 6.656 3.66 6.688 6.168 ;
  LAYER M1 ;
        RECT 6.72 3.66 6.752 6.168 ;
  LAYER M1 ;
        RECT 6.784 3.66 6.816 6.168 ;
  LAYER M1 ;
        RECT 6.848 3.66 6.88 6.168 ;
  LAYER M1 ;
        RECT 6.912 3.66 6.944 6.168 ;
  LAYER M1 ;
        RECT 6.976 3.66 7.008 6.168 ;
  LAYER M1 ;
        RECT 7.04 3.66 7.072 6.168 ;
  LAYER M1 ;
        RECT 7.104 3.66 7.136 6.168 ;
  LAYER M1 ;
        RECT 7.168 3.66 7.2 6.168 ;
  LAYER M1 ;
        RECT 7.232 3.66 7.264 6.168 ;
  LAYER M1 ;
        RECT 7.296 3.66 7.328 6.168 ;
  LAYER M1 ;
        RECT 7.36 3.66 7.392 6.168 ;
  LAYER M1 ;
        RECT 7.424 3.66 7.456 6.168 ;
  LAYER M1 ;
        RECT 7.488 3.66 7.52 6.168 ;
  LAYER M1 ;
        RECT 7.552 3.66 7.584 6.168 ;
  LAYER M1 ;
        RECT 7.616 3.66 7.648 6.168 ;
  LAYER M1 ;
        RECT 7.68 3.66 7.712 6.168 ;
  LAYER M1 ;
        RECT 7.744 3.66 7.776 6.168 ;
  LAYER M1 ;
        RECT 7.808 3.66 7.84 6.168 ;
  LAYER M1 ;
        RECT 7.872 3.66 7.904 6.168 ;
  LAYER M1 ;
        RECT 7.936 3.66 7.968 6.168 ;
  LAYER M1 ;
        RECT 8 3.66 8.032 6.168 ;
  LAYER M1 ;
        RECT 8.064 3.66 8.096 6.168 ;
  LAYER M1 ;
        RECT 8.128 3.66 8.16 6.168 ;
  LAYER M1 ;
        RECT 8.192 3.66 8.224 6.168 ;
  LAYER M1 ;
        RECT 8.256 3.66 8.288 6.168 ;
  LAYER M1 ;
        RECT 8.32 3.66 8.352 6.168 ;
  LAYER M1 ;
        RECT 8.384 3.66 8.416 6.168 ;
  LAYER M1 ;
        RECT 8.448 3.66 8.48 6.168 ;
  LAYER M2 ;
        RECT 6.124 3.744 8.596 3.776 ;
  LAYER M2 ;
        RECT 6.124 3.808 8.596 3.84 ;
  LAYER M2 ;
        RECT 6.124 3.872 8.596 3.904 ;
  LAYER M2 ;
        RECT 6.124 3.936 8.596 3.968 ;
  LAYER M2 ;
        RECT 6.124 4 8.596 4.032 ;
  LAYER M2 ;
        RECT 6.124 4.064 8.596 4.096 ;
  LAYER M2 ;
        RECT 6.124 4.128 8.596 4.16 ;
  LAYER M2 ;
        RECT 6.124 4.192 8.596 4.224 ;
  LAYER M2 ;
        RECT 6.124 4.256 8.596 4.288 ;
  LAYER M2 ;
        RECT 6.124 4.32 8.596 4.352 ;
  LAYER M2 ;
        RECT 6.124 4.384 8.596 4.416 ;
  LAYER M2 ;
        RECT 6.124 4.448 8.596 4.48 ;
  LAYER M2 ;
        RECT 6.124 4.512 8.596 4.544 ;
  LAYER M2 ;
        RECT 6.124 4.576 8.596 4.608 ;
  LAYER M2 ;
        RECT 6.124 4.64 8.596 4.672 ;
  LAYER M2 ;
        RECT 6.124 4.704 8.596 4.736 ;
  LAYER M2 ;
        RECT 6.124 4.768 8.596 4.8 ;
  LAYER M2 ;
        RECT 6.124 4.832 8.596 4.864 ;
  LAYER M2 ;
        RECT 6.124 4.896 8.596 4.928 ;
  LAYER M2 ;
        RECT 6.124 4.96 8.596 4.992 ;
  LAYER M2 ;
        RECT 6.124 5.024 8.596 5.056 ;
  LAYER M2 ;
        RECT 6.124 5.088 8.596 5.12 ;
  LAYER M2 ;
        RECT 6.124 5.152 8.596 5.184 ;
  LAYER M2 ;
        RECT 6.124 5.216 8.596 5.248 ;
  LAYER M2 ;
        RECT 6.124 5.28 8.596 5.312 ;
  LAYER M2 ;
        RECT 6.124 5.344 8.596 5.376 ;
  LAYER M2 ;
        RECT 6.124 5.408 8.596 5.44 ;
  LAYER M2 ;
        RECT 6.124 5.472 8.596 5.504 ;
  LAYER M2 ;
        RECT 6.124 5.536 8.596 5.568 ;
  LAYER M2 ;
        RECT 6.124 5.6 8.596 5.632 ;
  LAYER M2 ;
        RECT 6.124 5.664 8.596 5.696 ;
  LAYER M2 ;
        RECT 6.124 5.728 8.596 5.76 ;
  LAYER M2 ;
        RECT 6.124 5.792 8.596 5.824 ;
  LAYER M2 ;
        RECT 6.124 5.856 8.596 5.888 ;
  LAYER M2 ;
        RECT 6.124 5.92 8.596 5.952 ;
  LAYER M2 ;
        RECT 6.124 5.984 8.596 6.016 ;
  LAYER M3 ;
        RECT 6.144 3.66 6.176 6.168 ;
  LAYER M3 ;
        RECT 6.208 3.66 6.24 6.168 ;
  LAYER M3 ;
        RECT 6.272 3.66 6.304 6.168 ;
  LAYER M3 ;
        RECT 6.336 3.66 6.368 6.168 ;
  LAYER M3 ;
        RECT 6.4 3.66 6.432 6.168 ;
  LAYER M3 ;
        RECT 6.464 3.66 6.496 6.168 ;
  LAYER M3 ;
        RECT 6.528 3.66 6.56 6.168 ;
  LAYER M3 ;
        RECT 6.592 3.66 6.624 6.168 ;
  LAYER M3 ;
        RECT 6.656 3.66 6.688 6.168 ;
  LAYER M3 ;
        RECT 6.72 3.66 6.752 6.168 ;
  LAYER M3 ;
        RECT 6.784 3.66 6.816 6.168 ;
  LAYER M3 ;
        RECT 6.848 3.66 6.88 6.168 ;
  LAYER M3 ;
        RECT 6.912 3.66 6.944 6.168 ;
  LAYER M3 ;
        RECT 6.976 3.66 7.008 6.168 ;
  LAYER M3 ;
        RECT 7.04 3.66 7.072 6.168 ;
  LAYER M3 ;
        RECT 7.104 3.66 7.136 6.168 ;
  LAYER M3 ;
        RECT 7.168 3.66 7.2 6.168 ;
  LAYER M3 ;
        RECT 7.232 3.66 7.264 6.168 ;
  LAYER M3 ;
        RECT 7.296 3.66 7.328 6.168 ;
  LAYER M3 ;
        RECT 7.36 3.66 7.392 6.168 ;
  LAYER M3 ;
        RECT 7.424 3.66 7.456 6.168 ;
  LAYER M3 ;
        RECT 7.488 3.66 7.52 6.168 ;
  LAYER M3 ;
        RECT 7.552 3.66 7.584 6.168 ;
  LAYER M3 ;
        RECT 7.616 3.66 7.648 6.168 ;
  LAYER M3 ;
        RECT 7.68 3.66 7.712 6.168 ;
  LAYER M3 ;
        RECT 7.744 3.66 7.776 6.168 ;
  LAYER M3 ;
        RECT 7.808 3.66 7.84 6.168 ;
  LAYER M3 ;
        RECT 7.872 3.66 7.904 6.168 ;
  LAYER M3 ;
        RECT 7.936 3.66 7.968 6.168 ;
  LAYER M3 ;
        RECT 8 3.66 8.032 6.168 ;
  LAYER M3 ;
        RECT 8.064 3.66 8.096 6.168 ;
  LAYER M3 ;
        RECT 8.128 3.66 8.16 6.168 ;
  LAYER M3 ;
        RECT 8.192 3.66 8.224 6.168 ;
  LAYER M3 ;
        RECT 8.256 3.66 8.288 6.168 ;
  LAYER M3 ;
        RECT 8.32 3.66 8.352 6.168 ;
  LAYER M3 ;
        RECT 8.384 3.66 8.416 6.168 ;
  LAYER M3 ;
        RECT 8.448 3.66 8.48 6.168 ;
  LAYER M3 ;
        RECT 8.544 3.66 8.576 6.168 ;
  LAYER M1 ;
        RECT 6.159 3.696 6.161 6.132 ;
  LAYER M1 ;
        RECT 6.239 3.696 6.241 6.132 ;
  LAYER M1 ;
        RECT 6.319 3.696 6.321 6.132 ;
  LAYER M1 ;
        RECT 6.399 3.696 6.401 6.132 ;
  LAYER M1 ;
        RECT 6.479 3.696 6.481 6.132 ;
  LAYER M1 ;
        RECT 6.559 3.696 6.561 6.132 ;
  LAYER M1 ;
        RECT 6.639 3.696 6.641 6.132 ;
  LAYER M1 ;
        RECT 6.719 3.696 6.721 6.132 ;
  LAYER M1 ;
        RECT 6.799 3.696 6.801 6.132 ;
  LAYER M1 ;
        RECT 6.879 3.696 6.881 6.132 ;
  LAYER M1 ;
        RECT 6.959 3.696 6.961 6.132 ;
  LAYER M1 ;
        RECT 7.039 3.696 7.041 6.132 ;
  LAYER M1 ;
        RECT 7.119 3.696 7.121 6.132 ;
  LAYER M1 ;
        RECT 7.199 3.696 7.201 6.132 ;
  LAYER M1 ;
        RECT 7.279 3.696 7.281 6.132 ;
  LAYER M1 ;
        RECT 7.359 3.696 7.361 6.132 ;
  LAYER M1 ;
        RECT 7.439 3.696 7.441 6.132 ;
  LAYER M1 ;
        RECT 7.519 3.696 7.521 6.132 ;
  LAYER M1 ;
        RECT 7.599 3.696 7.601 6.132 ;
  LAYER M1 ;
        RECT 7.679 3.696 7.681 6.132 ;
  LAYER M1 ;
        RECT 7.759 3.696 7.761 6.132 ;
  LAYER M1 ;
        RECT 7.839 3.696 7.841 6.132 ;
  LAYER M1 ;
        RECT 7.919 3.696 7.921 6.132 ;
  LAYER M1 ;
        RECT 7.999 3.696 8.001 6.132 ;
  LAYER M1 ;
        RECT 8.079 3.696 8.081 6.132 ;
  LAYER M1 ;
        RECT 8.159 3.696 8.161 6.132 ;
  LAYER M1 ;
        RECT 8.239 3.696 8.241 6.132 ;
  LAYER M1 ;
        RECT 8.319 3.696 8.321 6.132 ;
  LAYER M1 ;
        RECT 8.399 3.696 8.401 6.132 ;
  LAYER M1 ;
        RECT 8.479 3.696 8.481 6.132 ;
  LAYER M2 ;
        RECT 6.16 3.695 8.56 3.697 ;
  LAYER M2 ;
        RECT 6.16 3.779 8.56 3.781 ;
  LAYER M2 ;
        RECT 6.16 3.863 8.56 3.865 ;
  LAYER M2 ;
        RECT 6.16 3.947 8.56 3.949 ;
  LAYER M2 ;
        RECT 6.16 4.031 8.56 4.033 ;
  LAYER M2 ;
        RECT 6.16 4.115 8.56 4.117 ;
  LAYER M2 ;
        RECT 6.16 4.199 8.56 4.201 ;
  LAYER M2 ;
        RECT 6.16 4.283 8.56 4.285 ;
  LAYER M2 ;
        RECT 6.16 4.367 8.56 4.369 ;
  LAYER M2 ;
        RECT 6.16 4.451 8.56 4.453 ;
  LAYER M2 ;
        RECT 6.16 4.535 8.56 4.537 ;
  LAYER M2 ;
        RECT 6.16 4.619 8.56 4.621 ;
  LAYER M2 ;
        RECT 6.16 4.7025 8.56 4.7045 ;
  LAYER M2 ;
        RECT 6.16 4.787 8.56 4.789 ;
  LAYER M2 ;
        RECT 6.16 4.871 8.56 4.873 ;
  LAYER M2 ;
        RECT 6.16 4.955 8.56 4.957 ;
  LAYER M2 ;
        RECT 6.16 5.039 8.56 5.041 ;
  LAYER M2 ;
        RECT 6.16 5.123 8.56 5.125 ;
  LAYER M2 ;
        RECT 6.16 5.207 8.56 5.209 ;
  LAYER M2 ;
        RECT 6.16 5.291 8.56 5.293 ;
  LAYER M2 ;
        RECT 6.16 5.375 8.56 5.377 ;
  LAYER M2 ;
        RECT 6.16 5.459 8.56 5.461 ;
  LAYER M2 ;
        RECT 6.16 5.543 8.56 5.545 ;
  LAYER M2 ;
        RECT 6.16 5.627 8.56 5.629 ;
  LAYER M2 ;
        RECT 6.16 5.711 8.56 5.713 ;
  LAYER M2 ;
        RECT 6.16 5.795 8.56 5.797 ;
  LAYER M2 ;
        RECT 6.16 5.879 8.56 5.881 ;
  LAYER M2 ;
        RECT 6.16 5.963 8.56 5.965 ;
  LAYER M2 ;
        RECT 6.16 6.047 8.56 6.049 ;
  LAYER M1 ;
        RECT 6.144 6.6 6.176 9.108 ;
  LAYER M1 ;
        RECT 6.208 6.6 6.24 9.108 ;
  LAYER M1 ;
        RECT 6.272 6.6 6.304 9.108 ;
  LAYER M1 ;
        RECT 6.336 6.6 6.368 9.108 ;
  LAYER M1 ;
        RECT 6.4 6.6 6.432 9.108 ;
  LAYER M1 ;
        RECT 6.464 6.6 6.496 9.108 ;
  LAYER M1 ;
        RECT 6.528 6.6 6.56 9.108 ;
  LAYER M1 ;
        RECT 6.592 6.6 6.624 9.108 ;
  LAYER M1 ;
        RECT 6.656 6.6 6.688 9.108 ;
  LAYER M1 ;
        RECT 6.72 6.6 6.752 9.108 ;
  LAYER M1 ;
        RECT 6.784 6.6 6.816 9.108 ;
  LAYER M1 ;
        RECT 6.848 6.6 6.88 9.108 ;
  LAYER M1 ;
        RECT 6.912 6.6 6.944 9.108 ;
  LAYER M1 ;
        RECT 6.976 6.6 7.008 9.108 ;
  LAYER M1 ;
        RECT 7.04 6.6 7.072 9.108 ;
  LAYER M1 ;
        RECT 7.104 6.6 7.136 9.108 ;
  LAYER M1 ;
        RECT 7.168 6.6 7.2 9.108 ;
  LAYER M1 ;
        RECT 7.232 6.6 7.264 9.108 ;
  LAYER M1 ;
        RECT 7.296 6.6 7.328 9.108 ;
  LAYER M1 ;
        RECT 7.36 6.6 7.392 9.108 ;
  LAYER M1 ;
        RECT 7.424 6.6 7.456 9.108 ;
  LAYER M1 ;
        RECT 7.488 6.6 7.52 9.108 ;
  LAYER M1 ;
        RECT 7.552 6.6 7.584 9.108 ;
  LAYER M1 ;
        RECT 7.616 6.6 7.648 9.108 ;
  LAYER M1 ;
        RECT 7.68 6.6 7.712 9.108 ;
  LAYER M1 ;
        RECT 7.744 6.6 7.776 9.108 ;
  LAYER M1 ;
        RECT 7.808 6.6 7.84 9.108 ;
  LAYER M1 ;
        RECT 7.872 6.6 7.904 9.108 ;
  LAYER M1 ;
        RECT 7.936 6.6 7.968 9.108 ;
  LAYER M1 ;
        RECT 8 6.6 8.032 9.108 ;
  LAYER M1 ;
        RECT 8.064 6.6 8.096 9.108 ;
  LAYER M1 ;
        RECT 8.128 6.6 8.16 9.108 ;
  LAYER M1 ;
        RECT 8.192 6.6 8.224 9.108 ;
  LAYER M1 ;
        RECT 8.256 6.6 8.288 9.108 ;
  LAYER M1 ;
        RECT 8.32 6.6 8.352 9.108 ;
  LAYER M1 ;
        RECT 8.384 6.6 8.416 9.108 ;
  LAYER M1 ;
        RECT 8.448 6.6 8.48 9.108 ;
  LAYER M2 ;
        RECT 6.124 6.684 8.596 6.716 ;
  LAYER M2 ;
        RECT 6.124 6.748 8.596 6.78 ;
  LAYER M2 ;
        RECT 6.124 6.812 8.596 6.844 ;
  LAYER M2 ;
        RECT 6.124 6.876 8.596 6.908 ;
  LAYER M2 ;
        RECT 6.124 6.94 8.596 6.972 ;
  LAYER M2 ;
        RECT 6.124 7.004 8.596 7.036 ;
  LAYER M2 ;
        RECT 6.124 7.068 8.596 7.1 ;
  LAYER M2 ;
        RECT 6.124 7.132 8.596 7.164 ;
  LAYER M2 ;
        RECT 6.124 7.196 8.596 7.228 ;
  LAYER M2 ;
        RECT 6.124 7.26 8.596 7.292 ;
  LAYER M2 ;
        RECT 6.124 7.324 8.596 7.356 ;
  LAYER M2 ;
        RECT 6.124 7.388 8.596 7.42 ;
  LAYER M2 ;
        RECT 6.124 7.452 8.596 7.484 ;
  LAYER M2 ;
        RECT 6.124 7.516 8.596 7.548 ;
  LAYER M2 ;
        RECT 6.124 7.58 8.596 7.612 ;
  LAYER M2 ;
        RECT 6.124 7.644 8.596 7.676 ;
  LAYER M2 ;
        RECT 6.124 7.708 8.596 7.74 ;
  LAYER M2 ;
        RECT 6.124 7.772 8.596 7.804 ;
  LAYER M2 ;
        RECT 6.124 7.836 8.596 7.868 ;
  LAYER M2 ;
        RECT 6.124 7.9 8.596 7.932 ;
  LAYER M2 ;
        RECT 6.124 7.964 8.596 7.996 ;
  LAYER M2 ;
        RECT 6.124 8.028 8.596 8.06 ;
  LAYER M2 ;
        RECT 6.124 8.092 8.596 8.124 ;
  LAYER M2 ;
        RECT 6.124 8.156 8.596 8.188 ;
  LAYER M2 ;
        RECT 6.124 8.22 8.596 8.252 ;
  LAYER M2 ;
        RECT 6.124 8.284 8.596 8.316 ;
  LAYER M2 ;
        RECT 6.124 8.348 8.596 8.38 ;
  LAYER M2 ;
        RECT 6.124 8.412 8.596 8.444 ;
  LAYER M2 ;
        RECT 6.124 8.476 8.596 8.508 ;
  LAYER M2 ;
        RECT 6.124 8.54 8.596 8.572 ;
  LAYER M2 ;
        RECT 6.124 8.604 8.596 8.636 ;
  LAYER M2 ;
        RECT 6.124 8.668 8.596 8.7 ;
  LAYER M2 ;
        RECT 6.124 8.732 8.596 8.764 ;
  LAYER M2 ;
        RECT 6.124 8.796 8.596 8.828 ;
  LAYER M2 ;
        RECT 6.124 8.86 8.596 8.892 ;
  LAYER M2 ;
        RECT 6.124 8.924 8.596 8.956 ;
  LAYER M3 ;
        RECT 6.144 6.6 6.176 9.108 ;
  LAYER M3 ;
        RECT 6.208 6.6 6.24 9.108 ;
  LAYER M3 ;
        RECT 6.272 6.6 6.304 9.108 ;
  LAYER M3 ;
        RECT 6.336 6.6 6.368 9.108 ;
  LAYER M3 ;
        RECT 6.4 6.6 6.432 9.108 ;
  LAYER M3 ;
        RECT 6.464 6.6 6.496 9.108 ;
  LAYER M3 ;
        RECT 6.528 6.6 6.56 9.108 ;
  LAYER M3 ;
        RECT 6.592 6.6 6.624 9.108 ;
  LAYER M3 ;
        RECT 6.656 6.6 6.688 9.108 ;
  LAYER M3 ;
        RECT 6.72 6.6 6.752 9.108 ;
  LAYER M3 ;
        RECT 6.784 6.6 6.816 9.108 ;
  LAYER M3 ;
        RECT 6.848 6.6 6.88 9.108 ;
  LAYER M3 ;
        RECT 6.912 6.6 6.944 9.108 ;
  LAYER M3 ;
        RECT 6.976 6.6 7.008 9.108 ;
  LAYER M3 ;
        RECT 7.04 6.6 7.072 9.108 ;
  LAYER M3 ;
        RECT 7.104 6.6 7.136 9.108 ;
  LAYER M3 ;
        RECT 7.168 6.6 7.2 9.108 ;
  LAYER M3 ;
        RECT 7.232 6.6 7.264 9.108 ;
  LAYER M3 ;
        RECT 7.296 6.6 7.328 9.108 ;
  LAYER M3 ;
        RECT 7.36 6.6 7.392 9.108 ;
  LAYER M3 ;
        RECT 7.424 6.6 7.456 9.108 ;
  LAYER M3 ;
        RECT 7.488 6.6 7.52 9.108 ;
  LAYER M3 ;
        RECT 7.552 6.6 7.584 9.108 ;
  LAYER M3 ;
        RECT 7.616 6.6 7.648 9.108 ;
  LAYER M3 ;
        RECT 7.68 6.6 7.712 9.108 ;
  LAYER M3 ;
        RECT 7.744 6.6 7.776 9.108 ;
  LAYER M3 ;
        RECT 7.808 6.6 7.84 9.108 ;
  LAYER M3 ;
        RECT 7.872 6.6 7.904 9.108 ;
  LAYER M3 ;
        RECT 7.936 6.6 7.968 9.108 ;
  LAYER M3 ;
        RECT 8 6.6 8.032 9.108 ;
  LAYER M3 ;
        RECT 8.064 6.6 8.096 9.108 ;
  LAYER M3 ;
        RECT 8.128 6.6 8.16 9.108 ;
  LAYER M3 ;
        RECT 8.192 6.6 8.224 9.108 ;
  LAYER M3 ;
        RECT 8.256 6.6 8.288 9.108 ;
  LAYER M3 ;
        RECT 8.32 6.6 8.352 9.108 ;
  LAYER M3 ;
        RECT 8.384 6.6 8.416 9.108 ;
  LAYER M3 ;
        RECT 8.448 6.6 8.48 9.108 ;
  LAYER M3 ;
        RECT 8.544 6.6 8.576 9.108 ;
  LAYER M1 ;
        RECT 6.159 6.636 6.161 9.072 ;
  LAYER M1 ;
        RECT 6.239 6.636 6.241 9.072 ;
  LAYER M1 ;
        RECT 6.319 6.636 6.321 9.072 ;
  LAYER M1 ;
        RECT 6.399 6.636 6.401 9.072 ;
  LAYER M1 ;
        RECT 6.479 6.636 6.481 9.072 ;
  LAYER M1 ;
        RECT 6.559 6.636 6.561 9.072 ;
  LAYER M1 ;
        RECT 6.639 6.636 6.641 9.072 ;
  LAYER M1 ;
        RECT 6.719 6.636 6.721 9.072 ;
  LAYER M1 ;
        RECT 6.799 6.636 6.801 9.072 ;
  LAYER M1 ;
        RECT 6.879 6.636 6.881 9.072 ;
  LAYER M1 ;
        RECT 6.959 6.636 6.961 9.072 ;
  LAYER M1 ;
        RECT 7.039 6.636 7.041 9.072 ;
  LAYER M1 ;
        RECT 7.119 6.636 7.121 9.072 ;
  LAYER M1 ;
        RECT 7.199 6.636 7.201 9.072 ;
  LAYER M1 ;
        RECT 7.279 6.636 7.281 9.072 ;
  LAYER M1 ;
        RECT 7.359 6.636 7.361 9.072 ;
  LAYER M1 ;
        RECT 7.439 6.636 7.441 9.072 ;
  LAYER M1 ;
        RECT 7.519 6.636 7.521 9.072 ;
  LAYER M1 ;
        RECT 7.599 6.636 7.601 9.072 ;
  LAYER M1 ;
        RECT 7.679 6.636 7.681 9.072 ;
  LAYER M1 ;
        RECT 7.759 6.636 7.761 9.072 ;
  LAYER M1 ;
        RECT 7.839 6.636 7.841 9.072 ;
  LAYER M1 ;
        RECT 7.919 6.636 7.921 9.072 ;
  LAYER M1 ;
        RECT 7.999 6.636 8.001 9.072 ;
  LAYER M1 ;
        RECT 8.079 6.636 8.081 9.072 ;
  LAYER M1 ;
        RECT 8.159 6.636 8.161 9.072 ;
  LAYER M1 ;
        RECT 8.239 6.636 8.241 9.072 ;
  LAYER M1 ;
        RECT 8.319 6.636 8.321 9.072 ;
  LAYER M1 ;
        RECT 8.399 6.636 8.401 9.072 ;
  LAYER M1 ;
        RECT 8.479 6.636 8.481 9.072 ;
  LAYER M2 ;
        RECT 6.16 6.635 8.56 6.637 ;
  LAYER M2 ;
        RECT 6.16 6.719 8.56 6.721 ;
  LAYER M2 ;
        RECT 6.16 6.803 8.56 6.805 ;
  LAYER M2 ;
        RECT 6.16 6.887 8.56 6.889 ;
  LAYER M2 ;
        RECT 6.16 6.971 8.56 6.973 ;
  LAYER M2 ;
        RECT 6.16 7.055 8.56 7.057 ;
  LAYER M2 ;
        RECT 6.16 7.139 8.56 7.141 ;
  LAYER M2 ;
        RECT 6.16 7.223 8.56 7.225 ;
  LAYER M2 ;
        RECT 6.16 7.307 8.56 7.309 ;
  LAYER M2 ;
        RECT 6.16 7.391 8.56 7.393 ;
  LAYER M2 ;
        RECT 6.16 7.475 8.56 7.477 ;
  LAYER M2 ;
        RECT 6.16 7.559 8.56 7.561 ;
  LAYER M2 ;
        RECT 6.16 7.6425 8.56 7.6445 ;
  LAYER M2 ;
        RECT 6.16 7.727 8.56 7.729 ;
  LAYER M2 ;
        RECT 6.16 7.811 8.56 7.813 ;
  LAYER M2 ;
        RECT 6.16 7.895 8.56 7.897 ;
  LAYER M2 ;
        RECT 6.16 7.979 8.56 7.981 ;
  LAYER M2 ;
        RECT 6.16 8.063 8.56 8.065 ;
  LAYER M2 ;
        RECT 6.16 8.147 8.56 8.149 ;
  LAYER M2 ;
        RECT 6.16 8.231 8.56 8.233 ;
  LAYER M2 ;
        RECT 6.16 8.315 8.56 8.317 ;
  LAYER M2 ;
        RECT 6.16 8.399 8.56 8.401 ;
  LAYER M2 ;
        RECT 6.16 8.483 8.56 8.485 ;
  LAYER M2 ;
        RECT 6.16 8.567 8.56 8.569 ;
  LAYER M2 ;
        RECT 6.16 8.651 8.56 8.653 ;
  LAYER M2 ;
        RECT 6.16 8.735 8.56 8.737 ;
  LAYER M2 ;
        RECT 6.16 8.819 8.56 8.821 ;
  LAYER M2 ;
        RECT 6.16 8.903 8.56 8.905 ;
  LAYER M2 ;
        RECT 6.16 8.987 8.56 8.989 ;
  LAYER M1 ;
        RECT 6.144 9.54 6.176 12.048 ;
  LAYER M1 ;
        RECT 6.208 9.54 6.24 12.048 ;
  LAYER M1 ;
        RECT 6.272 9.54 6.304 12.048 ;
  LAYER M1 ;
        RECT 6.336 9.54 6.368 12.048 ;
  LAYER M1 ;
        RECT 6.4 9.54 6.432 12.048 ;
  LAYER M1 ;
        RECT 6.464 9.54 6.496 12.048 ;
  LAYER M1 ;
        RECT 6.528 9.54 6.56 12.048 ;
  LAYER M1 ;
        RECT 6.592 9.54 6.624 12.048 ;
  LAYER M1 ;
        RECT 6.656 9.54 6.688 12.048 ;
  LAYER M1 ;
        RECT 6.72 9.54 6.752 12.048 ;
  LAYER M1 ;
        RECT 6.784 9.54 6.816 12.048 ;
  LAYER M1 ;
        RECT 6.848 9.54 6.88 12.048 ;
  LAYER M1 ;
        RECT 6.912 9.54 6.944 12.048 ;
  LAYER M1 ;
        RECT 6.976 9.54 7.008 12.048 ;
  LAYER M1 ;
        RECT 7.04 9.54 7.072 12.048 ;
  LAYER M1 ;
        RECT 7.104 9.54 7.136 12.048 ;
  LAYER M1 ;
        RECT 7.168 9.54 7.2 12.048 ;
  LAYER M1 ;
        RECT 7.232 9.54 7.264 12.048 ;
  LAYER M1 ;
        RECT 7.296 9.54 7.328 12.048 ;
  LAYER M1 ;
        RECT 7.36 9.54 7.392 12.048 ;
  LAYER M1 ;
        RECT 7.424 9.54 7.456 12.048 ;
  LAYER M1 ;
        RECT 7.488 9.54 7.52 12.048 ;
  LAYER M1 ;
        RECT 7.552 9.54 7.584 12.048 ;
  LAYER M1 ;
        RECT 7.616 9.54 7.648 12.048 ;
  LAYER M1 ;
        RECT 7.68 9.54 7.712 12.048 ;
  LAYER M1 ;
        RECT 7.744 9.54 7.776 12.048 ;
  LAYER M1 ;
        RECT 7.808 9.54 7.84 12.048 ;
  LAYER M1 ;
        RECT 7.872 9.54 7.904 12.048 ;
  LAYER M1 ;
        RECT 7.936 9.54 7.968 12.048 ;
  LAYER M1 ;
        RECT 8 9.54 8.032 12.048 ;
  LAYER M1 ;
        RECT 8.064 9.54 8.096 12.048 ;
  LAYER M1 ;
        RECT 8.128 9.54 8.16 12.048 ;
  LAYER M1 ;
        RECT 8.192 9.54 8.224 12.048 ;
  LAYER M1 ;
        RECT 8.256 9.54 8.288 12.048 ;
  LAYER M1 ;
        RECT 8.32 9.54 8.352 12.048 ;
  LAYER M1 ;
        RECT 8.384 9.54 8.416 12.048 ;
  LAYER M1 ;
        RECT 8.448 9.54 8.48 12.048 ;
  LAYER M2 ;
        RECT 6.124 9.624 8.596 9.656 ;
  LAYER M2 ;
        RECT 6.124 9.688 8.596 9.72 ;
  LAYER M2 ;
        RECT 6.124 9.752 8.596 9.784 ;
  LAYER M2 ;
        RECT 6.124 9.816 8.596 9.848 ;
  LAYER M2 ;
        RECT 6.124 9.88 8.596 9.912 ;
  LAYER M2 ;
        RECT 6.124 9.944 8.596 9.976 ;
  LAYER M2 ;
        RECT 6.124 10.008 8.596 10.04 ;
  LAYER M2 ;
        RECT 6.124 10.072 8.596 10.104 ;
  LAYER M2 ;
        RECT 6.124 10.136 8.596 10.168 ;
  LAYER M2 ;
        RECT 6.124 10.2 8.596 10.232 ;
  LAYER M2 ;
        RECT 6.124 10.264 8.596 10.296 ;
  LAYER M2 ;
        RECT 6.124 10.328 8.596 10.36 ;
  LAYER M2 ;
        RECT 6.124 10.392 8.596 10.424 ;
  LAYER M2 ;
        RECT 6.124 10.456 8.596 10.488 ;
  LAYER M2 ;
        RECT 6.124 10.52 8.596 10.552 ;
  LAYER M2 ;
        RECT 6.124 10.584 8.596 10.616 ;
  LAYER M2 ;
        RECT 6.124 10.648 8.596 10.68 ;
  LAYER M2 ;
        RECT 6.124 10.712 8.596 10.744 ;
  LAYER M2 ;
        RECT 6.124 10.776 8.596 10.808 ;
  LAYER M2 ;
        RECT 6.124 10.84 8.596 10.872 ;
  LAYER M2 ;
        RECT 6.124 10.904 8.596 10.936 ;
  LAYER M2 ;
        RECT 6.124 10.968 8.596 11 ;
  LAYER M2 ;
        RECT 6.124 11.032 8.596 11.064 ;
  LAYER M2 ;
        RECT 6.124 11.096 8.596 11.128 ;
  LAYER M2 ;
        RECT 6.124 11.16 8.596 11.192 ;
  LAYER M2 ;
        RECT 6.124 11.224 8.596 11.256 ;
  LAYER M2 ;
        RECT 6.124 11.288 8.596 11.32 ;
  LAYER M2 ;
        RECT 6.124 11.352 8.596 11.384 ;
  LAYER M2 ;
        RECT 6.124 11.416 8.596 11.448 ;
  LAYER M2 ;
        RECT 6.124 11.48 8.596 11.512 ;
  LAYER M2 ;
        RECT 6.124 11.544 8.596 11.576 ;
  LAYER M2 ;
        RECT 6.124 11.608 8.596 11.64 ;
  LAYER M2 ;
        RECT 6.124 11.672 8.596 11.704 ;
  LAYER M2 ;
        RECT 6.124 11.736 8.596 11.768 ;
  LAYER M2 ;
        RECT 6.124 11.8 8.596 11.832 ;
  LAYER M2 ;
        RECT 6.124 11.864 8.596 11.896 ;
  LAYER M3 ;
        RECT 6.144 9.54 6.176 12.048 ;
  LAYER M3 ;
        RECT 6.208 9.54 6.24 12.048 ;
  LAYER M3 ;
        RECT 6.272 9.54 6.304 12.048 ;
  LAYER M3 ;
        RECT 6.336 9.54 6.368 12.048 ;
  LAYER M3 ;
        RECT 6.4 9.54 6.432 12.048 ;
  LAYER M3 ;
        RECT 6.464 9.54 6.496 12.048 ;
  LAYER M3 ;
        RECT 6.528 9.54 6.56 12.048 ;
  LAYER M3 ;
        RECT 6.592 9.54 6.624 12.048 ;
  LAYER M3 ;
        RECT 6.656 9.54 6.688 12.048 ;
  LAYER M3 ;
        RECT 6.72 9.54 6.752 12.048 ;
  LAYER M3 ;
        RECT 6.784 9.54 6.816 12.048 ;
  LAYER M3 ;
        RECT 6.848 9.54 6.88 12.048 ;
  LAYER M3 ;
        RECT 6.912 9.54 6.944 12.048 ;
  LAYER M3 ;
        RECT 6.976 9.54 7.008 12.048 ;
  LAYER M3 ;
        RECT 7.04 9.54 7.072 12.048 ;
  LAYER M3 ;
        RECT 7.104 9.54 7.136 12.048 ;
  LAYER M3 ;
        RECT 7.168 9.54 7.2 12.048 ;
  LAYER M3 ;
        RECT 7.232 9.54 7.264 12.048 ;
  LAYER M3 ;
        RECT 7.296 9.54 7.328 12.048 ;
  LAYER M3 ;
        RECT 7.36 9.54 7.392 12.048 ;
  LAYER M3 ;
        RECT 7.424 9.54 7.456 12.048 ;
  LAYER M3 ;
        RECT 7.488 9.54 7.52 12.048 ;
  LAYER M3 ;
        RECT 7.552 9.54 7.584 12.048 ;
  LAYER M3 ;
        RECT 7.616 9.54 7.648 12.048 ;
  LAYER M3 ;
        RECT 7.68 9.54 7.712 12.048 ;
  LAYER M3 ;
        RECT 7.744 9.54 7.776 12.048 ;
  LAYER M3 ;
        RECT 7.808 9.54 7.84 12.048 ;
  LAYER M3 ;
        RECT 7.872 9.54 7.904 12.048 ;
  LAYER M3 ;
        RECT 7.936 9.54 7.968 12.048 ;
  LAYER M3 ;
        RECT 8 9.54 8.032 12.048 ;
  LAYER M3 ;
        RECT 8.064 9.54 8.096 12.048 ;
  LAYER M3 ;
        RECT 8.128 9.54 8.16 12.048 ;
  LAYER M3 ;
        RECT 8.192 9.54 8.224 12.048 ;
  LAYER M3 ;
        RECT 8.256 9.54 8.288 12.048 ;
  LAYER M3 ;
        RECT 8.32 9.54 8.352 12.048 ;
  LAYER M3 ;
        RECT 8.384 9.54 8.416 12.048 ;
  LAYER M3 ;
        RECT 8.448 9.54 8.48 12.048 ;
  LAYER M3 ;
        RECT 8.544 9.54 8.576 12.048 ;
  LAYER M1 ;
        RECT 6.159 9.576 6.161 12.012 ;
  LAYER M1 ;
        RECT 6.239 9.576 6.241 12.012 ;
  LAYER M1 ;
        RECT 6.319 9.576 6.321 12.012 ;
  LAYER M1 ;
        RECT 6.399 9.576 6.401 12.012 ;
  LAYER M1 ;
        RECT 6.479 9.576 6.481 12.012 ;
  LAYER M1 ;
        RECT 6.559 9.576 6.561 12.012 ;
  LAYER M1 ;
        RECT 6.639 9.576 6.641 12.012 ;
  LAYER M1 ;
        RECT 6.719 9.576 6.721 12.012 ;
  LAYER M1 ;
        RECT 6.799 9.576 6.801 12.012 ;
  LAYER M1 ;
        RECT 6.879 9.576 6.881 12.012 ;
  LAYER M1 ;
        RECT 6.959 9.576 6.961 12.012 ;
  LAYER M1 ;
        RECT 7.039 9.576 7.041 12.012 ;
  LAYER M1 ;
        RECT 7.119 9.576 7.121 12.012 ;
  LAYER M1 ;
        RECT 7.199 9.576 7.201 12.012 ;
  LAYER M1 ;
        RECT 7.279 9.576 7.281 12.012 ;
  LAYER M1 ;
        RECT 7.359 9.576 7.361 12.012 ;
  LAYER M1 ;
        RECT 7.439 9.576 7.441 12.012 ;
  LAYER M1 ;
        RECT 7.519 9.576 7.521 12.012 ;
  LAYER M1 ;
        RECT 7.599 9.576 7.601 12.012 ;
  LAYER M1 ;
        RECT 7.679 9.576 7.681 12.012 ;
  LAYER M1 ;
        RECT 7.759 9.576 7.761 12.012 ;
  LAYER M1 ;
        RECT 7.839 9.576 7.841 12.012 ;
  LAYER M1 ;
        RECT 7.919 9.576 7.921 12.012 ;
  LAYER M1 ;
        RECT 7.999 9.576 8.001 12.012 ;
  LAYER M1 ;
        RECT 8.079 9.576 8.081 12.012 ;
  LAYER M1 ;
        RECT 8.159 9.576 8.161 12.012 ;
  LAYER M1 ;
        RECT 8.239 9.576 8.241 12.012 ;
  LAYER M1 ;
        RECT 8.319 9.576 8.321 12.012 ;
  LAYER M1 ;
        RECT 8.399 9.576 8.401 12.012 ;
  LAYER M1 ;
        RECT 8.479 9.576 8.481 12.012 ;
  LAYER M2 ;
        RECT 6.16 9.575 8.56 9.577 ;
  LAYER M2 ;
        RECT 6.16 9.659 8.56 9.661 ;
  LAYER M2 ;
        RECT 6.16 9.743 8.56 9.745 ;
  LAYER M2 ;
        RECT 6.16 9.827 8.56 9.829 ;
  LAYER M2 ;
        RECT 6.16 9.911 8.56 9.913 ;
  LAYER M2 ;
        RECT 6.16 9.995 8.56 9.997 ;
  LAYER M2 ;
        RECT 6.16 10.079 8.56 10.081 ;
  LAYER M2 ;
        RECT 6.16 10.163 8.56 10.165 ;
  LAYER M2 ;
        RECT 6.16 10.247 8.56 10.249 ;
  LAYER M2 ;
        RECT 6.16 10.331 8.56 10.333 ;
  LAYER M2 ;
        RECT 6.16 10.415 8.56 10.417 ;
  LAYER M2 ;
        RECT 6.16 10.499 8.56 10.501 ;
  LAYER M2 ;
        RECT 6.16 10.5825 8.56 10.5845 ;
  LAYER M2 ;
        RECT 6.16 10.667 8.56 10.669 ;
  LAYER M2 ;
        RECT 6.16 10.751 8.56 10.753 ;
  LAYER M2 ;
        RECT 6.16 10.835 8.56 10.837 ;
  LAYER M2 ;
        RECT 6.16 10.919 8.56 10.921 ;
  LAYER M2 ;
        RECT 6.16 11.003 8.56 11.005 ;
  LAYER M2 ;
        RECT 6.16 11.087 8.56 11.089 ;
  LAYER M2 ;
        RECT 6.16 11.171 8.56 11.173 ;
  LAYER M2 ;
        RECT 6.16 11.255 8.56 11.257 ;
  LAYER M2 ;
        RECT 6.16 11.339 8.56 11.341 ;
  LAYER M2 ;
        RECT 6.16 11.423 8.56 11.425 ;
  LAYER M2 ;
        RECT 6.16 11.507 8.56 11.509 ;
  LAYER M2 ;
        RECT 6.16 11.591 8.56 11.593 ;
  LAYER M2 ;
        RECT 6.16 11.675 8.56 11.677 ;
  LAYER M2 ;
        RECT 6.16 11.759 8.56 11.761 ;
  LAYER M2 ;
        RECT 6.16 11.843 8.56 11.845 ;
  LAYER M2 ;
        RECT 6.16 11.927 8.56 11.929 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 14.988 ;
  LAYER M1 ;
        RECT 6.208 12.48 6.24 14.988 ;
  LAYER M1 ;
        RECT 6.272 12.48 6.304 14.988 ;
  LAYER M1 ;
        RECT 6.336 12.48 6.368 14.988 ;
  LAYER M1 ;
        RECT 6.4 12.48 6.432 14.988 ;
  LAYER M1 ;
        RECT 6.464 12.48 6.496 14.988 ;
  LAYER M1 ;
        RECT 6.528 12.48 6.56 14.988 ;
  LAYER M1 ;
        RECT 6.592 12.48 6.624 14.988 ;
  LAYER M1 ;
        RECT 6.656 12.48 6.688 14.988 ;
  LAYER M1 ;
        RECT 6.72 12.48 6.752 14.988 ;
  LAYER M1 ;
        RECT 6.784 12.48 6.816 14.988 ;
  LAYER M1 ;
        RECT 6.848 12.48 6.88 14.988 ;
  LAYER M1 ;
        RECT 6.912 12.48 6.944 14.988 ;
  LAYER M1 ;
        RECT 6.976 12.48 7.008 14.988 ;
  LAYER M1 ;
        RECT 7.04 12.48 7.072 14.988 ;
  LAYER M1 ;
        RECT 7.104 12.48 7.136 14.988 ;
  LAYER M1 ;
        RECT 7.168 12.48 7.2 14.988 ;
  LAYER M1 ;
        RECT 7.232 12.48 7.264 14.988 ;
  LAYER M1 ;
        RECT 7.296 12.48 7.328 14.988 ;
  LAYER M1 ;
        RECT 7.36 12.48 7.392 14.988 ;
  LAYER M1 ;
        RECT 7.424 12.48 7.456 14.988 ;
  LAYER M1 ;
        RECT 7.488 12.48 7.52 14.988 ;
  LAYER M1 ;
        RECT 7.552 12.48 7.584 14.988 ;
  LAYER M1 ;
        RECT 7.616 12.48 7.648 14.988 ;
  LAYER M1 ;
        RECT 7.68 12.48 7.712 14.988 ;
  LAYER M1 ;
        RECT 7.744 12.48 7.776 14.988 ;
  LAYER M1 ;
        RECT 7.808 12.48 7.84 14.988 ;
  LAYER M1 ;
        RECT 7.872 12.48 7.904 14.988 ;
  LAYER M1 ;
        RECT 7.936 12.48 7.968 14.988 ;
  LAYER M1 ;
        RECT 8 12.48 8.032 14.988 ;
  LAYER M1 ;
        RECT 8.064 12.48 8.096 14.988 ;
  LAYER M1 ;
        RECT 8.128 12.48 8.16 14.988 ;
  LAYER M1 ;
        RECT 8.192 12.48 8.224 14.988 ;
  LAYER M1 ;
        RECT 8.256 12.48 8.288 14.988 ;
  LAYER M1 ;
        RECT 8.32 12.48 8.352 14.988 ;
  LAYER M1 ;
        RECT 8.384 12.48 8.416 14.988 ;
  LAYER M1 ;
        RECT 8.448 12.48 8.48 14.988 ;
  LAYER M2 ;
        RECT 6.124 12.564 8.596 12.596 ;
  LAYER M2 ;
        RECT 6.124 12.628 8.596 12.66 ;
  LAYER M2 ;
        RECT 6.124 12.692 8.596 12.724 ;
  LAYER M2 ;
        RECT 6.124 12.756 8.596 12.788 ;
  LAYER M2 ;
        RECT 6.124 12.82 8.596 12.852 ;
  LAYER M2 ;
        RECT 6.124 12.884 8.596 12.916 ;
  LAYER M2 ;
        RECT 6.124 12.948 8.596 12.98 ;
  LAYER M2 ;
        RECT 6.124 13.012 8.596 13.044 ;
  LAYER M2 ;
        RECT 6.124 13.076 8.596 13.108 ;
  LAYER M2 ;
        RECT 6.124 13.14 8.596 13.172 ;
  LAYER M2 ;
        RECT 6.124 13.204 8.596 13.236 ;
  LAYER M2 ;
        RECT 6.124 13.268 8.596 13.3 ;
  LAYER M2 ;
        RECT 6.124 13.332 8.596 13.364 ;
  LAYER M2 ;
        RECT 6.124 13.396 8.596 13.428 ;
  LAYER M2 ;
        RECT 6.124 13.46 8.596 13.492 ;
  LAYER M2 ;
        RECT 6.124 13.524 8.596 13.556 ;
  LAYER M2 ;
        RECT 6.124 13.588 8.596 13.62 ;
  LAYER M2 ;
        RECT 6.124 13.652 8.596 13.684 ;
  LAYER M2 ;
        RECT 6.124 13.716 8.596 13.748 ;
  LAYER M2 ;
        RECT 6.124 13.78 8.596 13.812 ;
  LAYER M2 ;
        RECT 6.124 13.844 8.596 13.876 ;
  LAYER M2 ;
        RECT 6.124 13.908 8.596 13.94 ;
  LAYER M2 ;
        RECT 6.124 13.972 8.596 14.004 ;
  LAYER M2 ;
        RECT 6.124 14.036 8.596 14.068 ;
  LAYER M2 ;
        RECT 6.124 14.1 8.596 14.132 ;
  LAYER M2 ;
        RECT 6.124 14.164 8.596 14.196 ;
  LAYER M2 ;
        RECT 6.124 14.228 8.596 14.26 ;
  LAYER M2 ;
        RECT 6.124 14.292 8.596 14.324 ;
  LAYER M2 ;
        RECT 6.124 14.356 8.596 14.388 ;
  LAYER M2 ;
        RECT 6.124 14.42 8.596 14.452 ;
  LAYER M2 ;
        RECT 6.124 14.484 8.596 14.516 ;
  LAYER M2 ;
        RECT 6.124 14.548 8.596 14.58 ;
  LAYER M2 ;
        RECT 6.124 14.612 8.596 14.644 ;
  LAYER M2 ;
        RECT 6.124 14.676 8.596 14.708 ;
  LAYER M2 ;
        RECT 6.124 14.74 8.596 14.772 ;
  LAYER M2 ;
        RECT 6.124 14.804 8.596 14.836 ;
  LAYER M3 ;
        RECT 6.144 12.48 6.176 14.988 ;
  LAYER M3 ;
        RECT 6.208 12.48 6.24 14.988 ;
  LAYER M3 ;
        RECT 6.272 12.48 6.304 14.988 ;
  LAYER M3 ;
        RECT 6.336 12.48 6.368 14.988 ;
  LAYER M3 ;
        RECT 6.4 12.48 6.432 14.988 ;
  LAYER M3 ;
        RECT 6.464 12.48 6.496 14.988 ;
  LAYER M3 ;
        RECT 6.528 12.48 6.56 14.988 ;
  LAYER M3 ;
        RECT 6.592 12.48 6.624 14.988 ;
  LAYER M3 ;
        RECT 6.656 12.48 6.688 14.988 ;
  LAYER M3 ;
        RECT 6.72 12.48 6.752 14.988 ;
  LAYER M3 ;
        RECT 6.784 12.48 6.816 14.988 ;
  LAYER M3 ;
        RECT 6.848 12.48 6.88 14.988 ;
  LAYER M3 ;
        RECT 6.912 12.48 6.944 14.988 ;
  LAYER M3 ;
        RECT 6.976 12.48 7.008 14.988 ;
  LAYER M3 ;
        RECT 7.04 12.48 7.072 14.988 ;
  LAYER M3 ;
        RECT 7.104 12.48 7.136 14.988 ;
  LAYER M3 ;
        RECT 7.168 12.48 7.2 14.988 ;
  LAYER M3 ;
        RECT 7.232 12.48 7.264 14.988 ;
  LAYER M3 ;
        RECT 7.296 12.48 7.328 14.988 ;
  LAYER M3 ;
        RECT 7.36 12.48 7.392 14.988 ;
  LAYER M3 ;
        RECT 7.424 12.48 7.456 14.988 ;
  LAYER M3 ;
        RECT 7.488 12.48 7.52 14.988 ;
  LAYER M3 ;
        RECT 7.552 12.48 7.584 14.988 ;
  LAYER M3 ;
        RECT 7.616 12.48 7.648 14.988 ;
  LAYER M3 ;
        RECT 7.68 12.48 7.712 14.988 ;
  LAYER M3 ;
        RECT 7.744 12.48 7.776 14.988 ;
  LAYER M3 ;
        RECT 7.808 12.48 7.84 14.988 ;
  LAYER M3 ;
        RECT 7.872 12.48 7.904 14.988 ;
  LAYER M3 ;
        RECT 7.936 12.48 7.968 14.988 ;
  LAYER M3 ;
        RECT 8 12.48 8.032 14.988 ;
  LAYER M3 ;
        RECT 8.064 12.48 8.096 14.988 ;
  LAYER M3 ;
        RECT 8.128 12.48 8.16 14.988 ;
  LAYER M3 ;
        RECT 8.192 12.48 8.224 14.988 ;
  LAYER M3 ;
        RECT 8.256 12.48 8.288 14.988 ;
  LAYER M3 ;
        RECT 8.32 12.48 8.352 14.988 ;
  LAYER M3 ;
        RECT 8.384 12.48 8.416 14.988 ;
  LAYER M3 ;
        RECT 8.448 12.48 8.48 14.988 ;
  LAYER M3 ;
        RECT 8.544 12.48 8.576 14.988 ;
  LAYER M1 ;
        RECT 6.159 12.516 6.161 14.952 ;
  LAYER M1 ;
        RECT 6.239 12.516 6.241 14.952 ;
  LAYER M1 ;
        RECT 6.319 12.516 6.321 14.952 ;
  LAYER M1 ;
        RECT 6.399 12.516 6.401 14.952 ;
  LAYER M1 ;
        RECT 6.479 12.516 6.481 14.952 ;
  LAYER M1 ;
        RECT 6.559 12.516 6.561 14.952 ;
  LAYER M1 ;
        RECT 6.639 12.516 6.641 14.952 ;
  LAYER M1 ;
        RECT 6.719 12.516 6.721 14.952 ;
  LAYER M1 ;
        RECT 6.799 12.516 6.801 14.952 ;
  LAYER M1 ;
        RECT 6.879 12.516 6.881 14.952 ;
  LAYER M1 ;
        RECT 6.959 12.516 6.961 14.952 ;
  LAYER M1 ;
        RECT 7.039 12.516 7.041 14.952 ;
  LAYER M1 ;
        RECT 7.119 12.516 7.121 14.952 ;
  LAYER M1 ;
        RECT 7.199 12.516 7.201 14.952 ;
  LAYER M1 ;
        RECT 7.279 12.516 7.281 14.952 ;
  LAYER M1 ;
        RECT 7.359 12.516 7.361 14.952 ;
  LAYER M1 ;
        RECT 7.439 12.516 7.441 14.952 ;
  LAYER M1 ;
        RECT 7.519 12.516 7.521 14.952 ;
  LAYER M1 ;
        RECT 7.599 12.516 7.601 14.952 ;
  LAYER M1 ;
        RECT 7.679 12.516 7.681 14.952 ;
  LAYER M1 ;
        RECT 7.759 12.516 7.761 14.952 ;
  LAYER M1 ;
        RECT 7.839 12.516 7.841 14.952 ;
  LAYER M1 ;
        RECT 7.919 12.516 7.921 14.952 ;
  LAYER M1 ;
        RECT 7.999 12.516 8.001 14.952 ;
  LAYER M1 ;
        RECT 8.079 12.516 8.081 14.952 ;
  LAYER M1 ;
        RECT 8.159 12.516 8.161 14.952 ;
  LAYER M1 ;
        RECT 8.239 12.516 8.241 14.952 ;
  LAYER M1 ;
        RECT 8.319 12.516 8.321 14.952 ;
  LAYER M1 ;
        RECT 8.399 12.516 8.401 14.952 ;
  LAYER M1 ;
        RECT 8.479 12.516 8.481 14.952 ;
  LAYER M2 ;
        RECT 6.16 12.515 8.56 12.517 ;
  LAYER M2 ;
        RECT 6.16 12.599 8.56 12.601 ;
  LAYER M2 ;
        RECT 6.16 12.683 8.56 12.685 ;
  LAYER M2 ;
        RECT 6.16 12.767 8.56 12.769 ;
  LAYER M2 ;
        RECT 6.16 12.851 8.56 12.853 ;
  LAYER M2 ;
        RECT 6.16 12.935 8.56 12.937 ;
  LAYER M2 ;
        RECT 6.16 13.019 8.56 13.021 ;
  LAYER M2 ;
        RECT 6.16 13.103 8.56 13.105 ;
  LAYER M2 ;
        RECT 6.16 13.187 8.56 13.189 ;
  LAYER M2 ;
        RECT 6.16 13.271 8.56 13.273 ;
  LAYER M2 ;
        RECT 6.16 13.355 8.56 13.357 ;
  LAYER M2 ;
        RECT 6.16 13.439 8.56 13.441 ;
  LAYER M2 ;
        RECT 6.16 13.5225 8.56 13.5245 ;
  LAYER M2 ;
        RECT 6.16 13.607 8.56 13.609 ;
  LAYER M2 ;
        RECT 6.16 13.691 8.56 13.693 ;
  LAYER M2 ;
        RECT 6.16 13.775 8.56 13.777 ;
  LAYER M2 ;
        RECT 6.16 13.859 8.56 13.861 ;
  LAYER M2 ;
        RECT 6.16 13.943 8.56 13.945 ;
  LAYER M2 ;
        RECT 6.16 14.027 8.56 14.029 ;
  LAYER M2 ;
        RECT 6.16 14.111 8.56 14.113 ;
  LAYER M2 ;
        RECT 6.16 14.195 8.56 14.197 ;
  LAYER M2 ;
        RECT 6.16 14.279 8.56 14.281 ;
  LAYER M2 ;
        RECT 6.16 14.363 8.56 14.365 ;
  LAYER M2 ;
        RECT 6.16 14.447 8.56 14.449 ;
  LAYER M2 ;
        RECT 6.16 14.531 8.56 14.533 ;
  LAYER M2 ;
        RECT 6.16 14.615 8.56 14.617 ;
  LAYER M2 ;
        RECT 6.16 14.699 8.56 14.701 ;
  LAYER M2 ;
        RECT 6.16 14.783 8.56 14.785 ;
  LAYER M2 ;
        RECT 6.16 14.867 8.56 14.869 ;
  LAYER M1 ;
        RECT 6.144 15.42 6.176 17.928 ;
  LAYER M1 ;
        RECT 6.208 15.42 6.24 17.928 ;
  LAYER M1 ;
        RECT 6.272 15.42 6.304 17.928 ;
  LAYER M1 ;
        RECT 6.336 15.42 6.368 17.928 ;
  LAYER M1 ;
        RECT 6.4 15.42 6.432 17.928 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 17.928 ;
  LAYER M1 ;
        RECT 6.528 15.42 6.56 17.928 ;
  LAYER M1 ;
        RECT 6.592 15.42 6.624 17.928 ;
  LAYER M1 ;
        RECT 6.656 15.42 6.688 17.928 ;
  LAYER M1 ;
        RECT 6.72 15.42 6.752 17.928 ;
  LAYER M1 ;
        RECT 6.784 15.42 6.816 17.928 ;
  LAYER M1 ;
        RECT 6.848 15.42 6.88 17.928 ;
  LAYER M1 ;
        RECT 6.912 15.42 6.944 17.928 ;
  LAYER M1 ;
        RECT 6.976 15.42 7.008 17.928 ;
  LAYER M1 ;
        RECT 7.04 15.42 7.072 17.928 ;
  LAYER M1 ;
        RECT 7.104 15.42 7.136 17.928 ;
  LAYER M1 ;
        RECT 7.168 15.42 7.2 17.928 ;
  LAYER M1 ;
        RECT 7.232 15.42 7.264 17.928 ;
  LAYER M1 ;
        RECT 7.296 15.42 7.328 17.928 ;
  LAYER M1 ;
        RECT 7.36 15.42 7.392 17.928 ;
  LAYER M1 ;
        RECT 7.424 15.42 7.456 17.928 ;
  LAYER M1 ;
        RECT 7.488 15.42 7.52 17.928 ;
  LAYER M1 ;
        RECT 7.552 15.42 7.584 17.928 ;
  LAYER M1 ;
        RECT 7.616 15.42 7.648 17.928 ;
  LAYER M1 ;
        RECT 7.68 15.42 7.712 17.928 ;
  LAYER M1 ;
        RECT 7.744 15.42 7.776 17.928 ;
  LAYER M1 ;
        RECT 7.808 15.42 7.84 17.928 ;
  LAYER M1 ;
        RECT 7.872 15.42 7.904 17.928 ;
  LAYER M1 ;
        RECT 7.936 15.42 7.968 17.928 ;
  LAYER M1 ;
        RECT 8 15.42 8.032 17.928 ;
  LAYER M1 ;
        RECT 8.064 15.42 8.096 17.928 ;
  LAYER M1 ;
        RECT 8.128 15.42 8.16 17.928 ;
  LAYER M1 ;
        RECT 8.192 15.42 8.224 17.928 ;
  LAYER M1 ;
        RECT 8.256 15.42 8.288 17.928 ;
  LAYER M1 ;
        RECT 8.32 15.42 8.352 17.928 ;
  LAYER M1 ;
        RECT 8.384 15.42 8.416 17.928 ;
  LAYER M1 ;
        RECT 8.448 15.42 8.48 17.928 ;
  LAYER M2 ;
        RECT 6.124 15.504 8.596 15.536 ;
  LAYER M2 ;
        RECT 6.124 15.568 8.596 15.6 ;
  LAYER M2 ;
        RECT 6.124 15.632 8.596 15.664 ;
  LAYER M2 ;
        RECT 6.124 15.696 8.596 15.728 ;
  LAYER M2 ;
        RECT 6.124 15.76 8.596 15.792 ;
  LAYER M2 ;
        RECT 6.124 15.824 8.596 15.856 ;
  LAYER M2 ;
        RECT 6.124 15.888 8.596 15.92 ;
  LAYER M2 ;
        RECT 6.124 15.952 8.596 15.984 ;
  LAYER M2 ;
        RECT 6.124 16.016 8.596 16.048 ;
  LAYER M2 ;
        RECT 6.124 16.08 8.596 16.112 ;
  LAYER M2 ;
        RECT 6.124 16.144 8.596 16.176 ;
  LAYER M2 ;
        RECT 6.124 16.208 8.596 16.24 ;
  LAYER M2 ;
        RECT 6.124 16.272 8.596 16.304 ;
  LAYER M2 ;
        RECT 6.124 16.336 8.596 16.368 ;
  LAYER M2 ;
        RECT 6.124 16.4 8.596 16.432 ;
  LAYER M2 ;
        RECT 6.124 16.464 8.596 16.496 ;
  LAYER M2 ;
        RECT 6.124 16.528 8.596 16.56 ;
  LAYER M2 ;
        RECT 6.124 16.592 8.596 16.624 ;
  LAYER M2 ;
        RECT 6.124 16.656 8.596 16.688 ;
  LAYER M2 ;
        RECT 6.124 16.72 8.596 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.784 8.596 16.816 ;
  LAYER M2 ;
        RECT 6.124 16.848 8.596 16.88 ;
  LAYER M2 ;
        RECT 6.124 16.912 8.596 16.944 ;
  LAYER M2 ;
        RECT 6.124 16.976 8.596 17.008 ;
  LAYER M2 ;
        RECT 6.124 17.04 8.596 17.072 ;
  LAYER M2 ;
        RECT 6.124 17.104 8.596 17.136 ;
  LAYER M2 ;
        RECT 6.124 17.168 8.596 17.2 ;
  LAYER M2 ;
        RECT 6.124 17.232 8.596 17.264 ;
  LAYER M2 ;
        RECT 6.124 17.296 8.596 17.328 ;
  LAYER M2 ;
        RECT 6.124 17.36 8.596 17.392 ;
  LAYER M2 ;
        RECT 6.124 17.424 8.596 17.456 ;
  LAYER M2 ;
        RECT 6.124 17.488 8.596 17.52 ;
  LAYER M2 ;
        RECT 6.124 17.552 8.596 17.584 ;
  LAYER M2 ;
        RECT 6.124 17.616 8.596 17.648 ;
  LAYER M2 ;
        RECT 6.124 17.68 8.596 17.712 ;
  LAYER M2 ;
        RECT 6.124 17.744 8.596 17.776 ;
  LAYER M3 ;
        RECT 6.144 15.42 6.176 17.928 ;
  LAYER M3 ;
        RECT 6.208 15.42 6.24 17.928 ;
  LAYER M3 ;
        RECT 6.272 15.42 6.304 17.928 ;
  LAYER M3 ;
        RECT 6.336 15.42 6.368 17.928 ;
  LAYER M3 ;
        RECT 6.4 15.42 6.432 17.928 ;
  LAYER M3 ;
        RECT 6.464 15.42 6.496 17.928 ;
  LAYER M3 ;
        RECT 6.528 15.42 6.56 17.928 ;
  LAYER M3 ;
        RECT 6.592 15.42 6.624 17.928 ;
  LAYER M3 ;
        RECT 6.656 15.42 6.688 17.928 ;
  LAYER M3 ;
        RECT 6.72 15.42 6.752 17.928 ;
  LAYER M3 ;
        RECT 6.784 15.42 6.816 17.928 ;
  LAYER M3 ;
        RECT 6.848 15.42 6.88 17.928 ;
  LAYER M3 ;
        RECT 6.912 15.42 6.944 17.928 ;
  LAYER M3 ;
        RECT 6.976 15.42 7.008 17.928 ;
  LAYER M3 ;
        RECT 7.04 15.42 7.072 17.928 ;
  LAYER M3 ;
        RECT 7.104 15.42 7.136 17.928 ;
  LAYER M3 ;
        RECT 7.168 15.42 7.2 17.928 ;
  LAYER M3 ;
        RECT 7.232 15.42 7.264 17.928 ;
  LAYER M3 ;
        RECT 7.296 15.42 7.328 17.928 ;
  LAYER M3 ;
        RECT 7.36 15.42 7.392 17.928 ;
  LAYER M3 ;
        RECT 7.424 15.42 7.456 17.928 ;
  LAYER M3 ;
        RECT 7.488 15.42 7.52 17.928 ;
  LAYER M3 ;
        RECT 7.552 15.42 7.584 17.928 ;
  LAYER M3 ;
        RECT 7.616 15.42 7.648 17.928 ;
  LAYER M3 ;
        RECT 7.68 15.42 7.712 17.928 ;
  LAYER M3 ;
        RECT 7.744 15.42 7.776 17.928 ;
  LAYER M3 ;
        RECT 7.808 15.42 7.84 17.928 ;
  LAYER M3 ;
        RECT 7.872 15.42 7.904 17.928 ;
  LAYER M3 ;
        RECT 7.936 15.42 7.968 17.928 ;
  LAYER M3 ;
        RECT 8 15.42 8.032 17.928 ;
  LAYER M3 ;
        RECT 8.064 15.42 8.096 17.928 ;
  LAYER M3 ;
        RECT 8.128 15.42 8.16 17.928 ;
  LAYER M3 ;
        RECT 8.192 15.42 8.224 17.928 ;
  LAYER M3 ;
        RECT 8.256 15.42 8.288 17.928 ;
  LAYER M3 ;
        RECT 8.32 15.42 8.352 17.928 ;
  LAYER M3 ;
        RECT 8.384 15.42 8.416 17.928 ;
  LAYER M3 ;
        RECT 8.448 15.42 8.48 17.928 ;
  LAYER M3 ;
        RECT 8.544 15.42 8.576 17.928 ;
  LAYER M1 ;
        RECT 6.159 15.456 6.161 17.892 ;
  LAYER M1 ;
        RECT 6.239 15.456 6.241 17.892 ;
  LAYER M1 ;
        RECT 6.319 15.456 6.321 17.892 ;
  LAYER M1 ;
        RECT 6.399 15.456 6.401 17.892 ;
  LAYER M1 ;
        RECT 6.479 15.456 6.481 17.892 ;
  LAYER M1 ;
        RECT 6.559 15.456 6.561 17.892 ;
  LAYER M1 ;
        RECT 6.639 15.456 6.641 17.892 ;
  LAYER M1 ;
        RECT 6.719 15.456 6.721 17.892 ;
  LAYER M1 ;
        RECT 6.799 15.456 6.801 17.892 ;
  LAYER M1 ;
        RECT 6.879 15.456 6.881 17.892 ;
  LAYER M1 ;
        RECT 6.959 15.456 6.961 17.892 ;
  LAYER M1 ;
        RECT 7.039 15.456 7.041 17.892 ;
  LAYER M1 ;
        RECT 7.119 15.456 7.121 17.892 ;
  LAYER M1 ;
        RECT 7.199 15.456 7.201 17.892 ;
  LAYER M1 ;
        RECT 7.279 15.456 7.281 17.892 ;
  LAYER M1 ;
        RECT 7.359 15.456 7.361 17.892 ;
  LAYER M1 ;
        RECT 7.439 15.456 7.441 17.892 ;
  LAYER M1 ;
        RECT 7.519 15.456 7.521 17.892 ;
  LAYER M1 ;
        RECT 7.599 15.456 7.601 17.892 ;
  LAYER M1 ;
        RECT 7.679 15.456 7.681 17.892 ;
  LAYER M1 ;
        RECT 7.759 15.456 7.761 17.892 ;
  LAYER M1 ;
        RECT 7.839 15.456 7.841 17.892 ;
  LAYER M1 ;
        RECT 7.919 15.456 7.921 17.892 ;
  LAYER M1 ;
        RECT 7.999 15.456 8.001 17.892 ;
  LAYER M1 ;
        RECT 8.079 15.456 8.081 17.892 ;
  LAYER M1 ;
        RECT 8.159 15.456 8.161 17.892 ;
  LAYER M1 ;
        RECT 8.239 15.456 8.241 17.892 ;
  LAYER M1 ;
        RECT 8.319 15.456 8.321 17.892 ;
  LAYER M1 ;
        RECT 8.399 15.456 8.401 17.892 ;
  LAYER M1 ;
        RECT 8.479 15.456 8.481 17.892 ;
  LAYER M2 ;
        RECT 6.16 15.455 8.56 15.457 ;
  LAYER M2 ;
        RECT 6.16 15.539 8.56 15.541 ;
  LAYER M2 ;
        RECT 6.16 15.623 8.56 15.625 ;
  LAYER M2 ;
        RECT 6.16 15.707 8.56 15.709 ;
  LAYER M2 ;
        RECT 6.16 15.791 8.56 15.793 ;
  LAYER M2 ;
        RECT 6.16 15.875 8.56 15.877 ;
  LAYER M2 ;
        RECT 6.16 15.959 8.56 15.961 ;
  LAYER M2 ;
        RECT 6.16 16.043 8.56 16.045 ;
  LAYER M2 ;
        RECT 6.16 16.127 8.56 16.129 ;
  LAYER M2 ;
        RECT 6.16 16.211 8.56 16.213 ;
  LAYER M2 ;
        RECT 6.16 16.295 8.56 16.297 ;
  LAYER M2 ;
        RECT 6.16 16.379 8.56 16.381 ;
  LAYER M2 ;
        RECT 6.16 16.4625 8.56 16.4645 ;
  LAYER M2 ;
        RECT 6.16 16.547 8.56 16.549 ;
  LAYER M2 ;
        RECT 6.16 16.631 8.56 16.633 ;
  LAYER M2 ;
        RECT 6.16 16.715 8.56 16.717 ;
  LAYER M2 ;
        RECT 6.16 16.799 8.56 16.801 ;
  LAYER M2 ;
        RECT 6.16 16.883 8.56 16.885 ;
  LAYER M2 ;
        RECT 6.16 16.967 8.56 16.969 ;
  LAYER M2 ;
        RECT 6.16 17.051 8.56 17.053 ;
  LAYER M2 ;
        RECT 6.16 17.135 8.56 17.137 ;
  LAYER M2 ;
        RECT 6.16 17.219 8.56 17.221 ;
  LAYER M2 ;
        RECT 6.16 17.303 8.56 17.305 ;
  LAYER M2 ;
        RECT 6.16 17.387 8.56 17.389 ;
  LAYER M2 ;
        RECT 6.16 17.471 8.56 17.473 ;
  LAYER M2 ;
        RECT 6.16 17.555 8.56 17.557 ;
  LAYER M2 ;
        RECT 6.16 17.639 8.56 17.641 ;
  LAYER M2 ;
        RECT 6.16 17.723 8.56 17.725 ;
  LAYER M2 ;
        RECT 6.16 17.807 8.56 17.809 ;
  LAYER M1 ;
        RECT 9.024 0.72 9.056 3.228 ;
  LAYER M1 ;
        RECT 9.088 0.72 9.12 3.228 ;
  LAYER M1 ;
        RECT 9.152 0.72 9.184 3.228 ;
  LAYER M1 ;
        RECT 9.216 0.72 9.248 3.228 ;
  LAYER M1 ;
        RECT 9.28 0.72 9.312 3.228 ;
  LAYER M1 ;
        RECT 9.344 0.72 9.376 3.228 ;
  LAYER M1 ;
        RECT 9.408 0.72 9.44 3.228 ;
  LAYER M1 ;
        RECT 9.472 0.72 9.504 3.228 ;
  LAYER M1 ;
        RECT 9.536 0.72 9.568 3.228 ;
  LAYER M1 ;
        RECT 9.6 0.72 9.632 3.228 ;
  LAYER M1 ;
        RECT 9.664 0.72 9.696 3.228 ;
  LAYER M1 ;
        RECT 9.728 0.72 9.76 3.228 ;
  LAYER M1 ;
        RECT 9.792 0.72 9.824 3.228 ;
  LAYER M1 ;
        RECT 9.856 0.72 9.888 3.228 ;
  LAYER M1 ;
        RECT 9.92 0.72 9.952 3.228 ;
  LAYER M1 ;
        RECT 9.984 0.72 10.016 3.228 ;
  LAYER M1 ;
        RECT 10.048 0.72 10.08 3.228 ;
  LAYER M1 ;
        RECT 10.112 0.72 10.144 3.228 ;
  LAYER M1 ;
        RECT 10.176 0.72 10.208 3.228 ;
  LAYER M1 ;
        RECT 10.24 0.72 10.272 3.228 ;
  LAYER M1 ;
        RECT 10.304 0.72 10.336 3.228 ;
  LAYER M1 ;
        RECT 10.368 0.72 10.4 3.228 ;
  LAYER M1 ;
        RECT 10.432 0.72 10.464 3.228 ;
  LAYER M1 ;
        RECT 10.496 0.72 10.528 3.228 ;
  LAYER M1 ;
        RECT 10.56 0.72 10.592 3.228 ;
  LAYER M1 ;
        RECT 10.624 0.72 10.656 3.228 ;
  LAYER M1 ;
        RECT 10.688 0.72 10.72 3.228 ;
  LAYER M1 ;
        RECT 10.752 0.72 10.784 3.228 ;
  LAYER M1 ;
        RECT 10.816 0.72 10.848 3.228 ;
  LAYER M1 ;
        RECT 10.88 0.72 10.912 3.228 ;
  LAYER M1 ;
        RECT 10.944 0.72 10.976 3.228 ;
  LAYER M1 ;
        RECT 11.008 0.72 11.04 3.228 ;
  LAYER M1 ;
        RECT 11.072 0.72 11.104 3.228 ;
  LAYER M1 ;
        RECT 11.136 0.72 11.168 3.228 ;
  LAYER M1 ;
        RECT 11.2 0.72 11.232 3.228 ;
  LAYER M1 ;
        RECT 11.264 0.72 11.296 3.228 ;
  LAYER M1 ;
        RECT 11.328 0.72 11.36 3.228 ;
  LAYER M2 ;
        RECT 9.004 0.804 11.476 0.836 ;
  LAYER M2 ;
        RECT 9.004 0.868 11.476 0.9 ;
  LAYER M2 ;
        RECT 9.004 0.932 11.476 0.964 ;
  LAYER M2 ;
        RECT 9.004 0.996 11.476 1.028 ;
  LAYER M2 ;
        RECT 9.004 1.06 11.476 1.092 ;
  LAYER M2 ;
        RECT 9.004 1.124 11.476 1.156 ;
  LAYER M2 ;
        RECT 9.004 1.188 11.476 1.22 ;
  LAYER M2 ;
        RECT 9.004 1.252 11.476 1.284 ;
  LAYER M2 ;
        RECT 9.004 1.316 11.476 1.348 ;
  LAYER M2 ;
        RECT 9.004 1.38 11.476 1.412 ;
  LAYER M2 ;
        RECT 9.004 1.444 11.476 1.476 ;
  LAYER M2 ;
        RECT 9.004 1.508 11.476 1.54 ;
  LAYER M2 ;
        RECT 9.004 1.572 11.476 1.604 ;
  LAYER M2 ;
        RECT 9.004 1.636 11.476 1.668 ;
  LAYER M2 ;
        RECT 9.004 1.7 11.476 1.732 ;
  LAYER M2 ;
        RECT 9.004 1.764 11.476 1.796 ;
  LAYER M2 ;
        RECT 9.004 1.828 11.476 1.86 ;
  LAYER M2 ;
        RECT 9.004 1.892 11.476 1.924 ;
  LAYER M2 ;
        RECT 9.004 1.956 11.476 1.988 ;
  LAYER M2 ;
        RECT 9.004 2.02 11.476 2.052 ;
  LAYER M2 ;
        RECT 9.004 2.084 11.476 2.116 ;
  LAYER M2 ;
        RECT 9.004 2.148 11.476 2.18 ;
  LAYER M2 ;
        RECT 9.004 2.212 11.476 2.244 ;
  LAYER M2 ;
        RECT 9.004 2.276 11.476 2.308 ;
  LAYER M2 ;
        RECT 9.004 2.34 11.476 2.372 ;
  LAYER M2 ;
        RECT 9.004 2.404 11.476 2.436 ;
  LAYER M2 ;
        RECT 9.004 2.468 11.476 2.5 ;
  LAYER M2 ;
        RECT 9.004 2.532 11.476 2.564 ;
  LAYER M2 ;
        RECT 9.004 2.596 11.476 2.628 ;
  LAYER M2 ;
        RECT 9.004 2.66 11.476 2.692 ;
  LAYER M2 ;
        RECT 9.004 2.724 11.476 2.756 ;
  LAYER M2 ;
        RECT 9.004 2.788 11.476 2.82 ;
  LAYER M2 ;
        RECT 9.004 2.852 11.476 2.884 ;
  LAYER M2 ;
        RECT 9.004 2.916 11.476 2.948 ;
  LAYER M2 ;
        RECT 9.004 2.98 11.476 3.012 ;
  LAYER M2 ;
        RECT 9.004 3.044 11.476 3.076 ;
  LAYER M3 ;
        RECT 9.024 0.72 9.056 3.228 ;
  LAYER M3 ;
        RECT 9.088 0.72 9.12 3.228 ;
  LAYER M3 ;
        RECT 9.152 0.72 9.184 3.228 ;
  LAYER M3 ;
        RECT 9.216 0.72 9.248 3.228 ;
  LAYER M3 ;
        RECT 9.28 0.72 9.312 3.228 ;
  LAYER M3 ;
        RECT 9.344 0.72 9.376 3.228 ;
  LAYER M3 ;
        RECT 9.408 0.72 9.44 3.228 ;
  LAYER M3 ;
        RECT 9.472 0.72 9.504 3.228 ;
  LAYER M3 ;
        RECT 9.536 0.72 9.568 3.228 ;
  LAYER M3 ;
        RECT 9.6 0.72 9.632 3.228 ;
  LAYER M3 ;
        RECT 9.664 0.72 9.696 3.228 ;
  LAYER M3 ;
        RECT 9.728 0.72 9.76 3.228 ;
  LAYER M3 ;
        RECT 9.792 0.72 9.824 3.228 ;
  LAYER M3 ;
        RECT 9.856 0.72 9.888 3.228 ;
  LAYER M3 ;
        RECT 9.92 0.72 9.952 3.228 ;
  LAYER M3 ;
        RECT 9.984 0.72 10.016 3.228 ;
  LAYER M3 ;
        RECT 10.048 0.72 10.08 3.228 ;
  LAYER M3 ;
        RECT 10.112 0.72 10.144 3.228 ;
  LAYER M3 ;
        RECT 10.176 0.72 10.208 3.228 ;
  LAYER M3 ;
        RECT 10.24 0.72 10.272 3.228 ;
  LAYER M3 ;
        RECT 10.304 0.72 10.336 3.228 ;
  LAYER M3 ;
        RECT 10.368 0.72 10.4 3.228 ;
  LAYER M3 ;
        RECT 10.432 0.72 10.464 3.228 ;
  LAYER M3 ;
        RECT 10.496 0.72 10.528 3.228 ;
  LAYER M3 ;
        RECT 10.56 0.72 10.592 3.228 ;
  LAYER M3 ;
        RECT 10.624 0.72 10.656 3.228 ;
  LAYER M3 ;
        RECT 10.688 0.72 10.72 3.228 ;
  LAYER M3 ;
        RECT 10.752 0.72 10.784 3.228 ;
  LAYER M3 ;
        RECT 10.816 0.72 10.848 3.228 ;
  LAYER M3 ;
        RECT 10.88 0.72 10.912 3.228 ;
  LAYER M3 ;
        RECT 10.944 0.72 10.976 3.228 ;
  LAYER M3 ;
        RECT 11.008 0.72 11.04 3.228 ;
  LAYER M3 ;
        RECT 11.072 0.72 11.104 3.228 ;
  LAYER M3 ;
        RECT 11.136 0.72 11.168 3.228 ;
  LAYER M3 ;
        RECT 11.2 0.72 11.232 3.228 ;
  LAYER M3 ;
        RECT 11.264 0.72 11.296 3.228 ;
  LAYER M3 ;
        RECT 11.328 0.72 11.36 3.228 ;
  LAYER M3 ;
        RECT 11.424 0.72 11.456 3.228 ;
  LAYER M1 ;
        RECT 9.039 0.756 9.041 3.192 ;
  LAYER M1 ;
        RECT 9.119 0.756 9.121 3.192 ;
  LAYER M1 ;
        RECT 9.199 0.756 9.201 3.192 ;
  LAYER M1 ;
        RECT 9.279 0.756 9.281 3.192 ;
  LAYER M1 ;
        RECT 9.359 0.756 9.361 3.192 ;
  LAYER M1 ;
        RECT 9.439 0.756 9.441 3.192 ;
  LAYER M1 ;
        RECT 9.519 0.756 9.521 3.192 ;
  LAYER M1 ;
        RECT 9.599 0.756 9.601 3.192 ;
  LAYER M1 ;
        RECT 9.679 0.756 9.681 3.192 ;
  LAYER M1 ;
        RECT 9.759 0.756 9.761 3.192 ;
  LAYER M1 ;
        RECT 9.839 0.756 9.841 3.192 ;
  LAYER M1 ;
        RECT 9.919 0.756 9.921 3.192 ;
  LAYER M1 ;
        RECT 9.999 0.756 10.001 3.192 ;
  LAYER M1 ;
        RECT 10.079 0.756 10.081 3.192 ;
  LAYER M1 ;
        RECT 10.159 0.756 10.161 3.192 ;
  LAYER M1 ;
        RECT 10.239 0.756 10.241 3.192 ;
  LAYER M1 ;
        RECT 10.319 0.756 10.321 3.192 ;
  LAYER M1 ;
        RECT 10.399 0.756 10.401 3.192 ;
  LAYER M1 ;
        RECT 10.479 0.756 10.481 3.192 ;
  LAYER M1 ;
        RECT 10.559 0.756 10.561 3.192 ;
  LAYER M1 ;
        RECT 10.639 0.756 10.641 3.192 ;
  LAYER M1 ;
        RECT 10.719 0.756 10.721 3.192 ;
  LAYER M1 ;
        RECT 10.799 0.756 10.801 3.192 ;
  LAYER M1 ;
        RECT 10.879 0.756 10.881 3.192 ;
  LAYER M1 ;
        RECT 10.959 0.756 10.961 3.192 ;
  LAYER M1 ;
        RECT 11.039 0.756 11.041 3.192 ;
  LAYER M1 ;
        RECT 11.119 0.756 11.121 3.192 ;
  LAYER M1 ;
        RECT 11.199 0.756 11.201 3.192 ;
  LAYER M1 ;
        RECT 11.279 0.756 11.281 3.192 ;
  LAYER M1 ;
        RECT 11.359 0.756 11.361 3.192 ;
  LAYER M2 ;
        RECT 9.04 0.755 11.44 0.757 ;
  LAYER M2 ;
        RECT 9.04 0.839 11.44 0.841 ;
  LAYER M2 ;
        RECT 9.04 0.923 11.44 0.925 ;
  LAYER M2 ;
        RECT 9.04 1.007 11.44 1.009 ;
  LAYER M2 ;
        RECT 9.04 1.091 11.44 1.093 ;
  LAYER M2 ;
        RECT 9.04 1.175 11.44 1.177 ;
  LAYER M2 ;
        RECT 9.04 1.259 11.44 1.261 ;
  LAYER M2 ;
        RECT 9.04 1.343 11.44 1.345 ;
  LAYER M2 ;
        RECT 9.04 1.427 11.44 1.429 ;
  LAYER M2 ;
        RECT 9.04 1.511 11.44 1.513 ;
  LAYER M2 ;
        RECT 9.04 1.595 11.44 1.597 ;
  LAYER M2 ;
        RECT 9.04 1.679 11.44 1.681 ;
  LAYER M2 ;
        RECT 9.04 1.7625 11.44 1.7645 ;
  LAYER M2 ;
        RECT 9.04 1.847 11.44 1.849 ;
  LAYER M2 ;
        RECT 9.04 1.931 11.44 1.933 ;
  LAYER M2 ;
        RECT 9.04 2.015 11.44 2.017 ;
  LAYER M2 ;
        RECT 9.04 2.099 11.44 2.101 ;
  LAYER M2 ;
        RECT 9.04 2.183 11.44 2.185 ;
  LAYER M2 ;
        RECT 9.04 2.267 11.44 2.269 ;
  LAYER M2 ;
        RECT 9.04 2.351 11.44 2.353 ;
  LAYER M2 ;
        RECT 9.04 2.435 11.44 2.437 ;
  LAYER M2 ;
        RECT 9.04 2.519 11.44 2.521 ;
  LAYER M2 ;
        RECT 9.04 2.603 11.44 2.605 ;
  LAYER M2 ;
        RECT 9.04 2.687 11.44 2.689 ;
  LAYER M2 ;
        RECT 9.04 2.771 11.44 2.773 ;
  LAYER M2 ;
        RECT 9.04 2.855 11.44 2.857 ;
  LAYER M2 ;
        RECT 9.04 2.939 11.44 2.941 ;
  LAYER M2 ;
        RECT 9.04 3.023 11.44 3.025 ;
  LAYER M2 ;
        RECT 9.04 3.107 11.44 3.109 ;
  LAYER M1 ;
        RECT 9.024 3.66 9.056 6.168 ;
  LAYER M1 ;
        RECT 9.088 3.66 9.12 6.168 ;
  LAYER M1 ;
        RECT 9.152 3.66 9.184 6.168 ;
  LAYER M1 ;
        RECT 9.216 3.66 9.248 6.168 ;
  LAYER M1 ;
        RECT 9.28 3.66 9.312 6.168 ;
  LAYER M1 ;
        RECT 9.344 3.66 9.376 6.168 ;
  LAYER M1 ;
        RECT 9.408 3.66 9.44 6.168 ;
  LAYER M1 ;
        RECT 9.472 3.66 9.504 6.168 ;
  LAYER M1 ;
        RECT 9.536 3.66 9.568 6.168 ;
  LAYER M1 ;
        RECT 9.6 3.66 9.632 6.168 ;
  LAYER M1 ;
        RECT 9.664 3.66 9.696 6.168 ;
  LAYER M1 ;
        RECT 9.728 3.66 9.76 6.168 ;
  LAYER M1 ;
        RECT 9.792 3.66 9.824 6.168 ;
  LAYER M1 ;
        RECT 9.856 3.66 9.888 6.168 ;
  LAYER M1 ;
        RECT 9.92 3.66 9.952 6.168 ;
  LAYER M1 ;
        RECT 9.984 3.66 10.016 6.168 ;
  LAYER M1 ;
        RECT 10.048 3.66 10.08 6.168 ;
  LAYER M1 ;
        RECT 10.112 3.66 10.144 6.168 ;
  LAYER M1 ;
        RECT 10.176 3.66 10.208 6.168 ;
  LAYER M1 ;
        RECT 10.24 3.66 10.272 6.168 ;
  LAYER M1 ;
        RECT 10.304 3.66 10.336 6.168 ;
  LAYER M1 ;
        RECT 10.368 3.66 10.4 6.168 ;
  LAYER M1 ;
        RECT 10.432 3.66 10.464 6.168 ;
  LAYER M1 ;
        RECT 10.496 3.66 10.528 6.168 ;
  LAYER M1 ;
        RECT 10.56 3.66 10.592 6.168 ;
  LAYER M1 ;
        RECT 10.624 3.66 10.656 6.168 ;
  LAYER M1 ;
        RECT 10.688 3.66 10.72 6.168 ;
  LAYER M1 ;
        RECT 10.752 3.66 10.784 6.168 ;
  LAYER M1 ;
        RECT 10.816 3.66 10.848 6.168 ;
  LAYER M1 ;
        RECT 10.88 3.66 10.912 6.168 ;
  LAYER M1 ;
        RECT 10.944 3.66 10.976 6.168 ;
  LAYER M1 ;
        RECT 11.008 3.66 11.04 6.168 ;
  LAYER M1 ;
        RECT 11.072 3.66 11.104 6.168 ;
  LAYER M1 ;
        RECT 11.136 3.66 11.168 6.168 ;
  LAYER M1 ;
        RECT 11.2 3.66 11.232 6.168 ;
  LAYER M1 ;
        RECT 11.264 3.66 11.296 6.168 ;
  LAYER M1 ;
        RECT 11.328 3.66 11.36 6.168 ;
  LAYER M2 ;
        RECT 9.004 3.744 11.476 3.776 ;
  LAYER M2 ;
        RECT 9.004 3.808 11.476 3.84 ;
  LAYER M2 ;
        RECT 9.004 3.872 11.476 3.904 ;
  LAYER M2 ;
        RECT 9.004 3.936 11.476 3.968 ;
  LAYER M2 ;
        RECT 9.004 4 11.476 4.032 ;
  LAYER M2 ;
        RECT 9.004 4.064 11.476 4.096 ;
  LAYER M2 ;
        RECT 9.004 4.128 11.476 4.16 ;
  LAYER M2 ;
        RECT 9.004 4.192 11.476 4.224 ;
  LAYER M2 ;
        RECT 9.004 4.256 11.476 4.288 ;
  LAYER M2 ;
        RECT 9.004 4.32 11.476 4.352 ;
  LAYER M2 ;
        RECT 9.004 4.384 11.476 4.416 ;
  LAYER M2 ;
        RECT 9.004 4.448 11.476 4.48 ;
  LAYER M2 ;
        RECT 9.004 4.512 11.476 4.544 ;
  LAYER M2 ;
        RECT 9.004 4.576 11.476 4.608 ;
  LAYER M2 ;
        RECT 9.004 4.64 11.476 4.672 ;
  LAYER M2 ;
        RECT 9.004 4.704 11.476 4.736 ;
  LAYER M2 ;
        RECT 9.004 4.768 11.476 4.8 ;
  LAYER M2 ;
        RECT 9.004 4.832 11.476 4.864 ;
  LAYER M2 ;
        RECT 9.004 4.896 11.476 4.928 ;
  LAYER M2 ;
        RECT 9.004 4.96 11.476 4.992 ;
  LAYER M2 ;
        RECT 9.004 5.024 11.476 5.056 ;
  LAYER M2 ;
        RECT 9.004 5.088 11.476 5.12 ;
  LAYER M2 ;
        RECT 9.004 5.152 11.476 5.184 ;
  LAYER M2 ;
        RECT 9.004 5.216 11.476 5.248 ;
  LAYER M2 ;
        RECT 9.004 5.28 11.476 5.312 ;
  LAYER M2 ;
        RECT 9.004 5.344 11.476 5.376 ;
  LAYER M2 ;
        RECT 9.004 5.408 11.476 5.44 ;
  LAYER M2 ;
        RECT 9.004 5.472 11.476 5.504 ;
  LAYER M2 ;
        RECT 9.004 5.536 11.476 5.568 ;
  LAYER M2 ;
        RECT 9.004 5.6 11.476 5.632 ;
  LAYER M2 ;
        RECT 9.004 5.664 11.476 5.696 ;
  LAYER M2 ;
        RECT 9.004 5.728 11.476 5.76 ;
  LAYER M2 ;
        RECT 9.004 5.792 11.476 5.824 ;
  LAYER M2 ;
        RECT 9.004 5.856 11.476 5.888 ;
  LAYER M2 ;
        RECT 9.004 5.92 11.476 5.952 ;
  LAYER M2 ;
        RECT 9.004 5.984 11.476 6.016 ;
  LAYER M3 ;
        RECT 9.024 3.66 9.056 6.168 ;
  LAYER M3 ;
        RECT 9.088 3.66 9.12 6.168 ;
  LAYER M3 ;
        RECT 9.152 3.66 9.184 6.168 ;
  LAYER M3 ;
        RECT 9.216 3.66 9.248 6.168 ;
  LAYER M3 ;
        RECT 9.28 3.66 9.312 6.168 ;
  LAYER M3 ;
        RECT 9.344 3.66 9.376 6.168 ;
  LAYER M3 ;
        RECT 9.408 3.66 9.44 6.168 ;
  LAYER M3 ;
        RECT 9.472 3.66 9.504 6.168 ;
  LAYER M3 ;
        RECT 9.536 3.66 9.568 6.168 ;
  LAYER M3 ;
        RECT 9.6 3.66 9.632 6.168 ;
  LAYER M3 ;
        RECT 9.664 3.66 9.696 6.168 ;
  LAYER M3 ;
        RECT 9.728 3.66 9.76 6.168 ;
  LAYER M3 ;
        RECT 9.792 3.66 9.824 6.168 ;
  LAYER M3 ;
        RECT 9.856 3.66 9.888 6.168 ;
  LAYER M3 ;
        RECT 9.92 3.66 9.952 6.168 ;
  LAYER M3 ;
        RECT 9.984 3.66 10.016 6.168 ;
  LAYER M3 ;
        RECT 10.048 3.66 10.08 6.168 ;
  LAYER M3 ;
        RECT 10.112 3.66 10.144 6.168 ;
  LAYER M3 ;
        RECT 10.176 3.66 10.208 6.168 ;
  LAYER M3 ;
        RECT 10.24 3.66 10.272 6.168 ;
  LAYER M3 ;
        RECT 10.304 3.66 10.336 6.168 ;
  LAYER M3 ;
        RECT 10.368 3.66 10.4 6.168 ;
  LAYER M3 ;
        RECT 10.432 3.66 10.464 6.168 ;
  LAYER M3 ;
        RECT 10.496 3.66 10.528 6.168 ;
  LAYER M3 ;
        RECT 10.56 3.66 10.592 6.168 ;
  LAYER M3 ;
        RECT 10.624 3.66 10.656 6.168 ;
  LAYER M3 ;
        RECT 10.688 3.66 10.72 6.168 ;
  LAYER M3 ;
        RECT 10.752 3.66 10.784 6.168 ;
  LAYER M3 ;
        RECT 10.816 3.66 10.848 6.168 ;
  LAYER M3 ;
        RECT 10.88 3.66 10.912 6.168 ;
  LAYER M3 ;
        RECT 10.944 3.66 10.976 6.168 ;
  LAYER M3 ;
        RECT 11.008 3.66 11.04 6.168 ;
  LAYER M3 ;
        RECT 11.072 3.66 11.104 6.168 ;
  LAYER M3 ;
        RECT 11.136 3.66 11.168 6.168 ;
  LAYER M3 ;
        RECT 11.2 3.66 11.232 6.168 ;
  LAYER M3 ;
        RECT 11.264 3.66 11.296 6.168 ;
  LAYER M3 ;
        RECT 11.328 3.66 11.36 6.168 ;
  LAYER M3 ;
        RECT 11.424 3.66 11.456 6.168 ;
  LAYER M1 ;
        RECT 9.039 3.696 9.041 6.132 ;
  LAYER M1 ;
        RECT 9.119 3.696 9.121 6.132 ;
  LAYER M1 ;
        RECT 9.199 3.696 9.201 6.132 ;
  LAYER M1 ;
        RECT 9.279 3.696 9.281 6.132 ;
  LAYER M1 ;
        RECT 9.359 3.696 9.361 6.132 ;
  LAYER M1 ;
        RECT 9.439 3.696 9.441 6.132 ;
  LAYER M1 ;
        RECT 9.519 3.696 9.521 6.132 ;
  LAYER M1 ;
        RECT 9.599 3.696 9.601 6.132 ;
  LAYER M1 ;
        RECT 9.679 3.696 9.681 6.132 ;
  LAYER M1 ;
        RECT 9.759 3.696 9.761 6.132 ;
  LAYER M1 ;
        RECT 9.839 3.696 9.841 6.132 ;
  LAYER M1 ;
        RECT 9.919 3.696 9.921 6.132 ;
  LAYER M1 ;
        RECT 9.999 3.696 10.001 6.132 ;
  LAYER M1 ;
        RECT 10.079 3.696 10.081 6.132 ;
  LAYER M1 ;
        RECT 10.159 3.696 10.161 6.132 ;
  LAYER M1 ;
        RECT 10.239 3.696 10.241 6.132 ;
  LAYER M1 ;
        RECT 10.319 3.696 10.321 6.132 ;
  LAYER M1 ;
        RECT 10.399 3.696 10.401 6.132 ;
  LAYER M1 ;
        RECT 10.479 3.696 10.481 6.132 ;
  LAYER M1 ;
        RECT 10.559 3.696 10.561 6.132 ;
  LAYER M1 ;
        RECT 10.639 3.696 10.641 6.132 ;
  LAYER M1 ;
        RECT 10.719 3.696 10.721 6.132 ;
  LAYER M1 ;
        RECT 10.799 3.696 10.801 6.132 ;
  LAYER M1 ;
        RECT 10.879 3.696 10.881 6.132 ;
  LAYER M1 ;
        RECT 10.959 3.696 10.961 6.132 ;
  LAYER M1 ;
        RECT 11.039 3.696 11.041 6.132 ;
  LAYER M1 ;
        RECT 11.119 3.696 11.121 6.132 ;
  LAYER M1 ;
        RECT 11.199 3.696 11.201 6.132 ;
  LAYER M1 ;
        RECT 11.279 3.696 11.281 6.132 ;
  LAYER M1 ;
        RECT 11.359 3.696 11.361 6.132 ;
  LAYER M2 ;
        RECT 9.04 3.695 11.44 3.697 ;
  LAYER M2 ;
        RECT 9.04 3.779 11.44 3.781 ;
  LAYER M2 ;
        RECT 9.04 3.863 11.44 3.865 ;
  LAYER M2 ;
        RECT 9.04 3.947 11.44 3.949 ;
  LAYER M2 ;
        RECT 9.04 4.031 11.44 4.033 ;
  LAYER M2 ;
        RECT 9.04 4.115 11.44 4.117 ;
  LAYER M2 ;
        RECT 9.04 4.199 11.44 4.201 ;
  LAYER M2 ;
        RECT 9.04 4.283 11.44 4.285 ;
  LAYER M2 ;
        RECT 9.04 4.367 11.44 4.369 ;
  LAYER M2 ;
        RECT 9.04 4.451 11.44 4.453 ;
  LAYER M2 ;
        RECT 9.04 4.535 11.44 4.537 ;
  LAYER M2 ;
        RECT 9.04 4.619 11.44 4.621 ;
  LAYER M2 ;
        RECT 9.04 4.7025 11.44 4.7045 ;
  LAYER M2 ;
        RECT 9.04 4.787 11.44 4.789 ;
  LAYER M2 ;
        RECT 9.04 4.871 11.44 4.873 ;
  LAYER M2 ;
        RECT 9.04 4.955 11.44 4.957 ;
  LAYER M2 ;
        RECT 9.04 5.039 11.44 5.041 ;
  LAYER M2 ;
        RECT 9.04 5.123 11.44 5.125 ;
  LAYER M2 ;
        RECT 9.04 5.207 11.44 5.209 ;
  LAYER M2 ;
        RECT 9.04 5.291 11.44 5.293 ;
  LAYER M2 ;
        RECT 9.04 5.375 11.44 5.377 ;
  LAYER M2 ;
        RECT 9.04 5.459 11.44 5.461 ;
  LAYER M2 ;
        RECT 9.04 5.543 11.44 5.545 ;
  LAYER M2 ;
        RECT 9.04 5.627 11.44 5.629 ;
  LAYER M2 ;
        RECT 9.04 5.711 11.44 5.713 ;
  LAYER M2 ;
        RECT 9.04 5.795 11.44 5.797 ;
  LAYER M2 ;
        RECT 9.04 5.879 11.44 5.881 ;
  LAYER M2 ;
        RECT 9.04 5.963 11.44 5.965 ;
  LAYER M2 ;
        RECT 9.04 6.047 11.44 6.049 ;
  LAYER M1 ;
        RECT 9.024 6.6 9.056 9.108 ;
  LAYER M1 ;
        RECT 9.088 6.6 9.12 9.108 ;
  LAYER M1 ;
        RECT 9.152 6.6 9.184 9.108 ;
  LAYER M1 ;
        RECT 9.216 6.6 9.248 9.108 ;
  LAYER M1 ;
        RECT 9.28 6.6 9.312 9.108 ;
  LAYER M1 ;
        RECT 9.344 6.6 9.376 9.108 ;
  LAYER M1 ;
        RECT 9.408 6.6 9.44 9.108 ;
  LAYER M1 ;
        RECT 9.472 6.6 9.504 9.108 ;
  LAYER M1 ;
        RECT 9.536 6.6 9.568 9.108 ;
  LAYER M1 ;
        RECT 9.6 6.6 9.632 9.108 ;
  LAYER M1 ;
        RECT 9.664 6.6 9.696 9.108 ;
  LAYER M1 ;
        RECT 9.728 6.6 9.76 9.108 ;
  LAYER M1 ;
        RECT 9.792 6.6 9.824 9.108 ;
  LAYER M1 ;
        RECT 9.856 6.6 9.888 9.108 ;
  LAYER M1 ;
        RECT 9.92 6.6 9.952 9.108 ;
  LAYER M1 ;
        RECT 9.984 6.6 10.016 9.108 ;
  LAYER M1 ;
        RECT 10.048 6.6 10.08 9.108 ;
  LAYER M1 ;
        RECT 10.112 6.6 10.144 9.108 ;
  LAYER M1 ;
        RECT 10.176 6.6 10.208 9.108 ;
  LAYER M1 ;
        RECT 10.24 6.6 10.272 9.108 ;
  LAYER M1 ;
        RECT 10.304 6.6 10.336 9.108 ;
  LAYER M1 ;
        RECT 10.368 6.6 10.4 9.108 ;
  LAYER M1 ;
        RECT 10.432 6.6 10.464 9.108 ;
  LAYER M1 ;
        RECT 10.496 6.6 10.528 9.108 ;
  LAYER M1 ;
        RECT 10.56 6.6 10.592 9.108 ;
  LAYER M1 ;
        RECT 10.624 6.6 10.656 9.108 ;
  LAYER M1 ;
        RECT 10.688 6.6 10.72 9.108 ;
  LAYER M1 ;
        RECT 10.752 6.6 10.784 9.108 ;
  LAYER M1 ;
        RECT 10.816 6.6 10.848 9.108 ;
  LAYER M1 ;
        RECT 10.88 6.6 10.912 9.108 ;
  LAYER M1 ;
        RECT 10.944 6.6 10.976 9.108 ;
  LAYER M1 ;
        RECT 11.008 6.6 11.04 9.108 ;
  LAYER M1 ;
        RECT 11.072 6.6 11.104 9.108 ;
  LAYER M1 ;
        RECT 11.136 6.6 11.168 9.108 ;
  LAYER M1 ;
        RECT 11.2 6.6 11.232 9.108 ;
  LAYER M1 ;
        RECT 11.264 6.6 11.296 9.108 ;
  LAYER M1 ;
        RECT 11.328 6.6 11.36 9.108 ;
  LAYER M2 ;
        RECT 9.004 6.684 11.476 6.716 ;
  LAYER M2 ;
        RECT 9.004 6.748 11.476 6.78 ;
  LAYER M2 ;
        RECT 9.004 6.812 11.476 6.844 ;
  LAYER M2 ;
        RECT 9.004 6.876 11.476 6.908 ;
  LAYER M2 ;
        RECT 9.004 6.94 11.476 6.972 ;
  LAYER M2 ;
        RECT 9.004 7.004 11.476 7.036 ;
  LAYER M2 ;
        RECT 9.004 7.068 11.476 7.1 ;
  LAYER M2 ;
        RECT 9.004 7.132 11.476 7.164 ;
  LAYER M2 ;
        RECT 9.004 7.196 11.476 7.228 ;
  LAYER M2 ;
        RECT 9.004 7.26 11.476 7.292 ;
  LAYER M2 ;
        RECT 9.004 7.324 11.476 7.356 ;
  LAYER M2 ;
        RECT 9.004 7.388 11.476 7.42 ;
  LAYER M2 ;
        RECT 9.004 7.452 11.476 7.484 ;
  LAYER M2 ;
        RECT 9.004 7.516 11.476 7.548 ;
  LAYER M2 ;
        RECT 9.004 7.58 11.476 7.612 ;
  LAYER M2 ;
        RECT 9.004 7.644 11.476 7.676 ;
  LAYER M2 ;
        RECT 9.004 7.708 11.476 7.74 ;
  LAYER M2 ;
        RECT 9.004 7.772 11.476 7.804 ;
  LAYER M2 ;
        RECT 9.004 7.836 11.476 7.868 ;
  LAYER M2 ;
        RECT 9.004 7.9 11.476 7.932 ;
  LAYER M2 ;
        RECT 9.004 7.964 11.476 7.996 ;
  LAYER M2 ;
        RECT 9.004 8.028 11.476 8.06 ;
  LAYER M2 ;
        RECT 9.004 8.092 11.476 8.124 ;
  LAYER M2 ;
        RECT 9.004 8.156 11.476 8.188 ;
  LAYER M2 ;
        RECT 9.004 8.22 11.476 8.252 ;
  LAYER M2 ;
        RECT 9.004 8.284 11.476 8.316 ;
  LAYER M2 ;
        RECT 9.004 8.348 11.476 8.38 ;
  LAYER M2 ;
        RECT 9.004 8.412 11.476 8.444 ;
  LAYER M2 ;
        RECT 9.004 8.476 11.476 8.508 ;
  LAYER M2 ;
        RECT 9.004 8.54 11.476 8.572 ;
  LAYER M2 ;
        RECT 9.004 8.604 11.476 8.636 ;
  LAYER M2 ;
        RECT 9.004 8.668 11.476 8.7 ;
  LAYER M2 ;
        RECT 9.004 8.732 11.476 8.764 ;
  LAYER M2 ;
        RECT 9.004 8.796 11.476 8.828 ;
  LAYER M2 ;
        RECT 9.004 8.86 11.476 8.892 ;
  LAYER M2 ;
        RECT 9.004 8.924 11.476 8.956 ;
  LAYER M3 ;
        RECT 9.024 6.6 9.056 9.108 ;
  LAYER M3 ;
        RECT 9.088 6.6 9.12 9.108 ;
  LAYER M3 ;
        RECT 9.152 6.6 9.184 9.108 ;
  LAYER M3 ;
        RECT 9.216 6.6 9.248 9.108 ;
  LAYER M3 ;
        RECT 9.28 6.6 9.312 9.108 ;
  LAYER M3 ;
        RECT 9.344 6.6 9.376 9.108 ;
  LAYER M3 ;
        RECT 9.408 6.6 9.44 9.108 ;
  LAYER M3 ;
        RECT 9.472 6.6 9.504 9.108 ;
  LAYER M3 ;
        RECT 9.536 6.6 9.568 9.108 ;
  LAYER M3 ;
        RECT 9.6 6.6 9.632 9.108 ;
  LAYER M3 ;
        RECT 9.664 6.6 9.696 9.108 ;
  LAYER M3 ;
        RECT 9.728 6.6 9.76 9.108 ;
  LAYER M3 ;
        RECT 9.792 6.6 9.824 9.108 ;
  LAYER M3 ;
        RECT 9.856 6.6 9.888 9.108 ;
  LAYER M3 ;
        RECT 9.92 6.6 9.952 9.108 ;
  LAYER M3 ;
        RECT 9.984 6.6 10.016 9.108 ;
  LAYER M3 ;
        RECT 10.048 6.6 10.08 9.108 ;
  LAYER M3 ;
        RECT 10.112 6.6 10.144 9.108 ;
  LAYER M3 ;
        RECT 10.176 6.6 10.208 9.108 ;
  LAYER M3 ;
        RECT 10.24 6.6 10.272 9.108 ;
  LAYER M3 ;
        RECT 10.304 6.6 10.336 9.108 ;
  LAYER M3 ;
        RECT 10.368 6.6 10.4 9.108 ;
  LAYER M3 ;
        RECT 10.432 6.6 10.464 9.108 ;
  LAYER M3 ;
        RECT 10.496 6.6 10.528 9.108 ;
  LAYER M3 ;
        RECT 10.56 6.6 10.592 9.108 ;
  LAYER M3 ;
        RECT 10.624 6.6 10.656 9.108 ;
  LAYER M3 ;
        RECT 10.688 6.6 10.72 9.108 ;
  LAYER M3 ;
        RECT 10.752 6.6 10.784 9.108 ;
  LAYER M3 ;
        RECT 10.816 6.6 10.848 9.108 ;
  LAYER M3 ;
        RECT 10.88 6.6 10.912 9.108 ;
  LAYER M3 ;
        RECT 10.944 6.6 10.976 9.108 ;
  LAYER M3 ;
        RECT 11.008 6.6 11.04 9.108 ;
  LAYER M3 ;
        RECT 11.072 6.6 11.104 9.108 ;
  LAYER M3 ;
        RECT 11.136 6.6 11.168 9.108 ;
  LAYER M3 ;
        RECT 11.2 6.6 11.232 9.108 ;
  LAYER M3 ;
        RECT 11.264 6.6 11.296 9.108 ;
  LAYER M3 ;
        RECT 11.328 6.6 11.36 9.108 ;
  LAYER M3 ;
        RECT 11.424 6.6 11.456 9.108 ;
  LAYER M1 ;
        RECT 9.039 6.636 9.041 9.072 ;
  LAYER M1 ;
        RECT 9.119 6.636 9.121 9.072 ;
  LAYER M1 ;
        RECT 9.199 6.636 9.201 9.072 ;
  LAYER M1 ;
        RECT 9.279 6.636 9.281 9.072 ;
  LAYER M1 ;
        RECT 9.359 6.636 9.361 9.072 ;
  LAYER M1 ;
        RECT 9.439 6.636 9.441 9.072 ;
  LAYER M1 ;
        RECT 9.519 6.636 9.521 9.072 ;
  LAYER M1 ;
        RECT 9.599 6.636 9.601 9.072 ;
  LAYER M1 ;
        RECT 9.679 6.636 9.681 9.072 ;
  LAYER M1 ;
        RECT 9.759 6.636 9.761 9.072 ;
  LAYER M1 ;
        RECT 9.839 6.636 9.841 9.072 ;
  LAYER M1 ;
        RECT 9.919 6.636 9.921 9.072 ;
  LAYER M1 ;
        RECT 9.999 6.636 10.001 9.072 ;
  LAYER M1 ;
        RECT 10.079 6.636 10.081 9.072 ;
  LAYER M1 ;
        RECT 10.159 6.636 10.161 9.072 ;
  LAYER M1 ;
        RECT 10.239 6.636 10.241 9.072 ;
  LAYER M1 ;
        RECT 10.319 6.636 10.321 9.072 ;
  LAYER M1 ;
        RECT 10.399 6.636 10.401 9.072 ;
  LAYER M1 ;
        RECT 10.479 6.636 10.481 9.072 ;
  LAYER M1 ;
        RECT 10.559 6.636 10.561 9.072 ;
  LAYER M1 ;
        RECT 10.639 6.636 10.641 9.072 ;
  LAYER M1 ;
        RECT 10.719 6.636 10.721 9.072 ;
  LAYER M1 ;
        RECT 10.799 6.636 10.801 9.072 ;
  LAYER M1 ;
        RECT 10.879 6.636 10.881 9.072 ;
  LAYER M1 ;
        RECT 10.959 6.636 10.961 9.072 ;
  LAYER M1 ;
        RECT 11.039 6.636 11.041 9.072 ;
  LAYER M1 ;
        RECT 11.119 6.636 11.121 9.072 ;
  LAYER M1 ;
        RECT 11.199 6.636 11.201 9.072 ;
  LAYER M1 ;
        RECT 11.279 6.636 11.281 9.072 ;
  LAYER M1 ;
        RECT 11.359 6.636 11.361 9.072 ;
  LAYER M2 ;
        RECT 9.04 6.635 11.44 6.637 ;
  LAYER M2 ;
        RECT 9.04 6.719 11.44 6.721 ;
  LAYER M2 ;
        RECT 9.04 6.803 11.44 6.805 ;
  LAYER M2 ;
        RECT 9.04 6.887 11.44 6.889 ;
  LAYER M2 ;
        RECT 9.04 6.971 11.44 6.973 ;
  LAYER M2 ;
        RECT 9.04 7.055 11.44 7.057 ;
  LAYER M2 ;
        RECT 9.04 7.139 11.44 7.141 ;
  LAYER M2 ;
        RECT 9.04 7.223 11.44 7.225 ;
  LAYER M2 ;
        RECT 9.04 7.307 11.44 7.309 ;
  LAYER M2 ;
        RECT 9.04 7.391 11.44 7.393 ;
  LAYER M2 ;
        RECT 9.04 7.475 11.44 7.477 ;
  LAYER M2 ;
        RECT 9.04 7.559 11.44 7.561 ;
  LAYER M2 ;
        RECT 9.04 7.6425 11.44 7.6445 ;
  LAYER M2 ;
        RECT 9.04 7.727 11.44 7.729 ;
  LAYER M2 ;
        RECT 9.04 7.811 11.44 7.813 ;
  LAYER M2 ;
        RECT 9.04 7.895 11.44 7.897 ;
  LAYER M2 ;
        RECT 9.04 7.979 11.44 7.981 ;
  LAYER M2 ;
        RECT 9.04 8.063 11.44 8.065 ;
  LAYER M2 ;
        RECT 9.04 8.147 11.44 8.149 ;
  LAYER M2 ;
        RECT 9.04 8.231 11.44 8.233 ;
  LAYER M2 ;
        RECT 9.04 8.315 11.44 8.317 ;
  LAYER M2 ;
        RECT 9.04 8.399 11.44 8.401 ;
  LAYER M2 ;
        RECT 9.04 8.483 11.44 8.485 ;
  LAYER M2 ;
        RECT 9.04 8.567 11.44 8.569 ;
  LAYER M2 ;
        RECT 9.04 8.651 11.44 8.653 ;
  LAYER M2 ;
        RECT 9.04 8.735 11.44 8.737 ;
  LAYER M2 ;
        RECT 9.04 8.819 11.44 8.821 ;
  LAYER M2 ;
        RECT 9.04 8.903 11.44 8.905 ;
  LAYER M2 ;
        RECT 9.04 8.987 11.44 8.989 ;
  LAYER M1 ;
        RECT 9.024 9.54 9.056 12.048 ;
  LAYER M1 ;
        RECT 9.088 9.54 9.12 12.048 ;
  LAYER M1 ;
        RECT 9.152 9.54 9.184 12.048 ;
  LAYER M1 ;
        RECT 9.216 9.54 9.248 12.048 ;
  LAYER M1 ;
        RECT 9.28 9.54 9.312 12.048 ;
  LAYER M1 ;
        RECT 9.344 9.54 9.376 12.048 ;
  LAYER M1 ;
        RECT 9.408 9.54 9.44 12.048 ;
  LAYER M1 ;
        RECT 9.472 9.54 9.504 12.048 ;
  LAYER M1 ;
        RECT 9.536 9.54 9.568 12.048 ;
  LAYER M1 ;
        RECT 9.6 9.54 9.632 12.048 ;
  LAYER M1 ;
        RECT 9.664 9.54 9.696 12.048 ;
  LAYER M1 ;
        RECT 9.728 9.54 9.76 12.048 ;
  LAYER M1 ;
        RECT 9.792 9.54 9.824 12.048 ;
  LAYER M1 ;
        RECT 9.856 9.54 9.888 12.048 ;
  LAYER M1 ;
        RECT 9.92 9.54 9.952 12.048 ;
  LAYER M1 ;
        RECT 9.984 9.54 10.016 12.048 ;
  LAYER M1 ;
        RECT 10.048 9.54 10.08 12.048 ;
  LAYER M1 ;
        RECT 10.112 9.54 10.144 12.048 ;
  LAYER M1 ;
        RECT 10.176 9.54 10.208 12.048 ;
  LAYER M1 ;
        RECT 10.24 9.54 10.272 12.048 ;
  LAYER M1 ;
        RECT 10.304 9.54 10.336 12.048 ;
  LAYER M1 ;
        RECT 10.368 9.54 10.4 12.048 ;
  LAYER M1 ;
        RECT 10.432 9.54 10.464 12.048 ;
  LAYER M1 ;
        RECT 10.496 9.54 10.528 12.048 ;
  LAYER M1 ;
        RECT 10.56 9.54 10.592 12.048 ;
  LAYER M1 ;
        RECT 10.624 9.54 10.656 12.048 ;
  LAYER M1 ;
        RECT 10.688 9.54 10.72 12.048 ;
  LAYER M1 ;
        RECT 10.752 9.54 10.784 12.048 ;
  LAYER M1 ;
        RECT 10.816 9.54 10.848 12.048 ;
  LAYER M1 ;
        RECT 10.88 9.54 10.912 12.048 ;
  LAYER M1 ;
        RECT 10.944 9.54 10.976 12.048 ;
  LAYER M1 ;
        RECT 11.008 9.54 11.04 12.048 ;
  LAYER M1 ;
        RECT 11.072 9.54 11.104 12.048 ;
  LAYER M1 ;
        RECT 11.136 9.54 11.168 12.048 ;
  LAYER M1 ;
        RECT 11.2 9.54 11.232 12.048 ;
  LAYER M1 ;
        RECT 11.264 9.54 11.296 12.048 ;
  LAYER M1 ;
        RECT 11.328 9.54 11.36 12.048 ;
  LAYER M2 ;
        RECT 9.004 9.624 11.476 9.656 ;
  LAYER M2 ;
        RECT 9.004 9.688 11.476 9.72 ;
  LAYER M2 ;
        RECT 9.004 9.752 11.476 9.784 ;
  LAYER M2 ;
        RECT 9.004 9.816 11.476 9.848 ;
  LAYER M2 ;
        RECT 9.004 9.88 11.476 9.912 ;
  LAYER M2 ;
        RECT 9.004 9.944 11.476 9.976 ;
  LAYER M2 ;
        RECT 9.004 10.008 11.476 10.04 ;
  LAYER M2 ;
        RECT 9.004 10.072 11.476 10.104 ;
  LAYER M2 ;
        RECT 9.004 10.136 11.476 10.168 ;
  LAYER M2 ;
        RECT 9.004 10.2 11.476 10.232 ;
  LAYER M2 ;
        RECT 9.004 10.264 11.476 10.296 ;
  LAYER M2 ;
        RECT 9.004 10.328 11.476 10.36 ;
  LAYER M2 ;
        RECT 9.004 10.392 11.476 10.424 ;
  LAYER M2 ;
        RECT 9.004 10.456 11.476 10.488 ;
  LAYER M2 ;
        RECT 9.004 10.52 11.476 10.552 ;
  LAYER M2 ;
        RECT 9.004 10.584 11.476 10.616 ;
  LAYER M2 ;
        RECT 9.004 10.648 11.476 10.68 ;
  LAYER M2 ;
        RECT 9.004 10.712 11.476 10.744 ;
  LAYER M2 ;
        RECT 9.004 10.776 11.476 10.808 ;
  LAYER M2 ;
        RECT 9.004 10.84 11.476 10.872 ;
  LAYER M2 ;
        RECT 9.004 10.904 11.476 10.936 ;
  LAYER M2 ;
        RECT 9.004 10.968 11.476 11 ;
  LAYER M2 ;
        RECT 9.004 11.032 11.476 11.064 ;
  LAYER M2 ;
        RECT 9.004 11.096 11.476 11.128 ;
  LAYER M2 ;
        RECT 9.004 11.16 11.476 11.192 ;
  LAYER M2 ;
        RECT 9.004 11.224 11.476 11.256 ;
  LAYER M2 ;
        RECT 9.004 11.288 11.476 11.32 ;
  LAYER M2 ;
        RECT 9.004 11.352 11.476 11.384 ;
  LAYER M2 ;
        RECT 9.004 11.416 11.476 11.448 ;
  LAYER M2 ;
        RECT 9.004 11.48 11.476 11.512 ;
  LAYER M2 ;
        RECT 9.004 11.544 11.476 11.576 ;
  LAYER M2 ;
        RECT 9.004 11.608 11.476 11.64 ;
  LAYER M2 ;
        RECT 9.004 11.672 11.476 11.704 ;
  LAYER M2 ;
        RECT 9.004 11.736 11.476 11.768 ;
  LAYER M2 ;
        RECT 9.004 11.8 11.476 11.832 ;
  LAYER M2 ;
        RECT 9.004 11.864 11.476 11.896 ;
  LAYER M3 ;
        RECT 9.024 9.54 9.056 12.048 ;
  LAYER M3 ;
        RECT 9.088 9.54 9.12 12.048 ;
  LAYER M3 ;
        RECT 9.152 9.54 9.184 12.048 ;
  LAYER M3 ;
        RECT 9.216 9.54 9.248 12.048 ;
  LAYER M3 ;
        RECT 9.28 9.54 9.312 12.048 ;
  LAYER M3 ;
        RECT 9.344 9.54 9.376 12.048 ;
  LAYER M3 ;
        RECT 9.408 9.54 9.44 12.048 ;
  LAYER M3 ;
        RECT 9.472 9.54 9.504 12.048 ;
  LAYER M3 ;
        RECT 9.536 9.54 9.568 12.048 ;
  LAYER M3 ;
        RECT 9.6 9.54 9.632 12.048 ;
  LAYER M3 ;
        RECT 9.664 9.54 9.696 12.048 ;
  LAYER M3 ;
        RECT 9.728 9.54 9.76 12.048 ;
  LAYER M3 ;
        RECT 9.792 9.54 9.824 12.048 ;
  LAYER M3 ;
        RECT 9.856 9.54 9.888 12.048 ;
  LAYER M3 ;
        RECT 9.92 9.54 9.952 12.048 ;
  LAYER M3 ;
        RECT 9.984 9.54 10.016 12.048 ;
  LAYER M3 ;
        RECT 10.048 9.54 10.08 12.048 ;
  LAYER M3 ;
        RECT 10.112 9.54 10.144 12.048 ;
  LAYER M3 ;
        RECT 10.176 9.54 10.208 12.048 ;
  LAYER M3 ;
        RECT 10.24 9.54 10.272 12.048 ;
  LAYER M3 ;
        RECT 10.304 9.54 10.336 12.048 ;
  LAYER M3 ;
        RECT 10.368 9.54 10.4 12.048 ;
  LAYER M3 ;
        RECT 10.432 9.54 10.464 12.048 ;
  LAYER M3 ;
        RECT 10.496 9.54 10.528 12.048 ;
  LAYER M3 ;
        RECT 10.56 9.54 10.592 12.048 ;
  LAYER M3 ;
        RECT 10.624 9.54 10.656 12.048 ;
  LAYER M3 ;
        RECT 10.688 9.54 10.72 12.048 ;
  LAYER M3 ;
        RECT 10.752 9.54 10.784 12.048 ;
  LAYER M3 ;
        RECT 10.816 9.54 10.848 12.048 ;
  LAYER M3 ;
        RECT 10.88 9.54 10.912 12.048 ;
  LAYER M3 ;
        RECT 10.944 9.54 10.976 12.048 ;
  LAYER M3 ;
        RECT 11.008 9.54 11.04 12.048 ;
  LAYER M3 ;
        RECT 11.072 9.54 11.104 12.048 ;
  LAYER M3 ;
        RECT 11.136 9.54 11.168 12.048 ;
  LAYER M3 ;
        RECT 11.2 9.54 11.232 12.048 ;
  LAYER M3 ;
        RECT 11.264 9.54 11.296 12.048 ;
  LAYER M3 ;
        RECT 11.328 9.54 11.36 12.048 ;
  LAYER M3 ;
        RECT 11.424 9.54 11.456 12.048 ;
  LAYER M1 ;
        RECT 9.039 9.576 9.041 12.012 ;
  LAYER M1 ;
        RECT 9.119 9.576 9.121 12.012 ;
  LAYER M1 ;
        RECT 9.199 9.576 9.201 12.012 ;
  LAYER M1 ;
        RECT 9.279 9.576 9.281 12.012 ;
  LAYER M1 ;
        RECT 9.359 9.576 9.361 12.012 ;
  LAYER M1 ;
        RECT 9.439 9.576 9.441 12.012 ;
  LAYER M1 ;
        RECT 9.519 9.576 9.521 12.012 ;
  LAYER M1 ;
        RECT 9.599 9.576 9.601 12.012 ;
  LAYER M1 ;
        RECT 9.679 9.576 9.681 12.012 ;
  LAYER M1 ;
        RECT 9.759 9.576 9.761 12.012 ;
  LAYER M1 ;
        RECT 9.839 9.576 9.841 12.012 ;
  LAYER M1 ;
        RECT 9.919 9.576 9.921 12.012 ;
  LAYER M1 ;
        RECT 9.999 9.576 10.001 12.012 ;
  LAYER M1 ;
        RECT 10.079 9.576 10.081 12.012 ;
  LAYER M1 ;
        RECT 10.159 9.576 10.161 12.012 ;
  LAYER M1 ;
        RECT 10.239 9.576 10.241 12.012 ;
  LAYER M1 ;
        RECT 10.319 9.576 10.321 12.012 ;
  LAYER M1 ;
        RECT 10.399 9.576 10.401 12.012 ;
  LAYER M1 ;
        RECT 10.479 9.576 10.481 12.012 ;
  LAYER M1 ;
        RECT 10.559 9.576 10.561 12.012 ;
  LAYER M1 ;
        RECT 10.639 9.576 10.641 12.012 ;
  LAYER M1 ;
        RECT 10.719 9.576 10.721 12.012 ;
  LAYER M1 ;
        RECT 10.799 9.576 10.801 12.012 ;
  LAYER M1 ;
        RECT 10.879 9.576 10.881 12.012 ;
  LAYER M1 ;
        RECT 10.959 9.576 10.961 12.012 ;
  LAYER M1 ;
        RECT 11.039 9.576 11.041 12.012 ;
  LAYER M1 ;
        RECT 11.119 9.576 11.121 12.012 ;
  LAYER M1 ;
        RECT 11.199 9.576 11.201 12.012 ;
  LAYER M1 ;
        RECT 11.279 9.576 11.281 12.012 ;
  LAYER M1 ;
        RECT 11.359 9.576 11.361 12.012 ;
  LAYER M2 ;
        RECT 9.04 9.575 11.44 9.577 ;
  LAYER M2 ;
        RECT 9.04 9.659 11.44 9.661 ;
  LAYER M2 ;
        RECT 9.04 9.743 11.44 9.745 ;
  LAYER M2 ;
        RECT 9.04 9.827 11.44 9.829 ;
  LAYER M2 ;
        RECT 9.04 9.911 11.44 9.913 ;
  LAYER M2 ;
        RECT 9.04 9.995 11.44 9.997 ;
  LAYER M2 ;
        RECT 9.04 10.079 11.44 10.081 ;
  LAYER M2 ;
        RECT 9.04 10.163 11.44 10.165 ;
  LAYER M2 ;
        RECT 9.04 10.247 11.44 10.249 ;
  LAYER M2 ;
        RECT 9.04 10.331 11.44 10.333 ;
  LAYER M2 ;
        RECT 9.04 10.415 11.44 10.417 ;
  LAYER M2 ;
        RECT 9.04 10.499 11.44 10.501 ;
  LAYER M2 ;
        RECT 9.04 10.5825 11.44 10.5845 ;
  LAYER M2 ;
        RECT 9.04 10.667 11.44 10.669 ;
  LAYER M2 ;
        RECT 9.04 10.751 11.44 10.753 ;
  LAYER M2 ;
        RECT 9.04 10.835 11.44 10.837 ;
  LAYER M2 ;
        RECT 9.04 10.919 11.44 10.921 ;
  LAYER M2 ;
        RECT 9.04 11.003 11.44 11.005 ;
  LAYER M2 ;
        RECT 9.04 11.087 11.44 11.089 ;
  LAYER M2 ;
        RECT 9.04 11.171 11.44 11.173 ;
  LAYER M2 ;
        RECT 9.04 11.255 11.44 11.257 ;
  LAYER M2 ;
        RECT 9.04 11.339 11.44 11.341 ;
  LAYER M2 ;
        RECT 9.04 11.423 11.44 11.425 ;
  LAYER M2 ;
        RECT 9.04 11.507 11.44 11.509 ;
  LAYER M2 ;
        RECT 9.04 11.591 11.44 11.593 ;
  LAYER M2 ;
        RECT 9.04 11.675 11.44 11.677 ;
  LAYER M2 ;
        RECT 9.04 11.759 11.44 11.761 ;
  LAYER M2 ;
        RECT 9.04 11.843 11.44 11.845 ;
  LAYER M2 ;
        RECT 9.04 11.927 11.44 11.929 ;
  LAYER M1 ;
        RECT 9.024 12.48 9.056 14.988 ;
  LAYER M1 ;
        RECT 9.088 12.48 9.12 14.988 ;
  LAYER M1 ;
        RECT 9.152 12.48 9.184 14.988 ;
  LAYER M1 ;
        RECT 9.216 12.48 9.248 14.988 ;
  LAYER M1 ;
        RECT 9.28 12.48 9.312 14.988 ;
  LAYER M1 ;
        RECT 9.344 12.48 9.376 14.988 ;
  LAYER M1 ;
        RECT 9.408 12.48 9.44 14.988 ;
  LAYER M1 ;
        RECT 9.472 12.48 9.504 14.988 ;
  LAYER M1 ;
        RECT 9.536 12.48 9.568 14.988 ;
  LAYER M1 ;
        RECT 9.6 12.48 9.632 14.988 ;
  LAYER M1 ;
        RECT 9.664 12.48 9.696 14.988 ;
  LAYER M1 ;
        RECT 9.728 12.48 9.76 14.988 ;
  LAYER M1 ;
        RECT 9.792 12.48 9.824 14.988 ;
  LAYER M1 ;
        RECT 9.856 12.48 9.888 14.988 ;
  LAYER M1 ;
        RECT 9.92 12.48 9.952 14.988 ;
  LAYER M1 ;
        RECT 9.984 12.48 10.016 14.988 ;
  LAYER M1 ;
        RECT 10.048 12.48 10.08 14.988 ;
  LAYER M1 ;
        RECT 10.112 12.48 10.144 14.988 ;
  LAYER M1 ;
        RECT 10.176 12.48 10.208 14.988 ;
  LAYER M1 ;
        RECT 10.24 12.48 10.272 14.988 ;
  LAYER M1 ;
        RECT 10.304 12.48 10.336 14.988 ;
  LAYER M1 ;
        RECT 10.368 12.48 10.4 14.988 ;
  LAYER M1 ;
        RECT 10.432 12.48 10.464 14.988 ;
  LAYER M1 ;
        RECT 10.496 12.48 10.528 14.988 ;
  LAYER M1 ;
        RECT 10.56 12.48 10.592 14.988 ;
  LAYER M1 ;
        RECT 10.624 12.48 10.656 14.988 ;
  LAYER M1 ;
        RECT 10.688 12.48 10.72 14.988 ;
  LAYER M1 ;
        RECT 10.752 12.48 10.784 14.988 ;
  LAYER M1 ;
        RECT 10.816 12.48 10.848 14.988 ;
  LAYER M1 ;
        RECT 10.88 12.48 10.912 14.988 ;
  LAYER M1 ;
        RECT 10.944 12.48 10.976 14.988 ;
  LAYER M1 ;
        RECT 11.008 12.48 11.04 14.988 ;
  LAYER M1 ;
        RECT 11.072 12.48 11.104 14.988 ;
  LAYER M1 ;
        RECT 11.136 12.48 11.168 14.988 ;
  LAYER M1 ;
        RECT 11.2 12.48 11.232 14.988 ;
  LAYER M1 ;
        RECT 11.264 12.48 11.296 14.988 ;
  LAYER M1 ;
        RECT 11.328 12.48 11.36 14.988 ;
  LAYER M2 ;
        RECT 9.004 12.564 11.476 12.596 ;
  LAYER M2 ;
        RECT 9.004 12.628 11.476 12.66 ;
  LAYER M2 ;
        RECT 9.004 12.692 11.476 12.724 ;
  LAYER M2 ;
        RECT 9.004 12.756 11.476 12.788 ;
  LAYER M2 ;
        RECT 9.004 12.82 11.476 12.852 ;
  LAYER M2 ;
        RECT 9.004 12.884 11.476 12.916 ;
  LAYER M2 ;
        RECT 9.004 12.948 11.476 12.98 ;
  LAYER M2 ;
        RECT 9.004 13.012 11.476 13.044 ;
  LAYER M2 ;
        RECT 9.004 13.076 11.476 13.108 ;
  LAYER M2 ;
        RECT 9.004 13.14 11.476 13.172 ;
  LAYER M2 ;
        RECT 9.004 13.204 11.476 13.236 ;
  LAYER M2 ;
        RECT 9.004 13.268 11.476 13.3 ;
  LAYER M2 ;
        RECT 9.004 13.332 11.476 13.364 ;
  LAYER M2 ;
        RECT 9.004 13.396 11.476 13.428 ;
  LAYER M2 ;
        RECT 9.004 13.46 11.476 13.492 ;
  LAYER M2 ;
        RECT 9.004 13.524 11.476 13.556 ;
  LAYER M2 ;
        RECT 9.004 13.588 11.476 13.62 ;
  LAYER M2 ;
        RECT 9.004 13.652 11.476 13.684 ;
  LAYER M2 ;
        RECT 9.004 13.716 11.476 13.748 ;
  LAYER M2 ;
        RECT 9.004 13.78 11.476 13.812 ;
  LAYER M2 ;
        RECT 9.004 13.844 11.476 13.876 ;
  LAYER M2 ;
        RECT 9.004 13.908 11.476 13.94 ;
  LAYER M2 ;
        RECT 9.004 13.972 11.476 14.004 ;
  LAYER M2 ;
        RECT 9.004 14.036 11.476 14.068 ;
  LAYER M2 ;
        RECT 9.004 14.1 11.476 14.132 ;
  LAYER M2 ;
        RECT 9.004 14.164 11.476 14.196 ;
  LAYER M2 ;
        RECT 9.004 14.228 11.476 14.26 ;
  LAYER M2 ;
        RECT 9.004 14.292 11.476 14.324 ;
  LAYER M2 ;
        RECT 9.004 14.356 11.476 14.388 ;
  LAYER M2 ;
        RECT 9.004 14.42 11.476 14.452 ;
  LAYER M2 ;
        RECT 9.004 14.484 11.476 14.516 ;
  LAYER M2 ;
        RECT 9.004 14.548 11.476 14.58 ;
  LAYER M2 ;
        RECT 9.004 14.612 11.476 14.644 ;
  LAYER M2 ;
        RECT 9.004 14.676 11.476 14.708 ;
  LAYER M2 ;
        RECT 9.004 14.74 11.476 14.772 ;
  LAYER M2 ;
        RECT 9.004 14.804 11.476 14.836 ;
  LAYER M3 ;
        RECT 9.024 12.48 9.056 14.988 ;
  LAYER M3 ;
        RECT 9.088 12.48 9.12 14.988 ;
  LAYER M3 ;
        RECT 9.152 12.48 9.184 14.988 ;
  LAYER M3 ;
        RECT 9.216 12.48 9.248 14.988 ;
  LAYER M3 ;
        RECT 9.28 12.48 9.312 14.988 ;
  LAYER M3 ;
        RECT 9.344 12.48 9.376 14.988 ;
  LAYER M3 ;
        RECT 9.408 12.48 9.44 14.988 ;
  LAYER M3 ;
        RECT 9.472 12.48 9.504 14.988 ;
  LAYER M3 ;
        RECT 9.536 12.48 9.568 14.988 ;
  LAYER M3 ;
        RECT 9.6 12.48 9.632 14.988 ;
  LAYER M3 ;
        RECT 9.664 12.48 9.696 14.988 ;
  LAYER M3 ;
        RECT 9.728 12.48 9.76 14.988 ;
  LAYER M3 ;
        RECT 9.792 12.48 9.824 14.988 ;
  LAYER M3 ;
        RECT 9.856 12.48 9.888 14.988 ;
  LAYER M3 ;
        RECT 9.92 12.48 9.952 14.988 ;
  LAYER M3 ;
        RECT 9.984 12.48 10.016 14.988 ;
  LAYER M3 ;
        RECT 10.048 12.48 10.08 14.988 ;
  LAYER M3 ;
        RECT 10.112 12.48 10.144 14.988 ;
  LAYER M3 ;
        RECT 10.176 12.48 10.208 14.988 ;
  LAYER M3 ;
        RECT 10.24 12.48 10.272 14.988 ;
  LAYER M3 ;
        RECT 10.304 12.48 10.336 14.988 ;
  LAYER M3 ;
        RECT 10.368 12.48 10.4 14.988 ;
  LAYER M3 ;
        RECT 10.432 12.48 10.464 14.988 ;
  LAYER M3 ;
        RECT 10.496 12.48 10.528 14.988 ;
  LAYER M3 ;
        RECT 10.56 12.48 10.592 14.988 ;
  LAYER M3 ;
        RECT 10.624 12.48 10.656 14.988 ;
  LAYER M3 ;
        RECT 10.688 12.48 10.72 14.988 ;
  LAYER M3 ;
        RECT 10.752 12.48 10.784 14.988 ;
  LAYER M3 ;
        RECT 10.816 12.48 10.848 14.988 ;
  LAYER M3 ;
        RECT 10.88 12.48 10.912 14.988 ;
  LAYER M3 ;
        RECT 10.944 12.48 10.976 14.988 ;
  LAYER M3 ;
        RECT 11.008 12.48 11.04 14.988 ;
  LAYER M3 ;
        RECT 11.072 12.48 11.104 14.988 ;
  LAYER M3 ;
        RECT 11.136 12.48 11.168 14.988 ;
  LAYER M3 ;
        RECT 11.2 12.48 11.232 14.988 ;
  LAYER M3 ;
        RECT 11.264 12.48 11.296 14.988 ;
  LAYER M3 ;
        RECT 11.328 12.48 11.36 14.988 ;
  LAYER M3 ;
        RECT 11.424 12.48 11.456 14.988 ;
  LAYER M1 ;
        RECT 9.039 12.516 9.041 14.952 ;
  LAYER M1 ;
        RECT 9.119 12.516 9.121 14.952 ;
  LAYER M1 ;
        RECT 9.199 12.516 9.201 14.952 ;
  LAYER M1 ;
        RECT 9.279 12.516 9.281 14.952 ;
  LAYER M1 ;
        RECT 9.359 12.516 9.361 14.952 ;
  LAYER M1 ;
        RECT 9.439 12.516 9.441 14.952 ;
  LAYER M1 ;
        RECT 9.519 12.516 9.521 14.952 ;
  LAYER M1 ;
        RECT 9.599 12.516 9.601 14.952 ;
  LAYER M1 ;
        RECT 9.679 12.516 9.681 14.952 ;
  LAYER M1 ;
        RECT 9.759 12.516 9.761 14.952 ;
  LAYER M1 ;
        RECT 9.839 12.516 9.841 14.952 ;
  LAYER M1 ;
        RECT 9.919 12.516 9.921 14.952 ;
  LAYER M1 ;
        RECT 9.999 12.516 10.001 14.952 ;
  LAYER M1 ;
        RECT 10.079 12.516 10.081 14.952 ;
  LAYER M1 ;
        RECT 10.159 12.516 10.161 14.952 ;
  LAYER M1 ;
        RECT 10.239 12.516 10.241 14.952 ;
  LAYER M1 ;
        RECT 10.319 12.516 10.321 14.952 ;
  LAYER M1 ;
        RECT 10.399 12.516 10.401 14.952 ;
  LAYER M1 ;
        RECT 10.479 12.516 10.481 14.952 ;
  LAYER M1 ;
        RECT 10.559 12.516 10.561 14.952 ;
  LAYER M1 ;
        RECT 10.639 12.516 10.641 14.952 ;
  LAYER M1 ;
        RECT 10.719 12.516 10.721 14.952 ;
  LAYER M1 ;
        RECT 10.799 12.516 10.801 14.952 ;
  LAYER M1 ;
        RECT 10.879 12.516 10.881 14.952 ;
  LAYER M1 ;
        RECT 10.959 12.516 10.961 14.952 ;
  LAYER M1 ;
        RECT 11.039 12.516 11.041 14.952 ;
  LAYER M1 ;
        RECT 11.119 12.516 11.121 14.952 ;
  LAYER M1 ;
        RECT 11.199 12.516 11.201 14.952 ;
  LAYER M1 ;
        RECT 11.279 12.516 11.281 14.952 ;
  LAYER M1 ;
        RECT 11.359 12.516 11.361 14.952 ;
  LAYER M2 ;
        RECT 9.04 12.515 11.44 12.517 ;
  LAYER M2 ;
        RECT 9.04 12.599 11.44 12.601 ;
  LAYER M2 ;
        RECT 9.04 12.683 11.44 12.685 ;
  LAYER M2 ;
        RECT 9.04 12.767 11.44 12.769 ;
  LAYER M2 ;
        RECT 9.04 12.851 11.44 12.853 ;
  LAYER M2 ;
        RECT 9.04 12.935 11.44 12.937 ;
  LAYER M2 ;
        RECT 9.04 13.019 11.44 13.021 ;
  LAYER M2 ;
        RECT 9.04 13.103 11.44 13.105 ;
  LAYER M2 ;
        RECT 9.04 13.187 11.44 13.189 ;
  LAYER M2 ;
        RECT 9.04 13.271 11.44 13.273 ;
  LAYER M2 ;
        RECT 9.04 13.355 11.44 13.357 ;
  LAYER M2 ;
        RECT 9.04 13.439 11.44 13.441 ;
  LAYER M2 ;
        RECT 9.04 13.5225 11.44 13.5245 ;
  LAYER M2 ;
        RECT 9.04 13.607 11.44 13.609 ;
  LAYER M2 ;
        RECT 9.04 13.691 11.44 13.693 ;
  LAYER M2 ;
        RECT 9.04 13.775 11.44 13.777 ;
  LAYER M2 ;
        RECT 9.04 13.859 11.44 13.861 ;
  LAYER M2 ;
        RECT 9.04 13.943 11.44 13.945 ;
  LAYER M2 ;
        RECT 9.04 14.027 11.44 14.029 ;
  LAYER M2 ;
        RECT 9.04 14.111 11.44 14.113 ;
  LAYER M2 ;
        RECT 9.04 14.195 11.44 14.197 ;
  LAYER M2 ;
        RECT 9.04 14.279 11.44 14.281 ;
  LAYER M2 ;
        RECT 9.04 14.363 11.44 14.365 ;
  LAYER M2 ;
        RECT 9.04 14.447 11.44 14.449 ;
  LAYER M2 ;
        RECT 9.04 14.531 11.44 14.533 ;
  LAYER M2 ;
        RECT 9.04 14.615 11.44 14.617 ;
  LAYER M2 ;
        RECT 9.04 14.699 11.44 14.701 ;
  LAYER M2 ;
        RECT 9.04 14.783 11.44 14.785 ;
  LAYER M2 ;
        RECT 9.04 14.867 11.44 14.869 ;
  LAYER M1 ;
        RECT 9.024 15.42 9.056 17.928 ;
  LAYER M1 ;
        RECT 9.088 15.42 9.12 17.928 ;
  LAYER M1 ;
        RECT 9.152 15.42 9.184 17.928 ;
  LAYER M1 ;
        RECT 9.216 15.42 9.248 17.928 ;
  LAYER M1 ;
        RECT 9.28 15.42 9.312 17.928 ;
  LAYER M1 ;
        RECT 9.344 15.42 9.376 17.928 ;
  LAYER M1 ;
        RECT 9.408 15.42 9.44 17.928 ;
  LAYER M1 ;
        RECT 9.472 15.42 9.504 17.928 ;
  LAYER M1 ;
        RECT 9.536 15.42 9.568 17.928 ;
  LAYER M1 ;
        RECT 9.6 15.42 9.632 17.928 ;
  LAYER M1 ;
        RECT 9.664 15.42 9.696 17.928 ;
  LAYER M1 ;
        RECT 9.728 15.42 9.76 17.928 ;
  LAYER M1 ;
        RECT 9.792 15.42 9.824 17.928 ;
  LAYER M1 ;
        RECT 9.856 15.42 9.888 17.928 ;
  LAYER M1 ;
        RECT 9.92 15.42 9.952 17.928 ;
  LAYER M1 ;
        RECT 9.984 15.42 10.016 17.928 ;
  LAYER M1 ;
        RECT 10.048 15.42 10.08 17.928 ;
  LAYER M1 ;
        RECT 10.112 15.42 10.144 17.928 ;
  LAYER M1 ;
        RECT 10.176 15.42 10.208 17.928 ;
  LAYER M1 ;
        RECT 10.24 15.42 10.272 17.928 ;
  LAYER M1 ;
        RECT 10.304 15.42 10.336 17.928 ;
  LAYER M1 ;
        RECT 10.368 15.42 10.4 17.928 ;
  LAYER M1 ;
        RECT 10.432 15.42 10.464 17.928 ;
  LAYER M1 ;
        RECT 10.496 15.42 10.528 17.928 ;
  LAYER M1 ;
        RECT 10.56 15.42 10.592 17.928 ;
  LAYER M1 ;
        RECT 10.624 15.42 10.656 17.928 ;
  LAYER M1 ;
        RECT 10.688 15.42 10.72 17.928 ;
  LAYER M1 ;
        RECT 10.752 15.42 10.784 17.928 ;
  LAYER M1 ;
        RECT 10.816 15.42 10.848 17.928 ;
  LAYER M1 ;
        RECT 10.88 15.42 10.912 17.928 ;
  LAYER M1 ;
        RECT 10.944 15.42 10.976 17.928 ;
  LAYER M1 ;
        RECT 11.008 15.42 11.04 17.928 ;
  LAYER M1 ;
        RECT 11.072 15.42 11.104 17.928 ;
  LAYER M1 ;
        RECT 11.136 15.42 11.168 17.928 ;
  LAYER M1 ;
        RECT 11.2 15.42 11.232 17.928 ;
  LAYER M1 ;
        RECT 11.264 15.42 11.296 17.928 ;
  LAYER M1 ;
        RECT 11.328 15.42 11.36 17.928 ;
  LAYER M2 ;
        RECT 9.004 15.504 11.476 15.536 ;
  LAYER M2 ;
        RECT 9.004 15.568 11.476 15.6 ;
  LAYER M2 ;
        RECT 9.004 15.632 11.476 15.664 ;
  LAYER M2 ;
        RECT 9.004 15.696 11.476 15.728 ;
  LAYER M2 ;
        RECT 9.004 15.76 11.476 15.792 ;
  LAYER M2 ;
        RECT 9.004 15.824 11.476 15.856 ;
  LAYER M2 ;
        RECT 9.004 15.888 11.476 15.92 ;
  LAYER M2 ;
        RECT 9.004 15.952 11.476 15.984 ;
  LAYER M2 ;
        RECT 9.004 16.016 11.476 16.048 ;
  LAYER M2 ;
        RECT 9.004 16.08 11.476 16.112 ;
  LAYER M2 ;
        RECT 9.004 16.144 11.476 16.176 ;
  LAYER M2 ;
        RECT 9.004 16.208 11.476 16.24 ;
  LAYER M2 ;
        RECT 9.004 16.272 11.476 16.304 ;
  LAYER M2 ;
        RECT 9.004 16.336 11.476 16.368 ;
  LAYER M2 ;
        RECT 9.004 16.4 11.476 16.432 ;
  LAYER M2 ;
        RECT 9.004 16.464 11.476 16.496 ;
  LAYER M2 ;
        RECT 9.004 16.528 11.476 16.56 ;
  LAYER M2 ;
        RECT 9.004 16.592 11.476 16.624 ;
  LAYER M2 ;
        RECT 9.004 16.656 11.476 16.688 ;
  LAYER M2 ;
        RECT 9.004 16.72 11.476 16.752 ;
  LAYER M2 ;
        RECT 9.004 16.784 11.476 16.816 ;
  LAYER M2 ;
        RECT 9.004 16.848 11.476 16.88 ;
  LAYER M2 ;
        RECT 9.004 16.912 11.476 16.944 ;
  LAYER M2 ;
        RECT 9.004 16.976 11.476 17.008 ;
  LAYER M2 ;
        RECT 9.004 17.04 11.476 17.072 ;
  LAYER M2 ;
        RECT 9.004 17.104 11.476 17.136 ;
  LAYER M2 ;
        RECT 9.004 17.168 11.476 17.2 ;
  LAYER M2 ;
        RECT 9.004 17.232 11.476 17.264 ;
  LAYER M2 ;
        RECT 9.004 17.296 11.476 17.328 ;
  LAYER M2 ;
        RECT 9.004 17.36 11.476 17.392 ;
  LAYER M2 ;
        RECT 9.004 17.424 11.476 17.456 ;
  LAYER M2 ;
        RECT 9.004 17.488 11.476 17.52 ;
  LAYER M2 ;
        RECT 9.004 17.552 11.476 17.584 ;
  LAYER M2 ;
        RECT 9.004 17.616 11.476 17.648 ;
  LAYER M2 ;
        RECT 9.004 17.68 11.476 17.712 ;
  LAYER M2 ;
        RECT 9.004 17.744 11.476 17.776 ;
  LAYER M3 ;
        RECT 9.024 15.42 9.056 17.928 ;
  LAYER M3 ;
        RECT 9.088 15.42 9.12 17.928 ;
  LAYER M3 ;
        RECT 9.152 15.42 9.184 17.928 ;
  LAYER M3 ;
        RECT 9.216 15.42 9.248 17.928 ;
  LAYER M3 ;
        RECT 9.28 15.42 9.312 17.928 ;
  LAYER M3 ;
        RECT 9.344 15.42 9.376 17.928 ;
  LAYER M3 ;
        RECT 9.408 15.42 9.44 17.928 ;
  LAYER M3 ;
        RECT 9.472 15.42 9.504 17.928 ;
  LAYER M3 ;
        RECT 9.536 15.42 9.568 17.928 ;
  LAYER M3 ;
        RECT 9.6 15.42 9.632 17.928 ;
  LAYER M3 ;
        RECT 9.664 15.42 9.696 17.928 ;
  LAYER M3 ;
        RECT 9.728 15.42 9.76 17.928 ;
  LAYER M3 ;
        RECT 9.792 15.42 9.824 17.928 ;
  LAYER M3 ;
        RECT 9.856 15.42 9.888 17.928 ;
  LAYER M3 ;
        RECT 9.92 15.42 9.952 17.928 ;
  LAYER M3 ;
        RECT 9.984 15.42 10.016 17.928 ;
  LAYER M3 ;
        RECT 10.048 15.42 10.08 17.928 ;
  LAYER M3 ;
        RECT 10.112 15.42 10.144 17.928 ;
  LAYER M3 ;
        RECT 10.176 15.42 10.208 17.928 ;
  LAYER M3 ;
        RECT 10.24 15.42 10.272 17.928 ;
  LAYER M3 ;
        RECT 10.304 15.42 10.336 17.928 ;
  LAYER M3 ;
        RECT 10.368 15.42 10.4 17.928 ;
  LAYER M3 ;
        RECT 10.432 15.42 10.464 17.928 ;
  LAYER M3 ;
        RECT 10.496 15.42 10.528 17.928 ;
  LAYER M3 ;
        RECT 10.56 15.42 10.592 17.928 ;
  LAYER M3 ;
        RECT 10.624 15.42 10.656 17.928 ;
  LAYER M3 ;
        RECT 10.688 15.42 10.72 17.928 ;
  LAYER M3 ;
        RECT 10.752 15.42 10.784 17.928 ;
  LAYER M3 ;
        RECT 10.816 15.42 10.848 17.928 ;
  LAYER M3 ;
        RECT 10.88 15.42 10.912 17.928 ;
  LAYER M3 ;
        RECT 10.944 15.42 10.976 17.928 ;
  LAYER M3 ;
        RECT 11.008 15.42 11.04 17.928 ;
  LAYER M3 ;
        RECT 11.072 15.42 11.104 17.928 ;
  LAYER M3 ;
        RECT 11.136 15.42 11.168 17.928 ;
  LAYER M3 ;
        RECT 11.2 15.42 11.232 17.928 ;
  LAYER M3 ;
        RECT 11.264 15.42 11.296 17.928 ;
  LAYER M3 ;
        RECT 11.328 15.42 11.36 17.928 ;
  LAYER M3 ;
        RECT 11.424 15.42 11.456 17.928 ;
  LAYER M1 ;
        RECT 9.039 15.456 9.041 17.892 ;
  LAYER M1 ;
        RECT 9.119 15.456 9.121 17.892 ;
  LAYER M1 ;
        RECT 9.199 15.456 9.201 17.892 ;
  LAYER M1 ;
        RECT 9.279 15.456 9.281 17.892 ;
  LAYER M1 ;
        RECT 9.359 15.456 9.361 17.892 ;
  LAYER M1 ;
        RECT 9.439 15.456 9.441 17.892 ;
  LAYER M1 ;
        RECT 9.519 15.456 9.521 17.892 ;
  LAYER M1 ;
        RECT 9.599 15.456 9.601 17.892 ;
  LAYER M1 ;
        RECT 9.679 15.456 9.681 17.892 ;
  LAYER M1 ;
        RECT 9.759 15.456 9.761 17.892 ;
  LAYER M1 ;
        RECT 9.839 15.456 9.841 17.892 ;
  LAYER M1 ;
        RECT 9.919 15.456 9.921 17.892 ;
  LAYER M1 ;
        RECT 9.999 15.456 10.001 17.892 ;
  LAYER M1 ;
        RECT 10.079 15.456 10.081 17.892 ;
  LAYER M1 ;
        RECT 10.159 15.456 10.161 17.892 ;
  LAYER M1 ;
        RECT 10.239 15.456 10.241 17.892 ;
  LAYER M1 ;
        RECT 10.319 15.456 10.321 17.892 ;
  LAYER M1 ;
        RECT 10.399 15.456 10.401 17.892 ;
  LAYER M1 ;
        RECT 10.479 15.456 10.481 17.892 ;
  LAYER M1 ;
        RECT 10.559 15.456 10.561 17.892 ;
  LAYER M1 ;
        RECT 10.639 15.456 10.641 17.892 ;
  LAYER M1 ;
        RECT 10.719 15.456 10.721 17.892 ;
  LAYER M1 ;
        RECT 10.799 15.456 10.801 17.892 ;
  LAYER M1 ;
        RECT 10.879 15.456 10.881 17.892 ;
  LAYER M1 ;
        RECT 10.959 15.456 10.961 17.892 ;
  LAYER M1 ;
        RECT 11.039 15.456 11.041 17.892 ;
  LAYER M1 ;
        RECT 11.119 15.456 11.121 17.892 ;
  LAYER M1 ;
        RECT 11.199 15.456 11.201 17.892 ;
  LAYER M1 ;
        RECT 11.279 15.456 11.281 17.892 ;
  LAYER M1 ;
        RECT 11.359 15.456 11.361 17.892 ;
  LAYER M2 ;
        RECT 9.04 15.455 11.44 15.457 ;
  LAYER M2 ;
        RECT 9.04 15.539 11.44 15.541 ;
  LAYER M2 ;
        RECT 9.04 15.623 11.44 15.625 ;
  LAYER M2 ;
        RECT 9.04 15.707 11.44 15.709 ;
  LAYER M2 ;
        RECT 9.04 15.791 11.44 15.793 ;
  LAYER M2 ;
        RECT 9.04 15.875 11.44 15.877 ;
  LAYER M2 ;
        RECT 9.04 15.959 11.44 15.961 ;
  LAYER M2 ;
        RECT 9.04 16.043 11.44 16.045 ;
  LAYER M2 ;
        RECT 9.04 16.127 11.44 16.129 ;
  LAYER M2 ;
        RECT 9.04 16.211 11.44 16.213 ;
  LAYER M2 ;
        RECT 9.04 16.295 11.44 16.297 ;
  LAYER M2 ;
        RECT 9.04 16.379 11.44 16.381 ;
  LAYER M2 ;
        RECT 9.04 16.4625 11.44 16.4645 ;
  LAYER M2 ;
        RECT 9.04 16.547 11.44 16.549 ;
  LAYER M2 ;
        RECT 9.04 16.631 11.44 16.633 ;
  LAYER M2 ;
        RECT 9.04 16.715 11.44 16.717 ;
  LAYER M2 ;
        RECT 9.04 16.799 11.44 16.801 ;
  LAYER M2 ;
        RECT 9.04 16.883 11.44 16.885 ;
  LAYER M2 ;
        RECT 9.04 16.967 11.44 16.969 ;
  LAYER M2 ;
        RECT 9.04 17.051 11.44 17.053 ;
  LAYER M2 ;
        RECT 9.04 17.135 11.44 17.137 ;
  LAYER M2 ;
        RECT 9.04 17.219 11.44 17.221 ;
  LAYER M2 ;
        RECT 9.04 17.303 11.44 17.305 ;
  LAYER M2 ;
        RECT 9.04 17.387 11.44 17.389 ;
  LAYER M2 ;
        RECT 9.04 17.471 11.44 17.473 ;
  LAYER M2 ;
        RECT 9.04 17.555 11.44 17.557 ;
  LAYER M2 ;
        RECT 9.04 17.639 11.44 17.641 ;
  LAYER M2 ;
        RECT 9.04 17.723 11.44 17.725 ;
  LAYER M2 ;
        RECT 9.04 17.807 11.44 17.809 ;
  END 
END Cap_60fF
