MACRO Cap_12f
  ORIGIN 0 0 ;
  FOREIGN Cap_12f 0 0 ;
  SIZE 2.4000 BY 2.4360 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 -0.0160 2.4360 0.0160 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 2.4200 2.4360 2.4520 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
  END
END Cap_12f
MACRO Res_r20000
  ORIGIN 0 0 ;
  FOREIGN Res_r20000 0 0 ;
  SIZE 1.0400 BY 1.7640 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.3560 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6040 0.0680 0.9320 0.1000 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 1.7160 ;
    LAYER M1 ;
      RECT 0.3040 1.6640 0.4000 1.6960 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 1.7160 ;
    LAYER M1 ;
      RECT 0.3680 0.0680 0.4640 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 1.7160 ;
    LAYER M1 ;
      RECT 0.4320 1.6640 0.5280 1.6960 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 1.7160 ;
    LAYER M1 ;
      RECT 0.4960 0.0680 0.5920 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 1.7160 ;
    LAYER M1 ;
      RECT 0.5600 1.6640 0.6560 1.6960 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 1.7160 ;
    LAYER V1 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
  END
END Res_r20000
MACRO Switch_NMOS_nfin48_n12_X2_Y2_ST2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin48_n12_X2_Y2_ST2 0 0 ;
  SIZE 1.1200 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.8880 0.5000 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.7560 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 0.7560 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 2.6720 0.7560 2.7040 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 0.7560 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 0.7560 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
  END
END Switch_NMOS_nfin48_n12_X2_Y2_ST2
MACRO Res_r500
  ORIGIN 0 0 ;
  FOREIGN Res_r500 0 0 ;
  SIZE 1.0400 BY 1.7640 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.3560 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6040 0.0680 0.9320 0.1000 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 1.7160 ;
    LAYER M1 ;
      RECT 0.3040 1.6640 0.4000 1.6960 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 1.7160 ;
    LAYER M1 ;
      RECT 0.3680 0.0680 0.4640 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 1.7160 ;
    LAYER M1 ;
      RECT 0.4320 1.6640 0.5280 1.6960 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 1.7160 ;
    LAYER M1 ;
      RECT 0.4960 0.0680 0.5920 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 1.7160 ;
    LAYER M1 ;
      RECT 0.5600 1.6640 0.6560 1.6960 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 1.7160 ;
    LAYER V1 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
  END
END Res_r500
MACRO Switch_PMOS_nfin48_n12_X2_Y2_ST2
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin48_n12_X2_Y2_ST2 0 0 ;
  SIZE 1.1200 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.8880 0.5000 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.7560 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 0.7560 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 2.6720 0.7560 2.7040 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 0.7560 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 0.7560 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V2 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
  END
END Switch_PMOS_nfin48_n12_X2_Y2_ST2
