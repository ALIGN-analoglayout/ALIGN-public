MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 15.76 BY 23.1 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.844 22.644 2.876 22.716 ;
      LAYER M2 ;
        RECT 2.824 22.664 2.896 22.696 ;
      LAYER M1 ;
        RECT 12.796 22.644 12.828 22.716 ;
      LAYER M2 ;
        RECT 12.776 22.664 12.848 22.696 ;
      LAYER M2 ;
        RECT 2.86 22.664 12.812 22.696 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.98 0.384 6.012 0.456 ;
      LAYER M2 ;
        RECT 5.96 0.404 6.032 0.436 ;
      LAYER M1 ;
        RECT 9.276 0.384 9.308 0.456 ;
      LAYER M2 ;
        RECT 9.256 0.404 9.328 0.436 ;
      LAYER M2 ;
        RECT 5.996 0.404 9.292 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.364 22.812 6.396 22.884 ;
      LAYER M2 ;
        RECT 6.344 22.832 6.416 22.864 ;
      LAYER M1 ;
        RECT 9.596 22.812 9.628 22.884 ;
      LAYER M2 ;
        RECT 9.576 22.832 9.648 22.864 ;
      LAYER M2 ;
        RECT 6.38 22.832 9.612 22.864 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.684 0.216 2.716 0.288 ;
      LAYER M2 ;
        RECT 2.664 0.236 2.736 0.268 ;
      LAYER M1 ;
        RECT 12.572 0.216 12.604 0.288 ;
      LAYER M2 ;
        RECT 12.552 0.236 12.624 0.268 ;
      LAYER M2 ;
        RECT 2.7 0.236 12.588 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 9.052 7.188 9.084 7.26 ;
  LAYER M2 ;
        RECT 9.032 7.208 9.104 7.24 ;
  LAYER M2 ;
        RECT 5.996 7.208 9.068 7.24 ;
  LAYER M1 ;
        RECT 5.98 7.188 6.012 7.26 ;
  LAYER M2 ;
        RECT 5.96 7.208 6.032 7.24 ;
  LAYER M1 ;
        RECT 9.052 13.404 9.084 13.476 ;
  LAYER M2 ;
        RECT 9.032 13.424 9.104 13.456 ;
  LAYER M2 ;
        RECT 5.996 13.424 9.068 13.456 ;
  LAYER M1 ;
        RECT 5.98 13.404 6.012 13.476 ;
  LAYER M2 ;
        RECT 5.96 13.424 6.032 13.456 ;
  LAYER M1 ;
        RECT 5.756 10.296 5.788 10.368 ;
  LAYER M2 ;
        RECT 5.736 10.316 5.808 10.348 ;
  LAYER M1 ;
        RECT 5.756 10.164 5.788 10.332 ;
  LAYER M1 ;
        RECT 5.756 10.128 5.788 10.2 ;
  LAYER M2 ;
        RECT 5.736 10.148 5.808 10.18 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.996 10.18 ;
  LAYER M1 ;
        RECT 5.98 10.128 6.012 10.2 ;
  LAYER M2 ;
        RECT 5.96 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 5.756 7.188 5.788 7.26 ;
  LAYER M2 ;
        RECT 5.736 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 5.756 7.056 5.788 7.224 ;
  LAYER M1 ;
        RECT 5.756 7.02 5.788 7.092 ;
  LAYER M2 ;
        RECT 5.736 7.04 5.808 7.072 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.996 7.072 ;
  LAYER M1 ;
        RECT 5.98 7.02 6.012 7.092 ;
  LAYER M2 ;
        RECT 5.96 7.04 6.032 7.072 ;
  LAYER M1 ;
        RECT 5.98 0.384 6.012 0.456 ;
  LAYER M2 ;
        RECT 5.96 0.404 6.032 0.436 ;
  LAYER M1 ;
        RECT 5.98 0.42 6.012 0.672 ;
  LAYER M1 ;
        RECT 5.98 0.672 6.012 13.44 ;
  LAYER M1 ;
        RECT 12.348 10.296 12.38 10.368 ;
  LAYER M2 ;
        RECT 12.328 10.316 12.4 10.348 ;
  LAYER M2 ;
        RECT 9.292 10.316 12.364 10.348 ;
  LAYER M1 ;
        RECT 9.276 10.296 9.308 10.368 ;
  LAYER M2 ;
        RECT 9.256 10.316 9.328 10.348 ;
  LAYER M1 ;
        RECT 12.348 13.404 12.38 13.476 ;
  LAYER M2 ;
        RECT 12.328 13.424 12.4 13.456 ;
  LAYER M2 ;
        RECT 9.292 13.424 12.364 13.456 ;
  LAYER M1 ;
        RECT 9.276 13.404 9.308 13.476 ;
  LAYER M2 ;
        RECT 9.256 13.424 9.328 13.456 ;
  LAYER M1 ;
        RECT 9.276 0.384 9.308 0.456 ;
  LAYER M2 ;
        RECT 9.256 0.404 9.328 0.436 ;
  LAYER M1 ;
        RECT 9.276 0.42 9.308 0.672 ;
  LAYER M1 ;
        RECT 9.276 0.672 9.308 13.44 ;
  LAYER M2 ;
        RECT 5.996 0.404 9.292 0.436 ;
  LAYER M1 ;
        RECT 5.756 13.404 5.788 13.476 ;
  LAYER M2 ;
        RECT 5.736 13.424 5.808 13.456 ;
  LAYER M2 ;
        RECT 2.7 13.424 5.772 13.456 ;
  LAYER M1 ;
        RECT 2.684 13.404 2.716 13.476 ;
  LAYER M2 ;
        RECT 2.664 13.424 2.736 13.456 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 16.584 ;
  LAYER M2 ;
        RECT 5.736 16.532 5.808 16.564 ;
  LAYER M2 ;
        RECT 2.7 16.532 5.772 16.564 ;
  LAYER M1 ;
        RECT 2.684 16.512 2.716 16.584 ;
  LAYER M2 ;
        RECT 2.664 16.532 2.736 16.564 ;
  LAYER M1 ;
        RECT 2.684 0.216 2.716 0.288 ;
  LAYER M2 ;
        RECT 2.664 0.236 2.736 0.268 ;
  LAYER M1 ;
        RECT 2.684 0.252 2.716 0.672 ;
  LAYER M1 ;
        RECT 2.684 0.672 2.716 16.548 ;
  LAYER M1 ;
        RECT 12.348 7.188 12.38 7.26 ;
  LAYER M2 ;
        RECT 12.328 7.208 12.4 7.24 ;
  LAYER M1 ;
        RECT 12.348 7.056 12.38 7.224 ;
  LAYER M1 ;
        RECT 12.348 7.02 12.38 7.092 ;
  LAYER M2 ;
        RECT 12.328 7.04 12.4 7.072 ;
  LAYER M2 ;
        RECT 12.364 7.04 12.588 7.072 ;
  LAYER M1 ;
        RECT 12.572 7.02 12.604 7.092 ;
  LAYER M2 ;
        RECT 12.552 7.04 12.624 7.072 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 4.152 ;
  LAYER M2 ;
        RECT 12.328 4.1 12.4 4.132 ;
  LAYER M1 ;
        RECT 12.348 3.948 12.38 4.116 ;
  LAYER M1 ;
        RECT 12.348 3.912 12.38 3.984 ;
  LAYER M2 ;
        RECT 12.328 3.932 12.4 3.964 ;
  LAYER M2 ;
        RECT 12.364 3.932 12.588 3.964 ;
  LAYER M1 ;
        RECT 12.572 3.912 12.604 3.984 ;
  LAYER M2 ;
        RECT 12.552 3.932 12.624 3.964 ;
  LAYER M1 ;
        RECT 12.572 0.216 12.604 0.288 ;
  LAYER M2 ;
        RECT 12.552 0.236 12.624 0.268 ;
  LAYER M1 ;
        RECT 12.572 0.252 12.604 0.672 ;
  LAYER M1 ;
        RECT 12.572 0.672 12.604 7.056 ;
  LAYER M2 ;
        RECT 2.7 0.236 12.588 0.268 ;
  LAYER M1 ;
        RECT 9.052 16.512 9.084 16.584 ;
  LAYER M2 ;
        RECT 9.032 16.532 9.104 16.564 ;
  LAYER M2 ;
        RECT 5.772 16.532 9.068 16.564 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 16.584 ;
  LAYER M2 ;
        RECT 5.736 16.532 5.808 16.564 ;
  LAYER M1 ;
        RECT 9.052 4.08 9.084 4.152 ;
  LAYER M2 ;
        RECT 9.032 4.1 9.104 4.132 ;
  LAYER M2 ;
        RECT 9.068 4.1 12.364 4.132 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 4.152 ;
  LAYER M2 ;
        RECT 12.328 4.1 12.4 4.132 ;
  LAYER M1 ;
        RECT 5.756 0.972 5.788 1.044 ;
  LAYER M2 ;
        RECT 5.736 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 5.756 0.84 5.788 1.008 ;
  LAYER M1 ;
        RECT 5.756 0.804 5.788 0.876 ;
  LAYER M2 ;
        RECT 5.736 0.824 5.808 0.856 ;
  LAYER M2 ;
        RECT 5.772 0.824 6.156 0.856 ;
  LAYER M1 ;
        RECT 6.14 0.804 6.172 0.876 ;
  LAYER M2 ;
        RECT 6.12 0.824 6.192 0.856 ;
  LAYER M1 ;
        RECT 5.756 4.08 5.788 4.152 ;
  LAYER M2 ;
        RECT 5.736 4.1 5.808 4.132 ;
  LAYER M1 ;
        RECT 5.756 3.948 5.788 4.116 ;
  LAYER M1 ;
        RECT 5.756 3.912 5.788 3.984 ;
  LAYER M2 ;
        RECT 5.736 3.932 5.808 3.964 ;
  LAYER M2 ;
        RECT 5.772 3.932 6.156 3.964 ;
  LAYER M1 ;
        RECT 6.14 3.912 6.172 3.984 ;
  LAYER M2 ;
        RECT 6.12 3.932 6.192 3.964 ;
  LAYER M1 ;
        RECT 5.756 19.62 5.788 19.692 ;
  LAYER M2 ;
        RECT 5.736 19.64 5.808 19.672 ;
  LAYER M1 ;
        RECT 5.756 19.488 5.788 19.656 ;
  LAYER M1 ;
        RECT 5.756 19.452 5.788 19.524 ;
  LAYER M2 ;
        RECT 5.736 19.472 5.808 19.504 ;
  LAYER M2 ;
        RECT 5.772 19.472 6.156 19.504 ;
  LAYER M1 ;
        RECT 6.14 19.452 6.172 19.524 ;
  LAYER M2 ;
        RECT 6.12 19.472 6.192 19.504 ;
  LAYER M1 ;
        RECT 9.052 0.972 9.084 1.044 ;
  LAYER M2 ;
        RECT 9.032 0.992 9.104 1.024 ;
  LAYER M2 ;
        RECT 6.156 0.992 9.068 1.024 ;
  LAYER M1 ;
        RECT 6.14 0.972 6.172 1.044 ;
  LAYER M2 ;
        RECT 6.12 0.992 6.192 1.024 ;
  LAYER M1 ;
        RECT 9.052 10.296 9.084 10.368 ;
  LAYER M2 ;
        RECT 9.032 10.316 9.104 10.348 ;
  LAYER M2 ;
        RECT 6.156 10.316 9.068 10.348 ;
  LAYER M1 ;
        RECT 6.14 10.296 6.172 10.368 ;
  LAYER M2 ;
        RECT 6.12 10.316 6.192 10.348 ;
  LAYER M1 ;
        RECT 9.052 19.62 9.084 19.692 ;
  LAYER M2 ;
        RECT 9.032 19.64 9.104 19.672 ;
  LAYER M2 ;
        RECT 6.156 19.64 9.068 19.672 ;
  LAYER M1 ;
        RECT 6.14 19.62 6.172 19.692 ;
  LAYER M2 ;
        RECT 6.12 19.64 6.192 19.672 ;
  LAYER M1 ;
        RECT 6.14 0.048 6.172 0.12 ;
  LAYER M2 ;
        RECT 6.12 0.068 6.192 0.1 ;
  LAYER M1 ;
        RECT 6.14 0.084 6.172 0.672 ;
  LAYER M1 ;
        RECT 6.14 0.672 6.172 19.656 ;
  LAYER M1 ;
        RECT 12.348 0.972 12.38 1.044 ;
  LAYER M2 ;
        RECT 12.328 0.992 12.4 1.024 ;
  LAYER M2 ;
        RECT 9.452 0.992 12.364 1.024 ;
  LAYER M1 ;
        RECT 9.436 0.972 9.468 1.044 ;
  LAYER M2 ;
        RECT 9.416 0.992 9.488 1.024 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 16.584 ;
  LAYER M2 ;
        RECT 12.328 16.532 12.4 16.564 ;
  LAYER M2 ;
        RECT 9.452 16.532 12.364 16.564 ;
  LAYER M1 ;
        RECT 9.436 16.512 9.468 16.584 ;
  LAYER M2 ;
        RECT 9.416 16.532 9.488 16.564 ;
  LAYER M1 ;
        RECT 12.348 19.62 12.38 19.692 ;
  LAYER M2 ;
        RECT 12.328 19.64 12.4 19.672 ;
  LAYER M2 ;
        RECT 9.452 19.64 12.364 19.672 ;
  LAYER M1 ;
        RECT 9.436 19.62 9.468 19.692 ;
  LAYER M2 ;
        RECT 9.416 19.64 9.488 19.672 ;
  LAYER M1 ;
        RECT 9.436 0.048 9.468 0.12 ;
  LAYER M2 ;
        RECT 9.416 0.068 9.488 0.1 ;
  LAYER M1 ;
        RECT 9.436 0.084 9.468 0.672 ;
  LAYER M1 ;
        RECT 9.436 0.672 9.468 19.656 ;
  LAYER M2 ;
        RECT 6.156 0.068 9.452 0.1 ;
  LAYER M1 ;
        RECT 2.46 19.62 2.492 19.692 ;
  LAYER M2 ;
        RECT 2.44 19.64 2.512 19.672 ;
  LAYER M2 ;
        RECT 2.476 19.64 5.772 19.672 ;
  LAYER M1 ;
        RECT 5.756 19.62 5.788 19.692 ;
  LAYER M2 ;
        RECT 5.736 19.64 5.808 19.672 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 16.548 2.492 19.656 ;
  LAYER M1 ;
        RECT 2.46 19.62 2.492 19.692 ;
  LAYER M2 ;
        RECT 2.44 19.64 2.512 19.672 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 13.44 2.492 16.548 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 10.332 2.492 13.44 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 7.224 2.492 10.332 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 2.46 4.116 2.492 7.224 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 1.044 ;
  LAYER M2 ;
        RECT 2.44 0.992 2.512 1.024 ;
  LAYER M1 ;
        RECT 2.46 1.008 2.492 4.116 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 15.644 19.62 15.676 19.692 ;
  LAYER M2 ;
        RECT 15.624 19.64 15.696 19.672 ;
  LAYER M2 ;
        RECT 12.364 19.64 15.66 19.672 ;
  LAYER M1 ;
        RECT 12.348 19.62 12.38 19.692 ;
  LAYER M2 ;
        RECT 12.328 19.64 12.4 19.672 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 16.584 ;
  LAYER M2 ;
        RECT 15.624 16.532 15.696 16.564 ;
  LAYER M2 ;
        RECT 12.364 16.532 15.66 16.564 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 16.584 ;
  LAYER M2 ;
        RECT 12.328 16.532 12.4 16.564 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 13.476 ;
  LAYER M2 ;
        RECT 15.624 13.424 15.696 13.456 ;
  LAYER M1 ;
        RECT 15.644 13.44 15.676 16.548 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 16.584 ;
  LAYER M2 ;
        RECT 15.624 16.532 15.696 16.564 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 10.368 ;
  LAYER M2 ;
        RECT 15.624 10.316 15.696 10.348 ;
  LAYER M1 ;
        RECT 15.644 10.332 15.676 13.44 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 13.476 ;
  LAYER M2 ;
        RECT 15.624 13.424 15.696 13.456 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 7.26 ;
  LAYER M2 ;
        RECT 15.624 7.208 15.696 7.24 ;
  LAYER M1 ;
        RECT 15.644 7.224 15.676 10.332 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 10.368 ;
  LAYER M2 ;
        RECT 15.624 10.316 15.696 10.348 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 4.152 ;
  LAYER M2 ;
        RECT 15.624 4.1 15.696 4.132 ;
  LAYER M1 ;
        RECT 15.644 4.116 15.676 7.224 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 7.26 ;
  LAYER M2 ;
        RECT 15.624 7.208 15.696 7.24 ;
  LAYER M1 ;
        RECT 15.644 0.972 15.676 1.044 ;
  LAYER M2 ;
        RECT 15.624 0.992 15.696 1.024 ;
  LAYER M1 ;
        RECT 15.644 1.008 15.676 4.116 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 4.152 ;
  LAYER M2 ;
        RECT 15.624 4.1 15.696 4.132 ;
  LAYER M1 ;
        RECT 3.388 12.732 3.42 12.804 ;
  LAYER M2 ;
        RECT 3.368 12.752 3.44 12.784 ;
  LAYER M2 ;
        RECT 2.86 12.752 3.404 12.784 ;
  LAYER M1 ;
        RECT 2.844 12.732 2.876 12.804 ;
  LAYER M2 ;
        RECT 2.824 12.752 2.896 12.784 ;
  LAYER M1 ;
        RECT 3.388 9.624 3.42 9.696 ;
  LAYER M2 ;
        RECT 3.368 9.644 3.44 9.676 ;
  LAYER M2 ;
        RECT 2.86 9.644 3.404 9.676 ;
  LAYER M1 ;
        RECT 2.844 9.624 2.876 9.696 ;
  LAYER M2 ;
        RECT 2.824 9.644 2.896 9.676 ;
  LAYER M1 ;
        RECT 2.844 22.644 2.876 22.716 ;
  LAYER M2 ;
        RECT 2.824 22.664 2.896 22.696 ;
  LAYER M1 ;
        RECT 2.844 22.428 2.876 22.68 ;
  LAYER M1 ;
        RECT 2.844 9.66 2.876 22.428 ;
  LAYER M1 ;
        RECT 9.98 12.732 10.012 12.804 ;
  LAYER M2 ;
        RECT 9.96 12.752 10.032 12.784 ;
  LAYER M1 ;
        RECT 9.996 12.752 12.748 12.784 ;
  LAYER M1 ;
        RECT 12.732 12.732 12.764 12.804 ;
  LAYER M2 ;
        RECT 12.712 12.752 12.784 12.784 ;
  LAYER M2 ;
        RECT 12.748 12.752 12.812 12.784 ;
  LAYER M1 ;
        RECT 12.796 12.732 12.828 12.804 ;
  LAYER M2 ;
        RECT 12.776 12.752 12.848 12.784 ;
  LAYER M1 ;
        RECT 9.98 15.84 10.012 15.912 ;
  LAYER M2 ;
        RECT 9.96 15.86 10.032 15.892 ;
  LAYER M1 ;
        RECT 9.996 15.86 12.748 15.892 ;
  LAYER M1 ;
        RECT 12.732 15.84 12.764 15.912 ;
  LAYER M2 ;
        RECT 12.712 15.86 12.784 15.892 ;
  LAYER M2 ;
        RECT 12.748 15.86 12.812 15.892 ;
  LAYER M1 ;
        RECT 12.796 15.84 12.828 15.912 ;
  LAYER M2 ;
        RECT 12.776 15.86 12.848 15.892 ;
  LAYER M1 ;
        RECT 12.796 22.644 12.828 22.716 ;
  LAYER M2 ;
        RECT 12.776 22.664 12.848 22.696 ;
  LAYER M1 ;
        RECT 12.796 22.428 12.828 22.68 ;
  LAYER M1 ;
        RECT 12.796 12.936 12.828 22.428 ;
  LAYER M2 ;
        RECT 2.86 22.664 12.812 22.696 ;
  LAYER M1 ;
        RECT 6.684 9.624 6.716 9.696 ;
  LAYER M2 ;
        RECT 6.664 9.644 6.736 9.676 ;
  LAYER M2 ;
        RECT 3.404 9.644 6.7 9.676 ;
  LAYER M1 ;
        RECT 3.388 9.624 3.42 9.696 ;
  LAYER M2 ;
        RECT 3.368 9.644 3.44 9.676 ;
  LAYER M1 ;
        RECT 6.684 15.84 6.716 15.912 ;
  LAYER M2 ;
        RECT 6.664 15.86 6.736 15.892 ;
  LAYER M2 ;
        RECT 6.7 15.86 9.996 15.892 ;
  LAYER M1 ;
        RECT 9.98 15.84 10.012 15.912 ;
  LAYER M2 ;
        RECT 9.96 15.86 10.032 15.892 ;
  LAYER M1 ;
        RECT 3.388 15.84 3.42 15.912 ;
  LAYER M2 ;
        RECT 3.368 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 3.404 15.86 6.316 15.892 ;
  LAYER M1 ;
        RECT 6.3 15.84 6.332 15.912 ;
  LAYER M2 ;
        RECT 6.28 15.86 6.352 15.892 ;
  LAYER M2 ;
        RECT 6.316 15.86 6.38 15.892 ;
  LAYER M1 ;
        RECT 6.364 15.84 6.396 15.912 ;
  LAYER M2 ;
        RECT 6.344 15.86 6.416 15.892 ;
  LAYER M1 ;
        RECT 6.684 6.516 6.716 6.588 ;
  LAYER M2 ;
        RECT 6.664 6.536 6.736 6.568 ;
  LAYER M2 ;
        RECT 6.316 6.536 6.7 6.568 ;
  LAYER M1 ;
        RECT 6.3 6.516 6.332 6.588 ;
  LAYER M2 ;
        RECT 6.28 6.536 6.352 6.568 ;
  LAYER M1 ;
        RECT 6.684 18.948 6.716 19.02 ;
  LAYER M2 ;
        RECT 6.664 18.968 6.736 19 ;
  LAYER M2 ;
        RECT 6.316 18.968 6.7 19 ;
  LAYER M1 ;
        RECT 6.3 18.948 6.332 19.02 ;
  LAYER M2 ;
        RECT 6.28 18.968 6.352 19 ;
  LAYER M1 ;
        RECT 3.388 18.948 3.42 19.02 ;
  LAYER M2 ;
        RECT 3.368 18.968 3.44 19 ;
  LAYER M1 ;
        RECT 3.404 18.968 6.316 19 ;
  LAYER M1 ;
        RECT 6.3 18.948 6.332 19.02 ;
  LAYER M2 ;
        RECT 6.28 18.968 6.352 19 ;
  LAYER M2 ;
        RECT 6.316 18.968 6.38 19 ;
  LAYER M1 ;
        RECT 6.364 18.948 6.396 19.02 ;
  LAYER M2 ;
        RECT 6.344 18.968 6.416 19 ;
  LAYER M1 ;
        RECT 6.364 22.812 6.396 22.884 ;
  LAYER M2 ;
        RECT 6.344 22.832 6.416 22.864 ;
  LAYER M1 ;
        RECT 6.364 22.428 6.396 22.848 ;
  LAYER M1 ;
        RECT 6.364 6.552 6.396 22.428 ;
  LAYER M1 ;
        RECT 9.98 9.624 10.012 9.696 ;
  LAYER M2 ;
        RECT 9.96 9.644 10.032 9.676 ;
  LAYER M2 ;
        RECT 9.612 9.644 9.996 9.676 ;
  LAYER M1 ;
        RECT 9.596 9.624 9.628 9.696 ;
  LAYER M2 ;
        RECT 9.576 9.644 9.648 9.676 ;
  LAYER M1 ;
        RECT 9.98 6.516 10.012 6.588 ;
  LAYER M2 ;
        RECT 9.96 6.536 10.032 6.568 ;
  LAYER M2 ;
        RECT 9.612 6.536 9.996 6.568 ;
  LAYER M1 ;
        RECT 9.596 6.516 9.628 6.588 ;
  LAYER M2 ;
        RECT 9.576 6.536 9.648 6.568 ;
  LAYER M1 ;
        RECT 9.596 22.812 9.628 22.884 ;
  LAYER M2 ;
        RECT 9.576 22.832 9.648 22.864 ;
  LAYER M1 ;
        RECT 9.596 22.428 9.628 22.848 ;
  LAYER M1 ;
        RECT 9.596 6.552 9.628 22.428 ;
  LAYER M2 ;
        RECT 6.38 22.832 9.612 22.864 ;
  LAYER M1 ;
        RECT 3.388 3.408 3.42 3.48 ;
  LAYER M2 ;
        RECT 3.368 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 3.404 3.428 6.476 3.46 ;
  LAYER M1 ;
        RECT 6.46 3.408 6.492 3.48 ;
  LAYER M2 ;
        RECT 6.44 3.428 6.512 3.46 ;
  LAYER M2 ;
        RECT 6.476 3.428 6.54 3.46 ;
  LAYER M1 ;
        RECT 6.524 3.408 6.556 3.48 ;
  LAYER M2 ;
        RECT 6.504 3.428 6.576 3.46 ;
  LAYER M1 ;
        RECT 3.388 6.516 3.42 6.588 ;
  LAYER M2 ;
        RECT 3.368 6.536 3.44 6.568 ;
  LAYER M1 ;
        RECT 3.404 6.536 6.476 6.568 ;
  LAYER M1 ;
        RECT 6.46 6.516 6.492 6.588 ;
  LAYER M2 ;
        RECT 6.44 6.536 6.512 6.568 ;
  LAYER M2 ;
        RECT 6.476 6.536 6.54 6.568 ;
  LAYER M1 ;
        RECT 6.524 6.516 6.556 6.588 ;
  LAYER M2 ;
        RECT 6.504 6.536 6.576 6.568 ;
  LAYER M1 ;
        RECT 3.388 22.056 3.42 22.128 ;
  LAYER M2 ;
        RECT 3.368 22.076 3.44 22.108 ;
  LAYER M1 ;
        RECT 3.404 22.076 6.476 22.108 ;
  LAYER M1 ;
        RECT 6.46 22.056 6.492 22.128 ;
  LAYER M2 ;
        RECT 6.44 22.076 6.512 22.108 ;
  LAYER M2 ;
        RECT 6.476 22.076 6.54 22.108 ;
  LAYER M1 ;
        RECT 6.524 22.056 6.556 22.128 ;
  LAYER M2 ;
        RECT 6.504 22.076 6.576 22.108 ;
  LAYER M1 ;
        RECT 6.684 3.408 6.716 3.48 ;
  LAYER M2 ;
        RECT 6.664 3.428 6.736 3.46 ;
  LAYER M2 ;
        RECT 6.476 3.428 6.7 3.46 ;
  LAYER M1 ;
        RECT 6.46 3.408 6.492 3.48 ;
  LAYER M2 ;
        RECT 6.44 3.428 6.512 3.46 ;
  LAYER M1 ;
        RECT 6.684 12.732 6.716 12.804 ;
  LAYER M2 ;
        RECT 6.664 12.752 6.736 12.784 ;
  LAYER M2 ;
        RECT 6.476 12.752 6.7 12.784 ;
  LAYER M1 ;
        RECT 6.46 12.732 6.492 12.804 ;
  LAYER M2 ;
        RECT 6.44 12.752 6.512 12.784 ;
  LAYER M1 ;
        RECT 6.684 22.056 6.716 22.128 ;
  LAYER M2 ;
        RECT 6.664 22.076 6.736 22.108 ;
  LAYER M2 ;
        RECT 6.476 22.076 6.7 22.108 ;
  LAYER M1 ;
        RECT 6.46 22.056 6.492 22.128 ;
  LAYER M2 ;
        RECT 6.44 22.076 6.512 22.108 ;
  LAYER M1 ;
        RECT 6.46 22.98 6.492 23.052 ;
  LAYER M2 ;
        RECT 6.44 23 6.512 23.032 ;
  LAYER M1 ;
        RECT 6.46 22.428 6.492 23.016 ;
  LAYER M1 ;
        RECT 6.46 3.444 6.492 22.428 ;
  LAYER M1 ;
        RECT 9.98 3.408 10.012 3.48 ;
  LAYER M2 ;
        RECT 9.96 3.428 10.032 3.46 ;
  LAYER M2 ;
        RECT 9.772 3.428 9.996 3.46 ;
  LAYER M1 ;
        RECT 9.756 3.408 9.788 3.48 ;
  LAYER M2 ;
        RECT 9.736 3.428 9.808 3.46 ;
  LAYER M1 ;
        RECT 9.98 18.948 10.012 19.02 ;
  LAYER M2 ;
        RECT 9.96 18.968 10.032 19 ;
  LAYER M2 ;
        RECT 9.772 18.968 9.996 19 ;
  LAYER M1 ;
        RECT 9.756 18.948 9.788 19.02 ;
  LAYER M2 ;
        RECT 9.736 18.968 9.808 19 ;
  LAYER M1 ;
        RECT 9.98 22.056 10.012 22.128 ;
  LAYER M2 ;
        RECT 9.96 22.076 10.032 22.108 ;
  LAYER M2 ;
        RECT 9.772 22.076 9.996 22.108 ;
  LAYER M1 ;
        RECT 9.756 22.056 9.788 22.128 ;
  LAYER M2 ;
        RECT 9.736 22.076 9.808 22.108 ;
  LAYER M1 ;
        RECT 9.756 22.98 9.788 23.052 ;
  LAYER M2 ;
        RECT 9.736 23 9.808 23.032 ;
  LAYER M1 ;
        RECT 9.756 22.428 9.788 23.016 ;
  LAYER M1 ;
        RECT 9.756 3.444 9.788 22.428 ;
  LAYER M2 ;
        RECT 6.476 23 9.772 23.032 ;
  LAYER M1 ;
        RECT 0.092 22.056 0.124 22.128 ;
  LAYER M2 ;
        RECT 0.072 22.076 0.144 22.108 ;
  LAYER M2 ;
        RECT 0.108 22.076 3.404 22.108 ;
  LAYER M1 ;
        RECT 3.388 22.056 3.42 22.128 ;
  LAYER M2 ;
        RECT 3.368 22.076 3.44 22.108 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 18.984 0.124 22.092 ;
  LAYER M1 ;
        RECT 0.092 22.056 0.124 22.128 ;
  LAYER M2 ;
        RECT 0.072 22.076 0.144 22.108 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 15.876 0.124 18.984 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 12.768 0.124 15.876 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 9.66 0.124 12.768 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 0.092 6.552 0.124 9.66 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 3.408 0.124 3.48 ;
  LAYER M2 ;
        RECT 0.072 3.428 0.144 3.46 ;
  LAYER M1 ;
        RECT 0.092 3.444 0.124 6.552 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 13.276 22.056 13.308 22.128 ;
  LAYER M2 ;
        RECT 13.256 22.076 13.328 22.108 ;
  LAYER M2 ;
        RECT 9.996 22.076 13.292 22.108 ;
  LAYER M1 ;
        RECT 9.98 22.056 10.012 22.128 ;
  LAYER M2 ;
        RECT 9.96 22.076 10.032 22.108 ;
  LAYER M1 ;
        RECT 13.276 18.948 13.308 19.02 ;
  LAYER M2 ;
        RECT 13.256 18.968 13.328 19 ;
  LAYER M2 ;
        RECT 9.996 18.968 13.292 19 ;
  LAYER M1 ;
        RECT 9.98 18.948 10.012 19.02 ;
  LAYER M2 ;
        RECT 9.96 18.968 10.032 19 ;
  LAYER M1 ;
        RECT 13.276 15.84 13.308 15.912 ;
  LAYER M2 ;
        RECT 13.256 15.86 13.328 15.892 ;
  LAYER M1 ;
        RECT 13.276 15.876 13.308 18.984 ;
  LAYER M1 ;
        RECT 13.276 18.948 13.308 19.02 ;
  LAYER M2 ;
        RECT 13.256 18.968 13.328 19 ;
  LAYER M1 ;
        RECT 13.276 12.732 13.308 12.804 ;
  LAYER M2 ;
        RECT 13.256 12.752 13.328 12.784 ;
  LAYER M1 ;
        RECT 13.276 12.768 13.308 15.876 ;
  LAYER M1 ;
        RECT 13.276 15.84 13.308 15.912 ;
  LAYER M2 ;
        RECT 13.256 15.86 13.328 15.892 ;
  LAYER M1 ;
        RECT 13.276 9.624 13.308 9.696 ;
  LAYER M2 ;
        RECT 13.256 9.644 13.328 9.676 ;
  LAYER M1 ;
        RECT 13.276 9.66 13.308 12.768 ;
  LAYER M1 ;
        RECT 13.276 12.732 13.308 12.804 ;
  LAYER M2 ;
        RECT 13.256 12.752 13.328 12.784 ;
  LAYER M1 ;
        RECT 13.276 6.516 13.308 6.588 ;
  LAYER M2 ;
        RECT 13.256 6.536 13.328 6.568 ;
  LAYER M1 ;
        RECT 13.276 6.552 13.308 9.66 ;
  LAYER M1 ;
        RECT 13.276 9.624 13.308 9.696 ;
  LAYER M2 ;
        RECT 13.256 9.644 13.328 9.676 ;
  LAYER M1 ;
        RECT 13.276 3.408 13.308 3.48 ;
  LAYER M2 ;
        RECT 13.256 3.428 13.328 3.46 ;
  LAYER M1 ;
        RECT 13.276 3.444 13.308 6.552 ;
  LAYER M1 ;
        RECT 13.276 6.516 13.308 6.588 ;
  LAYER M2 ;
        RECT 13.256 6.536 13.328 6.568 ;
  LAYER M1 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M3 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M2 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M1 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M3 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M2 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M1 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M3 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M2 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M1 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M3 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M2 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M1 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M3 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M2 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M1 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M3 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M2 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M1 ;
        RECT 0.044 19.572 2.54 22.176 ;
  LAYER M3 ;
        RECT 0.044 19.572 2.54 22.176 ;
  LAYER M2 ;
        RECT 0.044 19.572 2.54 22.176 ;
  LAYER M1 ;
        RECT 3.34 0.924 5.836 3.528 ;
  LAYER M3 ;
        RECT 3.34 0.924 5.836 3.528 ;
  LAYER M2 ;
        RECT 3.34 0.924 5.836 3.528 ;
  LAYER M1 ;
        RECT 3.34 4.032 5.836 6.636 ;
  LAYER M3 ;
        RECT 3.34 4.032 5.836 6.636 ;
  LAYER M2 ;
        RECT 3.34 4.032 5.836 6.636 ;
  LAYER M1 ;
        RECT 3.34 7.14 5.836 9.744 ;
  LAYER M3 ;
        RECT 3.34 7.14 5.836 9.744 ;
  LAYER M2 ;
        RECT 3.34 7.14 5.836 9.744 ;
  LAYER M1 ;
        RECT 3.34 10.248 5.836 12.852 ;
  LAYER M3 ;
        RECT 3.34 10.248 5.836 12.852 ;
  LAYER M2 ;
        RECT 3.34 10.248 5.836 12.852 ;
  LAYER M1 ;
        RECT 3.34 13.356 5.836 15.96 ;
  LAYER M3 ;
        RECT 3.34 13.356 5.836 15.96 ;
  LAYER M2 ;
        RECT 3.34 13.356 5.836 15.96 ;
  LAYER M1 ;
        RECT 3.34 16.464 5.836 19.068 ;
  LAYER M3 ;
        RECT 3.34 16.464 5.836 19.068 ;
  LAYER M2 ;
        RECT 3.34 16.464 5.836 19.068 ;
  LAYER M1 ;
        RECT 3.34 19.572 5.836 22.176 ;
  LAYER M3 ;
        RECT 3.34 19.572 5.836 22.176 ;
  LAYER M2 ;
        RECT 3.34 19.572 5.836 22.176 ;
  LAYER M1 ;
        RECT 6.636 0.924 9.132 3.528 ;
  LAYER M3 ;
        RECT 6.636 0.924 9.132 3.528 ;
  LAYER M2 ;
        RECT 6.636 0.924 9.132 3.528 ;
  LAYER M1 ;
        RECT 6.636 4.032 9.132 6.636 ;
  LAYER M3 ;
        RECT 6.636 4.032 9.132 6.636 ;
  LAYER M2 ;
        RECT 6.636 4.032 9.132 6.636 ;
  LAYER M1 ;
        RECT 6.636 7.14 9.132 9.744 ;
  LAYER M3 ;
        RECT 6.636 7.14 9.132 9.744 ;
  LAYER M2 ;
        RECT 6.636 7.14 9.132 9.744 ;
  LAYER M1 ;
        RECT 6.636 10.248 9.132 12.852 ;
  LAYER M3 ;
        RECT 6.636 10.248 9.132 12.852 ;
  LAYER M2 ;
        RECT 6.636 10.248 9.132 12.852 ;
  LAYER M1 ;
        RECT 6.636 13.356 9.132 15.96 ;
  LAYER M3 ;
        RECT 6.636 13.356 9.132 15.96 ;
  LAYER M2 ;
        RECT 6.636 13.356 9.132 15.96 ;
  LAYER M1 ;
        RECT 6.636 16.464 9.132 19.068 ;
  LAYER M3 ;
        RECT 6.636 16.464 9.132 19.068 ;
  LAYER M2 ;
        RECT 6.636 16.464 9.132 19.068 ;
  LAYER M1 ;
        RECT 6.636 19.572 9.132 22.176 ;
  LAYER M3 ;
        RECT 6.636 19.572 9.132 22.176 ;
  LAYER M2 ;
        RECT 6.636 19.572 9.132 22.176 ;
  LAYER M1 ;
        RECT 9.932 0.924 12.428 3.528 ;
  LAYER M3 ;
        RECT 9.932 0.924 12.428 3.528 ;
  LAYER M2 ;
        RECT 9.932 0.924 12.428 3.528 ;
  LAYER M1 ;
        RECT 9.932 4.032 12.428 6.636 ;
  LAYER M3 ;
        RECT 9.932 4.032 12.428 6.636 ;
  LAYER M2 ;
        RECT 9.932 4.032 12.428 6.636 ;
  LAYER M1 ;
        RECT 9.932 7.14 12.428 9.744 ;
  LAYER M3 ;
        RECT 9.932 7.14 12.428 9.744 ;
  LAYER M2 ;
        RECT 9.932 7.14 12.428 9.744 ;
  LAYER M1 ;
        RECT 9.932 10.248 12.428 12.852 ;
  LAYER M3 ;
        RECT 9.932 10.248 12.428 12.852 ;
  LAYER M2 ;
        RECT 9.932 10.248 12.428 12.852 ;
  LAYER M1 ;
        RECT 9.932 13.356 12.428 15.96 ;
  LAYER M3 ;
        RECT 9.932 13.356 12.428 15.96 ;
  LAYER M2 ;
        RECT 9.932 13.356 12.428 15.96 ;
  LAYER M1 ;
        RECT 9.932 16.464 12.428 19.068 ;
  LAYER M3 ;
        RECT 9.932 16.464 12.428 19.068 ;
  LAYER M2 ;
        RECT 9.932 16.464 12.428 19.068 ;
  LAYER M1 ;
        RECT 9.932 19.572 12.428 22.176 ;
  LAYER M3 ;
        RECT 9.932 19.572 12.428 22.176 ;
  LAYER M2 ;
        RECT 9.932 19.572 12.428 22.176 ;
  LAYER M1 ;
        RECT 13.228 0.924 15.724 3.528 ;
  LAYER M3 ;
        RECT 13.228 0.924 15.724 3.528 ;
  LAYER M2 ;
        RECT 13.228 0.924 15.724 3.528 ;
  LAYER M1 ;
        RECT 13.228 4.032 15.724 6.636 ;
  LAYER M3 ;
        RECT 13.228 4.032 15.724 6.636 ;
  LAYER M2 ;
        RECT 13.228 4.032 15.724 6.636 ;
  LAYER M1 ;
        RECT 13.228 7.14 15.724 9.744 ;
  LAYER M3 ;
        RECT 13.228 7.14 15.724 9.744 ;
  LAYER M2 ;
        RECT 13.228 7.14 15.724 9.744 ;
  LAYER M1 ;
        RECT 13.228 10.248 15.724 12.852 ;
  LAYER M3 ;
        RECT 13.228 10.248 15.724 12.852 ;
  LAYER M2 ;
        RECT 13.228 10.248 15.724 12.852 ;
  LAYER M1 ;
        RECT 13.228 13.356 15.724 15.96 ;
  LAYER M3 ;
        RECT 13.228 13.356 15.724 15.96 ;
  LAYER M2 ;
        RECT 13.228 13.356 15.724 15.96 ;
  LAYER M1 ;
        RECT 13.228 16.464 15.724 19.068 ;
  LAYER M3 ;
        RECT 13.228 16.464 15.724 19.068 ;
  LAYER M2 ;
        RECT 13.228 16.464 15.724 19.068 ;
  LAYER M1 ;
        RECT 13.228 19.572 15.724 22.176 ;
  LAYER M3 ;
        RECT 13.228 19.572 15.724 22.176 ;
  LAYER M2 ;
        RECT 13.228 19.572 15.724 22.176 ;
  END 
END Cap_60fF_Cap_60fF
