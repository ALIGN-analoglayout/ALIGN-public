.model n nmos nfin=1 w=1 nf=1 l=1 m=1
.model p pmos nfin=1 w=1 nf=1 l=1 m=1
.model npv nmos nfin=1 w=1 nf=1 l=1 m=1 source=sig drain=sig dv=0
.model ppv pmos nfin=1 w=1 nf=1 l=1 m=1 source=sig drain=sig dv=0
