************************************************************************
* auCdl Netlist:
* 
* Library Name:  OTA_class
* Top Cell Name: single_ended_telescopic
* View Name:     schematic
* Netlisted on:  Sep 11 21:39:36 2019
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: OTA_class
* Cell Name:    single_ended_telescopic
* View Name:    schematic
************************************************************************

.SUBCKT single_ended_telescopic Vbiasn Vbiasp2 Vinn Vinp Voutp
*.PININFO Vbiasn:I Vbiasp2:I Vinn:I Vinp:I Voutp:O
MM3 Voutp Vinp net11 gnd! nmos_rvt w=WA l=LA nfin=nA
MM0 net13 Vinn net11 gnd! nmos_rvt w=WA l=LA nfin=nA
MM4 net11 Vbiasn gnd! gnd! nmos_rvt w=WA l=LA nfin=nA
MM6 net13 Vbiasp2 net016 vdd! pmos_rvt w=WA l=LA nfin=nA
MM5 Voutp Vbiasp2 net014 vdd! pmos_rvt w=WA l=LA nfin=nA
MM1 net014 net13 vdd! vdd! pmos_rvt w=WA l=LA nfin=nA
MM2 net016 net13 vdd! vdd! pmos_rvt w=WA l=LA nfin=nA
.ENDS


.SUBCKT LG_load_biasp_LV Biasn Vbiasp2
*.PININFO Biasn:I Vbiasp2:O
MM0 Vbiasp2 Biasn gnd! gnd! nmos_rvt w=WA l=LA nfin=nA
MM3 net8 Vbiasp2 vdd! vdd! pmos_rvt w=WA l=LA nfin=nA
MM1 Vbiasp2 Vbiasp2 net8 vdd! pmos_rvt w=WA l=LA nfin=nA
.ENDS

.SUBCKT CR1_1 Vbiasn
*.PININFO Vbiasn:O
RRF vdd! Vbiasn res=rK
MM0 Vbiasn Vbiasn gnd! gnd! nmos_rvt w=WA l=LA nfin=nA
.ENDS


xiota LG_Vbiasn LG_Vbiasp2 Vinn Vinp Voutp single_ended_telescopic
xiLG_load_biasp_LV Biasn LG_Vbiasp2 LG_load_biasp_LV
xibCR1_1 Biasn CR1_1
.END