MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 1.2800 BY 1.7640 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
      LAYER M2 ;
        RECT 0.2040 0.9500 0.9160 0.9820 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2780 0.9960 0.3100 ;
      LAYER M2 ;
        RECT 0.2840 1.1180 0.9960 1.1500 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 1.0760 0.2260 ;
      LAYER M2 ;
        RECT 0.3640 1.0340 1.0760 1.0660 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER M3 ;
      RECT 0.5400 0.0900 0.5800 0.1620 ;
    LAYER M3 ;
      RECT 0.6200 0.1740 0.6600 0.2460 ;
    LAYER M3 ;
      RECT 0.4600 0.2580 0.5000 0.3300 ;
    LAYER M1 ;
      RECT 0.3040 0.9300 0.3360 1.5900 ;
    LAYER M1 ;
      RECT 0.9440 0.9300 0.9760 1.5900 ;
    LAYER M1 ;
      RECT 0.2240 0.9300 0.2560 1.5900 ;
    LAYER M1 ;
      RECT 0.8640 0.9300 0.8960 1.5900 ;
    LAYER M1 ;
      RECT 0.3840 0.9300 0.4160 1.5900 ;
    LAYER M1 ;
      RECT 1.0240 0.9300 1.0560 1.5900 ;
    LAYER M3 ;
      RECT 0.5400 0.0900 0.5800 1.0020 ;
    LAYER M3 ;
      RECT 0.6200 0.1740 0.6600 1.0860 ;
    LAYER M3 ;
      RECT 0.4600 0.2580 0.5000 1.1700 ;
  END
END test
