
.subckt SAR_ADC_6b_2GSPS CLK VDD VSS IN IP REFN REFP DOUT<5> DOUT<4> DOUT<3> DOUT<2> DOUT<1> DOUT<0>
I11 QE CLK QIP QSN QSP QD VDD VSS SUB3_CLK1
I18 DN<1> DN<2> DP<1> DP<2> ON OP LAT<1> LAT<2> RDY<1> RDY<2> RS<1> RS<2> VDD VSS SUB2_COMP_DUPLEX
I27 N_Nch<5> N_Nch<4> N_Nch<3> N_Nch<2> N_Nch<1> P_Nch<5> P_Nch<4> P_Nch<3> P_Nch<2> P_Nch<1> IN IP ON OP QSN QSP REFN REFP VDD VSS SUB1_CDAC_6b_diff
I20 DN<1> DN<2> DOUT<5> DOUT<4> DOUT<3> DOUT<2> DOUT<1> DOUT<0> DP<1> DP<2> ENV<2> ENV<3> ENV<4> QIP N_Nch<5> N_Nch<4> N_Nch<3> N_Nch<2> N_Nch<1> P_Nch<5> P_Nch<4> P_Nch<3> P_Nch<2> P_Nch<1> QE RDY<1> RDY<2> VDD VSS SUB5_SEQ_TOP_6b_v2
I10 ENV<2> ENV<3> ENV<4> LAT<1> LAT<2> QD RDY<1> RDY<2> RS<1> RS<2> VDD VSS SUB3_CLK2
.ends SAR_ADC_6b_2GSPS

.subckt SUB3_CLK1 CK_E I QIP QSN QSP QS_DEL_more
I25 net073 VDD VDD VSS VSS QS_DEL BUF_X4
I43 net025 VDD VDD VSS VSS QS_DEL_more INV_X4
I27 QS_DEL_more VDD VDD VSS VSS net062 INV_X4
I108 QS_DEL VDD VDD VSS VSS net062 INV_X6
I100 net37 VDD VDD VSS VSS net35 INV_X6
I121 CK_E VDD VDD VSS VSS net074 BUF_X12
I97 net033 VDD VDD VSS VSS I BUF_X12
C13 VSS QS_DEL Cap_4f
C10 net060 VSS Cap_4f
C11 net061 VSS Cap_4f
C12 net062 VSS Cap_4f
C5 net35 VSS Cap_6f
C15 net37 VSS Cap_6f
C7 net011 VSS Cap_6f
I41 net026 VDD VDD VSS VSS net019 DLY2_X2
I104 net061 VDD VDD VSS VSS net060 DLY2_X2
I102 net062 VDD VDD VSS VSS net061 DLY2_X2
I18 net35 VDD VDD VSS VSS net011 DLY2_X2
I46 net011 VDD VDD VSS VSS net033 DLY2_X2
I109 QSP VDD VDD VSS VSS net076 INV_X16
I111 QSN VDD VDD VSS VSS net057 INV_X16
I120 QIP VDD VDD VSS VSS net025 INV_X8
I110 net076 VDD VDD VSS VSS net057 INV_X8
I112 net057 VDD VDD VSS VSS net073 BUF_X6
I40 net074 VDD VDD VSS VSS net019 net026 NAND2_X4
I101 net069 VDD VDD VSS VSS net37 net033 NAND2_X4
I29 net019 VDD VDD VSS VSS net060 DLY4_X4
I22 net060 VDD VDD VSS VSS net069 DLY4_X4
.ends SUB3_CLK1
