MACRO Switch_NMOS_n12_X3_Y3
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y3 0 0 ;
  SIZE 1.9200 BY 2.5200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.5560 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 1.5560 0.9400 ;
      LAYER M2 ;
        RECT 0.2040 1.7480 1.5560 1.7800 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.7160 0.1840 ;
      LAYER M2 ;
        RECT 0.3640 0.9920 1.7160 1.0240 ;
      LAYER M2 ;
        RECT 0.3640 1.8320 1.7160 1.8640 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 1.6360 0.2680 ;
      LAYER M2 ;
        RECT 0.2840 1.0760 1.6360 1.1080 ;
      LAYER M2 ;
        RECT 0.2840 1.9160 1.6360 1.9480 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.3040 1.7280 0.3360 2.3880 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 1.7280 0.9760 2.3880 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 1.7280 1.6160 2.3880 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 1.7280 0.2560 2.3880 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 0.8640 1.7280 0.8960 2.3880 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.5040 1.7280 1.5360 2.3880 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 1.7280 0.4160 2.3880 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 1.7280 1.0560 2.3880 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 1.7280 1.6960 2.3880 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 1.7480 0.2560 1.7800 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 1.7480 0.8960 1.7800 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.9080 1.5360 0.9400 ;
    LAYER V1 ;
      RECT 1.5040 1.7480 1.5360 1.7800 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9920 0.4160 1.0240 ;
    LAYER V1 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.9920 1.6960 1.0240 ;
    LAYER V1 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 1.0760 0.3360 1.1080 ;
    LAYER V1 ;
      RECT 0.3040 1.9160 0.3360 1.9480 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 1.0760 0.9760 1.1080 ;
    LAYER V1 ;
      RECT 0.9440 1.9160 0.9760 1.9480 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 1.0760 1.6160 1.1080 ;
    LAYER V1 ;
      RECT 1.5840 1.9160 1.6160 1.9480 ;
    LAYER M3 ;
      RECT 0.8600 0.0480 0.9000 1.8000 ;
    LAYER M3 ;
      RECT 0.9400 0.1320 0.9800 1.8840 ;
    LAYER M3 ;
      RECT 0.7800 0.2160 0.8200 1.9680 ;
    LAYER V2 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V2 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V2 ;
      RECT 0.8640 1.7480 0.8960 1.7800 ;
    LAYER V2 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V2 ;
      RECT 0.9440 0.9920 0.9760 1.0240 ;
    LAYER V2 ;
      RECT 0.9440 1.8320 0.9760 1.8640 ;
    LAYER V2 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V2 ;
      RECT 0.7840 1.0760 0.8160 1.1080 ;
    LAYER V2 ;
      RECT 0.7840 1.9160 0.8160 1.9480 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER V0 ;
      RECT 0.2240 1.9160 0.2560 1.9480 ;
    LAYER V0 ;
      RECT 0.2240 2.0420 0.2560 2.0740 ;
    LAYER V0 ;
      RECT 0.2240 2.1680 0.2560 2.2000 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER V0 ;
      RECT 0.8640 1.9160 0.8960 1.9480 ;
    LAYER V0 ;
      RECT 0.8640 2.0420 0.8960 2.0740 ;
    LAYER V0 ;
      RECT 0.8640 2.1680 0.8960 2.2000 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER V0 ;
      RECT 1.5040 1.9160 1.5360 1.9480 ;
    LAYER V0 ;
      RECT 1.5040 2.0420 1.5360 2.0740 ;
    LAYER V0 ;
      RECT 1.5040 2.1680 1.5360 2.2000 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V0 ;
      RECT 0.3840 1.9160 0.4160 1.9480 ;
    LAYER V0 ;
      RECT 0.3840 2.0420 0.4160 2.0740 ;
    LAYER V0 ;
      RECT 0.3840 2.1680 0.4160 2.2000 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER V0 ;
      RECT 1.0240 1.9160 1.0560 1.9480 ;
    LAYER V0 ;
      RECT 1.0240 2.0420 1.0560 2.0740 ;
    LAYER V0 ;
      RECT 1.0240 2.1680 1.0560 2.2000 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER V0 ;
      RECT 1.6640 1.9160 1.6960 1.9480 ;
    LAYER V0 ;
      RECT 1.6640 2.0420 1.6960 2.0740 ;
    LAYER V0 ;
      RECT 1.6640 2.1680 1.6960 2.2000 ;
  END
END Switch_NMOS_n12_X3_Y3
