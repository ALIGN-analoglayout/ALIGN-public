MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 1.5560 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 2.2760 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.3200 1.0560 0.3520 ;
    LAYER V1 ;
      RECT 1.5040 0.3200 1.5360 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
  END
END CMC_PMOS_n12_X2_Y1
