MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 15.2 BY 13.776 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.24 13.32 6.272 13.392 ;
      LAYER M2 ;
        RECT 6.22 13.34 6.292 13.372 ;
      LAYER M1 ;
        RECT 9.152 13.32 9.184 13.392 ;
      LAYER M2 ;
        RECT 9.132 13.34 9.204 13.372 ;
      LAYER M2 ;
        RECT 6.256 13.34 9.168 13.372 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
      LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
      LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
      LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
      LAYER M2 ;
        RECT 6.032 0.404 9.008 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 13.488 3.232 13.56 ;
      LAYER M2 ;
        RECT 3.18 13.508 3.252 13.54 ;
      LAYER M1 ;
        RECT 12.192 13.488 12.224 13.56 ;
      LAYER M2 ;
        RECT 12.172 13.508 12.244 13.54 ;
      LAYER M2 ;
        RECT 3.216 13.508 12.208 13.54 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
      LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 11.984 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M2 ;
        RECT 6.032 7.208 8.784 7.24 ;
  LAYER M1 ;
        RECT 6.016 7.188 6.048 7.26 ;
  LAYER M2 ;
        RECT 5.996 7.208 6.068 7.24 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M1 ;
        RECT 5.792 3.948 5.824 4.116 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M2 ;
        RECT 5.808 3.932 6.032 3.964 ;
  LAYER M1 ;
        RECT 6.016 3.912 6.048 3.984 ;
  LAYER M2 ;
        RECT 5.996 3.932 6.068 3.964 ;
  LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
  LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
  LAYER M1 ;
        RECT 6.016 0.42 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 7.224 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M2 ;
        RECT 9.008 7.208 11.76 7.24 ;
  LAYER M1 ;
        RECT 8.992 7.188 9.024 7.26 ;
  LAYER M2 ;
        RECT 8.972 7.208 9.044 7.24 ;
  LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
  LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
  LAYER M1 ;
        RECT 8.992 0.42 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 7.224 ;
  LAYER M2 ;
        RECT 6.032 0.404 9.008 0.436 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M2 ;
        RECT 3.056 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 3.04 7.188 3.072 7.26 ;
  LAYER M2 ;
        RECT 3.02 7.208 3.092 7.24 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 7.224 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M1 ;
        RECT 11.744 3.948 11.776 4.116 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 11.76 3.932 11.984 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
  LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
  LAYER M1 ;
        RECT 11.968 0.252 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 3.948 ;
  LAYER M2 ;
        RECT 3.056 0.236 11.984 0.268 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M2 ;
        RECT 8.784 4.1 11.76 4.132 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 2.832 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 2.832 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 2.832 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 2.832 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 10.332 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.84 14.752 1.008 ;
  LAYER M1 ;
        RECT 14.72 0.804 14.752 0.876 ;
  LAYER M2 ;
        RECT 14.7 0.824 14.772 0.856 ;
  LAYER M2 ;
        RECT 14.736 0.824 14.96 0.856 ;
  LAYER M1 ;
        RECT 14.944 0.804 14.976 0.876 ;
  LAYER M2 ;
        RECT 14.924 0.824 14.996 0.856 ;
  LAYER M1 ;
        RECT 14.72 4.08 14.752 4.152 ;
  LAYER M2 ;
        RECT 14.7 4.1 14.772 4.132 ;
  LAYER M1 ;
        RECT 14.72 3.948 14.752 4.116 ;
  LAYER M1 ;
        RECT 14.72 3.912 14.752 3.984 ;
  LAYER M2 ;
        RECT 14.7 3.932 14.772 3.964 ;
  LAYER M2 ;
        RECT 14.736 3.932 14.96 3.964 ;
  LAYER M1 ;
        RECT 14.944 3.912 14.976 3.984 ;
  LAYER M2 ;
        RECT 14.924 3.932 14.996 3.964 ;
  LAYER M1 ;
        RECT 14.72 7.188 14.752 7.26 ;
  LAYER M2 ;
        RECT 14.7 7.208 14.772 7.24 ;
  LAYER M1 ;
        RECT 14.72 7.056 14.752 7.224 ;
  LAYER M1 ;
        RECT 14.72 7.02 14.752 7.092 ;
  LAYER M2 ;
        RECT 14.7 7.04 14.772 7.072 ;
  LAYER M2 ;
        RECT 14.736 7.04 14.96 7.072 ;
  LAYER M1 ;
        RECT 14.944 7.02 14.976 7.092 ;
  LAYER M2 ;
        RECT 14.924 7.04 14.996 7.072 ;
  LAYER M1 ;
        RECT 14.72 10.296 14.752 10.368 ;
  LAYER M2 ;
        RECT 14.7 10.316 14.772 10.348 ;
  LAYER M1 ;
        RECT 14.72 10.164 14.752 10.332 ;
  LAYER M1 ;
        RECT 14.72 10.128 14.752 10.2 ;
  LAYER M2 ;
        RECT 14.7 10.148 14.772 10.18 ;
  LAYER M2 ;
        RECT 14.736 10.148 14.96 10.18 ;
  LAYER M1 ;
        RECT 14.944 10.128 14.976 10.2 ;
  LAYER M2 ;
        RECT 14.924 10.148 14.996 10.18 ;
  LAYER M1 ;
        RECT 14.944 0.048 14.976 0.12 ;
  LAYER M2 ;
        RECT 14.924 0.068 14.996 0.1 ;
  LAYER M1 ;
        RECT 14.944 0.084 14.976 0.672 ;
  LAYER M1 ;
        RECT 14.944 0.672 14.976 10.164 ;
  LAYER M2 ;
        RECT 0.08 0.068 14.96 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 2.832 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M2 ;
        RECT 2.832 10.316 5.808 10.348 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M2 ;
        RECT 5.808 10.316 8.784 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M2 ;
        RECT 8.784 10.316 11.76 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M2 ;
        RECT 11.76 0.992 14.736 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M2 ;
        RECT 6.192 9.644 6.416 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M1 ;
        RECT 3.44 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.256 6.568 ;
  LAYER M1 ;
        RECT 6.24 6.516 6.272 6.588 ;
  LAYER M2 ;
        RECT 6.22 6.536 6.292 6.568 ;
  LAYER M1 ;
        RECT 6.24 13.32 6.272 13.392 ;
  LAYER M2 ;
        RECT 6.22 13.34 6.292 13.372 ;
  LAYER M1 ;
        RECT 6.24 13.104 6.272 13.356 ;
  LAYER M1 ;
        RECT 6.24 6.72 6.272 13.104 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M2 ;
        RECT 9.168 9.644 9.392 9.676 ;
  LAYER M1 ;
        RECT 9.152 9.624 9.184 9.696 ;
  LAYER M2 ;
        RECT 9.132 9.644 9.204 9.676 ;
  LAYER M1 ;
        RECT 9.152 13.32 9.184 13.392 ;
  LAYER M2 ;
        RECT 9.132 13.34 9.204 13.372 ;
  LAYER M1 ;
        RECT 9.152 13.104 9.184 13.356 ;
  LAYER M1 ;
        RECT 9.152 9.66 9.184 13.104 ;
  LAYER M2 ;
        RECT 6.256 13.34 9.168 13.372 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.216 9.644 3.44 9.676 ;
  LAYER M1 ;
        RECT 3.2 9.624 3.232 9.696 ;
  LAYER M2 ;
        RECT 3.18 9.644 3.252 9.676 ;
  LAYER M1 ;
        RECT 3.2 13.488 3.232 13.56 ;
  LAYER M2 ;
        RECT 3.18 13.508 3.252 13.54 ;
  LAYER M1 ;
        RECT 3.2 13.104 3.232 13.524 ;
  LAYER M1 ;
        RECT 3.2 9.66 3.232 13.104 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.392 6.536 12.144 6.568 ;
  LAYER M1 ;
        RECT 12.128 6.516 12.16 6.588 ;
  LAYER M2 ;
        RECT 12.108 6.536 12.18 6.568 ;
  LAYER M2 ;
        RECT 12.144 6.536 12.208 6.568 ;
  LAYER M1 ;
        RECT 12.192 6.516 12.224 6.588 ;
  LAYER M2 ;
        RECT 12.172 6.536 12.244 6.568 ;
  LAYER M1 ;
        RECT 12.192 13.488 12.224 13.56 ;
  LAYER M2 ;
        RECT 12.172 13.508 12.244 13.54 ;
  LAYER M1 ;
        RECT 12.192 13.104 12.224 13.524 ;
  LAYER M1 ;
        RECT 12.192 6.72 12.224 13.104 ;
  LAYER M2 ;
        RECT 3.216 13.508 12.208 13.54 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.416 6.536 9.392 6.568 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.224 13.656 0.256 13.728 ;
  LAYER M2 ;
        RECT 0.204 13.676 0.276 13.708 ;
  LAYER M1 ;
        RECT 0.224 13.104 0.256 13.692 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 13.104 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M1 ;
        RECT 12.368 3.428 15.12 3.46 ;
  LAYER M1 ;
        RECT 15.104 3.408 15.136 3.48 ;
  LAYER M2 ;
        RECT 15.084 3.428 15.156 3.46 ;
  LAYER M2 ;
        RECT 15.12 3.428 15.184 3.46 ;
  LAYER M1 ;
        RECT 15.168 3.408 15.2 3.48 ;
  LAYER M2 ;
        RECT 15.148 3.428 15.22 3.46 ;
  LAYER M1 ;
        RECT 12.352 6.516 12.384 6.588 ;
  LAYER M2 ;
        RECT 12.332 6.536 12.404 6.568 ;
  LAYER M1 ;
        RECT 12.368 6.536 15.12 6.568 ;
  LAYER M1 ;
        RECT 15.104 6.516 15.136 6.588 ;
  LAYER M2 ;
        RECT 15.084 6.536 15.156 6.568 ;
  LAYER M2 ;
        RECT 15.12 6.536 15.184 6.568 ;
  LAYER M1 ;
        RECT 15.168 6.516 15.2 6.588 ;
  LAYER M2 ;
        RECT 15.148 6.536 15.22 6.568 ;
  LAYER M1 ;
        RECT 12.352 9.624 12.384 9.696 ;
  LAYER M2 ;
        RECT 12.332 9.644 12.404 9.676 ;
  LAYER M1 ;
        RECT 12.368 9.644 15.12 9.676 ;
  LAYER M1 ;
        RECT 15.104 9.624 15.136 9.696 ;
  LAYER M2 ;
        RECT 15.084 9.644 15.156 9.676 ;
  LAYER M2 ;
        RECT 15.12 9.644 15.184 9.676 ;
  LAYER M1 ;
        RECT 15.168 9.624 15.2 9.696 ;
  LAYER M2 ;
        RECT 15.148 9.644 15.22 9.676 ;
  LAYER M1 ;
        RECT 12.352 12.732 12.384 12.804 ;
  LAYER M2 ;
        RECT 12.332 12.752 12.404 12.784 ;
  LAYER M1 ;
        RECT 12.368 12.752 15.12 12.784 ;
  LAYER M1 ;
        RECT 15.104 12.732 15.136 12.804 ;
  LAYER M2 ;
        RECT 15.084 12.752 15.156 12.784 ;
  LAYER M2 ;
        RECT 15.12 12.752 15.184 12.784 ;
  LAYER M1 ;
        RECT 15.168 12.732 15.2 12.804 ;
  LAYER M2 ;
        RECT 15.148 12.752 15.22 12.784 ;
  LAYER M1 ;
        RECT 15.168 13.656 15.2 13.728 ;
  LAYER M2 ;
        RECT 15.148 13.676 15.22 13.708 ;
  LAYER M1 ;
        RECT 15.168 13.104 15.2 13.692 ;
  LAYER M1 ;
        RECT 15.168 3.612 15.2 13.104 ;
  LAYER M2 ;
        RECT 0.24 13.676 15.184 13.708 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 0.464 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 3.44 12.752 6.416 12.784 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M2 ;
        RECT 6.416 12.752 9.392 12.784 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M2 ;
        RECT 9.392 3.428 12.368 3.46 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M3 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M3 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M3 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M3 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M3 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M3 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M3 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M3 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M3 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M3 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M3 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M3 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M3 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M3 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M3 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M3 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M2 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M1 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M3 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M2 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M1 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M3 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M2 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M1 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M3 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M2 ;
        RECT 12.304 10.248 14.8 12.852 ;
  END 
END Cap_30fF_Cap_30fF
