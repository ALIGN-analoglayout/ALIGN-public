MACRO Switch_PMOS_B_nfin5_nf6_m1_n12_X3_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_B_nfin5_nf6_m1_n12_X3_Y1_SLVT 0 0 ;
  SIZE 0.9600 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.7560 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.6760 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.6760 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.6760 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
  END
END Switch_PMOS_B_nfin5_nf6_m1_n12_X3_Y1_SLVT
MACRO Switch_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_NMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT
MACRO Res_958p82
  ORIGIN 0 0 ;
  FOREIGN Res_958p82 0 0 ;
  SIZE 0.9600 BY 3.2760 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.3560 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.5400 3.1760 0.8680 3.2080 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 3.2280 ;
    LAYER M1 ;
      RECT 0.3040 3.1760 0.4000 3.2080 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 3.2280 ;
    LAYER M1 ;
      RECT 0.3680 0.0680 0.4640 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 3.2280 ;
    LAYER M1 ;
      RECT 0.4320 3.1760 0.5280 3.2080 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 3.2280 ;
    LAYER M1 ;
      RECT 0.4960 0.0680 0.5920 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 3.2280 ;
    LAYER V1 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.5600 3.1760 0.5920 3.2080 ;
  END
END Res_958p82
MACRO DP_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN DP_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9920 0.5160 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END DP_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
MACRO Dcap_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Dcap_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 0.2880 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.5160 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 0.1520 0.1760 0.1840 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Dcap_NMOS_B_nfin4_nf6_m1_n12_X2_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf8_m1_n12_X2_Y2_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf8_m1_n12_X2_Y2_SLVT 0 0 ;
  SIZE 0.8000 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.8880 0.3400 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 1.2440 0.5960 1.2760 ;
    LAYER M2 ;
      RECT 0.1240 2.6720 0.5160 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.3280 0.5160 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.5160 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.2440 0.1760 1.2760 ;
    LAYER V2 ;
      RECT 0.1440 2.6720 0.1760 2.7040 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER V2 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
  END
END Switch_PMOS_nfin5_nf8_m1_n12_X2_Y2_SLVT
MACRO CMC_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END CMC_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO CMC_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END CMC_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf5_m1_n12_X3_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf5_m1_n12_X3_Y1_SLVT 0 0 ;
  SIZE 0.9600 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.6760 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.6760 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 1.4960 0.6760 1.5280 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V2 ;
      RECT 0.2240 1.4960 0.2560 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
  END
END Switch_PMOS_nfin5_nf5_m1_n12_X3_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf3_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf3_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_nfin4_nf3_m1_n12_X1_Y1_SLVT
MACRO CCP_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 1.0440 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER M2 ;
      RECT 0.1240 0.9920 0.3560 1.0240 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.5160 0.2680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V2 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END CCP_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
MACRO Cap_12f
  ORIGIN 0 0 ;
  FOREIGN Cap_12f 0 0 ;
  SIZE 2.4000 BY 2.4360 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 -0.0160 2.4360 0.0160 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 2.4200 2.4360 2.4520 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
  END
END Cap_12f
MACRO CCP_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 1.0440 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER M2 ;
      RECT 0.1240 0.9920 0.3560 1.0240 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.5160 0.2680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V2 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END CCP_NMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_PMOS_nfin4_nf4_m1_n12_X2_Y1_SLVT
MACRO Switch_PMOS_B_nfin5_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_B_nfin5_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 1.4960 0.3560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_B_nfin5_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 1.4960 0.3560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf2_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf2_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_nfin4_nf2_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf2_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf2_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_nfin5_nf2_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 1.4960 0.3560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_NMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 1.4960 0.3560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_B_nfin4_nf2_m1_n12_X1_Y1_SLVT
MACRO CMC_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT 0 0 ;
  SIZE 1.4400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 1.1560 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 1.1560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 1.4960 1.1560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
  END
END CMC_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT
MACRO DP_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 1.1200 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.8360 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 0.6760 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.8360 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.9920 0.6760 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.8360 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9920 0.6560 1.0240 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
  END
END DP_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
MACRO Dummy_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Dummy_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.9080 0.3560 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 0.9080 0.1760 0.9400 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Dummy_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf6_m1_n12_X3_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf6_m1_n12_X3_Y1_SLVT 0 0 ;
  SIZE 0.9600 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.6760 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.6760 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 1.4960 0.6760 1.5280 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V2 ;
      RECT 0.2240 1.4960 0.2560 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
  END
END Switch_PMOS_nfin5_nf6_m1_n12_X3_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_nfin5_nf1_m1_n12_X1_Y1_SLVT
MACRO Res_1917p65
  ORIGIN 0 0 ;
  FOREIGN Res_1917p65 0 0 ;
  SIZE 1.2800 BY 3.2760 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 0.3560 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7960 3.1760 1.1240 3.2080 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 3.2280 ;
    LAYER M1 ;
      RECT 0.3040 3.1760 0.4000 3.2080 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 3.2280 ;
    LAYER M1 ;
      RECT 0.3680 0.0680 0.4640 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 3.2280 ;
    LAYER M1 ;
      RECT 0.4320 3.1760 0.5280 3.2080 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 3.2280 ;
    LAYER M1 ;
      RECT 0.4960 0.0680 0.5920 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 3.2280 ;
    LAYER M1 ;
      RECT 0.5600 3.1760 0.6560 3.2080 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 3.2280 ;
    LAYER M1 ;
      RECT 0.6240 0.0680 0.7200 0.1000 ;
    LAYER M1 ;
      RECT 0.6880 0.0480 0.7200 3.2280 ;
    LAYER M1 ;
      RECT 0.6880 3.1760 0.7840 3.2080 ;
    LAYER M1 ;
      RECT 0.7520 0.0480 0.7840 3.2280 ;
    LAYER M1 ;
      RECT 0.7520 0.0680 0.8480 0.1000 ;
    LAYER M1 ;
      RECT 0.8160 0.0480 0.8480 3.2280 ;
    LAYER V1 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.8160 3.1760 0.8480 3.2080 ;
  END
END Res_1917p65
MACRO Switch_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
MACRO Switch_NMOS_B_nfin4_nf11_m1_n12_X2_Y2_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_B_nfin4_nf11_m1_n12_X2_Y2_SLVT 0 0 ;
  SIZE 0.8000 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.2960 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.8880 0.3400 2.1360 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 2.6720 0.5160 2.7040 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.2240 0.3360 1.9680 ;
    LAYER M1 ;
      RECT 0.3040 2.0640 0.3360 2.3040 ;
    LAYER M1 ;
      RECT 0.3040 2.5680 0.3360 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.2240 0.4960 1.9680 ;
    LAYER M1 ;
      RECT 0.4640 2.0640 0.4960 2.3040 ;
    LAYER M1 ;
      RECT 0.4640 2.5680 0.4960 2.8080 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 1.2440 0.5960 1.2760 ;
    LAYER M2 ;
      RECT 0.2040 1.3280 0.5160 1.3600 ;
    LAYER M2 ;
      RECT 0.2840 2.0840 0.5160 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.3280 0.3360 1.3600 ;
    LAYER V1 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V1 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V1 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V1 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.2440 0.1760 1.2760 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER V2 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.5800 0.3360 1.6120 ;
    LAYER V0 ;
      RECT 0.3040 1.7060 0.3360 1.7380 ;
    LAYER V0 ;
      RECT 0.3040 1.8320 0.3360 1.8640 ;
    LAYER V0 ;
      RECT 0.3040 2.0840 0.3360 2.1160 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.3040 2.6720 0.3360 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.5800 0.4960 1.6120 ;
    LAYER V0 ;
      RECT 0.4640 1.7060 0.4960 1.7380 ;
    LAYER V0 ;
      RECT 0.4640 1.8320 0.4960 1.8640 ;
    LAYER V0 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.4640 2.6720 0.4960 2.7040 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
  END
END Switch_NMOS_B_nfin4_nf11_m1_n12_X2_Y2_SLVT
MACRO Switch_PMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0600 0.0480 0.1000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.0440 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.0440 1.4960 0.3560 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.0640 0.0680 0.0960 0.1000 ;
    LAYER V2 ;
      RECT 0.0640 1.4960 0.0960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf5_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf5_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_NMOS_nfin4_nf5_m1_n12_X2_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf3_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf3_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_PMOS_nfin5_nf3_m1_n12_X2_Y1_SLVT
MACRO CCP_S_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CCP_S_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 2.5600 BY 1.8480 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.1520 1.7160 0.1840 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2600 0.2160 1.3000 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3400 0.3000 1.3800 1.0440 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 2.2760 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.3920 1.6160 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.3920 2.2560 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M2 ;
      RECT 0.9240 0.9080 1.6360 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 2.2760 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.9920 2.2760 1.0240 ;
    LAYER M2 ;
      RECT 0.9240 0.3200 1.6360 0.3520 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.1520 0.8960 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.5040 0.1520 1.5360 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.3200 1.6160 0.3520 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 2.2240 0.2360 2.2560 0.2680 ;
    LAYER V1 ;
      RECT 2.2240 0.9920 2.2560 1.0240 ;
    LAYER V1 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 1.2640 0.2360 1.2960 0.2680 ;
    LAYER V2 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V2 ;
      RECT 1.3440 0.3200 1.3760 0.3520 ;
    LAYER V2 ;
      RECT 1.3440 0.9920 1.3760 1.0240 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
  END
END CCP_S_NMOS_B_nfin4_nf4_m1_n12_X2_Y1_SLVT
MACRO DP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN DP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9920 0.5160 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END DP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf6_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf6_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_NMOS_nfin4_nf6_m1_n12_X2_Y1_SLVT
MACRO CCP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 1.0440 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER M2 ;
      RECT 0.1240 0.9920 0.3560 1.0240 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.5160 0.2680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V2 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V2 ;
      RECT 0.3040 0.9920 0.3360 1.0240 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END CCP_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 1.4960 0.3560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Switch_PMOS_B_nfin4_nf1_m1_n12_X1_Y1_SLVT
MACRO Switch_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT 0 0 ;
  SIZE 0.9600 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.6760 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.6760 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 1.4960 0.6760 1.5280 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V2 ;
      RECT 0.2240 1.4960 0.2560 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
  END
END Switch_NMOS_nfin4_nf8_m1_n12_X3_Y1_SLVT
MACRO Switch_PMOS_nfin5_nf4_m1_n12_X2_Y1_SLVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin5_nf4_m1_n12_X2_Y1_SLVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.5160 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END Switch_PMOS_nfin5_nf4_m1_n12_X2_Y1_SLVT
