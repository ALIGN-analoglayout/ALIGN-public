MACRO SCM_PMOS_nfin5_n12_X1_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN SCM_PMOS_nfin5_n12_X1_Y1_RVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END SCM_PMOS_nfin5_n12_X1_Y1_RVT
MACRO SCM_NMOS_nfin5_n12_X1_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin5_n12_X1_Y1_RVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END SCM_NMOS_nfin5_n12_X1_Y1_RVT
MACRO DP_NMOS_B_nfin5_n12_X1_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin5_n12_X1_Y1_RVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.5960 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.9080 0.3560 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9920 0.5160 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.5160 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END DP_NMOS_B_nfin5_n12_X1_Y1_RVT
