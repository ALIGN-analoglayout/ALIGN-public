MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 10.32 BY 35.532 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.808 35.076 3.84 35.148 ;
      LAYER M2 ;
        RECT 3.788 35.096 3.86 35.128 ;
      LAYER M1 ;
        RECT 7.104 35.076 7.136 35.148 ;
      LAYER M2 ;
        RECT 7.084 35.096 7.156 35.128 ;
      LAYER M2 ;
        RECT 3.824 35.096 7.12 35.128 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
      LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
      LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
      LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
      LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.968 35.244 4 35.316 ;
      LAYER M2 ;
        RECT 3.948 35.264 4.02 35.296 ;
      LAYER M1 ;
        RECT 7.264 35.244 7.296 35.316 ;
      LAYER M2 ;
        RECT 7.244 35.264 7.316 35.296 ;
      LAYER M2 ;
        RECT 3.984 35.264 7.28 35.296 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
      LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
      LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
      LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
      LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.496 16.512 6.528 16.584 ;
  LAYER M2 ;
        RECT 6.476 16.532 6.548 16.564 ;
  LAYER M2 ;
        RECT 3.376 16.532 6.512 16.564 ;
  LAYER M1 ;
        RECT 3.36 16.512 3.392 16.584 ;
  LAYER M2 ;
        RECT 3.34 16.532 3.412 16.564 ;
  LAYER M1 ;
        RECT 6.496 4.08 6.528 4.152 ;
  LAYER M2 ;
        RECT 6.476 4.1 6.548 4.132 ;
  LAYER M2 ;
        RECT 3.376 4.1 6.512 4.132 ;
  LAYER M1 ;
        RECT 3.36 4.08 3.392 4.152 ;
  LAYER M2 ;
        RECT 3.34 4.1 3.412 4.132 ;
  LAYER M1 ;
        RECT 6.496 28.944 6.528 29.016 ;
  LAYER M2 ;
        RECT 6.476 28.964 6.548 28.996 ;
  LAYER M2 ;
        RECT 3.376 28.964 6.512 28.996 ;
  LAYER M1 ;
        RECT 3.36 28.944 3.392 29.016 ;
  LAYER M2 ;
        RECT 3.34 28.964 3.412 28.996 ;
  LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
  LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
  LAYER M1 ;
        RECT 3.36 0.42 3.392 0.672 ;
  LAYER M1 ;
        RECT 3.36 0.672 3.392 28.98 ;
  LAYER M1 ;
        RECT 6.496 16.512 6.528 16.584 ;
  LAYER M2 ;
        RECT 6.476 16.532 6.548 16.564 ;
  LAYER M1 ;
        RECT 6.496 16.38 6.528 16.548 ;
  LAYER M1 ;
        RECT 6.496 16.344 6.528 16.416 ;
  LAYER M2 ;
        RECT 6.476 16.364 6.548 16.396 ;
  LAYER M2 ;
        RECT 6.512 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 16.416 ;
  LAYER M2 ;
        RECT 6.636 16.364 6.708 16.396 ;
  LAYER M1 ;
        RECT 6.496 4.08 6.528 4.152 ;
  LAYER M2 ;
        RECT 6.476 4.1 6.548 4.132 ;
  LAYER M1 ;
        RECT 6.496 3.948 6.528 4.116 ;
  LAYER M1 ;
        RECT 6.496 3.912 6.528 3.984 ;
  LAYER M2 ;
        RECT 6.476 3.932 6.548 3.964 ;
  LAYER M2 ;
        RECT 6.512 3.932 6.672 3.964 ;
  LAYER M1 ;
        RECT 6.656 3.912 6.688 3.984 ;
  LAYER M2 ;
        RECT 6.636 3.932 6.708 3.964 ;
  LAYER M1 ;
        RECT 6.496 28.944 6.528 29.016 ;
  LAYER M2 ;
        RECT 6.476 28.964 6.548 28.996 ;
  LAYER M1 ;
        RECT 6.496 28.812 6.528 28.98 ;
  LAYER M1 ;
        RECT 6.496 28.776 6.528 28.848 ;
  LAYER M2 ;
        RECT 6.476 28.796 6.548 28.828 ;
  LAYER M2 ;
        RECT 6.512 28.796 6.672 28.828 ;
  LAYER M1 ;
        RECT 6.656 28.776 6.688 28.848 ;
  LAYER M2 ;
        RECT 6.636 28.796 6.708 28.828 ;
  LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
  LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
  LAYER M1 ;
        RECT 6.656 0.42 6.688 0.672 ;
  LAYER M1 ;
        RECT 6.656 0.672 6.688 28.812 ;
  LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
  LAYER M1 ;
        RECT 6.496 13.404 6.528 13.476 ;
  LAYER M2 ;
        RECT 6.476 13.424 6.548 13.456 ;
  LAYER M2 ;
        RECT 3.536 13.424 6.512 13.456 ;
  LAYER M1 ;
        RECT 3.52 13.404 3.552 13.476 ;
  LAYER M2 ;
        RECT 3.5 13.424 3.572 13.456 ;
  LAYER M1 ;
        RECT 6.496 19.62 6.528 19.692 ;
  LAYER M2 ;
        RECT 6.476 19.64 6.548 19.672 ;
  LAYER M2 ;
        RECT 3.536 19.64 6.512 19.672 ;
  LAYER M1 ;
        RECT 3.52 19.62 3.552 19.692 ;
  LAYER M2 ;
        RECT 3.5 19.64 3.572 19.672 ;
  LAYER M1 ;
        RECT 6.496 10.296 6.528 10.368 ;
  LAYER M2 ;
        RECT 6.476 10.316 6.548 10.348 ;
  LAYER M2 ;
        RECT 3.536 10.316 6.512 10.348 ;
  LAYER M1 ;
        RECT 3.52 10.296 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.5 10.316 3.572 10.348 ;
  LAYER M1 ;
        RECT 6.496 22.728 6.528 22.8 ;
  LAYER M2 ;
        RECT 6.476 22.748 6.548 22.78 ;
  LAYER M2 ;
        RECT 3.536 22.748 6.512 22.78 ;
  LAYER M1 ;
        RECT 3.52 22.728 3.552 22.8 ;
  LAYER M2 ;
        RECT 3.5 22.748 3.572 22.78 ;
  LAYER M1 ;
        RECT 6.496 7.188 6.528 7.26 ;
  LAYER M2 ;
        RECT 6.476 7.208 6.548 7.24 ;
  LAYER M2 ;
        RECT 3.536 7.208 6.512 7.24 ;
  LAYER M1 ;
        RECT 3.52 7.188 3.552 7.26 ;
  LAYER M2 ;
        RECT 3.5 7.208 3.572 7.24 ;
  LAYER M1 ;
        RECT 6.496 25.836 6.528 25.908 ;
  LAYER M2 ;
        RECT 6.476 25.856 6.548 25.888 ;
  LAYER M2 ;
        RECT 3.536 25.856 6.512 25.888 ;
  LAYER M1 ;
        RECT 3.52 25.836 3.552 25.908 ;
  LAYER M2 ;
        RECT 3.5 25.856 3.572 25.888 ;
  LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
  LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
  LAYER M1 ;
        RECT 3.52 0.252 3.552 0.672 ;
  LAYER M1 ;
        RECT 3.52 0.672 3.552 25.872 ;
  LAYER M1 ;
        RECT 6.496 13.404 6.528 13.476 ;
  LAYER M2 ;
        RECT 6.476 13.424 6.548 13.456 ;
  LAYER M1 ;
        RECT 6.496 13.272 6.528 13.44 ;
  LAYER M1 ;
        RECT 6.496 13.236 6.528 13.308 ;
  LAYER M2 ;
        RECT 6.476 13.256 6.548 13.288 ;
  LAYER M2 ;
        RECT 6.512 13.256 6.832 13.288 ;
  LAYER M1 ;
        RECT 6.816 13.236 6.848 13.308 ;
  LAYER M2 ;
        RECT 6.796 13.256 6.868 13.288 ;
  LAYER M1 ;
        RECT 6.496 19.62 6.528 19.692 ;
  LAYER M2 ;
        RECT 6.476 19.64 6.548 19.672 ;
  LAYER M1 ;
        RECT 6.496 19.488 6.528 19.656 ;
  LAYER M1 ;
        RECT 6.496 19.452 6.528 19.524 ;
  LAYER M2 ;
        RECT 6.476 19.472 6.548 19.504 ;
  LAYER M2 ;
        RECT 6.512 19.472 6.832 19.504 ;
  LAYER M1 ;
        RECT 6.816 19.452 6.848 19.524 ;
  LAYER M2 ;
        RECT 6.796 19.472 6.868 19.504 ;
  LAYER M1 ;
        RECT 6.496 10.296 6.528 10.368 ;
  LAYER M2 ;
        RECT 6.476 10.316 6.548 10.348 ;
  LAYER M1 ;
        RECT 6.496 10.164 6.528 10.332 ;
  LAYER M1 ;
        RECT 6.496 10.128 6.528 10.2 ;
  LAYER M2 ;
        RECT 6.476 10.148 6.548 10.18 ;
  LAYER M2 ;
        RECT 6.512 10.148 6.832 10.18 ;
  LAYER M1 ;
        RECT 6.816 10.128 6.848 10.2 ;
  LAYER M2 ;
        RECT 6.796 10.148 6.868 10.18 ;
  LAYER M1 ;
        RECT 6.496 22.728 6.528 22.8 ;
  LAYER M2 ;
        RECT 6.476 22.748 6.548 22.78 ;
  LAYER M1 ;
        RECT 6.496 22.596 6.528 22.764 ;
  LAYER M1 ;
        RECT 6.496 22.56 6.528 22.632 ;
  LAYER M2 ;
        RECT 6.476 22.58 6.548 22.612 ;
  LAYER M2 ;
        RECT 6.512 22.58 6.832 22.612 ;
  LAYER M1 ;
        RECT 6.816 22.56 6.848 22.632 ;
  LAYER M2 ;
        RECT 6.796 22.58 6.868 22.612 ;
  LAYER M1 ;
        RECT 6.496 7.188 6.528 7.26 ;
  LAYER M2 ;
        RECT 6.476 7.208 6.548 7.24 ;
  LAYER M1 ;
        RECT 6.496 7.056 6.528 7.224 ;
  LAYER M1 ;
        RECT 6.496 7.02 6.528 7.092 ;
  LAYER M2 ;
        RECT 6.476 7.04 6.548 7.072 ;
  LAYER M2 ;
        RECT 6.512 7.04 6.832 7.072 ;
  LAYER M1 ;
        RECT 6.816 7.02 6.848 7.092 ;
  LAYER M2 ;
        RECT 6.796 7.04 6.868 7.072 ;
  LAYER M1 ;
        RECT 6.496 25.836 6.528 25.908 ;
  LAYER M2 ;
        RECT 6.476 25.856 6.548 25.888 ;
  LAYER M1 ;
        RECT 6.496 25.704 6.528 25.872 ;
  LAYER M1 ;
        RECT 6.496 25.668 6.528 25.74 ;
  LAYER M2 ;
        RECT 6.476 25.688 6.548 25.72 ;
  LAYER M2 ;
        RECT 6.512 25.688 6.832 25.72 ;
  LAYER M1 ;
        RECT 6.816 25.668 6.848 25.74 ;
  LAYER M2 ;
        RECT 6.796 25.688 6.868 25.72 ;
  LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
  LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
  LAYER M1 ;
        RECT 6.816 0.252 6.848 0.672 ;
  LAYER M1 ;
        RECT 6.816 0.672 6.848 25.704 ;
  LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
  LAYER M1 ;
        RECT 3.2 0.972 3.232 1.044 ;
  LAYER M2 ;
        RECT 3.18 0.992 3.252 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 3.216 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 3.2 4.08 3.232 4.152 ;
  LAYER M2 ;
        RECT 3.18 4.1 3.252 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 3.216 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 3.2 7.188 3.232 7.26 ;
  LAYER M2 ;
        RECT 3.18 7.208 3.252 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 3.216 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 3.2 10.296 3.232 10.368 ;
  LAYER M2 ;
        RECT 3.18 10.316 3.252 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 3.216 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 3.2 13.404 3.232 13.476 ;
  LAYER M2 ;
        RECT 3.18 13.424 3.252 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 3.216 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 3.2 16.512 3.232 16.584 ;
  LAYER M2 ;
        RECT 3.18 16.532 3.252 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 3.216 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 3.2 19.62 3.232 19.692 ;
  LAYER M2 ;
        RECT 3.18 19.64 3.252 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 3.216 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 3.2 22.728 3.232 22.8 ;
  LAYER M2 ;
        RECT 3.18 22.748 3.252 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 3.216 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 3.2 25.836 3.232 25.908 ;
  LAYER M2 ;
        RECT 3.18 25.856 3.252 25.888 ;
  LAYER M2 ;
        RECT 0.08 25.856 3.216 25.888 ;
  LAYER M1 ;
        RECT 0.064 25.836 0.096 25.908 ;
  LAYER M2 ;
        RECT 0.044 25.856 0.116 25.888 ;
  LAYER M1 ;
        RECT 3.2 28.944 3.232 29.016 ;
  LAYER M2 ;
        RECT 3.18 28.964 3.252 28.996 ;
  LAYER M2 ;
        RECT 0.08 28.964 3.216 28.996 ;
  LAYER M1 ;
        RECT 0.064 28.944 0.096 29.016 ;
  LAYER M2 ;
        RECT 0.044 28.964 0.116 28.996 ;
  LAYER M1 ;
        RECT 3.2 32.052 3.232 32.124 ;
  LAYER M2 ;
        RECT 3.18 32.072 3.252 32.104 ;
  LAYER M2 ;
        RECT 0.08 32.072 3.216 32.104 ;
  LAYER M1 ;
        RECT 0.064 32.052 0.096 32.124 ;
  LAYER M2 ;
        RECT 0.044 32.072 0.116 32.104 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 32.088 ;
  LAYER M1 ;
        RECT 9.792 0.972 9.824 1.044 ;
  LAYER M2 ;
        RECT 9.772 0.992 9.844 1.024 ;
  LAYER M1 ;
        RECT 9.792 0.84 9.824 1.008 ;
  LAYER M1 ;
        RECT 9.792 0.804 9.824 0.876 ;
  LAYER M2 ;
        RECT 9.772 0.824 9.844 0.856 ;
  LAYER M2 ;
        RECT 9.808 0.824 9.968 0.856 ;
  LAYER M1 ;
        RECT 9.952 0.804 9.984 0.876 ;
  LAYER M2 ;
        RECT 9.932 0.824 10.004 0.856 ;
  LAYER M1 ;
        RECT 9.792 4.08 9.824 4.152 ;
  LAYER M2 ;
        RECT 9.772 4.1 9.844 4.132 ;
  LAYER M1 ;
        RECT 9.792 3.948 9.824 4.116 ;
  LAYER M1 ;
        RECT 9.792 3.912 9.824 3.984 ;
  LAYER M2 ;
        RECT 9.772 3.932 9.844 3.964 ;
  LAYER M2 ;
        RECT 9.808 3.932 9.968 3.964 ;
  LAYER M1 ;
        RECT 9.952 3.912 9.984 3.984 ;
  LAYER M2 ;
        RECT 9.932 3.932 10.004 3.964 ;
  LAYER M1 ;
        RECT 9.792 7.188 9.824 7.26 ;
  LAYER M2 ;
        RECT 9.772 7.208 9.844 7.24 ;
  LAYER M1 ;
        RECT 9.792 7.056 9.824 7.224 ;
  LAYER M1 ;
        RECT 9.792 7.02 9.824 7.092 ;
  LAYER M2 ;
        RECT 9.772 7.04 9.844 7.072 ;
  LAYER M2 ;
        RECT 9.808 7.04 9.968 7.072 ;
  LAYER M1 ;
        RECT 9.952 7.02 9.984 7.092 ;
  LAYER M2 ;
        RECT 9.932 7.04 10.004 7.072 ;
  LAYER M1 ;
        RECT 9.792 10.296 9.824 10.368 ;
  LAYER M2 ;
        RECT 9.772 10.316 9.844 10.348 ;
  LAYER M1 ;
        RECT 9.792 10.164 9.824 10.332 ;
  LAYER M1 ;
        RECT 9.792 10.128 9.824 10.2 ;
  LAYER M2 ;
        RECT 9.772 10.148 9.844 10.18 ;
  LAYER M2 ;
        RECT 9.808 10.148 9.968 10.18 ;
  LAYER M1 ;
        RECT 9.952 10.128 9.984 10.2 ;
  LAYER M2 ;
        RECT 9.932 10.148 10.004 10.18 ;
  LAYER M1 ;
        RECT 9.792 13.404 9.824 13.476 ;
  LAYER M2 ;
        RECT 9.772 13.424 9.844 13.456 ;
  LAYER M1 ;
        RECT 9.792 13.272 9.824 13.44 ;
  LAYER M1 ;
        RECT 9.792 13.236 9.824 13.308 ;
  LAYER M2 ;
        RECT 9.772 13.256 9.844 13.288 ;
  LAYER M2 ;
        RECT 9.808 13.256 9.968 13.288 ;
  LAYER M1 ;
        RECT 9.952 13.236 9.984 13.308 ;
  LAYER M2 ;
        RECT 9.932 13.256 10.004 13.288 ;
  LAYER M1 ;
        RECT 9.792 16.512 9.824 16.584 ;
  LAYER M2 ;
        RECT 9.772 16.532 9.844 16.564 ;
  LAYER M1 ;
        RECT 9.792 16.38 9.824 16.548 ;
  LAYER M1 ;
        RECT 9.792 16.344 9.824 16.416 ;
  LAYER M2 ;
        RECT 9.772 16.364 9.844 16.396 ;
  LAYER M2 ;
        RECT 9.808 16.364 9.968 16.396 ;
  LAYER M1 ;
        RECT 9.952 16.344 9.984 16.416 ;
  LAYER M2 ;
        RECT 9.932 16.364 10.004 16.396 ;
  LAYER M1 ;
        RECT 9.792 19.62 9.824 19.692 ;
  LAYER M2 ;
        RECT 9.772 19.64 9.844 19.672 ;
  LAYER M1 ;
        RECT 9.792 19.488 9.824 19.656 ;
  LAYER M1 ;
        RECT 9.792 19.452 9.824 19.524 ;
  LAYER M2 ;
        RECT 9.772 19.472 9.844 19.504 ;
  LAYER M2 ;
        RECT 9.808 19.472 9.968 19.504 ;
  LAYER M1 ;
        RECT 9.952 19.452 9.984 19.524 ;
  LAYER M2 ;
        RECT 9.932 19.472 10.004 19.504 ;
  LAYER M1 ;
        RECT 9.792 22.728 9.824 22.8 ;
  LAYER M2 ;
        RECT 9.772 22.748 9.844 22.78 ;
  LAYER M1 ;
        RECT 9.792 22.596 9.824 22.764 ;
  LAYER M1 ;
        RECT 9.792 22.56 9.824 22.632 ;
  LAYER M2 ;
        RECT 9.772 22.58 9.844 22.612 ;
  LAYER M2 ;
        RECT 9.808 22.58 9.968 22.612 ;
  LAYER M1 ;
        RECT 9.952 22.56 9.984 22.632 ;
  LAYER M2 ;
        RECT 9.932 22.58 10.004 22.612 ;
  LAYER M1 ;
        RECT 9.792 25.836 9.824 25.908 ;
  LAYER M2 ;
        RECT 9.772 25.856 9.844 25.888 ;
  LAYER M1 ;
        RECT 9.792 25.704 9.824 25.872 ;
  LAYER M1 ;
        RECT 9.792 25.668 9.824 25.74 ;
  LAYER M2 ;
        RECT 9.772 25.688 9.844 25.72 ;
  LAYER M2 ;
        RECT 9.808 25.688 9.968 25.72 ;
  LAYER M1 ;
        RECT 9.952 25.668 9.984 25.74 ;
  LAYER M2 ;
        RECT 9.932 25.688 10.004 25.72 ;
  LAYER M1 ;
        RECT 9.792 28.944 9.824 29.016 ;
  LAYER M2 ;
        RECT 9.772 28.964 9.844 28.996 ;
  LAYER M1 ;
        RECT 9.792 28.812 9.824 28.98 ;
  LAYER M1 ;
        RECT 9.792 28.776 9.824 28.848 ;
  LAYER M2 ;
        RECT 9.772 28.796 9.844 28.828 ;
  LAYER M2 ;
        RECT 9.808 28.796 9.968 28.828 ;
  LAYER M1 ;
        RECT 9.952 28.776 9.984 28.848 ;
  LAYER M2 ;
        RECT 9.932 28.796 10.004 28.828 ;
  LAYER M1 ;
        RECT 9.792 32.052 9.824 32.124 ;
  LAYER M2 ;
        RECT 9.772 32.072 9.844 32.104 ;
  LAYER M1 ;
        RECT 9.792 31.92 9.824 32.088 ;
  LAYER M1 ;
        RECT 9.792 31.884 9.824 31.956 ;
  LAYER M2 ;
        RECT 9.772 31.904 9.844 31.936 ;
  LAYER M2 ;
        RECT 9.808 31.904 9.968 31.936 ;
  LAYER M1 ;
        RECT 9.952 31.884 9.984 31.956 ;
  LAYER M2 ;
        RECT 9.932 31.904 10.004 31.936 ;
  LAYER M1 ;
        RECT 9.952 0.048 9.984 0.12 ;
  LAYER M2 ;
        RECT 9.932 0.068 10.004 0.1 ;
  LAYER M1 ;
        RECT 9.952 0.084 9.984 0.672 ;
  LAYER M1 ;
        RECT 9.952 0.672 9.984 31.92 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.968 0.1 ;
  LAYER M1 ;
        RECT 6.496 0.972 6.528 1.044 ;
  LAYER M2 ;
        RECT 6.476 0.992 6.548 1.024 ;
  LAYER M2 ;
        RECT 3.216 0.992 6.512 1.024 ;
  LAYER M1 ;
        RECT 3.2 0.972 3.232 1.044 ;
  LAYER M2 ;
        RECT 3.18 0.992 3.252 1.024 ;
  LAYER M1 ;
        RECT 6.496 32.052 6.528 32.124 ;
  LAYER M2 ;
        RECT 6.476 32.072 6.548 32.104 ;
  LAYER M2 ;
        RECT 3.216 32.072 6.512 32.104 ;
  LAYER M1 ;
        RECT 3.2 32.052 3.232 32.124 ;
  LAYER M2 ;
        RECT 3.18 32.072 3.252 32.104 ;
  LAYER M1 ;
        RECT 4.128 18.948 4.16 19.02 ;
  LAYER M2 ;
        RECT 4.108 18.968 4.18 19 ;
  LAYER M2 ;
        RECT 3.824 18.968 4.144 19 ;
  LAYER M1 ;
        RECT 3.808 18.948 3.84 19.02 ;
  LAYER M2 ;
        RECT 3.788 18.968 3.86 19 ;
  LAYER M1 ;
        RECT 4.128 6.516 4.16 6.588 ;
  LAYER M2 ;
        RECT 4.108 6.536 4.18 6.568 ;
  LAYER M2 ;
        RECT 3.824 6.536 4.144 6.568 ;
  LAYER M1 ;
        RECT 3.808 6.516 3.84 6.588 ;
  LAYER M2 ;
        RECT 3.788 6.536 3.86 6.568 ;
  LAYER M1 ;
        RECT 4.128 31.38 4.16 31.452 ;
  LAYER M2 ;
        RECT 4.108 31.4 4.18 31.432 ;
  LAYER M2 ;
        RECT 3.824 31.4 4.144 31.432 ;
  LAYER M1 ;
        RECT 3.808 31.38 3.84 31.452 ;
  LAYER M2 ;
        RECT 3.788 31.4 3.86 31.432 ;
  LAYER M1 ;
        RECT 3.808 35.076 3.84 35.148 ;
  LAYER M2 ;
        RECT 3.788 35.096 3.86 35.128 ;
  LAYER M1 ;
        RECT 3.808 34.86 3.84 35.112 ;
  LAYER M1 ;
        RECT 3.808 6.552 3.84 34.86 ;
  LAYER M1 ;
        RECT 4.128 18.948 4.16 19.02 ;
  LAYER M2 ;
        RECT 4.108 18.968 4.18 19 ;
  LAYER M1 ;
        RECT 4.128 18.984 4.16 19.152 ;
  LAYER M1 ;
        RECT 4.128 19.116 4.16 19.188 ;
  LAYER M2 ;
        RECT 4.108 19.136 4.18 19.168 ;
  LAYER M2 ;
        RECT 4.144 19.136 7.12 19.168 ;
  LAYER M1 ;
        RECT 7.104 19.116 7.136 19.188 ;
  LAYER M2 ;
        RECT 7.084 19.136 7.156 19.168 ;
  LAYER M1 ;
        RECT 4.128 6.516 4.16 6.588 ;
  LAYER M2 ;
        RECT 4.108 6.536 4.18 6.568 ;
  LAYER M1 ;
        RECT 4.128 6.552 4.16 6.72 ;
  LAYER M1 ;
        RECT 4.128 6.684 4.16 6.756 ;
  LAYER M2 ;
        RECT 4.108 6.704 4.18 6.736 ;
  LAYER M2 ;
        RECT 4.144 6.704 7.12 6.736 ;
  LAYER M1 ;
        RECT 7.104 6.684 7.136 6.756 ;
  LAYER M2 ;
        RECT 7.084 6.704 7.156 6.736 ;
  LAYER M1 ;
        RECT 4.128 31.38 4.16 31.452 ;
  LAYER M2 ;
        RECT 4.108 31.4 4.18 31.432 ;
  LAYER M1 ;
        RECT 4.128 31.416 4.16 31.584 ;
  LAYER M1 ;
        RECT 4.128 31.548 4.16 31.62 ;
  LAYER M2 ;
        RECT 4.108 31.568 4.18 31.6 ;
  LAYER M2 ;
        RECT 4.144 31.568 7.12 31.6 ;
  LAYER M1 ;
        RECT 7.104 31.548 7.136 31.62 ;
  LAYER M2 ;
        RECT 7.084 31.568 7.156 31.6 ;
  LAYER M1 ;
        RECT 7.104 35.076 7.136 35.148 ;
  LAYER M2 ;
        RECT 7.084 35.096 7.156 35.128 ;
  LAYER M1 ;
        RECT 7.104 34.86 7.136 35.112 ;
  LAYER M1 ;
        RECT 7.104 6.72 7.136 34.86 ;
  LAYER M2 ;
        RECT 3.824 35.096 7.12 35.128 ;
  LAYER M1 ;
        RECT 4.128 15.84 4.16 15.912 ;
  LAYER M2 ;
        RECT 4.108 15.86 4.18 15.892 ;
  LAYER M2 ;
        RECT 3.984 15.86 4.144 15.892 ;
  LAYER M1 ;
        RECT 3.968 15.84 4 15.912 ;
  LAYER M2 ;
        RECT 3.948 15.86 4.02 15.892 ;
  LAYER M1 ;
        RECT 4.128 22.056 4.16 22.128 ;
  LAYER M2 ;
        RECT 4.108 22.076 4.18 22.108 ;
  LAYER M2 ;
        RECT 3.984 22.076 4.144 22.108 ;
  LAYER M1 ;
        RECT 3.968 22.056 4 22.128 ;
  LAYER M2 ;
        RECT 3.948 22.076 4.02 22.108 ;
  LAYER M1 ;
        RECT 4.128 12.732 4.16 12.804 ;
  LAYER M2 ;
        RECT 4.108 12.752 4.18 12.784 ;
  LAYER M2 ;
        RECT 3.984 12.752 4.144 12.784 ;
  LAYER M1 ;
        RECT 3.968 12.732 4 12.804 ;
  LAYER M2 ;
        RECT 3.948 12.752 4.02 12.784 ;
  LAYER M1 ;
        RECT 4.128 25.164 4.16 25.236 ;
  LAYER M2 ;
        RECT 4.108 25.184 4.18 25.216 ;
  LAYER M2 ;
        RECT 3.984 25.184 4.144 25.216 ;
  LAYER M1 ;
        RECT 3.968 25.164 4 25.236 ;
  LAYER M2 ;
        RECT 3.948 25.184 4.02 25.216 ;
  LAYER M1 ;
        RECT 4.128 9.624 4.16 9.696 ;
  LAYER M2 ;
        RECT 4.108 9.644 4.18 9.676 ;
  LAYER M2 ;
        RECT 3.984 9.644 4.144 9.676 ;
  LAYER M1 ;
        RECT 3.968 9.624 4 9.696 ;
  LAYER M2 ;
        RECT 3.948 9.644 4.02 9.676 ;
  LAYER M1 ;
        RECT 4.128 28.272 4.16 28.344 ;
  LAYER M2 ;
        RECT 4.108 28.292 4.18 28.324 ;
  LAYER M2 ;
        RECT 3.984 28.292 4.144 28.324 ;
  LAYER M1 ;
        RECT 3.968 28.272 4 28.344 ;
  LAYER M2 ;
        RECT 3.948 28.292 4.02 28.324 ;
  LAYER M1 ;
        RECT 3.968 35.244 4 35.316 ;
  LAYER M2 ;
        RECT 3.948 35.264 4.02 35.296 ;
  LAYER M1 ;
        RECT 3.968 34.86 4 35.28 ;
  LAYER M1 ;
        RECT 3.968 9.66 4 34.86 ;
  LAYER M1 ;
        RECT 4.128 15.84 4.16 15.912 ;
  LAYER M2 ;
        RECT 4.108 15.86 4.18 15.892 ;
  LAYER M1 ;
        RECT 4.128 15.876 4.16 16.044 ;
  LAYER M1 ;
        RECT 4.128 16.008 4.16 16.08 ;
  LAYER M2 ;
        RECT 4.108 16.028 4.18 16.06 ;
  LAYER M2 ;
        RECT 4.144 16.028 7.28 16.06 ;
  LAYER M1 ;
        RECT 7.264 16.008 7.296 16.08 ;
  LAYER M2 ;
        RECT 7.244 16.028 7.316 16.06 ;
  LAYER M1 ;
        RECT 4.128 22.056 4.16 22.128 ;
  LAYER M2 ;
        RECT 4.108 22.076 4.18 22.108 ;
  LAYER M1 ;
        RECT 4.128 22.092 4.16 22.26 ;
  LAYER M1 ;
        RECT 4.128 22.224 4.16 22.296 ;
  LAYER M2 ;
        RECT 4.108 22.244 4.18 22.276 ;
  LAYER M2 ;
        RECT 4.144 22.244 7.28 22.276 ;
  LAYER M1 ;
        RECT 7.264 22.224 7.296 22.296 ;
  LAYER M2 ;
        RECT 7.244 22.244 7.316 22.276 ;
  LAYER M1 ;
        RECT 4.128 12.732 4.16 12.804 ;
  LAYER M2 ;
        RECT 4.108 12.752 4.18 12.784 ;
  LAYER M1 ;
        RECT 4.128 12.768 4.16 12.936 ;
  LAYER M1 ;
        RECT 4.128 12.9 4.16 12.972 ;
  LAYER M2 ;
        RECT 4.108 12.92 4.18 12.952 ;
  LAYER M2 ;
        RECT 4.144 12.92 7.28 12.952 ;
  LAYER M1 ;
        RECT 7.264 12.9 7.296 12.972 ;
  LAYER M2 ;
        RECT 7.244 12.92 7.316 12.952 ;
  LAYER M1 ;
        RECT 4.128 25.164 4.16 25.236 ;
  LAYER M2 ;
        RECT 4.108 25.184 4.18 25.216 ;
  LAYER M1 ;
        RECT 4.128 25.2 4.16 25.368 ;
  LAYER M1 ;
        RECT 4.128 25.332 4.16 25.404 ;
  LAYER M2 ;
        RECT 4.108 25.352 4.18 25.384 ;
  LAYER M2 ;
        RECT 4.144 25.352 7.28 25.384 ;
  LAYER M1 ;
        RECT 7.264 25.332 7.296 25.404 ;
  LAYER M2 ;
        RECT 7.244 25.352 7.316 25.384 ;
  LAYER M1 ;
        RECT 4.128 9.624 4.16 9.696 ;
  LAYER M2 ;
        RECT 4.108 9.644 4.18 9.676 ;
  LAYER M1 ;
        RECT 4.128 9.66 4.16 9.828 ;
  LAYER M1 ;
        RECT 4.128 9.792 4.16 9.864 ;
  LAYER M2 ;
        RECT 4.108 9.812 4.18 9.844 ;
  LAYER M2 ;
        RECT 4.144 9.812 7.28 9.844 ;
  LAYER M1 ;
        RECT 7.264 9.792 7.296 9.864 ;
  LAYER M2 ;
        RECT 7.244 9.812 7.316 9.844 ;
  LAYER M1 ;
        RECT 4.128 28.272 4.16 28.344 ;
  LAYER M2 ;
        RECT 4.108 28.292 4.18 28.324 ;
  LAYER M1 ;
        RECT 4.128 28.308 4.16 28.476 ;
  LAYER M1 ;
        RECT 4.128 28.44 4.16 28.512 ;
  LAYER M2 ;
        RECT 4.108 28.46 4.18 28.492 ;
  LAYER M2 ;
        RECT 4.144 28.46 7.28 28.492 ;
  LAYER M1 ;
        RECT 7.264 28.44 7.296 28.512 ;
  LAYER M2 ;
        RECT 7.244 28.46 7.316 28.492 ;
  LAYER M1 ;
        RECT 7.264 35.244 7.296 35.316 ;
  LAYER M2 ;
        RECT 7.244 35.264 7.316 35.296 ;
  LAYER M1 ;
        RECT 7.264 34.86 7.296 35.28 ;
  LAYER M1 ;
        RECT 7.264 9.828 7.296 34.86 ;
  LAYER M2 ;
        RECT 3.984 35.264 7.28 35.296 ;
  LAYER M1 ;
        RECT 0.832 3.408 0.864 3.48 ;
  LAYER M2 ;
        RECT 0.812 3.428 0.884 3.46 ;
  LAYER M2 ;
        RECT 0.368 3.428 0.848 3.46 ;
  LAYER M1 ;
        RECT 0.352 3.408 0.384 3.48 ;
  LAYER M2 ;
        RECT 0.332 3.428 0.404 3.46 ;
  LAYER M1 ;
        RECT 0.832 6.516 0.864 6.588 ;
  LAYER M2 ;
        RECT 0.812 6.536 0.884 6.568 ;
  LAYER M2 ;
        RECT 0.368 6.536 0.848 6.568 ;
  LAYER M1 ;
        RECT 0.352 6.516 0.384 6.588 ;
  LAYER M2 ;
        RECT 0.332 6.536 0.404 6.568 ;
  LAYER M1 ;
        RECT 0.832 9.624 0.864 9.696 ;
  LAYER M2 ;
        RECT 0.812 9.644 0.884 9.676 ;
  LAYER M2 ;
        RECT 0.368 9.644 0.848 9.676 ;
  LAYER M1 ;
        RECT 0.352 9.624 0.384 9.696 ;
  LAYER M2 ;
        RECT 0.332 9.644 0.404 9.676 ;
  LAYER M1 ;
        RECT 0.832 12.732 0.864 12.804 ;
  LAYER M2 ;
        RECT 0.812 12.752 0.884 12.784 ;
  LAYER M2 ;
        RECT 0.368 12.752 0.848 12.784 ;
  LAYER M1 ;
        RECT 0.352 12.732 0.384 12.804 ;
  LAYER M2 ;
        RECT 0.332 12.752 0.404 12.784 ;
  LAYER M1 ;
        RECT 0.832 15.84 0.864 15.912 ;
  LAYER M2 ;
        RECT 0.812 15.86 0.884 15.892 ;
  LAYER M2 ;
        RECT 0.368 15.86 0.848 15.892 ;
  LAYER M1 ;
        RECT 0.352 15.84 0.384 15.912 ;
  LAYER M2 ;
        RECT 0.332 15.86 0.404 15.892 ;
  LAYER M1 ;
        RECT 0.832 18.948 0.864 19.02 ;
  LAYER M2 ;
        RECT 0.812 18.968 0.884 19 ;
  LAYER M2 ;
        RECT 0.368 18.968 0.848 19 ;
  LAYER M1 ;
        RECT 0.352 18.948 0.384 19.02 ;
  LAYER M2 ;
        RECT 0.332 18.968 0.404 19 ;
  LAYER M1 ;
        RECT 0.832 22.056 0.864 22.128 ;
  LAYER M2 ;
        RECT 0.812 22.076 0.884 22.108 ;
  LAYER M2 ;
        RECT 0.368 22.076 0.848 22.108 ;
  LAYER M1 ;
        RECT 0.352 22.056 0.384 22.128 ;
  LAYER M2 ;
        RECT 0.332 22.076 0.404 22.108 ;
  LAYER M1 ;
        RECT 0.832 25.164 0.864 25.236 ;
  LAYER M2 ;
        RECT 0.812 25.184 0.884 25.216 ;
  LAYER M2 ;
        RECT 0.368 25.184 0.848 25.216 ;
  LAYER M1 ;
        RECT 0.352 25.164 0.384 25.236 ;
  LAYER M2 ;
        RECT 0.332 25.184 0.404 25.216 ;
  LAYER M1 ;
        RECT 0.832 28.272 0.864 28.344 ;
  LAYER M2 ;
        RECT 0.812 28.292 0.884 28.324 ;
  LAYER M2 ;
        RECT 0.368 28.292 0.848 28.324 ;
  LAYER M1 ;
        RECT 0.352 28.272 0.384 28.344 ;
  LAYER M2 ;
        RECT 0.332 28.292 0.404 28.324 ;
  LAYER M1 ;
        RECT 0.832 31.38 0.864 31.452 ;
  LAYER M2 ;
        RECT 0.812 31.4 0.884 31.432 ;
  LAYER M2 ;
        RECT 0.368 31.4 0.848 31.432 ;
  LAYER M1 ;
        RECT 0.352 31.38 0.384 31.452 ;
  LAYER M2 ;
        RECT 0.332 31.4 0.404 31.432 ;
  LAYER M1 ;
        RECT 0.832 34.488 0.864 34.56 ;
  LAYER M2 ;
        RECT 0.812 34.508 0.884 34.54 ;
  LAYER M2 ;
        RECT 0.368 34.508 0.848 34.54 ;
  LAYER M1 ;
        RECT 0.352 34.488 0.384 34.56 ;
  LAYER M2 ;
        RECT 0.332 34.508 0.404 34.54 ;
  LAYER M1 ;
        RECT 0.352 35.412 0.384 35.484 ;
  LAYER M2 ;
        RECT 0.332 35.432 0.404 35.464 ;
  LAYER M1 ;
        RECT 0.352 34.86 0.384 35.448 ;
  LAYER M1 ;
        RECT 0.352 3.444 0.384 34.86 ;
  LAYER M1 ;
        RECT 7.424 3.408 7.456 3.48 ;
  LAYER M2 ;
        RECT 7.404 3.428 7.476 3.46 ;
  LAYER M1 ;
        RECT 7.424 3.444 7.456 3.612 ;
  LAYER M1 ;
        RECT 7.424 3.576 7.456 3.648 ;
  LAYER M2 ;
        RECT 7.404 3.596 7.476 3.628 ;
  LAYER M2 ;
        RECT 7.44 3.596 10.256 3.628 ;
  LAYER M1 ;
        RECT 10.24 3.576 10.272 3.648 ;
  LAYER M2 ;
        RECT 10.22 3.596 10.292 3.628 ;
  LAYER M1 ;
        RECT 7.424 6.516 7.456 6.588 ;
  LAYER M2 ;
        RECT 7.404 6.536 7.476 6.568 ;
  LAYER M1 ;
        RECT 7.424 6.552 7.456 6.72 ;
  LAYER M1 ;
        RECT 7.424 6.684 7.456 6.756 ;
  LAYER M2 ;
        RECT 7.404 6.704 7.476 6.736 ;
  LAYER M2 ;
        RECT 7.44 6.704 10.256 6.736 ;
  LAYER M1 ;
        RECT 10.24 6.684 10.272 6.756 ;
  LAYER M2 ;
        RECT 10.22 6.704 10.292 6.736 ;
  LAYER M1 ;
        RECT 7.424 9.624 7.456 9.696 ;
  LAYER M2 ;
        RECT 7.404 9.644 7.476 9.676 ;
  LAYER M1 ;
        RECT 7.424 9.66 7.456 9.828 ;
  LAYER M1 ;
        RECT 7.424 9.792 7.456 9.864 ;
  LAYER M2 ;
        RECT 7.404 9.812 7.476 9.844 ;
  LAYER M2 ;
        RECT 7.44 9.812 10.256 9.844 ;
  LAYER M1 ;
        RECT 10.24 9.792 10.272 9.864 ;
  LAYER M2 ;
        RECT 10.22 9.812 10.292 9.844 ;
  LAYER M1 ;
        RECT 7.424 12.732 7.456 12.804 ;
  LAYER M2 ;
        RECT 7.404 12.752 7.476 12.784 ;
  LAYER M1 ;
        RECT 7.424 12.768 7.456 12.936 ;
  LAYER M1 ;
        RECT 7.424 12.9 7.456 12.972 ;
  LAYER M2 ;
        RECT 7.404 12.92 7.476 12.952 ;
  LAYER M2 ;
        RECT 7.44 12.92 10.256 12.952 ;
  LAYER M1 ;
        RECT 10.24 12.9 10.272 12.972 ;
  LAYER M2 ;
        RECT 10.22 12.92 10.292 12.952 ;
  LAYER M1 ;
        RECT 7.424 15.84 7.456 15.912 ;
  LAYER M2 ;
        RECT 7.404 15.86 7.476 15.892 ;
  LAYER M1 ;
        RECT 7.424 15.876 7.456 16.044 ;
  LAYER M1 ;
        RECT 7.424 16.008 7.456 16.08 ;
  LAYER M2 ;
        RECT 7.404 16.028 7.476 16.06 ;
  LAYER M2 ;
        RECT 7.44 16.028 10.256 16.06 ;
  LAYER M1 ;
        RECT 10.24 16.008 10.272 16.08 ;
  LAYER M2 ;
        RECT 10.22 16.028 10.292 16.06 ;
  LAYER M1 ;
        RECT 7.424 18.948 7.456 19.02 ;
  LAYER M2 ;
        RECT 7.404 18.968 7.476 19 ;
  LAYER M1 ;
        RECT 7.424 18.984 7.456 19.152 ;
  LAYER M1 ;
        RECT 7.424 19.116 7.456 19.188 ;
  LAYER M2 ;
        RECT 7.404 19.136 7.476 19.168 ;
  LAYER M2 ;
        RECT 7.44 19.136 10.256 19.168 ;
  LAYER M1 ;
        RECT 10.24 19.116 10.272 19.188 ;
  LAYER M2 ;
        RECT 10.22 19.136 10.292 19.168 ;
  LAYER M1 ;
        RECT 7.424 22.056 7.456 22.128 ;
  LAYER M2 ;
        RECT 7.404 22.076 7.476 22.108 ;
  LAYER M1 ;
        RECT 7.424 22.092 7.456 22.26 ;
  LAYER M1 ;
        RECT 7.424 22.224 7.456 22.296 ;
  LAYER M2 ;
        RECT 7.404 22.244 7.476 22.276 ;
  LAYER M2 ;
        RECT 7.44 22.244 10.256 22.276 ;
  LAYER M1 ;
        RECT 10.24 22.224 10.272 22.296 ;
  LAYER M2 ;
        RECT 10.22 22.244 10.292 22.276 ;
  LAYER M1 ;
        RECT 7.424 25.164 7.456 25.236 ;
  LAYER M2 ;
        RECT 7.404 25.184 7.476 25.216 ;
  LAYER M1 ;
        RECT 7.424 25.2 7.456 25.368 ;
  LAYER M1 ;
        RECT 7.424 25.332 7.456 25.404 ;
  LAYER M2 ;
        RECT 7.404 25.352 7.476 25.384 ;
  LAYER M2 ;
        RECT 7.44 25.352 10.256 25.384 ;
  LAYER M1 ;
        RECT 10.24 25.332 10.272 25.404 ;
  LAYER M2 ;
        RECT 10.22 25.352 10.292 25.384 ;
  LAYER M1 ;
        RECT 7.424 28.272 7.456 28.344 ;
  LAYER M2 ;
        RECT 7.404 28.292 7.476 28.324 ;
  LAYER M1 ;
        RECT 7.424 28.308 7.456 28.476 ;
  LAYER M1 ;
        RECT 7.424 28.44 7.456 28.512 ;
  LAYER M2 ;
        RECT 7.404 28.46 7.476 28.492 ;
  LAYER M2 ;
        RECT 7.44 28.46 10.256 28.492 ;
  LAYER M1 ;
        RECT 10.24 28.44 10.272 28.512 ;
  LAYER M2 ;
        RECT 10.22 28.46 10.292 28.492 ;
  LAYER M1 ;
        RECT 7.424 31.38 7.456 31.452 ;
  LAYER M2 ;
        RECT 7.404 31.4 7.476 31.432 ;
  LAYER M1 ;
        RECT 7.424 31.416 7.456 31.584 ;
  LAYER M1 ;
        RECT 7.424 31.548 7.456 31.62 ;
  LAYER M2 ;
        RECT 7.404 31.568 7.476 31.6 ;
  LAYER M2 ;
        RECT 7.44 31.568 10.256 31.6 ;
  LAYER M1 ;
        RECT 10.24 31.548 10.272 31.62 ;
  LAYER M2 ;
        RECT 10.22 31.568 10.292 31.6 ;
  LAYER M1 ;
        RECT 7.424 34.488 7.456 34.56 ;
  LAYER M2 ;
        RECT 7.404 34.508 7.476 34.54 ;
  LAYER M1 ;
        RECT 7.424 34.524 7.456 34.692 ;
  LAYER M1 ;
        RECT 7.424 34.656 7.456 34.728 ;
  LAYER M2 ;
        RECT 7.404 34.676 7.476 34.708 ;
  LAYER M2 ;
        RECT 7.44 34.676 10.256 34.708 ;
  LAYER M1 ;
        RECT 10.24 34.656 10.272 34.728 ;
  LAYER M2 ;
        RECT 10.22 34.676 10.292 34.708 ;
  LAYER M1 ;
        RECT 10.24 35.412 10.272 35.484 ;
  LAYER M2 ;
        RECT 10.22 35.432 10.292 35.464 ;
  LAYER M1 ;
        RECT 10.24 34.86 10.272 35.448 ;
  LAYER M1 ;
        RECT 10.24 3.612 10.272 34.86 ;
  LAYER M2 ;
        RECT 0.368 35.432 10.256 35.464 ;
  LAYER M1 ;
        RECT 4.128 3.408 4.16 3.48 ;
  LAYER M2 ;
        RECT 4.108 3.428 4.18 3.46 ;
  LAYER M2 ;
        RECT 0.848 3.428 4.144 3.46 ;
  LAYER M1 ;
        RECT 0.832 3.408 0.864 3.48 ;
  LAYER M2 ;
        RECT 0.812 3.428 0.884 3.46 ;
  LAYER M1 ;
        RECT 4.128 34.488 4.16 34.56 ;
  LAYER M2 ;
        RECT 4.108 34.508 4.18 34.54 ;
  LAYER M2 ;
        RECT 0.848 34.508 4.144 34.54 ;
  LAYER M1 ;
        RECT 0.832 34.488 0.864 34.56 ;
  LAYER M2 ;
        RECT 0.812 34.508 0.884 34.54 ;
  LAYER M1 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M3 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M2 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M1 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M3 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M2 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M1 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M3 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M2 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M1 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M3 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M2 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M1 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M3 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M2 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M1 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M3 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M2 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M1 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M3 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M2 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M1 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M3 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M2 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M1 ;
        RECT 0.784 25.788 3.28 28.392 ;
  LAYER M3 ;
        RECT 0.784 25.788 3.28 28.392 ;
  LAYER M2 ;
        RECT 0.784 25.788 3.28 28.392 ;
  LAYER M1 ;
        RECT 0.784 28.896 3.28 31.5 ;
  LAYER M3 ;
        RECT 0.784 28.896 3.28 31.5 ;
  LAYER M2 ;
        RECT 0.784 28.896 3.28 31.5 ;
  LAYER M1 ;
        RECT 0.784 32.004 3.28 34.608 ;
  LAYER M3 ;
        RECT 0.784 32.004 3.28 34.608 ;
  LAYER M2 ;
        RECT 0.784 32.004 3.28 34.608 ;
  LAYER M1 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M3 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M2 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M1 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M3 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M2 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M1 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M3 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M2 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M1 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M3 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M2 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M1 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M3 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M2 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M1 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M3 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M2 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M1 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M3 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M2 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M1 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M3 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M2 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M1 ;
        RECT 4.08 25.788 6.576 28.392 ;
  LAYER M3 ;
        RECT 4.08 25.788 6.576 28.392 ;
  LAYER M2 ;
        RECT 4.08 25.788 6.576 28.392 ;
  LAYER M1 ;
        RECT 4.08 28.896 6.576 31.5 ;
  LAYER M3 ;
        RECT 4.08 28.896 6.576 31.5 ;
  LAYER M2 ;
        RECT 4.08 28.896 6.576 31.5 ;
  LAYER M1 ;
        RECT 4.08 32.004 6.576 34.608 ;
  LAYER M3 ;
        RECT 4.08 32.004 6.576 34.608 ;
  LAYER M2 ;
        RECT 4.08 32.004 6.576 34.608 ;
  LAYER M1 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M3 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M2 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M1 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M3 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M2 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M1 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M3 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M2 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M1 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M3 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M2 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M1 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M3 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M2 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M1 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M3 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M2 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M1 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M3 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M2 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M1 ;
        RECT 7.376 22.68 9.872 25.284 ;
  LAYER M3 ;
        RECT 7.376 22.68 9.872 25.284 ;
  LAYER M2 ;
        RECT 7.376 22.68 9.872 25.284 ;
  LAYER M1 ;
        RECT 7.376 25.788 9.872 28.392 ;
  LAYER M3 ;
        RECT 7.376 25.788 9.872 28.392 ;
  LAYER M2 ;
        RECT 7.376 25.788 9.872 28.392 ;
  LAYER M1 ;
        RECT 7.376 28.896 9.872 31.5 ;
  LAYER M3 ;
        RECT 7.376 28.896 9.872 31.5 ;
  LAYER M2 ;
        RECT 7.376 28.896 9.872 31.5 ;
  LAYER M1 ;
        RECT 7.376 32.004 9.872 34.608 ;
  LAYER M3 ;
        RECT 7.376 32.004 9.872 34.608 ;
  LAYER M2 ;
        RECT 7.376 32.004 9.872 34.608 ;
  END 
END Cap_30fF_Cap_60fF
