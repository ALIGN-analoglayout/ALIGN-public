MACRO CMC_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.8440 0.2360 3.4760 0.2680 ;
    LAYER M2 ;
      RECT 1.0040 0.3200 3.6360 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.4040 3.5560 0.4360 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
  END
END CMC_NMOS_n12_X3_Y1
MACRO CMC_PMOS_S_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.0760 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.5960 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 0.9960 0.3520 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END CMC_PMOS_S_n12_X1_Y1
MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.3560 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.1960 0.1840 ;
    LAYER M2 ;
      RECT 0.8440 0.2360 1.7160 0.2680 ;
    LAYER M2 ;
      RECT 1.0040 0.3200 1.5560 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.4040 2.2760 0.4360 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
  END
END CMC_PMOS_n12_X2_Y1
MACRO CMFB_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMFB_NMOS_n12_X3_Y1 0 0 ;
  SIZE 5.1200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END DB
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M1 ;
      RECT 4.1440 0.0480 4.1760 0.7080 ;
    LAYER M1 ;
      RECT 4.0640 0.0480 4.0960 0.7080 ;
    LAYER M1 ;
      RECT 4.2240 0.0480 4.2560 0.7080 ;
    LAYER M1 ;
      RECT 4.7840 0.0480 4.8160 0.7080 ;
    LAYER M1 ;
      RECT 4.7040 0.0480 4.7360 0.7080 ;
    LAYER M1 ;
      RECT 4.8640 0.0480 4.8960 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 4.7560 0.1000 ;
    LAYER M2 ;
      RECT 2.2040 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.2360 4.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 4.8360 0.3520 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
    LAYER pc ;
      RECT 4.1110 0.0680 4.2090 0.1000 ;
    LAYER pc ;
      RECT 4.7510 0.0680 4.8490 0.1000 ;
  END
END CMFB_NMOS_n12_X3_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 1.0760 0.1840 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DP_NMOS_n12_X3_Y3
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X3_Y3 0 0 ;
  SIZE 3.8400 BY 2.5200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.7400 0.0480 1.7800 1.8000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.8200 0.1320 1.8600 1.8840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9000 0.2160 1.9400 1.9680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9800 0.3000 2.0200 2.0520 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.0600 0.3840 2.1000 2.1360 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.3040 1.7280 0.3360 2.3880 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 1.7280 0.2560 2.3880 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 1.7280 0.4160 2.3880 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 1.7280 0.9760 2.3880 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 0.8640 1.7280 0.8960 2.3880 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 1.7280 1.0560 2.3880 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 1.7280 1.6160 2.3880 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.5040 1.7280 1.5360 2.3880 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 1.7280 1.6960 2.3880 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 1.7280 2.2560 2.3880 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER M1 ;
      RECT 2.1440 1.7280 2.1760 2.3880 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER M1 ;
      RECT 2.3040 1.7280 2.3360 2.3880 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 1.7280 2.8960 2.3880 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER M1 ;
      RECT 2.7840 1.7280 2.8160 2.3880 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER M1 ;
      RECT 2.9440 1.7280 2.9760 2.3880 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.8880 3.5360 1.5480 ;
    LAYER M1 ;
      RECT 3.5040 1.7280 3.5360 2.3880 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.8880 3.4560 1.5480 ;
    LAYER M1 ;
      RECT 3.4240 1.7280 3.4560 2.3880 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.8880 3.6160 1.5480 ;
    LAYER M1 ;
      RECT 3.5840 1.7280 3.6160 2.3880 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 3.4760 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 1.0040 0.2360 3.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 2.9160 0.3520 ;
    LAYER M2 ;
      RECT 0.9240 0.4040 3.5560 0.4360 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 3.4760 0.9400 ;
    LAYER M2 ;
      RECT 1.0040 0.9920 3.6360 1.0240 ;
    LAYER M2 ;
      RECT 0.3640 1.0760 2.9960 1.1080 ;
    LAYER M2 ;
      RECT 0.9240 1.1600 3.5560 1.1920 ;
    LAYER M2 ;
      RECT 0.2840 1.2440 2.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.2040 1.7480 3.4760 1.7800 ;
    LAYER M2 ;
      RECT 0.3640 1.8320 2.9960 1.8640 ;
    LAYER M2 ;
      RECT 1.0040 1.9160 3.6360 1.9480 ;
    LAYER M2 ;
      RECT 0.2840 2.0000 2.9160 2.0320 ;
    LAYER M2 ;
      RECT 0.9240 2.0840 3.5560 2.1160 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
    LAYER pc ;
      RECT 0.2710 0.9080 0.3690 0.9400 ;
    LAYER pc ;
      RECT 0.9110 0.9080 1.0090 0.9400 ;
    LAYER pc ;
      RECT 1.5510 0.9080 1.6490 0.9400 ;
    LAYER pc ;
      RECT 2.1910 0.9080 2.2890 0.9400 ;
    LAYER pc ;
      RECT 2.8310 0.9080 2.9290 0.9400 ;
    LAYER pc ;
      RECT 3.4710 0.9080 3.5690 0.9400 ;
    LAYER pc ;
      RECT 0.2710 1.7480 0.3690 1.7800 ;
    LAYER pc ;
      RECT 0.9110 1.7480 1.0090 1.7800 ;
    LAYER pc ;
      RECT 1.5510 1.7480 1.6490 1.7800 ;
    LAYER pc ;
      RECT 2.1910 1.7480 2.2890 1.7800 ;
    LAYER pc ;
      RECT 2.8310 1.7480 2.9290 1.7800 ;
    LAYER pc ;
      RECT 3.4710 1.7480 3.5690 1.7800 ;
  END
END DP_NMOS_n12_X3_Y3
MACRO Switch_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y1 0 0 ;
  SIZE 1.9200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 1.6360 0.2680 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
  END
END Switch_NMOS_n12_X3_Y1
MACRO Switch_NMOS_n12_X3_Y3
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y3 0 0 ;
  SIZE 1.9200 BY 2.5200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8600 0.0480 0.9000 1.8000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9400 0.1320 0.9800 1.8840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.0200 0.2160 1.0600 1.9680 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.3040 1.7280 0.3360 2.3880 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 1.7280 0.2560 2.3880 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 1.7280 0.4160 2.3880 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 1.7280 0.9760 2.3880 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 0.8640 1.7280 0.8960 2.3880 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 1.7280 1.0560 2.3880 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 1.7280 1.6160 2.3880 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.5040 1.7280 1.5360 2.3880 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 1.7280 1.6960 2.3880 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 1.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 1.5560 0.9400 ;
    LAYER M2 ;
      RECT 0.3640 0.9920 1.7160 1.0240 ;
    LAYER M2 ;
      RECT 0.2840 1.0760 1.6360 1.1080 ;
    LAYER M2 ;
      RECT 0.2040 1.7480 1.5560 1.7800 ;
    LAYER M2 ;
      RECT 0.3640 1.8320 1.7160 1.8640 ;
    LAYER M2 ;
      RECT 0.2840 1.9160 1.6360 1.9480 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 0.2710 0.9080 0.3690 0.9400 ;
    LAYER pc ;
      RECT 0.9110 0.9080 1.0090 0.9400 ;
    LAYER pc ;
      RECT 1.5510 0.9080 1.6490 0.9400 ;
    LAYER pc ;
      RECT 0.2710 1.7480 0.3690 1.7800 ;
    LAYER pc ;
      RECT 0.9110 1.7480 1.0090 1.7800 ;
    LAYER pc ;
      RECT 1.5510 1.7480 1.6490 1.7800 ;
  END
END Switch_NMOS_n12_X3_Y3
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1520 0.4360 0.1840 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.5160 0.2680 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.0760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.9960 0.2680 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END Switch_PMOS_n12_X2_Y1
