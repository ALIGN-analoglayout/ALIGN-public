MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 9.28 BY 25.872 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 25.584 3.232 25.656 ;
      LAYER M2 ;
        RECT 3.18 25.604 3.252 25.636 ;
      LAYER M1 ;
        RECT 6.176 25.584 6.208 25.656 ;
      LAYER M2 ;
        RECT 6.156 25.604 6.228 25.636 ;
      LAYER M2 ;
        RECT 3.216 25.604 6.192 25.636 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 3.056 10.148 5.808 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M2 ;
        RECT 3.056 13.256 5.808 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M2 ;
        RECT 3.056 7.04 5.808 7.072 ;
  LAYER M1 ;
        RECT 3.04 7.02 3.072 7.092 ;
  LAYER M2 ;
        RECT 3.02 7.04 3.092 7.072 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 16.416 ;
  LAYER M2 ;
        RECT 5.772 16.364 5.844 16.396 ;
  LAYER M2 ;
        RECT 3.056 16.364 5.808 16.396 ;
  LAYER M1 ;
        RECT 3.04 16.344 3.072 16.416 ;
  LAYER M2 ;
        RECT 3.02 16.364 3.092 16.396 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M2 ;
        RECT 3.056 3.932 5.808 3.964 ;
  LAYER M1 ;
        RECT 3.04 3.912 3.072 3.984 ;
  LAYER M2 ;
        RECT 3.02 3.932 3.092 3.964 ;
  LAYER M1 ;
        RECT 5.792 19.452 5.824 19.524 ;
  LAYER M2 ;
        RECT 5.772 19.472 5.844 19.504 ;
  LAYER M2 ;
        RECT 3.056 19.472 5.808 19.504 ;
  LAYER M1 ;
        RECT 3.04 19.452 3.072 19.524 ;
  LAYER M2 ;
        RECT 3.02 19.472 3.092 19.504 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.504 ;
  LAYER M1 ;
        RECT 3.04 0.504 3.072 19.488 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M1 ;
        RECT 5.792 9.996 5.824 10.164 ;
  LAYER M1 ;
        RECT 5.792 9.96 5.824 10.032 ;
  LAYER M2 ;
        RECT 5.772 9.98 5.844 10.012 ;
  LAYER M2 ;
        RECT 5.808 9.98 6.032 10.012 ;
  LAYER M1 ;
        RECT 6.016 9.96 6.048 10.032 ;
  LAYER M2 ;
        RECT 5.996 9.98 6.068 10.012 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M1 ;
        RECT 5.792 13.104 5.824 13.272 ;
  LAYER M1 ;
        RECT 5.792 13.068 5.824 13.14 ;
  LAYER M2 ;
        RECT 5.772 13.088 5.844 13.12 ;
  LAYER M2 ;
        RECT 5.808 13.088 6.032 13.12 ;
  LAYER M1 ;
        RECT 6.016 13.068 6.048 13.14 ;
  LAYER M2 ;
        RECT 5.996 13.088 6.068 13.12 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M1 ;
        RECT 5.792 6.888 5.824 7.056 ;
  LAYER M1 ;
        RECT 5.792 6.852 5.824 6.924 ;
  LAYER M2 ;
        RECT 5.772 6.872 5.844 6.904 ;
  LAYER M2 ;
        RECT 5.808 6.872 6.032 6.904 ;
  LAYER M1 ;
        RECT 6.016 6.852 6.048 6.924 ;
  LAYER M2 ;
        RECT 5.996 6.872 6.068 6.904 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 16.416 ;
  LAYER M2 ;
        RECT 5.772 16.364 5.844 16.396 ;
  LAYER M1 ;
        RECT 5.792 16.212 5.824 16.38 ;
  LAYER M1 ;
        RECT 5.792 16.176 5.824 16.248 ;
  LAYER M2 ;
        RECT 5.772 16.196 5.844 16.228 ;
  LAYER M2 ;
        RECT 5.808 16.196 6.032 16.228 ;
  LAYER M1 ;
        RECT 6.016 16.176 6.048 16.248 ;
  LAYER M2 ;
        RECT 5.996 16.196 6.068 16.228 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M1 ;
        RECT 5.792 3.78 5.824 3.948 ;
  LAYER M1 ;
        RECT 5.792 3.744 5.824 3.816 ;
  LAYER M2 ;
        RECT 5.772 3.764 5.844 3.796 ;
  LAYER M2 ;
        RECT 5.808 3.764 6.032 3.796 ;
  LAYER M1 ;
        RECT 6.016 3.744 6.048 3.816 ;
  LAYER M2 ;
        RECT 5.996 3.764 6.068 3.796 ;
  LAYER M1 ;
        RECT 5.792 19.452 5.824 19.524 ;
  LAYER M2 ;
        RECT 5.772 19.472 5.844 19.504 ;
  LAYER M1 ;
        RECT 5.792 19.32 5.824 19.488 ;
  LAYER M1 ;
        RECT 5.792 19.284 5.824 19.356 ;
  LAYER M2 ;
        RECT 5.772 19.304 5.844 19.336 ;
  LAYER M2 ;
        RECT 5.808 19.304 6.032 19.336 ;
  LAYER M1 ;
        RECT 6.016 19.284 6.048 19.356 ;
  LAYER M2 ;
        RECT 5.996 19.304 6.068 19.336 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.504 ;
  LAYER M1 ;
        RECT 6.016 0.504 6.048 19.32 ;
  LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M2 ;
        RECT 0.08 0.824 2.832 0.856 ;
  LAYER M1 ;
        RECT 0.064 0.804 0.096 0.876 ;
  LAYER M2 ;
        RECT 0.044 0.824 0.116 0.856 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M2 ;
        RECT 0.08 3.932 2.832 3.964 ;
  LAYER M1 ;
        RECT 0.064 3.912 0.096 3.984 ;
  LAYER M2 ;
        RECT 0.044 3.932 0.116 3.964 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M2 ;
        RECT 0.08 7.04 2.832 7.072 ;
  LAYER M1 ;
        RECT 0.064 7.02 0.096 7.092 ;
  LAYER M2 ;
        RECT 0.044 7.04 0.116 7.072 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M2 ;
        RECT 0.08 10.148 2.832 10.18 ;
  LAYER M1 ;
        RECT 0.064 10.128 0.096 10.2 ;
  LAYER M2 ;
        RECT 0.044 10.148 0.116 10.18 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 13.308 ;
  LAYER M2 ;
        RECT 2.796 13.256 2.868 13.288 ;
  LAYER M2 ;
        RECT 0.08 13.256 2.832 13.288 ;
  LAYER M1 ;
        RECT 0.064 13.236 0.096 13.308 ;
  LAYER M2 ;
        RECT 0.044 13.256 0.116 13.288 ;
  LAYER M1 ;
        RECT 2.816 16.344 2.848 16.416 ;
  LAYER M2 ;
        RECT 2.796 16.364 2.868 16.396 ;
  LAYER M2 ;
        RECT 0.08 16.364 2.832 16.396 ;
  LAYER M1 ;
        RECT 0.064 16.344 0.096 16.416 ;
  LAYER M2 ;
        RECT 0.044 16.364 0.116 16.396 ;
  LAYER M1 ;
        RECT 2.816 19.452 2.848 19.524 ;
  LAYER M2 ;
        RECT 2.796 19.472 2.868 19.504 ;
  LAYER M2 ;
        RECT 0.08 19.472 2.832 19.504 ;
  LAYER M1 ;
        RECT 0.064 19.452 0.096 19.524 ;
  LAYER M2 ;
        RECT 0.044 19.472 0.116 19.504 ;
  LAYER M1 ;
        RECT 2.816 22.56 2.848 22.632 ;
  LAYER M2 ;
        RECT 2.796 22.58 2.868 22.612 ;
  LAYER M2 ;
        RECT 0.08 22.58 2.832 22.612 ;
  LAYER M1 ;
        RECT 0.064 22.56 0.096 22.632 ;
  LAYER M2 ;
        RECT 0.044 22.58 0.116 22.612 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.504 ;
  LAYER M1 ;
        RECT 0.064 0.504 0.096 22.596 ;
  LAYER M1 ;
        RECT 8.768 0.804 8.8 0.876 ;
  LAYER M2 ;
        RECT 8.748 0.824 8.82 0.856 ;
  LAYER M1 ;
        RECT 8.768 0.672 8.8 0.84 ;
  LAYER M1 ;
        RECT 8.768 0.636 8.8 0.708 ;
  LAYER M2 ;
        RECT 8.748 0.656 8.82 0.688 ;
  LAYER M2 ;
        RECT 8.784 0.656 9.008 0.688 ;
  LAYER M1 ;
        RECT 8.992 0.636 9.024 0.708 ;
  LAYER M2 ;
        RECT 8.972 0.656 9.044 0.688 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M1 ;
        RECT 8.768 3.78 8.8 3.948 ;
  LAYER M1 ;
        RECT 8.768 3.744 8.8 3.816 ;
  LAYER M2 ;
        RECT 8.748 3.764 8.82 3.796 ;
  LAYER M2 ;
        RECT 8.784 3.764 9.008 3.796 ;
  LAYER M1 ;
        RECT 8.992 3.744 9.024 3.816 ;
  LAYER M2 ;
        RECT 8.972 3.764 9.044 3.796 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M1 ;
        RECT 8.768 6.888 8.8 7.056 ;
  LAYER M1 ;
        RECT 8.768 6.852 8.8 6.924 ;
  LAYER M2 ;
        RECT 8.748 6.872 8.82 6.904 ;
  LAYER M2 ;
        RECT 8.784 6.872 9.008 6.904 ;
  LAYER M1 ;
        RECT 8.992 6.852 9.024 6.924 ;
  LAYER M2 ;
        RECT 8.972 6.872 9.044 6.904 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M1 ;
        RECT 8.768 9.996 8.8 10.164 ;
  LAYER M1 ;
        RECT 8.768 9.96 8.8 10.032 ;
  LAYER M2 ;
        RECT 8.748 9.98 8.82 10.012 ;
  LAYER M2 ;
        RECT 8.784 9.98 9.008 10.012 ;
  LAYER M1 ;
        RECT 8.992 9.96 9.024 10.032 ;
  LAYER M2 ;
        RECT 8.972 9.98 9.044 10.012 ;
  LAYER M1 ;
        RECT 8.768 13.236 8.8 13.308 ;
  LAYER M2 ;
        RECT 8.748 13.256 8.82 13.288 ;
  LAYER M1 ;
        RECT 8.768 13.104 8.8 13.272 ;
  LAYER M1 ;
        RECT 8.768 13.068 8.8 13.14 ;
  LAYER M2 ;
        RECT 8.748 13.088 8.82 13.12 ;
  LAYER M2 ;
        RECT 8.784 13.088 9.008 13.12 ;
  LAYER M1 ;
        RECT 8.992 13.068 9.024 13.14 ;
  LAYER M2 ;
        RECT 8.972 13.088 9.044 13.12 ;
  LAYER M1 ;
        RECT 8.768 16.344 8.8 16.416 ;
  LAYER M2 ;
        RECT 8.748 16.364 8.82 16.396 ;
  LAYER M1 ;
        RECT 8.768 16.212 8.8 16.38 ;
  LAYER M1 ;
        RECT 8.768 16.176 8.8 16.248 ;
  LAYER M2 ;
        RECT 8.748 16.196 8.82 16.228 ;
  LAYER M2 ;
        RECT 8.784 16.196 9.008 16.228 ;
  LAYER M1 ;
        RECT 8.992 16.176 9.024 16.248 ;
  LAYER M2 ;
        RECT 8.972 16.196 9.044 16.228 ;
  LAYER M1 ;
        RECT 8.768 19.452 8.8 19.524 ;
  LAYER M2 ;
        RECT 8.748 19.472 8.82 19.504 ;
  LAYER M1 ;
        RECT 8.768 19.32 8.8 19.488 ;
  LAYER M1 ;
        RECT 8.768 19.284 8.8 19.356 ;
  LAYER M2 ;
        RECT 8.748 19.304 8.82 19.336 ;
  LAYER M2 ;
        RECT 8.784 19.304 9.008 19.336 ;
  LAYER M1 ;
        RECT 8.992 19.284 9.024 19.356 ;
  LAYER M2 ;
        RECT 8.972 19.304 9.044 19.336 ;
  LAYER M1 ;
        RECT 8.768 22.56 8.8 22.632 ;
  LAYER M2 ;
        RECT 8.748 22.58 8.82 22.612 ;
  LAYER M1 ;
        RECT 8.768 22.428 8.8 22.596 ;
  LAYER M1 ;
        RECT 8.768 22.392 8.8 22.464 ;
  LAYER M2 ;
        RECT 8.748 22.412 8.82 22.444 ;
  LAYER M2 ;
        RECT 8.784 22.412 9.008 22.444 ;
  LAYER M1 ;
        RECT 8.992 22.392 9.024 22.464 ;
  LAYER M2 ;
        RECT 8.972 22.412 9.044 22.444 ;
  LAYER M1 ;
        RECT 8.992 0.048 9.024 0.12 ;
  LAYER M2 ;
        RECT 8.972 0.068 9.044 0.1 ;
  LAYER M1 ;
        RECT 8.992 0.084 9.024 0.504 ;
  LAYER M1 ;
        RECT 8.992 0.504 9.024 22.428 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.008 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.804 5.824 0.876 ;
  LAYER M2 ;
        RECT 5.772 0.824 5.844 0.856 ;
  LAYER M2 ;
        RECT 2.832 0.824 5.808 0.856 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M1 ;
        RECT 5.792 22.56 5.824 22.632 ;
  LAYER M2 ;
        RECT 5.772 22.58 5.844 22.612 ;
  LAYER M2 ;
        RECT 2.832 22.58 5.808 22.612 ;
  LAYER M1 ;
        RECT 2.816 22.56 2.848 22.632 ;
  LAYER M2 ;
        RECT 2.796 22.58 2.868 22.612 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M2 ;
        RECT 3.216 12.584 3.44 12.616 ;
  LAYER M1 ;
        RECT 3.2 12.564 3.232 12.636 ;
  LAYER M2 ;
        RECT 3.18 12.584 3.252 12.616 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M2 ;
        RECT 3.216 15.692 3.44 15.724 ;
  LAYER M1 ;
        RECT 3.2 15.672 3.232 15.744 ;
  LAYER M2 ;
        RECT 3.18 15.692 3.252 15.724 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M2 ;
        RECT 3.216 9.476 3.44 9.508 ;
  LAYER M1 ;
        RECT 3.2 9.456 3.232 9.528 ;
  LAYER M2 ;
        RECT 3.18 9.476 3.252 9.508 ;
  LAYER M1 ;
        RECT 3.424 18.78 3.456 18.852 ;
  LAYER M2 ;
        RECT 3.404 18.8 3.476 18.832 ;
  LAYER M2 ;
        RECT 3.216 18.8 3.44 18.832 ;
  LAYER M1 ;
        RECT 3.2 18.78 3.232 18.852 ;
  LAYER M2 ;
        RECT 3.18 18.8 3.252 18.832 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M2 ;
        RECT 3.216 6.368 3.44 6.4 ;
  LAYER M1 ;
        RECT 3.2 6.348 3.232 6.42 ;
  LAYER M2 ;
        RECT 3.18 6.368 3.252 6.4 ;
  LAYER M1 ;
        RECT 3.424 21.888 3.456 21.96 ;
  LAYER M2 ;
        RECT 3.404 21.908 3.476 21.94 ;
  LAYER M2 ;
        RECT 3.216 21.908 3.44 21.94 ;
  LAYER M1 ;
        RECT 3.2 21.888 3.232 21.96 ;
  LAYER M2 ;
        RECT 3.18 21.908 3.252 21.94 ;
  LAYER M1 ;
        RECT 3.2 25.584 3.232 25.656 ;
  LAYER M2 ;
        RECT 3.18 25.604 3.252 25.636 ;
  LAYER M1 ;
        RECT 3.2 25.368 3.232 25.62 ;
  LAYER M1 ;
        RECT 3.2 6.384 3.232 25.368 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M1 ;
        RECT 3.424 12.6 3.456 12.768 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.44 12.752 6.192 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M1 ;
        RECT 3.424 15.708 3.456 15.876 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 3.44 15.86 6.192 15.892 ;
  LAYER M1 ;
        RECT 6.176 15.84 6.208 15.912 ;
  LAYER M2 ;
        RECT 6.156 15.86 6.228 15.892 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M1 ;
        RECT 3.424 9.492 3.456 9.66 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.44 9.644 6.192 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 3.424 18.78 3.456 18.852 ;
  LAYER M2 ;
        RECT 3.404 18.8 3.476 18.832 ;
  LAYER M1 ;
        RECT 3.424 18.816 3.456 18.984 ;
  LAYER M1 ;
        RECT 3.424 18.948 3.456 19.02 ;
  LAYER M2 ;
        RECT 3.404 18.968 3.476 19 ;
  LAYER M2 ;
        RECT 3.44 18.968 6.192 19 ;
  LAYER M1 ;
        RECT 6.176 18.948 6.208 19.02 ;
  LAYER M2 ;
        RECT 6.156 18.968 6.228 19 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M1 ;
        RECT 3.424 6.384 3.456 6.552 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 3.44 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 3.424 21.888 3.456 21.96 ;
  LAYER M2 ;
        RECT 3.404 21.908 3.476 21.94 ;
  LAYER M1 ;
        RECT 3.424 21.924 3.456 22.092 ;
  LAYER M1 ;
        RECT 3.424 22.056 3.456 22.128 ;
  LAYER M2 ;
        RECT 3.404 22.076 3.476 22.108 ;
  LAYER M2 ;
        RECT 3.44 22.076 6.192 22.108 ;
  LAYER M1 ;
        RECT 6.176 22.056 6.208 22.128 ;
  LAYER M2 ;
        RECT 6.156 22.076 6.228 22.108 ;
  LAYER M1 ;
        RECT 6.176 25.584 6.208 25.656 ;
  LAYER M2 ;
        RECT 6.156 25.604 6.228 25.636 ;
  LAYER M1 ;
        RECT 6.176 25.368 6.208 25.62 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 25.368 ;
  LAYER M2 ;
        RECT 3.216 25.604 6.192 25.636 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M2 ;
        RECT 0.24 3.26 0.464 3.292 ;
  LAYER M1 ;
        RECT 0.224 3.24 0.256 3.312 ;
  LAYER M2 ;
        RECT 0.204 3.26 0.276 3.292 ;
  LAYER M1 ;
        RECT 0.448 6.348 0.48 6.42 ;
  LAYER M2 ;
        RECT 0.428 6.368 0.5 6.4 ;
  LAYER M2 ;
        RECT 0.24 6.368 0.464 6.4 ;
  LAYER M1 ;
        RECT 0.224 6.348 0.256 6.42 ;
  LAYER M2 ;
        RECT 0.204 6.368 0.276 6.4 ;
  LAYER M1 ;
        RECT 0.448 9.456 0.48 9.528 ;
  LAYER M2 ;
        RECT 0.428 9.476 0.5 9.508 ;
  LAYER M2 ;
        RECT 0.24 9.476 0.464 9.508 ;
  LAYER M1 ;
        RECT 0.224 9.456 0.256 9.528 ;
  LAYER M2 ;
        RECT 0.204 9.476 0.276 9.508 ;
  LAYER M1 ;
        RECT 0.448 12.564 0.48 12.636 ;
  LAYER M2 ;
        RECT 0.428 12.584 0.5 12.616 ;
  LAYER M2 ;
        RECT 0.24 12.584 0.464 12.616 ;
  LAYER M1 ;
        RECT 0.224 12.564 0.256 12.636 ;
  LAYER M2 ;
        RECT 0.204 12.584 0.276 12.616 ;
  LAYER M1 ;
        RECT 0.448 15.672 0.48 15.744 ;
  LAYER M2 ;
        RECT 0.428 15.692 0.5 15.724 ;
  LAYER M2 ;
        RECT 0.24 15.692 0.464 15.724 ;
  LAYER M1 ;
        RECT 0.224 15.672 0.256 15.744 ;
  LAYER M2 ;
        RECT 0.204 15.692 0.276 15.724 ;
  LAYER M1 ;
        RECT 0.448 18.78 0.48 18.852 ;
  LAYER M2 ;
        RECT 0.428 18.8 0.5 18.832 ;
  LAYER M2 ;
        RECT 0.24 18.8 0.464 18.832 ;
  LAYER M1 ;
        RECT 0.224 18.78 0.256 18.852 ;
  LAYER M2 ;
        RECT 0.204 18.8 0.276 18.832 ;
  LAYER M1 ;
        RECT 0.448 21.888 0.48 21.96 ;
  LAYER M2 ;
        RECT 0.428 21.908 0.5 21.94 ;
  LAYER M2 ;
        RECT 0.24 21.908 0.464 21.94 ;
  LAYER M1 ;
        RECT 0.224 21.888 0.256 21.96 ;
  LAYER M2 ;
        RECT 0.204 21.908 0.276 21.94 ;
  LAYER M1 ;
        RECT 0.448 24.996 0.48 25.068 ;
  LAYER M2 ;
        RECT 0.428 25.016 0.5 25.048 ;
  LAYER M2 ;
        RECT 0.24 25.016 0.464 25.048 ;
  LAYER M1 ;
        RECT 0.224 24.996 0.256 25.068 ;
  LAYER M2 ;
        RECT 0.204 25.016 0.276 25.048 ;
  LAYER M1 ;
        RECT 0.224 25.752 0.256 25.824 ;
  LAYER M2 ;
        RECT 0.204 25.772 0.276 25.804 ;
  LAYER M1 ;
        RECT 0.224 25.368 0.256 25.788 ;
  LAYER M1 ;
        RECT 0.224 3.276 0.256 25.368 ;
  LAYER M1 ;
        RECT 6.4 3.24 6.432 3.312 ;
  LAYER M2 ;
        RECT 6.38 3.26 6.452 3.292 ;
  LAYER M1 ;
        RECT 6.416 3.26 9.168 3.292 ;
  LAYER M1 ;
        RECT 9.152 3.24 9.184 3.312 ;
  LAYER M2 ;
        RECT 9.132 3.26 9.204 3.292 ;
  LAYER M2 ;
        RECT 9.168 3.26 9.232 3.292 ;
  LAYER M1 ;
        RECT 9.216 3.24 9.248 3.312 ;
  LAYER M2 ;
        RECT 9.196 3.26 9.268 3.292 ;
  LAYER M1 ;
        RECT 6.4 6.348 6.432 6.42 ;
  LAYER M2 ;
        RECT 6.38 6.368 6.452 6.4 ;
  LAYER M1 ;
        RECT 6.416 6.368 9.168 6.4 ;
  LAYER M1 ;
        RECT 9.152 6.348 9.184 6.42 ;
  LAYER M2 ;
        RECT 9.132 6.368 9.204 6.4 ;
  LAYER M2 ;
        RECT 9.168 6.368 9.232 6.4 ;
  LAYER M1 ;
        RECT 9.216 6.348 9.248 6.42 ;
  LAYER M2 ;
        RECT 9.196 6.368 9.268 6.4 ;
  LAYER M1 ;
        RECT 6.4 9.456 6.432 9.528 ;
  LAYER M2 ;
        RECT 6.38 9.476 6.452 9.508 ;
  LAYER M1 ;
        RECT 6.416 9.476 9.168 9.508 ;
  LAYER M1 ;
        RECT 9.152 9.456 9.184 9.528 ;
  LAYER M2 ;
        RECT 9.132 9.476 9.204 9.508 ;
  LAYER M2 ;
        RECT 9.168 9.476 9.232 9.508 ;
  LAYER M1 ;
        RECT 9.216 9.456 9.248 9.528 ;
  LAYER M2 ;
        RECT 9.196 9.476 9.268 9.508 ;
  LAYER M1 ;
        RECT 6.4 12.564 6.432 12.636 ;
  LAYER M2 ;
        RECT 6.38 12.584 6.452 12.616 ;
  LAYER M1 ;
        RECT 6.416 12.584 9.168 12.616 ;
  LAYER M1 ;
        RECT 9.152 12.564 9.184 12.636 ;
  LAYER M2 ;
        RECT 9.132 12.584 9.204 12.616 ;
  LAYER M2 ;
        RECT 9.168 12.584 9.232 12.616 ;
  LAYER M1 ;
        RECT 9.216 12.564 9.248 12.636 ;
  LAYER M2 ;
        RECT 9.196 12.584 9.268 12.616 ;
  LAYER M1 ;
        RECT 6.4 15.672 6.432 15.744 ;
  LAYER M2 ;
        RECT 6.38 15.692 6.452 15.724 ;
  LAYER M1 ;
        RECT 6.416 15.692 9.168 15.724 ;
  LAYER M1 ;
        RECT 9.152 15.672 9.184 15.744 ;
  LAYER M2 ;
        RECT 9.132 15.692 9.204 15.724 ;
  LAYER M2 ;
        RECT 9.168 15.692 9.232 15.724 ;
  LAYER M1 ;
        RECT 9.216 15.672 9.248 15.744 ;
  LAYER M2 ;
        RECT 9.196 15.692 9.268 15.724 ;
  LAYER M1 ;
        RECT 6.4 18.78 6.432 18.852 ;
  LAYER M2 ;
        RECT 6.38 18.8 6.452 18.832 ;
  LAYER M1 ;
        RECT 6.416 18.8 9.168 18.832 ;
  LAYER M1 ;
        RECT 9.152 18.78 9.184 18.852 ;
  LAYER M2 ;
        RECT 9.132 18.8 9.204 18.832 ;
  LAYER M2 ;
        RECT 9.168 18.8 9.232 18.832 ;
  LAYER M1 ;
        RECT 9.216 18.78 9.248 18.852 ;
  LAYER M2 ;
        RECT 9.196 18.8 9.268 18.832 ;
  LAYER M1 ;
        RECT 6.4 21.888 6.432 21.96 ;
  LAYER M2 ;
        RECT 6.38 21.908 6.452 21.94 ;
  LAYER M1 ;
        RECT 6.416 21.908 9.168 21.94 ;
  LAYER M1 ;
        RECT 9.152 21.888 9.184 21.96 ;
  LAYER M2 ;
        RECT 9.132 21.908 9.204 21.94 ;
  LAYER M2 ;
        RECT 9.168 21.908 9.232 21.94 ;
  LAYER M1 ;
        RECT 9.216 21.888 9.248 21.96 ;
  LAYER M2 ;
        RECT 9.196 21.908 9.268 21.94 ;
  LAYER M1 ;
        RECT 6.4 24.996 6.432 25.068 ;
  LAYER M2 ;
        RECT 6.38 25.016 6.452 25.048 ;
  LAYER M1 ;
        RECT 6.416 25.016 9.168 25.048 ;
  LAYER M1 ;
        RECT 9.152 24.996 9.184 25.068 ;
  LAYER M2 ;
        RECT 9.132 25.016 9.204 25.048 ;
  LAYER M2 ;
        RECT 9.168 25.016 9.232 25.048 ;
  LAYER M1 ;
        RECT 9.216 24.996 9.248 25.068 ;
  LAYER M2 ;
        RECT 9.196 25.016 9.268 25.048 ;
  LAYER M1 ;
        RECT 9.216 25.752 9.248 25.824 ;
  LAYER M2 ;
        RECT 9.196 25.772 9.268 25.804 ;
  LAYER M1 ;
        RECT 9.216 25.368 9.248 25.788 ;
  LAYER M1 ;
        RECT 9.216 3.444 9.248 25.368 ;
  LAYER M2 ;
        RECT 0.24 25.772 9.232 25.804 ;
  LAYER M1 ;
        RECT 3.424 3.24 3.456 3.312 ;
  LAYER M2 ;
        RECT 3.404 3.26 3.476 3.292 ;
  LAYER M2 ;
        RECT 0.464 3.26 3.44 3.292 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M1 ;
        RECT 3.424 24.996 3.456 25.068 ;
  LAYER M2 ;
        RECT 3.404 25.016 3.476 25.048 ;
  LAYER M2 ;
        RECT 0.464 25.016 3.44 25.048 ;
  LAYER M1 ;
        RECT 0.448 24.996 0.48 25.068 ;
  LAYER M2 ;
        RECT 0.428 25.016 0.5 25.048 ;
  LAYER M1 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M3 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M1 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M3 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M1 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M3 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M2 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M1 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M3 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M2 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M1 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M3 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M2 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M1 ;
        RECT 0.4 16.296 2.896 18.9 ;
  LAYER M3 ;
        RECT 0.4 16.296 2.896 18.9 ;
  LAYER M2 ;
        RECT 0.4 16.296 2.896 18.9 ;
  LAYER M1 ;
        RECT 0.4 19.404 2.896 22.008 ;
  LAYER M3 ;
        RECT 0.4 19.404 2.896 22.008 ;
  LAYER M2 ;
        RECT 0.4 19.404 2.896 22.008 ;
  LAYER M1 ;
        RECT 0.4 22.512 2.896 25.116 ;
  LAYER M3 ;
        RECT 0.4 22.512 2.896 25.116 ;
  LAYER M2 ;
        RECT 0.4 22.512 2.896 25.116 ;
  LAYER M1 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M3 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M2 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M1 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M3 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M2 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M1 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M3 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M2 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M1 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M3 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M2 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M1 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M3 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M2 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M1 ;
        RECT 3.376 16.296 5.872 18.9 ;
  LAYER M3 ;
        RECT 3.376 16.296 5.872 18.9 ;
  LAYER M2 ;
        RECT 3.376 16.296 5.872 18.9 ;
  LAYER M1 ;
        RECT 3.376 19.404 5.872 22.008 ;
  LAYER M3 ;
        RECT 3.376 19.404 5.872 22.008 ;
  LAYER M2 ;
        RECT 3.376 19.404 5.872 22.008 ;
  LAYER M1 ;
        RECT 3.376 22.512 5.872 25.116 ;
  LAYER M3 ;
        RECT 3.376 22.512 5.872 25.116 ;
  LAYER M2 ;
        RECT 3.376 22.512 5.872 25.116 ;
  LAYER M1 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M3 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M2 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M1 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M3 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M2 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M1 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M3 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M2 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M1 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M3 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M2 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M1 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M3 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M2 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M1 ;
        RECT 6.352 16.296 8.848 18.9 ;
  LAYER M3 ;
        RECT 6.352 16.296 8.848 18.9 ;
  LAYER M2 ;
        RECT 6.352 16.296 8.848 18.9 ;
  LAYER M1 ;
        RECT 6.352 19.404 8.848 22.008 ;
  LAYER M3 ;
        RECT 6.352 19.404 8.848 22.008 ;
  LAYER M2 ;
        RECT 6.352 19.404 8.848 22.008 ;
  LAYER M1 ;
        RECT 6.352 22.512 8.848 25.116 ;
  LAYER M3 ;
        RECT 6.352 22.512 8.848 25.116 ;
  LAYER M2 ;
        RECT 6.352 22.512 8.848 25.116 ;
  END 
END Cap_60fF
