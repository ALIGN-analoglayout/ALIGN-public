MACRO CMC_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.8360 0.1000 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 3.4760 0.2680 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 3.6360 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 3.5560 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER V0 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V0 ;
      RECT 3.4240 0.3620 3.4560 0.3940 ;
    LAYER V0 ;
      RECT 3.4240 0.4880 3.4560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER V0 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V0 ;
      RECT 3.5840 0.3620 3.6160 0.3940 ;
    LAYER V0 ;
      RECT 3.5840 0.4880 3.6160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V1 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.3200 1.0560 0.3520 ;
    LAYER V1 ;
      RECT 2.3040 0.3200 2.3360 0.3520 ;
    LAYER V1 ;
      RECT 3.5840 0.3200 3.6160 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V1 ;
      RECT 2.8640 0.4040 2.8960 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 3.5040 0.4040 3.5360 0.4360 ;
  END
END CMC_NMOS_n12_X3_Y1
MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 1.5560 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 2.2760 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.3200 1.0560 0.3520 ;
    LAYER V1 ;
      RECT 1.5040 0.3200 1.5360 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
  END
END CMC_PMOS_n12_X2_Y1
MACRO CMC_PMOS_S_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 0.4360 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 1.0760 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 0.9960 0.3520 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
  END
END CMC_PMOS_S_n12_X1_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 1.0760 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DP_NMOS_n12_X3_Y3
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X3_Y3 0 0 ;
  SIZE 3.8400 BY 2.5200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 3.4760 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 3.4760 0.9400 ;
      LAYER M2 ;
        RECT 0.2040 1.7480 3.4760 1.7800 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
      LAYER M2 ;
        RECT 1.0040 0.9920 3.6360 1.0240 ;
      LAYER M2 ;
        RECT 0.3640 1.8320 2.9960 1.8640 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 3.6360 0.2680 ;
      LAYER M2 ;
        RECT 0.3640 1.0760 2.9960 1.1080 ;
      LAYER M2 ;
        RECT 1.0040 1.9160 3.6360 1.9480 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 2.9160 0.3520 ;
      LAYER M2 ;
        RECT 0.9240 1.1600 3.5560 1.1920 ;
      LAYER M2 ;
        RECT 0.2840 2.0000 2.9160 2.0320 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4040 3.5560 0.4360 ;
      LAYER M2 ;
        RECT 0.2840 1.2440 2.9160 1.2760 ;
      LAYER M2 ;
        RECT 0.9240 2.0840 3.5560 2.1160 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER V0 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V0 ;
      RECT 3.4240 0.3620 3.4560 0.3940 ;
    LAYER V0 ;
      RECT 3.4240 0.4880 3.4560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER V0 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V0 ;
      RECT 3.5840 0.3620 3.6160 0.3940 ;
    LAYER V0 ;
      RECT 3.5840 0.4880 3.6160 0.5200 ;
    LAYER M3 ;
      RECT 1.8200 0.0480 1.8600 0.1200 ;
    LAYER V2 ;
      RECT 1.8200 0.0680 1.8600 0.1000 ;
    LAYER V2 ;
      RECT 1.8200 0.0680 1.8600 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 3.4240 0.0680 3.4560 0.1000 ;
    LAYER M3 ;
      RECT 1.7400 0.1320 1.7800 0.2040 ;
    LAYER V2 ;
      RECT 1.7400 0.1520 1.7800 0.1840 ;
    LAYER V2 ;
      RECT 1.7400 0.1520 1.7800 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER M3 ;
      RECT 1.9000 0.2160 1.9400 0.2880 ;
    LAYER V2 ;
      RECT 1.9000 0.2360 1.9400 0.2680 ;
    LAYER V2 ;
      RECT 1.9000 0.2360 1.9400 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V1 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER M3 ;
      RECT 1.6600 0.3000 1.7000 0.3720 ;
    LAYER V2 ;
      RECT 1.6600 0.3200 1.7000 0.3520 ;
    LAYER V2 ;
      RECT 1.6600 0.3200 1.7000 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 1.5840 0.3200 1.6160 0.3520 ;
    LAYER V1 ;
      RECT 2.8640 0.3200 2.8960 0.3520 ;
    LAYER M3 ;
      RECT 1.9800 0.3840 2.0200 0.4560 ;
    LAYER V2 ;
      RECT 1.9800 0.4040 2.0200 0.4360 ;
    LAYER V2 ;
      RECT 1.9800 0.4040 2.0200 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 3.5040 0.4040 3.5360 0.4360 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 3.5040 0.8880 3.5360 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER V0 ;
      RECT 2.7840 1.0760 2.8160 1.1080 ;
    LAYER V0 ;
      RECT 2.7840 1.2020 2.8160 1.2340 ;
    LAYER V0 ;
      RECT 2.7840 1.3280 2.8160 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER V0 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER V0 ;
      RECT 2.1440 1.2020 2.1760 1.2340 ;
    LAYER V0 ;
      RECT 2.1440 1.3280 2.1760 1.3600 ;
    LAYER M1 ;
      RECT 3.4240 0.8880 3.4560 1.5480 ;
    LAYER V0 ;
      RECT 3.4240 1.0760 3.4560 1.1080 ;
    LAYER V0 ;
      RECT 3.4240 1.2020 3.4560 1.2340 ;
    LAYER V0 ;
      RECT 3.4240 1.3280 3.4560 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER V0 ;
      RECT 2.9440 1.0760 2.9760 1.1080 ;
    LAYER V0 ;
      RECT 2.9440 1.2020 2.9760 1.2340 ;
    LAYER V0 ;
      RECT 2.9440 1.3280 2.9760 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER V0 ;
      RECT 2.3040 1.0760 2.3360 1.1080 ;
    LAYER V0 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER V0 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER M1 ;
      RECT 3.5840 0.8880 3.6160 1.5480 ;
    LAYER V0 ;
      RECT 3.5840 1.0760 3.6160 1.1080 ;
    LAYER V0 ;
      RECT 3.5840 1.2020 3.6160 1.2340 ;
    LAYER V0 ;
      RECT 3.5840 1.3280 3.6160 1.3600 ;
    LAYER M3 ;
      RECT 1.8200 0.0480 1.8600 0.9600 ;
    LAYER V2 ;
      RECT 1.8200 0.0680 1.8600 0.1000 ;
    LAYER V2 ;
      RECT 1.8200 0.9080 1.8600 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 1.5040 0.9080 1.5360 0.9400 ;
    LAYER V1 ;
      RECT 2.7840 0.9080 2.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 2.1440 0.9080 2.1760 0.9400 ;
    LAYER V1 ;
      RECT 3.4240 0.9080 3.4560 0.9400 ;
    LAYER M3 ;
      RECT 1.7400 0.1320 1.7800 1.0440 ;
    LAYER V2 ;
      RECT 1.7400 0.1520 1.7800 0.1840 ;
    LAYER V2 ;
      RECT 1.7400 0.9920 1.7800 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 2.3040 0.9920 2.3360 1.0240 ;
    LAYER V1 ;
      RECT 3.5840 0.9920 3.6160 1.0240 ;
    LAYER M3 ;
      RECT 1.9000 0.2160 1.9400 1.1280 ;
    LAYER V2 ;
      RECT 1.9000 0.2360 1.9400 0.2680 ;
    LAYER V2 ;
      RECT 1.9000 1.0760 1.9400 1.1080 ;
    LAYER V1 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V1 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V1 ;
      RECT 2.9440 1.0760 2.9760 1.1080 ;
    LAYER M3 ;
      RECT 1.6600 0.3000 1.7000 1.2120 ;
    LAYER V2 ;
      RECT 1.6600 0.3200 1.7000 0.3520 ;
    LAYER V2 ;
      RECT 1.6600 1.1600 1.7000 1.1920 ;
    LAYER V1 ;
      RECT 0.9440 1.1600 0.9760 1.1920 ;
    LAYER V1 ;
      RECT 2.2240 1.1600 2.2560 1.1920 ;
    LAYER V1 ;
      RECT 3.5040 1.1600 3.5360 1.1920 ;
    LAYER M3 ;
      RECT 1.9800 0.3840 2.0200 1.2960 ;
    LAYER V2 ;
      RECT 1.9800 0.4040 2.0200 0.4360 ;
    LAYER V2 ;
      RECT 1.9800 1.2440 2.0200 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V1 ;
      RECT 1.5840 1.2440 1.6160 1.2760 ;
    LAYER V1 ;
      RECT 2.8640 1.2440 2.8960 1.2760 ;
    LAYER M1 ;
      RECT 0.3040 1.7280 0.3360 2.3880 ;
    LAYER M1 ;
      RECT 1.5840 1.7280 1.6160 2.3880 ;
    LAYER M1 ;
      RECT 2.8640 1.7280 2.8960 2.3880 ;
    LAYER M1 ;
      RECT 0.9440 1.7280 0.9760 2.3880 ;
    LAYER M1 ;
      RECT 2.2240 1.7280 2.2560 2.3880 ;
    LAYER M1 ;
      RECT 3.5040 1.7280 3.5360 2.3880 ;
    LAYER M1 ;
      RECT 0.2240 1.7280 0.2560 2.3880 ;
    LAYER V0 ;
      RECT 0.2240 1.9160 0.2560 1.9480 ;
    LAYER V0 ;
      RECT 0.2240 2.0420 0.2560 2.0740 ;
    LAYER V0 ;
      RECT 0.2240 2.1680 0.2560 2.2000 ;
    LAYER M1 ;
      RECT 1.5040 1.7280 1.5360 2.3880 ;
    LAYER V0 ;
      RECT 1.5040 1.9160 1.5360 1.9480 ;
    LAYER V0 ;
      RECT 1.5040 2.0420 1.5360 2.0740 ;
    LAYER V0 ;
      RECT 1.5040 2.1680 1.5360 2.2000 ;
    LAYER M1 ;
      RECT 2.7840 1.7280 2.8160 2.3880 ;
    LAYER V0 ;
      RECT 2.7840 1.9160 2.8160 1.9480 ;
    LAYER V0 ;
      RECT 2.7840 2.0420 2.8160 2.0740 ;
    LAYER V0 ;
      RECT 2.7840 2.1680 2.8160 2.2000 ;
    LAYER M1 ;
      RECT 0.8640 1.7280 0.8960 2.3880 ;
    LAYER V0 ;
      RECT 0.8640 1.9160 0.8960 1.9480 ;
    LAYER V0 ;
      RECT 0.8640 2.0420 0.8960 2.0740 ;
    LAYER V0 ;
      RECT 0.8640 2.1680 0.8960 2.2000 ;
    LAYER M1 ;
      RECT 2.1440 1.7280 2.1760 2.3880 ;
    LAYER V0 ;
      RECT 2.1440 1.9160 2.1760 1.9480 ;
    LAYER V0 ;
      RECT 2.1440 2.0420 2.1760 2.0740 ;
    LAYER V0 ;
      RECT 2.1440 2.1680 2.1760 2.2000 ;
    LAYER M1 ;
      RECT 3.4240 1.7280 3.4560 2.3880 ;
    LAYER V0 ;
      RECT 3.4240 1.9160 3.4560 1.9480 ;
    LAYER V0 ;
      RECT 3.4240 2.0420 3.4560 2.0740 ;
    LAYER V0 ;
      RECT 3.4240 2.1680 3.4560 2.2000 ;
    LAYER M1 ;
      RECT 0.3840 1.7280 0.4160 2.3880 ;
    LAYER V0 ;
      RECT 0.3840 1.9160 0.4160 1.9480 ;
    LAYER V0 ;
      RECT 0.3840 2.0420 0.4160 2.0740 ;
    LAYER V0 ;
      RECT 0.3840 2.1680 0.4160 2.2000 ;
    LAYER M1 ;
      RECT 1.6640 1.7280 1.6960 2.3880 ;
    LAYER V0 ;
      RECT 1.6640 1.9160 1.6960 1.9480 ;
    LAYER V0 ;
      RECT 1.6640 2.0420 1.6960 2.0740 ;
    LAYER V0 ;
      RECT 1.6640 2.1680 1.6960 2.2000 ;
    LAYER M1 ;
      RECT 2.9440 1.7280 2.9760 2.3880 ;
    LAYER V0 ;
      RECT 2.9440 1.9160 2.9760 1.9480 ;
    LAYER V0 ;
      RECT 2.9440 2.0420 2.9760 2.0740 ;
    LAYER V0 ;
      RECT 2.9440 2.1680 2.9760 2.2000 ;
    LAYER M1 ;
      RECT 1.0240 1.7280 1.0560 2.3880 ;
    LAYER V0 ;
      RECT 1.0240 1.9160 1.0560 1.9480 ;
    LAYER V0 ;
      RECT 1.0240 2.0420 1.0560 2.0740 ;
    LAYER V0 ;
      RECT 1.0240 2.1680 1.0560 2.2000 ;
    LAYER M1 ;
      RECT 2.3040 1.7280 2.3360 2.3880 ;
    LAYER V0 ;
      RECT 2.3040 1.9160 2.3360 1.9480 ;
    LAYER V0 ;
      RECT 2.3040 2.0420 2.3360 2.0740 ;
    LAYER V0 ;
      RECT 2.3040 2.1680 2.3360 2.2000 ;
    LAYER M1 ;
      RECT 3.5840 1.7280 3.6160 2.3880 ;
    LAYER V0 ;
      RECT 3.5840 1.9160 3.6160 1.9480 ;
    LAYER V0 ;
      RECT 3.5840 2.0420 3.6160 2.0740 ;
    LAYER V0 ;
      RECT 3.5840 2.1680 3.6160 2.2000 ;
    LAYER M3 ;
      RECT 1.8200 0.0480 1.8600 1.8000 ;
    LAYER V2 ;
      RECT 1.8200 0.0680 1.8600 0.1000 ;
    LAYER V2 ;
      RECT 1.8200 1.7480 1.8600 1.7800 ;
    LAYER V1 ;
      RECT 0.2240 1.7480 0.2560 1.7800 ;
    LAYER V1 ;
      RECT 1.5040 1.7480 1.5360 1.7800 ;
    LAYER V1 ;
      RECT 2.7840 1.7480 2.8160 1.7800 ;
    LAYER V1 ;
      RECT 0.8640 1.7480 0.8960 1.7800 ;
    LAYER V1 ;
      RECT 2.1440 1.7480 2.1760 1.7800 ;
    LAYER V1 ;
      RECT 3.4240 1.7480 3.4560 1.7800 ;
    LAYER M3 ;
      RECT 1.7400 0.1320 1.7800 1.8840 ;
    LAYER V2 ;
      RECT 1.7400 0.1520 1.7800 0.1840 ;
    LAYER V2 ;
      RECT 1.7400 1.8320 1.7800 1.8640 ;
    LAYER V1 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V1 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V1 ;
      RECT 2.9440 1.8320 2.9760 1.8640 ;
    LAYER M3 ;
      RECT 1.9000 0.2160 1.9400 1.9680 ;
    LAYER V2 ;
      RECT 1.9000 0.2360 1.9400 0.2680 ;
    LAYER V2 ;
      RECT 1.9000 1.9160 1.9400 1.9480 ;
    LAYER V1 ;
      RECT 1.0240 1.9160 1.0560 1.9480 ;
    LAYER V1 ;
      RECT 2.3040 1.9160 2.3360 1.9480 ;
    LAYER V1 ;
      RECT 3.5840 1.9160 3.6160 1.9480 ;
    LAYER M3 ;
      RECT 1.6600 0.3000 1.7000 2.0520 ;
    LAYER V2 ;
      RECT 1.6600 0.3200 1.7000 0.3520 ;
    LAYER V2 ;
      RECT 1.6600 2.0000 1.7000 2.0320 ;
    LAYER V1 ;
      RECT 0.3040 2.0000 0.3360 2.0320 ;
    LAYER V1 ;
      RECT 1.5840 2.0000 1.6160 2.0320 ;
    LAYER V1 ;
      RECT 2.8640 2.0000 2.8960 2.0320 ;
    LAYER M3 ;
      RECT 1.9800 0.3840 2.0200 2.1360 ;
    LAYER V2 ;
      RECT 1.9800 0.4040 2.0200 0.4360 ;
    LAYER V2 ;
      RECT 1.9800 2.0840 2.0200 2.1160 ;
    LAYER V1 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V1 ;
      RECT 2.2240 2.0840 2.2560 2.1160 ;
    LAYER V1 ;
      RECT 3.5040 2.0840 3.5360 2.1160 ;
  END
END DP_NMOS_n12_X3_Y3
MACRO Switch_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y1 0 0 ;
  SIZE 1.9200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.5560 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 1.6360 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.7160 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
  END
END Switch_NMOS_n12_X3_Y1
MACRO Switch_NMOS_n12_X3_Y3
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y3 0 0 ;
  SIZE 1.9200 BY 2.5200 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.5560 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 1.5560 0.9400 ;
      LAYER M2 ;
        RECT 0.2040 1.7480 1.5560 1.7800 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 1.6360 0.2680 ;
      LAYER M2 ;
        RECT 0.2840 1.0760 1.6360 1.1080 ;
      LAYER M2 ;
        RECT 0.2840 1.9160 1.6360 1.9480 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.7160 0.1840 ;
      LAYER M2 ;
        RECT 0.3640 0.9920 1.7160 1.0240 ;
      LAYER M2 ;
        RECT 0.3640 1.8320 1.7160 1.8640 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M3 ;
      RECT 0.8600 0.0480 0.9000 0.1200 ;
    LAYER V2 ;
      RECT 0.8600 0.0680 0.9000 0.1000 ;
    LAYER V2 ;
      RECT 0.8600 0.0680 0.9000 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER M3 ;
      RECT 0.9400 0.1320 0.9800 0.2040 ;
    LAYER V2 ;
      RECT 0.9400 0.1520 0.9800 0.1840 ;
    LAYER V2 ;
      RECT 0.9400 0.1520 0.9800 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER M3 ;
      RECT 0.7800 0.2160 0.8200 0.2880 ;
    LAYER V2 ;
      RECT 0.7800 0.2360 0.8200 0.2680 ;
    LAYER V2 ;
      RECT 0.7800 0.2360 0.8200 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M3 ;
      RECT 0.8600 0.0480 0.9000 0.9600 ;
    LAYER V2 ;
      RECT 0.8600 0.0680 0.9000 0.1000 ;
    LAYER V2 ;
      RECT 0.8600 0.9080 0.9000 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 1.5040 0.9080 1.5360 0.9400 ;
    LAYER M3 ;
      RECT 0.9400 0.1320 0.9800 1.0440 ;
    LAYER V2 ;
      RECT 0.9400 0.1520 0.9800 0.1840 ;
    LAYER V2 ;
      RECT 0.9400 0.9920 0.9800 1.0240 ;
    LAYER V1 ;
      RECT 0.3840 0.9920 0.4160 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.6640 0.9920 1.6960 1.0240 ;
    LAYER M3 ;
      RECT 0.7800 0.2160 0.8200 1.1280 ;
    LAYER V2 ;
      RECT 0.7800 0.2360 0.8200 0.2680 ;
    LAYER V2 ;
      RECT 0.7800 1.0760 0.8200 1.1080 ;
    LAYER V1 ;
      RECT 0.3040 1.0760 0.3360 1.1080 ;
    LAYER V1 ;
      RECT 0.9440 1.0760 0.9760 1.1080 ;
    LAYER V1 ;
      RECT 1.5840 1.0760 1.6160 1.1080 ;
    LAYER M1 ;
      RECT 0.3040 1.7280 0.3360 2.3880 ;
    LAYER M1 ;
      RECT 0.9440 1.7280 0.9760 2.3880 ;
    LAYER M1 ;
      RECT 1.5840 1.7280 1.6160 2.3880 ;
    LAYER M1 ;
      RECT 0.2240 1.7280 0.2560 2.3880 ;
    LAYER V0 ;
      RECT 0.2240 1.9160 0.2560 1.9480 ;
    LAYER V0 ;
      RECT 0.2240 2.0420 0.2560 2.0740 ;
    LAYER V0 ;
      RECT 0.2240 2.1680 0.2560 2.2000 ;
    LAYER M1 ;
      RECT 0.8640 1.7280 0.8960 2.3880 ;
    LAYER V0 ;
      RECT 0.8640 1.9160 0.8960 1.9480 ;
    LAYER V0 ;
      RECT 0.8640 2.0420 0.8960 2.0740 ;
    LAYER V0 ;
      RECT 0.8640 2.1680 0.8960 2.2000 ;
    LAYER M1 ;
      RECT 1.5040 1.7280 1.5360 2.3880 ;
    LAYER V0 ;
      RECT 1.5040 1.9160 1.5360 1.9480 ;
    LAYER V0 ;
      RECT 1.5040 2.0420 1.5360 2.0740 ;
    LAYER V0 ;
      RECT 1.5040 2.1680 1.5360 2.2000 ;
    LAYER M1 ;
      RECT 0.3840 1.7280 0.4160 2.3880 ;
    LAYER V0 ;
      RECT 0.3840 1.9160 0.4160 1.9480 ;
    LAYER V0 ;
      RECT 0.3840 2.0420 0.4160 2.0740 ;
    LAYER V0 ;
      RECT 0.3840 2.1680 0.4160 2.2000 ;
    LAYER M1 ;
      RECT 1.0240 1.7280 1.0560 2.3880 ;
    LAYER V0 ;
      RECT 1.0240 1.9160 1.0560 1.9480 ;
    LAYER V0 ;
      RECT 1.0240 2.0420 1.0560 2.0740 ;
    LAYER V0 ;
      RECT 1.0240 2.1680 1.0560 2.2000 ;
    LAYER M1 ;
      RECT 1.6640 1.7280 1.6960 2.3880 ;
    LAYER V0 ;
      RECT 1.6640 1.9160 1.6960 1.9480 ;
    LAYER V0 ;
      RECT 1.6640 2.0420 1.6960 2.0740 ;
    LAYER V0 ;
      RECT 1.6640 2.1680 1.6960 2.2000 ;
    LAYER M3 ;
      RECT 0.8600 0.0480 0.9000 1.8000 ;
    LAYER V2 ;
      RECT 0.8600 0.0680 0.9000 0.1000 ;
    LAYER V2 ;
      RECT 0.8600 1.7480 0.9000 1.7800 ;
    LAYER V1 ;
      RECT 0.2240 1.7480 0.2560 1.7800 ;
    LAYER V1 ;
      RECT 0.8640 1.7480 0.8960 1.7800 ;
    LAYER V1 ;
      RECT 1.5040 1.7480 1.5360 1.7800 ;
    LAYER M3 ;
      RECT 0.9400 0.1320 0.9800 1.8840 ;
    LAYER V2 ;
      RECT 0.9400 0.1520 0.9800 0.1840 ;
    LAYER V2 ;
      RECT 0.9400 1.8320 0.9800 1.8640 ;
    LAYER V1 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V1 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V1 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER M3 ;
      RECT 0.7800 0.2160 0.8200 1.9680 ;
    LAYER V2 ;
      RECT 0.7800 0.2360 0.8200 0.2680 ;
    LAYER V2 ;
      RECT 0.7800 1.9160 0.8200 1.9480 ;
    LAYER V1 ;
      RECT 0.3040 1.9160 0.3360 1.9480 ;
    LAYER V1 ;
      RECT 0.9440 1.9160 0.9760 1.9480 ;
    LAYER V1 ;
      RECT 1.5840 1.9160 1.6160 1.9480 ;
  END
END Switch_NMOS_n12_X3_Y3
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.2760 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.3560 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 0.4360 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.9960 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.0760 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
  END
END Switch_PMOS_n12_X2_Y1
MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 2.5600 BY 1.6800 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 2.3560 0.9400 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
      LAYER M2 ;
        RECT 1.0040 0.9920 1.5560 1.0240 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 1.5560 0.2680 ;
      LAYER M2 ;
        RECT 0.3640 1.0760 2.1960 1.1080 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 2.2760 0.3520 ;
      LAYER M2 ;
        RECT 0.9240 1.1600 1.6360 1.1920 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4040 1.6360 0.4360 ;
      LAYER M2 ;
        RECT 0.2840 1.2440 2.2760 1.2760 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M3 ;
      RECT 1.2600 0.0480 1.3000 0.1200 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER M3 ;
      RECT 1.1800 0.1320 1.2200 0.2040 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER M3 ;
      RECT 1.3400 0.2160 1.3800 0.2880 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER M3 ;
      RECT 1.1000 0.3000 1.1400 0.3720 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 2.2240 0.3200 2.2560 0.3520 ;
    LAYER M3 ;
      RECT 1.4200 0.3840 1.4600 0.4560 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER V0 ;
      RECT 2.3040 1.0760 2.3360 1.1080 ;
    LAYER V0 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER V0 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER V0 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER V0 ;
      RECT 2.1440 1.2020 2.1760 1.2340 ;
    LAYER V0 ;
      RECT 2.1440 1.3280 2.1760 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M3 ;
      RECT 1.2600 0.0480 1.3000 0.9600 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V2 ;
      RECT 1.2600 0.9080 1.3000 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.3040 0.9080 2.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER M3 ;
      RECT 1.1800 0.1320 1.2200 1.0440 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V2 ;
      RECT 1.1800 0.9920 1.2200 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.5040 0.9920 1.5360 1.0240 ;
    LAYER M3 ;
      RECT 1.3400 0.2160 1.3800 1.1280 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V2 ;
      RECT 1.3400 1.0760 1.3800 1.1080 ;
    LAYER V1 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V1 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER M3 ;
      RECT 1.1000 0.3000 1.1400 1.2120 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V2 ;
      RECT 1.1000 1.1600 1.1400 1.1920 ;
    LAYER V1 ;
      RECT 0.9440 1.1600 0.9760 1.1920 ;
    LAYER V1 ;
      RECT 1.5840 1.1600 1.6160 1.1920 ;
    LAYER M3 ;
      RECT 1.4200 0.3840 1.4600 1.2960 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V2 ;
      RECT 1.4200 1.2440 1.4600 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V1 ;
      RECT 2.2240 1.2440 2.2560 1.2760 ;
  END
END test
