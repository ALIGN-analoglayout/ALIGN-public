.model n nmos nfin=1 w=1 nf=1 l=1 m=1
.model p pmos nfin=1 w=1 nf=1 l=1 m=1
.model nlvt nmos nfin=1 w=1 nf=1 l=1 m=1
.model plvt pmos nfin=1 w=1 nf=1 l=1 m=1
.model npv nmos nfin=1 w=1 nf=1 l=1 m=1 source=sig drain=sig dv=0
.model ppv pmos nfin=1 w=1 nf=1 l=1 m=1 source=sig drain=sig dv=0
.model tfr_flat tfr w=1 l=1
.model tfr_prim tfr w=1 l=1
