MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 14.72 BY 16.044 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.984 15.588 6.016 15.66 ;
      LAYER M2 ;
        RECT 5.964 15.608 6.036 15.64 ;
      LAYER M1 ;
        RECT 8.864 15.588 8.896 15.66 ;
      LAYER M2 ;
        RECT 8.844 15.608 8.916 15.64 ;
      LAYER M2 ;
        RECT 6 15.608 8.88 15.64 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
      LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
      LAYER M1 ;
        RECT 8.704 0.384 8.736 0.456 ;
      LAYER M2 ;
        RECT 8.684 0.404 8.756 0.436 ;
      LAYER M2 ;
        RECT 5.84 0.404 8.72 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 15.756 3.136 15.828 ;
      LAYER M2 ;
        RECT 3.084 15.776 3.156 15.808 ;
      LAYER M1 ;
        RECT 11.744 15.756 11.776 15.828 ;
      LAYER M2 ;
        RECT 11.724 15.776 11.796 15.808 ;
      LAYER M2 ;
        RECT 3.12 15.776 11.76 15.808 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
      LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
      LAYER M1 ;
        RECT 11.584 0.216 11.616 0.288 ;
      LAYER M2 ;
        RECT 11.564 0.236 11.636 0.268 ;
      LAYER M2 ;
        RECT 2.96 0.236 11.6 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.544 6.768 8.576 6.84 ;
  LAYER M2 ;
        RECT 8.524 6.788 8.596 6.82 ;
  LAYER M2 ;
        RECT 5.84 6.788 8.56 6.82 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 6.84 ;
  LAYER M2 ;
        RECT 5.804 6.788 5.876 6.82 ;
  LAYER M1 ;
        RECT 5.664 9.708 5.696 9.78 ;
  LAYER M2 ;
        RECT 5.644 9.728 5.716 9.76 ;
  LAYER M1 ;
        RECT 5.664 9.576 5.696 9.744 ;
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M2 ;
        RECT 5.68 9.56 5.84 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
  LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 0.588 ;
  LAYER M1 ;
        RECT 5.824 0.588 5.856 9.576 ;
  LAYER M1 ;
        RECT 11.424 3.828 11.456 3.9 ;
  LAYER M2 ;
        RECT 11.404 3.848 11.476 3.88 ;
  LAYER M2 ;
        RECT 8.72 3.848 11.44 3.88 ;
  LAYER M1 ;
        RECT 8.704 3.828 8.736 3.9 ;
  LAYER M2 ;
        RECT 8.684 3.848 8.756 3.88 ;
  LAYER M1 ;
        RECT 8.704 0.384 8.736 0.456 ;
  LAYER M2 ;
        RECT 8.684 0.404 8.756 0.436 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 0.588 ;
  LAYER M1 ;
        RECT 8.704 0.588 8.736 3.864 ;
  LAYER M2 ;
        RECT 5.84 0.404 8.72 0.436 ;
  LAYER M1 ;
        RECT 5.664 6.768 5.696 6.84 ;
  LAYER M2 ;
        RECT 5.644 6.788 5.716 6.82 ;
  LAYER M2 ;
        RECT 2.96 6.788 5.68 6.82 ;
  LAYER M1 ;
        RECT 2.944 6.768 2.976 6.84 ;
  LAYER M2 ;
        RECT 2.924 6.788 2.996 6.82 ;
  LAYER M1 ;
        RECT 5.664 3.828 5.696 3.9 ;
  LAYER M2 ;
        RECT 5.644 3.848 5.716 3.88 ;
  LAYER M2 ;
        RECT 2.96 3.848 5.68 3.88 ;
  LAYER M1 ;
        RECT 2.944 3.828 2.976 3.9 ;
  LAYER M2 ;
        RECT 2.924 3.848 2.996 3.88 ;
  LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
  LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
  LAYER M1 ;
        RECT 2.944 0.252 2.976 0.588 ;
  LAYER M1 ;
        RECT 2.944 0.588 2.976 6.804 ;
  LAYER M1 ;
        RECT 11.424 6.768 11.456 6.84 ;
  LAYER M2 ;
        RECT 11.404 6.788 11.476 6.82 ;
  LAYER M1 ;
        RECT 11.424 6.636 11.456 6.804 ;
  LAYER M1 ;
        RECT 11.424 6.6 11.456 6.672 ;
  LAYER M2 ;
        RECT 11.404 6.62 11.476 6.652 ;
  LAYER M2 ;
        RECT 11.44 6.62 11.6 6.652 ;
  LAYER M1 ;
        RECT 11.584 6.6 11.616 6.672 ;
  LAYER M2 ;
        RECT 11.564 6.62 11.636 6.652 ;
  LAYER M1 ;
        RECT 11.424 9.708 11.456 9.78 ;
  LAYER M2 ;
        RECT 11.404 9.728 11.476 9.76 ;
  LAYER M1 ;
        RECT 11.424 9.576 11.456 9.744 ;
  LAYER M1 ;
        RECT 11.424 9.54 11.456 9.612 ;
  LAYER M2 ;
        RECT 11.404 9.56 11.476 9.592 ;
  LAYER M2 ;
        RECT 11.44 9.56 11.6 9.592 ;
  LAYER M1 ;
        RECT 11.584 9.54 11.616 9.612 ;
  LAYER M2 ;
        RECT 11.564 9.56 11.636 9.592 ;
  LAYER M1 ;
        RECT 11.584 0.216 11.616 0.288 ;
  LAYER M2 ;
        RECT 11.564 0.236 11.636 0.268 ;
  LAYER M1 ;
        RECT 11.584 0.252 11.616 0.588 ;
  LAYER M1 ;
        RECT 11.584 0.588 11.616 9.576 ;
  LAYER M2 ;
        RECT 2.96 0.236 11.6 0.268 ;
  LAYER M1 ;
        RECT 8.544 3.828 8.576 3.9 ;
  LAYER M2 ;
        RECT 8.524 3.848 8.596 3.88 ;
  LAYER M2 ;
        RECT 5.68 3.848 8.56 3.88 ;
  LAYER M1 ;
        RECT 5.664 3.828 5.696 3.9 ;
  LAYER M2 ;
        RECT 5.644 3.848 5.716 3.88 ;
  LAYER M1 ;
        RECT 8.544 9.708 8.576 9.78 ;
  LAYER M2 ;
        RECT 8.524 9.728 8.596 9.76 ;
  LAYER M2 ;
        RECT 8.56 9.728 11.44 9.76 ;
  LAYER M1 ;
        RECT 11.424 9.708 11.456 9.78 ;
  LAYER M2 ;
        RECT 11.404 9.728 11.476 9.76 ;
  LAYER M1 ;
        RECT 2.784 0.888 2.816 0.96 ;
  LAYER M2 ;
        RECT 2.764 0.908 2.836 0.94 ;
  LAYER M2 ;
        RECT 0.08 0.908 2.8 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 2.784 3.828 2.816 3.9 ;
  LAYER M2 ;
        RECT 2.764 3.848 2.836 3.88 ;
  LAYER M2 ;
        RECT 0.08 3.848 2.8 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 2.784 6.768 2.816 6.84 ;
  LAYER M2 ;
        RECT 2.764 6.788 2.836 6.82 ;
  LAYER M2 ;
        RECT 0.08 6.788 2.8 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 2.784 9.708 2.816 9.78 ;
  LAYER M2 ;
        RECT 2.764 9.728 2.836 9.76 ;
  LAYER M2 ;
        RECT 0.08 9.728 2.8 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 2.784 12.648 2.816 12.72 ;
  LAYER M2 ;
        RECT 2.764 12.668 2.836 12.7 ;
  LAYER M2 ;
        RECT 0.08 12.668 2.8 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.588 ;
  LAYER M1 ;
        RECT 0.064 0.588 0.096 12.684 ;
  LAYER M1 ;
        RECT 14.304 0.888 14.336 0.96 ;
  LAYER M2 ;
        RECT 14.284 0.908 14.356 0.94 ;
  LAYER M1 ;
        RECT 14.304 0.756 14.336 0.924 ;
  LAYER M1 ;
        RECT 14.304 0.72 14.336 0.792 ;
  LAYER M2 ;
        RECT 14.284 0.74 14.356 0.772 ;
  LAYER M2 ;
        RECT 14.32 0.74 14.48 0.772 ;
  LAYER M1 ;
        RECT 14.464 0.72 14.496 0.792 ;
  LAYER M2 ;
        RECT 14.444 0.74 14.516 0.772 ;
  LAYER M1 ;
        RECT 14.304 3.828 14.336 3.9 ;
  LAYER M2 ;
        RECT 14.284 3.848 14.356 3.88 ;
  LAYER M1 ;
        RECT 14.304 3.696 14.336 3.864 ;
  LAYER M1 ;
        RECT 14.304 3.66 14.336 3.732 ;
  LAYER M2 ;
        RECT 14.284 3.68 14.356 3.712 ;
  LAYER M2 ;
        RECT 14.32 3.68 14.48 3.712 ;
  LAYER M1 ;
        RECT 14.464 3.66 14.496 3.732 ;
  LAYER M2 ;
        RECT 14.444 3.68 14.516 3.712 ;
  LAYER M1 ;
        RECT 14.304 6.768 14.336 6.84 ;
  LAYER M2 ;
        RECT 14.284 6.788 14.356 6.82 ;
  LAYER M1 ;
        RECT 14.304 6.636 14.336 6.804 ;
  LAYER M1 ;
        RECT 14.304 6.6 14.336 6.672 ;
  LAYER M2 ;
        RECT 14.284 6.62 14.356 6.652 ;
  LAYER M2 ;
        RECT 14.32 6.62 14.48 6.652 ;
  LAYER M1 ;
        RECT 14.464 6.6 14.496 6.672 ;
  LAYER M2 ;
        RECT 14.444 6.62 14.516 6.652 ;
  LAYER M1 ;
        RECT 14.304 9.708 14.336 9.78 ;
  LAYER M2 ;
        RECT 14.284 9.728 14.356 9.76 ;
  LAYER M1 ;
        RECT 14.304 9.576 14.336 9.744 ;
  LAYER M1 ;
        RECT 14.304 9.54 14.336 9.612 ;
  LAYER M2 ;
        RECT 14.284 9.56 14.356 9.592 ;
  LAYER M2 ;
        RECT 14.32 9.56 14.48 9.592 ;
  LAYER M1 ;
        RECT 14.464 9.54 14.496 9.612 ;
  LAYER M2 ;
        RECT 14.444 9.56 14.516 9.592 ;
  LAYER M1 ;
        RECT 14.304 12.648 14.336 12.72 ;
  LAYER M2 ;
        RECT 14.284 12.668 14.356 12.7 ;
  LAYER M1 ;
        RECT 14.304 12.516 14.336 12.684 ;
  LAYER M1 ;
        RECT 14.304 12.48 14.336 12.552 ;
  LAYER M2 ;
        RECT 14.284 12.5 14.356 12.532 ;
  LAYER M2 ;
        RECT 14.32 12.5 14.48 12.532 ;
  LAYER M1 ;
        RECT 14.464 12.48 14.496 12.552 ;
  LAYER M2 ;
        RECT 14.444 12.5 14.516 12.532 ;
  LAYER M1 ;
        RECT 14.464 0.048 14.496 0.12 ;
  LAYER M2 ;
        RECT 14.444 0.068 14.516 0.1 ;
  LAYER M1 ;
        RECT 14.464 0.084 14.496 0.588 ;
  LAYER M1 ;
        RECT 14.464 0.588 14.496 12.516 ;
  LAYER M2 ;
        RECT 0.08 0.068 14.48 0.1 ;
  LAYER M1 ;
        RECT 5.664 0.888 5.696 0.96 ;
  LAYER M2 ;
        RECT 5.644 0.908 5.716 0.94 ;
  LAYER M2 ;
        RECT 2.8 0.908 5.68 0.94 ;
  LAYER M1 ;
        RECT 2.784 0.888 2.816 0.96 ;
  LAYER M2 ;
        RECT 2.764 0.908 2.836 0.94 ;
  LAYER M1 ;
        RECT 5.664 12.648 5.696 12.72 ;
  LAYER M2 ;
        RECT 5.644 12.668 5.716 12.7 ;
  LAYER M2 ;
        RECT 2.8 12.668 5.68 12.7 ;
  LAYER M1 ;
        RECT 2.784 12.648 2.816 12.72 ;
  LAYER M2 ;
        RECT 2.764 12.668 2.836 12.7 ;
  LAYER M1 ;
        RECT 8.544 12.648 8.576 12.72 ;
  LAYER M2 ;
        RECT 8.524 12.668 8.596 12.7 ;
  LAYER M2 ;
        RECT 5.68 12.668 8.56 12.7 ;
  LAYER M1 ;
        RECT 5.664 12.648 5.696 12.72 ;
  LAYER M2 ;
        RECT 5.644 12.668 5.716 12.7 ;
  LAYER M1 ;
        RECT 11.424 12.648 11.456 12.72 ;
  LAYER M2 ;
        RECT 11.404 12.668 11.476 12.7 ;
  LAYER M2 ;
        RECT 8.56 12.668 11.44 12.7 ;
  LAYER M1 ;
        RECT 8.544 12.648 8.576 12.72 ;
  LAYER M2 ;
        RECT 8.524 12.668 8.596 12.7 ;
  LAYER M1 ;
        RECT 11.424 0.888 11.456 0.96 ;
  LAYER M2 ;
        RECT 11.404 0.908 11.476 0.94 ;
  LAYER M2 ;
        RECT 11.44 0.908 14.32 0.94 ;
  LAYER M1 ;
        RECT 14.304 0.888 14.336 0.96 ;
  LAYER M2 ;
        RECT 14.284 0.908 14.356 0.94 ;
  LAYER M1 ;
        RECT 8.544 0.888 8.576 0.96 ;
  LAYER M2 ;
        RECT 8.524 0.908 8.596 0.94 ;
  LAYER M2 ;
        RECT 8.56 0.908 11.44 0.94 ;
  LAYER M1 ;
        RECT 11.424 0.888 11.456 0.96 ;
  LAYER M2 ;
        RECT 11.404 0.908 11.476 0.94 ;
  LAYER M1 ;
        RECT 6.144 9.204 6.176 9.276 ;
  LAYER M2 ;
        RECT 6.124 9.224 6.196 9.256 ;
  LAYER M2 ;
        RECT 6 9.224 6.16 9.256 ;
  LAYER M1 ;
        RECT 5.984 9.204 6.016 9.276 ;
  LAYER M2 ;
        RECT 5.964 9.224 6.036 9.256 ;
  LAYER M1 ;
        RECT 3.264 12.144 3.296 12.216 ;
  LAYER M2 ;
        RECT 3.244 12.164 3.316 12.196 ;
  LAYER M1 ;
        RECT 3.264 12.18 3.296 12.348 ;
  LAYER M1 ;
        RECT 3.264 12.312 3.296 12.384 ;
  LAYER M2 ;
        RECT 3.244 12.332 3.316 12.364 ;
  LAYER M2 ;
        RECT 3.28 12.332 6 12.364 ;
  LAYER M1 ;
        RECT 5.984 12.312 6.016 12.384 ;
  LAYER M2 ;
        RECT 5.964 12.332 6.036 12.364 ;
  LAYER M1 ;
        RECT 5.984 15.588 6.016 15.66 ;
  LAYER M2 ;
        RECT 5.964 15.608 6.036 15.64 ;
  LAYER M1 ;
        RECT 5.984 15.456 6.016 15.624 ;
  LAYER M1 ;
        RECT 5.984 9.24 6.016 15.456 ;
  LAYER M1 ;
        RECT 9.024 6.264 9.056 6.336 ;
  LAYER M2 ;
        RECT 9.004 6.284 9.076 6.316 ;
  LAYER M2 ;
        RECT 8.88 6.284 9.04 6.316 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M1 ;
        RECT 8.864 15.588 8.896 15.66 ;
  LAYER M2 ;
        RECT 8.844 15.608 8.916 15.64 ;
  LAYER M1 ;
        RECT 8.864 15.456 8.896 15.624 ;
  LAYER M1 ;
        RECT 8.864 6.3 8.896 15.456 ;
  LAYER M2 ;
        RECT 6 15.608 8.88 15.64 ;
  LAYER M1 ;
        RECT 3.264 9.204 3.296 9.276 ;
  LAYER M2 ;
        RECT 3.244 9.224 3.316 9.256 ;
  LAYER M2 ;
        RECT 3.12 9.224 3.28 9.256 ;
  LAYER M1 ;
        RECT 3.104 9.204 3.136 9.276 ;
  LAYER M2 ;
        RECT 3.084 9.224 3.156 9.256 ;
  LAYER M1 ;
        RECT 3.264 6.264 3.296 6.336 ;
  LAYER M2 ;
        RECT 3.244 6.284 3.316 6.316 ;
  LAYER M2 ;
        RECT 3.12 6.284 3.28 6.316 ;
  LAYER M1 ;
        RECT 3.104 6.264 3.136 6.336 ;
  LAYER M2 ;
        RECT 3.084 6.284 3.156 6.316 ;
  LAYER M1 ;
        RECT 3.104 15.756 3.136 15.828 ;
  LAYER M2 ;
        RECT 3.084 15.776 3.156 15.808 ;
  LAYER M1 ;
        RECT 3.104 15.456 3.136 15.792 ;
  LAYER M1 ;
        RECT 3.104 6.3 3.136 15.456 ;
  LAYER M1 ;
        RECT 9.024 9.204 9.056 9.276 ;
  LAYER M2 ;
        RECT 9.004 9.224 9.076 9.256 ;
  LAYER M1 ;
        RECT 9.024 9.24 9.056 9.408 ;
  LAYER M1 ;
        RECT 9.024 9.372 9.056 9.444 ;
  LAYER M2 ;
        RECT 9.004 9.392 9.076 9.424 ;
  LAYER M2 ;
        RECT 9.04 9.392 11.76 9.424 ;
  LAYER M1 ;
        RECT 11.744 9.372 11.776 9.444 ;
  LAYER M2 ;
        RECT 11.724 9.392 11.796 9.424 ;
  LAYER M1 ;
        RECT 9.024 12.144 9.056 12.216 ;
  LAYER M2 ;
        RECT 9.004 12.164 9.076 12.196 ;
  LAYER M1 ;
        RECT 9.024 12.18 9.056 12.348 ;
  LAYER M1 ;
        RECT 9.024 12.312 9.056 12.384 ;
  LAYER M2 ;
        RECT 9.004 12.332 9.076 12.364 ;
  LAYER M2 ;
        RECT 9.04 12.332 11.76 12.364 ;
  LAYER M1 ;
        RECT 11.744 12.312 11.776 12.384 ;
  LAYER M2 ;
        RECT 11.724 12.332 11.796 12.364 ;
  LAYER M1 ;
        RECT 11.744 15.756 11.776 15.828 ;
  LAYER M2 ;
        RECT 11.724 15.776 11.796 15.808 ;
  LAYER M1 ;
        RECT 11.744 15.456 11.776 15.792 ;
  LAYER M1 ;
        RECT 11.744 9.408 11.776 15.456 ;
  LAYER M2 ;
        RECT 3.12 15.776 11.76 15.808 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M2 ;
        RECT 3.28 6.284 6.16 6.316 ;
  LAYER M1 ;
        RECT 3.264 6.264 3.296 6.336 ;
  LAYER M2 ;
        RECT 3.244 6.284 3.316 6.316 ;
  LAYER M1 ;
        RECT 6.144 12.144 6.176 12.216 ;
  LAYER M2 ;
        RECT 6.124 12.164 6.196 12.196 ;
  LAYER M2 ;
        RECT 6.16 12.164 9.04 12.196 ;
  LAYER M1 ;
        RECT 9.024 12.144 9.056 12.216 ;
  LAYER M2 ;
        RECT 9.004 12.164 9.076 12.196 ;
  LAYER M1 ;
        RECT 0.384 3.324 0.416 3.396 ;
  LAYER M2 ;
        RECT 0.364 3.344 0.436 3.376 ;
  LAYER M2 ;
        RECT 0.24 3.344 0.4 3.376 ;
  LAYER M1 ;
        RECT 0.224 3.324 0.256 3.396 ;
  LAYER M2 ;
        RECT 0.204 3.344 0.276 3.376 ;
  LAYER M1 ;
        RECT 0.384 6.264 0.416 6.336 ;
  LAYER M2 ;
        RECT 0.364 6.284 0.436 6.316 ;
  LAYER M2 ;
        RECT 0.24 6.284 0.4 6.316 ;
  LAYER M1 ;
        RECT 0.224 6.264 0.256 6.336 ;
  LAYER M2 ;
        RECT 0.204 6.284 0.276 6.316 ;
  LAYER M1 ;
        RECT 0.384 9.204 0.416 9.276 ;
  LAYER M2 ;
        RECT 0.364 9.224 0.436 9.256 ;
  LAYER M2 ;
        RECT 0.24 9.224 0.4 9.256 ;
  LAYER M1 ;
        RECT 0.224 9.204 0.256 9.276 ;
  LAYER M2 ;
        RECT 0.204 9.224 0.276 9.256 ;
  LAYER M1 ;
        RECT 0.384 12.144 0.416 12.216 ;
  LAYER M2 ;
        RECT 0.364 12.164 0.436 12.196 ;
  LAYER M2 ;
        RECT 0.24 12.164 0.4 12.196 ;
  LAYER M1 ;
        RECT 0.224 12.144 0.256 12.216 ;
  LAYER M2 ;
        RECT 0.204 12.164 0.276 12.196 ;
  LAYER M1 ;
        RECT 0.384 15.084 0.416 15.156 ;
  LAYER M2 ;
        RECT 0.364 15.104 0.436 15.136 ;
  LAYER M2 ;
        RECT 0.24 15.104 0.4 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.084 0.256 15.156 ;
  LAYER M2 ;
        RECT 0.204 15.104 0.276 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.924 0.256 15.996 ;
  LAYER M2 ;
        RECT 0.204 15.944 0.276 15.976 ;
  LAYER M1 ;
        RECT 0.224 15.456 0.256 15.96 ;
  LAYER M1 ;
        RECT 0.224 3.36 0.256 15.456 ;
  LAYER M1 ;
        RECT 11.904 3.324 11.936 3.396 ;
  LAYER M2 ;
        RECT 11.884 3.344 11.956 3.376 ;
  LAYER M1 ;
        RECT 11.904 3.36 11.936 3.528 ;
  LAYER M1 ;
        RECT 11.904 3.492 11.936 3.564 ;
  LAYER M2 ;
        RECT 11.884 3.512 11.956 3.544 ;
  LAYER M2 ;
        RECT 11.92 3.512 14.64 3.544 ;
  LAYER M1 ;
        RECT 14.624 3.492 14.656 3.564 ;
  LAYER M2 ;
        RECT 14.604 3.512 14.676 3.544 ;
  LAYER M1 ;
        RECT 11.904 6.264 11.936 6.336 ;
  LAYER M2 ;
        RECT 11.884 6.284 11.956 6.316 ;
  LAYER M1 ;
        RECT 11.904 6.3 11.936 6.468 ;
  LAYER M1 ;
        RECT 11.904 6.432 11.936 6.504 ;
  LAYER M2 ;
        RECT 11.884 6.452 11.956 6.484 ;
  LAYER M2 ;
        RECT 11.92 6.452 14.64 6.484 ;
  LAYER M1 ;
        RECT 14.624 6.432 14.656 6.504 ;
  LAYER M2 ;
        RECT 14.604 6.452 14.676 6.484 ;
  LAYER M1 ;
        RECT 11.904 9.204 11.936 9.276 ;
  LAYER M2 ;
        RECT 11.884 9.224 11.956 9.256 ;
  LAYER M1 ;
        RECT 11.904 9.24 11.936 9.408 ;
  LAYER M1 ;
        RECT 11.904 9.372 11.936 9.444 ;
  LAYER M2 ;
        RECT 11.884 9.392 11.956 9.424 ;
  LAYER M2 ;
        RECT 11.92 9.392 14.64 9.424 ;
  LAYER M1 ;
        RECT 14.624 9.372 14.656 9.444 ;
  LAYER M2 ;
        RECT 14.604 9.392 14.676 9.424 ;
  LAYER M1 ;
        RECT 11.904 12.144 11.936 12.216 ;
  LAYER M2 ;
        RECT 11.884 12.164 11.956 12.196 ;
  LAYER M1 ;
        RECT 11.904 12.18 11.936 12.348 ;
  LAYER M1 ;
        RECT 11.904 12.312 11.936 12.384 ;
  LAYER M2 ;
        RECT 11.884 12.332 11.956 12.364 ;
  LAYER M2 ;
        RECT 11.92 12.332 14.64 12.364 ;
  LAYER M1 ;
        RECT 14.624 12.312 14.656 12.384 ;
  LAYER M2 ;
        RECT 14.604 12.332 14.676 12.364 ;
  LAYER M1 ;
        RECT 11.904 15.084 11.936 15.156 ;
  LAYER M2 ;
        RECT 11.884 15.104 11.956 15.136 ;
  LAYER M1 ;
        RECT 11.904 15.12 11.936 15.288 ;
  LAYER M1 ;
        RECT 11.904 15.252 11.936 15.324 ;
  LAYER M2 ;
        RECT 11.884 15.272 11.956 15.304 ;
  LAYER M2 ;
        RECT 11.92 15.272 14.64 15.304 ;
  LAYER M1 ;
        RECT 14.624 15.252 14.656 15.324 ;
  LAYER M2 ;
        RECT 14.604 15.272 14.676 15.304 ;
  LAYER M1 ;
        RECT 14.624 15.924 14.656 15.996 ;
  LAYER M2 ;
        RECT 14.604 15.944 14.676 15.976 ;
  LAYER M1 ;
        RECT 14.624 15.456 14.656 15.96 ;
  LAYER M1 ;
        RECT 14.624 3.528 14.656 15.456 ;
  LAYER M2 ;
        RECT 0.24 15.944 14.64 15.976 ;
  LAYER M1 ;
        RECT 3.264 3.324 3.296 3.396 ;
  LAYER M2 ;
        RECT 3.244 3.344 3.316 3.376 ;
  LAYER M2 ;
        RECT 0.4 3.344 3.28 3.376 ;
  LAYER M1 ;
        RECT 0.384 3.324 0.416 3.396 ;
  LAYER M2 ;
        RECT 0.364 3.344 0.436 3.376 ;
  LAYER M1 ;
        RECT 3.264 15.084 3.296 15.156 ;
  LAYER M2 ;
        RECT 3.244 15.104 3.316 15.136 ;
  LAYER M2 ;
        RECT 0.4 15.104 3.28 15.136 ;
  LAYER M1 ;
        RECT 0.384 15.084 0.416 15.156 ;
  LAYER M2 ;
        RECT 0.364 15.104 0.436 15.136 ;
  LAYER M1 ;
        RECT 6.144 15.084 6.176 15.156 ;
  LAYER M2 ;
        RECT 6.124 15.104 6.196 15.136 ;
  LAYER M2 ;
        RECT 3.28 15.104 6.16 15.136 ;
  LAYER M1 ;
        RECT 3.264 15.084 3.296 15.156 ;
  LAYER M2 ;
        RECT 3.244 15.104 3.316 15.136 ;
  LAYER M1 ;
        RECT 9.024 15.084 9.056 15.156 ;
  LAYER M2 ;
        RECT 9.004 15.104 9.076 15.136 ;
  LAYER M2 ;
        RECT 6.16 15.104 9.04 15.136 ;
  LAYER M1 ;
        RECT 6.144 15.084 6.176 15.156 ;
  LAYER M2 ;
        RECT 6.124 15.104 6.196 15.136 ;
  LAYER M1 ;
        RECT 9.024 3.324 9.056 3.396 ;
  LAYER M2 ;
        RECT 9.004 3.344 9.076 3.376 ;
  LAYER M2 ;
        RECT 9.04 3.344 11.92 3.376 ;
  LAYER M1 ;
        RECT 11.904 3.324 11.936 3.396 ;
  LAYER M2 ;
        RECT 11.884 3.344 11.956 3.376 ;
  LAYER M1 ;
        RECT 6.144 3.324 6.176 3.396 ;
  LAYER M2 ;
        RECT 6.124 3.344 6.196 3.376 ;
  LAYER M2 ;
        RECT 6.16 3.344 9.04 3.376 ;
  LAYER M1 ;
        RECT 9.024 3.324 9.056 3.396 ;
  LAYER M2 ;
        RECT 9.004 3.344 9.076 3.376 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M1 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M3 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M1 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M2 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M3 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M1 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M2 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M3 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M1 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M2 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M3 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M1 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M2 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M3 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M1 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M2 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M3 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M1 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M2 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M3 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M1 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M2 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M3 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M1 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M2 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M3 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M1 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M2 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M3 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M1 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M2 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M3 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M1 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M2 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M3 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M1 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M2 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M3 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M1 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M2 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M3 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M1 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M2 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M3 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M1 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M2 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M3 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M1 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M2 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M3 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M1 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M2 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M3 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M1 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M2 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M3 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M1 ;
        RECT 11.92 0.924 14.32 3.36 ;
  LAYER M2 ;
        RECT 11.92 0.924 14.32 3.36 ;
  LAYER M3 ;
        RECT 11.92 0.924 14.32 3.36 ;
  LAYER M1 ;
        RECT 11.92 3.864 14.32 6.3 ;
  LAYER M2 ;
        RECT 11.92 3.864 14.32 6.3 ;
  LAYER M3 ;
        RECT 11.92 3.864 14.32 6.3 ;
  LAYER M1 ;
        RECT 11.92 6.804 14.32 9.24 ;
  LAYER M2 ;
        RECT 11.92 6.804 14.32 9.24 ;
  LAYER M3 ;
        RECT 11.92 6.804 14.32 9.24 ;
  LAYER M1 ;
        RECT 11.92 9.744 14.32 12.18 ;
  LAYER M2 ;
        RECT 11.92 9.744 14.32 12.18 ;
  LAYER M3 ;
        RECT 11.92 9.744 14.32 12.18 ;
  LAYER M1 ;
        RECT 11.92 12.684 14.32 15.12 ;
  LAYER M2 ;
        RECT 11.92 12.684 14.32 15.12 ;
  LAYER M3 ;
        RECT 11.92 12.684 14.32 15.12 ;
  END 
END Cap_30fF_Cap_60fF
