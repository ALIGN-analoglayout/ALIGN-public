MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 2.5600 BY 3.4440 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
      LAYER M2 ;
        RECT 0.2040 0.9500 2.1960 0.9820 ;
      LAYER M2 ;
        RECT 0.2040 1.7900 2.1960 1.8220 ;
      LAYER M2 ;
        RECT 0.2040 2.6300 2.1960 2.6620 ;
    END
  END S
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1940 2.3560 0.2260 ;
      LAYER M2 ;
        RECT 0.2840 1.0340 2.2760 1.0660 ;
      LAYER M2 ;
        RECT 0.2840 1.8740 2.3560 1.9060 ;
      LAYER M2 ;
        RECT 0.2840 2.7140 2.2760 2.7460 ;
    END
  END D0
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
      LAYER M2 ;
        RECT 0.3640 1.1180 2.3560 1.1500 ;
      LAYER M2 ;
        RECT 1.0040 1.9580 1.7160 1.9900 ;
      LAYER M2 ;
        RECT 0.3640 2.7980 2.3560 2.8300 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3620 1.7160 0.3940 ;
      LAYER M2 ;
        RECT 0.3640 1.2020 2.3560 1.2340 ;
      LAYER M2 ;
        RECT 1.0040 2.0420 1.7160 2.0740 ;
      LAYER M2 ;
        RECT 0.3640 2.8820 2.3560 2.9140 ;
    END
  END D2
  PIN D3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.4460 2.3560 0.4780 ;
      LAYER M2 ;
        RECT 1.0040 1.2860 1.7160 1.3180 ;
      LAYER M2 ;
        RECT 0.3640 2.1260 2.3560 2.1580 ;
      LAYER M2 ;
        RECT 1.0040 2.9660 1.7160 2.9980 ;
    END
  END D3
  PIN D4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.5300 2.3560 0.5620 ;
      LAYER M2 ;
        RECT 1.0040 1.3700 1.7160 1.4020 ;
      LAYER M2 ;
        RECT 0.3640 2.2100 2.3560 2.2420 ;
      LAYER M2 ;
        RECT 1.0040 3.0500 1.7160 3.0820 ;
    END
  END D4
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 0.1620 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER M3 ;
      RECT 1.1000 0.1740 1.1400 0.2460 ;
    LAYER V2 ;
      RECT 1.1000 0.1940 1.1400 0.2260 ;
    LAYER V2 ;
      RECT 1.1000 0.1940 1.1400 0.2260 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.3040 0.1940 0.3360 0.2260 ;
    LAYER V1 ;
      RECT 2.2240 0.1940 2.2560 0.2260 ;
    LAYER V1 ;
      RECT 0.9440 0.1940 0.9760 0.2260 ;
    LAYER V1 ;
      RECT 1.5840 0.1940 1.6160 0.2260 ;
    LAYER M3 ;
      RECT 1.2600 0.2580 1.3000 0.3300 ;
    LAYER V2 ;
      RECT 1.2600 0.2780 1.3000 0.3100 ;
    LAYER V2 ;
      RECT 1.2600 0.2780 1.3000 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER M3 ;
      RECT 1.3400 0.3420 1.3800 0.4140 ;
    LAYER V2 ;
      RECT 1.3400 0.3620 1.3800 0.3940 ;
    LAYER V2 ;
      RECT 1.3400 0.3620 1.3800 0.3940 ;
    LAYER V1 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V1 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER M3 ;
      RECT 1.3400 0.4260 1.3800 0.4980 ;
    LAYER V2 ;
      RECT 1.3400 0.4460 1.3800 0.4780 ;
    LAYER V2 ;
      RECT 1.3400 0.4460 1.3800 0.4780 ;
    LAYER V1 ;
      RECT 0.3840 0.4460 0.4160 0.4780 ;
    LAYER V1 ;
      RECT 2.3040 0.4460 2.3360 0.4780 ;
    LAYER M3 ;
      RECT 1.4200 0.5100 1.4600 0.5820 ;
    LAYER V2 ;
      RECT 1.4200 0.5300 1.4600 0.5620 ;
    LAYER V2 ;
      RECT 1.4200 0.5300 1.4600 0.5620 ;
    LAYER V1 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V1 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 0.3040 0.9300 0.3360 1.5900 ;
    LAYER M1 ;
      RECT 2.2240 0.9300 2.2560 1.5900 ;
    LAYER M1 ;
      RECT 0.9440 0.9300 0.9760 1.5900 ;
    LAYER M1 ;
      RECT 1.5840 0.9300 1.6160 1.5900 ;
    LAYER M1 ;
      RECT 0.2240 0.9300 0.2560 1.5900 ;
    LAYER V0 ;
      RECT 0.2240 1.1180 0.2560 1.1500 ;
    LAYER V0 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V0 ;
      RECT 0.2240 1.3700 0.2560 1.4020 ;
    LAYER M1 ;
      RECT 2.1440 0.9300 2.1760 1.5900 ;
    LAYER V0 ;
      RECT 2.1440 1.1180 2.1760 1.1500 ;
    LAYER V0 ;
      RECT 2.1440 1.2440 2.1760 1.2760 ;
    LAYER V0 ;
      RECT 2.1440 1.3700 2.1760 1.4020 ;
    LAYER M1 ;
      RECT 0.8640 0.9300 0.8960 1.5900 ;
    LAYER V0 ;
      RECT 0.8640 1.1180 0.8960 1.1500 ;
    LAYER V0 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V0 ;
      RECT 0.8640 1.3700 0.8960 1.4020 ;
    LAYER M1 ;
      RECT 1.5040 0.9300 1.5360 1.5900 ;
    LAYER V0 ;
      RECT 1.5040 1.1180 1.5360 1.1500 ;
    LAYER V0 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V0 ;
      RECT 1.5040 1.3700 1.5360 1.4020 ;
    LAYER M1 ;
      RECT 0.3840 0.9300 0.4160 1.5900 ;
    LAYER V0 ;
      RECT 0.3840 1.1180 0.4160 1.1500 ;
    LAYER V0 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V0 ;
      RECT 0.3840 1.3700 0.4160 1.4020 ;
    LAYER M1 ;
      RECT 2.3040 0.9300 2.3360 1.5900 ;
    LAYER V0 ;
      RECT 2.3040 1.1180 2.3360 1.1500 ;
    LAYER V0 ;
      RECT 2.3040 1.2440 2.3360 1.2760 ;
    LAYER V0 ;
      RECT 2.3040 1.3700 2.3360 1.4020 ;
    LAYER M1 ;
      RECT 1.0240 0.9300 1.0560 1.5900 ;
    LAYER V0 ;
      RECT 1.0240 1.1180 1.0560 1.1500 ;
    LAYER V0 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V0 ;
      RECT 1.0240 1.3700 1.0560 1.4020 ;
    LAYER M1 ;
      RECT 1.6640 0.9300 1.6960 1.5900 ;
    LAYER V0 ;
      RECT 1.6640 1.1180 1.6960 1.1500 ;
    LAYER V0 ;
      RECT 1.6640 1.2440 1.6960 1.2760 ;
    LAYER V0 ;
      RECT 1.6640 1.3700 1.6960 1.4020 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 1.0020 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 0.9500 1.2200 0.9820 ;
    LAYER V1 ;
      RECT 0.2240 0.9500 0.2560 0.9820 ;
    LAYER V1 ;
      RECT 2.1440 0.9500 2.1760 0.9820 ;
    LAYER V1 ;
      RECT 0.8640 0.9500 0.8960 0.9820 ;
    LAYER V1 ;
      RECT 1.5040 0.9500 1.5360 0.9820 ;
    LAYER M3 ;
      RECT 1.1000 0.1740 1.1400 1.0860 ;
    LAYER V2 ;
      RECT 1.1000 0.1940 1.1400 0.2260 ;
    LAYER V2 ;
      RECT 1.1000 1.0340 1.1400 1.0660 ;
    LAYER V1 ;
      RECT 1.0240 1.0340 1.0560 1.0660 ;
    LAYER V1 ;
      RECT 1.6640 1.0340 1.6960 1.0660 ;
    LAYER V1 ;
      RECT 0.3040 1.0340 0.3360 1.0660 ;
    LAYER V1 ;
      RECT 2.2240 1.0340 2.2560 1.0660 ;
    LAYER V1 ;
      RECT 0.9440 1.0340 0.9760 1.0660 ;
    LAYER V1 ;
      RECT 1.5840 1.0340 1.6160 1.0660 ;
    LAYER M3 ;
      RECT 1.2600 0.2580 1.3000 1.1700 ;
    LAYER V2 ;
      RECT 1.2600 0.2780 1.3000 0.3100 ;
    LAYER V2 ;
      RECT 1.2600 1.1180 1.3000 1.1500 ;
    LAYER V1 ;
      RECT 0.3840 1.1180 0.4160 1.1500 ;
    LAYER V1 ;
      RECT 2.3040 1.1180 2.3360 1.1500 ;
    LAYER M3 ;
      RECT 1.3400 0.3420 1.3800 1.2540 ;
    LAYER V2 ;
      RECT 1.3400 0.3620 1.3800 0.3940 ;
    LAYER V2 ;
      RECT 1.3400 1.2020 1.3800 1.2340 ;
    LAYER V1 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V1 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER M3 ;
      RECT 1.3400 0.4260 1.3800 1.3380 ;
    LAYER V2 ;
      RECT 1.3400 0.4460 1.3800 0.4780 ;
    LAYER V2 ;
      RECT 1.3400 1.2860 1.3800 1.3180 ;
    LAYER V1 ;
      RECT 1.0240 1.2860 1.0560 1.3180 ;
    LAYER V1 ;
      RECT 1.6640 1.2860 1.6960 1.3180 ;
    LAYER M3 ;
      RECT 1.4200 0.5100 1.4600 1.4220 ;
    LAYER V2 ;
      RECT 1.4200 0.5300 1.4600 0.5620 ;
    LAYER V2 ;
      RECT 1.4200 1.3700 1.4600 1.4020 ;
    LAYER V1 ;
      RECT 1.0240 1.3700 1.0560 1.4020 ;
    LAYER V1 ;
      RECT 1.6640 1.3700 1.6960 1.4020 ;
    LAYER M1 ;
      RECT 0.3040 1.7700 0.3360 2.4300 ;
    LAYER M1 ;
      RECT 2.2240 1.7700 2.2560 2.4300 ;
    LAYER M1 ;
      RECT 0.9440 1.7700 0.9760 2.4300 ;
    LAYER M1 ;
      RECT 1.5840 1.7700 1.6160 2.4300 ;
    LAYER M1 ;
      RECT 0.2240 1.7700 0.2560 2.4300 ;
    LAYER V0 ;
      RECT 0.2240 1.9580 0.2560 1.9900 ;
    LAYER V0 ;
      RECT 0.2240 2.0840 0.2560 2.1160 ;
    LAYER V0 ;
      RECT 0.2240 2.2100 0.2560 2.2420 ;
    LAYER M1 ;
      RECT 2.1440 1.7700 2.1760 2.4300 ;
    LAYER V0 ;
      RECT 2.1440 1.9580 2.1760 1.9900 ;
    LAYER V0 ;
      RECT 2.1440 2.0840 2.1760 2.1160 ;
    LAYER V0 ;
      RECT 2.1440 2.2100 2.1760 2.2420 ;
    LAYER M1 ;
      RECT 0.8640 1.7700 0.8960 2.4300 ;
    LAYER V0 ;
      RECT 0.8640 1.9580 0.8960 1.9900 ;
    LAYER V0 ;
      RECT 0.8640 2.0840 0.8960 2.1160 ;
    LAYER V0 ;
      RECT 0.8640 2.2100 0.8960 2.2420 ;
    LAYER M1 ;
      RECT 1.5040 1.7700 1.5360 2.4300 ;
    LAYER V0 ;
      RECT 1.5040 1.9580 1.5360 1.9900 ;
    LAYER V0 ;
      RECT 1.5040 2.0840 1.5360 2.1160 ;
    LAYER V0 ;
      RECT 1.5040 2.2100 1.5360 2.2420 ;
    LAYER M1 ;
      RECT 0.3840 1.7700 0.4160 2.4300 ;
    LAYER V0 ;
      RECT 0.3840 1.9580 0.4160 1.9900 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.2100 0.4160 2.2420 ;
    LAYER M1 ;
      RECT 2.3040 1.7700 2.3360 2.4300 ;
    LAYER V0 ;
      RECT 2.3040 1.9580 2.3360 1.9900 ;
    LAYER V0 ;
      RECT 2.3040 2.0840 2.3360 2.1160 ;
    LAYER V0 ;
      RECT 2.3040 2.2100 2.3360 2.2420 ;
    LAYER M1 ;
      RECT 1.0240 1.7700 1.0560 2.4300 ;
    LAYER V0 ;
      RECT 1.0240 1.9580 1.0560 1.9900 ;
    LAYER V0 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V0 ;
      RECT 1.0240 2.2100 1.0560 2.2420 ;
    LAYER M1 ;
      RECT 1.6640 1.7700 1.6960 2.4300 ;
    LAYER V0 ;
      RECT 1.6640 1.9580 1.6960 1.9900 ;
    LAYER V0 ;
      RECT 1.6640 2.0840 1.6960 2.1160 ;
    LAYER V0 ;
      RECT 1.6640 2.2100 1.6960 2.2420 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 1.8420 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 1.7900 1.2200 1.8220 ;
    LAYER V1 ;
      RECT 0.2240 1.7900 0.2560 1.8220 ;
    LAYER V1 ;
      RECT 2.1440 1.7900 2.1760 1.8220 ;
    LAYER V1 ;
      RECT 0.8640 1.7900 0.8960 1.8220 ;
    LAYER V1 ;
      RECT 1.5040 1.7900 1.5360 1.8220 ;
    LAYER M3 ;
      RECT 1.1000 0.1740 1.1400 1.9260 ;
    LAYER V2 ;
      RECT 1.1000 0.1940 1.1400 0.2260 ;
    LAYER V2 ;
      RECT 1.1000 1.8740 1.1400 1.9060 ;
    LAYER V1 ;
      RECT 0.3840 1.8740 0.4160 1.9060 ;
    LAYER V1 ;
      RECT 2.3040 1.8740 2.3360 1.9060 ;
    LAYER V1 ;
      RECT 0.3040 1.8740 0.3360 1.9060 ;
    LAYER V1 ;
      RECT 2.2240 1.8740 2.2560 1.9060 ;
    LAYER V1 ;
      RECT 0.9440 1.8740 0.9760 1.9060 ;
    LAYER V1 ;
      RECT 1.5840 1.8740 1.6160 1.9060 ;
    LAYER M3 ;
      RECT 1.2600 0.2580 1.3000 2.0100 ;
    LAYER V2 ;
      RECT 1.2600 0.2780 1.3000 0.3100 ;
    LAYER V2 ;
      RECT 1.2600 1.9580 1.3000 1.9900 ;
    LAYER V1 ;
      RECT 1.0240 1.9580 1.0560 1.9900 ;
    LAYER V1 ;
      RECT 1.6640 1.9580 1.6960 1.9900 ;
    LAYER M3 ;
      RECT 1.3400 0.3420 1.3800 2.0940 ;
    LAYER V2 ;
      RECT 1.3400 0.3620 1.3800 0.3940 ;
    LAYER V2 ;
      RECT 1.3400 2.0420 1.3800 2.0740 ;
    LAYER V1 ;
      RECT 1.0240 2.0420 1.0560 2.0740 ;
    LAYER V1 ;
      RECT 1.6640 2.0420 1.6960 2.0740 ;
    LAYER M3 ;
      RECT 1.3400 0.4260 1.3800 2.1780 ;
    LAYER V2 ;
      RECT 1.3400 0.4460 1.3800 0.4780 ;
    LAYER V2 ;
      RECT 1.3400 2.1260 1.3800 2.1580 ;
    LAYER V1 ;
      RECT 0.3840 2.1260 0.4160 2.1580 ;
    LAYER V1 ;
      RECT 2.3040 2.1260 2.3360 2.1580 ;
    LAYER M3 ;
      RECT 1.4200 0.5100 1.4600 2.2620 ;
    LAYER V2 ;
      RECT 1.4200 0.5300 1.4600 0.5620 ;
    LAYER V2 ;
      RECT 1.4200 2.2100 1.4600 2.2420 ;
    LAYER V1 ;
      RECT 0.3840 2.2100 0.4160 2.2420 ;
    LAYER V1 ;
      RECT 2.3040 2.2100 2.3360 2.2420 ;
    LAYER M1 ;
      RECT 0.3040 2.6100 0.3360 3.2700 ;
    LAYER M1 ;
      RECT 2.2240 2.6100 2.2560 3.2700 ;
    LAYER M1 ;
      RECT 0.9440 2.6100 0.9760 3.2700 ;
    LAYER M1 ;
      RECT 1.5840 2.6100 1.6160 3.2700 ;
    LAYER M1 ;
      RECT 0.2240 2.6100 0.2560 3.2700 ;
    LAYER V0 ;
      RECT 0.2240 2.7980 0.2560 2.8300 ;
    LAYER V0 ;
      RECT 0.2240 2.9240 0.2560 2.9560 ;
    LAYER V0 ;
      RECT 0.2240 3.0500 0.2560 3.0820 ;
    LAYER M1 ;
      RECT 2.1440 2.6100 2.1760 3.2700 ;
    LAYER V0 ;
      RECT 2.1440 2.7980 2.1760 2.8300 ;
    LAYER V0 ;
      RECT 2.1440 2.9240 2.1760 2.9560 ;
    LAYER V0 ;
      RECT 2.1440 3.0500 2.1760 3.0820 ;
    LAYER M1 ;
      RECT 0.8640 2.6100 0.8960 3.2700 ;
    LAYER V0 ;
      RECT 0.8640 2.7980 0.8960 2.8300 ;
    LAYER V0 ;
      RECT 0.8640 2.9240 0.8960 2.9560 ;
    LAYER V0 ;
      RECT 0.8640 3.0500 0.8960 3.0820 ;
    LAYER M1 ;
      RECT 1.5040 2.6100 1.5360 3.2700 ;
    LAYER V0 ;
      RECT 1.5040 2.7980 1.5360 2.8300 ;
    LAYER V0 ;
      RECT 1.5040 2.9240 1.5360 2.9560 ;
    LAYER V0 ;
      RECT 1.5040 3.0500 1.5360 3.0820 ;
    LAYER M1 ;
      RECT 0.3840 2.6100 0.4160 3.2700 ;
    LAYER V0 ;
      RECT 0.3840 2.7980 0.4160 2.8300 ;
    LAYER V0 ;
      RECT 0.3840 2.9240 0.4160 2.9560 ;
    LAYER V0 ;
      RECT 0.3840 3.0500 0.4160 3.0820 ;
    LAYER M1 ;
      RECT 2.3040 2.6100 2.3360 3.2700 ;
    LAYER V0 ;
      RECT 2.3040 2.7980 2.3360 2.8300 ;
    LAYER V0 ;
      RECT 2.3040 2.9240 2.3360 2.9560 ;
    LAYER V0 ;
      RECT 2.3040 3.0500 2.3360 3.0820 ;
    LAYER M1 ;
      RECT 1.0240 2.6100 1.0560 3.2700 ;
    LAYER V0 ;
      RECT 1.0240 2.7980 1.0560 2.8300 ;
    LAYER V0 ;
      RECT 1.0240 2.9240 1.0560 2.9560 ;
    LAYER V0 ;
      RECT 1.0240 3.0500 1.0560 3.0820 ;
    LAYER M1 ;
      RECT 1.6640 2.6100 1.6960 3.2700 ;
    LAYER V0 ;
      RECT 1.6640 2.7980 1.6960 2.8300 ;
    LAYER V0 ;
      RECT 1.6640 2.9240 1.6960 2.9560 ;
    LAYER V0 ;
      RECT 1.6640 3.0500 1.6960 3.0820 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 2.6820 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 2.6300 1.2200 2.6620 ;
    LAYER V1 ;
      RECT 0.2240 2.6300 0.2560 2.6620 ;
    LAYER V1 ;
      RECT 2.1440 2.6300 2.1760 2.6620 ;
    LAYER V1 ;
      RECT 0.8640 2.6300 0.8960 2.6620 ;
    LAYER V1 ;
      RECT 1.5040 2.6300 1.5360 2.6620 ;
    LAYER M3 ;
      RECT 1.1000 0.1740 1.1400 2.7660 ;
    LAYER V2 ;
      RECT 1.1000 0.1940 1.1400 0.2260 ;
    LAYER V2 ;
      RECT 1.1000 2.7140 1.1400 2.7460 ;
    LAYER V1 ;
      RECT 1.0240 2.7140 1.0560 2.7460 ;
    LAYER V1 ;
      RECT 1.6640 2.7140 1.6960 2.7460 ;
    LAYER V1 ;
      RECT 0.3040 2.7140 0.3360 2.7460 ;
    LAYER V1 ;
      RECT 2.2240 2.7140 2.2560 2.7460 ;
    LAYER V1 ;
      RECT 0.9440 2.7140 0.9760 2.7460 ;
    LAYER V1 ;
      RECT 1.5840 2.7140 1.6160 2.7460 ;
    LAYER M3 ;
      RECT 1.2600 0.2580 1.3000 2.8500 ;
    LAYER V2 ;
      RECT 1.2600 0.2780 1.3000 0.3100 ;
    LAYER V2 ;
      RECT 1.2600 2.7980 1.3000 2.8300 ;
    LAYER V1 ;
      RECT 0.3840 2.7980 0.4160 2.8300 ;
    LAYER V1 ;
      RECT 2.3040 2.7980 2.3360 2.8300 ;
    LAYER M3 ;
      RECT 1.3400 0.3420 1.3800 2.9340 ;
    LAYER V2 ;
      RECT 1.3400 0.3620 1.3800 0.3940 ;
    LAYER V2 ;
      RECT 1.3400 2.8820 1.3800 2.9140 ;
    LAYER V1 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V1 ;
      RECT 2.3040 2.8820 2.3360 2.9140 ;
    LAYER M3 ;
      RECT 1.3400 0.4260 1.3800 3.0180 ;
    LAYER V2 ;
      RECT 1.3400 0.4460 1.3800 0.4780 ;
    LAYER V2 ;
      RECT 1.3400 2.9660 1.3800 2.9980 ;
    LAYER V1 ;
      RECT 1.0240 2.9660 1.0560 2.9980 ;
    LAYER V1 ;
      RECT 1.6640 2.9660 1.6960 2.9980 ;
    LAYER M3 ;
      RECT 1.4200 0.5100 1.4600 3.1020 ;
    LAYER V2 ;
      RECT 1.4200 0.5300 1.4600 0.5620 ;
    LAYER V2 ;
      RECT 1.4200 3.0500 1.4600 3.0820 ;
    LAYER V1 ;
      RECT 1.0240 3.0500 1.0560 3.0820 ;
    LAYER V1 ;
      RECT 1.6640 3.0500 1.6960 3.0820 ;
  END
END test
