MACRO switched_capacitor_combination
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_combination 0 0 ;
  SIZE 16 BY 31.416 ;
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.684 0.32 10.756 0.352 ;
      LAYER M2 ;
        RECT 9.964 0.488 10.036 0.52 ;
      LAYER M2 ;
        RECT 8.604 0.488 8.676 0.52 ;
      LAYER M2 ;
        RECT 10.24 0.32 10.72 0.352 ;
      LAYER M3 ;
        RECT 10.22 0.316 10.26 0.356 ;
      LAYER M4 ;
        RECT 10.08 0.316 10.24 0.356 ;
      LAYER M5 ;
        RECT 10.048 0.336 10.112 0.504 ;
      LAYER M4 ;
        RECT 10.08 0.484 10.24 0.524 ;
      LAYER M3 ;
        RECT 10.22 0.484 10.26 0.524 ;
      LAYER M2 ;
        RECT 10 0.488 10.24 0.52 ;
      LAYER M2 ;
        RECT 8.64 0.488 10.08 0.52 ;
    END
  END phi2
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.764 0.152 10.836 0.184 ;
      LAYER M2 ;
        RECT 10.044 0.656 10.116 0.688 ;
      LAYER M2 ;
        RECT 8.684 0.656 8.756 0.688 ;
      LAYER M2 ;
        RECT 10.08 0.152 10.8 0.184 ;
      LAYER M3 ;
        RECT 10.06 0.168 10.1 0.672 ;
      LAYER M2 ;
        RECT 10.064 0.656 10.096 0.688 ;
      LAYER M2 ;
        RECT 8.88 0.656 10.08 0.688 ;
      LAYER M3 ;
        RECT 8.86 0.652 8.9 0.692 ;
      LAYER M4 ;
        RECT 8.72 0.652 8.88 0.692 ;
      LAYER M3 ;
        RECT 8.7 0.652 8.74 0.692 ;
      LAYER M2 ;
        RECT 8.704 0.656 8.736 0.688 ;
    END
  END agnd
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 0.32 0.436 0.352 ;
      LAYER M2 ;
        RECT 9.324 0.572 9.396 0.604 ;
      LAYER M2 ;
        RECT 7.964 0.572 8.036 0.604 ;
      LAYER M2 ;
        RECT 0.4 0.32 7.84 0.352 ;
      LAYER M3 ;
        RECT 7.82 0.336 7.86 0.588 ;
      LAYER M4 ;
        RECT 7.84 0.568 8 0.608 ;
      LAYER M3 ;
        RECT 7.98 0.568 8.02 0.608 ;
      LAYER M2 ;
        RECT 7.984 0.572 8.016 0.604 ;
      LAYER M4 ;
        RECT 8 0.568 8.16 0.608 ;
      LAYER M3 ;
        RECT 8.14 0.568 8.18 0.608 ;
      LAYER M2 ;
        RECT 8.16 0.572 9.36 0.604 ;
    END
  END phi1
  PIN Vin
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.284 0.152 0.356 0.184 ;
    END
  END Vin
  PIN Vin_ota
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.404 0.74 9.476 0.772 ;
      LAYER M1 ;
        RECT 3.76 31.128 3.792 31.2 ;
      LAYER M2 ;
        RECT 3.74 31.148 3.812 31.18 ;
      LAYER M1 ;
        RECT 12.688 31.128 12.72 31.2 ;
      LAYER M2 ;
        RECT 12.668 31.148 12.74 31.18 ;
      LAYER M2 ;
        RECT 3.776 31.148 12.704 31.18 ;
      LAYER M2 ;
        RECT 9.44 0.74 9.68 0.772 ;
      LAYER M3 ;
        RECT 9.66 0.756 9.7 30.996 ;
      LAYER M4 ;
        RECT 9.36 30.976 9.68 31.016 ;
      LAYER M5 ;
        RECT 9.328 30.996 9.392 31.164 ;
      LAYER M4 ;
        RECT 9.34 31.144 9.38 31.184 ;
      LAYER M3 ;
        RECT 9.34 31.144 9.38 31.184 ;
      LAYER M2 ;
        RECT 9.344 31.148 9.376 31.18 ;
    END
  END Vin_ota
  PIN Voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.044 0.74 8.116 0.772 ;
      LAYER M1 ;
        RECT 3.92 14.748 3.952 14.82 ;
      LAYER M2 ;
        RECT 3.9 14.768 3.972 14.8 ;
      LAYER M1 ;
        RECT 12.848 14.748 12.88 14.82 ;
      LAYER M2 ;
        RECT 12.828 14.768 12.9 14.8 ;
      LAYER M2 ;
        RECT 3.936 14.768 12.864 14.8 ;
      LAYER M2 ;
        RECT 8.064 0.74 8.096 0.772 ;
      LAYER M3 ;
        RECT 8.06 0.756 8.1 1.008 ;
      LAYER M4 ;
        RECT 7.92 0.988 8.08 1.028 ;
      LAYER M5 ;
        RECT 7.888 1.008 7.952 14.784 ;
      LAYER M4 ;
        RECT 7.9 14.764 7.94 14.804 ;
      LAYER M3 ;
        RECT 7.9 14.764 7.94 14.804 ;
      LAYER M2 ;
        RECT 7.904 14.768 7.936 14.8 ;
    END
  END Voutn
  OBS 
  LAYER M1 ;
        RECT 9.632 14.16 9.664 14.232 ;
  LAYER M2 ;
        RECT 9.612 14.18 9.684 14.212 ;
  LAYER M1 ;
        RECT 6.656 14.16 6.688 14.232 ;
  LAYER M2 ;
        RECT 6.636 14.18 6.708 14.212 ;
  LAYER M2 ;
        RECT 6.672 14.18 9.648 14.212 ;
  LAYER M2 ;
        RECT 9.244 0.824 9.956 0.856 ;
  LAYER M1 ;
        RECT 6.736 30.96 6.768 31.032 ;
  LAYER M2 ;
        RECT 6.716 30.98 6.788 31.012 ;
  LAYER M1 ;
        RECT 9.712 30.96 9.744 31.032 ;
  LAYER M2 ;
        RECT 9.692 30.98 9.764 31.012 ;
  LAYER M2 ;
        RECT 6.752 30.98 9.728 31.012 ;
  LAYER M2 ;
        RECT 9.504 14.18 9.536 14.212 ;
  LAYER M3 ;
        RECT 9.5 0.84 9.54 14.196 ;
  LAYER M2 ;
        RECT 9.504 0.824 9.536 0.856 ;
  LAYER M2 ;
        RECT 7.184 14.18 7.216 14.212 ;
  LAYER M3 ;
        RECT 7.18 14.196 7.22 14.7 ;
  LAYER M4 ;
        RECT 7.18 14.68 7.22 14.72 ;
  LAYER M5 ;
        RECT 7.168 14.7 7.232 30.996 ;
  LAYER M4 ;
        RECT 7.18 30.976 7.22 31.016 ;
  LAYER M3 ;
        RECT 7.18 30.976 7.22 31.016 ;
  LAYER M2 ;
        RECT 7.184 30.98 7.216 31.012 ;
  LAYER M1 ;
        RECT 9.792 1.224 9.824 1.296 ;
  LAYER M2 ;
        RECT 9.772 1.244 9.844 1.276 ;
  LAYER M1 ;
        RECT 6.816 1.224 6.848 1.296 ;
  LAYER M2 ;
        RECT 6.796 1.244 6.868 1.276 ;
  LAYER M2 ;
        RECT 6.832 1.244 9.808 1.276 ;
  LAYER M2 ;
        RECT 10.604 0.236 10.676 0.268 ;
  LAYER M2 ;
        RECT 0.444 0.236 0.516 0.268 ;
  LAYER M2 ;
        RECT 9.84 1.244 10.32 1.276 ;
  LAYER M3 ;
        RECT 10.3 0.252 10.34 1.26 ;
  LAYER M4 ;
        RECT 10.32 0.232 10.64 0.272 ;
  LAYER M3 ;
        RECT 10.62 0.232 10.66 0.272 ;
  LAYER M2 ;
        RECT 10.624 0.236 10.656 0.268 ;
  LAYER M2 ;
        RECT 0.8 1.244 6.8 1.276 ;
  LAYER M3 ;
        RECT 0.78 0.252 0.82 1.26 ;
  LAYER M4 ;
        RECT 0.48 0.232 0.8 0.272 ;
  LAYER M3 ;
        RECT 0.46 0.232 0.5 0.272 ;
  LAYER M2 ;
        RECT 0.464 0.236 0.496 0.268 ;
  LAYER M2 ;
        RECT 7.884 0.824 8.596 0.856 ;
  LAYER M1 ;
        RECT 6.896 14.916 6.928 14.988 ;
  LAYER M2 ;
        RECT 6.876 14.936 6.948 14.968 ;
  LAYER M1 ;
        RECT 9.872 14.916 9.904 14.988 ;
  LAYER M2 ;
        RECT 9.852 14.936 9.924 14.968 ;
  LAYER M2 ;
        RECT 6.912 14.936 9.888 14.968 ;
  LAYER M2 ;
        RECT 7.904 0.824 7.936 0.856 ;
  LAYER M3 ;
        RECT 7.9 0.84 7.94 1.596 ;
  LAYER M4 ;
        RECT 7.776 1.576 7.92 1.616 ;
  LAYER M5 ;
        RECT 7.744 1.596 7.808 14.952 ;
  LAYER M4 ;
        RECT 7.776 14.932 7.92 14.972 ;
  LAYER M3 ;
        RECT 7.9 14.932 7.94 14.972 ;
  LAYER M2 ;
        RECT 7.904 14.936 7.936 14.968 ;
  LAYER M1 ;
        RECT 7.04 4.92 7.072 4.992 ;
  LAYER M2 ;
        RECT 7.02 4.94 7.092 4.972 ;
  LAYER M2 ;
        RECT 7.056 4.94 9.808 4.972 ;
  LAYER M1 ;
        RECT 9.792 4.92 9.824 4.992 ;
  LAYER M2 ;
        RECT 9.772 4.94 9.844 4.972 ;
  LAYER M1 ;
        RECT 7.04 8.028 7.072 8.1 ;
  LAYER M2 ;
        RECT 7.02 8.048 7.092 8.08 ;
  LAYER M2 ;
        RECT 7.056 8.048 9.808 8.08 ;
  LAYER M1 ;
        RECT 9.792 8.028 9.824 8.1 ;
  LAYER M2 ;
        RECT 9.772 8.048 9.844 8.08 ;
  LAYER M1 ;
        RECT 10.016 4.92 10.048 4.992 ;
  LAYER M2 ;
        RECT 9.996 4.94 10.068 4.972 ;
  LAYER M1 ;
        RECT 10.016 4.788 10.048 4.956 ;
  LAYER M1 ;
        RECT 10.016 4.752 10.048 4.824 ;
  LAYER M2 ;
        RECT 9.996 4.772 10.068 4.804 ;
  LAYER M2 ;
        RECT 9.808 4.772 10.032 4.804 ;
  LAYER M1 ;
        RECT 9.792 4.752 9.824 4.824 ;
  LAYER M2 ;
        RECT 9.772 4.772 9.844 4.804 ;
  LAYER M1 ;
        RECT 10.016 8.028 10.048 8.1 ;
  LAYER M2 ;
        RECT 9.996 8.048 10.068 8.08 ;
  LAYER M1 ;
        RECT 10.016 7.896 10.048 8.064 ;
  LAYER M1 ;
        RECT 10.016 7.86 10.048 7.932 ;
  LAYER M2 ;
        RECT 9.996 7.88 10.068 7.912 ;
  LAYER M2 ;
        RECT 9.808 7.88 10.032 7.912 ;
  LAYER M1 ;
        RECT 9.792 7.86 9.824 7.932 ;
  LAYER M2 ;
        RECT 9.772 7.88 9.844 7.912 ;
  LAYER M1 ;
        RECT 9.792 1.224 9.824 1.296 ;
  LAYER M2 ;
        RECT 9.772 1.244 9.844 1.276 ;
  LAYER M1 ;
        RECT 9.792 1.26 9.824 1.512 ;
  LAYER M1 ;
        RECT 9.792 1.512 9.824 8.064 ;
  LAYER M1 ;
        RECT 4.064 8.028 4.096 8.1 ;
  LAYER M2 ;
        RECT 4.044 8.048 4.116 8.08 ;
  LAYER M2 ;
        RECT 4.08 8.048 6.832 8.08 ;
  LAYER M1 ;
        RECT 6.816 8.028 6.848 8.1 ;
  LAYER M2 ;
        RECT 6.796 8.048 6.868 8.08 ;
  LAYER M1 ;
        RECT 4.064 4.92 4.096 4.992 ;
  LAYER M2 ;
        RECT 4.044 4.94 4.116 4.972 ;
  LAYER M2 ;
        RECT 4.08 4.94 6.832 4.972 ;
  LAYER M1 ;
        RECT 6.816 4.92 6.848 4.992 ;
  LAYER M2 ;
        RECT 6.796 4.94 6.868 4.972 ;
  LAYER M1 ;
        RECT 6.816 1.224 6.848 1.296 ;
  LAYER M2 ;
        RECT 6.796 1.244 6.868 1.276 ;
  LAYER M1 ;
        RECT 6.816 1.26 6.848 1.512 ;
  LAYER M1 ;
        RECT 6.816 1.512 6.848 8.064 ;
  LAYER M2 ;
        RECT 6.832 1.244 9.808 1.276 ;
  LAYER M1 ;
        RECT 12.992 1.812 13.024 1.884 ;
  LAYER M2 ;
        RECT 12.972 1.832 13.044 1.864 ;
  LAYER M1 ;
        RECT 12.992 1.68 13.024 1.848 ;
  LAYER M1 ;
        RECT 12.992 1.644 13.024 1.716 ;
  LAYER M2 ;
        RECT 12.972 1.664 13.044 1.696 ;
  LAYER M2 ;
        RECT 12.784 1.664 13.008 1.696 ;
  LAYER M1 ;
        RECT 12.768 1.644 12.8 1.716 ;
  LAYER M2 ;
        RECT 12.748 1.664 12.82 1.696 ;
  LAYER M1 ;
        RECT 12.992 4.92 13.024 4.992 ;
  LAYER M2 ;
        RECT 12.972 4.94 13.044 4.972 ;
  LAYER M1 ;
        RECT 12.992 4.788 13.024 4.956 ;
  LAYER M1 ;
        RECT 12.992 4.752 13.024 4.824 ;
  LAYER M2 ;
        RECT 12.972 4.772 13.044 4.804 ;
  LAYER M2 ;
        RECT 12.784 4.772 13.008 4.804 ;
  LAYER M1 ;
        RECT 12.768 4.752 12.8 4.824 ;
  LAYER M2 ;
        RECT 12.748 4.772 12.82 4.804 ;
  LAYER M1 ;
        RECT 12.992 8.028 13.024 8.1 ;
  LAYER M2 ;
        RECT 12.972 8.048 13.044 8.08 ;
  LAYER M1 ;
        RECT 12.992 7.896 13.024 8.064 ;
  LAYER M1 ;
        RECT 12.992 7.86 13.024 7.932 ;
  LAYER M2 ;
        RECT 12.972 7.88 13.044 7.912 ;
  LAYER M2 ;
        RECT 12.784 7.88 13.008 7.912 ;
  LAYER M1 ;
        RECT 12.768 7.86 12.8 7.932 ;
  LAYER M2 ;
        RECT 12.748 7.88 12.82 7.912 ;
  LAYER M1 ;
        RECT 12.992 11.136 13.024 11.208 ;
  LAYER M2 ;
        RECT 12.972 11.156 13.044 11.188 ;
  LAYER M1 ;
        RECT 12.992 11.004 13.024 11.172 ;
  LAYER M1 ;
        RECT 12.992 10.968 13.024 11.04 ;
  LAYER M2 ;
        RECT 12.972 10.988 13.044 11.02 ;
  LAYER M2 ;
        RECT 12.784 10.988 13.008 11.02 ;
  LAYER M1 ;
        RECT 12.768 10.968 12.8 11.04 ;
  LAYER M2 ;
        RECT 12.748 10.988 12.82 11.02 ;
  LAYER M1 ;
        RECT 10.016 1.812 10.048 1.884 ;
  LAYER M2 ;
        RECT 9.996 1.832 10.068 1.864 ;
  LAYER M2 ;
        RECT 10.032 1.832 12.784 1.864 ;
  LAYER M1 ;
        RECT 12.768 1.812 12.8 1.884 ;
  LAYER M2 ;
        RECT 12.748 1.832 12.82 1.864 ;
  LAYER M1 ;
        RECT 10.016 11.136 10.048 11.208 ;
  LAYER M2 ;
        RECT 9.996 11.156 10.068 11.188 ;
  LAYER M2 ;
        RECT 10.032 11.156 12.784 11.188 ;
  LAYER M1 ;
        RECT 12.768 11.136 12.8 11.208 ;
  LAYER M2 ;
        RECT 12.748 11.156 12.82 11.188 ;
  LAYER M1 ;
        RECT 12.768 1.056 12.8 1.128 ;
  LAYER M2 ;
        RECT 12.748 1.076 12.82 1.108 ;
  LAYER M1 ;
        RECT 12.768 1.092 12.8 1.512 ;
  LAYER M1 ;
        RECT 12.768 1.512 12.8 11.172 ;
  LAYER M1 ;
        RECT 4.064 1.812 4.096 1.884 ;
  LAYER M2 ;
        RECT 4.044 1.832 4.116 1.864 ;
  LAYER M1 ;
        RECT 4.064 1.68 4.096 1.848 ;
  LAYER M1 ;
        RECT 4.064 1.644 4.096 1.716 ;
  LAYER M2 ;
        RECT 4.044 1.664 4.116 1.696 ;
  LAYER M2 ;
        RECT 3.856 1.664 4.08 1.696 ;
  LAYER M1 ;
        RECT 3.84 1.644 3.872 1.716 ;
  LAYER M2 ;
        RECT 3.82 1.664 3.892 1.696 ;
  LAYER M1 ;
        RECT 4.064 11.136 4.096 11.208 ;
  LAYER M2 ;
        RECT 4.044 11.156 4.116 11.188 ;
  LAYER M1 ;
        RECT 4.064 11.004 4.096 11.172 ;
  LAYER M1 ;
        RECT 4.064 10.968 4.096 11.04 ;
  LAYER M2 ;
        RECT 4.044 10.988 4.116 11.02 ;
  LAYER M2 ;
        RECT 3.856 10.988 4.08 11.02 ;
  LAYER M1 ;
        RECT 3.84 10.968 3.872 11.04 ;
  LAYER M2 ;
        RECT 3.82 10.988 3.892 11.02 ;
  LAYER M1 ;
        RECT 1.088 1.812 1.12 1.884 ;
  LAYER M2 ;
        RECT 1.068 1.832 1.14 1.864 ;
  LAYER M2 ;
        RECT 1.104 1.832 3.856 1.864 ;
  LAYER M1 ;
        RECT 3.84 1.812 3.872 1.884 ;
  LAYER M2 ;
        RECT 3.82 1.832 3.892 1.864 ;
  LAYER M1 ;
        RECT 1.088 4.92 1.12 4.992 ;
  LAYER M2 ;
        RECT 1.068 4.94 1.14 4.972 ;
  LAYER M2 ;
        RECT 1.104 4.94 3.856 4.972 ;
  LAYER M1 ;
        RECT 3.84 4.92 3.872 4.992 ;
  LAYER M2 ;
        RECT 3.82 4.94 3.892 4.972 ;
  LAYER M1 ;
        RECT 1.088 8.028 1.12 8.1 ;
  LAYER M2 ;
        RECT 1.068 8.048 1.14 8.08 ;
  LAYER M2 ;
        RECT 1.104 8.048 3.856 8.08 ;
  LAYER M1 ;
        RECT 3.84 8.028 3.872 8.1 ;
  LAYER M2 ;
        RECT 3.82 8.048 3.892 8.08 ;
  LAYER M1 ;
        RECT 1.088 11.136 1.12 11.208 ;
  LAYER M2 ;
        RECT 1.068 11.156 1.14 11.188 ;
  LAYER M2 ;
        RECT 1.104 11.156 3.856 11.188 ;
  LAYER M1 ;
        RECT 3.84 11.136 3.872 11.208 ;
  LAYER M2 ;
        RECT 3.82 11.156 3.892 11.188 ;
  LAYER M1 ;
        RECT 3.84 1.056 3.872 1.128 ;
  LAYER M2 ;
        RECT 3.82 1.076 3.892 1.108 ;
  LAYER M1 ;
        RECT 3.84 1.092 3.872 1.512 ;
  LAYER M1 ;
        RECT 3.84 1.512 3.872 11.172 ;
  LAYER M2 ;
        RECT 3.856 1.076 12.784 1.108 ;
  LAYER M1 ;
        RECT 7.04 11.136 7.072 11.208 ;
  LAYER M2 ;
        RECT 7.02 11.156 7.092 11.188 ;
  LAYER M2 ;
        RECT 7.056 11.156 10.032 11.188 ;
  LAYER M1 ;
        RECT 10.016 11.136 10.048 11.208 ;
  LAYER M2 ;
        RECT 9.996 11.156 10.068 11.188 ;
  LAYER M1 ;
        RECT 7.04 1.812 7.072 1.884 ;
  LAYER M2 ;
        RECT 7.02 1.832 7.092 1.864 ;
  LAYER M2 ;
        RECT 4.08 1.832 7.056 1.864 ;
  LAYER M1 ;
        RECT 4.064 1.812 4.096 1.884 ;
  LAYER M2 ;
        RECT 4.044 1.832 4.116 1.864 ;
  LAYER M1 ;
        RECT 9.408 7.356 9.44 7.428 ;
  LAYER M2 ;
        RECT 9.388 7.376 9.46 7.408 ;
  LAYER M2 ;
        RECT 9.424 7.376 9.648 7.408 ;
  LAYER M1 ;
        RECT 9.632 7.356 9.664 7.428 ;
  LAYER M2 ;
        RECT 9.612 7.376 9.684 7.408 ;
  LAYER M1 ;
        RECT 9.408 10.464 9.44 10.536 ;
  LAYER M2 ;
        RECT 9.388 10.484 9.46 10.516 ;
  LAYER M2 ;
        RECT 9.424 10.484 9.648 10.516 ;
  LAYER M1 ;
        RECT 9.632 10.464 9.664 10.536 ;
  LAYER M2 ;
        RECT 9.612 10.484 9.684 10.516 ;
  LAYER M1 ;
        RECT 12.384 7.356 12.416 7.428 ;
  LAYER M2 ;
        RECT 12.364 7.376 12.436 7.408 ;
  LAYER M1 ;
        RECT 12.384 7.392 12.416 7.56 ;
  LAYER M1 ;
        RECT 12.384 7.524 12.416 7.596 ;
  LAYER M2 ;
        RECT 12.364 7.544 12.436 7.576 ;
  LAYER M2 ;
        RECT 9.648 7.544 12.4 7.576 ;
  LAYER M1 ;
        RECT 9.632 7.524 9.664 7.596 ;
  LAYER M2 ;
        RECT 9.612 7.544 9.684 7.576 ;
  LAYER M1 ;
        RECT 12.384 10.464 12.416 10.536 ;
  LAYER M2 ;
        RECT 12.364 10.484 12.436 10.516 ;
  LAYER M1 ;
        RECT 12.384 10.5 12.416 10.668 ;
  LAYER M1 ;
        RECT 12.384 10.632 12.416 10.704 ;
  LAYER M2 ;
        RECT 12.364 10.652 12.436 10.684 ;
  LAYER M2 ;
        RECT 9.648 10.652 12.4 10.684 ;
  LAYER M1 ;
        RECT 9.632 10.632 9.664 10.704 ;
  LAYER M2 ;
        RECT 9.612 10.652 9.684 10.684 ;
  LAYER M1 ;
        RECT 9.632 14.16 9.664 14.232 ;
  LAYER M2 ;
        RECT 9.612 14.18 9.684 14.212 ;
  LAYER M1 ;
        RECT 9.632 13.944 9.664 14.196 ;
  LAYER M1 ;
        RECT 9.632 7.392 9.664 13.944 ;
  LAYER M1 ;
        RECT 6.432 10.464 6.464 10.536 ;
  LAYER M2 ;
        RECT 6.412 10.484 6.484 10.516 ;
  LAYER M2 ;
        RECT 6.448 10.484 6.672 10.516 ;
  LAYER M1 ;
        RECT 6.656 10.464 6.688 10.536 ;
  LAYER M2 ;
        RECT 6.636 10.484 6.708 10.516 ;
  LAYER M1 ;
        RECT 6.432 7.356 6.464 7.428 ;
  LAYER M2 ;
        RECT 6.412 7.376 6.484 7.408 ;
  LAYER M2 ;
        RECT 6.448 7.376 6.672 7.408 ;
  LAYER M1 ;
        RECT 6.656 7.356 6.688 7.428 ;
  LAYER M2 ;
        RECT 6.636 7.376 6.708 7.408 ;
  LAYER M1 ;
        RECT 6.656 14.16 6.688 14.232 ;
  LAYER M2 ;
        RECT 6.636 14.18 6.708 14.212 ;
  LAYER M1 ;
        RECT 6.656 13.944 6.688 14.196 ;
  LAYER M1 ;
        RECT 6.656 7.392 6.688 13.944 ;
  LAYER M2 ;
        RECT 6.672 14.18 9.648 14.212 ;
  LAYER M1 ;
        RECT 15.36 4.248 15.392 4.32 ;
  LAYER M2 ;
        RECT 15.34 4.268 15.412 4.3 ;
  LAYER M2 ;
        RECT 15.376 4.268 15.76 4.3 ;
  LAYER M1 ;
        RECT 15.744 4.248 15.776 4.32 ;
  LAYER M2 ;
        RECT 15.724 4.268 15.796 4.3 ;
  LAYER M1 ;
        RECT 15.36 7.356 15.392 7.428 ;
  LAYER M2 ;
        RECT 15.34 7.376 15.412 7.408 ;
  LAYER M2 ;
        RECT 15.376 7.376 15.76 7.408 ;
  LAYER M1 ;
        RECT 15.744 7.356 15.776 7.428 ;
  LAYER M2 ;
        RECT 15.724 7.376 15.796 7.408 ;
  LAYER M1 ;
        RECT 15.36 10.464 15.392 10.536 ;
  LAYER M2 ;
        RECT 15.34 10.484 15.412 10.516 ;
  LAYER M2 ;
        RECT 15.376 10.484 15.76 10.516 ;
  LAYER M1 ;
        RECT 15.744 10.464 15.776 10.536 ;
  LAYER M2 ;
        RECT 15.724 10.484 15.796 10.516 ;
  LAYER M1 ;
        RECT 15.36 13.572 15.392 13.644 ;
  LAYER M2 ;
        RECT 15.34 13.592 15.412 13.624 ;
  LAYER M2 ;
        RECT 15.376 13.592 15.76 13.624 ;
  LAYER M1 ;
        RECT 15.744 13.572 15.776 13.644 ;
  LAYER M2 ;
        RECT 15.724 13.592 15.796 13.624 ;
  LAYER M1 ;
        RECT 15.744 14.328 15.776 14.4 ;
  LAYER M2 ;
        RECT 15.724 14.348 15.796 14.38 ;
  LAYER M1 ;
        RECT 15.744 13.944 15.776 14.364 ;
  LAYER M1 ;
        RECT 15.744 4.284 15.776 13.944 ;
  LAYER M1 ;
        RECT 3.456 4.248 3.488 4.32 ;
  LAYER M2 ;
        RECT 3.436 4.268 3.508 4.3 ;
  LAYER M1 ;
        RECT 3.456 4.284 3.488 4.452 ;
  LAYER M1 ;
        RECT 3.456 4.416 3.488 4.488 ;
  LAYER M2 ;
        RECT 3.436 4.436 3.508 4.468 ;
  LAYER M2 ;
        RECT 0.88 4.436 3.472 4.468 ;
  LAYER M1 ;
        RECT 0.864 4.416 0.896 4.488 ;
  LAYER M2 ;
        RECT 0.844 4.436 0.916 4.468 ;
  LAYER M1 ;
        RECT 3.456 7.356 3.488 7.428 ;
  LAYER M2 ;
        RECT 3.436 7.376 3.508 7.408 ;
  LAYER M1 ;
        RECT 3.456 7.392 3.488 7.56 ;
  LAYER M1 ;
        RECT 3.456 7.524 3.488 7.596 ;
  LAYER M2 ;
        RECT 3.436 7.544 3.508 7.576 ;
  LAYER M2 ;
        RECT 0.88 7.544 3.472 7.576 ;
  LAYER M1 ;
        RECT 0.864 7.524 0.896 7.596 ;
  LAYER M2 ;
        RECT 0.844 7.544 0.916 7.576 ;
  LAYER M1 ;
        RECT 3.456 10.464 3.488 10.536 ;
  LAYER M2 ;
        RECT 3.436 10.484 3.508 10.516 ;
  LAYER M1 ;
        RECT 3.456 10.5 3.488 10.668 ;
  LAYER M1 ;
        RECT 3.456 10.632 3.488 10.704 ;
  LAYER M2 ;
        RECT 3.436 10.652 3.508 10.684 ;
  LAYER M2 ;
        RECT 0.88 10.652 3.472 10.684 ;
  LAYER M1 ;
        RECT 0.864 10.632 0.896 10.704 ;
  LAYER M2 ;
        RECT 0.844 10.652 0.916 10.684 ;
  LAYER M1 ;
        RECT 3.456 13.572 3.488 13.644 ;
  LAYER M2 ;
        RECT 3.436 13.592 3.508 13.624 ;
  LAYER M1 ;
        RECT 3.456 13.608 3.488 13.776 ;
  LAYER M1 ;
        RECT 3.456 13.74 3.488 13.812 ;
  LAYER M2 ;
        RECT 3.436 13.76 3.508 13.792 ;
  LAYER M2 ;
        RECT 0.88 13.76 3.472 13.792 ;
  LAYER M1 ;
        RECT 0.864 13.74 0.896 13.812 ;
  LAYER M2 ;
        RECT 0.844 13.76 0.916 13.792 ;
  LAYER M1 ;
        RECT 0.864 14.328 0.896 14.4 ;
  LAYER M2 ;
        RECT 0.844 14.348 0.916 14.38 ;
  LAYER M1 ;
        RECT 0.864 13.944 0.896 14.364 ;
  LAYER M1 ;
        RECT 0.864 4.452 0.896 13.944 ;
  LAYER M2 ;
        RECT 0.88 14.348 15.76 14.38 ;
  LAYER M1 ;
        RECT 12.384 4.248 12.416 4.32 ;
  LAYER M2 ;
        RECT 12.364 4.268 12.436 4.3 ;
  LAYER M2 ;
        RECT 12.4 4.268 15.376 4.3 ;
  LAYER M1 ;
        RECT 15.36 4.248 15.392 4.32 ;
  LAYER M2 ;
        RECT 15.34 4.268 15.412 4.3 ;
  LAYER M1 ;
        RECT 12.384 13.572 12.416 13.644 ;
  LAYER M2 ;
        RECT 12.364 13.592 12.436 13.624 ;
  LAYER M2 ;
        RECT 12.4 13.592 15.376 13.624 ;
  LAYER M1 ;
        RECT 15.36 13.572 15.392 13.644 ;
  LAYER M2 ;
        RECT 15.34 13.592 15.412 13.624 ;
  LAYER M1 ;
        RECT 9.408 13.572 9.44 13.644 ;
  LAYER M2 ;
        RECT 9.388 13.592 9.46 13.624 ;
  LAYER M2 ;
        RECT 9.424 13.592 12.4 13.624 ;
  LAYER M1 ;
        RECT 12.384 13.572 12.416 13.644 ;
  LAYER M2 ;
        RECT 12.364 13.592 12.436 13.624 ;
  LAYER M1 ;
        RECT 6.432 13.572 6.464 13.644 ;
  LAYER M2 ;
        RECT 6.412 13.592 6.484 13.624 ;
  LAYER M2 ;
        RECT 6.448 13.592 9.424 13.624 ;
  LAYER M1 ;
        RECT 9.408 13.572 9.44 13.644 ;
  LAYER M2 ;
        RECT 9.388 13.592 9.46 13.624 ;
  LAYER M1 ;
        RECT 6.432 4.248 6.464 4.32 ;
  LAYER M2 ;
        RECT 6.412 4.268 6.484 4.3 ;
  LAYER M2 ;
        RECT 3.472 4.268 6.448 4.3 ;
  LAYER M1 ;
        RECT 3.456 4.248 3.488 4.32 ;
  LAYER M2 ;
        RECT 3.436 4.268 3.508 4.3 ;
  LAYER M1 ;
        RECT 9.408 4.248 9.44 4.32 ;
  LAYER M2 ;
        RECT 9.388 4.268 9.46 4.3 ;
  LAYER M2 ;
        RECT 6.448 4.268 9.424 4.3 ;
  LAYER M1 ;
        RECT 6.432 4.248 6.464 4.32 ;
  LAYER M2 ;
        RECT 6.412 4.268 6.484 4.3 ;
  LAYER M1 ;
        RECT 12.944 1.764 15.44 4.368 ;
  LAYER M3 ;
        RECT 12.944 1.764 15.44 4.368 ;
  LAYER M2 ;
        RECT 12.944 1.764 15.44 4.368 ;
  LAYER M1 ;
        RECT 12.944 4.872 15.44 7.476 ;
  LAYER M3 ;
        RECT 12.944 4.872 15.44 7.476 ;
  LAYER M2 ;
        RECT 12.944 4.872 15.44 7.476 ;
  LAYER M1 ;
        RECT 12.944 7.98 15.44 10.584 ;
  LAYER M3 ;
        RECT 12.944 7.98 15.44 10.584 ;
  LAYER M2 ;
        RECT 12.944 7.98 15.44 10.584 ;
  LAYER M1 ;
        RECT 12.944 11.088 15.44 13.692 ;
  LAYER M3 ;
        RECT 12.944 11.088 15.44 13.692 ;
  LAYER M2 ;
        RECT 12.944 11.088 15.44 13.692 ;
  LAYER M1 ;
        RECT 9.968 1.764 12.464 4.368 ;
  LAYER M3 ;
        RECT 9.968 1.764 12.464 4.368 ;
  LAYER M2 ;
        RECT 9.968 1.764 12.464 4.368 ;
  LAYER M1 ;
        RECT 9.968 4.872 12.464 7.476 ;
  LAYER M3 ;
        RECT 9.968 4.872 12.464 7.476 ;
  LAYER M2 ;
        RECT 9.968 4.872 12.464 7.476 ;
  LAYER M1 ;
        RECT 9.968 7.98 12.464 10.584 ;
  LAYER M3 ;
        RECT 9.968 7.98 12.464 10.584 ;
  LAYER M2 ;
        RECT 9.968 7.98 12.464 10.584 ;
  LAYER M1 ;
        RECT 9.968 11.088 12.464 13.692 ;
  LAYER M3 ;
        RECT 9.968 11.088 12.464 13.692 ;
  LAYER M2 ;
        RECT 9.968 11.088 12.464 13.692 ;
  LAYER M1 ;
        RECT 6.992 1.764 9.488 4.368 ;
  LAYER M3 ;
        RECT 6.992 1.764 9.488 4.368 ;
  LAYER M2 ;
        RECT 6.992 1.764 9.488 4.368 ;
  LAYER M1 ;
        RECT 6.992 4.872 9.488 7.476 ;
  LAYER M3 ;
        RECT 6.992 4.872 9.488 7.476 ;
  LAYER M2 ;
        RECT 6.992 4.872 9.488 7.476 ;
  LAYER M1 ;
        RECT 6.992 7.98 9.488 10.584 ;
  LAYER M3 ;
        RECT 6.992 7.98 9.488 10.584 ;
  LAYER M2 ;
        RECT 6.992 7.98 9.488 10.584 ;
  LAYER M1 ;
        RECT 6.992 11.088 9.488 13.692 ;
  LAYER M3 ;
        RECT 6.992 11.088 9.488 13.692 ;
  LAYER M2 ;
        RECT 6.992 11.088 9.488 13.692 ;
  LAYER M1 ;
        RECT 4.016 1.764 6.512 4.368 ;
  LAYER M3 ;
        RECT 4.016 1.764 6.512 4.368 ;
  LAYER M2 ;
        RECT 4.016 1.764 6.512 4.368 ;
  LAYER M1 ;
        RECT 4.016 4.872 6.512 7.476 ;
  LAYER M3 ;
        RECT 4.016 4.872 6.512 7.476 ;
  LAYER M2 ;
        RECT 4.016 4.872 6.512 7.476 ;
  LAYER M1 ;
        RECT 4.016 7.98 6.512 10.584 ;
  LAYER M3 ;
        RECT 4.016 7.98 6.512 10.584 ;
  LAYER M2 ;
        RECT 4.016 7.98 6.512 10.584 ;
  LAYER M1 ;
        RECT 4.016 11.088 6.512 13.692 ;
  LAYER M3 ;
        RECT 4.016 11.088 6.512 13.692 ;
  LAYER M2 ;
        RECT 4.016 11.088 6.512 13.692 ;
  LAYER M1 ;
        RECT 1.04 1.764 3.536 4.368 ;
  LAYER M3 ;
        RECT 1.04 1.764 3.536 4.368 ;
  LAYER M2 ;
        RECT 1.04 1.764 3.536 4.368 ;
  LAYER M1 ;
        RECT 1.04 4.872 3.536 7.476 ;
  LAYER M3 ;
        RECT 1.04 4.872 3.536 7.476 ;
  LAYER M2 ;
        RECT 1.04 4.872 3.536 7.476 ;
  LAYER M1 ;
        RECT 1.04 7.98 3.536 10.584 ;
  LAYER M3 ;
        RECT 1.04 7.98 3.536 10.584 ;
  LAYER M2 ;
        RECT 1.04 7.98 3.536 10.584 ;
  LAYER M1 ;
        RECT 1.04 11.088 3.536 13.692 ;
  LAYER M3 ;
        RECT 1.04 11.088 3.536 13.692 ;
  LAYER M2 ;
        RECT 1.04 11.088 3.536 13.692 ;
  LAYER M1 ;
        RECT 10.704 0.132 10.736 0.792 ;
  LAYER M1 ;
        RECT 10.784 0.132 10.816 0.792 ;
  LAYER M1 ;
        RECT 10.624 0.572 10.656 0.604 ;
  LAYER M1 ;
        RECT 0.384 0.132 0.416 0.792 ;
  LAYER M1 ;
        RECT 0.304 0.132 0.336 0.792 ;
  LAYER M1 ;
        RECT 0.464 0.572 0.496 0.604 ;
  LAYER M1 ;
        RECT 9.344 0.216 9.376 0.876 ;
  LAYER M1 ;
        RECT 9.984 0.216 10.016 0.876 ;
  LAYER M1 ;
        RECT 9.264 0.216 9.296 0.876 ;
  LAYER M1 ;
        RECT 9.904 0.216 9.936 0.876 ;
  LAYER M1 ;
        RECT 9.424 0.216 9.456 0.876 ;
  LAYER M1 ;
        RECT 10.064 0.404 10.096 0.436 ;
  LAYER M1 ;
        RECT 7.984 0.216 8.016 0.876 ;
  LAYER M1 ;
        RECT 8.624 0.216 8.656 0.876 ;
  LAYER M1 ;
        RECT 7.904 0.216 7.936 0.876 ;
  LAYER M1 ;
        RECT 8.544 0.216 8.576 0.876 ;
  LAYER M1 ;
        RECT 8.064 0.216 8.096 0.876 ;
  LAYER M1 ;
        RECT 8.704 0.404 8.736 0.436 ;
  LAYER M1 ;
        RECT 9.488 24.156 9.52 24.228 ;
  LAYER M2 ;
        RECT 9.468 24.176 9.54 24.208 ;
  LAYER M2 ;
        RECT 6.752 24.176 9.504 24.208 ;
  LAYER M1 ;
        RECT 6.736 24.156 6.768 24.228 ;
  LAYER M2 ;
        RECT 6.716 24.176 6.788 24.208 ;
  LAYER M1 ;
        RECT 6.512 21.048 6.544 21.12 ;
  LAYER M2 ;
        RECT 6.492 21.068 6.564 21.1 ;
  LAYER M1 ;
        RECT 6.512 21.084 6.544 21.252 ;
  LAYER M1 ;
        RECT 6.512 21.216 6.544 21.288 ;
  LAYER M2 ;
        RECT 6.492 21.236 6.564 21.268 ;
  LAYER M2 ;
        RECT 6.528 21.236 6.752 21.268 ;
  LAYER M1 ;
        RECT 6.736 21.216 6.768 21.288 ;
  LAYER M2 ;
        RECT 6.716 21.236 6.788 21.268 ;
  LAYER M1 ;
        RECT 6.736 30.96 6.768 31.032 ;
  LAYER M2 ;
        RECT 6.716 30.98 6.788 31.012 ;
  LAYER M1 ;
        RECT 6.736 30.744 6.768 30.996 ;
  LAYER M1 ;
        RECT 6.736 21.252 6.768 30.744 ;
  LAYER M1 ;
        RECT 12.464 27.264 12.496 27.336 ;
  LAYER M2 ;
        RECT 12.444 27.284 12.516 27.316 ;
  LAYER M2 ;
        RECT 9.728 27.284 12.48 27.316 ;
  LAYER M1 ;
        RECT 9.712 27.264 9.744 27.336 ;
  LAYER M2 ;
        RECT 9.692 27.284 9.764 27.316 ;
  LAYER M1 ;
        RECT 9.712 30.96 9.744 31.032 ;
  LAYER M2 ;
        RECT 9.692 30.98 9.764 31.012 ;
  LAYER M1 ;
        RECT 9.712 30.744 9.744 30.996 ;
  LAYER M1 ;
        RECT 9.712 27.3 9.744 30.744 ;
  LAYER M2 ;
        RECT 6.752 30.98 9.728 31.012 ;
  LAYER M1 ;
        RECT 6.512 24.156 6.544 24.228 ;
  LAYER M2 ;
        RECT 6.492 24.176 6.564 24.208 ;
  LAYER M2 ;
        RECT 3.776 24.176 6.528 24.208 ;
  LAYER M1 ;
        RECT 3.76 24.156 3.792 24.228 ;
  LAYER M2 ;
        RECT 3.74 24.176 3.812 24.208 ;
  LAYER M1 ;
        RECT 6.512 27.264 6.544 27.336 ;
  LAYER M2 ;
        RECT 6.492 27.284 6.564 27.316 ;
  LAYER M2 ;
        RECT 3.776 27.284 6.528 27.316 ;
  LAYER M1 ;
        RECT 3.76 27.264 3.792 27.336 ;
  LAYER M2 ;
        RECT 3.74 27.284 3.812 27.316 ;
  LAYER M1 ;
        RECT 3.76 31.128 3.792 31.2 ;
  LAYER M2 ;
        RECT 3.74 31.148 3.812 31.18 ;
  LAYER M1 ;
        RECT 3.76 30.744 3.792 31.164 ;
  LAYER M1 ;
        RECT 3.76 24.192 3.792 30.744 ;
  LAYER M1 ;
        RECT 12.464 24.156 12.496 24.228 ;
  LAYER M2 ;
        RECT 12.444 24.176 12.516 24.208 ;
  LAYER M1 ;
        RECT 12.464 24.192 12.496 24.36 ;
  LAYER M1 ;
        RECT 12.464 24.324 12.496 24.396 ;
  LAYER M2 ;
        RECT 12.444 24.344 12.516 24.376 ;
  LAYER M2 ;
        RECT 12.48 24.344 12.704 24.376 ;
  LAYER M1 ;
        RECT 12.688 24.324 12.72 24.396 ;
  LAYER M2 ;
        RECT 12.668 24.344 12.74 24.376 ;
  LAYER M1 ;
        RECT 12.464 21.048 12.496 21.12 ;
  LAYER M2 ;
        RECT 12.444 21.068 12.516 21.1 ;
  LAYER M1 ;
        RECT 12.464 21.084 12.496 21.252 ;
  LAYER M1 ;
        RECT 12.464 21.216 12.496 21.288 ;
  LAYER M2 ;
        RECT 12.444 21.236 12.516 21.268 ;
  LAYER M2 ;
        RECT 12.48 21.236 12.704 21.268 ;
  LAYER M1 ;
        RECT 12.688 21.216 12.72 21.288 ;
  LAYER M2 ;
        RECT 12.668 21.236 12.74 21.268 ;
  LAYER M1 ;
        RECT 12.688 31.128 12.72 31.2 ;
  LAYER M2 ;
        RECT 12.668 31.148 12.74 31.18 ;
  LAYER M1 ;
        RECT 12.688 30.744 12.72 31.164 ;
  LAYER M1 ;
        RECT 12.688 21.252 12.72 30.744 ;
  LAYER M2 ;
        RECT 3.776 31.148 12.704 31.18 ;
  LAYER M1 ;
        RECT 9.488 27.264 9.52 27.336 ;
  LAYER M2 ;
        RECT 9.468 27.284 9.54 27.316 ;
  LAYER M2 ;
        RECT 6.528 27.284 9.504 27.316 ;
  LAYER M1 ;
        RECT 6.512 27.264 6.544 27.336 ;
  LAYER M2 ;
        RECT 6.492 27.284 6.564 27.316 ;
  LAYER M1 ;
        RECT 9.488 21.048 9.52 21.12 ;
  LAYER M2 ;
        RECT 9.468 21.068 9.54 21.1 ;
  LAYER M2 ;
        RECT 9.504 21.068 12.48 21.1 ;
  LAYER M1 ;
        RECT 12.464 21.048 12.496 21.12 ;
  LAYER M2 ;
        RECT 12.444 21.068 12.516 21.1 ;
  LAYER M1 ;
        RECT 3.536 30.372 3.568 30.444 ;
  LAYER M2 ;
        RECT 3.516 30.392 3.588 30.424 ;
  LAYER M2 ;
        RECT 0.8 30.392 3.552 30.424 ;
  LAYER M1 ;
        RECT 0.784 30.372 0.816 30.444 ;
  LAYER M2 ;
        RECT 0.764 30.392 0.836 30.424 ;
  LAYER M1 ;
        RECT 3.536 27.264 3.568 27.336 ;
  LAYER M2 ;
        RECT 3.516 27.284 3.588 27.316 ;
  LAYER M2 ;
        RECT 0.8 27.284 3.552 27.316 ;
  LAYER M1 ;
        RECT 0.784 27.264 0.816 27.336 ;
  LAYER M2 ;
        RECT 0.764 27.284 0.836 27.316 ;
  LAYER M1 ;
        RECT 3.536 24.156 3.568 24.228 ;
  LAYER M2 ;
        RECT 3.516 24.176 3.588 24.208 ;
  LAYER M2 ;
        RECT 0.8 24.176 3.552 24.208 ;
  LAYER M1 ;
        RECT 0.784 24.156 0.816 24.228 ;
  LAYER M2 ;
        RECT 0.764 24.176 0.836 24.208 ;
  LAYER M1 ;
        RECT 3.536 21.048 3.568 21.12 ;
  LAYER M2 ;
        RECT 3.516 21.068 3.588 21.1 ;
  LAYER M2 ;
        RECT 0.8 21.068 3.552 21.1 ;
  LAYER M1 ;
        RECT 0.784 21.048 0.816 21.12 ;
  LAYER M2 ;
        RECT 0.764 21.068 0.836 21.1 ;
  LAYER M1 ;
        RECT 3.536 17.94 3.568 18.012 ;
  LAYER M2 ;
        RECT 3.516 17.96 3.588 17.992 ;
  LAYER M2 ;
        RECT 0.8 17.96 3.552 17.992 ;
  LAYER M1 ;
        RECT 0.784 17.94 0.816 18.012 ;
  LAYER M2 ;
        RECT 0.764 17.96 0.836 17.992 ;
  LAYER M1 ;
        RECT 0.784 31.296 0.816 31.368 ;
  LAYER M2 ;
        RECT 0.764 31.316 0.836 31.348 ;
  LAYER M1 ;
        RECT 0.784 30.744 0.816 31.332 ;
  LAYER M1 ;
        RECT 0.784 17.976 0.816 30.744 ;
  LAYER M1 ;
        RECT 15.44 30.372 15.472 30.444 ;
  LAYER M2 ;
        RECT 15.42 30.392 15.492 30.424 ;
  LAYER M1 ;
        RECT 15.44 30.408 15.472 30.576 ;
  LAYER M1 ;
        RECT 15.44 30.54 15.472 30.612 ;
  LAYER M2 ;
        RECT 15.42 30.56 15.492 30.592 ;
  LAYER M2 ;
        RECT 15.456 30.56 15.68 30.592 ;
  LAYER M1 ;
        RECT 15.664 30.54 15.696 30.612 ;
  LAYER M2 ;
        RECT 15.644 30.56 15.716 30.592 ;
  LAYER M1 ;
        RECT 15.44 27.264 15.472 27.336 ;
  LAYER M2 ;
        RECT 15.42 27.284 15.492 27.316 ;
  LAYER M1 ;
        RECT 15.44 27.3 15.472 27.468 ;
  LAYER M1 ;
        RECT 15.44 27.432 15.472 27.504 ;
  LAYER M2 ;
        RECT 15.42 27.452 15.492 27.484 ;
  LAYER M2 ;
        RECT 15.456 27.452 15.68 27.484 ;
  LAYER M1 ;
        RECT 15.664 27.432 15.696 27.504 ;
  LAYER M2 ;
        RECT 15.644 27.452 15.716 27.484 ;
  LAYER M1 ;
        RECT 15.44 24.156 15.472 24.228 ;
  LAYER M2 ;
        RECT 15.42 24.176 15.492 24.208 ;
  LAYER M1 ;
        RECT 15.44 24.192 15.472 24.36 ;
  LAYER M1 ;
        RECT 15.44 24.324 15.472 24.396 ;
  LAYER M2 ;
        RECT 15.42 24.344 15.492 24.376 ;
  LAYER M2 ;
        RECT 15.456 24.344 15.68 24.376 ;
  LAYER M1 ;
        RECT 15.664 24.324 15.696 24.396 ;
  LAYER M2 ;
        RECT 15.644 24.344 15.716 24.376 ;
  LAYER M1 ;
        RECT 15.44 21.048 15.472 21.12 ;
  LAYER M2 ;
        RECT 15.42 21.068 15.492 21.1 ;
  LAYER M1 ;
        RECT 15.44 21.084 15.472 21.252 ;
  LAYER M1 ;
        RECT 15.44 21.216 15.472 21.288 ;
  LAYER M2 ;
        RECT 15.42 21.236 15.492 21.268 ;
  LAYER M2 ;
        RECT 15.456 21.236 15.68 21.268 ;
  LAYER M1 ;
        RECT 15.664 21.216 15.696 21.288 ;
  LAYER M2 ;
        RECT 15.644 21.236 15.716 21.268 ;
  LAYER M1 ;
        RECT 15.44 17.94 15.472 18.012 ;
  LAYER M2 ;
        RECT 15.42 17.96 15.492 17.992 ;
  LAYER M1 ;
        RECT 15.44 17.976 15.472 18.144 ;
  LAYER M1 ;
        RECT 15.44 18.108 15.472 18.18 ;
  LAYER M2 ;
        RECT 15.42 18.128 15.492 18.16 ;
  LAYER M2 ;
        RECT 15.456 18.128 15.68 18.16 ;
  LAYER M1 ;
        RECT 15.664 18.108 15.696 18.18 ;
  LAYER M2 ;
        RECT 15.644 18.128 15.716 18.16 ;
  LAYER M1 ;
        RECT 15.664 31.296 15.696 31.368 ;
  LAYER M2 ;
        RECT 15.644 31.316 15.716 31.348 ;
  LAYER M1 ;
        RECT 15.664 30.744 15.696 31.332 ;
  LAYER M1 ;
        RECT 15.664 18.144 15.696 30.744 ;
  LAYER M2 ;
        RECT 0.8 31.316 15.68 31.348 ;
  LAYER M1 ;
        RECT 6.512 30.372 6.544 30.444 ;
  LAYER M2 ;
        RECT 6.492 30.392 6.564 30.424 ;
  LAYER M2 ;
        RECT 3.552 30.392 6.528 30.424 ;
  LAYER M1 ;
        RECT 3.536 30.372 3.568 30.444 ;
  LAYER M2 ;
        RECT 3.516 30.392 3.588 30.424 ;
  LAYER M1 ;
        RECT 6.512 17.94 6.544 18.012 ;
  LAYER M2 ;
        RECT 6.492 17.96 6.564 17.992 ;
  LAYER M2 ;
        RECT 3.552 17.96 6.528 17.992 ;
  LAYER M1 ;
        RECT 3.536 17.94 3.568 18.012 ;
  LAYER M2 ;
        RECT 3.516 17.96 3.588 17.992 ;
  LAYER M1 ;
        RECT 9.488 17.94 9.52 18.012 ;
  LAYER M2 ;
        RECT 9.468 17.96 9.54 17.992 ;
  LAYER M2 ;
        RECT 6.528 17.96 9.504 17.992 ;
  LAYER M1 ;
        RECT 6.512 17.94 6.544 18.012 ;
  LAYER M2 ;
        RECT 6.492 17.96 6.564 17.992 ;
  LAYER M1 ;
        RECT 12.464 17.94 12.496 18.012 ;
  LAYER M2 ;
        RECT 12.444 17.96 12.516 17.992 ;
  LAYER M2 ;
        RECT 9.504 17.96 12.48 17.992 ;
  LAYER M1 ;
        RECT 9.488 17.94 9.52 18.012 ;
  LAYER M2 ;
        RECT 9.468 17.96 9.54 17.992 ;
  LAYER M1 ;
        RECT 12.464 30.372 12.496 30.444 ;
  LAYER M2 ;
        RECT 12.444 30.392 12.516 30.424 ;
  LAYER M2 ;
        RECT 12.48 30.392 15.456 30.424 ;
  LAYER M1 ;
        RECT 15.44 30.372 15.472 30.444 ;
  LAYER M2 ;
        RECT 15.42 30.392 15.492 30.424 ;
  LAYER M1 ;
        RECT 9.488 30.372 9.52 30.444 ;
  LAYER M2 ;
        RECT 9.468 30.392 9.54 30.424 ;
  LAYER M2 ;
        RECT 9.504 30.392 12.48 30.424 ;
  LAYER M1 ;
        RECT 12.464 30.372 12.496 30.444 ;
  LAYER M2 ;
        RECT 12.444 30.392 12.516 30.424 ;
  LAYER M1 ;
        RECT 7.12 21.72 7.152 21.792 ;
  LAYER M2 ;
        RECT 7.1 21.74 7.172 21.772 ;
  LAYER M2 ;
        RECT 6.912 21.74 7.136 21.772 ;
  LAYER M1 ;
        RECT 6.896 21.72 6.928 21.792 ;
  LAYER M2 ;
        RECT 6.876 21.74 6.948 21.772 ;
  LAYER M1 ;
        RECT 4.144 18.612 4.176 18.684 ;
  LAYER M2 ;
        RECT 4.124 18.632 4.196 18.664 ;
  LAYER M1 ;
        RECT 4.144 18.48 4.176 18.648 ;
  LAYER M1 ;
        RECT 4.144 18.444 4.176 18.516 ;
  LAYER M2 ;
        RECT 4.124 18.464 4.196 18.496 ;
  LAYER M2 ;
        RECT 4.16 18.464 6.912 18.496 ;
  LAYER M1 ;
        RECT 6.896 18.444 6.928 18.516 ;
  LAYER M2 ;
        RECT 6.876 18.464 6.948 18.496 ;
  LAYER M1 ;
        RECT 6.896 14.916 6.928 14.988 ;
  LAYER M2 ;
        RECT 6.876 14.936 6.948 14.968 ;
  LAYER M1 ;
        RECT 6.896 14.952 6.928 15.204 ;
  LAYER M1 ;
        RECT 6.896 15.204 6.928 21.756 ;
  LAYER M1 ;
        RECT 10.096 24.828 10.128 24.9 ;
  LAYER M2 ;
        RECT 10.076 24.848 10.148 24.88 ;
  LAYER M2 ;
        RECT 9.888 24.848 10.112 24.88 ;
  LAYER M1 ;
        RECT 9.872 24.828 9.904 24.9 ;
  LAYER M2 ;
        RECT 9.852 24.848 9.924 24.88 ;
  LAYER M1 ;
        RECT 9.872 14.916 9.904 14.988 ;
  LAYER M2 ;
        RECT 9.852 14.936 9.924 14.968 ;
  LAYER M1 ;
        RECT 9.872 14.952 9.904 15.204 ;
  LAYER M1 ;
        RECT 9.872 15.204 9.904 24.864 ;
  LAYER M2 ;
        RECT 6.912 14.936 9.888 14.968 ;
  LAYER M1 ;
        RECT 4.144 21.72 4.176 21.792 ;
  LAYER M2 ;
        RECT 4.124 21.74 4.196 21.772 ;
  LAYER M2 ;
        RECT 3.936 21.74 4.16 21.772 ;
  LAYER M1 ;
        RECT 3.92 21.72 3.952 21.792 ;
  LAYER M2 ;
        RECT 3.9 21.74 3.972 21.772 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 24.9 ;
  LAYER M2 ;
        RECT 4.124 24.848 4.196 24.88 ;
  LAYER M2 ;
        RECT 3.936 24.848 4.16 24.88 ;
  LAYER M1 ;
        RECT 3.92 24.828 3.952 24.9 ;
  LAYER M2 ;
        RECT 3.9 24.848 3.972 24.88 ;
  LAYER M1 ;
        RECT 3.92 14.748 3.952 14.82 ;
  LAYER M2 ;
        RECT 3.9 14.768 3.972 14.8 ;
  LAYER M1 ;
        RECT 3.92 14.784 3.952 15.204 ;
  LAYER M1 ;
        RECT 3.92 15.204 3.952 24.864 ;
  LAYER M1 ;
        RECT 10.096 21.72 10.128 21.792 ;
  LAYER M2 ;
        RECT 10.076 21.74 10.148 21.772 ;
  LAYER M1 ;
        RECT 10.096 21.588 10.128 21.756 ;
  LAYER M1 ;
        RECT 10.096 21.552 10.128 21.624 ;
  LAYER M2 ;
        RECT 10.076 21.572 10.148 21.604 ;
  LAYER M2 ;
        RECT 10.112 21.572 12.864 21.604 ;
  LAYER M1 ;
        RECT 12.848 21.552 12.88 21.624 ;
  LAYER M2 ;
        RECT 12.828 21.572 12.9 21.604 ;
  LAYER M1 ;
        RECT 10.096 18.612 10.128 18.684 ;
  LAYER M2 ;
        RECT 10.076 18.632 10.148 18.664 ;
  LAYER M1 ;
        RECT 10.096 18.48 10.128 18.648 ;
  LAYER M1 ;
        RECT 10.096 18.444 10.128 18.516 ;
  LAYER M2 ;
        RECT 10.076 18.464 10.148 18.496 ;
  LAYER M2 ;
        RECT 10.112 18.464 12.864 18.496 ;
  LAYER M1 ;
        RECT 12.848 18.444 12.88 18.516 ;
  LAYER M2 ;
        RECT 12.828 18.464 12.9 18.496 ;
  LAYER M1 ;
        RECT 12.848 14.748 12.88 14.82 ;
  LAYER M2 ;
        RECT 12.828 14.768 12.9 14.8 ;
  LAYER M1 ;
        RECT 12.848 14.784 12.88 15.204 ;
  LAYER M1 ;
        RECT 12.848 15.204 12.88 21.588 ;
  LAYER M2 ;
        RECT 3.936 14.768 12.864 14.8 ;
  LAYER M1 ;
        RECT 7.12 24.828 7.152 24.9 ;
  LAYER M2 ;
        RECT 7.1 24.848 7.172 24.88 ;
  LAYER M2 ;
        RECT 4.16 24.848 7.136 24.88 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 24.9 ;
  LAYER M2 ;
        RECT 4.124 24.848 4.196 24.88 ;
  LAYER M1 ;
        RECT 7.12 18.612 7.152 18.684 ;
  LAYER M2 ;
        RECT 7.1 18.632 7.172 18.664 ;
  LAYER M2 ;
        RECT 7.136 18.632 10.112 18.664 ;
  LAYER M1 ;
        RECT 10.096 18.612 10.128 18.684 ;
  LAYER M2 ;
        RECT 10.076 18.632 10.148 18.664 ;
  LAYER M1 ;
        RECT 1.168 27.936 1.2 28.008 ;
  LAYER M2 ;
        RECT 1.148 27.956 1.22 27.988 ;
  LAYER M2 ;
        RECT 0.96 27.956 1.184 27.988 ;
  LAYER M1 ;
        RECT 0.944 27.936 0.976 28.008 ;
  LAYER M2 ;
        RECT 0.924 27.956 0.996 27.988 ;
  LAYER M1 ;
        RECT 1.168 24.828 1.2 24.9 ;
  LAYER M2 ;
        RECT 1.148 24.848 1.22 24.88 ;
  LAYER M2 ;
        RECT 0.96 24.848 1.184 24.88 ;
  LAYER M1 ;
        RECT 0.944 24.828 0.976 24.9 ;
  LAYER M2 ;
        RECT 0.924 24.848 0.996 24.88 ;
  LAYER M1 ;
        RECT 1.168 21.72 1.2 21.792 ;
  LAYER M2 ;
        RECT 1.148 21.74 1.22 21.772 ;
  LAYER M2 ;
        RECT 0.96 21.74 1.184 21.772 ;
  LAYER M1 ;
        RECT 0.944 21.72 0.976 21.792 ;
  LAYER M2 ;
        RECT 0.924 21.74 0.996 21.772 ;
  LAYER M1 ;
        RECT 1.168 18.612 1.2 18.684 ;
  LAYER M2 ;
        RECT 1.148 18.632 1.22 18.664 ;
  LAYER M2 ;
        RECT 0.96 18.632 1.184 18.664 ;
  LAYER M1 ;
        RECT 0.944 18.612 0.976 18.684 ;
  LAYER M2 ;
        RECT 0.924 18.632 0.996 18.664 ;
  LAYER M1 ;
        RECT 1.168 15.504 1.2 15.576 ;
  LAYER M2 ;
        RECT 1.148 15.524 1.22 15.556 ;
  LAYER M2 ;
        RECT 0.96 15.524 1.184 15.556 ;
  LAYER M1 ;
        RECT 0.944 15.504 0.976 15.576 ;
  LAYER M2 ;
        RECT 0.924 15.524 0.996 15.556 ;
  LAYER M1 ;
        RECT 0.944 14.58 0.976 14.652 ;
  LAYER M2 ;
        RECT 0.924 14.6 0.996 14.632 ;
  LAYER M1 ;
        RECT 0.944 14.616 0.976 15.204 ;
  LAYER M1 ;
        RECT 0.944 15.204 0.976 27.972 ;
  LAYER M1 ;
        RECT 13.072 27.936 13.104 28.008 ;
  LAYER M2 ;
        RECT 13.052 27.956 13.124 27.988 ;
  LAYER M1 ;
        RECT 13.072 27.804 13.104 27.972 ;
  LAYER M1 ;
        RECT 13.072 27.768 13.104 27.84 ;
  LAYER M2 ;
        RECT 13.052 27.788 13.124 27.82 ;
  LAYER M2 ;
        RECT 13.088 27.788 15.84 27.82 ;
  LAYER M1 ;
        RECT 15.824 27.768 15.856 27.84 ;
  LAYER M2 ;
        RECT 15.804 27.788 15.876 27.82 ;
  LAYER M1 ;
        RECT 13.072 24.828 13.104 24.9 ;
  LAYER M2 ;
        RECT 13.052 24.848 13.124 24.88 ;
  LAYER M1 ;
        RECT 13.072 24.696 13.104 24.864 ;
  LAYER M1 ;
        RECT 13.072 24.66 13.104 24.732 ;
  LAYER M2 ;
        RECT 13.052 24.68 13.124 24.712 ;
  LAYER M2 ;
        RECT 13.088 24.68 15.84 24.712 ;
  LAYER M1 ;
        RECT 15.824 24.66 15.856 24.732 ;
  LAYER M2 ;
        RECT 15.804 24.68 15.876 24.712 ;
  LAYER M1 ;
        RECT 13.072 21.72 13.104 21.792 ;
  LAYER M2 ;
        RECT 13.052 21.74 13.124 21.772 ;
  LAYER M1 ;
        RECT 13.072 21.588 13.104 21.756 ;
  LAYER M1 ;
        RECT 13.072 21.552 13.104 21.624 ;
  LAYER M2 ;
        RECT 13.052 21.572 13.124 21.604 ;
  LAYER M2 ;
        RECT 13.088 21.572 15.84 21.604 ;
  LAYER M1 ;
        RECT 15.824 21.552 15.856 21.624 ;
  LAYER M2 ;
        RECT 15.804 21.572 15.876 21.604 ;
  LAYER M1 ;
        RECT 13.072 18.612 13.104 18.684 ;
  LAYER M2 ;
        RECT 13.052 18.632 13.124 18.664 ;
  LAYER M1 ;
        RECT 13.072 18.48 13.104 18.648 ;
  LAYER M1 ;
        RECT 13.072 18.444 13.104 18.516 ;
  LAYER M2 ;
        RECT 13.052 18.464 13.124 18.496 ;
  LAYER M2 ;
        RECT 13.088 18.464 15.84 18.496 ;
  LAYER M1 ;
        RECT 15.824 18.444 15.856 18.516 ;
  LAYER M2 ;
        RECT 15.804 18.464 15.876 18.496 ;
  LAYER M1 ;
        RECT 13.072 15.504 13.104 15.576 ;
  LAYER M2 ;
        RECT 13.052 15.524 13.124 15.556 ;
  LAYER M1 ;
        RECT 13.072 15.372 13.104 15.54 ;
  LAYER M1 ;
        RECT 13.072 15.336 13.104 15.408 ;
  LAYER M2 ;
        RECT 13.052 15.356 13.124 15.388 ;
  LAYER M2 ;
        RECT 13.088 15.356 15.84 15.388 ;
  LAYER M1 ;
        RECT 15.824 15.336 15.856 15.408 ;
  LAYER M2 ;
        RECT 15.804 15.356 15.876 15.388 ;
  LAYER M1 ;
        RECT 15.824 14.58 15.856 14.652 ;
  LAYER M2 ;
        RECT 15.804 14.6 15.876 14.632 ;
  LAYER M1 ;
        RECT 15.824 14.616 15.856 15.204 ;
  LAYER M1 ;
        RECT 15.824 15.204 15.856 27.804 ;
  LAYER M2 ;
        RECT 0.96 14.6 15.84 14.632 ;
  LAYER M1 ;
        RECT 4.144 27.936 4.176 28.008 ;
  LAYER M2 ;
        RECT 4.124 27.956 4.196 27.988 ;
  LAYER M2 ;
        RECT 1.184 27.956 4.16 27.988 ;
  LAYER M1 ;
        RECT 1.168 27.936 1.2 28.008 ;
  LAYER M2 ;
        RECT 1.148 27.956 1.22 27.988 ;
  LAYER M1 ;
        RECT 4.144 15.504 4.176 15.576 ;
  LAYER M2 ;
        RECT 4.124 15.524 4.196 15.556 ;
  LAYER M2 ;
        RECT 1.184 15.524 4.16 15.556 ;
  LAYER M1 ;
        RECT 1.168 15.504 1.2 15.576 ;
  LAYER M2 ;
        RECT 1.148 15.524 1.22 15.556 ;
  LAYER M1 ;
        RECT 7.12 15.504 7.152 15.576 ;
  LAYER M2 ;
        RECT 7.1 15.524 7.172 15.556 ;
  LAYER M2 ;
        RECT 4.16 15.524 7.136 15.556 ;
  LAYER M1 ;
        RECT 4.144 15.504 4.176 15.576 ;
  LAYER M2 ;
        RECT 4.124 15.524 4.196 15.556 ;
  LAYER M1 ;
        RECT 10.096 15.504 10.128 15.576 ;
  LAYER M2 ;
        RECT 10.076 15.524 10.148 15.556 ;
  LAYER M2 ;
        RECT 7.136 15.524 10.112 15.556 ;
  LAYER M1 ;
        RECT 7.12 15.504 7.152 15.576 ;
  LAYER M2 ;
        RECT 7.1 15.524 7.172 15.556 ;
  LAYER M1 ;
        RECT 10.096 27.936 10.128 28.008 ;
  LAYER M2 ;
        RECT 10.076 27.956 10.148 27.988 ;
  LAYER M2 ;
        RECT 10.112 27.956 13.088 27.988 ;
  LAYER M1 ;
        RECT 13.072 27.936 13.104 28.008 ;
  LAYER M2 ;
        RECT 13.052 27.956 13.124 27.988 ;
  LAYER M1 ;
        RECT 7.12 27.936 7.152 28.008 ;
  LAYER M2 ;
        RECT 7.1 27.956 7.172 27.988 ;
  LAYER M2 ;
        RECT 7.136 27.956 10.112 27.988 ;
  LAYER M1 ;
        RECT 10.096 27.936 10.128 28.008 ;
  LAYER M2 ;
        RECT 10.076 27.956 10.148 27.988 ;
  LAYER M1 ;
        RECT 1.12 27.888 3.616 30.492 ;
  LAYER M3 ;
        RECT 1.12 27.888 3.616 30.492 ;
  LAYER M2 ;
        RECT 1.12 27.888 3.616 30.492 ;
  LAYER M1 ;
        RECT 1.12 24.78 3.616 27.384 ;
  LAYER M3 ;
        RECT 1.12 24.78 3.616 27.384 ;
  LAYER M2 ;
        RECT 1.12 24.78 3.616 27.384 ;
  LAYER M1 ;
        RECT 1.12 21.672 3.616 24.276 ;
  LAYER M3 ;
        RECT 1.12 21.672 3.616 24.276 ;
  LAYER M2 ;
        RECT 1.12 21.672 3.616 24.276 ;
  LAYER M1 ;
        RECT 1.12 18.564 3.616 21.168 ;
  LAYER M3 ;
        RECT 1.12 18.564 3.616 21.168 ;
  LAYER M2 ;
        RECT 1.12 18.564 3.616 21.168 ;
  LAYER M1 ;
        RECT 1.12 15.456 3.616 18.06 ;
  LAYER M3 ;
        RECT 1.12 15.456 3.616 18.06 ;
  LAYER M2 ;
        RECT 1.12 15.456 3.616 18.06 ;
  LAYER M1 ;
        RECT 4.096 27.888 6.592 30.492 ;
  LAYER M3 ;
        RECT 4.096 27.888 6.592 30.492 ;
  LAYER M2 ;
        RECT 4.096 27.888 6.592 30.492 ;
  LAYER M1 ;
        RECT 4.096 24.78 6.592 27.384 ;
  LAYER M3 ;
        RECT 4.096 24.78 6.592 27.384 ;
  LAYER M2 ;
        RECT 4.096 24.78 6.592 27.384 ;
  LAYER M1 ;
        RECT 4.096 21.672 6.592 24.276 ;
  LAYER M3 ;
        RECT 4.096 21.672 6.592 24.276 ;
  LAYER M2 ;
        RECT 4.096 21.672 6.592 24.276 ;
  LAYER M1 ;
        RECT 4.096 18.564 6.592 21.168 ;
  LAYER M3 ;
        RECT 4.096 18.564 6.592 21.168 ;
  LAYER M2 ;
        RECT 4.096 18.564 6.592 21.168 ;
  LAYER M1 ;
        RECT 4.096 15.456 6.592 18.06 ;
  LAYER M3 ;
        RECT 4.096 15.456 6.592 18.06 ;
  LAYER M2 ;
        RECT 4.096 15.456 6.592 18.06 ;
  LAYER M1 ;
        RECT 7.072 27.888 9.568 30.492 ;
  LAYER M3 ;
        RECT 7.072 27.888 9.568 30.492 ;
  LAYER M2 ;
        RECT 7.072 27.888 9.568 30.492 ;
  LAYER M1 ;
        RECT 7.072 24.78 9.568 27.384 ;
  LAYER M3 ;
        RECT 7.072 24.78 9.568 27.384 ;
  LAYER M2 ;
        RECT 7.072 24.78 9.568 27.384 ;
  LAYER M1 ;
        RECT 7.072 21.672 9.568 24.276 ;
  LAYER M3 ;
        RECT 7.072 21.672 9.568 24.276 ;
  LAYER M2 ;
        RECT 7.072 21.672 9.568 24.276 ;
  LAYER M1 ;
        RECT 7.072 18.564 9.568 21.168 ;
  LAYER M3 ;
        RECT 7.072 18.564 9.568 21.168 ;
  LAYER M2 ;
        RECT 7.072 18.564 9.568 21.168 ;
  LAYER M1 ;
        RECT 7.072 15.456 9.568 18.06 ;
  LAYER M3 ;
        RECT 7.072 15.456 9.568 18.06 ;
  LAYER M2 ;
        RECT 7.072 15.456 9.568 18.06 ;
  LAYER M1 ;
        RECT 10.048 27.888 12.544 30.492 ;
  LAYER M3 ;
        RECT 10.048 27.888 12.544 30.492 ;
  LAYER M2 ;
        RECT 10.048 27.888 12.544 30.492 ;
  LAYER M1 ;
        RECT 10.048 24.78 12.544 27.384 ;
  LAYER M3 ;
        RECT 10.048 24.78 12.544 27.384 ;
  LAYER M2 ;
        RECT 10.048 24.78 12.544 27.384 ;
  LAYER M1 ;
        RECT 10.048 21.672 12.544 24.276 ;
  LAYER M3 ;
        RECT 10.048 21.672 12.544 24.276 ;
  LAYER M2 ;
        RECT 10.048 21.672 12.544 24.276 ;
  LAYER M1 ;
        RECT 10.048 18.564 12.544 21.168 ;
  LAYER M3 ;
        RECT 10.048 18.564 12.544 21.168 ;
  LAYER M2 ;
        RECT 10.048 18.564 12.544 21.168 ;
  LAYER M1 ;
        RECT 10.048 15.456 12.544 18.06 ;
  LAYER M3 ;
        RECT 10.048 15.456 12.544 18.06 ;
  LAYER M2 ;
        RECT 10.048 15.456 12.544 18.06 ;
  LAYER M1 ;
        RECT 13.024 27.888 15.52 30.492 ;
  LAYER M3 ;
        RECT 13.024 27.888 15.52 30.492 ;
  LAYER M2 ;
        RECT 13.024 27.888 15.52 30.492 ;
  LAYER M1 ;
        RECT 13.024 24.78 15.52 27.384 ;
  LAYER M3 ;
        RECT 13.024 24.78 15.52 27.384 ;
  LAYER M2 ;
        RECT 13.024 24.78 15.52 27.384 ;
  LAYER M1 ;
        RECT 13.024 21.672 15.52 24.276 ;
  LAYER M3 ;
        RECT 13.024 21.672 15.52 24.276 ;
  LAYER M2 ;
        RECT 13.024 21.672 15.52 24.276 ;
  LAYER M1 ;
        RECT 13.024 18.564 15.52 21.168 ;
  LAYER M3 ;
        RECT 13.024 18.564 15.52 21.168 ;
  LAYER M2 ;
        RECT 13.024 18.564 15.52 21.168 ;
  LAYER M1 ;
        RECT 13.024 15.456 15.52 18.06 ;
  LAYER M3 ;
        RECT 13.024 15.456 15.52 18.06 ;
  LAYER M2 ;
        RECT 13.024 15.456 15.52 18.06 ;
  END 
END switched_capacitor_combination
