.subckt common_source vin vop vcc vss
mp0 vop vop vcc vcc p w=720e-9 nf=4 m=4
mn0 vop vin vss vss n w=720e-9 nf=4 m=4
.ends common_source
