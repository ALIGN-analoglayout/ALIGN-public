MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 18.08 BY 16.884 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
      LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
      LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
      LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
      LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
      LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
      LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
      LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
      LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
      LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
      LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
      LAYER M2 ;
        RECT 6.032 0.236 11.984 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M1 ;
        RECT 8.768 7.056 8.8 7.224 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M2 ;
        RECT 8.784 7.04 9.008 7.072 ;
  LAYER M1 ;
        RECT 8.992 7.02 9.024 7.092 ;
  LAYER M2 ;
        RECT 8.972 7.04 9.044 7.072 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M2 ;
        RECT 9.008 7.208 11.76 7.24 ;
  LAYER M1 ;
        RECT 8.992 7.188 9.024 7.26 ;
  LAYER M2 ;
        RECT 8.972 7.208 9.044 7.24 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.164 8.8 10.332 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M2 ;
        RECT 8.784 10.148 9.008 10.18 ;
  LAYER M1 ;
        RECT 8.992 10.128 9.024 10.2 ;
  LAYER M2 ;
        RECT 8.972 10.148 9.044 10.18 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M2 ;
        RECT 9.008 4.1 11.76 4.132 ;
  LAYER M1 ;
        RECT 8.992 4.08 9.024 4.152 ;
  LAYER M2 ;
        RECT 8.972 4.1 9.044 4.132 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M1 ;
        RECT 8.768 3.948 8.8 4.116 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 8.784 3.932 9.008 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M2 ;
        RECT 9.008 10.316 11.76 10.348 ;
  LAYER M1 ;
        RECT 8.992 10.296 9.024 10.368 ;
  LAYER M2 ;
        RECT 8.972 10.316 9.044 10.348 ;
  LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
  LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
  LAYER M1 ;
        RECT 8.992 0.42 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 10.332 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M1 ;
        RECT 5.792 7.056 5.824 7.224 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M2 ;
        RECT 5.808 7.04 6.032 7.072 ;
  LAYER M1 ;
        RECT 6.016 7.02 6.048 7.092 ;
  LAYER M2 ;
        RECT 5.996 7.04 6.068 7.072 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.164 5.824 10.332 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M1 ;
        RECT 5.792 3.948 5.824 4.116 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M2 ;
        RECT 5.808 3.932 6.032 3.964 ;
  LAYER M1 ;
        RECT 6.016 3.912 6.048 3.984 ;
  LAYER M2 ;
        RECT 5.996 3.932 6.068 3.964 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 10.164 ;
  LAYER M1 ;
        RECT 14.72 7.188 14.752 7.26 ;
  LAYER M2 ;
        RECT 14.7 7.208 14.772 7.24 ;
  LAYER M2 ;
        RECT 11.984 7.208 14.736 7.24 ;
  LAYER M1 ;
        RECT 11.968 7.188 12 7.26 ;
  LAYER M2 ;
        RECT 11.948 7.208 12.02 7.24 ;
  LAYER M1 ;
        RECT 14.72 4.08 14.752 4.152 ;
  LAYER M2 ;
        RECT 14.7 4.1 14.772 4.132 ;
  LAYER M2 ;
        RECT 11.984 4.1 14.736 4.132 ;
  LAYER M1 ;
        RECT 11.968 4.08 12 4.152 ;
  LAYER M2 ;
        RECT 11.948 4.1 12.02 4.132 ;
  LAYER M1 ;
        RECT 14.72 10.296 14.752 10.368 ;
  LAYER M2 ;
        RECT 14.7 10.316 14.772 10.348 ;
  LAYER M2 ;
        RECT 11.984 10.316 14.736 10.348 ;
  LAYER M1 ;
        RECT 11.968 10.296 12 10.368 ;
  LAYER M2 ;
        RECT 11.948 10.316 12.02 10.348 ;
  LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
  LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
  LAYER M1 ;
        RECT 11.968 0.252 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 10.332 ;
  LAYER M2 ;
        RECT 6.032 0.236 11.984 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.84 2.848 1.008 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M2 ;
        RECT 2.832 0.824 3.056 0.856 ;
  LAYER M1 ;
        RECT 3.04 0.804 3.072 0.876 ;
  LAYER M2 ;
        RECT 3.02 0.824 3.092 0.856 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M1 ;
        RECT 2.816 3.948 2.848 4.116 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M2 ;
        RECT 2.832 3.932 3.056 3.964 ;
  LAYER M1 ;
        RECT 3.04 3.912 3.072 3.984 ;
  LAYER M2 ;
        RECT 3.02 3.932 3.092 3.964 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M1 ;
        RECT 2.816 7.056 2.848 7.224 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M2 ;
        RECT 2.832 7.04 3.056 7.072 ;
  LAYER M1 ;
        RECT 3.04 7.02 3.072 7.092 ;
  LAYER M2 ;
        RECT 3.02 7.04 3.092 7.072 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M1 ;
        RECT 2.816 10.164 2.848 10.332 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M2 ;
        RECT 2.832 10.148 3.056 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M1 ;
        RECT 2.816 13.272 2.848 13.44 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 13.308 ;
  LAYER M2 ;
        RECT 2.796 13.256 2.868 13.288 ;
  LAYER M2 ;
        RECT 2.832 13.256 3.056 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 3.056 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 3.04 0.972 3.072 1.044 ;
  LAYER M2 ;
        RECT 3.02 0.992 3.092 1.024 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M2 ;
        RECT 3.056 13.424 5.808 13.456 ;
  LAYER M1 ;
        RECT 3.04 13.404 3.072 13.476 ;
  LAYER M2 ;
        RECT 3.02 13.424 3.092 13.456 ;
  LAYER M1 ;
        RECT 3.04 0.048 3.072 0.12 ;
  LAYER M2 ;
        RECT 3.02 0.068 3.092 0.1 ;
  LAYER M1 ;
        RECT 3.04 0.084 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 13.44 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.84 14.752 1.008 ;
  LAYER M1 ;
        RECT 14.72 0.804 14.752 0.876 ;
  LAYER M2 ;
        RECT 14.7 0.824 14.772 0.856 ;
  LAYER M2 ;
        RECT 14.736 0.824 14.96 0.856 ;
  LAYER M1 ;
        RECT 14.944 0.804 14.976 0.876 ;
  LAYER M2 ;
        RECT 14.924 0.824 14.996 0.856 ;
  LAYER M1 ;
        RECT 14.72 13.404 14.752 13.476 ;
  LAYER M2 ;
        RECT 14.7 13.424 14.772 13.456 ;
  LAYER M1 ;
        RECT 14.72 13.272 14.752 13.44 ;
  LAYER M1 ;
        RECT 14.72 13.236 14.752 13.308 ;
  LAYER M2 ;
        RECT 14.7 13.256 14.772 13.288 ;
  LAYER M2 ;
        RECT 14.736 13.256 14.96 13.288 ;
  LAYER M1 ;
        RECT 14.944 13.236 14.976 13.308 ;
  LAYER M2 ;
        RECT 14.924 13.256 14.996 13.288 ;
  LAYER M1 ;
        RECT 17.696 0.972 17.728 1.044 ;
  LAYER M2 ;
        RECT 17.676 0.992 17.748 1.024 ;
  LAYER M2 ;
        RECT 14.96 0.992 17.712 1.024 ;
  LAYER M1 ;
        RECT 14.944 0.972 14.976 1.044 ;
  LAYER M2 ;
        RECT 14.924 0.992 14.996 1.024 ;
  LAYER M1 ;
        RECT 17.696 4.08 17.728 4.152 ;
  LAYER M2 ;
        RECT 17.676 4.1 17.748 4.132 ;
  LAYER M2 ;
        RECT 14.96 4.1 17.712 4.132 ;
  LAYER M1 ;
        RECT 14.944 4.08 14.976 4.152 ;
  LAYER M2 ;
        RECT 14.924 4.1 14.996 4.132 ;
  LAYER M1 ;
        RECT 17.696 7.188 17.728 7.26 ;
  LAYER M2 ;
        RECT 17.676 7.208 17.748 7.24 ;
  LAYER M2 ;
        RECT 14.96 7.208 17.712 7.24 ;
  LAYER M1 ;
        RECT 14.944 7.188 14.976 7.26 ;
  LAYER M2 ;
        RECT 14.924 7.208 14.996 7.24 ;
  LAYER M1 ;
        RECT 17.696 10.296 17.728 10.368 ;
  LAYER M2 ;
        RECT 17.676 10.316 17.748 10.348 ;
  LAYER M2 ;
        RECT 14.96 10.316 17.712 10.348 ;
  LAYER M1 ;
        RECT 14.944 10.296 14.976 10.368 ;
  LAYER M2 ;
        RECT 14.924 10.316 14.996 10.348 ;
  LAYER M1 ;
        RECT 17.696 13.404 17.728 13.476 ;
  LAYER M2 ;
        RECT 17.676 13.424 17.748 13.456 ;
  LAYER M2 ;
        RECT 14.96 13.424 17.712 13.456 ;
  LAYER M1 ;
        RECT 14.944 13.404 14.976 13.476 ;
  LAYER M2 ;
        RECT 14.924 13.424 14.996 13.456 ;
  LAYER M1 ;
        RECT 14.944 0.048 14.976 0.12 ;
  LAYER M2 ;
        RECT 14.924 0.068 14.996 0.1 ;
  LAYER M1 ;
        RECT 14.944 0.084 14.976 0.672 ;
  LAYER M1 ;
        RECT 14.944 0.672 14.976 13.44 ;
  LAYER M2 ;
        RECT 3.056 0.068 14.96 0.1 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M2 ;
        RECT 5.808 13.424 8.784 13.456 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 13.476 ;
  LAYER M2 ;
        RECT 11.724 13.424 11.796 13.456 ;
  LAYER M2 ;
        RECT 8.784 13.424 11.76 13.456 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M2 ;
        RECT 11.76 0.992 14.736 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M2 ;
        RECT 6.192 9.644 6.416 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 6.192 12.752 6.416 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.416 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
  LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
  LAYER M1 ;
        RECT 6.176 16.212 6.208 16.464 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 16.212 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M1 ;
        RECT 9.376 9.66 9.408 9.828 ;
  LAYER M1 ;
        RECT 9.376 9.792 9.408 9.864 ;
  LAYER M2 ;
        RECT 9.356 9.812 9.428 9.844 ;
  LAYER M2 ;
        RECT 9.392 9.812 12.144 9.844 ;
  LAYER M1 ;
        RECT 12.128 9.792 12.16 9.864 ;
  LAYER M2 ;
        RECT 12.108 9.812 12.18 9.844 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.376 6.552 9.408 6.72 ;
  LAYER M1 ;
        RECT 9.376 6.684 9.408 6.756 ;
  LAYER M2 ;
        RECT 9.356 6.704 9.428 6.736 ;
  LAYER M2 ;
        RECT 9.392 6.704 12.144 6.736 ;
  LAYER M1 ;
        RECT 12.128 6.684 12.16 6.756 ;
  LAYER M2 ;
        RECT 12.108 6.704 12.18 6.736 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M1 ;
        RECT 9.376 12.768 9.408 12.936 ;
  LAYER M1 ;
        RECT 9.376 12.9 9.408 12.972 ;
  LAYER M2 ;
        RECT 9.356 12.92 9.428 12.952 ;
  LAYER M2 ;
        RECT 9.392 12.92 12.144 12.952 ;
  LAYER M1 ;
        RECT 12.128 12.9 12.16 12.972 ;
  LAYER M2 ;
        RECT 12.108 12.92 12.18 12.952 ;
  LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
  LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
  LAYER M1 ;
        RECT 12.128 16.212 12.16 16.464 ;
  LAYER M1 ;
        RECT 12.128 6.72 12.16 16.212 ;
  LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.216 9.644 3.44 9.676 ;
  LAYER M1 ;
        RECT 3.2 9.624 3.232 9.696 ;
  LAYER M2 ;
        RECT 3.18 9.644 3.252 9.676 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 3.216 6.536 3.44 6.568 ;
  LAYER M1 ;
        RECT 3.2 6.516 3.232 6.588 ;
  LAYER M2 ;
        RECT 3.18 6.536 3.252 6.568 ;
  LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
  LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
  LAYER M1 ;
        RECT 3.2 16.212 3.232 16.632 ;
  LAYER M1 ;
        RECT 3.2 6.552 3.232 16.212 ;
  LAYER M1 ;
        RECT 12.352 9.624 12.384 9.696 ;
  LAYER M2 ;
        RECT 12.332 9.644 12.404 9.676 ;
  LAYER M1 ;
        RECT 12.352 9.66 12.384 9.828 ;
  LAYER M1 ;
        RECT 12.352 9.792 12.384 9.864 ;
  LAYER M2 ;
        RECT 12.332 9.812 12.404 9.844 ;
  LAYER M2 ;
        RECT 12.368 9.812 15.12 9.844 ;
  LAYER M1 ;
        RECT 15.104 9.792 15.136 9.864 ;
  LAYER M2 ;
        RECT 15.084 9.812 15.156 9.844 ;
  LAYER M1 ;
        RECT 12.352 6.516 12.384 6.588 ;
  LAYER M2 ;
        RECT 12.332 6.536 12.404 6.568 ;
  LAYER M1 ;
        RECT 12.352 6.552 12.384 6.72 ;
  LAYER M1 ;
        RECT 12.352 6.684 12.384 6.756 ;
  LAYER M2 ;
        RECT 12.332 6.704 12.404 6.736 ;
  LAYER M2 ;
        RECT 12.368 6.704 15.12 6.736 ;
  LAYER M1 ;
        RECT 15.104 6.684 15.136 6.756 ;
  LAYER M2 ;
        RECT 15.084 6.704 15.156 6.736 ;
  LAYER M1 ;
        RECT 12.352 12.732 12.384 12.804 ;
  LAYER M2 ;
        RECT 12.332 12.752 12.404 12.784 ;
  LAYER M1 ;
        RECT 12.352 12.768 12.384 12.936 ;
  LAYER M1 ;
        RECT 12.352 12.9 12.384 12.972 ;
  LAYER M2 ;
        RECT 12.332 12.92 12.404 12.952 ;
  LAYER M2 ;
        RECT 12.368 12.92 15.12 12.952 ;
  LAYER M1 ;
        RECT 15.104 12.9 15.136 12.972 ;
  LAYER M2 ;
        RECT 15.084 12.92 15.156 12.952 ;
  LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
  LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
  LAYER M1 ;
        RECT 15.104 16.212 15.136 16.632 ;
  LAYER M1 ;
        RECT 15.104 6.72 15.136 16.212 ;
  LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.08 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.064 3.408 0.096 3.48 ;
  LAYER M2 ;
        RECT 0.044 3.428 0.116 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.08 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.064 6.516 0.096 6.588 ;
  LAYER M2 ;
        RECT 0.044 6.536 0.116 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.08 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.064 9.624 0.096 9.696 ;
  LAYER M2 ;
        RECT 0.044 9.644 0.116 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.08 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.064 12.732 0.096 12.804 ;
  LAYER M2 ;
        RECT 0.044 12.752 0.116 12.784 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M2 ;
        RECT 0.08 15.86 0.464 15.892 ;
  LAYER M1 ;
        RECT 0.064 15.84 0.096 15.912 ;
  LAYER M2 ;
        RECT 0.044 15.86 0.116 15.892 ;
  LAYER M1 ;
        RECT 0.064 16.764 0.096 16.836 ;
  LAYER M2 ;
        RECT 0.044 16.784 0.116 16.816 ;
  LAYER M1 ;
        RECT 0.064 16.212 0.096 16.8 ;
  LAYER M1 ;
        RECT 0.064 3.444 0.096 16.212 ;
  LAYER M1 ;
        RECT 15.328 3.408 15.36 3.48 ;
  LAYER M2 ;
        RECT 15.308 3.428 15.38 3.46 ;
  LAYER M1 ;
        RECT 15.328 3.444 15.36 3.612 ;
  LAYER M1 ;
        RECT 15.328 3.576 15.36 3.648 ;
  LAYER M2 ;
        RECT 15.308 3.596 15.38 3.628 ;
  LAYER M2 ;
        RECT 15.344 3.596 17.936 3.628 ;
  LAYER M1 ;
        RECT 17.92 3.576 17.952 3.648 ;
  LAYER M2 ;
        RECT 17.9 3.596 17.972 3.628 ;
  LAYER M1 ;
        RECT 15.328 6.516 15.36 6.588 ;
  LAYER M2 ;
        RECT 15.308 6.536 15.38 6.568 ;
  LAYER M1 ;
        RECT 15.328 6.552 15.36 6.72 ;
  LAYER M1 ;
        RECT 15.328 6.684 15.36 6.756 ;
  LAYER M2 ;
        RECT 15.308 6.704 15.38 6.736 ;
  LAYER M2 ;
        RECT 15.344 6.704 17.936 6.736 ;
  LAYER M1 ;
        RECT 17.92 6.684 17.952 6.756 ;
  LAYER M2 ;
        RECT 17.9 6.704 17.972 6.736 ;
  LAYER M1 ;
        RECT 15.328 9.624 15.36 9.696 ;
  LAYER M2 ;
        RECT 15.308 9.644 15.38 9.676 ;
  LAYER M1 ;
        RECT 15.328 9.66 15.36 9.828 ;
  LAYER M1 ;
        RECT 15.328 9.792 15.36 9.864 ;
  LAYER M2 ;
        RECT 15.308 9.812 15.38 9.844 ;
  LAYER M2 ;
        RECT 15.344 9.812 17.936 9.844 ;
  LAYER M1 ;
        RECT 17.92 9.792 17.952 9.864 ;
  LAYER M2 ;
        RECT 17.9 9.812 17.972 9.844 ;
  LAYER M1 ;
        RECT 15.328 12.732 15.36 12.804 ;
  LAYER M2 ;
        RECT 15.308 12.752 15.38 12.784 ;
  LAYER M1 ;
        RECT 15.328 12.768 15.36 12.936 ;
  LAYER M1 ;
        RECT 15.328 12.9 15.36 12.972 ;
  LAYER M2 ;
        RECT 15.308 12.92 15.38 12.952 ;
  LAYER M2 ;
        RECT 15.344 12.92 17.936 12.952 ;
  LAYER M1 ;
        RECT 17.92 12.9 17.952 12.972 ;
  LAYER M2 ;
        RECT 17.9 12.92 17.972 12.952 ;
  LAYER M1 ;
        RECT 15.328 15.84 15.36 15.912 ;
  LAYER M2 ;
        RECT 15.308 15.86 15.38 15.892 ;
  LAYER M1 ;
        RECT 15.328 15.876 15.36 16.044 ;
  LAYER M1 ;
        RECT 15.328 16.008 15.36 16.08 ;
  LAYER M2 ;
        RECT 15.308 16.028 15.38 16.06 ;
  LAYER M2 ;
        RECT 15.344 16.028 17.936 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.008 17.952 16.08 ;
  LAYER M2 ;
        RECT 17.9 16.028 17.972 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.764 17.952 16.836 ;
  LAYER M2 ;
        RECT 17.9 16.784 17.972 16.816 ;
  LAYER M1 ;
        RECT 17.92 16.212 17.952 16.8 ;
  LAYER M1 ;
        RECT 17.92 3.612 17.952 16.212 ;
  LAYER M2 ;
        RECT 0.08 16.784 17.936 16.816 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 0.464 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M2 ;
        RECT 3.44 15.86 6.416 15.892 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M2 ;
        RECT 6.416 15.86 9.392 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M1 ;
        RECT 12.352 15.84 12.384 15.912 ;
  LAYER M2 ;
        RECT 12.332 15.86 12.404 15.892 ;
  LAYER M2 ;
        RECT 9.392 15.86 12.368 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M2 ;
        RECT 12.368 3.428 15.344 3.46 ;
  LAYER M1 ;
        RECT 15.328 3.408 15.36 3.48 ;
  LAYER M2 ;
        RECT 15.308 3.428 15.38 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M2 ;
        RECT 9.392 3.428 12.368 3.46 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.448 0.972 0.48 3.48 ;
  LAYER M3 ;
        RECT 0.448 3.428 0.48 3.46 ;
  LAYER M1 ;
        RECT 0.512 0.972 0.544 3.48 ;
  LAYER M3 ;
        RECT 0.512 0.992 0.544 1.024 ;
  LAYER M1 ;
        RECT 0.576 0.972 0.608 3.48 ;
  LAYER M3 ;
        RECT 0.576 3.428 0.608 3.46 ;
  LAYER M1 ;
        RECT 0.64 0.972 0.672 3.48 ;
  LAYER M3 ;
        RECT 0.64 0.992 0.672 1.024 ;
  LAYER M1 ;
        RECT 0.704 0.972 0.736 3.48 ;
  LAYER M3 ;
        RECT 0.704 3.428 0.736 3.46 ;
  LAYER M1 ;
        RECT 0.768 0.972 0.8 3.48 ;
  LAYER M3 ;
        RECT 0.768 0.992 0.8 1.024 ;
  LAYER M1 ;
        RECT 0.832 0.972 0.864 3.48 ;
  LAYER M3 ;
        RECT 0.832 3.428 0.864 3.46 ;
  LAYER M1 ;
        RECT 0.896 0.972 0.928 3.48 ;
  LAYER M3 ;
        RECT 0.896 0.992 0.928 1.024 ;
  LAYER M1 ;
        RECT 0.96 0.972 0.992 3.48 ;
  LAYER M3 ;
        RECT 0.96 3.428 0.992 3.46 ;
  LAYER M1 ;
        RECT 1.024 0.972 1.056 3.48 ;
  LAYER M3 ;
        RECT 1.024 0.992 1.056 1.024 ;
  LAYER M1 ;
        RECT 1.088 0.972 1.12 3.48 ;
  LAYER M3 ;
        RECT 1.088 3.428 1.12 3.46 ;
  LAYER M1 ;
        RECT 1.152 0.972 1.184 3.48 ;
  LAYER M3 ;
        RECT 1.152 0.992 1.184 1.024 ;
  LAYER M1 ;
        RECT 1.216 0.972 1.248 3.48 ;
  LAYER M3 ;
        RECT 1.216 3.428 1.248 3.46 ;
  LAYER M1 ;
        RECT 1.28 0.972 1.312 3.48 ;
  LAYER M3 ;
        RECT 1.28 0.992 1.312 1.024 ;
  LAYER M1 ;
        RECT 1.344 0.972 1.376 3.48 ;
  LAYER M3 ;
        RECT 1.344 3.428 1.376 3.46 ;
  LAYER M1 ;
        RECT 1.408 0.972 1.44 3.48 ;
  LAYER M3 ;
        RECT 1.408 0.992 1.44 1.024 ;
  LAYER M1 ;
        RECT 1.472 0.972 1.504 3.48 ;
  LAYER M3 ;
        RECT 1.472 3.428 1.504 3.46 ;
  LAYER M1 ;
        RECT 1.536 0.972 1.568 3.48 ;
  LAYER M3 ;
        RECT 1.536 0.992 1.568 1.024 ;
  LAYER M1 ;
        RECT 1.6 0.972 1.632 3.48 ;
  LAYER M3 ;
        RECT 1.6 3.428 1.632 3.46 ;
  LAYER M1 ;
        RECT 1.664 0.972 1.696 3.48 ;
  LAYER M3 ;
        RECT 1.664 0.992 1.696 1.024 ;
  LAYER M1 ;
        RECT 1.728 0.972 1.76 3.48 ;
  LAYER M3 ;
        RECT 1.728 3.428 1.76 3.46 ;
  LAYER M1 ;
        RECT 1.792 0.972 1.824 3.48 ;
  LAYER M3 ;
        RECT 1.792 0.992 1.824 1.024 ;
  LAYER M1 ;
        RECT 1.856 0.972 1.888 3.48 ;
  LAYER M3 ;
        RECT 1.856 3.428 1.888 3.46 ;
  LAYER M1 ;
        RECT 1.92 0.972 1.952 3.48 ;
  LAYER M3 ;
        RECT 1.92 0.992 1.952 1.024 ;
  LAYER M1 ;
        RECT 1.984 0.972 2.016 3.48 ;
  LAYER M3 ;
        RECT 1.984 3.428 2.016 3.46 ;
  LAYER M1 ;
        RECT 2.048 0.972 2.08 3.48 ;
  LAYER M3 ;
        RECT 2.048 0.992 2.08 1.024 ;
  LAYER M1 ;
        RECT 2.112 0.972 2.144 3.48 ;
  LAYER M3 ;
        RECT 2.112 3.428 2.144 3.46 ;
  LAYER M1 ;
        RECT 2.176 0.972 2.208 3.48 ;
  LAYER M3 ;
        RECT 2.176 0.992 2.208 1.024 ;
  LAYER M1 ;
        RECT 2.24 0.972 2.272 3.48 ;
  LAYER M3 ;
        RECT 2.24 3.428 2.272 3.46 ;
  LAYER M1 ;
        RECT 2.304 0.972 2.336 3.48 ;
  LAYER M3 ;
        RECT 2.304 0.992 2.336 1.024 ;
  LAYER M1 ;
        RECT 2.368 0.972 2.4 3.48 ;
  LAYER M3 ;
        RECT 2.368 3.428 2.4 3.46 ;
  LAYER M1 ;
        RECT 2.432 0.972 2.464 3.48 ;
  LAYER M3 ;
        RECT 2.432 0.992 2.464 1.024 ;
  LAYER M1 ;
        RECT 2.496 0.972 2.528 3.48 ;
  LAYER M3 ;
        RECT 2.496 3.428 2.528 3.46 ;
  LAYER M1 ;
        RECT 2.56 0.972 2.592 3.48 ;
  LAYER M3 ;
        RECT 2.56 0.992 2.592 1.024 ;
  LAYER M1 ;
        RECT 2.624 0.972 2.656 3.48 ;
  LAYER M3 ;
        RECT 2.624 3.428 2.656 3.46 ;
  LAYER M1 ;
        RECT 2.688 0.972 2.72 3.48 ;
  LAYER M3 ;
        RECT 2.688 0.992 2.72 1.024 ;
  LAYER M1 ;
        RECT 2.752 0.972 2.784 3.48 ;
  LAYER M3 ;
        RECT 2.752 3.428 2.784 3.46 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 3.48 ;
  LAYER M3 ;
        RECT 0.448 1.056 0.48 1.088 ;
  LAYER M2 ;
        RECT 2.816 1.12 2.848 1.152 ;
  LAYER M2 ;
        RECT 0.448 1.184 0.48 1.216 ;
  LAYER M2 ;
        RECT 2.816 1.248 2.848 1.28 ;
  LAYER M2 ;
        RECT 0.448 1.312 0.48 1.344 ;
  LAYER M2 ;
        RECT 2.816 1.376 2.848 1.408 ;
  LAYER M2 ;
        RECT 0.448 1.44 0.48 1.472 ;
  LAYER M2 ;
        RECT 2.816 1.504 2.848 1.536 ;
  LAYER M2 ;
        RECT 0.448 1.568 0.48 1.6 ;
  LAYER M2 ;
        RECT 2.816 1.632 2.848 1.664 ;
  LAYER M2 ;
        RECT 0.448 1.696 0.48 1.728 ;
  LAYER M2 ;
        RECT 2.816 1.76 2.848 1.792 ;
  LAYER M2 ;
        RECT 0.448 1.824 0.48 1.856 ;
  LAYER M2 ;
        RECT 2.816 1.888 2.848 1.92 ;
  LAYER M2 ;
        RECT 0.448 1.952 0.48 1.984 ;
  LAYER M2 ;
        RECT 2.816 2.016 2.848 2.048 ;
  LAYER M2 ;
        RECT 0.448 2.08 0.48 2.112 ;
  LAYER M2 ;
        RECT 2.816 2.144 2.848 2.176 ;
  LAYER M2 ;
        RECT 0.448 2.208 0.48 2.24 ;
  LAYER M2 ;
        RECT 2.816 2.272 2.848 2.304 ;
  LAYER M2 ;
        RECT 0.448 2.336 0.48 2.368 ;
  LAYER M2 ;
        RECT 2.816 2.4 2.848 2.432 ;
  LAYER M2 ;
        RECT 0.448 2.464 0.48 2.496 ;
  LAYER M2 ;
        RECT 2.816 2.528 2.848 2.56 ;
  LAYER M2 ;
        RECT 0.448 2.592 0.48 2.624 ;
  LAYER M2 ;
        RECT 2.816 2.656 2.848 2.688 ;
  LAYER M2 ;
        RECT 0.448 2.72 0.48 2.752 ;
  LAYER M2 ;
        RECT 2.816 2.784 2.848 2.816 ;
  LAYER M2 ;
        RECT 0.448 2.848 0.48 2.88 ;
  LAYER M2 ;
        RECT 2.816 2.912 2.848 2.944 ;
  LAYER M2 ;
        RECT 0.448 2.976 0.48 3.008 ;
  LAYER M2 ;
        RECT 2.816 3.04 2.848 3.072 ;
  LAYER M2 ;
        RECT 0.448 3.104 0.48 3.136 ;
  LAYER M2 ;
        RECT 2.816 3.168 2.848 3.2 ;
  LAYER M2 ;
        RECT 0.448 3.232 0.48 3.264 ;
  LAYER M2 ;
        RECT 2.816 3.296 2.848 3.328 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.448 4.08 0.48 6.588 ;
  LAYER M3 ;
        RECT 0.448 6.536 0.48 6.568 ;
  LAYER M1 ;
        RECT 0.512 4.08 0.544 6.588 ;
  LAYER M3 ;
        RECT 0.512 4.1 0.544 4.132 ;
  LAYER M1 ;
        RECT 0.576 4.08 0.608 6.588 ;
  LAYER M3 ;
        RECT 0.576 6.536 0.608 6.568 ;
  LAYER M1 ;
        RECT 0.64 4.08 0.672 6.588 ;
  LAYER M3 ;
        RECT 0.64 4.1 0.672 4.132 ;
  LAYER M1 ;
        RECT 0.704 4.08 0.736 6.588 ;
  LAYER M3 ;
        RECT 0.704 6.536 0.736 6.568 ;
  LAYER M1 ;
        RECT 0.768 4.08 0.8 6.588 ;
  LAYER M3 ;
        RECT 0.768 4.1 0.8 4.132 ;
  LAYER M1 ;
        RECT 0.832 4.08 0.864 6.588 ;
  LAYER M3 ;
        RECT 0.832 6.536 0.864 6.568 ;
  LAYER M1 ;
        RECT 0.896 4.08 0.928 6.588 ;
  LAYER M3 ;
        RECT 0.896 4.1 0.928 4.132 ;
  LAYER M1 ;
        RECT 0.96 4.08 0.992 6.588 ;
  LAYER M3 ;
        RECT 0.96 6.536 0.992 6.568 ;
  LAYER M1 ;
        RECT 1.024 4.08 1.056 6.588 ;
  LAYER M3 ;
        RECT 1.024 4.1 1.056 4.132 ;
  LAYER M1 ;
        RECT 1.088 4.08 1.12 6.588 ;
  LAYER M3 ;
        RECT 1.088 6.536 1.12 6.568 ;
  LAYER M1 ;
        RECT 1.152 4.08 1.184 6.588 ;
  LAYER M3 ;
        RECT 1.152 4.1 1.184 4.132 ;
  LAYER M1 ;
        RECT 1.216 4.08 1.248 6.588 ;
  LAYER M3 ;
        RECT 1.216 6.536 1.248 6.568 ;
  LAYER M1 ;
        RECT 1.28 4.08 1.312 6.588 ;
  LAYER M3 ;
        RECT 1.28 4.1 1.312 4.132 ;
  LAYER M1 ;
        RECT 1.344 4.08 1.376 6.588 ;
  LAYER M3 ;
        RECT 1.344 6.536 1.376 6.568 ;
  LAYER M1 ;
        RECT 1.408 4.08 1.44 6.588 ;
  LAYER M3 ;
        RECT 1.408 4.1 1.44 4.132 ;
  LAYER M1 ;
        RECT 1.472 4.08 1.504 6.588 ;
  LAYER M3 ;
        RECT 1.472 6.536 1.504 6.568 ;
  LAYER M1 ;
        RECT 1.536 4.08 1.568 6.588 ;
  LAYER M3 ;
        RECT 1.536 4.1 1.568 4.132 ;
  LAYER M1 ;
        RECT 1.6 4.08 1.632 6.588 ;
  LAYER M3 ;
        RECT 1.6 6.536 1.632 6.568 ;
  LAYER M1 ;
        RECT 1.664 4.08 1.696 6.588 ;
  LAYER M3 ;
        RECT 1.664 4.1 1.696 4.132 ;
  LAYER M1 ;
        RECT 1.728 4.08 1.76 6.588 ;
  LAYER M3 ;
        RECT 1.728 6.536 1.76 6.568 ;
  LAYER M1 ;
        RECT 1.792 4.08 1.824 6.588 ;
  LAYER M3 ;
        RECT 1.792 4.1 1.824 4.132 ;
  LAYER M1 ;
        RECT 1.856 4.08 1.888 6.588 ;
  LAYER M3 ;
        RECT 1.856 6.536 1.888 6.568 ;
  LAYER M1 ;
        RECT 1.92 4.08 1.952 6.588 ;
  LAYER M3 ;
        RECT 1.92 4.1 1.952 4.132 ;
  LAYER M1 ;
        RECT 1.984 4.08 2.016 6.588 ;
  LAYER M3 ;
        RECT 1.984 6.536 2.016 6.568 ;
  LAYER M1 ;
        RECT 2.048 4.08 2.08 6.588 ;
  LAYER M3 ;
        RECT 2.048 4.1 2.08 4.132 ;
  LAYER M1 ;
        RECT 2.112 4.08 2.144 6.588 ;
  LAYER M3 ;
        RECT 2.112 6.536 2.144 6.568 ;
  LAYER M1 ;
        RECT 2.176 4.08 2.208 6.588 ;
  LAYER M3 ;
        RECT 2.176 4.1 2.208 4.132 ;
  LAYER M1 ;
        RECT 2.24 4.08 2.272 6.588 ;
  LAYER M3 ;
        RECT 2.24 6.536 2.272 6.568 ;
  LAYER M1 ;
        RECT 2.304 4.08 2.336 6.588 ;
  LAYER M3 ;
        RECT 2.304 4.1 2.336 4.132 ;
  LAYER M1 ;
        RECT 2.368 4.08 2.4 6.588 ;
  LAYER M3 ;
        RECT 2.368 6.536 2.4 6.568 ;
  LAYER M1 ;
        RECT 2.432 4.08 2.464 6.588 ;
  LAYER M3 ;
        RECT 2.432 4.1 2.464 4.132 ;
  LAYER M1 ;
        RECT 2.496 4.08 2.528 6.588 ;
  LAYER M3 ;
        RECT 2.496 6.536 2.528 6.568 ;
  LAYER M1 ;
        RECT 2.56 4.08 2.592 6.588 ;
  LAYER M3 ;
        RECT 2.56 4.1 2.592 4.132 ;
  LAYER M1 ;
        RECT 2.624 4.08 2.656 6.588 ;
  LAYER M3 ;
        RECT 2.624 6.536 2.656 6.568 ;
  LAYER M1 ;
        RECT 2.688 4.08 2.72 6.588 ;
  LAYER M3 ;
        RECT 2.688 4.1 2.72 4.132 ;
  LAYER M1 ;
        RECT 2.752 4.08 2.784 6.588 ;
  LAYER M3 ;
        RECT 2.752 6.536 2.784 6.568 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 6.588 ;
  LAYER M3 ;
        RECT 0.448 4.164 0.48 4.196 ;
  LAYER M2 ;
        RECT 2.816 4.228 2.848 4.26 ;
  LAYER M2 ;
        RECT 0.448 4.292 0.48 4.324 ;
  LAYER M2 ;
        RECT 2.816 4.356 2.848 4.388 ;
  LAYER M2 ;
        RECT 0.448 4.42 0.48 4.452 ;
  LAYER M2 ;
        RECT 2.816 4.484 2.848 4.516 ;
  LAYER M2 ;
        RECT 0.448 4.548 0.48 4.58 ;
  LAYER M2 ;
        RECT 2.816 4.612 2.848 4.644 ;
  LAYER M2 ;
        RECT 0.448 4.676 0.48 4.708 ;
  LAYER M2 ;
        RECT 2.816 4.74 2.848 4.772 ;
  LAYER M2 ;
        RECT 0.448 4.804 0.48 4.836 ;
  LAYER M2 ;
        RECT 2.816 4.868 2.848 4.9 ;
  LAYER M2 ;
        RECT 0.448 4.932 0.48 4.964 ;
  LAYER M2 ;
        RECT 2.816 4.996 2.848 5.028 ;
  LAYER M2 ;
        RECT 0.448 5.06 0.48 5.092 ;
  LAYER M2 ;
        RECT 2.816 5.124 2.848 5.156 ;
  LAYER M2 ;
        RECT 0.448 5.188 0.48 5.22 ;
  LAYER M2 ;
        RECT 2.816 5.252 2.848 5.284 ;
  LAYER M2 ;
        RECT 0.448 5.316 0.48 5.348 ;
  LAYER M2 ;
        RECT 2.816 5.38 2.848 5.412 ;
  LAYER M2 ;
        RECT 0.448 5.444 0.48 5.476 ;
  LAYER M2 ;
        RECT 2.816 5.508 2.848 5.54 ;
  LAYER M2 ;
        RECT 0.448 5.572 0.48 5.604 ;
  LAYER M2 ;
        RECT 2.816 5.636 2.848 5.668 ;
  LAYER M2 ;
        RECT 0.448 5.7 0.48 5.732 ;
  LAYER M2 ;
        RECT 2.816 5.764 2.848 5.796 ;
  LAYER M2 ;
        RECT 0.448 5.828 0.48 5.86 ;
  LAYER M2 ;
        RECT 2.816 5.892 2.848 5.924 ;
  LAYER M2 ;
        RECT 0.448 5.956 0.48 5.988 ;
  LAYER M2 ;
        RECT 2.816 6.02 2.848 6.052 ;
  LAYER M2 ;
        RECT 0.448 6.084 0.48 6.116 ;
  LAYER M2 ;
        RECT 2.816 6.148 2.848 6.18 ;
  LAYER M2 ;
        RECT 0.448 6.212 0.48 6.244 ;
  LAYER M2 ;
        RECT 2.816 6.276 2.848 6.308 ;
  LAYER M2 ;
        RECT 0.448 6.34 0.48 6.372 ;
  LAYER M2 ;
        RECT 2.816 6.404 2.848 6.436 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.448 7.188 0.48 9.696 ;
  LAYER M3 ;
        RECT 0.448 9.644 0.48 9.676 ;
  LAYER M1 ;
        RECT 0.512 7.188 0.544 9.696 ;
  LAYER M3 ;
        RECT 0.512 7.208 0.544 7.24 ;
  LAYER M1 ;
        RECT 0.576 7.188 0.608 9.696 ;
  LAYER M3 ;
        RECT 0.576 9.644 0.608 9.676 ;
  LAYER M1 ;
        RECT 0.64 7.188 0.672 9.696 ;
  LAYER M3 ;
        RECT 0.64 7.208 0.672 7.24 ;
  LAYER M1 ;
        RECT 0.704 7.188 0.736 9.696 ;
  LAYER M3 ;
        RECT 0.704 9.644 0.736 9.676 ;
  LAYER M1 ;
        RECT 0.768 7.188 0.8 9.696 ;
  LAYER M3 ;
        RECT 0.768 7.208 0.8 7.24 ;
  LAYER M1 ;
        RECT 0.832 7.188 0.864 9.696 ;
  LAYER M3 ;
        RECT 0.832 9.644 0.864 9.676 ;
  LAYER M1 ;
        RECT 0.896 7.188 0.928 9.696 ;
  LAYER M3 ;
        RECT 0.896 7.208 0.928 7.24 ;
  LAYER M1 ;
        RECT 0.96 7.188 0.992 9.696 ;
  LAYER M3 ;
        RECT 0.96 9.644 0.992 9.676 ;
  LAYER M1 ;
        RECT 1.024 7.188 1.056 9.696 ;
  LAYER M3 ;
        RECT 1.024 7.208 1.056 7.24 ;
  LAYER M1 ;
        RECT 1.088 7.188 1.12 9.696 ;
  LAYER M3 ;
        RECT 1.088 9.644 1.12 9.676 ;
  LAYER M1 ;
        RECT 1.152 7.188 1.184 9.696 ;
  LAYER M3 ;
        RECT 1.152 7.208 1.184 7.24 ;
  LAYER M1 ;
        RECT 1.216 7.188 1.248 9.696 ;
  LAYER M3 ;
        RECT 1.216 9.644 1.248 9.676 ;
  LAYER M1 ;
        RECT 1.28 7.188 1.312 9.696 ;
  LAYER M3 ;
        RECT 1.28 7.208 1.312 7.24 ;
  LAYER M1 ;
        RECT 1.344 7.188 1.376 9.696 ;
  LAYER M3 ;
        RECT 1.344 9.644 1.376 9.676 ;
  LAYER M1 ;
        RECT 1.408 7.188 1.44 9.696 ;
  LAYER M3 ;
        RECT 1.408 7.208 1.44 7.24 ;
  LAYER M1 ;
        RECT 1.472 7.188 1.504 9.696 ;
  LAYER M3 ;
        RECT 1.472 9.644 1.504 9.676 ;
  LAYER M1 ;
        RECT 1.536 7.188 1.568 9.696 ;
  LAYER M3 ;
        RECT 1.536 7.208 1.568 7.24 ;
  LAYER M1 ;
        RECT 1.6 7.188 1.632 9.696 ;
  LAYER M3 ;
        RECT 1.6 9.644 1.632 9.676 ;
  LAYER M1 ;
        RECT 1.664 7.188 1.696 9.696 ;
  LAYER M3 ;
        RECT 1.664 7.208 1.696 7.24 ;
  LAYER M1 ;
        RECT 1.728 7.188 1.76 9.696 ;
  LAYER M3 ;
        RECT 1.728 9.644 1.76 9.676 ;
  LAYER M1 ;
        RECT 1.792 7.188 1.824 9.696 ;
  LAYER M3 ;
        RECT 1.792 7.208 1.824 7.24 ;
  LAYER M1 ;
        RECT 1.856 7.188 1.888 9.696 ;
  LAYER M3 ;
        RECT 1.856 9.644 1.888 9.676 ;
  LAYER M1 ;
        RECT 1.92 7.188 1.952 9.696 ;
  LAYER M3 ;
        RECT 1.92 7.208 1.952 7.24 ;
  LAYER M1 ;
        RECT 1.984 7.188 2.016 9.696 ;
  LAYER M3 ;
        RECT 1.984 9.644 2.016 9.676 ;
  LAYER M1 ;
        RECT 2.048 7.188 2.08 9.696 ;
  LAYER M3 ;
        RECT 2.048 7.208 2.08 7.24 ;
  LAYER M1 ;
        RECT 2.112 7.188 2.144 9.696 ;
  LAYER M3 ;
        RECT 2.112 9.644 2.144 9.676 ;
  LAYER M1 ;
        RECT 2.176 7.188 2.208 9.696 ;
  LAYER M3 ;
        RECT 2.176 7.208 2.208 7.24 ;
  LAYER M1 ;
        RECT 2.24 7.188 2.272 9.696 ;
  LAYER M3 ;
        RECT 2.24 9.644 2.272 9.676 ;
  LAYER M1 ;
        RECT 2.304 7.188 2.336 9.696 ;
  LAYER M3 ;
        RECT 2.304 7.208 2.336 7.24 ;
  LAYER M1 ;
        RECT 2.368 7.188 2.4 9.696 ;
  LAYER M3 ;
        RECT 2.368 9.644 2.4 9.676 ;
  LAYER M1 ;
        RECT 2.432 7.188 2.464 9.696 ;
  LAYER M3 ;
        RECT 2.432 7.208 2.464 7.24 ;
  LAYER M1 ;
        RECT 2.496 7.188 2.528 9.696 ;
  LAYER M3 ;
        RECT 2.496 9.644 2.528 9.676 ;
  LAYER M1 ;
        RECT 2.56 7.188 2.592 9.696 ;
  LAYER M3 ;
        RECT 2.56 7.208 2.592 7.24 ;
  LAYER M1 ;
        RECT 2.624 7.188 2.656 9.696 ;
  LAYER M3 ;
        RECT 2.624 9.644 2.656 9.676 ;
  LAYER M1 ;
        RECT 2.688 7.188 2.72 9.696 ;
  LAYER M3 ;
        RECT 2.688 7.208 2.72 7.24 ;
  LAYER M1 ;
        RECT 2.752 7.188 2.784 9.696 ;
  LAYER M3 ;
        RECT 2.752 9.644 2.784 9.676 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 9.696 ;
  LAYER M3 ;
        RECT 0.448 7.272 0.48 7.304 ;
  LAYER M2 ;
        RECT 2.816 7.336 2.848 7.368 ;
  LAYER M2 ;
        RECT 0.448 7.4 0.48 7.432 ;
  LAYER M2 ;
        RECT 2.816 7.464 2.848 7.496 ;
  LAYER M2 ;
        RECT 0.448 7.528 0.48 7.56 ;
  LAYER M2 ;
        RECT 2.816 7.592 2.848 7.624 ;
  LAYER M2 ;
        RECT 0.448 7.656 0.48 7.688 ;
  LAYER M2 ;
        RECT 2.816 7.72 2.848 7.752 ;
  LAYER M2 ;
        RECT 0.448 7.784 0.48 7.816 ;
  LAYER M2 ;
        RECT 2.816 7.848 2.848 7.88 ;
  LAYER M2 ;
        RECT 0.448 7.912 0.48 7.944 ;
  LAYER M2 ;
        RECT 2.816 7.976 2.848 8.008 ;
  LAYER M2 ;
        RECT 0.448 8.04 0.48 8.072 ;
  LAYER M2 ;
        RECT 2.816 8.104 2.848 8.136 ;
  LAYER M2 ;
        RECT 0.448 8.168 0.48 8.2 ;
  LAYER M2 ;
        RECT 2.816 8.232 2.848 8.264 ;
  LAYER M2 ;
        RECT 0.448 8.296 0.48 8.328 ;
  LAYER M2 ;
        RECT 2.816 8.36 2.848 8.392 ;
  LAYER M2 ;
        RECT 0.448 8.424 0.48 8.456 ;
  LAYER M2 ;
        RECT 2.816 8.488 2.848 8.52 ;
  LAYER M2 ;
        RECT 0.448 8.552 0.48 8.584 ;
  LAYER M2 ;
        RECT 2.816 8.616 2.848 8.648 ;
  LAYER M2 ;
        RECT 0.448 8.68 0.48 8.712 ;
  LAYER M2 ;
        RECT 2.816 8.744 2.848 8.776 ;
  LAYER M2 ;
        RECT 0.448 8.808 0.48 8.84 ;
  LAYER M2 ;
        RECT 2.816 8.872 2.848 8.904 ;
  LAYER M2 ;
        RECT 0.448 8.936 0.48 8.968 ;
  LAYER M2 ;
        RECT 2.816 9 2.848 9.032 ;
  LAYER M2 ;
        RECT 0.448 9.064 0.48 9.096 ;
  LAYER M2 ;
        RECT 2.816 9.128 2.848 9.16 ;
  LAYER M2 ;
        RECT 0.448 9.192 0.48 9.224 ;
  LAYER M2 ;
        RECT 2.816 9.256 2.848 9.288 ;
  LAYER M2 ;
        RECT 0.448 9.32 0.48 9.352 ;
  LAYER M2 ;
        RECT 2.816 9.384 2.848 9.416 ;
  LAYER M2 ;
        RECT 0.448 9.448 0.48 9.48 ;
  LAYER M2 ;
        RECT 2.816 9.512 2.848 9.544 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.448 10.296 0.48 12.804 ;
  LAYER M3 ;
        RECT 0.448 12.752 0.48 12.784 ;
  LAYER M1 ;
        RECT 0.512 10.296 0.544 12.804 ;
  LAYER M3 ;
        RECT 0.512 10.316 0.544 10.348 ;
  LAYER M1 ;
        RECT 0.576 10.296 0.608 12.804 ;
  LAYER M3 ;
        RECT 0.576 12.752 0.608 12.784 ;
  LAYER M1 ;
        RECT 0.64 10.296 0.672 12.804 ;
  LAYER M3 ;
        RECT 0.64 10.316 0.672 10.348 ;
  LAYER M1 ;
        RECT 0.704 10.296 0.736 12.804 ;
  LAYER M3 ;
        RECT 0.704 12.752 0.736 12.784 ;
  LAYER M1 ;
        RECT 0.768 10.296 0.8 12.804 ;
  LAYER M3 ;
        RECT 0.768 10.316 0.8 10.348 ;
  LAYER M1 ;
        RECT 0.832 10.296 0.864 12.804 ;
  LAYER M3 ;
        RECT 0.832 12.752 0.864 12.784 ;
  LAYER M1 ;
        RECT 0.896 10.296 0.928 12.804 ;
  LAYER M3 ;
        RECT 0.896 10.316 0.928 10.348 ;
  LAYER M1 ;
        RECT 0.96 10.296 0.992 12.804 ;
  LAYER M3 ;
        RECT 0.96 12.752 0.992 12.784 ;
  LAYER M1 ;
        RECT 1.024 10.296 1.056 12.804 ;
  LAYER M3 ;
        RECT 1.024 10.316 1.056 10.348 ;
  LAYER M1 ;
        RECT 1.088 10.296 1.12 12.804 ;
  LAYER M3 ;
        RECT 1.088 12.752 1.12 12.784 ;
  LAYER M1 ;
        RECT 1.152 10.296 1.184 12.804 ;
  LAYER M3 ;
        RECT 1.152 10.316 1.184 10.348 ;
  LAYER M1 ;
        RECT 1.216 10.296 1.248 12.804 ;
  LAYER M3 ;
        RECT 1.216 12.752 1.248 12.784 ;
  LAYER M1 ;
        RECT 1.28 10.296 1.312 12.804 ;
  LAYER M3 ;
        RECT 1.28 10.316 1.312 10.348 ;
  LAYER M1 ;
        RECT 1.344 10.296 1.376 12.804 ;
  LAYER M3 ;
        RECT 1.344 12.752 1.376 12.784 ;
  LAYER M1 ;
        RECT 1.408 10.296 1.44 12.804 ;
  LAYER M3 ;
        RECT 1.408 10.316 1.44 10.348 ;
  LAYER M1 ;
        RECT 1.472 10.296 1.504 12.804 ;
  LAYER M3 ;
        RECT 1.472 12.752 1.504 12.784 ;
  LAYER M1 ;
        RECT 1.536 10.296 1.568 12.804 ;
  LAYER M3 ;
        RECT 1.536 10.316 1.568 10.348 ;
  LAYER M1 ;
        RECT 1.6 10.296 1.632 12.804 ;
  LAYER M3 ;
        RECT 1.6 12.752 1.632 12.784 ;
  LAYER M1 ;
        RECT 1.664 10.296 1.696 12.804 ;
  LAYER M3 ;
        RECT 1.664 10.316 1.696 10.348 ;
  LAYER M1 ;
        RECT 1.728 10.296 1.76 12.804 ;
  LAYER M3 ;
        RECT 1.728 12.752 1.76 12.784 ;
  LAYER M1 ;
        RECT 1.792 10.296 1.824 12.804 ;
  LAYER M3 ;
        RECT 1.792 10.316 1.824 10.348 ;
  LAYER M1 ;
        RECT 1.856 10.296 1.888 12.804 ;
  LAYER M3 ;
        RECT 1.856 12.752 1.888 12.784 ;
  LAYER M1 ;
        RECT 1.92 10.296 1.952 12.804 ;
  LAYER M3 ;
        RECT 1.92 10.316 1.952 10.348 ;
  LAYER M1 ;
        RECT 1.984 10.296 2.016 12.804 ;
  LAYER M3 ;
        RECT 1.984 12.752 2.016 12.784 ;
  LAYER M1 ;
        RECT 2.048 10.296 2.08 12.804 ;
  LAYER M3 ;
        RECT 2.048 10.316 2.08 10.348 ;
  LAYER M1 ;
        RECT 2.112 10.296 2.144 12.804 ;
  LAYER M3 ;
        RECT 2.112 12.752 2.144 12.784 ;
  LAYER M1 ;
        RECT 2.176 10.296 2.208 12.804 ;
  LAYER M3 ;
        RECT 2.176 10.316 2.208 10.348 ;
  LAYER M1 ;
        RECT 2.24 10.296 2.272 12.804 ;
  LAYER M3 ;
        RECT 2.24 12.752 2.272 12.784 ;
  LAYER M1 ;
        RECT 2.304 10.296 2.336 12.804 ;
  LAYER M3 ;
        RECT 2.304 10.316 2.336 10.348 ;
  LAYER M1 ;
        RECT 2.368 10.296 2.4 12.804 ;
  LAYER M3 ;
        RECT 2.368 12.752 2.4 12.784 ;
  LAYER M1 ;
        RECT 2.432 10.296 2.464 12.804 ;
  LAYER M3 ;
        RECT 2.432 10.316 2.464 10.348 ;
  LAYER M1 ;
        RECT 2.496 10.296 2.528 12.804 ;
  LAYER M3 ;
        RECT 2.496 12.752 2.528 12.784 ;
  LAYER M1 ;
        RECT 2.56 10.296 2.592 12.804 ;
  LAYER M3 ;
        RECT 2.56 10.316 2.592 10.348 ;
  LAYER M1 ;
        RECT 2.624 10.296 2.656 12.804 ;
  LAYER M3 ;
        RECT 2.624 12.752 2.656 12.784 ;
  LAYER M1 ;
        RECT 2.688 10.296 2.72 12.804 ;
  LAYER M3 ;
        RECT 2.688 10.316 2.72 10.348 ;
  LAYER M1 ;
        RECT 2.752 10.296 2.784 12.804 ;
  LAYER M3 ;
        RECT 2.752 12.752 2.784 12.784 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 12.804 ;
  LAYER M3 ;
        RECT 0.448 10.38 0.48 10.412 ;
  LAYER M2 ;
        RECT 2.816 10.444 2.848 10.476 ;
  LAYER M2 ;
        RECT 0.448 10.508 0.48 10.54 ;
  LAYER M2 ;
        RECT 2.816 10.572 2.848 10.604 ;
  LAYER M2 ;
        RECT 0.448 10.636 0.48 10.668 ;
  LAYER M2 ;
        RECT 2.816 10.7 2.848 10.732 ;
  LAYER M2 ;
        RECT 0.448 10.764 0.48 10.796 ;
  LAYER M2 ;
        RECT 2.816 10.828 2.848 10.86 ;
  LAYER M2 ;
        RECT 0.448 10.892 0.48 10.924 ;
  LAYER M2 ;
        RECT 2.816 10.956 2.848 10.988 ;
  LAYER M2 ;
        RECT 0.448 11.02 0.48 11.052 ;
  LAYER M2 ;
        RECT 2.816 11.084 2.848 11.116 ;
  LAYER M2 ;
        RECT 0.448 11.148 0.48 11.18 ;
  LAYER M2 ;
        RECT 2.816 11.212 2.848 11.244 ;
  LAYER M2 ;
        RECT 0.448 11.276 0.48 11.308 ;
  LAYER M2 ;
        RECT 2.816 11.34 2.848 11.372 ;
  LAYER M2 ;
        RECT 0.448 11.404 0.48 11.436 ;
  LAYER M2 ;
        RECT 2.816 11.468 2.848 11.5 ;
  LAYER M2 ;
        RECT 0.448 11.532 0.48 11.564 ;
  LAYER M2 ;
        RECT 2.816 11.596 2.848 11.628 ;
  LAYER M2 ;
        RECT 0.448 11.66 0.48 11.692 ;
  LAYER M2 ;
        RECT 2.816 11.724 2.848 11.756 ;
  LAYER M2 ;
        RECT 0.448 11.788 0.48 11.82 ;
  LAYER M2 ;
        RECT 2.816 11.852 2.848 11.884 ;
  LAYER M2 ;
        RECT 0.448 11.916 0.48 11.948 ;
  LAYER M2 ;
        RECT 2.816 11.98 2.848 12.012 ;
  LAYER M2 ;
        RECT 0.448 12.044 0.48 12.076 ;
  LAYER M2 ;
        RECT 2.816 12.108 2.848 12.14 ;
  LAYER M2 ;
        RECT 0.448 12.172 0.48 12.204 ;
  LAYER M2 ;
        RECT 2.816 12.236 2.848 12.268 ;
  LAYER M2 ;
        RECT 0.448 12.3 0.48 12.332 ;
  LAYER M2 ;
        RECT 2.816 12.364 2.848 12.396 ;
  LAYER M2 ;
        RECT 0.448 12.428 0.48 12.46 ;
  LAYER M2 ;
        RECT 2.816 12.492 2.848 12.524 ;
  LAYER M2 ;
        RECT 0.448 12.556 0.48 12.588 ;
  LAYER M2 ;
        RECT 2.816 12.62 2.848 12.652 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 0.448 13.404 0.48 15.912 ;
  LAYER M3 ;
        RECT 0.448 15.86 0.48 15.892 ;
  LAYER M1 ;
        RECT 0.512 13.404 0.544 15.912 ;
  LAYER M3 ;
        RECT 0.512 13.424 0.544 13.456 ;
  LAYER M1 ;
        RECT 0.576 13.404 0.608 15.912 ;
  LAYER M3 ;
        RECT 0.576 15.86 0.608 15.892 ;
  LAYER M1 ;
        RECT 0.64 13.404 0.672 15.912 ;
  LAYER M3 ;
        RECT 0.64 13.424 0.672 13.456 ;
  LAYER M1 ;
        RECT 0.704 13.404 0.736 15.912 ;
  LAYER M3 ;
        RECT 0.704 15.86 0.736 15.892 ;
  LAYER M1 ;
        RECT 0.768 13.404 0.8 15.912 ;
  LAYER M3 ;
        RECT 0.768 13.424 0.8 13.456 ;
  LAYER M1 ;
        RECT 0.832 13.404 0.864 15.912 ;
  LAYER M3 ;
        RECT 0.832 15.86 0.864 15.892 ;
  LAYER M1 ;
        RECT 0.896 13.404 0.928 15.912 ;
  LAYER M3 ;
        RECT 0.896 13.424 0.928 13.456 ;
  LAYER M1 ;
        RECT 0.96 13.404 0.992 15.912 ;
  LAYER M3 ;
        RECT 0.96 15.86 0.992 15.892 ;
  LAYER M1 ;
        RECT 1.024 13.404 1.056 15.912 ;
  LAYER M3 ;
        RECT 1.024 13.424 1.056 13.456 ;
  LAYER M1 ;
        RECT 1.088 13.404 1.12 15.912 ;
  LAYER M3 ;
        RECT 1.088 15.86 1.12 15.892 ;
  LAYER M1 ;
        RECT 1.152 13.404 1.184 15.912 ;
  LAYER M3 ;
        RECT 1.152 13.424 1.184 13.456 ;
  LAYER M1 ;
        RECT 1.216 13.404 1.248 15.912 ;
  LAYER M3 ;
        RECT 1.216 15.86 1.248 15.892 ;
  LAYER M1 ;
        RECT 1.28 13.404 1.312 15.912 ;
  LAYER M3 ;
        RECT 1.28 13.424 1.312 13.456 ;
  LAYER M1 ;
        RECT 1.344 13.404 1.376 15.912 ;
  LAYER M3 ;
        RECT 1.344 15.86 1.376 15.892 ;
  LAYER M1 ;
        RECT 1.408 13.404 1.44 15.912 ;
  LAYER M3 ;
        RECT 1.408 13.424 1.44 13.456 ;
  LAYER M1 ;
        RECT 1.472 13.404 1.504 15.912 ;
  LAYER M3 ;
        RECT 1.472 15.86 1.504 15.892 ;
  LAYER M1 ;
        RECT 1.536 13.404 1.568 15.912 ;
  LAYER M3 ;
        RECT 1.536 13.424 1.568 13.456 ;
  LAYER M1 ;
        RECT 1.6 13.404 1.632 15.912 ;
  LAYER M3 ;
        RECT 1.6 15.86 1.632 15.892 ;
  LAYER M1 ;
        RECT 1.664 13.404 1.696 15.912 ;
  LAYER M3 ;
        RECT 1.664 13.424 1.696 13.456 ;
  LAYER M1 ;
        RECT 1.728 13.404 1.76 15.912 ;
  LAYER M3 ;
        RECT 1.728 15.86 1.76 15.892 ;
  LAYER M1 ;
        RECT 1.792 13.404 1.824 15.912 ;
  LAYER M3 ;
        RECT 1.792 13.424 1.824 13.456 ;
  LAYER M1 ;
        RECT 1.856 13.404 1.888 15.912 ;
  LAYER M3 ;
        RECT 1.856 15.86 1.888 15.892 ;
  LAYER M1 ;
        RECT 1.92 13.404 1.952 15.912 ;
  LAYER M3 ;
        RECT 1.92 13.424 1.952 13.456 ;
  LAYER M1 ;
        RECT 1.984 13.404 2.016 15.912 ;
  LAYER M3 ;
        RECT 1.984 15.86 2.016 15.892 ;
  LAYER M1 ;
        RECT 2.048 13.404 2.08 15.912 ;
  LAYER M3 ;
        RECT 2.048 13.424 2.08 13.456 ;
  LAYER M1 ;
        RECT 2.112 13.404 2.144 15.912 ;
  LAYER M3 ;
        RECT 2.112 15.86 2.144 15.892 ;
  LAYER M1 ;
        RECT 2.176 13.404 2.208 15.912 ;
  LAYER M3 ;
        RECT 2.176 13.424 2.208 13.456 ;
  LAYER M1 ;
        RECT 2.24 13.404 2.272 15.912 ;
  LAYER M3 ;
        RECT 2.24 15.86 2.272 15.892 ;
  LAYER M1 ;
        RECT 2.304 13.404 2.336 15.912 ;
  LAYER M3 ;
        RECT 2.304 13.424 2.336 13.456 ;
  LAYER M1 ;
        RECT 2.368 13.404 2.4 15.912 ;
  LAYER M3 ;
        RECT 2.368 15.86 2.4 15.892 ;
  LAYER M1 ;
        RECT 2.432 13.404 2.464 15.912 ;
  LAYER M3 ;
        RECT 2.432 13.424 2.464 13.456 ;
  LAYER M1 ;
        RECT 2.496 13.404 2.528 15.912 ;
  LAYER M3 ;
        RECT 2.496 15.86 2.528 15.892 ;
  LAYER M1 ;
        RECT 2.56 13.404 2.592 15.912 ;
  LAYER M3 ;
        RECT 2.56 13.424 2.592 13.456 ;
  LAYER M1 ;
        RECT 2.624 13.404 2.656 15.912 ;
  LAYER M3 ;
        RECT 2.624 15.86 2.656 15.892 ;
  LAYER M1 ;
        RECT 2.688 13.404 2.72 15.912 ;
  LAYER M3 ;
        RECT 2.688 13.424 2.72 13.456 ;
  LAYER M1 ;
        RECT 2.752 13.404 2.784 15.912 ;
  LAYER M3 ;
        RECT 2.752 15.86 2.784 15.892 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 15.912 ;
  LAYER M3 ;
        RECT 0.448 13.488 0.48 13.52 ;
  LAYER M2 ;
        RECT 2.816 13.552 2.848 13.584 ;
  LAYER M2 ;
        RECT 0.448 13.616 0.48 13.648 ;
  LAYER M2 ;
        RECT 2.816 13.68 2.848 13.712 ;
  LAYER M2 ;
        RECT 0.448 13.744 0.48 13.776 ;
  LAYER M2 ;
        RECT 2.816 13.808 2.848 13.84 ;
  LAYER M2 ;
        RECT 0.448 13.872 0.48 13.904 ;
  LAYER M2 ;
        RECT 2.816 13.936 2.848 13.968 ;
  LAYER M2 ;
        RECT 0.448 14 0.48 14.032 ;
  LAYER M2 ;
        RECT 2.816 14.064 2.848 14.096 ;
  LAYER M2 ;
        RECT 0.448 14.128 0.48 14.16 ;
  LAYER M2 ;
        RECT 2.816 14.192 2.848 14.224 ;
  LAYER M2 ;
        RECT 0.448 14.256 0.48 14.288 ;
  LAYER M2 ;
        RECT 2.816 14.32 2.848 14.352 ;
  LAYER M2 ;
        RECT 0.448 14.384 0.48 14.416 ;
  LAYER M2 ;
        RECT 2.816 14.448 2.848 14.48 ;
  LAYER M2 ;
        RECT 0.448 14.512 0.48 14.544 ;
  LAYER M2 ;
        RECT 2.816 14.576 2.848 14.608 ;
  LAYER M2 ;
        RECT 0.448 14.64 0.48 14.672 ;
  LAYER M2 ;
        RECT 2.816 14.704 2.848 14.736 ;
  LAYER M2 ;
        RECT 0.448 14.768 0.48 14.8 ;
  LAYER M2 ;
        RECT 2.816 14.832 2.848 14.864 ;
  LAYER M2 ;
        RECT 0.448 14.896 0.48 14.928 ;
  LAYER M2 ;
        RECT 2.816 14.96 2.848 14.992 ;
  LAYER M2 ;
        RECT 0.448 15.024 0.48 15.056 ;
  LAYER M2 ;
        RECT 2.816 15.088 2.848 15.12 ;
  LAYER M2 ;
        RECT 0.448 15.152 0.48 15.184 ;
  LAYER M2 ;
        RECT 2.816 15.216 2.848 15.248 ;
  LAYER M2 ;
        RECT 0.448 15.28 0.48 15.312 ;
  LAYER M2 ;
        RECT 2.816 15.344 2.848 15.376 ;
  LAYER M2 ;
        RECT 0.448 15.408 0.48 15.44 ;
  LAYER M2 ;
        RECT 2.816 15.472 2.848 15.504 ;
  LAYER M2 ;
        RECT 0.448 15.536 0.48 15.568 ;
  LAYER M2 ;
        RECT 2.816 15.6 2.848 15.632 ;
  LAYER M2 ;
        RECT 0.448 15.664 0.48 15.696 ;
  LAYER M2 ;
        RECT 2.816 15.728 2.848 15.76 ;
  LAYER M2 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M1 ;
        RECT 3.424 0.972 3.456 3.48 ;
  LAYER M3 ;
        RECT 3.424 3.428 3.456 3.46 ;
  LAYER M1 ;
        RECT 3.488 0.972 3.52 3.48 ;
  LAYER M3 ;
        RECT 3.488 0.992 3.52 1.024 ;
  LAYER M1 ;
        RECT 3.552 0.972 3.584 3.48 ;
  LAYER M3 ;
        RECT 3.552 3.428 3.584 3.46 ;
  LAYER M1 ;
        RECT 3.616 0.972 3.648 3.48 ;
  LAYER M3 ;
        RECT 3.616 0.992 3.648 1.024 ;
  LAYER M1 ;
        RECT 3.68 0.972 3.712 3.48 ;
  LAYER M3 ;
        RECT 3.68 3.428 3.712 3.46 ;
  LAYER M1 ;
        RECT 3.744 0.972 3.776 3.48 ;
  LAYER M3 ;
        RECT 3.744 0.992 3.776 1.024 ;
  LAYER M1 ;
        RECT 3.808 0.972 3.84 3.48 ;
  LAYER M3 ;
        RECT 3.808 3.428 3.84 3.46 ;
  LAYER M1 ;
        RECT 3.872 0.972 3.904 3.48 ;
  LAYER M3 ;
        RECT 3.872 0.992 3.904 1.024 ;
  LAYER M1 ;
        RECT 3.936 0.972 3.968 3.48 ;
  LAYER M3 ;
        RECT 3.936 3.428 3.968 3.46 ;
  LAYER M1 ;
        RECT 4 0.972 4.032 3.48 ;
  LAYER M3 ;
        RECT 4 0.992 4.032 1.024 ;
  LAYER M1 ;
        RECT 4.064 0.972 4.096 3.48 ;
  LAYER M3 ;
        RECT 4.064 3.428 4.096 3.46 ;
  LAYER M1 ;
        RECT 4.128 0.972 4.16 3.48 ;
  LAYER M3 ;
        RECT 4.128 0.992 4.16 1.024 ;
  LAYER M1 ;
        RECT 4.192 0.972 4.224 3.48 ;
  LAYER M3 ;
        RECT 4.192 3.428 4.224 3.46 ;
  LAYER M1 ;
        RECT 4.256 0.972 4.288 3.48 ;
  LAYER M3 ;
        RECT 4.256 0.992 4.288 1.024 ;
  LAYER M1 ;
        RECT 4.32 0.972 4.352 3.48 ;
  LAYER M3 ;
        RECT 4.32 3.428 4.352 3.46 ;
  LAYER M1 ;
        RECT 4.384 0.972 4.416 3.48 ;
  LAYER M3 ;
        RECT 4.384 0.992 4.416 1.024 ;
  LAYER M1 ;
        RECT 4.448 0.972 4.48 3.48 ;
  LAYER M3 ;
        RECT 4.448 3.428 4.48 3.46 ;
  LAYER M1 ;
        RECT 4.512 0.972 4.544 3.48 ;
  LAYER M3 ;
        RECT 4.512 0.992 4.544 1.024 ;
  LAYER M1 ;
        RECT 4.576 0.972 4.608 3.48 ;
  LAYER M3 ;
        RECT 4.576 3.428 4.608 3.46 ;
  LAYER M1 ;
        RECT 4.64 0.972 4.672 3.48 ;
  LAYER M3 ;
        RECT 4.64 0.992 4.672 1.024 ;
  LAYER M1 ;
        RECT 4.704 0.972 4.736 3.48 ;
  LAYER M3 ;
        RECT 4.704 3.428 4.736 3.46 ;
  LAYER M1 ;
        RECT 4.768 0.972 4.8 3.48 ;
  LAYER M3 ;
        RECT 4.768 0.992 4.8 1.024 ;
  LAYER M1 ;
        RECT 4.832 0.972 4.864 3.48 ;
  LAYER M3 ;
        RECT 4.832 3.428 4.864 3.46 ;
  LAYER M1 ;
        RECT 4.896 0.972 4.928 3.48 ;
  LAYER M3 ;
        RECT 4.896 0.992 4.928 1.024 ;
  LAYER M1 ;
        RECT 4.96 0.972 4.992 3.48 ;
  LAYER M3 ;
        RECT 4.96 3.428 4.992 3.46 ;
  LAYER M1 ;
        RECT 5.024 0.972 5.056 3.48 ;
  LAYER M3 ;
        RECT 5.024 0.992 5.056 1.024 ;
  LAYER M1 ;
        RECT 5.088 0.972 5.12 3.48 ;
  LAYER M3 ;
        RECT 5.088 3.428 5.12 3.46 ;
  LAYER M1 ;
        RECT 5.152 0.972 5.184 3.48 ;
  LAYER M3 ;
        RECT 5.152 0.992 5.184 1.024 ;
  LAYER M1 ;
        RECT 5.216 0.972 5.248 3.48 ;
  LAYER M3 ;
        RECT 5.216 3.428 5.248 3.46 ;
  LAYER M1 ;
        RECT 5.28 0.972 5.312 3.48 ;
  LAYER M3 ;
        RECT 5.28 0.992 5.312 1.024 ;
  LAYER M1 ;
        RECT 5.344 0.972 5.376 3.48 ;
  LAYER M3 ;
        RECT 5.344 3.428 5.376 3.46 ;
  LAYER M1 ;
        RECT 5.408 0.972 5.44 3.48 ;
  LAYER M3 ;
        RECT 5.408 0.992 5.44 1.024 ;
  LAYER M1 ;
        RECT 5.472 0.972 5.504 3.48 ;
  LAYER M3 ;
        RECT 5.472 3.428 5.504 3.46 ;
  LAYER M1 ;
        RECT 5.536 0.972 5.568 3.48 ;
  LAYER M3 ;
        RECT 5.536 0.992 5.568 1.024 ;
  LAYER M1 ;
        RECT 5.6 0.972 5.632 3.48 ;
  LAYER M3 ;
        RECT 5.6 3.428 5.632 3.46 ;
  LAYER M1 ;
        RECT 5.664 0.972 5.696 3.48 ;
  LAYER M3 ;
        RECT 5.664 0.992 5.696 1.024 ;
  LAYER M1 ;
        RECT 5.728 0.972 5.76 3.48 ;
  LAYER M3 ;
        RECT 5.728 3.428 5.76 3.46 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 3.48 ;
  LAYER M3 ;
        RECT 3.424 1.056 3.456 1.088 ;
  LAYER M2 ;
        RECT 5.792 1.12 5.824 1.152 ;
  LAYER M2 ;
        RECT 3.424 1.184 3.456 1.216 ;
  LAYER M2 ;
        RECT 5.792 1.248 5.824 1.28 ;
  LAYER M2 ;
        RECT 3.424 1.312 3.456 1.344 ;
  LAYER M2 ;
        RECT 5.792 1.376 5.824 1.408 ;
  LAYER M2 ;
        RECT 3.424 1.44 3.456 1.472 ;
  LAYER M2 ;
        RECT 5.792 1.504 5.824 1.536 ;
  LAYER M2 ;
        RECT 3.424 1.568 3.456 1.6 ;
  LAYER M2 ;
        RECT 5.792 1.632 5.824 1.664 ;
  LAYER M2 ;
        RECT 3.424 1.696 3.456 1.728 ;
  LAYER M2 ;
        RECT 5.792 1.76 5.824 1.792 ;
  LAYER M2 ;
        RECT 3.424 1.824 3.456 1.856 ;
  LAYER M2 ;
        RECT 5.792 1.888 5.824 1.92 ;
  LAYER M2 ;
        RECT 3.424 1.952 3.456 1.984 ;
  LAYER M2 ;
        RECT 5.792 2.016 5.824 2.048 ;
  LAYER M2 ;
        RECT 3.424 2.08 3.456 2.112 ;
  LAYER M2 ;
        RECT 5.792 2.144 5.824 2.176 ;
  LAYER M2 ;
        RECT 3.424 2.208 3.456 2.24 ;
  LAYER M2 ;
        RECT 5.792 2.272 5.824 2.304 ;
  LAYER M2 ;
        RECT 3.424 2.336 3.456 2.368 ;
  LAYER M2 ;
        RECT 5.792 2.4 5.824 2.432 ;
  LAYER M2 ;
        RECT 3.424 2.464 3.456 2.496 ;
  LAYER M2 ;
        RECT 5.792 2.528 5.824 2.56 ;
  LAYER M2 ;
        RECT 3.424 2.592 3.456 2.624 ;
  LAYER M2 ;
        RECT 5.792 2.656 5.824 2.688 ;
  LAYER M2 ;
        RECT 3.424 2.72 3.456 2.752 ;
  LAYER M2 ;
        RECT 5.792 2.784 5.824 2.816 ;
  LAYER M2 ;
        RECT 3.424 2.848 3.456 2.88 ;
  LAYER M2 ;
        RECT 5.792 2.912 5.824 2.944 ;
  LAYER M2 ;
        RECT 3.424 2.976 3.456 3.008 ;
  LAYER M2 ;
        RECT 5.792 3.04 5.824 3.072 ;
  LAYER M2 ;
        RECT 3.424 3.104 3.456 3.136 ;
  LAYER M2 ;
        RECT 5.792 3.168 5.824 3.2 ;
  LAYER M2 ;
        RECT 3.424 3.232 3.456 3.264 ;
  LAYER M2 ;
        RECT 5.792 3.296 5.824 3.328 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.424 4.08 3.456 6.588 ;
  LAYER M3 ;
        RECT 3.424 6.536 3.456 6.568 ;
  LAYER M1 ;
        RECT 3.488 4.08 3.52 6.588 ;
  LAYER M3 ;
        RECT 3.488 4.1 3.52 4.132 ;
  LAYER M1 ;
        RECT 3.552 4.08 3.584 6.588 ;
  LAYER M3 ;
        RECT 3.552 6.536 3.584 6.568 ;
  LAYER M1 ;
        RECT 3.616 4.08 3.648 6.588 ;
  LAYER M3 ;
        RECT 3.616 4.1 3.648 4.132 ;
  LAYER M1 ;
        RECT 3.68 4.08 3.712 6.588 ;
  LAYER M3 ;
        RECT 3.68 6.536 3.712 6.568 ;
  LAYER M1 ;
        RECT 3.744 4.08 3.776 6.588 ;
  LAYER M3 ;
        RECT 3.744 4.1 3.776 4.132 ;
  LAYER M1 ;
        RECT 3.808 4.08 3.84 6.588 ;
  LAYER M3 ;
        RECT 3.808 6.536 3.84 6.568 ;
  LAYER M1 ;
        RECT 3.872 4.08 3.904 6.588 ;
  LAYER M3 ;
        RECT 3.872 4.1 3.904 4.132 ;
  LAYER M1 ;
        RECT 3.936 4.08 3.968 6.588 ;
  LAYER M3 ;
        RECT 3.936 6.536 3.968 6.568 ;
  LAYER M1 ;
        RECT 4 4.08 4.032 6.588 ;
  LAYER M3 ;
        RECT 4 4.1 4.032 4.132 ;
  LAYER M1 ;
        RECT 4.064 4.08 4.096 6.588 ;
  LAYER M3 ;
        RECT 4.064 6.536 4.096 6.568 ;
  LAYER M1 ;
        RECT 4.128 4.08 4.16 6.588 ;
  LAYER M3 ;
        RECT 4.128 4.1 4.16 4.132 ;
  LAYER M1 ;
        RECT 4.192 4.08 4.224 6.588 ;
  LAYER M3 ;
        RECT 4.192 6.536 4.224 6.568 ;
  LAYER M1 ;
        RECT 4.256 4.08 4.288 6.588 ;
  LAYER M3 ;
        RECT 4.256 4.1 4.288 4.132 ;
  LAYER M1 ;
        RECT 4.32 4.08 4.352 6.588 ;
  LAYER M3 ;
        RECT 4.32 6.536 4.352 6.568 ;
  LAYER M1 ;
        RECT 4.384 4.08 4.416 6.588 ;
  LAYER M3 ;
        RECT 4.384 4.1 4.416 4.132 ;
  LAYER M1 ;
        RECT 4.448 4.08 4.48 6.588 ;
  LAYER M3 ;
        RECT 4.448 6.536 4.48 6.568 ;
  LAYER M1 ;
        RECT 4.512 4.08 4.544 6.588 ;
  LAYER M3 ;
        RECT 4.512 4.1 4.544 4.132 ;
  LAYER M1 ;
        RECT 4.576 4.08 4.608 6.588 ;
  LAYER M3 ;
        RECT 4.576 6.536 4.608 6.568 ;
  LAYER M1 ;
        RECT 4.64 4.08 4.672 6.588 ;
  LAYER M3 ;
        RECT 4.64 4.1 4.672 4.132 ;
  LAYER M1 ;
        RECT 4.704 4.08 4.736 6.588 ;
  LAYER M3 ;
        RECT 4.704 6.536 4.736 6.568 ;
  LAYER M1 ;
        RECT 4.768 4.08 4.8 6.588 ;
  LAYER M3 ;
        RECT 4.768 4.1 4.8 4.132 ;
  LAYER M1 ;
        RECT 4.832 4.08 4.864 6.588 ;
  LAYER M3 ;
        RECT 4.832 6.536 4.864 6.568 ;
  LAYER M1 ;
        RECT 4.896 4.08 4.928 6.588 ;
  LAYER M3 ;
        RECT 4.896 4.1 4.928 4.132 ;
  LAYER M1 ;
        RECT 4.96 4.08 4.992 6.588 ;
  LAYER M3 ;
        RECT 4.96 6.536 4.992 6.568 ;
  LAYER M1 ;
        RECT 5.024 4.08 5.056 6.588 ;
  LAYER M3 ;
        RECT 5.024 4.1 5.056 4.132 ;
  LAYER M1 ;
        RECT 5.088 4.08 5.12 6.588 ;
  LAYER M3 ;
        RECT 5.088 6.536 5.12 6.568 ;
  LAYER M1 ;
        RECT 5.152 4.08 5.184 6.588 ;
  LAYER M3 ;
        RECT 5.152 4.1 5.184 4.132 ;
  LAYER M1 ;
        RECT 5.216 4.08 5.248 6.588 ;
  LAYER M3 ;
        RECT 5.216 6.536 5.248 6.568 ;
  LAYER M1 ;
        RECT 5.28 4.08 5.312 6.588 ;
  LAYER M3 ;
        RECT 5.28 4.1 5.312 4.132 ;
  LAYER M1 ;
        RECT 5.344 4.08 5.376 6.588 ;
  LAYER M3 ;
        RECT 5.344 6.536 5.376 6.568 ;
  LAYER M1 ;
        RECT 5.408 4.08 5.44 6.588 ;
  LAYER M3 ;
        RECT 5.408 4.1 5.44 4.132 ;
  LAYER M1 ;
        RECT 5.472 4.08 5.504 6.588 ;
  LAYER M3 ;
        RECT 5.472 6.536 5.504 6.568 ;
  LAYER M1 ;
        RECT 5.536 4.08 5.568 6.588 ;
  LAYER M3 ;
        RECT 5.536 4.1 5.568 4.132 ;
  LAYER M1 ;
        RECT 5.6 4.08 5.632 6.588 ;
  LAYER M3 ;
        RECT 5.6 6.536 5.632 6.568 ;
  LAYER M1 ;
        RECT 5.664 4.08 5.696 6.588 ;
  LAYER M3 ;
        RECT 5.664 4.1 5.696 4.132 ;
  LAYER M1 ;
        RECT 5.728 4.08 5.76 6.588 ;
  LAYER M3 ;
        RECT 5.728 6.536 5.76 6.568 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 6.588 ;
  LAYER M3 ;
        RECT 3.424 4.164 3.456 4.196 ;
  LAYER M2 ;
        RECT 5.792 4.228 5.824 4.26 ;
  LAYER M2 ;
        RECT 3.424 4.292 3.456 4.324 ;
  LAYER M2 ;
        RECT 5.792 4.356 5.824 4.388 ;
  LAYER M2 ;
        RECT 3.424 4.42 3.456 4.452 ;
  LAYER M2 ;
        RECT 5.792 4.484 5.824 4.516 ;
  LAYER M2 ;
        RECT 3.424 4.548 3.456 4.58 ;
  LAYER M2 ;
        RECT 5.792 4.612 5.824 4.644 ;
  LAYER M2 ;
        RECT 3.424 4.676 3.456 4.708 ;
  LAYER M2 ;
        RECT 5.792 4.74 5.824 4.772 ;
  LAYER M2 ;
        RECT 3.424 4.804 3.456 4.836 ;
  LAYER M2 ;
        RECT 5.792 4.868 5.824 4.9 ;
  LAYER M2 ;
        RECT 3.424 4.932 3.456 4.964 ;
  LAYER M2 ;
        RECT 5.792 4.996 5.824 5.028 ;
  LAYER M2 ;
        RECT 3.424 5.06 3.456 5.092 ;
  LAYER M2 ;
        RECT 5.792 5.124 5.824 5.156 ;
  LAYER M2 ;
        RECT 3.424 5.188 3.456 5.22 ;
  LAYER M2 ;
        RECT 5.792 5.252 5.824 5.284 ;
  LAYER M2 ;
        RECT 3.424 5.316 3.456 5.348 ;
  LAYER M2 ;
        RECT 5.792 5.38 5.824 5.412 ;
  LAYER M2 ;
        RECT 3.424 5.444 3.456 5.476 ;
  LAYER M2 ;
        RECT 5.792 5.508 5.824 5.54 ;
  LAYER M2 ;
        RECT 3.424 5.572 3.456 5.604 ;
  LAYER M2 ;
        RECT 5.792 5.636 5.824 5.668 ;
  LAYER M2 ;
        RECT 3.424 5.7 3.456 5.732 ;
  LAYER M2 ;
        RECT 5.792 5.764 5.824 5.796 ;
  LAYER M2 ;
        RECT 3.424 5.828 3.456 5.86 ;
  LAYER M2 ;
        RECT 5.792 5.892 5.824 5.924 ;
  LAYER M2 ;
        RECT 3.424 5.956 3.456 5.988 ;
  LAYER M2 ;
        RECT 5.792 6.02 5.824 6.052 ;
  LAYER M2 ;
        RECT 3.424 6.084 3.456 6.116 ;
  LAYER M2 ;
        RECT 5.792 6.148 5.824 6.18 ;
  LAYER M2 ;
        RECT 3.424 6.212 3.456 6.244 ;
  LAYER M2 ;
        RECT 5.792 6.276 5.824 6.308 ;
  LAYER M2 ;
        RECT 3.424 6.34 3.456 6.372 ;
  LAYER M2 ;
        RECT 5.792 6.404 5.824 6.436 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.424 7.188 3.456 9.696 ;
  LAYER M3 ;
        RECT 3.424 9.644 3.456 9.676 ;
  LAYER M1 ;
        RECT 3.488 7.188 3.52 9.696 ;
  LAYER M3 ;
        RECT 3.488 7.208 3.52 7.24 ;
  LAYER M1 ;
        RECT 3.552 7.188 3.584 9.696 ;
  LAYER M3 ;
        RECT 3.552 9.644 3.584 9.676 ;
  LAYER M1 ;
        RECT 3.616 7.188 3.648 9.696 ;
  LAYER M3 ;
        RECT 3.616 7.208 3.648 7.24 ;
  LAYER M1 ;
        RECT 3.68 7.188 3.712 9.696 ;
  LAYER M3 ;
        RECT 3.68 9.644 3.712 9.676 ;
  LAYER M1 ;
        RECT 3.744 7.188 3.776 9.696 ;
  LAYER M3 ;
        RECT 3.744 7.208 3.776 7.24 ;
  LAYER M1 ;
        RECT 3.808 7.188 3.84 9.696 ;
  LAYER M3 ;
        RECT 3.808 9.644 3.84 9.676 ;
  LAYER M1 ;
        RECT 3.872 7.188 3.904 9.696 ;
  LAYER M3 ;
        RECT 3.872 7.208 3.904 7.24 ;
  LAYER M1 ;
        RECT 3.936 7.188 3.968 9.696 ;
  LAYER M3 ;
        RECT 3.936 9.644 3.968 9.676 ;
  LAYER M1 ;
        RECT 4 7.188 4.032 9.696 ;
  LAYER M3 ;
        RECT 4 7.208 4.032 7.24 ;
  LAYER M1 ;
        RECT 4.064 7.188 4.096 9.696 ;
  LAYER M3 ;
        RECT 4.064 9.644 4.096 9.676 ;
  LAYER M1 ;
        RECT 4.128 7.188 4.16 9.696 ;
  LAYER M3 ;
        RECT 4.128 7.208 4.16 7.24 ;
  LAYER M1 ;
        RECT 4.192 7.188 4.224 9.696 ;
  LAYER M3 ;
        RECT 4.192 9.644 4.224 9.676 ;
  LAYER M1 ;
        RECT 4.256 7.188 4.288 9.696 ;
  LAYER M3 ;
        RECT 4.256 7.208 4.288 7.24 ;
  LAYER M1 ;
        RECT 4.32 7.188 4.352 9.696 ;
  LAYER M3 ;
        RECT 4.32 9.644 4.352 9.676 ;
  LAYER M1 ;
        RECT 4.384 7.188 4.416 9.696 ;
  LAYER M3 ;
        RECT 4.384 7.208 4.416 7.24 ;
  LAYER M1 ;
        RECT 4.448 7.188 4.48 9.696 ;
  LAYER M3 ;
        RECT 4.448 9.644 4.48 9.676 ;
  LAYER M1 ;
        RECT 4.512 7.188 4.544 9.696 ;
  LAYER M3 ;
        RECT 4.512 7.208 4.544 7.24 ;
  LAYER M1 ;
        RECT 4.576 7.188 4.608 9.696 ;
  LAYER M3 ;
        RECT 4.576 9.644 4.608 9.676 ;
  LAYER M1 ;
        RECT 4.64 7.188 4.672 9.696 ;
  LAYER M3 ;
        RECT 4.64 7.208 4.672 7.24 ;
  LAYER M1 ;
        RECT 4.704 7.188 4.736 9.696 ;
  LAYER M3 ;
        RECT 4.704 9.644 4.736 9.676 ;
  LAYER M1 ;
        RECT 4.768 7.188 4.8 9.696 ;
  LAYER M3 ;
        RECT 4.768 7.208 4.8 7.24 ;
  LAYER M1 ;
        RECT 4.832 7.188 4.864 9.696 ;
  LAYER M3 ;
        RECT 4.832 9.644 4.864 9.676 ;
  LAYER M1 ;
        RECT 4.896 7.188 4.928 9.696 ;
  LAYER M3 ;
        RECT 4.896 7.208 4.928 7.24 ;
  LAYER M1 ;
        RECT 4.96 7.188 4.992 9.696 ;
  LAYER M3 ;
        RECT 4.96 9.644 4.992 9.676 ;
  LAYER M1 ;
        RECT 5.024 7.188 5.056 9.696 ;
  LAYER M3 ;
        RECT 5.024 7.208 5.056 7.24 ;
  LAYER M1 ;
        RECT 5.088 7.188 5.12 9.696 ;
  LAYER M3 ;
        RECT 5.088 9.644 5.12 9.676 ;
  LAYER M1 ;
        RECT 5.152 7.188 5.184 9.696 ;
  LAYER M3 ;
        RECT 5.152 7.208 5.184 7.24 ;
  LAYER M1 ;
        RECT 5.216 7.188 5.248 9.696 ;
  LAYER M3 ;
        RECT 5.216 9.644 5.248 9.676 ;
  LAYER M1 ;
        RECT 5.28 7.188 5.312 9.696 ;
  LAYER M3 ;
        RECT 5.28 7.208 5.312 7.24 ;
  LAYER M1 ;
        RECT 5.344 7.188 5.376 9.696 ;
  LAYER M3 ;
        RECT 5.344 9.644 5.376 9.676 ;
  LAYER M1 ;
        RECT 5.408 7.188 5.44 9.696 ;
  LAYER M3 ;
        RECT 5.408 7.208 5.44 7.24 ;
  LAYER M1 ;
        RECT 5.472 7.188 5.504 9.696 ;
  LAYER M3 ;
        RECT 5.472 9.644 5.504 9.676 ;
  LAYER M1 ;
        RECT 5.536 7.188 5.568 9.696 ;
  LAYER M3 ;
        RECT 5.536 7.208 5.568 7.24 ;
  LAYER M1 ;
        RECT 5.6 7.188 5.632 9.696 ;
  LAYER M3 ;
        RECT 5.6 9.644 5.632 9.676 ;
  LAYER M1 ;
        RECT 5.664 7.188 5.696 9.696 ;
  LAYER M3 ;
        RECT 5.664 7.208 5.696 7.24 ;
  LAYER M1 ;
        RECT 5.728 7.188 5.76 9.696 ;
  LAYER M3 ;
        RECT 5.728 9.644 5.76 9.676 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 9.696 ;
  LAYER M3 ;
        RECT 3.424 7.272 3.456 7.304 ;
  LAYER M2 ;
        RECT 5.792 7.336 5.824 7.368 ;
  LAYER M2 ;
        RECT 3.424 7.4 3.456 7.432 ;
  LAYER M2 ;
        RECT 5.792 7.464 5.824 7.496 ;
  LAYER M2 ;
        RECT 3.424 7.528 3.456 7.56 ;
  LAYER M2 ;
        RECT 5.792 7.592 5.824 7.624 ;
  LAYER M2 ;
        RECT 3.424 7.656 3.456 7.688 ;
  LAYER M2 ;
        RECT 5.792 7.72 5.824 7.752 ;
  LAYER M2 ;
        RECT 3.424 7.784 3.456 7.816 ;
  LAYER M2 ;
        RECT 5.792 7.848 5.824 7.88 ;
  LAYER M2 ;
        RECT 3.424 7.912 3.456 7.944 ;
  LAYER M2 ;
        RECT 5.792 7.976 5.824 8.008 ;
  LAYER M2 ;
        RECT 3.424 8.04 3.456 8.072 ;
  LAYER M2 ;
        RECT 5.792 8.104 5.824 8.136 ;
  LAYER M2 ;
        RECT 3.424 8.168 3.456 8.2 ;
  LAYER M2 ;
        RECT 5.792 8.232 5.824 8.264 ;
  LAYER M2 ;
        RECT 3.424 8.296 3.456 8.328 ;
  LAYER M2 ;
        RECT 5.792 8.36 5.824 8.392 ;
  LAYER M2 ;
        RECT 3.424 8.424 3.456 8.456 ;
  LAYER M2 ;
        RECT 5.792 8.488 5.824 8.52 ;
  LAYER M2 ;
        RECT 3.424 8.552 3.456 8.584 ;
  LAYER M2 ;
        RECT 5.792 8.616 5.824 8.648 ;
  LAYER M2 ;
        RECT 3.424 8.68 3.456 8.712 ;
  LAYER M2 ;
        RECT 5.792 8.744 5.824 8.776 ;
  LAYER M2 ;
        RECT 3.424 8.808 3.456 8.84 ;
  LAYER M2 ;
        RECT 5.792 8.872 5.824 8.904 ;
  LAYER M2 ;
        RECT 3.424 8.936 3.456 8.968 ;
  LAYER M2 ;
        RECT 5.792 9 5.824 9.032 ;
  LAYER M2 ;
        RECT 3.424 9.064 3.456 9.096 ;
  LAYER M2 ;
        RECT 5.792 9.128 5.824 9.16 ;
  LAYER M2 ;
        RECT 3.424 9.192 3.456 9.224 ;
  LAYER M2 ;
        RECT 5.792 9.256 5.824 9.288 ;
  LAYER M2 ;
        RECT 3.424 9.32 3.456 9.352 ;
  LAYER M2 ;
        RECT 5.792 9.384 5.824 9.416 ;
  LAYER M2 ;
        RECT 3.424 9.448 3.456 9.48 ;
  LAYER M2 ;
        RECT 5.792 9.512 5.824 9.544 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.424 10.296 3.456 12.804 ;
  LAYER M3 ;
        RECT 3.424 12.752 3.456 12.784 ;
  LAYER M1 ;
        RECT 3.488 10.296 3.52 12.804 ;
  LAYER M3 ;
        RECT 3.488 10.316 3.52 10.348 ;
  LAYER M1 ;
        RECT 3.552 10.296 3.584 12.804 ;
  LAYER M3 ;
        RECT 3.552 12.752 3.584 12.784 ;
  LAYER M1 ;
        RECT 3.616 10.296 3.648 12.804 ;
  LAYER M3 ;
        RECT 3.616 10.316 3.648 10.348 ;
  LAYER M1 ;
        RECT 3.68 10.296 3.712 12.804 ;
  LAYER M3 ;
        RECT 3.68 12.752 3.712 12.784 ;
  LAYER M1 ;
        RECT 3.744 10.296 3.776 12.804 ;
  LAYER M3 ;
        RECT 3.744 10.316 3.776 10.348 ;
  LAYER M1 ;
        RECT 3.808 10.296 3.84 12.804 ;
  LAYER M3 ;
        RECT 3.808 12.752 3.84 12.784 ;
  LAYER M1 ;
        RECT 3.872 10.296 3.904 12.804 ;
  LAYER M3 ;
        RECT 3.872 10.316 3.904 10.348 ;
  LAYER M1 ;
        RECT 3.936 10.296 3.968 12.804 ;
  LAYER M3 ;
        RECT 3.936 12.752 3.968 12.784 ;
  LAYER M1 ;
        RECT 4 10.296 4.032 12.804 ;
  LAYER M3 ;
        RECT 4 10.316 4.032 10.348 ;
  LAYER M1 ;
        RECT 4.064 10.296 4.096 12.804 ;
  LAYER M3 ;
        RECT 4.064 12.752 4.096 12.784 ;
  LAYER M1 ;
        RECT 4.128 10.296 4.16 12.804 ;
  LAYER M3 ;
        RECT 4.128 10.316 4.16 10.348 ;
  LAYER M1 ;
        RECT 4.192 10.296 4.224 12.804 ;
  LAYER M3 ;
        RECT 4.192 12.752 4.224 12.784 ;
  LAYER M1 ;
        RECT 4.256 10.296 4.288 12.804 ;
  LAYER M3 ;
        RECT 4.256 10.316 4.288 10.348 ;
  LAYER M1 ;
        RECT 4.32 10.296 4.352 12.804 ;
  LAYER M3 ;
        RECT 4.32 12.752 4.352 12.784 ;
  LAYER M1 ;
        RECT 4.384 10.296 4.416 12.804 ;
  LAYER M3 ;
        RECT 4.384 10.316 4.416 10.348 ;
  LAYER M1 ;
        RECT 4.448 10.296 4.48 12.804 ;
  LAYER M3 ;
        RECT 4.448 12.752 4.48 12.784 ;
  LAYER M1 ;
        RECT 4.512 10.296 4.544 12.804 ;
  LAYER M3 ;
        RECT 4.512 10.316 4.544 10.348 ;
  LAYER M1 ;
        RECT 4.576 10.296 4.608 12.804 ;
  LAYER M3 ;
        RECT 4.576 12.752 4.608 12.784 ;
  LAYER M1 ;
        RECT 4.64 10.296 4.672 12.804 ;
  LAYER M3 ;
        RECT 4.64 10.316 4.672 10.348 ;
  LAYER M1 ;
        RECT 4.704 10.296 4.736 12.804 ;
  LAYER M3 ;
        RECT 4.704 12.752 4.736 12.784 ;
  LAYER M1 ;
        RECT 4.768 10.296 4.8 12.804 ;
  LAYER M3 ;
        RECT 4.768 10.316 4.8 10.348 ;
  LAYER M1 ;
        RECT 4.832 10.296 4.864 12.804 ;
  LAYER M3 ;
        RECT 4.832 12.752 4.864 12.784 ;
  LAYER M1 ;
        RECT 4.896 10.296 4.928 12.804 ;
  LAYER M3 ;
        RECT 4.896 10.316 4.928 10.348 ;
  LAYER M1 ;
        RECT 4.96 10.296 4.992 12.804 ;
  LAYER M3 ;
        RECT 4.96 12.752 4.992 12.784 ;
  LAYER M1 ;
        RECT 5.024 10.296 5.056 12.804 ;
  LAYER M3 ;
        RECT 5.024 10.316 5.056 10.348 ;
  LAYER M1 ;
        RECT 5.088 10.296 5.12 12.804 ;
  LAYER M3 ;
        RECT 5.088 12.752 5.12 12.784 ;
  LAYER M1 ;
        RECT 5.152 10.296 5.184 12.804 ;
  LAYER M3 ;
        RECT 5.152 10.316 5.184 10.348 ;
  LAYER M1 ;
        RECT 5.216 10.296 5.248 12.804 ;
  LAYER M3 ;
        RECT 5.216 12.752 5.248 12.784 ;
  LAYER M1 ;
        RECT 5.28 10.296 5.312 12.804 ;
  LAYER M3 ;
        RECT 5.28 10.316 5.312 10.348 ;
  LAYER M1 ;
        RECT 5.344 10.296 5.376 12.804 ;
  LAYER M3 ;
        RECT 5.344 12.752 5.376 12.784 ;
  LAYER M1 ;
        RECT 5.408 10.296 5.44 12.804 ;
  LAYER M3 ;
        RECT 5.408 10.316 5.44 10.348 ;
  LAYER M1 ;
        RECT 5.472 10.296 5.504 12.804 ;
  LAYER M3 ;
        RECT 5.472 12.752 5.504 12.784 ;
  LAYER M1 ;
        RECT 5.536 10.296 5.568 12.804 ;
  LAYER M3 ;
        RECT 5.536 10.316 5.568 10.348 ;
  LAYER M1 ;
        RECT 5.6 10.296 5.632 12.804 ;
  LAYER M3 ;
        RECT 5.6 12.752 5.632 12.784 ;
  LAYER M1 ;
        RECT 5.664 10.296 5.696 12.804 ;
  LAYER M3 ;
        RECT 5.664 10.316 5.696 10.348 ;
  LAYER M1 ;
        RECT 5.728 10.296 5.76 12.804 ;
  LAYER M3 ;
        RECT 5.728 12.752 5.76 12.784 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 12.804 ;
  LAYER M3 ;
        RECT 3.424 10.38 3.456 10.412 ;
  LAYER M2 ;
        RECT 5.792 10.444 5.824 10.476 ;
  LAYER M2 ;
        RECT 3.424 10.508 3.456 10.54 ;
  LAYER M2 ;
        RECT 5.792 10.572 5.824 10.604 ;
  LAYER M2 ;
        RECT 3.424 10.636 3.456 10.668 ;
  LAYER M2 ;
        RECT 5.792 10.7 5.824 10.732 ;
  LAYER M2 ;
        RECT 3.424 10.764 3.456 10.796 ;
  LAYER M2 ;
        RECT 5.792 10.828 5.824 10.86 ;
  LAYER M2 ;
        RECT 3.424 10.892 3.456 10.924 ;
  LAYER M2 ;
        RECT 5.792 10.956 5.824 10.988 ;
  LAYER M2 ;
        RECT 3.424 11.02 3.456 11.052 ;
  LAYER M2 ;
        RECT 5.792 11.084 5.824 11.116 ;
  LAYER M2 ;
        RECT 3.424 11.148 3.456 11.18 ;
  LAYER M2 ;
        RECT 5.792 11.212 5.824 11.244 ;
  LAYER M2 ;
        RECT 3.424 11.276 3.456 11.308 ;
  LAYER M2 ;
        RECT 5.792 11.34 5.824 11.372 ;
  LAYER M2 ;
        RECT 3.424 11.404 3.456 11.436 ;
  LAYER M2 ;
        RECT 5.792 11.468 5.824 11.5 ;
  LAYER M2 ;
        RECT 3.424 11.532 3.456 11.564 ;
  LAYER M2 ;
        RECT 5.792 11.596 5.824 11.628 ;
  LAYER M2 ;
        RECT 3.424 11.66 3.456 11.692 ;
  LAYER M2 ;
        RECT 5.792 11.724 5.824 11.756 ;
  LAYER M2 ;
        RECT 3.424 11.788 3.456 11.82 ;
  LAYER M2 ;
        RECT 5.792 11.852 5.824 11.884 ;
  LAYER M2 ;
        RECT 3.424 11.916 3.456 11.948 ;
  LAYER M2 ;
        RECT 5.792 11.98 5.824 12.012 ;
  LAYER M2 ;
        RECT 3.424 12.044 3.456 12.076 ;
  LAYER M2 ;
        RECT 5.792 12.108 5.824 12.14 ;
  LAYER M2 ;
        RECT 3.424 12.172 3.456 12.204 ;
  LAYER M2 ;
        RECT 5.792 12.236 5.824 12.268 ;
  LAYER M2 ;
        RECT 3.424 12.3 3.456 12.332 ;
  LAYER M2 ;
        RECT 5.792 12.364 5.824 12.396 ;
  LAYER M2 ;
        RECT 3.424 12.428 3.456 12.46 ;
  LAYER M2 ;
        RECT 5.792 12.492 5.824 12.524 ;
  LAYER M2 ;
        RECT 3.424 12.556 3.456 12.588 ;
  LAYER M2 ;
        RECT 5.792 12.62 5.824 12.652 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 3.424 13.404 3.456 15.912 ;
  LAYER M3 ;
        RECT 3.424 15.86 3.456 15.892 ;
  LAYER M1 ;
        RECT 3.488 13.404 3.52 15.912 ;
  LAYER M3 ;
        RECT 3.488 13.424 3.52 13.456 ;
  LAYER M1 ;
        RECT 3.552 13.404 3.584 15.912 ;
  LAYER M3 ;
        RECT 3.552 15.86 3.584 15.892 ;
  LAYER M1 ;
        RECT 3.616 13.404 3.648 15.912 ;
  LAYER M3 ;
        RECT 3.616 13.424 3.648 13.456 ;
  LAYER M1 ;
        RECT 3.68 13.404 3.712 15.912 ;
  LAYER M3 ;
        RECT 3.68 15.86 3.712 15.892 ;
  LAYER M1 ;
        RECT 3.744 13.404 3.776 15.912 ;
  LAYER M3 ;
        RECT 3.744 13.424 3.776 13.456 ;
  LAYER M1 ;
        RECT 3.808 13.404 3.84 15.912 ;
  LAYER M3 ;
        RECT 3.808 15.86 3.84 15.892 ;
  LAYER M1 ;
        RECT 3.872 13.404 3.904 15.912 ;
  LAYER M3 ;
        RECT 3.872 13.424 3.904 13.456 ;
  LAYER M1 ;
        RECT 3.936 13.404 3.968 15.912 ;
  LAYER M3 ;
        RECT 3.936 15.86 3.968 15.892 ;
  LAYER M1 ;
        RECT 4 13.404 4.032 15.912 ;
  LAYER M3 ;
        RECT 4 13.424 4.032 13.456 ;
  LAYER M1 ;
        RECT 4.064 13.404 4.096 15.912 ;
  LAYER M3 ;
        RECT 4.064 15.86 4.096 15.892 ;
  LAYER M1 ;
        RECT 4.128 13.404 4.16 15.912 ;
  LAYER M3 ;
        RECT 4.128 13.424 4.16 13.456 ;
  LAYER M1 ;
        RECT 4.192 13.404 4.224 15.912 ;
  LAYER M3 ;
        RECT 4.192 15.86 4.224 15.892 ;
  LAYER M1 ;
        RECT 4.256 13.404 4.288 15.912 ;
  LAYER M3 ;
        RECT 4.256 13.424 4.288 13.456 ;
  LAYER M1 ;
        RECT 4.32 13.404 4.352 15.912 ;
  LAYER M3 ;
        RECT 4.32 15.86 4.352 15.892 ;
  LAYER M1 ;
        RECT 4.384 13.404 4.416 15.912 ;
  LAYER M3 ;
        RECT 4.384 13.424 4.416 13.456 ;
  LAYER M1 ;
        RECT 4.448 13.404 4.48 15.912 ;
  LAYER M3 ;
        RECT 4.448 15.86 4.48 15.892 ;
  LAYER M1 ;
        RECT 4.512 13.404 4.544 15.912 ;
  LAYER M3 ;
        RECT 4.512 13.424 4.544 13.456 ;
  LAYER M1 ;
        RECT 4.576 13.404 4.608 15.912 ;
  LAYER M3 ;
        RECT 4.576 15.86 4.608 15.892 ;
  LAYER M1 ;
        RECT 4.64 13.404 4.672 15.912 ;
  LAYER M3 ;
        RECT 4.64 13.424 4.672 13.456 ;
  LAYER M1 ;
        RECT 4.704 13.404 4.736 15.912 ;
  LAYER M3 ;
        RECT 4.704 15.86 4.736 15.892 ;
  LAYER M1 ;
        RECT 4.768 13.404 4.8 15.912 ;
  LAYER M3 ;
        RECT 4.768 13.424 4.8 13.456 ;
  LAYER M1 ;
        RECT 4.832 13.404 4.864 15.912 ;
  LAYER M3 ;
        RECT 4.832 15.86 4.864 15.892 ;
  LAYER M1 ;
        RECT 4.896 13.404 4.928 15.912 ;
  LAYER M3 ;
        RECT 4.896 13.424 4.928 13.456 ;
  LAYER M1 ;
        RECT 4.96 13.404 4.992 15.912 ;
  LAYER M3 ;
        RECT 4.96 15.86 4.992 15.892 ;
  LAYER M1 ;
        RECT 5.024 13.404 5.056 15.912 ;
  LAYER M3 ;
        RECT 5.024 13.424 5.056 13.456 ;
  LAYER M1 ;
        RECT 5.088 13.404 5.12 15.912 ;
  LAYER M3 ;
        RECT 5.088 15.86 5.12 15.892 ;
  LAYER M1 ;
        RECT 5.152 13.404 5.184 15.912 ;
  LAYER M3 ;
        RECT 5.152 13.424 5.184 13.456 ;
  LAYER M1 ;
        RECT 5.216 13.404 5.248 15.912 ;
  LAYER M3 ;
        RECT 5.216 15.86 5.248 15.892 ;
  LAYER M1 ;
        RECT 5.28 13.404 5.312 15.912 ;
  LAYER M3 ;
        RECT 5.28 13.424 5.312 13.456 ;
  LAYER M1 ;
        RECT 5.344 13.404 5.376 15.912 ;
  LAYER M3 ;
        RECT 5.344 15.86 5.376 15.892 ;
  LAYER M1 ;
        RECT 5.408 13.404 5.44 15.912 ;
  LAYER M3 ;
        RECT 5.408 13.424 5.44 13.456 ;
  LAYER M1 ;
        RECT 5.472 13.404 5.504 15.912 ;
  LAYER M3 ;
        RECT 5.472 15.86 5.504 15.892 ;
  LAYER M1 ;
        RECT 5.536 13.404 5.568 15.912 ;
  LAYER M3 ;
        RECT 5.536 13.424 5.568 13.456 ;
  LAYER M1 ;
        RECT 5.6 13.404 5.632 15.912 ;
  LAYER M3 ;
        RECT 5.6 15.86 5.632 15.892 ;
  LAYER M1 ;
        RECT 5.664 13.404 5.696 15.912 ;
  LAYER M3 ;
        RECT 5.664 13.424 5.696 13.456 ;
  LAYER M1 ;
        RECT 5.728 13.404 5.76 15.912 ;
  LAYER M3 ;
        RECT 5.728 15.86 5.76 15.892 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 15.912 ;
  LAYER M3 ;
        RECT 3.424 13.488 3.456 13.52 ;
  LAYER M2 ;
        RECT 5.792 13.552 5.824 13.584 ;
  LAYER M2 ;
        RECT 3.424 13.616 3.456 13.648 ;
  LAYER M2 ;
        RECT 5.792 13.68 5.824 13.712 ;
  LAYER M2 ;
        RECT 3.424 13.744 3.456 13.776 ;
  LAYER M2 ;
        RECT 5.792 13.808 5.824 13.84 ;
  LAYER M2 ;
        RECT 3.424 13.872 3.456 13.904 ;
  LAYER M2 ;
        RECT 5.792 13.936 5.824 13.968 ;
  LAYER M2 ;
        RECT 3.424 14 3.456 14.032 ;
  LAYER M2 ;
        RECT 5.792 14.064 5.824 14.096 ;
  LAYER M2 ;
        RECT 3.424 14.128 3.456 14.16 ;
  LAYER M2 ;
        RECT 5.792 14.192 5.824 14.224 ;
  LAYER M2 ;
        RECT 3.424 14.256 3.456 14.288 ;
  LAYER M2 ;
        RECT 5.792 14.32 5.824 14.352 ;
  LAYER M2 ;
        RECT 3.424 14.384 3.456 14.416 ;
  LAYER M2 ;
        RECT 5.792 14.448 5.824 14.48 ;
  LAYER M2 ;
        RECT 3.424 14.512 3.456 14.544 ;
  LAYER M2 ;
        RECT 5.792 14.576 5.824 14.608 ;
  LAYER M2 ;
        RECT 3.424 14.64 3.456 14.672 ;
  LAYER M2 ;
        RECT 5.792 14.704 5.824 14.736 ;
  LAYER M2 ;
        RECT 3.424 14.768 3.456 14.8 ;
  LAYER M2 ;
        RECT 5.792 14.832 5.824 14.864 ;
  LAYER M2 ;
        RECT 3.424 14.896 3.456 14.928 ;
  LAYER M2 ;
        RECT 5.792 14.96 5.824 14.992 ;
  LAYER M2 ;
        RECT 3.424 15.024 3.456 15.056 ;
  LAYER M2 ;
        RECT 5.792 15.088 5.824 15.12 ;
  LAYER M2 ;
        RECT 3.424 15.152 3.456 15.184 ;
  LAYER M2 ;
        RECT 5.792 15.216 5.824 15.248 ;
  LAYER M2 ;
        RECT 3.424 15.28 3.456 15.312 ;
  LAYER M2 ;
        RECT 5.792 15.344 5.824 15.376 ;
  LAYER M2 ;
        RECT 3.424 15.408 3.456 15.44 ;
  LAYER M2 ;
        RECT 5.792 15.472 5.824 15.504 ;
  LAYER M2 ;
        RECT 3.424 15.536 3.456 15.568 ;
  LAYER M2 ;
        RECT 5.792 15.6 5.824 15.632 ;
  LAYER M2 ;
        RECT 3.424 15.664 3.456 15.696 ;
  LAYER M2 ;
        RECT 5.792 15.728 5.824 15.76 ;
  LAYER M2 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M1 ;
        RECT 6.4 0.972 6.432 3.48 ;
  LAYER M3 ;
        RECT 6.4 3.428 6.432 3.46 ;
  LAYER M1 ;
        RECT 6.464 0.972 6.496 3.48 ;
  LAYER M3 ;
        RECT 6.464 0.992 6.496 1.024 ;
  LAYER M1 ;
        RECT 6.528 0.972 6.56 3.48 ;
  LAYER M3 ;
        RECT 6.528 3.428 6.56 3.46 ;
  LAYER M1 ;
        RECT 6.592 0.972 6.624 3.48 ;
  LAYER M3 ;
        RECT 6.592 0.992 6.624 1.024 ;
  LAYER M1 ;
        RECT 6.656 0.972 6.688 3.48 ;
  LAYER M3 ;
        RECT 6.656 3.428 6.688 3.46 ;
  LAYER M1 ;
        RECT 6.72 0.972 6.752 3.48 ;
  LAYER M3 ;
        RECT 6.72 0.992 6.752 1.024 ;
  LAYER M1 ;
        RECT 6.784 0.972 6.816 3.48 ;
  LAYER M3 ;
        RECT 6.784 3.428 6.816 3.46 ;
  LAYER M1 ;
        RECT 6.848 0.972 6.88 3.48 ;
  LAYER M3 ;
        RECT 6.848 0.992 6.88 1.024 ;
  LAYER M1 ;
        RECT 6.912 0.972 6.944 3.48 ;
  LAYER M3 ;
        RECT 6.912 3.428 6.944 3.46 ;
  LAYER M1 ;
        RECT 6.976 0.972 7.008 3.48 ;
  LAYER M3 ;
        RECT 6.976 0.992 7.008 1.024 ;
  LAYER M1 ;
        RECT 7.04 0.972 7.072 3.48 ;
  LAYER M3 ;
        RECT 7.04 3.428 7.072 3.46 ;
  LAYER M1 ;
        RECT 7.104 0.972 7.136 3.48 ;
  LAYER M3 ;
        RECT 7.104 0.992 7.136 1.024 ;
  LAYER M1 ;
        RECT 7.168 0.972 7.2 3.48 ;
  LAYER M3 ;
        RECT 7.168 3.428 7.2 3.46 ;
  LAYER M1 ;
        RECT 7.232 0.972 7.264 3.48 ;
  LAYER M3 ;
        RECT 7.232 0.992 7.264 1.024 ;
  LAYER M1 ;
        RECT 7.296 0.972 7.328 3.48 ;
  LAYER M3 ;
        RECT 7.296 3.428 7.328 3.46 ;
  LAYER M1 ;
        RECT 7.36 0.972 7.392 3.48 ;
  LAYER M3 ;
        RECT 7.36 0.992 7.392 1.024 ;
  LAYER M1 ;
        RECT 7.424 0.972 7.456 3.48 ;
  LAYER M3 ;
        RECT 7.424 3.428 7.456 3.46 ;
  LAYER M1 ;
        RECT 7.488 0.972 7.52 3.48 ;
  LAYER M3 ;
        RECT 7.488 0.992 7.52 1.024 ;
  LAYER M1 ;
        RECT 7.552 0.972 7.584 3.48 ;
  LAYER M3 ;
        RECT 7.552 3.428 7.584 3.46 ;
  LAYER M1 ;
        RECT 7.616 0.972 7.648 3.48 ;
  LAYER M3 ;
        RECT 7.616 0.992 7.648 1.024 ;
  LAYER M1 ;
        RECT 7.68 0.972 7.712 3.48 ;
  LAYER M3 ;
        RECT 7.68 3.428 7.712 3.46 ;
  LAYER M1 ;
        RECT 7.744 0.972 7.776 3.48 ;
  LAYER M3 ;
        RECT 7.744 0.992 7.776 1.024 ;
  LAYER M1 ;
        RECT 7.808 0.972 7.84 3.48 ;
  LAYER M3 ;
        RECT 7.808 3.428 7.84 3.46 ;
  LAYER M1 ;
        RECT 7.872 0.972 7.904 3.48 ;
  LAYER M3 ;
        RECT 7.872 0.992 7.904 1.024 ;
  LAYER M1 ;
        RECT 7.936 0.972 7.968 3.48 ;
  LAYER M3 ;
        RECT 7.936 3.428 7.968 3.46 ;
  LAYER M1 ;
        RECT 8 0.972 8.032 3.48 ;
  LAYER M3 ;
        RECT 8 0.992 8.032 1.024 ;
  LAYER M1 ;
        RECT 8.064 0.972 8.096 3.48 ;
  LAYER M3 ;
        RECT 8.064 3.428 8.096 3.46 ;
  LAYER M1 ;
        RECT 8.128 0.972 8.16 3.48 ;
  LAYER M3 ;
        RECT 8.128 0.992 8.16 1.024 ;
  LAYER M1 ;
        RECT 8.192 0.972 8.224 3.48 ;
  LAYER M3 ;
        RECT 8.192 3.428 8.224 3.46 ;
  LAYER M1 ;
        RECT 8.256 0.972 8.288 3.48 ;
  LAYER M3 ;
        RECT 8.256 0.992 8.288 1.024 ;
  LAYER M1 ;
        RECT 8.32 0.972 8.352 3.48 ;
  LAYER M3 ;
        RECT 8.32 3.428 8.352 3.46 ;
  LAYER M1 ;
        RECT 8.384 0.972 8.416 3.48 ;
  LAYER M3 ;
        RECT 8.384 0.992 8.416 1.024 ;
  LAYER M1 ;
        RECT 8.448 0.972 8.48 3.48 ;
  LAYER M3 ;
        RECT 8.448 3.428 8.48 3.46 ;
  LAYER M1 ;
        RECT 8.512 0.972 8.544 3.48 ;
  LAYER M3 ;
        RECT 8.512 0.992 8.544 1.024 ;
  LAYER M1 ;
        RECT 8.576 0.972 8.608 3.48 ;
  LAYER M3 ;
        RECT 8.576 3.428 8.608 3.46 ;
  LAYER M1 ;
        RECT 8.64 0.972 8.672 3.48 ;
  LAYER M3 ;
        RECT 8.64 0.992 8.672 1.024 ;
  LAYER M1 ;
        RECT 8.704 0.972 8.736 3.48 ;
  LAYER M3 ;
        RECT 8.704 3.428 8.736 3.46 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 3.48 ;
  LAYER M3 ;
        RECT 6.4 1.056 6.432 1.088 ;
  LAYER M2 ;
        RECT 8.768 1.12 8.8 1.152 ;
  LAYER M2 ;
        RECT 6.4 1.184 6.432 1.216 ;
  LAYER M2 ;
        RECT 8.768 1.248 8.8 1.28 ;
  LAYER M2 ;
        RECT 6.4 1.312 6.432 1.344 ;
  LAYER M2 ;
        RECT 8.768 1.376 8.8 1.408 ;
  LAYER M2 ;
        RECT 6.4 1.44 6.432 1.472 ;
  LAYER M2 ;
        RECT 8.768 1.504 8.8 1.536 ;
  LAYER M2 ;
        RECT 6.4 1.568 6.432 1.6 ;
  LAYER M2 ;
        RECT 8.768 1.632 8.8 1.664 ;
  LAYER M2 ;
        RECT 6.4 1.696 6.432 1.728 ;
  LAYER M2 ;
        RECT 8.768 1.76 8.8 1.792 ;
  LAYER M2 ;
        RECT 6.4 1.824 6.432 1.856 ;
  LAYER M2 ;
        RECT 8.768 1.888 8.8 1.92 ;
  LAYER M2 ;
        RECT 6.4 1.952 6.432 1.984 ;
  LAYER M2 ;
        RECT 8.768 2.016 8.8 2.048 ;
  LAYER M2 ;
        RECT 6.4 2.08 6.432 2.112 ;
  LAYER M2 ;
        RECT 8.768 2.144 8.8 2.176 ;
  LAYER M2 ;
        RECT 6.4 2.208 6.432 2.24 ;
  LAYER M2 ;
        RECT 8.768 2.272 8.8 2.304 ;
  LAYER M2 ;
        RECT 6.4 2.336 6.432 2.368 ;
  LAYER M2 ;
        RECT 8.768 2.4 8.8 2.432 ;
  LAYER M2 ;
        RECT 6.4 2.464 6.432 2.496 ;
  LAYER M2 ;
        RECT 8.768 2.528 8.8 2.56 ;
  LAYER M2 ;
        RECT 6.4 2.592 6.432 2.624 ;
  LAYER M2 ;
        RECT 8.768 2.656 8.8 2.688 ;
  LAYER M2 ;
        RECT 6.4 2.72 6.432 2.752 ;
  LAYER M2 ;
        RECT 8.768 2.784 8.8 2.816 ;
  LAYER M2 ;
        RECT 6.4 2.848 6.432 2.88 ;
  LAYER M2 ;
        RECT 8.768 2.912 8.8 2.944 ;
  LAYER M2 ;
        RECT 6.4 2.976 6.432 3.008 ;
  LAYER M2 ;
        RECT 8.768 3.04 8.8 3.072 ;
  LAYER M2 ;
        RECT 6.4 3.104 6.432 3.136 ;
  LAYER M2 ;
        RECT 8.768 3.168 8.8 3.2 ;
  LAYER M2 ;
        RECT 6.4 3.232 6.432 3.264 ;
  LAYER M2 ;
        RECT 8.768 3.296 8.8 3.328 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.4 4.08 6.432 6.588 ;
  LAYER M3 ;
        RECT 6.4 6.536 6.432 6.568 ;
  LAYER M1 ;
        RECT 6.464 4.08 6.496 6.588 ;
  LAYER M3 ;
        RECT 6.464 4.1 6.496 4.132 ;
  LAYER M1 ;
        RECT 6.528 4.08 6.56 6.588 ;
  LAYER M3 ;
        RECT 6.528 6.536 6.56 6.568 ;
  LAYER M1 ;
        RECT 6.592 4.08 6.624 6.588 ;
  LAYER M3 ;
        RECT 6.592 4.1 6.624 4.132 ;
  LAYER M1 ;
        RECT 6.656 4.08 6.688 6.588 ;
  LAYER M3 ;
        RECT 6.656 6.536 6.688 6.568 ;
  LAYER M1 ;
        RECT 6.72 4.08 6.752 6.588 ;
  LAYER M3 ;
        RECT 6.72 4.1 6.752 4.132 ;
  LAYER M1 ;
        RECT 6.784 4.08 6.816 6.588 ;
  LAYER M3 ;
        RECT 6.784 6.536 6.816 6.568 ;
  LAYER M1 ;
        RECT 6.848 4.08 6.88 6.588 ;
  LAYER M3 ;
        RECT 6.848 4.1 6.88 4.132 ;
  LAYER M1 ;
        RECT 6.912 4.08 6.944 6.588 ;
  LAYER M3 ;
        RECT 6.912 6.536 6.944 6.568 ;
  LAYER M1 ;
        RECT 6.976 4.08 7.008 6.588 ;
  LAYER M3 ;
        RECT 6.976 4.1 7.008 4.132 ;
  LAYER M1 ;
        RECT 7.04 4.08 7.072 6.588 ;
  LAYER M3 ;
        RECT 7.04 6.536 7.072 6.568 ;
  LAYER M1 ;
        RECT 7.104 4.08 7.136 6.588 ;
  LAYER M3 ;
        RECT 7.104 4.1 7.136 4.132 ;
  LAYER M1 ;
        RECT 7.168 4.08 7.2 6.588 ;
  LAYER M3 ;
        RECT 7.168 6.536 7.2 6.568 ;
  LAYER M1 ;
        RECT 7.232 4.08 7.264 6.588 ;
  LAYER M3 ;
        RECT 7.232 4.1 7.264 4.132 ;
  LAYER M1 ;
        RECT 7.296 4.08 7.328 6.588 ;
  LAYER M3 ;
        RECT 7.296 6.536 7.328 6.568 ;
  LAYER M1 ;
        RECT 7.36 4.08 7.392 6.588 ;
  LAYER M3 ;
        RECT 7.36 4.1 7.392 4.132 ;
  LAYER M1 ;
        RECT 7.424 4.08 7.456 6.588 ;
  LAYER M3 ;
        RECT 7.424 6.536 7.456 6.568 ;
  LAYER M1 ;
        RECT 7.488 4.08 7.52 6.588 ;
  LAYER M3 ;
        RECT 7.488 4.1 7.52 4.132 ;
  LAYER M1 ;
        RECT 7.552 4.08 7.584 6.588 ;
  LAYER M3 ;
        RECT 7.552 6.536 7.584 6.568 ;
  LAYER M1 ;
        RECT 7.616 4.08 7.648 6.588 ;
  LAYER M3 ;
        RECT 7.616 4.1 7.648 4.132 ;
  LAYER M1 ;
        RECT 7.68 4.08 7.712 6.588 ;
  LAYER M3 ;
        RECT 7.68 6.536 7.712 6.568 ;
  LAYER M1 ;
        RECT 7.744 4.08 7.776 6.588 ;
  LAYER M3 ;
        RECT 7.744 4.1 7.776 4.132 ;
  LAYER M1 ;
        RECT 7.808 4.08 7.84 6.588 ;
  LAYER M3 ;
        RECT 7.808 6.536 7.84 6.568 ;
  LAYER M1 ;
        RECT 7.872 4.08 7.904 6.588 ;
  LAYER M3 ;
        RECT 7.872 4.1 7.904 4.132 ;
  LAYER M1 ;
        RECT 7.936 4.08 7.968 6.588 ;
  LAYER M3 ;
        RECT 7.936 6.536 7.968 6.568 ;
  LAYER M1 ;
        RECT 8 4.08 8.032 6.588 ;
  LAYER M3 ;
        RECT 8 4.1 8.032 4.132 ;
  LAYER M1 ;
        RECT 8.064 4.08 8.096 6.588 ;
  LAYER M3 ;
        RECT 8.064 6.536 8.096 6.568 ;
  LAYER M1 ;
        RECT 8.128 4.08 8.16 6.588 ;
  LAYER M3 ;
        RECT 8.128 4.1 8.16 4.132 ;
  LAYER M1 ;
        RECT 8.192 4.08 8.224 6.588 ;
  LAYER M3 ;
        RECT 8.192 6.536 8.224 6.568 ;
  LAYER M1 ;
        RECT 8.256 4.08 8.288 6.588 ;
  LAYER M3 ;
        RECT 8.256 4.1 8.288 4.132 ;
  LAYER M1 ;
        RECT 8.32 4.08 8.352 6.588 ;
  LAYER M3 ;
        RECT 8.32 6.536 8.352 6.568 ;
  LAYER M1 ;
        RECT 8.384 4.08 8.416 6.588 ;
  LAYER M3 ;
        RECT 8.384 4.1 8.416 4.132 ;
  LAYER M1 ;
        RECT 8.448 4.08 8.48 6.588 ;
  LAYER M3 ;
        RECT 8.448 6.536 8.48 6.568 ;
  LAYER M1 ;
        RECT 8.512 4.08 8.544 6.588 ;
  LAYER M3 ;
        RECT 8.512 4.1 8.544 4.132 ;
  LAYER M1 ;
        RECT 8.576 4.08 8.608 6.588 ;
  LAYER M3 ;
        RECT 8.576 6.536 8.608 6.568 ;
  LAYER M1 ;
        RECT 8.64 4.08 8.672 6.588 ;
  LAYER M3 ;
        RECT 8.64 4.1 8.672 4.132 ;
  LAYER M1 ;
        RECT 8.704 4.08 8.736 6.588 ;
  LAYER M3 ;
        RECT 8.704 6.536 8.736 6.568 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 6.588 ;
  LAYER M3 ;
        RECT 6.4 4.164 6.432 4.196 ;
  LAYER M2 ;
        RECT 8.768 4.228 8.8 4.26 ;
  LAYER M2 ;
        RECT 6.4 4.292 6.432 4.324 ;
  LAYER M2 ;
        RECT 8.768 4.356 8.8 4.388 ;
  LAYER M2 ;
        RECT 6.4 4.42 6.432 4.452 ;
  LAYER M2 ;
        RECT 8.768 4.484 8.8 4.516 ;
  LAYER M2 ;
        RECT 6.4 4.548 6.432 4.58 ;
  LAYER M2 ;
        RECT 8.768 4.612 8.8 4.644 ;
  LAYER M2 ;
        RECT 6.4 4.676 6.432 4.708 ;
  LAYER M2 ;
        RECT 8.768 4.74 8.8 4.772 ;
  LAYER M2 ;
        RECT 6.4 4.804 6.432 4.836 ;
  LAYER M2 ;
        RECT 8.768 4.868 8.8 4.9 ;
  LAYER M2 ;
        RECT 6.4 4.932 6.432 4.964 ;
  LAYER M2 ;
        RECT 8.768 4.996 8.8 5.028 ;
  LAYER M2 ;
        RECT 6.4 5.06 6.432 5.092 ;
  LAYER M2 ;
        RECT 8.768 5.124 8.8 5.156 ;
  LAYER M2 ;
        RECT 6.4 5.188 6.432 5.22 ;
  LAYER M2 ;
        RECT 8.768 5.252 8.8 5.284 ;
  LAYER M2 ;
        RECT 6.4 5.316 6.432 5.348 ;
  LAYER M2 ;
        RECT 8.768 5.38 8.8 5.412 ;
  LAYER M2 ;
        RECT 6.4 5.444 6.432 5.476 ;
  LAYER M2 ;
        RECT 8.768 5.508 8.8 5.54 ;
  LAYER M2 ;
        RECT 6.4 5.572 6.432 5.604 ;
  LAYER M2 ;
        RECT 8.768 5.636 8.8 5.668 ;
  LAYER M2 ;
        RECT 6.4 5.7 6.432 5.732 ;
  LAYER M2 ;
        RECT 8.768 5.764 8.8 5.796 ;
  LAYER M2 ;
        RECT 6.4 5.828 6.432 5.86 ;
  LAYER M2 ;
        RECT 8.768 5.892 8.8 5.924 ;
  LAYER M2 ;
        RECT 6.4 5.956 6.432 5.988 ;
  LAYER M2 ;
        RECT 8.768 6.02 8.8 6.052 ;
  LAYER M2 ;
        RECT 6.4 6.084 6.432 6.116 ;
  LAYER M2 ;
        RECT 8.768 6.148 8.8 6.18 ;
  LAYER M2 ;
        RECT 6.4 6.212 6.432 6.244 ;
  LAYER M2 ;
        RECT 8.768 6.276 8.8 6.308 ;
  LAYER M2 ;
        RECT 6.4 6.34 6.432 6.372 ;
  LAYER M2 ;
        RECT 8.768 6.404 8.8 6.436 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.4 7.188 6.432 9.696 ;
  LAYER M3 ;
        RECT 6.4 9.644 6.432 9.676 ;
  LAYER M1 ;
        RECT 6.464 7.188 6.496 9.696 ;
  LAYER M3 ;
        RECT 6.464 7.208 6.496 7.24 ;
  LAYER M1 ;
        RECT 6.528 7.188 6.56 9.696 ;
  LAYER M3 ;
        RECT 6.528 9.644 6.56 9.676 ;
  LAYER M1 ;
        RECT 6.592 7.188 6.624 9.696 ;
  LAYER M3 ;
        RECT 6.592 7.208 6.624 7.24 ;
  LAYER M1 ;
        RECT 6.656 7.188 6.688 9.696 ;
  LAYER M3 ;
        RECT 6.656 9.644 6.688 9.676 ;
  LAYER M1 ;
        RECT 6.72 7.188 6.752 9.696 ;
  LAYER M3 ;
        RECT 6.72 7.208 6.752 7.24 ;
  LAYER M1 ;
        RECT 6.784 7.188 6.816 9.696 ;
  LAYER M3 ;
        RECT 6.784 9.644 6.816 9.676 ;
  LAYER M1 ;
        RECT 6.848 7.188 6.88 9.696 ;
  LAYER M3 ;
        RECT 6.848 7.208 6.88 7.24 ;
  LAYER M1 ;
        RECT 6.912 7.188 6.944 9.696 ;
  LAYER M3 ;
        RECT 6.912 9.644 6.944 9.676 ;
  LAYER M1 ;
        RECT 6.976 7.188 7.008 9.696 ;
  LAYER M3 ;
        RECT 6.976 7.208 7.008 7.24 ;
  LAYER M1 ;
        RECT 7.04 7.188 7.072 9.696 ;
  LAYER M3 ;
        RECT 7.04 9.644 7.072 9.676 ;
  LAYER M1 ;
        RECT 7.104 7.188 7.136 9.696 ;
  LAYER M3 ;
        RECT 7.104 7.208 7.136 7.24 ;
  LAYER M1 ;
        RECT 7.168 7.188 7.2 9.696 ;
  LAYER M3 ;
        RECT 7.168 9.644 7.2 9.676 ;
  LAYER M1 ;
        RECT 7.232 7.188 7.264 9.696 ;
  LAYER M3 ;
        RECT 7.232 7.208 7.264 7.24 ;
  LAYER M1 ;
        RECT 7.296 7.188 7.328 9.696 ;
  LAYER M3 ;
        RECT 7.296 9.644 7.328 9.676 ;
  LAYER M1 ;
        RECT 7.36 7.188 7.392 9.696 ;
  LAYER M3 ;
        RECT 7.36 7.208 7.392 7.24 ;
  LAYER M1 ;
        RECT 7.424 7.188 7.456 9.696 ;
  LAYER M3 ;
        RECT 7.424 9.644 7.456 9.676 ;
  LAYER M1 ;
        RECT 7.488 7.188 7.52 9.696 ;
  LAYER M3 ;
        RECT 7.488 7.208 7.52 7.24 ;
  LAYER M1 ;
        RECT 7.552 7.188 7.584 9.696 ;
  LAYER M3 ;
        RECT 7.552 9.644 7.584 9.676 ;
  LAYER M1 ;
        RECT 7.616 7.188 7.648 9.696 ;
  LAYER M3 ;
        RECT 7.616 7.208 7.648 7.24 ;
  LAYER M1 ;
        RECT 7.68 7.188 7.712 9.696 ;
  LAYER M3 ;
        RECT 7.68 9.644 7.712 9.676 ;
  LAYER M1 ;
        RECT 7.744 7.188 7.776 9.696 ;
  LAYER M3 ;
        RECT 7.744 7.208 7.776 7.24 ;
  LAYER M1 ;
        RECT 7.808 7.188 7.84 9.696 ;
  LAYER M3 ;
        RECT 7.808 9.644 7.84 9.676 ;
  LAYER M1 ;
        RECT 7.872 7.188 7.904 9.696 ;
  LAYER M3 ;
        RECT 7.872 7.208 7.904 7.24 ;
  LAYER M1 ;
        RECT 7.936 7.188 7.968 9.696 ;
  LAYER M3 ;
        RECT 7.936 9.644 7.968 9.676 ;
  LAYER M1 ;
        RECT 8 7.188 8.032 9.696 ;
  LAYER M3 ;
        RECT 8 7.208 8.032 7.24 ;
  LAYER M1 ;
        RECT 8.064 7.188 8.096 9.696 ;
  LAYER M3 ;
        RECT 8.064 9.644 8.096 9.676 ;
  LAYER M1 ;
        RECT 8.128 7.188 8.16 9.696 ;
  LAYER M3 ;
        RECT 8.128 7.208 8.16 7.24 ;
  LAYER M1 ;
        RECT 8.192 7.188 8.224 9.696 ;
  LAYER M3 ;
        RECT 8.192 9.644 8.224 9.676 ;
  LAYER M1 ;
        RECT 8.256 7.188 8.288 9.696 ;
  LAYER M3 ;
        RECT 8.256 7.208 8.288 7.24 ;
  LAYER M1 ;
        RECT 8.32 7.188 8.352 9.696 ;
  LAYER M3 ;
        RECT 8.32 9.644 8.352 9.676 ;
  LAYER M1 ;
        RECT 8.384 7.188 8.416 9.696 ;
  LAYER M3 ;
        RECT 8.384 7.208 8.416 7.24 ;
  LAYER M1 ;
        RECT 8.448 7.188 8.48 9.696 ;
  LAYER M3 ;
        RECT 8.448 9.644 8.48 9.676 ;
  LAYER M1 ;
        RECT 8.512 7.188 8.544 9.696 ;
  LAYER M3 ;
        RECT 8.512 7.208 8.544 7.24 ;
  LAYER M1 ;
        RECT 8.576 7.188 8.608 9.696 ;
  LAYER M3 ;
        RECT 8.576 9.644 8.608 9.676 ;
  LAYER M1 ;
        RECT 8.64 7.188 8.672 9.696 ;
  LAYER M3 ;
        RECT 8.64 7.208 8.672 7.24 ;
  LAYER M1 ;
        RECT 8.704 7.188 8.736 9.696 ;
  LAYER M3 ;
        RECT 8.704 9.644 8.736 9.676 ;
  LAYER M1 ;
        RECT 8.768 7.188 8.8 9.696 ;
  LAYER M3 ;
        RECT 6.4 7.272 6.432 7.304 ;
  LAYER M2 ;
        RECT 8.768 7.336 8.8 7.368 ;
  LAYER M2 ;
        RECT 6.4 7.4 6.432 7.432 ;
  LAYER M2 ;
        RECT 8.768 7.464 8.8 7.496 ;
  LAYER M2 ;
        RECT 6.4 7.528 6.432 7.56 ;
  LAYER M2 ;
        RECT 8.768 7.592 8.8 7.624 ;
  LAYER M2 ;
        RECT 6.4 7.656 6.432 7.688 ;
  LAYER M2 ;
        RECT 8.768 7.72 8.8 7.752 ;
  LAYER M2 ;
        RECT 6.4 7.784 6.432 7.816 ;
  LAYER M2 ;
        RECT 8.768 7.848 8.8 7.88 ;
  LAYER M2 ;
        RECT 6.4 7.912 6.432 7.944 ;
  LAYER M2 ;
        RECT 8.768 7.976 8.8 8.008 ;
  LAYER M2 ;
        RECT 6.4 8.04 6.432 8.072 ;
  LAYER M2 ;
        RECT 8.768 8.104 8.8 8.136 ;
  LAYER M2 ;
        RECT 6.4 8.168 6.432 8.2 ;
  LAYER M2 ;
        RECT 8.768 8.232 8.8 8.264 ;
  LAYER M2 ;
        RECT 6.4 8.296 6.432 8.328 ;
  LAYER M2 ;
        RECT 8.768 8.36 8.8 8.392 ;
  LAYER M2 ;
        RECT 6.4 8.424 6.432 8.456 ;
  LAYER M2 ;
        RECT 8.768 8.488 8.8 8.52 ;
  LAYER M2 ;
        RECT 6.4 8.552 6.432 8.584 ;
  LAYER M2 ;
        RECT 8.768 8.616 8.8 8.648 ;
  LAYER M2 ;
        RECT 6.4 8.68 6.432 8.712 ;
  LAYER M2 ;
        RECT 8.768 8.744 8.8 8.776 ;
  LAYER M2 ;
        RECT 6.4 8.808 6.432 8.84 ;
  LAYER M2 ;
        RECT 8.768 8.872 8.8 8.904 ;
  LAYER M2 ;
        RECT 6.4 8.936 6.432 8.968 ;
  LAYER M2 ;
        RECT 8.768 9 8.8 9.032 ;
  LAYER M2 ;
        RECT 6.4 9.064 6.432 9.096 ;
  LAYER M2 ;
        RECT 8.768 9.128 8.8 9.16 ;
  LAYER M2 ;
        RECT 6.4 9.192 6.432 9.224 ;
  LAYER M2 ;
        RECT 8.768 9.256 8.8 9.288 ;
  LAYER M2 ;
        RECT 6.4 9.32 6.432 9.352 ;
  LAYER M2 ;
        RECT 8.768 9.384 8.8 9.416 ;
  LAYER M2 ;
        RECT 6.4 9.448 6.432 9.48 ;
  LAYER M2 ;
        RECT 8.768 9.512 8.8 9.544 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.4 10.296 6.432 12.804 ;
  LAYER M3 ;
        RECT 6.4 12.752 6.432 12.784 ;
  LAYER M1 ;
        RECT 6.464 10.296 6.496 12.804 ;
  LAYER M3 ;
        RECT 6.464 10.316 6.496 10.348 ;
  LAYER M1 ;
        RECT 6.528 10.296 6.56 12.804 ;
  LAYER M3 ;
        RECT 6.528 12.752 6.56 12.784 ;
  LAYER M1 ;
        RECT 6.592 10.296 6.624 12.804 ;
  LAYER M3 ;
        RECT 6.592 10.316 6.624 10.348 ;
  LAYER M1 ;
        RECT 6.656 10.296 6.688 12.804 ;
  LAYER M3 ;
        RECT 6.656 12.752 6.688 12.784 ;
  LAYER M1 ;
        RECT 6.72 10.296 6.752 12.804 ;
  LAYER M3 ;
        RECT 6.72 10.316 6.752 10.348 ;
  LAYER M1 ;
        RECT 6.784 10.296 6.816 12.804 ;
  LAYER M3 ;
        RECT 6.784 12.752 6.816 12.784 ;
  LAYER M1 ;
        RECT 6.848 10.296 6.88 12.804 ;
  LAYER M3 ;
        RECT 6.848 10.316 6.88 10.348 ;
  LAYER M1 ;
        RECT 6.912 10.296 6.944 12.804 ;
  LAYER M3 ;
        RECT 6.912 12.752 6.944 12.784 ;
  LAYER M1 ;
        RECT 6.976 10.296 7.008 12.804 ;
  LAYER M3 ;
        RECT 6.976 10.316 7.008 10.348 ;
  LAYER M1 ;
        RECT 7.04 10.296 7.072 12.804 ;
  LAYER M3 ;
        RECT 7.04 12.752 7.072 12.784 ;
  LAYER M1 ;
        RECT 7.104 10.296 7.136 12.804 ;
  LAYER M3 ;
        RECT 7.104 10.316 7.136 10.348 ;
  LAYER M1 ;
        RECT 7.168 10.296 7.2 12.804 ;
  LAYER M3 ;
        RECT 7.168 12.752 7.2 12.784 ;
  LAYER M1 ;
        RECT 7.232 10.296 7.264 12.804 ;
  LAYER M3 ;
        RECT 7.232 10.316 7.264 10.348 ;
  LAYER M1 ;
        RECT 7.296 10.296 7.328 12.804 ;
  LAYER M3 ;
        RECT 7.296 12.752 7.328 12.784 ;
  LAYER M1 ;
        RECT 7.36 10.296 7.392 12.804 ;
  LAYER M3 ;
        RECT 7.36 10.316 7.392 10.348 ;
  LAYER M1 ;
        RECT 7.424 10.296 7.456 12.804 ;
  LAYER M3 ;
        RECT 7.424 12.752 7.456 12.784 ;
  LAYER M1 ;
        RECT 7.488 10.296 7.52 12.804 ;
  LAYER M3 ;
        RECT 7.488 10.316 7.52 10.348 ;
  LAYER M1 ;
        RECT 7.552 10.296 7.584 12.804 ;
  LAYER M3 ;
        RECT 7.552 12.752 7.584 12.784 ;
  LAYER M1 ;
        RECT 7.616 10.296 7.648 12.804 ;
  LAYER M3 ;
        RECT 7.616 10.316 7.648 10.348 ;
  LAYER M1 ;
        RECT 7.68 10.296 7.712 12.804 ;
  LAYER M3 ;
        RECT 7.68 12.752 7.712 12.784 ;
  LAYER M1 ;
        RECT 7.744 10.296 7.776 12.804 ;
  LAYER M3 ;
        RECT 7.744 10.316 7.776 10.348 ;
  LAYER M1 ;
        RECT 7.808 10.296 7.84 12.804 ;
  LAYER M3 ;
        RECT 7.808 12.752 7.84 12.784 ;
  LAYER M1 ;
        RECT 7.872 10.296 7.904 12.804 ;
  LAYER M3 ;
        RECT 7.872 10.316 7.904 10.348 ;
  LAYER M1 ;
        RECT 7.936 10.296 7.968 12.804 ;
  LAYER M3 ;
        RECT 7.936 12.752 7.968 12.784 ;
  LAYER M1 ;
        RECT 8 10.296 8.032 12.804 ;
  LAYER M3 ;
        RECT 8 10.316 8.032 10.348 ;
  LAYER M1 ;
        RECT 8.064 10.296 8.096 12.804 ;
  LAYER M3 ;
        RECT 8.064 12.752 8.096 12.784 ;
  LAYER M1 ;
        RECT 8.128 10.296 8.16 12.804 ;
  LAYER M3 ;
        RECT 8.128 10.316 8.16 10.348 ;
  LAYER M1 ;
        RECT 8.192 10.296 8.224 12.804 ;
  LAYER M3 ;
        RECT 8.192 12.752 8.224 12.784 ;
  LAYER M1 ;
        RECT 8.256 10.296 8.288 12.804 ;
  LAYER M3 ;
        RECT 8.256 10.316 8.288 10.348 ;
  LAYER M1 ;
        RECT 8.32 10.296 8.352 12.804 ;
  LAYER M3 ;
        RECT 8.32 12.752 8.352 12.784 ;
  LAYER M1 ;
        RECT 8.384 10.296 8.416 12.804 ;
  LAYER M3 ;
        RECT 8.384 10.316 8.416 10.348 ;
  LAYER M1 ;
        RECT 8.448 10.296 8.48 12.804 ;
  LAYER M3 ;
        RECT 8.448 12.752 8.48 12.784 ;
  LAYER M1 ;
        RECT 8.512 10.296 8.544 12.804 ;
  LAYER M3 ;
        RECT 8.512 10.316 8.544 10.348 ;
  LAYER M1 ;
        RECT 8.576 10.296 8.608 12.804 ;
  LAYER M3 ;
        RECT 8.576 12.752 8.608 12.784 ;
  LAYER M1 ;
        RECT 8.64 10.296 8.672 12.804 ;
  LAYER M3 ;
        RECT 8.64 10.316 8.672 10.348 ;
  LAYER M1 ;
        RECT 8.704 10.296 8.736 12.804 ;
  LAYER M3 ;
        RECT 8.704 12.752 8.736 12.784 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 12.804 ;
  LAYER M3 ;
        RECT 6.4 10.38 6.432 10.412 ;
  LAYER M2 ;
        RECT 8.768 10.444 8.8 10.476 ;
  LAYER M2 ;
        RECT 6.4 10.508 6.432 10.54 ;
  LAYER M2 ;
        RECT 8.768 10.572 8.8 10.604 ;
  LAYER M2 ;
        RECT 6.4 10.636 6.432 10.668 ;
  LAYER M2 ;
        RECT 8.768 10.7 8.8 10.732 ;
  LAYER M2 ;
        RECT 6.4 10.764 6.432 10.796 ;
  LAYER M2 ;
        RECT 8.768 10.828 8.8 10.86 ;
  LAYER M2 ;
        RECT 6.4 10.892 6.432 10.924 ;
  LAYER M2 ;
        RECT 8.768 10.956 8.8 10.988 ;
  LAYER M2 ;
        RECT 6.4 11.02 6.432 11.052 ;
  LAYER M2 ;
        RECT 8.768 11.084 8.8 11.116 ;
  LAYER M2 ;
        RECT 6.4 11.148 6.432 11.18 ;
  LAYER M2 ;
        RECT 8.768 11.212 8.8 11.244 ;
  LAYER M2 ;
        RECT 6.4 11.276 6.432 11.308 ;
  LAYER M2 ;
        RECT 8.768 11.34 8.8 11.372 ;
  LAYER M2 ;
        RECT 6.4 11.404 6.432 11.436 ;
  LAYER M2 ;
        RECT 8.768 11.468 8.8 11.5 ;
  LAYER M2 ;
        RECT 6.4 11.532 6.432 11.564 ;
  LAYER M2 ;
        RECT 8.768 11.596 8.8 11.628 ;
  LAYER M2 ;
        RECT 6.4 11.66 6.432 11.692 ;
  LAYER M2 ;
        RECT 8.768 11.724 8.8 11.756 ;
  LAYER M2 ;
        RECT 6.4 11.788 6.432 11.82 ;
  LAYER M2 ;
        RECT 8.768 11.852 8.8 11.884 ;
  LAYER M2 ;
        RECT 6.4 11.916 6.432 11.948 ;
  LAYER M2 ;
        RECT 8.768 11.98 8.8 12.012 ;
  LAYER M2 ;
        RECT 6.4 12.044 6.432 12.076 ;
  LAYER M2 ;
        RECT 8.768 12.108 8.8 12.14 ;
  LAYER M2 ;
        RECT 6.4 12.172 6.432 12.204 ;
  LAYER M2 ;
        RECT 8.768 12.236 8.8 12.268 ;
  LAYER M2 ;
        RECT 6.4 12.3 6.432 12.332 ;
  LAYER M2 ;
        RECT 8.768 12.364 8.8 12.396 ;
  LAYER M2 ;
        RECT 6.4 12.428 6.432 12.46 ;
  LAYER M2 ;
        RECT 8.768 12.492 8.8 12.524 ;
  LAYER M2 ;
        RECT 6.4 12.556 6.432 12.588 ;
  LAYER M2 ;
        RECT 8.768 12.62 8.8 12.652 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 6.4 13.404 6.432 15.912 ;
  LAYER M3 ;
        RECT 6.4 15.86 6.432 15.892 ;
  LAYER M1 ;
        RECT 6.464 13.404 6.496 15.912 ;
  LAYER M3 ;
        RECT 6.464 13.424 6.496 13.456 ;
  LAYER M1 ;
        RECT 6.528 13.404 6.56 15.912 ;
  LAYER M3 ;
        RECT 6.528 15.86 6.56 15.892 ;
  LAYER M1 ;
        RECT 6.592 13.404 6.624 15.912 ;
  LAYER M3 ;
        RECT 6.592 13.424 6.624 13.456 ;
  LAYER M1 ;
        RECT 6.656 13.404 6.688 15.912 ;
  LAYER M3 ;
        RECT 6.656 15.86 6.688 15.892 ;
  LAYER M1 ;
        RECT 6.72 13.404 6.752 15.912 ;
  LAYER M3 ;
        RECT 6.72 13.424 6.752 13.456 ;
  LAYER M1 ;
        RECT 6.784 13.404 6.816 15.912 ;
  LAYER M3 ;
        RECT 6.784 15.86 6.816 15.892 ;
  LAYER M1 ;
        RECT 6.848 13.404 6.88 15.912 ;
  LAYER M3 ;
        RECT 6.848 13.424 6.88 13.456 ;
  LAYER M1 ;
        RECT 6.912 13.404 6.944 15.912 ;
  LAYER M3 ;
        RECT 6.912 15.86 6.944 15.892 ;
  LAYER M1 ;
        RECT 6.976 13.404 7.008 15.912 ;
  LAYER M3 ;
        RECT 6.976 13.424 7.008 13.456 ;
  LAYER M1 ;
        RECT 7.04 13.404 7.072 15.912 ;
  LAYER M3 ;
        RECT 7.04 15.86 7.072 15.892 ;
  LAYER M1 ;
        RECT 7.104 13.404 7.136 15.912 ;
  LAYER M3 ;
        RECT 7.104 13.424 7.136 13.456 ;
  LAYER M1 ;
        RECT 7.168 13.404 7.2 15.912 ;
  LAYER M3 ;
        RECT 7.168 15.86 7.2 15.892 ;
  LAYER M1 ;
        RECT 7.232 13.404 7.264 15.912 ;
  LAYER M3 ;
        RECT 7.232 13.424 7.264 13.456 ;
  LAYER M1 ;
        RECT 7.296 13.404 7.328 15.912 ;
  LAYER M3 ;
        RECT 7.296 15.86 7.328 15.892 ;
  LAYER M1 ;
        RECT 7.36 13.404 7.392 15.912 ;
  LAYER M3 ;
        RECT 7.36 13.424 7.392 13.456 ;
  LAYER M1 ;
        RECT 7.424 13.404 7.456 15.912 ;
  LAYER M3 ;
        RECT 7.424 15.86 7.456 15.892 ;
  LAYER M1 ;
        RECT 7.488 13.404 7.52 15.912 ;
  LAYER M3 ;
        RECT 7.488 13.424 7.52 13.456 ;
  LAYER M1 ;
        RECT 7.552 13.404 7.584 15.912 ;
  LAYER M3 ;
        RECT 7.552 15.86 7.584 15.892 ;
  LAYER M1 ;
        RECT 7.616 13.404 7.648 15.912 ;
  LAYER M3 ;
        RECT 7.616 13.424 7.648 13.456 ;
  LAYER M1 ;
        RECT 7.68 13.404 7.712 15.912 ;
  LAYER M3 ;
        RECT 7.68 15.86 7.712 15.892 ;
  LAYER M1 ;
        RECT 7.744 13.404 7.776 15.912 ;
  LAYER M3 ;
        RECT 7.744 13.424 7.776 13.456 ;
  LAYER M1 ;
        RECT 7.808 13.404 7.84 15.912 ;
  LAYER M3 ;
        RECT 7.808 15.86 7.84 15.892 ;
  LAYER M1 ;
        RECT 7.872 13.404 7.904 15.912 ;
  LAYER M3 ;
        RECT 7.872 13.424 7.904 13.456 ;
  LAYER M1 ;
        RECT 7.936 13.404 7.968 15.912 ;
  LAYER M3 ;
        RECT 7.936 15.86 7.968 15.892 ;
  LAYER M1 ;
        RECT 8 13.404 8.032 15.912 ;
  LAYER M3 ;
        RECT 8 13.424 8.032 13.456 ;
  LAYER M1 ;
        RECT 8.064 13.404 8.096 15.912 ;
  LAYER M3 ;
        RECT 8.064 15.86 8.096 15.892 ;
  LAYER M1 ;
        RECT 8.128 13.404 8.16 15.912 ;
  LAYER M3 ;
        RECT 8.128 13.424 8.16 13.456 ;
  LAYER M1 ;
        RECT 8.192 13.404 8.224 15.912 ;
  LAYER M3 ;
        RECT 8.192 15.86 8.224 15.892 ;
  LAYER M1 ;
        RECT 8.256 13.404 8.288 15.912 ;
  LAYER M3 ;
        RECT 8.256 13.424 8.288 13.456 ;
  LAYER M1 ;
        RECT 8.32 13.404 8.352 15.912 ;
  LAYER M3 ;
        RECT 8.32 15.86 8.352 15.892 ;
  LAYER M1 ;
        RECT 8.384 13.404 8.416 15.912 ;
  LAYER M3 ;
        RECT 8.384 13.424 8.416 13.456 ;
  LAYER M1 ;
        RECT 8.448 13.404 8.48 15.912 ;
  LAYER M3 ;
        RECT 8.448 15.86 8.48 15.892 ;
  LAYER M1 ;
        RECT 8.512 13.404 8.544 15.912 ;
  LAYER M3 ;
        RECT 8.512 13.424 8.544 13.456 ;
  LAYER M1 ;
        RECT 8.576 13.404 8.608 15.912 ;
  LAYER M3 ;
        RECT 8.576 15.86 8.608 15.892 ;
  LAYER M1 ;
        RECT 8.64 13.404 8.672 15.912 ;
  LAYER M3 ;
        RECT 8.64 13.424 8.672 13.456 ;
  LAYER M1 ;
        RECT 8.704 13.404 8.736 15.912 ;
  LAYER M3 ;
        RECT 8.704 15.86 8.736 15.892 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 15.912 ;
  LAYER M3 ;
        RECT 6.4 13.488 6.432 13.52 ;
  LAYER M2 ;
        RECT 8.768 13.552 8.8 13.584 ;
  LAYER M2 ;
        RECT 6.4 13.616 6.432 13.648 ;
  LAYER M2 ;
        RECT 8.768 13.68 8.8 13.712 ;
  LAYER M2 ;
        RECT 6.4 13.744 6.432 13.776 ;
  LAYER M2 ;
        RECT 8.768 13.808 8.8 13.84 ;
  LAYER M2 ;
        RECT 6.4 13.872 6.432 13.904 ;
  LAYER M2 ;
        RECT 8.768 13.936 8.8 13.968 ;
  LAYER M2 ;
        RECT 6.4 14 6.432 14.032 ;
  LAYER M2 ;
        RECT 8.768 14.064 8.8 14.096 ;
  LAYER M2 ;
        RECT 6.4 14.128 6.432 14.16 ;
  LAYER M2 ;
        RECT 8.768 14.192 8.8 14.224 ;
  LAYER M2 ;
        RECT 6.4 14.256 6.432 14.288 ;
  LAYER M2 ;
        RECT 8.768 14.32 8.8 14.352 ;
  LAYER M2 ;
        RECT 6.4 14.384 6.432 14.416 ;
  LAYER M2 ;
        RECT 8.768 14.448 8.8 14.48 ;
  LAYER M2 ;
        RECT 6.4 14.512 6.432 14.544 ;
  LAYER M2 ;
        RECT 8.768 14.576 8.8 14.608 ;
  LAYER M2 ;
        RECT 6.4 14.64 6.432 14.672 ;
  LAYER M2 ;
        RECT 8.768 14.704 8.8 14.736 ;
  LAYER M2 ;
        RECT 6.4 14.768 6.432 14.8 ;
  LAYER M2 ;
        RECT 8.768 14.832 8.8 14.864 ;
  LAYER M2 ;
        RECT 6.4 14.896 6.432 14.928 ;
  LAYER M2 ;
        RECT 8.768 14.96 8.8 14.992 ;
  LAYER M2 ;
        RECT 6.4 15.024 6.432 15.056 ;
  LAYER M2 ;
        RECT 8.768 15.088 8.8 15.12 ;
  LAYER M2 ;
        RECT 6.4 15.152 6.432 15.184 ;
  LAYER M2 ;
        RECT 8.768 15.216 8.8 15.248 ;
  LAYER M2 ;
        RECT 6.4 15.28 6.432 15.312 ;
  LAYER M2 ;
        RECT 8.768 15.344 8.8 15.376 ;
  LAYER M2 ;
        RECT 6.4 15.408 6.432 15.44 ;
  LAYER M2 ;
        RECT 8.768 15.472 8.8 15.504 ;
  LAYER M2 ;
        RECT 6.4 15.536 6.432 15.568 ;
  LAYER M2 ;
        RECT 8.768 15.6 8.8 15.632 ;
  LAYER M2 ;
        RECT 6.4 15.664 6.432 15.696 ;
  LAYER M2 ;
        RECT 8.768 15.728 8.8 15.76 ;
  LAYER M2 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M1 ;
        RECT 9.376 0.972 9.408 3.48 ;
  LAYER M3 ;
        RECT 9.376 3.428 9.408 3.46 ;
  LAYER M1 ;
        RECT 9.44 0.972 9.472 3.48 ;
  LAYER M3 ;
        RECT 9.44 0.992 9.472 1.024 ;
  LAYER M1 ;
        RECT 9.504 0.972 9.536 3.48 ;
  LAYER M3 ;
        RECT 9.504 3.428 9.536 3.46 ;
  LAYER M1 ;
        RECT 9.568 0.972 9.6 3.48 ;
  LAYER M3 ;
        RECT 9.568 0.992 9.6 1.024 ;
  LAYER M1 ;
        RECT 9.632 0.972 9.664 3.48 ;
  LAYER M3 ;
        RECT 9.632 3.428 9.664 3.46 ;
  LAYER M1 ;
        RECT 9.696 0.972 9.728 3.48 ;
  LAYER M3 ;
        RECT 9.696 0.992 9.728 1.024 ;
  LAYER M1 ;
        RECT 9.76 0.972 9.792 3.48 ;
  LAYER M3 ;
        RECT 9.76 3.428 9.792 3.46 ;
  LAYER M1 ;
        RECT 9.824 0.972 9.856 3.48 ;
  LAYER M3 ;
        RECT 9.824 0.992 9.856 1.024 ;
  LAYER M1 ;
        RECT 9.888 0.972 9.92 3.48 ;
  LAYER M3 ;
        RECT 9.888 3.428 9.92 3.46 ;
  LAYER M1 ;
        RECT 9.952 0.972 9.984 3.48 ;
  LAYER M3 ;
        RECT 9.952 0.992 9.984 1.024 ;
  LAYER M1 ;
        RECT 10.016 0.972 10.048 3.48 ;
  LAYER M3 ;
        RECT 10.016 3.428 10.048 3.46 ;
  LAYER M1 ;
        RECT 10.08 0.972 10.112 3.48 ;
  LAYER M3 ;
        RECT 10.08 0.992 10.112 1.024 ;
  LAYER M1 ;
        RECT 10.144 0.972 10.176 3.48 ;
  LAYER M3 ;
        RECT 10.144 3.428 10.176 3.46 ;
  LAYER M1 ;
        RECT 10.208 0.972 10.24 3.48 ;
  LAYER M3 ;
        RECT 10.208 0.992 10.24 1.024 ;
  LAYER M1 ;
        RECT 10.272 0.972 10.304 3.48 ;
  LAYER M3 ;
        RECT 10.272 3.428 10.304 3.46 ;
  LAYER M1 ;
        RECT 10.336 0.972 10.368 3.48 ;
  LAYER M3 ;
        RECT 10.336 0.992 10.368 1.024 ;
  LAYER M1 ;
        RECT 10.4 0.972 10.432 3.48 ;
  LAYER M3 ;
        RECT 10.4 3.428 10.432 3.46 ;
  LAYER M1 ;
        RECT 10.464 0.972 10.496 3.48 ;
  LAYER M3 ;
        RECT 10.464 0.992 10.496 1.024 ;
  LAYER M1 ;
        RECT 10.528 0.972 10.56 3.48 ;
  LAYER M3 ;
        RECT 10.528 3.428 10.56 3.46 ;
  LAYER M1 ;
        RECT 10.592 0.972 10.624 3.48 ;
  LAYER M3 ;
        RECT 10.592 0.992 10.624 1.024 ;
  LAYER M1 ;
        RECT 10.656 0.972 10.688 3.48 ;
  LAYER M3 ;
        RECT 10.656 3.428 10.688 3.46 ;
  LAYER M1 ;
        RECT 10.72 0.972 10.752 3.48 ;
  LAYER M3 ;
        RECT 10.72 0.992 10.752 1.024 ;
  LAYER M1 ;
        RECT 10.784 0.972 10.816 3.48 ;
  LAYER M3 ;
        RECT 10.784 3.428 10.816 3.46 ;
  LAYER M1 ;
        RECT 10.848 0.972 10.88 3.48 ;
  LAYER M3 ;
        RECT 10.848 0.992 10.88 1.024 ;
  LAYER M1 ;
        RECT 10.912 0.972 10.944 3.48 ;
  LAYER M3 ;
        RECT 10.912 3.428 10.944 3.46 ;
  LAYER M1 ;
        RECT 10.976 0.972 11.008 3.48 ;
  LAYER M3 ;
        RECT 10.976 0.992 11.008 1.024 ;
  LAYER M1 ;
        RECT 11.04 0.972 11.072 3.48 ;
  LAYER M3 ;
        RECT 11.04 3.428 11.072 3.46 ;
  LAYER M1 ;
        RECT 11.104 0.972 11.136 3.48 ;
  LAYER M3 ;
        RECT 11.104 0.992 11.136 1.024 ;
  LAYER M1 ;
        RECT 11.168 0.972 11.2 3.48 ;
  LAYER M3 ;
        RECT 11.168 3.428 11.2 3.46 ;
  LAYER M1 ;
        RECT 11.232 0.972 11.264 3.48 ;
  LAYER M3 ;
        RECT 11.232 0.992 11.264 1.024 ;
  LAYER M1 ;
        RECT 11.296 0.972 11.328 3.48 ;
  LAYER M3 ;
        RECT 11.296 3.428 11.328 3.46 ;
  LAYER M1 ;
        RECT 11.36 0.972 11.392 3.48 ;
  LAYER M3 ;
        RECT 11.36 0.992 11.392 1.024 ;
  LAYER M1 ;
        RECT 11.424 0.972 11.456 3.48 ;
  LAYER M3 ;
        RECT 11.424 3.428 11.456 3.46 ;
  LAYER M1 ;
        RECT 11.488 0.972 11.52 3.48 ;
  LAYER M3 ;
        RECT 11.488 0.992 11.52 1.024 ;
  LAYER M1 ;
        RECT 11.552 0.972 11.584 3.48 ;
  LAYER M3 ;
        RECT 11.552 3.428 11.584 3.46 ;
  LAYER M1 ;
        RECT 11.616 0.972 11.648 3.48 ;
  LAYER M3 ;
        RECT 11.616 0.992 11.648 1.024 ;
  LAYER M1 ;
        RECT 11.68 0.972 11.712 3.48 ;
  LAYER M3 ;
        RECT 11.68 3.428 11.712 3.46 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 3.48 ;
  LAYER M3 ;
        RECT 9.376 1.056 9.408 1.088 ;
  LAYER M2 ;
        RECT 11.744 1.12 11.776 1.152 ;
  LAYER M2 ;
        RECT 9.376 1.184 9.408 1.216 ;
  LAYER M2 ;
        RECT 11.744 1.248 11.776 1.28 ;
  LAYER M2 ;
        RECT 9.376 1.312 9.408 1.344 ;
  LAYER M2 ;
        RECT 11.744 1.376 11.776 1.408 ;
  LAYER M2 ;
        RECT 9.376 1.44 9.408 1.472 ;
  LAYER M2 ;
        RECT 11.744 1.504 11.776 1.536 ;
  LAYER M2 ;
        RECT 9.376 1.568 9.408 1.6 ;
  LAYER M2 ;
        RECT 11.744 1.632 11.776 1.664 ;
  LAYER M2 ;
        RECT 9.376 1.696 9.408 1.728 ;
  LAYER M2 ;
        RECT 11.744 1.76 11.776 1.792 ;
  LAYER M2 ;
        RECT 9.376 1.824 9.408 1.856 ;
  LAYER M2 ;
        RECT 11.744 1.888 11.776 1.92 ;
  LAYER M2 ;
        RECT 9.376 1.952 9.408 1.984 ;
  LAYER M2 ;
        RECT 11.744 2.016 11.776 2.048 ;
  LAYER M2 ;
        RECT 9.376 2.08 9.408 2.112 ;
  LAYER M2 ;
        RECT 11.744 2.144 11.776 2.176 ;
  LAYER M2 ;
        RECT 9.376 2.208 9.408 2.24 ;
  LAYER M2 ;
        RECT 11.744 2.272 11.776 2.304 ;
  LAYER M2 ;
        RECT 9.376 2.336 9.408 2.368 ;
  LAYER M2 ;
        RECT 11.744 2.4 11.776 2.432 ;
  LAYER M2 ;
        RECT 9.376 2.464 9.408 2.496 ;
  LAYER M2 ;
        RECT 11.744 2.528 11.776 2.56 ;
  LAYER M2 ;
        RECT 9.376 2.592 9.408 2.624 ;
  LAYER M2 ;
        RECT 11.744 2.656 11.776 2.688 ;
  LAYER M2 ;
        RECT 9.376 2.72 9.408 2.752 ;
  LAYER M2 ;
        RECT 11.744 2.784 11.776 2.816 ;
  LAYER M2 ;
        RECT 9.376 2.848 9.408 2.88 ;
  LAYER M2 ;
        RECT 11.744 2.912 11.776 2.944 ;
  LAYER M2 ;
        RECT 9.376 2.976 9.408 3.008 ;
  LAYER M2 ;
        RECT 11.744 3.04 11.776 3.072 ;
  LAYER M2 ;
        RECT 9.376 3.104 9.408 3.136 ;
  LAYER M2 ;
        RECT 11.744 3.168 11.776 3.2 ;
  LAYER M2 ;
        RECT 9.376 3.232 9.408 3.264 ;
  LAYER M2 ;
        RECT 11.744 3.296 11.776 3.328 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.376 4.08 9.408 6.588 ;
  LAYER M3 ;
        RECT 9.376 6.536 9.408 6.568 ;
  LAYER M1 ;
        RECT 9.44 4.08 9.472 6.588 ;
  LAYER M3 ;
        RECT 9.44 4.1 9.472 4.132 ;
  LAYER M1 ;
        RECT 9.504 4.08 9.536 6.588 ;
  LAYER M3 ;
        RECT 9.504 6.536 9.536 6.568 ;
  LAYER M1 ;
        RECT 9.568 4.08 9.6 6.588 ;
  LAYER M3 ;
        RECT 9.568 4.1 9.6 4.132 ;
  LAYER M1 ;
        RECT 9.632 4.08 9.664 6.588 ;
  LAYER M3 ;
        RECT 9.632 6.536 9.664 6.568 ;
  LAYER M1 ;
        RECT 9.696 4.08 9.728 6.588 ;
  LAYER M3 ;
        RECT 9.696 4.1 9.728 4.132 ;
  LAYER M1 ;
        RECT 9.76 4.08 9.792 6.588 ;
  LAYER M3 ;
        RECT 9.76 6.536 9.792 6.568 ;
  LAYER M1 ;
        RECT 9.824 4.08 9.856 6.588 ;
  LAYER M3 ;
        RECT 9.824 4.1 9.856 4.132 ;
  LAYER M1 ;
        RECT 9.888 4.08 9.92 6.588 ;
  LAYER M3 ;
        RECT 9.888 6.536 9.92 6.568 ;
  LAYER M1 ;
        RECT 9.952 4.08 9.984 6.588 ;
  LAYER M3 ;
        RECT 9.952 4.1 9.984 4.132 ;
  LAYER M1 ;
        RECT 10.016 4.08 10.048 6.588 ;
  LAYER M3 ;
        RECT 10.016 6.536 10.048 6.568 ;
  LAYER M1 ;
        RECT 10.08 4.08 10.112 6.588 ;
  LAYER M3 ;
        RECT 10.08 4.1 10.112 4.132 ;
  LAYER M1 ;
        RECT 10.144 4.08 10.176 6.588 ;
  LAYER M3 ;
        RECT 10.144 6.536 10.176 6.568 ;
  LAYER M1 ;
        RECT 10.208 4.08 10.24 6.588 ;
  LAYER M3 ;
        RECT 10.208 4.1 10.24 4.132 ;
  LAYER M1 ;
        RECT 10.272 4.08 10.304 6.588 ;
  LAYER M3 ;
        RECT 10.272 6.536 10.304 6.568 ;
  LAYER M1 ;
        RECT 10.336 4.08 10.368 6.588 ;
  LAYER M3 ;
        RECT 10.336 4.1 10.368 4.132 ;
  LAYER M1 ;
        RECT 10.4 4.08 10.432 6.588 ;
  LAYER M3 ;
        RECT 10.4 6.536 10.432 6.568 ;
  LAYER M1 ;
        RECT 10.464 4.08 10.496 6.588 ;
  LAYER M3 ;
        RECT 10.464 4.1 10.496 4.132 ;
  LAYER M1 ;
        RECT 10.528 4.08 10.56 6.588 ;
  LAYER M3 ;
        RECT 10.528 6.536 10.56 6.568 ;
  LAYER M1 ;
        RECT 10.592 4.08 10.624 6.588 ;
  LAYER M3 ;
        RECT 10.592 4.1 10.624 4.132 ;
  LAYER M1 ;
        RECT 10.656 4.08 10.688 6.588 ;
  LAYER M3 ;
        RECT 10.656 6.536 10.688 6.568 ;
  LAYER M1 ;
        RECT 10.72 4.08 10.752 6.588 ;
  LAYER M3 ;
        RECT 10.72 4.1 10.752 4.132 ;
  LAYER M1 ;
        RECT 10.784 4.08 10.816 6.588 ;
  LAYER M3 ;
        RECT 10.784 6.536 10.816 6.568 ;
  LAYER M1 ;
        RECT 10.848 4.08 10.88 6.588 ;
  LAYER M3 ;
        RECT 10.848 4.1 10.88 4.132 ;
  LAYER M1 ;
        RECT 10.912 4.08 10.944 6.588 ;
  LAYER M3 ;
        RECT 10.912 6.536 10.944 6.568 ;
  LAYER M1 ;
        RECT 10.976 4.08 11.008 6.588 ;
  LAYER M3 ;
        RECT 10.976 4.1 11.008 4.132 ;
  LAYER M1 ;
        RECT 11.04 4.08 11.072 6.588 ;
  LAYER M3 ;
        RECT 11.04 6.536 11.072 6.568 ;
  LAYER M1 ;
        RECT 11.104 4.08 11.136 6.588 ;
  LAYER M3 ;
        RECT 11.104 4.1 11.136 4.132 ;
  LAYER M1 ;
        RECT 11.168 4.08 11.2 6.588 ;
  LAYER M3 ;
        RECT 11.168 6.536 11.2 6.568 ;
  LAYER M1 ;
        RECT 11.232 4.08 11.264 6.588 ;
  LAYER M3 ;
        RECT 11.232 4.1 11.264 4.132 ;
  LAYER M1 ;
        RECT 11.296 4.08 11.328 6.588 ;
  LAYER M3 ;
        RECT 11.296 6.536 11.328 6.568 ;
  LAYER M1 ;
        RECT 11.36 4.08 11.392 6.588 ;
  LAYER M3 ;
        RECT 11.36 4.1 11.392 4.132 ;
  LAYER M1 ;
        RECT 11.424 4.08 11.456 6.588 ;
  LAYER M3 ;
        RECT 11.424 6.536 11.456 6.568 ;
  LAYER M1 ;
        RECT 11.488 4.08 11.52 6.588 ;
  LAYER M3 ;
        RECT 11.488 4.1 11.52 4.132 ;
  LAYER M1 ;
        RECT 11.552 4.08 11.584 6.588 ;
  LAYER M3 ;
        RECT 11.552 6.536 11.584 6.568 ;
  LAYER M1 ;
        RECT 11.616 4.08 11.648 6.588 ;
  LAYER M3 ;
        RECT 11.616 4.1 11.648 4.132 ;
  LAYER M1 ;
        RECT 11.68 4.08 11.712 6.588 ;
  LAYER M3 ;
        RECT 11.68 6.536 11.712 6.568 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 6.588 ;
  LAYER M3 ;
        RECT 9.376 4.164 9.408 4.196 ;
  LAYER M2 ;
        RECT 11.744 4.228 11.776 4.26 ;
  LAYER M2 ;
        RECT 9.376 4.292 9.408 4.324 ;
  LAYER M2 ;
        RECT 11.744 4.356 11.776 4.388 ;
  LAYER M2 ;
        RECT 9.376 4.42 9.408 4.452 ;
  LAYER M2 ;
        RECT 11.744 4.484 11.776 4.516 ;
  LAYER M2 ;
        RECT 9.376 4.548 9.408 4.58 ;
  LAYER M2 ;
        RECT 11.744 4.612 11.776 4.644 ;
  LAYER M2 ;
        RECT 9.376 4.676 9.408 4.708 ;
  LAYER M2 ;
        RECT 11.744 4.74 11.776 4.772 ;
  LAYER M2 ;
        RECT 9.376 4.804 9.408 4.836 ;
  LAYER M2 ;
        RECT 11.744 4.868 11.776 4.9 ;
  LAYER M2 ;
        RECT 9.376 4.932 9.408 4.964 ;
  LAYER M2 ;
        RECT 11.744 4.996 11.776 5.028 ;
  LAYER M2 ;
        RECT 9.376 5.06 9.408 5.092 ;
  LAYER M2 ;
        RECT 11.744 5.124 11.776 5.156 ;
  LAYER M2 ;
        RECT 9.376 5.188 9.408 5.22 ;
  LAYER M2 ;
        RECT 11.744 5.252 11.776 5.284 ;
  LAYER M2 ;
        RECT 9.376 5.316 9.408 5.348 ;
  LAYER M2 ;
        RECT 11.744 5.38 11.776 5.412 ;
  LAYER M2 ;
        RECT 9.376 5.444 9.408 5.476 ;
  LAYER M2 ;
        RECT 11.744 5.508 11.776 5.54 ;
  LAYER M2 ;
        RECT 9.376 5.572 9.408 5.604 ;
  LAYER M2 ;
        RECT 11.744 5.636 11.776 5.668 ;
  LAYER M2 ;
        RECT 9.376 5.7 9.408 5.732 ;
  LAYER M2 ;
        RECT 11.744 5.764 11.776 5.796 ;
  LAYER M2 ;
        RECT 9.376 5.828 9.408 5.86 ;
  LAYER M2 ;
        RECT 11.744 5.892 11.776 5.924 ;
  LAYER M2 ;
        RECT 9.376 5.956 9.408 5.988 ;
  LAYER M2 ;
        RECT 11.744 6.02 11.776 6.052 ;
  LAYER M2 ;
        RECT 9.376 6.084 9.408 6.116 ;
  LAYER M2 ;
        RECT 11.744 6.148 11.776 6.18 ;
  LAYER M2 ;
        RECT 9.376 6.212 9.408 6.244 ;
  LAYER M2 ;
        RECT 11.744 6.276 11.776 6.308 ;
  LAYER M2 ;
        RECT 9.376 6.34 9.408 6.372 ;
  LAYER M2 ;
        RECT 11.744 6.404 11.776 6.436 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.376 7.188 9.408 9.696 ;
  LAYER M3 ;
        RECT 9.376 9.644 9.408 9.676 ;
  LAYER M1 ;
        RECT 9.44 7.188 9.472 9.696 ;
  LAYER M3 ;
        RECT 9.44 7.208 9.472 7.24 ;
  LAYER M1 ;
        RECT 9.504 7.188 9.536 9.696 ;
  LAYER M3 ;
        RECT 9.504 9.644 9.536 9.676 ;
  LAYER M1 ;
        RECT 9.568 7.188 9.6 9.696 ;
  LAYER M3 ;
        RECT 9.568 7.208 9.6 7.24 ;
  LAYER M1 ;
        RECT 9.632 7.188 9.664 9.696 ;
  LAYER M3 ;
        RECT 9.632 9.644 9.664 9.676 ;
  LAYER M1 ;
        RECT 9.696 7.188 9.728 9.696 ;
  LAYER M3 ;
        RECT 9.696 7.208 9.728 7.24 ;
  LAYER M1 ;
        RECT 9.76 7.188 9.792 9.696 ;
  LAYER M3 ;
        RECT 9.76 9.644 9.792 9.676 ;
  LAYER M1 ;
        RECT 9.824 7.188 9.856 9.696 ;
  LAYER M3 ;
        RECT 9.824 7.208 9.856 7.24 ;
  LAYER M1 ;
        RECT 9.888 7.188 9.92 9.696 ;
  LAYER M3 ;
        RECT 9.888 9.644 9.92 9.676 ;
  LAYER M1 ;
        RECT 9.952 7.188 9.984 9.696 ;
  LAYER M3 ;
        RECT 9.952 7.208 9.984 7.24 ;
  LAYER M1 ;
        RECT 10.016 7.188 10.048 9.696 ;
  LAYER M3 ;
        RECT 10.016 9.644 10.048 9.676 ;
  LAYER M1 ;
        RECT 10.08 7.188 10.112 9.696 ;
  LAYER M3 ;
        RECT 10.08 7.208 10.112 7.24 ;
  LAYER M1 ;
        RECT 10.144 7.188 10.176 9.696 ;
  LAYER M3 ;
        RECT 10.144 9.644 10.176 9.676 ;
  LAYER M1 ;
        RECT 10.208 7.188 10.24 9.696 ;
  LAYER M3 ;
        RECT 10.208 7.208 10.24 7.24 ;
  LAYER M1 ;
        RECT 10.272 7.188 10.304 9.696 ;
  LAYER M3 ;
        RECT 10.272 9.644 10.304 9.676 ;
  LAYER M1 ;
        RECT 10.336 7.188 10.368 9.696 ;
  LAYER M3 ;
        RECT 10.336 7.208 10.368 7.24 ;
  LAYER M1 ;
        RECT 10.4 7.188 10.432 9.696 ;
  LAYER M3 ;
        RECT 10.4 9.644 10.432 9.676 ;
  LAYER M1 ;
        RECT 10.464 7.188 10.496 9.696 ;
  LAYER M3 ;
        RECT 10.464 7.208 10.496 7.24 ;
  LAYER M1 ;
        RECT 10.528 7.188 10.56 9.696 ;
  LAYER M3 ;
        RECT 10.528 9.644 10.56 9.676 ;
  LAYER M1 ;
        RECT 10.592 7.188 10.624 9.696 ;
  LAYER M3 ;
        RECT 10.592 7.208 10.624 7.24 ;
  LAYER M1 ;
        RECT 10.656 7.188 10.688 9.696 ;
  LAYER M3 ;
        RECT 10.656 9.644 10.688 9.676 ;
  LAYER M1 ;
        RECT 10.72 7.188 10.752 9.696 ;
  LAYER M3 ;
        RECT 10.72 7.208 10.752 7.24 ;
  LAYER M1 ;
        RECT 10.784 7.188 10.816 9.696 ;
  LAYER M3 ;
        RECT 10.784 9.644 10.816 9.676 ;
  LAYER M1 ;
        RECT 10.848 7.188 10.88 9.696 ;
  LAYER M3 ;
        RECT 10.848 7.208 10.88 7.24 ;
  LAYER M1 ;
        RECT 10.912 7.188 10.944 9.696 ;
  LAYER M3 ;
        RECT 10.912 9.644 10.944 9.676 ;
  LAYER M1 ;
        RECT 10.976 7.188 11.008 9.696 ;
  LAYER M3 ;
        RECT 10.976 7.208 11.008 7.24 ;
  LAYER M1 ;
        RECT 11.04 7.188 11.072 9.696 ;
  LAYER M3 ;
        RECT 11.04 9.644 11.072 9.676 ;
  LAYER M1 ;
        RECT 11.104 7.188 11.136 9.696 ;
  LAYER M3 ;
        RECT 11.104 7.208 11.136 7.24 ;
  LAYER M1 ;
        RECT 11.168 7.188 11.2 9.696 ;
  LAYER M3 ;
        RECT 11.168 9.644 11.2 9.676 ;
  LAYER M1 ;
        RECT 11.232 7.188 11.264 9.696 ;
  LAYER M3 ;
        RECT 11.232 7.208 11.264 7.24 ;
  LAYER M1 ;
        RECT 11.296 7.188 11.328 9.696 ;
  LAYER M3 ;
        RECT 11.296 9.644 11.328 9.676 ;
  LAYER M1 ;
        RECT 11.36 7.188 11.392 9.696 ;
  LAYER M3 ;
        RECT 11.36 7.208 11.392 7.24 ;
  LAYER M1 ;
        RECT 11.424 7.188 11.456 9.696 ;
  LAYER M3 ;
        RECT 11.424 9.644 11.456 9.676 ;
  LAYER M1 ;
        RECT 11.488 7.188 11.52 9.696 ;
  LAYER M3 ;
        RECT 11.488 7.208 11.52 7.24 ;
  LAYER M1 ;
        RECT 11.552 7.188 11.584 9.696 ;
  LAYER M3 ;
        RECT 11.552 9.644 11.584 9.676 ;
  LAYER M1 ;
        RECT 11.616 7.188 11.648 9.696 ;
  LAYER M3 ;
        RECT 11.616 7.208 11.648 7.24 ;
  LAYER M1 ;
        RECT 11.68 7.188 11.712 9.696 ;
  LAYER M3 ;
        RECT 11.68 9.644 11.712 9.676 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 9.696 ;
  LAYER M3 ;
        RECT 9.376 7.272 9.408 7.304 ;
  LAYER M2 ;
        RECT 11.744 7.336 11.776 7.368 ;
  LAYER M2 ;
        RECT 9.376 7.4 9.408 7.432 ;
  LAYER M2 ;
        RECT 11.744 7.464 11.776 7.496 ;
  LAYER M2 ;
        RECT 9.376 7.528 9.408 7.56 ;
  LAYER M2 ;
        RECT 11.744 7.592 11.776 7.624 ;
  LAYER M2 ;
        RECT 9.376 7.656 9.408 7.688 ;
  LAYER M2 ;
        RECT 11.744 7.72 11.776 7.752 ;
  LAYER M2 ;
        RECT 9.376 7.784 9.408 7.816 ;
  LAYER M2 ;
        RECT 11.744 7.848 11.776 7.88 ;
  LAYER M2 ;
        RECT 9.376 7.912 9.408 7.944 ;
  LAYER M2 ;
        RECT 11.744 7.976 11.776 8.008 ;
  LAYER M2 ;
        RECT 9.376 8.04 9.408 8.072 ;
  LAYER M2 ;
        RECT 11.744 8.104 11.776 8.136 ;
  LAYER M2 ;
        RECT 9.376 8.168 9.408 8.2 ;
  LAYER M2 ;
        RECT 11.744 8.232 11.776 8.264 ;
  LAYER M2 ;
        RECT 9.376 8.296 9.408 8.328 ;
  LAYER M2 ;
        RECT 11.744 8.36 11.776 8.392 ;
  LAYER M2 ;
        RECT 9.376 8.424 9.408 8.456 ;
  LAYER M2 ;
        RECT 11.744 8.488 11.776 8.52 ;
  LAYER M2 ;
        RECT 9.376 8.552 9.408 8.584 ;
  LAYER M2 ;
        RECT 11.744 8.616 11.776 8.648 ;
  LAYER M2 ;
        RECT 9.376 8.68 9.408 8.712 ;
  LAYER M2 ;
        RECT 11.744 8.744 11.776 8.776 ;
  LAYER M2 ;
        RECT 9.376 8.808 9.408 8.84 ;
  LAYER M2 ;
        RECT 11.744 8.872 11.776 8.904 ;
  LAYER M2 ;
        RECT 9.376 8.936 9.408 8.968 ;
  LAYER M2 ;
        RECT 11.744 9 11.776 9.032 ;
  LAYER M2 ;
        RECT 9.376 9.064 9.408 9.096 ;
  LAYER M2 ;
        RECT 11.744 9.128 11.776 9.16 ;
  LAYER M2 ;
        RECT 9.376 9.192 9.408 9.224 ;
  LAYER M2 ;
        RECT 11.744 9.256 11.776 9.288 ;
  LAYER M2 ;
        RECT 9.376 9.32 9.408 9.352 ;
  LAYER M2 ;
        RECT 11.744 9.384 11.776 9.416 ;
  LAYER M2 ;
        RECT 9.376 9.448 9.408 9.48 ;
  LAYER M2 ;
        RECT 11.744 9.512 11.776 9.544 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.376 10.296 9.408 12.804 ;
  LAYER M3 ;
        RECT 9.376 12.752 9.408 12.784 ;
  LAYER M1 ;
        RECT 9.44 10.296 9.472 12.804 ;
  LAYER M3 ;
        RECT 9.44 10.316 9.472 10.348 ;
  LAYER M1 ;
        RECT 9.504 10.296 9.536 12.804 ;
  LAYER M3 ;
        RECT 9.504 12.752 9.536 12.784 ;
  LAYER M1 ;
        RECT 9.568 10.296 9.6 12.804 ;
  LAYER M3 ;
        RECT 9.568 10.316 9.6 10.348 ;
  LAYER M1 ;
        RECT 9.632 10.296 9.664 12.804 ;
  LAYER M3 ;
        RECT 9.632 12.752 9.664 12.784 ;
  LAYER M1 ;
        RECT 9.696 10.296 9.728 12.804 ;
  LAYER M3 ;
        RECT 9.696 10.316 9.728 10.348 ;
  LAYER M1 ;
        RECT 9.76 10.296 9.792 12.804 ;
  LAYER M3 ;
        RECT 9.76 12.752 9.792 12.784 ;
  LAYER M1 ;
        RECT 9.824 10.296 9.856 12.804 ;
  LAYER M3 ;
        RECT 9.824 10.316 9.856 10.348 ;
  LAYER M1 ;
        RECT 9.888 10.296 9.92 12.804 ;
  LAYER M3 ;
        RECT 9.888 12.752 9.92 12.784 ;
  LAYER M1 ;
        RECT 9.952 10.296 9.984 12.804 ;
  LAYER M3 ;
        RECT 9.952 10.316 9.984 10.348 ;
  LAYER M1 ;
        RECT 10.016 10.296 10.048 12.804 ;
  LAYER M3 ;
        RECT 10.016 12.752 10.048 12.784 ;
  LAYER M1 ;
        RECT 10.08 10.296 10.112 12.804 ;
  LAYER M3 ;
        RECT 10.08 10.316 10.112 10.348 ;
  LAYER M1 ;
        RECT 10.144 10.296 10.176 12.804 ;
  LAYER M3 ;
        RECT 10.144 12.752 10.176 12.784 ;
  LAYER M1 ;
        RECT 10.208 10.296 10.24 12.804 ;
  LAYER M3 ;
        RECT 10.208 10.316 10.24 10.348 ;
  LAYER M1 ;
        RECT 10.272 10.296 10.304 12.804 ;
  LAYER M3 ;
        RECT 10.272 12.752 10.304 12.784 ;
  LAYER M1 ;
        RECT 10.336 10.296 10.368 12.804 ;
  LAYER M3 ;
        RECT 10.336 10.316 10.368 10.348 ;
  LAYER M1 ;
        RECT 10.4 10.296 10.432 12.804 ;
  LAYER M3 ;
        RECT 10.4 12.752 10.432 12.784 ;
  LAYER M1 ;
        RECT 10.464 10.296 10.496 12.804 ;
  LAYER M3 ;
        RECT 10.464 10.316 10.496 10.348 ;
  LAYER M1 ;
        RECT 10.528 10.296 10.56 12.804 ;
  LAYER M3 ;
        RECT 10.528 12.752 10.56 12.784 ;
  LAYER M1 ;
        RECT 10.592 10.296 10.624 12.804 ;
  LAYER M3 ;
        RECT 10.592 10.316 10.624 10.348 ;
  LAYER M1 ;
        RECT 10.656 10.296 10.688 12.804 ;
  LAYER M3 ;
        RECT 10.656 12.752 10.688 12.784 ;
  LAYER M1 ;
        RECT 10.72 10.296 10.752 12.804 ;
  LAYER M3 ;
        RECT 10.72 10.316 10.752 10.348 ;
  LAYER M1 ;
        RECT 10.784 10.296 10.816 12.804 ;
  LAYER M3 ;
        RECT 10.784 12.752 10.816 12.784 ;
  LAYER M1 ;
        RECT 10.848 10.296 10.88 12.804 ;
  LAYER M3 ;
        RECT 10.848 10.316 10.88 10.348 ;
  LAYER M1 ;
        RECT 10.912 10.296 10.944 12.804 ;
  LAYER M3 ;
        RECT 10.912 12.752 10.944 12.784 ;
  LAYER M1 ;
        RECT 10.976 10.296 11.008 12.804 ;
  LAYER M3 ;
        RECT 10.976 10.316 11.008 10.348 ;
  LAYER M1 ;
        RECT 11.04 10.296 11.072 12.804 ;
  LAYER M3 ;
        RECT 11.04 12.752 11.072 12.784 ;
  LAYER M1 ;
        RECT 11.104 10.296 11.136 12.804 ;
  LAYER M3 ;
        RECT 11.104 10.316 11.136 10.348 ;
  LAYER M1 ;
        RECT 11.168 10.296 11.2 12.804 ;
  LAYER M3 ;
        RECT 11.168 12.752 11.2 12.784 ;
  LAYER M1 ;
        RECT 11.232 10.296 11.264 12.804 ;
  LAYER M3 ;
        RECT 11.232 10.316 11.264 10.348 ;
  LAYER M1 ;
        RECT 11.296 10.296 11.328 12.804 ;
  LAYER M3 ;
        RECT 11.296 12.752 11.328 12.784 ;
  LAYER M1 ;
        RECT 11.36 10.296 11.392 12.804 ;
  LAYER M3 ;
        RECT 11.36 10.316 11.392 10.348 ;
  LAYER M1 ;
        RECT 11.424 10.296 11.456 12.804 ;
  LAYER M3 ;
        RECT 11.424 12.752 11.456 12.784 ;
  LAYER M1 ;
        RECT 11.488 10.296 11.52 12.804 ;
  LAYER M3 ;
        RECT 11.488 10.316 11.52 10.348 ;
  LAYER M1 ;
        RECT 11.552 10.296 11.584 12.804 ;
  LAYER M3 ;
        RECT 11.552 12.752 11.584 12.784 ;
  LAYER M1 ;
        RECT 11.616 10.296 11.648 12.804 ;
  LAYER M3 ;
        RECT 11.616 10.316 11.648 10.348 ;
  LAYER M1 ;
        RECT 11.68 10.296 11.712 12.804 ;
  LAYER M3 ;
        RECT 11.68 12.752 11.712 12.784 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 12.804 ;
  LAYER M3 ;
        RECT 9.376 10.38 9.408 10.412 ;
  LAYER M2 ;
        RECT 11.744 10.444 11.776 10.476 ;
  LAYER M2 ;
        RECT 9.376 10.508 9.408 10.54 ;
  LAYER M2 ;
        RECT 11.744 10.572 11.776 10.604 ;
  LAYER M2 ;
        RECT 9.376 10.636 9.408 10.668 ;
  LAYER M2 ;
        RECT 11.744 10.7 11.776 10.732 ;
  LAYER M2 ;
        RECT 9.376 10.764 9.408 10.796 ;
  LAYER M2 ;
        RECT 11.744 10.828 11.776 10.86 ;
  LAYER M2 ;
        RECT 9.376 10.892 9.408 10.924 ;
  LAYER M2 ;
        RECT 11.744 10.956 11.776 10.988 ;
  LAYER M2 ;
        RECT 9.376 11.02 9.408 11.052 ;
  LAYER M2 ;
        RECT 11.744 11.084 11.776 11.116 ;
  LAYER M2 ;
        RECT 9.376 11.148 9.408 11.18 ;
  LAYER M2 ;
        RECT 11.744 11.212 11.776 11.244 ;
  LAYER M2 ;
        RECT 9.376 11.276 9.408 11.308 ;
  LAYER M2 ;
        RECT 11.744 11.34 11.776 11.372 ;
  LAYER M2 ;
        RECT 9.376 11.404 9.408 11.436 ;
  LAYER M2 ;
        RECT 11.744 11.468 11.776 11.5 ;
  LAYER M2 ;
        RECT 9.376 11.532 9.408 11.564 ;
  LAYER M2 ;
        RECT 11.744 11.596 11.776 11.628 ;
  LAYER M2 ;
        RECT 9.376 11.66 9.408 11.692 ;
  LAYER M2 ;
        RECT 11.744 11.724 11.776 11.756 ;
  LAYER M2 ;
        RECT 9.376 11.788 9.408 11.82 ;
  LAYER M2 ;
        RECT 11.744 11.852 11.776 11.884 ;
  LAYER M2 ;
        RECT 9.376 11.916 9.408 11.948 ;
  LAYER M2 ;
        RECT 11.744 11.98 11.776 12.012 ;
  LAYER M2 ;
        RECT 9.376 12.044 9.408 12.076 ;
  LAYER M2 ;
        RECT 11.744 12.108 11.776 12.14 ;
  LAYER M2 ;
        RECT 9.376 12.172 9.408 12.204 ;
  LAYER M2 ;
        RECT 11.744 12.236 11.776 12.268 ;
  LAYER M2 ;
        RECT 9.376 12.3 9.408 12.332 ;
  LAYER M2 ;
        RECT 11.744 12.364 11.776 12.396 ;
  LAYER M2 ;
        RECT 9.376 12.428 9.408 12.46 ;
  LAYER M2 ;
        RECT 11.744 12.492 11.776 12.524 ;
  LAYER M2 ;
        RECT 9.376 12.556 9.408 12.588 ;
  LAYER M2 ;
        RECT 11.744 12.62 11.776 12.652 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 9.376 13.404 9.408 15.912 ;
  LAYER M3 ;
        RECT 9.376 15.86 9.408 15.892 ;
  LAYER M1 ;
        RECT 9.44 13.404 9.472 15.912 ;
  LAYER M3 ;
        RECT 9.44 13.424 9.472 13.456 ;
  LAYER M1 ;
        RECT 9.504 13.404 9.536 15.912 ;
  LAYER M3 ;
        RECT 9.504 15.86 9.536 15.892 ;
  LAYER M1 ;
        RECT 9.568 13.404 9.6 15.912 ;
  LAYER M3 ;
        RECT 9.568 13.424 9.6 13.456 ;
  LAYER M1 ;
        RECT 9.632 13.404 9.664 15.912 ;
  LAYER M3 ;
        RECT 9.632 15.86 9.664 15.892 ;
  LAYER M1 ;
        RECT 9.696 13.404 9.728 15.912 ;
  LAYER M3 ;
        RECT 9.696 13.424 9.728 13.456 ;
  LAYER M1 ;
        RECT 9.76 13.404 9.792 15.912 ;
  LAYER M3 ;
        RECT 9.76 15.86 9.792 15.892 ;
  LAYER M1 ;
        RECT 9.824 13.404 9.856 15.912 ;
  LAYER M3 ;
        RECT 9.824 13.424 9.856 13.456 ;
  LAYER M1 ;
        RECT 9.888 13.404 9.92 15.912 ;
  LAYER M3 ;
        RECT 9.888 15.86 9.92 15.892 ;
  LAYER M1 ;
        RECT 9.952 13.404 9.984 15.912 ;
  LAYER M3 ;
        RECT 9.952 13.424 9.984 13.456 ;
  LAYER M1 ;
        RECT 10.016 13.404 10.048 15.912 ;
  LAYER M3 ;
        RECT 10.016 15.86 10.048 15.892 ;
  LAYER M1 ;
        RECT 10.08 13.404 10.112 15.912 ;
  LAYER M3 ;
        RECT 10.08 13.424 10.112 13.456 ;
  LAYER M1 ;
        RECT 10.144 13.404 10.176 15.912 ;
  LAYER M3 ;
        RECT 10.144 15.86 10.176 15.892 ;
  LAYER M1 ;
        RECT 10.208 13.404 10.24 15.912 ;
  LAYER M3 ;
        RECT 10.208 13.424 10.24 13.456 ;
  LAYER M1 ;
        RECT 10.272 13.404 10.304 15.912 ;
  LAYER M3 ;
        RECT 10.272 15.86 10.304 15.892 ;
  LAYER M1 ;
        RECT 10.336 13.404 10.368 15.912 ;
  LAYER M3 ;
        RECT 10.336 13.424 10.368 13.456 ;
  LAYER M1 ;
        RECT 10.4 13.404 10.432 15.912 ;
  LAYER M3 ;
        RECT 10.4 15.86 10.432 15.892 ;
  LAYER M1 ;
        RECT 10.464 13.404 10.496 15.912 ;
  LAYER M3 ;
        RECT 10.464 13.424 10.496 13.456 ;
  LAYER M1 ;
        RECT 10.528 13.404 10.56 15.912 ;
  LAYER M3 ;
        RECT 10.528 15.86 10.56 15.892 ;
  LAYER M1 ;
        RECT 10.592 13.404 10.624 15.912 ;
  LAYER M3 ;
        RECT 10.592 13.424 10.624 13.456 ;
  LAYER M1 ;
        RECT 10.656 13.404 10.688 15.912 ;
  LAYER M3 ;
        RECT 10.656 15.86 10.688 15.892 ;
  LAYER M1 ;
        RECT 10.72 13.404 10.752 15.912 ;
  LAYER M3 ;
        RECT 10.72 13.424 10.752 13.456 ;
  LAYER M1 ;
        RECT 10.784 13.404 10.816 15.912 ;
  LAYER M3 ;
        RECT 10.784 15.86 10.816 15.892 ;
  LAYER M1 ;
        RECT 10.848 13.404 10.88 15.912 ;
  LAYER M3 ;
        RECT 10.848 13.424 10.88 13.456 ;
  LAYER M1 ;
        RECT 10.912 13.404 10.944 15.912 ;
  LAYER M3 ;
        RECT 10.912 15.86 10.944 15.892 ;
  LAYER M1 ;
        RECT 10.976 13.404 11.008 15.912 ;
  LAYER M3 ;
        RECT 10.976 13.424 11.008 13.456 ;
  LAYER M1 ;
        RECT 11.04 13.404 11.072 15.912 ;
  LAYER M3 ;
        RECT 11.04 15.86 11.072 15.892 ;
  LAYER M1 ;
        RECT 11.104 13.404 11.136 15.912 ;
  LAYER M3 ;
        RECT 11.104 13.424 11.136 13.456 ;
  LAYER M1 ;
        RECT 11.168 13.404 11.2 15.912 ;
  LAYER M3 ;
        RECT 11.168 15.86 11.2 15.892 ;
  LAYER M1 ;
        RECT 11.232 13.404 11.264 15.912 ;
  LAYER M3 ;
        RECT 11.232 13.424 11.264 13.456 ;
  LAYER M1 ;
        RECT 11.296 13.404 11.328 15.912 ;
  LAYER M3 ;
        RECT 11.296 15.86 11.328 15.892 ;
  LAYER M1 ;
        RECT 11.36 13.404 11.392 15.912 ;
  LAYER M3 ;
        RECT 11.36 13.424 11.392 13.456 ;
  LAYER M1 ;
        RECT 11.424 13.404 11.456 15.912 ;
  LAYER M3 ;
        RECT 11.424 15.86 11.456 15.892 ;
  LAYER M1 ;
        RECT 11.488 13.404 11.52 15.912 ;
  LAYER M3 ;
        RECT 11.488 13.424 11.52 13.456 ;
  LAYER M1 ;
        RECT 11.552 13.404 11.584 15.912 ;
  LAYER M3 ;
        RECT 11.552 15.86 11.584 15.892 ;
  LAYER M1 ;
        RECT 11.616 13.404 11.648 15.912 ;
  LAYER M3 ;
        RECT 11.616 13.424 11.648 13.456 ;
  LAYER M1 ;
        RECT 11.68 13.404 11.712 15.912 ;
  LAYER M3 ;
        RECT 11.68 15.86 11.712 15.892 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 15.912 ;
  LAYER M3 ;
        RECT 9.376 13.488 9.408 13.52 ;
  LAYER M2 ;
        RECT 11.744 13.552 11.776 13.584 ;
  LAYER M2 ;
        RECT 9.376 13.616 9.408 13.648 ;
  LAYER M2 ;
        RECT 11.744 13.68 11.776 13.712 ;
  LAYER M2 ;
        RECT 9.376 13.744 9.408 13.776 ;
  LAYER M2 ;
        RECT 11.744 13.808 11.776 13.84 ;
  LAYER M2 ;
        RECT 9.376 13.872 9.408 13.904 ;
  LAYER M2 ;
        RECT 11.744 13.936 11.776 13.968 ;
  LAYER M2 ;
        RECT 9.376 14 9.408 14.032 ;
  LAYER M2 ;
        RECT 11.744 14.064 11.776 14.096 ;
  LAYER M2 ;
        RECT 9.376 14.128 9.408 14.16 ;
  LAYER M2 ;
        RECT 11.744 14.192 11.776 14.224 ;
  LAYER M2 ;
        RECT 9.376 14.256 9.408 14.288 ;
  LAYER M2 ;
        RECT 11.744 14.32 11.776 14.352 ;
  LAYER M2 ;
        RECT 9.376 14.384 9.408 14.416 ;
  LAYER M2 ;
        RECT 11.744 14.448 11.776 14.48 ;
  LAYER M2 ;
        RECT 9.376 14.512 9.408 14.544 ;
  LAYER M2 ;
        RECT 11.744 14.576 11.776 14.608 ;
  LAYER M2 ;
        RECT 9.376 14.64 9.408 14.672 ;
  LAYER M2 ;
        RECT 11.744 14.704 11.776 14.736 ;
  LAYER M2 ;
        RECT 9.376 14.768 9.408 14.8 ;
  LAYER M2 ;
        RECT 11.744 14.832 11.776 14.864 ;
  LAYER M2 ;
        RECT 9.376 14.896 9.408 14.928 ;
  LAYER M2 ;
        RECT 11.744 14.96 11.776 14.992 ;
  LAYER M2 ;
        RECT 9.376 15.024 9.408 15.056 ;
  LAYER M2 ;
        RECT 11.744 15.088 11.776 15.12 ;
  LAYER M2 ;
        RECT 9.376 15.152 9.408 15.184 ;
  LAYER M2 ;
        RECT 11.744 15.216 11.776 15.248 ;
  LAYER M2 ;
        RECT 9.376 15.28 9.408 15.312 ;
  LAYER M2 ;
        RECT 11.744 15.344 11.776 15.376 ;
  LAYER M2 ;
        RECT 9.376 15.408 9.408 15.44 ;
  LAYER M2 ;
        RECT 11.744 15.472 11.776 15.504 ;
  LAYER M2 ;
        RECT 9.376 15.536 9.408 15.568 ;
  LAYER M2 ;
        RECT 11.744 15.6 11.776 15.632 ;
  LAYER M2 ;
        RECT 9.376 15.664 9.408 15.696 ;
  LAYER M2 ;
        RECT 11.744 15.728 11.776 15.76 ;
  LAYER M2 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M1 ;
        RECT 12.352 0.972 12.384 3.48 ;
  LAYER M3 ;
        RECT 12.352 3.428 12.384 3.46 ;
  LAYER M1 ;
        RECT 12.416 0.972 12.448 3.48 ;
  LAYER M3 ;
        RECT 12.416 0.992 12.448 1.024 ;
  LAYER M1 ;
        RECT 12.48 0.972 12.512 3.48 ;
  LAYER M3 ;
        RECT 12.48 3.428 12.512 3.46 ;
  LAYER M1 ;
        RECT 12.544 0.972 12.576 3.48 ;
  LAYER M3 ;
        RECT 12.544 0.992 12.576 1.024 ;
  LAYER M1 ;
        RECT 12.608 0.972 12.64 3.48 ;
  LAYER M3 ;
        RECT 12.608 3.428 12.64 3.46 ;
  LAYER M1 ;
        RECT 12.672 0.972 12.704 3.48 ;
  LAYER M3 ;
        RECT 12.672 0.992 12.704 1.024 ;
  LAYER M1 ;
        RECT 12.736 0.972 12.768 3.48 ;
  LAYER M3 ;
        RECT 12.736 3.428 12.768 3.46 ;
  LAYER M1 ;
        RECT 12.8 0.972 12.832 3.48 ;
  LAYER M3 ;
        RECT 12.8 0.992 12.832 1.024 ;
  LAYER M1 ;
        RECT 12.864 0.972 12.896 3.48 ;
  LAYER M3 ;
        RECT 12.864 3.428 12.896 3.46 ;
  LAYER M1 ;
        RECT 12.928 0.972 12.96 3.48 ;
  LAYER M3 ;
        RECT 12.928 0.992 12.96 1.024 ;
  LAYER M1 ;
        RECT 12.992 0.972 13.024 3.48 ;
  LAYER M3 ;
        RECT 12.992 3.428 13.024 3.46 ;
  LAYER M1 ;
        RECT 13.056 0.972 13.088 3.48 ;
  LAYER M3 ;
        RECT 13.056 0.992 13.088 1.024 ;
  LAYER M1 ;
        RECT 13.12 0.972 13.152 3.48 ;
  LAYER M3 ;
        RECT 13.12 3.428 13.152 3.46 ;
  LAYER M1 ;
        RECT 13.184 0.972 13.216 3.48 ;
  LAYER M3 ;
        RECT 13.184 0.992 13.216 1.024 ;
  LAYER M1 ;
        RECT 13.248 0.972 13.28 3.48 ;
  LAYER M3 ;
        RECT 13.248 3.428 13.28 3.46 ;
  LAYER M1 ;
        RECT 13.312 0.972 13.344 3.48 ;
  LAYER M3 ;
        RECT 13.312 0.992 13.344 1.024 ;
  LAYER M1 ;
        RECT 13.376 0.972 13.408 3.48 ;
  LAYER M3 ;
        RECT 13.376 3.428 13.408 3.46 ;
  LAYER M1 ;
        RECT 13.44 0.972 13.472 3.48 ;
  LAYER M3 ;
        RECT 13.44 0.992 13.472 1.024 ;
  LAYER M1 ;
        RECT 13.504 0.972 13.536 3.48 ;
  LAYER M3 ;
        RECT 13.504 3.428 13.536 3.46 ;
  LAYER M1 ;
        RECT 13.568 0.972 13.6 3.48 ;
  LAYER M3 ;
        RECT 13.568 0.992 13.6 1.024 ;
  LAYER M1 ;
        RECT 13.632 0.972 13.664 3.48 ;
  LAYER M3 ;
        RECT 13.632 3.428 13.664 3.46 ;
  LAYER M1 ;
        RECT 13.696 0.972 13.728 3.48 ;
  LAYER M3 ;
        RECT 13.696 0.992 13.728 1.024 ;
  LAYER M1 ;
        RECT 13.76 0.972 13.792 3.48 ;
  LAYER M3 ;
        RECT 13.76 3.428 13.792 3.46 ;
  LAYER M1 ;
        RECT 13.824 0.972 13.856 3.48 ;
  LAYER M3 ;
        RECT 13.824 0.992 13.856 1.024 ;
  LAYER M1 ;
        RECT 13.888 0.972 13.92 3.48 ;
  LAYER M3 ;
        RECT 13.888 3.428 13.92 3.46 ;
  LAYER M1 ;
        RECT 13.952 0.972 13.984 3.48 ;
  LAYER M3 ;
        RECT 13.952 0.992 13.984 1.024 ;
  LAYER M1 ;
        RECT 14.016 0.972 14.048 3.48 ;
  LAYER M3 ;
        RECT 14.016 3.428 14.048 3.46 ;
  LAYER M1 ;
        RECT 14.08 0.972 14.112 3.48 ;
  LAYER M3 ;
        RECT 14.08 0.992 14.112 1.024 ;
  LAYER M1 ;
        RECT 14.144 0.972 14.176 3.48 ;
  LAYER M3 ;
        RECT 14.144 3.428 14.176 3.46 ;
  LAYER M1 ;
        RECT 14.208 0.972 14.24 3.48 ;
  LAYER M3 ;
        RECT 14.208 0.992 14.24 1.024 ;
  LAYER M1 ;
        RECT 14.272 0.972 14.304 3.48 ;
  LAYER M3 ;
        RECT 14.272 3.428 14.304 3.46 ;
  LAYER M1 ;
        RECT 14.336 0.972 14.368 3.48 ;
  LAYER M3 ;
        RECT 14.336 0.992 14.368 1.024 ;
  LAYER M1 ;
        RECT 14.4 0.972 14.432 3.48 ;
  LAYER M3 ;
        RECT 14.4 3.428 14.432 3.46 ;
  LAYER M1 ;
        RECT 14.464 0.972 14.496 3.48 ;
  LAYER M3 ;
        RECT 14.464 0.992 14.496 1.024 ;
  LAYER M1 ;
        RECT 14.528 0.972 14.56 3.48 ;
  LAYER M3 ;
        RECT 14.528 3.428 14.56 3.46 ;
  LAYER M1 ;
        RECT 14.592 0.972 14.624 3.48 ;
  LAYER M3 ;
        RECT 14.592 0.992 14.624 1.024 ;
  LAYER M1 ;
        RECT 14.656 0.972 14.688 3.48 ;
  LAYER M3 ;
        RECT 14.656 3.428 14.688 3.46 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 3.48 ;
  LAYER M3 ;
        RECT 12.352 1.056 12.384 1.088 ;
  LAYER M2 ;
        RECT 14.72 1.12 14.752 1.152 ;
  LAYER M2 ;
        RECT 12.352 1.184 12.384 1.216 ;
  LAYER M2 ;
        RECT 14.72 1.248 14.752 1.28 ;
  LAYER M2 ;
        RECT 12.352 1.312 12.384 1.344 ;
  LAYER M2 ;
        RECT 14.72 1.376 14.752 1.408 ;
  LAYER M2 ;
        RECT 12.352 1.44 12.384 1.472 ;
  LAYER M2 ;
        RECT 14.72 1.504 14.752 1.536 ;
  LAYER M2 ;
        RECT 12.352 1.568 12.384 1.6 ;
  LAYER M2 ;
        RECT 14.72 1.632 14.752 1.664 ;
  LAYER M2 ;
        RECT 12.352 1.696 12.384 1.728 ;
  LAYER M2 ;
        RECT 14.72 1.76 14.752 1.792 ;
  LAYER M2 ;
        RECT 12.352 1.824 12.384 1.856 ;
  LAYER M2 ;
        RECT 14.72 1.888 14.752 1.92 ;
  LAYER M2 ;
        RECT 12.352 1.952 12.384 1.984 ;
  LAYER M2 ;
        RECT 14.72 2.016 14.752 2.048 ;
  LAYER M2 ;
        RECT 12.352 2.08 12.384 2.112 ;
  LAYER M2 ;
        RECT 14.72 2.144 14.752 2.176 ;
  LAYER M2 ;
        RECT 12.352 2.208 12.384 2.24 ;
  LAYER M2 ;
        RECT 14.72 2.272 14.752 2.304 ;
  LAYER M2 ;
        RECT 12.352 2.336 12.384 2.368 ;
  LAYER M2 ;
        RECT 14.72 2.4 14.752 2.432 ;
  LAYER M2 ;
        RECT 12.352 2.464 12.384 2.496 ;
  LAYER M2 ;
        RECT 14.72 2.528 14.752 2.56 ;
  LAYER M2 ;
        RECT 12.352 2.592 12.384 2.624 ;
  LAYER M2 ;
        RECT 14.72 2.656 14.752 2.688 ;
  LAYER M2 ;
        RECT 12.352 2.72 12.384 2.752 ;
  LAYER M2 ;
        RECT 14.72 2.784 14.752 2.816 ;
  LAYER M2 ;
        RECT 12.352 2.848 12.384 2.88 ;
  LAYER M2 ;
        RECT 14.72 2.912 14.752 2.944 ;
  LAYER M2 ;
        RECT 12.352 2.976 12.384 3.008 ;
  LAYER M2 ;
        RECT 14.72 3.04 14.752 3.072 ;
  LAYER M2 ;
        RECT 12.352 3.104 12.384 3.136 ;
  LAYER M2 ;
        RECT 14.72 3.168 14.752 3.2 ;
  LAYER M2 ;
        RECT 12.352 3.232 12.384 3.264 ;
  LAYER M2 ;
        RECT 14.72 3.296 14.752 3.328 ;
  LAYER M2 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M1 ;
        RECT 12.352 4.08 12.384 6.588 ;
  LAYER M3 ;
        RECT 12.352 6.536 12.384 6.568 ;
  LAYER M1 ;
        RECT 12.416 4.08 12.448 6.588 ;
  LAYER M3 ;
        RECT 12.416 4.1 12.448 4.132 ;
  LAYER M1 ;
        RECT 12.48 4.08 12.512 6.588 ;
  LAYER M3 ;
        RECT 12.48 6.536 12.512 6.568 ;
  LAYER M1 ;
        RECT 12.544 4.08 12.576 6.588 ;
  LAYER M3 ;
        RECT 12.544 4.1 12.576 4.132 ;
  LAYER M1 ;
        RECT 12.608 4.08 12.64 6.588 ;
  LAYER M3 ;
        RECT 12.608 6.536 12.64 6.568 ;
  LAYER M1 ;
        RECT 12.672 4.08 12.704 6.588 ;
  LAYER M3 ;
        RECT 12.672 4.1 12.704 4.132 ;
  LAYER M1 ;
        RECT 12.736 4.08 12.768 6.588 ;
  LAYER M3 ;
        RECT 12.736 6.536 12.768 6.568 ;
  LAYER M1 ;
        RECT 12.8 4.08 12.832 6.588 ;
  LAYER M3 ;
        RECT 12.8 4.1 12.832 4.132 ;
  LAYER M1 ;
        RECT 12.864 4.08 12.896 6.588 ;
  LAYER M3 ;
        RECT 12.864 6.536 12.896 6.568 ;
  LAYER M1 ;
        RECT 12.928 4.08 12.96 6.588 ;
  LAYER M3 ;
        RECT 12.928 4.1 12.96 4.132 ;
  LAYER M1 ;
        RECT 12.992 4.08 13.024 6.588 ;
  LAYER M3 ;
        RECT 12.992 6.536 13.024 6.568 ;
  LAYER M1 ;
        RECT 13.056 4.08 13.088 6.588 ;
  LAYER M3 ;
        RECT 13.056 4.1 13.088 4.132 ;
  LAYER M1 ;
        RECT 13.12 4.08 13.152 6.588 ;
  LAYER M3 ;
        RECT 13.12 6.536 13.152 6.568 ;
  LAYER M1 ;
        RECT 13.184 4.08 13.216 6.588 ;
  LAYER M3 ;
        RECT 13.184 4.1 13.216 4.132 ;
  LAYER M1 ;
        RECT 13.248 4.08 13.28 6.588 ;
  LAYER M3 ;
        RECT 13.248 6.536 13.28 6.568 ;
  LAYER M1 ;
        RECT 13.312 4.08 13.344 6.588 ;
  LAYER M3 ;
        RECT 13.312 4.1 13.344 4.132 ;
  LAYER M1 ;
        RECT 13.376 4.08 13.408 6.588 ;
  LAYER M3 ;
        RECT 13.376 6.536 13.408 6.568 ;
  LAYER M1 ;
        RECT 13.44 4.08 13.472 6.588 ;
  LAYER M3 ;
        RECT 13.44 4.1 13.472 4.132 ;
  LAYER M1 ;
        RECT 13.504 4.08 13.536 6.588 ;
  LAYER M3 ;
        RECT 13.504 6.536 13.536 6.568 ;
  LAYER M1 ;
        RECT 13.568 4.08 13.6 6.588 ;
  LAYER M3 ;
        RECT 13.568 4.1 13.6 4.132 ;
  LAYER M1 ;
        RECT 13.632 4.08 13.664 6.588 ;
  LAYER M3 ;
        RECT 13.632 6.536 13.664 6.568 ;
  LAYER M1 ;
        RECT 13.696 4.08 13.728 6.588 ;
  LAYER M3 ;
        RECT 13.696 4.1 13.728 4.132 ;
  LAYER M1 ;
        RECT 13.76 4.08 13.792 6.588 ;
  LAYER M3 ;
        RECT 13.76 6.536 13.792 6.568 ;
  LAYER M1 ;
        RECT 13.824 4.08 13.856 6.588 ;
  LAYER M3 ;
        RECT 13.824 4.1 13.856 4.132 ;
  LAYER M1 ;
        RECT 13.888 4.08 13.92 6.588 ;
  LAYER M3 ;
        RECT 13.888 6.536 13.92 6.568 ;
  LAYER M1 ;
        RECT 13.952 4.08 13.984 6.588 ;
  LAYER M3 ;
        RECT 13.952 4.1 13.984 4.132 ;
  LAYER M1 ;
        RECT 14.016 4.08 14.048 6.588 ;
  LAYER M3 ;
        RECT 14.016 6.536 14.048 6.568 ;
  LAYER M1 ;
        RECT 14.08 4.08 14.112 6.588 ;
  LAYER M3 ;
        RECT 14.08 4.1 14.112 4.132 ;
  LAYER M1 ;
        RECT 14.144 4.08 14.176 6.588 ;
  LAYER M3 ;
        RECT 14.144 6.536 14.176 6.568 ;
  LAYER M1 ;
        RECT 14.208 4.08 14.24 6.588 ;
  LAYER M3 ;
        RECT 14.208 4.1 14.24 4.132 ;
  LAYER M1 ;
        RECT 14.272 4.08 14.304 6.588 ;
  LAYER M3 ;
        RECT 14.272 6.536 14.304 6.568 ;
  LAYER M1 ;
        RECT 14.336 4.08 14.368 6.588 ;
  LAYER M3 ;
        RECT 14.336 4.1 14.368 4.132 ;
  LAYER M1 ;
        RECT 14.4 4.08 14.432 6.588 ;
  LAYER M3 ;
        RECT 14.4 6.536 14.432 6.568 ;
  LAYER M1 ;
        RECT 14.464 4.08 14.496 6.588 ;
  LAYER M3 ;
        RECT 14.464 4.1 14.496 4.132 ;
  LAYER M1 ;
        RECT 14.528 4.08 14.56 6.588 ;
  LAYER M3 ;
        RECT 14.528 6.536 14.56 6.568 ;
  LAYER M1 ;
        RECT 14.592 4.08 14.624 6.588 ;
  LAYER M3 ;
        RECT 14.592 4.1 14.624 4.132 ;
  LAYER M1 ;
        RECT 14.656 4.08 14.688 6.588 ;
  LAYER M3 ;
        RECT 14.656 6.536 14.688 6.568 ;
  LAYER M1 ;
        RECT 14.72 4.08 14.752 6.588 ;
  LAYER M3 ;
        RECT 12.352 4.164 12.384 4.196 ;
  LAYER M2 ;
        RECT 14.72 4.228 14.752 4.26 ;
  LAYER M2 ;
        RECT 12.352 4.292 12.384 4.324 ;
  LAYER M2 ;
        RECT 14.72 4.356 14.752 4.388 ;
  LAYER M2 ;
        RECT 12.352 4.42 12.384 4.452 ;
  LAYER M2 ;
        RECT 14.72 4.484 14.752 4.516 ;
  LAYER M2 ;
        RECT 12.352 4.548 12.384 4.58 ;
  LAYER M2 ;
        RECT 14.72 4.612 14.752 4.644 ;
  LAYER M2 ;
        RECT 12.352 4.676 12.384 4.708 ;
  LAYER M2 ;
        RECT 14.72 4.74 14.752 4.772 ;
  LAYER M2 ;
        RECT 12.352 4.804 12.384 4.836 ;
  LAYER M2 ;
        RECT 14.72 4.868 14.752 4.9 ;
  LAYER M2 ;
        RECT 12.352 4.932 12.384 4.964 ;
  LAYER M2 ;
        RECT 14.72 4.996 14.752 5.028 ;
  LAYER M2 ;
        RECT 12.352 5.06 12.384 5.092 ;
  LAYER M2 ;
        RECT 14.72 5.124 14.752 5.156 ;
  LAYER M2 ;
        RECT 12.352 5.188 12.384 5.22 ;
  LAYER M2 ;
        RECT 14.72 5.252 14.752 5.284 ;
  LAYER M2 ;
        RECT 12.352 5.316 12.384 5.348 ;
  LAYER M2 ;
        RECT 14.72 5.38 14.752 5.412 ;
  LAYER M2 ;
        RECT 12.352 5.444 12.384 5.476 ;
  LAYER M2 ;
        RECT 14.72 5.508 14.752 5.54 ;
  LAYER M2 ;
        RECT 12.352 5.572 12.384 5.604 ;
  LAYER M2 ;
        RECT 14.72 5.636 14.752 5.668 ;
  LAYER M2 ;
        RECT 12.352 5.7 12.384 5.732 ;
  LAYER M2 ;
        RECT 14.72 5.764 14.752 5.796 ;
  LAYER M2 ;
        RECT 12.352 5.828 12.384 5.86 ;
  LAYER M2 ;
        RECT 14.72 5.892 14.752 5.924 ;
  LAYER M2 ;
        RECT 12.352 5.956 12.384 5.988 ;
  LAYER M2 ;
        RECT 14.72 6.02 14.752 6.052 ;
  LAYER M2 ;
        RECT 12.352 6.084 12.384 6.116 ;
  LAYER M2 ;
        RECT 14.72 6.148 14.752 6.18 ;
  LAYER M2 ;
        RECT 12.352 6.212 12.384 6.244 ;
  LAYER M2 ;
        RECT 14.72 6.276 14.752 6.308 ;
  LAYER M2 ;
        RECT 12.352 6.34 12.384 6.372 ;
  LAYER M2 ;
        RECT 14.72 6.404 14.752 6.436 ;
  LAYER M2 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M1 ;
        RECT 12.352 7.188 12.384 9.696 ;
  LAYER M3 ;
        RECT 12.352 9.644 12.384 9.676 ;
  LAYER M1 ;
        RECT 12.416 7.188 12.448 9.696 ;
  LAYER M3 ;
        RECT 12.416 7.208 12.448 7.24 ;
  LAYER M1 ;
        RECT 12.48 7.188 12.512 9.696 ;
  LAYER M3 ;
        RECT 12.48 9.644 12.512 9.676 ;
  LAYER M1 ;
        RECT 12.544 7.188 12.576 9.696 ;
  LAYER M3 ;
        RECT 12.544 7.208 12.576 7.24 ;
  LAYER M1 ;
        RECT 12.608 7.188 12.64 9.696 ;
  LAYER M3 ;
        RECT 12.608 9.644 12.64 9.676 ;
  LAYER M1 ;
        RECT 12.672 7.188 12.704 9.696 ;
  LAYER M3 ;
        RECT 12.672 7.208 12.704 7.24 ;
  LAYER M1 ;
        RECT 12.736 7.188 12.768 9.696 ;
  LAYER M3 ;
        RECT 12.736 9.644 12.768 9.676 ;
  LAYER M1 ;
        RECT 12.8 7.188 12.832 9.696 ;
  LAYER M3 ;
        RECT 12.8 7.208 12.832 7.24 ;
  LAYER M1 ;
        RECT 12.864 7.188 12.896 9.696 ;
  LAYER M3 ;
        RECT 12.864 9.644 12.896 9.676 ;
  LAYER M1 ;
        RECT 12.928 7.188 12.96 9.696 ;
  LAYER M3 ;
        RECT 12.928 7.208 12.96 7.24 ;
  LAYER M1 ;
        RECT 12.992 7.188 13.024 9.696 ;
  LAYER M3 ;
        RECT 12.992 9.644 13.024 9.676 ;
  LAYER M1 ;
        RECT 13.056 7.188 13.088 9.696 ;
  LAYER M3 ;
        RECT 13.056 7.208 13.088 7.24 ;
  LAYER M1 ;
        RECT 13.12 7.188 13.152 9.696 ;
  LAYER M3 ;
        RECT 13.12 9.644 13.152 9.676 ;
  LAYER M1 ;
        RECT 13.184 7.188 13.216 9.696 ;
  LAYER M3 ;
        RECT 13.184 7.208 13.216 7.24 ;
  LAYER M1 ;
        RECT 13.248 7.188 13.28 9.696 ;
  LAYER M3 ;
        RECT 13.248 9.644 13.28 9.676 ;
  LAYER M1 ;
        RECT 13.312 7.188 13.344 9.696 ;
  LAYER M3 ;
        RECT 13.312 7.208 13.344 7.24 ;
  LAYER M1 ;
        RECT 13.376 7.188 13.408 9.696 ;
  LAYER M3 ;
        RECT 13.376 9.644 13.408 9.676 ;
  LAYER M1 ;
        RECT 13.44 7.188 13.472 9.696 ;
  LAYER M3 ;
        RECT 13.44 7.208 13.472 7.24 ;
  LAYER M1 ;
        RECT 13.504 7.188 13.536 9.696 ;
  LAYER M3 ;
        RECT 13.504 9.644 13.536 9.676 ;
  LAYER M1 ;
        RECT 13.568 7.188 13.6 9.696 ;
  LAYER M3 ;
        RECT 13.568 7.208 13.6 7.24 ;
  LAYER M1 ;
        RECT 13.632 7.188 13.664 9.696 ;
  LAYER M3 ;
        RECT 13.632 9.644 13.664 9.676 ;
  LAYER M1 ;
        RECT 13.696 7.188 13.728 9.696 ;
  LAYER M3 ;
        RECT 13.696 7.208 13.728 7.24 ;
  LAYER M1 ;
        RECT 13.76 7.188 13.792 9.696 ;
  LAYER M3 ;
        RECT 13.76 9.644 13.792 9.676 ;
  LAYER M1 ;
        RECT 13.824 7.188 13.856 9.696 ;
  LAYER M3 ;
        RECT 13.824 7.208 13.856 7.24 ;
  LAYER M1 ;
        RECT 13.888 7.188 13.92 9.696 ;
  LAYER M3 ;
        RECT 13.888 9.644 13.92 9.676 ;
  LAYER M1 ;
        RECT 13.952 7.188 13.984 9.696 ;
  LAYER M3 ;
        RECT 13.952 7.208 13.984 7.24 ;
  LAYER M1 ;
        RECT 14.016 7.188 14.048 9.696 ;
  LAYER M3 ;
        RECT 14.016 9.644 14.048 9.676 ;
  LAYER M1 ;
        RECT 14.08 7.188 14.112 9.696 ;
  LAYER M3 ;
        RECT 14.08 7.208 14.112 7.24 ;
  LAYER M1 ;
        RECT 14.144 7.188 14.176 9.696 ;
  LAYER M3 ;
        RECT 14.144 9.644 14.176 9.676 ;
  LAYER M1 ;
        RECT 14.208 7.188 14.24 9.696 ;
  LAYER M3 ;
        RECT 14.208 7.208 14.24 7.24 ;
  LAYER M1 ;
        RECT 14.272 7.188 14.304 9.696 ;
  LAYER M3 ;
        RECT 14.272 9.644 14.304 9.676 ;
  LAYER M1 ;
        RECT 14.336 7.188 14.368 9.696 ;
  LAYER M3 ;
        RECT 14.336 7.208 14.368 7.24 ;
  LAYER M1 ;
        RECT 14.4 7.188 14.432 9.696 ;
  LAYER M3 ;
        RECT 14.4 9.644 14.432 9.676 ;
  LAYER M1 ;
        RECT 14.464 7.188 14.496 9.696 ;
  LAYER M3 ;
        RECT 14.464 7.208 14.496 7.24 ;
  LAYER M1 ;
        RECT 14.528 7.188 14.56 9.696 ;
  LAYER M3 ;
        RECT 14.528 9.644 14.56 9.676 ;
  LAYER M1 ;
        RECT 14.592 7.188 14.624 9.696 ;
  LAYER M3 ;
        RECT 14.592 7.208 14.624 7.24 ;
  LAYER M1 ;
        RECT 14.656 7.188 14.688 9.696 ;
  LAYER M3 ;
        RECT 14.656 9.644 14.688 9.676 ;
  LAYER M1 ;
        RECT 14.72 7.188 14.752 9.696 ;
  LAYER M3 ;
        RECT 12.352 7.272 12.384 7.304 ;
  LAYER M2 ;
        RECT 14.72 7.336 14.752 7.368 ;
  LAYER M2 ;
        RECT 12.352 7.4 12.384 7.432 ;
  LAYER M2 ;
        RECT 14.72 7.464 14.752 7.496 ;
  LAYER M2 ;
        RECT 12.352 7.528 12.384 7.56 ;
  LAYER M2 ;
        RECT 14.72 7.592 14.752 7.624 ;
  LAYER M2 ;
        RECT 12.352 7.656 12.384 7.688 ;
  LAYER M2 ;
        RECT 14.72 7.72 14.752 7.752 ;
  LAYER M2 ;
        RECT 12.352 7.784 12.384 7.816 ;
  LAYER M2 ;
        RECT 14.72 7.848 14.752 7.88 ;
  LAYER M2 ;
        RECT 12.352 7.912 12.384 7.944 ;
  LAYER M2 ;
        RECT 14.72 7.976 14.752 8.008 ;
  LAYER M2 ;
        RECT 12.352 8.04 12.384 8.072 ;
  LAYER M2 ;
        RECT 14.72 8.104 14.752 8.136 ;
  LAYER M2 ;
        RECT 12.352 8.168 12.384 8.2 ;
  LAYER M2 ;
        RECT 14.72 8.232 14.752 8.264 ;
  LAYER M2 ;
        RECT 12.352 8.296 12.384 8.328 ;
  LAYER M2 ;
        RECT 14.72 8.36 14.752 8.392 ;
  LAYER M2 ;
        RECT 12.352 8.424 12.384 8.456 ;
  LAYER M2 ;
        RECT 14.72 8.488 14.752 8.52 ;
  LAYER M2 ;
        RECT 12.352 8.552 12.384 8.584 ;
  LAYER M2 ;
        RECT 14.72 8.616 14.752 8.648 ;
  LAYER M2 ;
        RECT 12.352 8.68 12.384 8.712 ;
  LAYER M2 ;
        RECT 14.72 8.744 14.752 8.776 ;
  LAYER M2 ;
        RECT 12.352 8.808 12.384 8.84 ;
  LAYER M2 ;
        RECT 14.72 8.872 14.752 8.904 ;
  LAYER M2 ;
        RECT 12.352 8.936 12.384 8.968 ;
  LAYER M2 ;
        RECT 14.72 9 14.752 9.032 ;
  LAYER M2 ;
        RECT 12.352 9.064 12.384 9.096 ;
  LAYER M2 ;
        RECT 14.72 9.128 14.752 9.16 ;
  LAYER M2 ;
        RECT 12.352 9.192 12.384 9.224 ;
  LAYER M2 ;
        RECT 14.72 9.256 14.752 9.288 ;
  LAYER M2 ;
        RECT 12.352 9.32 12.384 9.352 ;
  LAYER M2 ;
        RECT 14.72 9.384 14.752 9.416 ;
  LAYER M2 ;
        RECT 12.352 9.448 12.384 9.48 ;
  LAYER M2 ;
        RECT 14.72 9.512 14.752 9.544 ;
  LAYER M2 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M1 ;
        RECT 12.352 10.296 12.384 12.804 ;
  LAYER M3 ;
        RECT 12.352 12.752 12.384 12.784 ;
  LAYER M1 ;
        RECT 12.416 10.296 12.448 12.804 ;
  LAYER M3 ;
        RECT 12.416 10.316 12.448 10.348 ;
  LAYER M1 ;
        RECT 12.48 10.296 12.512 12.804 ;
  LAYER M3 ;
        RECT 12.48 12.752 12.512 12.784 ;
  LAYER M1 ;
        RECT 12.544 10.296 12.576 12.804 ;
  LAYER M3 ;
        RECT 12.544 10.316 12.576 10.348 ;
  LAYER M1 ;
        RECT 12.608 10.296 12.64 12.804 ;
  LAYER M3 ;
        RECT 12.608 12.752 12.64 12.784 ;
  LAYER M1 ;
        RECT 12.672 10.296 12.704 12.804 ;
  LAYER M3 ;
        RECT 12.672 10.316 12.704 10.348 ;
  LAYER M1 ;
        RECT 12.736 10.296 12.768 12.804 ;
  LAYER M3 ;
        RECT 12.736 12.752 12.768 12.784 ;
  LAYER M1 ;
        RECT 12.8 10.296 12.832 12.804 ;
  LAYER M3 ;
        RECT 12.8 10.316 12.832 10.348 ;
  LAYER M1 ;
        RECT 12.864 10.296 12.896 12.804 ;
  LAYER M3 ;
        RECT 12.864 12.752 12.896 12.784 ;
  LAYER M1 ;
        RECT 12.928 10.296 12.96 12.804 ;
  LAYER M3 ;
        RECT 12.928 10.316 12.96 10.348 ;
  LAYER M1 ;
        RECT 12.992 10.296 13.024 12.804 ;
  LAYER M3 ;
        RECT 12.992 12.752 13.024 12.784 ;
  LAYER M1 ;
        RECT 13.056 10.296 13.088 12.804 ;
  LAYER M3 ;
        RECT 13.056 10.316 13.088 10.348 ;
  LAYER M1 ;
        RECT 13.12 10.296 13.152 12.804 ;
  LAYER M3 ;
        RECT 13.12 12.752 13.152 12.784 ;
  LAYER M1 ;
        RECT 13.184 10.296 13.216 12.804 ;
  LAYER M3 ;
        RECT 13.184 10.316 13.216 10.348 ;
  LAYER M1 ;
        RECT 13.248 10.296 13.28 12.804 ;
  LAYER M3 ;
        RECT 13.248 12.752 13.28 12.784 ;
  LAYER M1 ;
        RECT 13.312 10.296 13.344 12.804 ;
  LAYER M3 ;
        RECT 13.312 10.316 13.344 10.348 ;
  LAYER M1 ;
        RECT 13.376 10.296 13.408 12.804 ;
  LAYER M3 ;
        RECT 13.376 12.752 13.408 12.784 ;
  LAYER M1 ;
        RECT 13.44 10.296 13.472 12.804 ;
  LAYER M3 ;
        RECT 13.44 10.316 13.472 10.348 ;
  LAYER M1 ;
        RECT 13.504 10.296 13.536 12.804 ;
  LAYER M3 ;
        RECT 13.504 12.752 13.536 12.784 ;
  LAYER M1 ;
        RECT 13.568 10.296 13.6 12.804 ;
  LAYER M3 ;
        RECT 13.568 10.316 13.6 10.348 ;
  LAYER M1 ;
        RECT 13.632 10.296 13.664 12.804 ;
  LAYER M3 ;
        RECT 13.632 12.752 13.664 12.784 ;
  LAYER M1 ;
        RECT 13.696 10.296 13.728 12.804 ;
  LAYER M3 ;
        RECT 13.696 10.316 13.728 10.348 ;
  LAYER M1 ;
        RECT 13.76 10.296 13.792 12.804 ;
  LAYER M3 ;
        RECT 13.76 12.752 13.792 12.784 ;
  LAYER M1 ;
        RECT 13.824 10.296 13.856 12.804 ;
  LAYER M3 ;
        RECT 13.824 10.316 13.856 10.348 ;
  LAYER M1 ;
        RECT 13.888 10.296 13.92 12.804 ;
  LAYER M3 ;
        RECT 13.888 12.752 13.92 12.784 ;
  LAYER M1 ;
        RECT 13.952 10.296 13.984 12.804 ;
  LAYER M3 ;
        RECT 13.952 10.316 13.984 10.348 ;
  LAYER M1 ;
        RECT 14.016 10.296 14.048 12.804 ;
  LAYER M3 ;
        RECT 14.016 12.752 14.048 12.784 ;
  LAYER M1 ;
        RECT 14.08 10.296 14.112 12.804 ;
  LAYER M3 ;
        RECT 14.08 10.316 14.112 10.348 ;
  LAYER M1 ;
        RECT 14.144 10.296 14.176 12.804 ;
  LAYER M3 ;
        RECT 14.144 12.752 14.176 12.784 ;
  LAYER M1 ;
        RECT 14.208 10.296 14.24 12.804 ;
  LAYER M3 ;
        RECT 14.208 10.316 14.24 10.348 ;
  LAYER M1 ;
        RECT 14.272 10.296 14.304 12.804 ;
  LAYER M3 ;
        RECT 14.272 12.752 14.304 12.784 ;
  LAYER M1 ;
        RECT 14.336 10.296 14.368 12.804 ;
  LAYER M3 ;
        RECT 14.336 10.316 14.368 10.348 ;
  LAYER M1 ;
        RECT 14.4 10.296 14.432 12.804 ;
  LAYER M3 ;
        RECT 14.4 12.752 14.432 12.784 ;
  LAYER M1 ;
        RECT 14.464 10.296 14.496 12.804 ;
  LAYER M3 ;
        RECT 14.464 10.316 14.496 10.348 ;
  LAYER M1 ;
        RECT 14.528 10.296 14.56 12.804 ;
  LAYER M3 ;
        RECT 14.528 12.752 14.56 12.784 ;
  LAYER M1 ;
        RECT 14.592 10.296 14.624 12.804 ;
  LAYER M3 ;
        RECT 14.592 10.316 14.624 10.348 ;
  LAYER M1 ;
        RECT 14.656 10.296 14.688 12.804 ;
  LAYER M3 ;
        RECT 14.656 12.752 14.688 12.784 ;
  LAYER M1 ;
        RECT 14.72 10.296 14.752 12.804 ;
  LAYER M3 ;
        RECT 12.352 10.38 12.384 10.412 ;
  LAYER M2 ;
        RECT 14.72 10.444 14.752 10.476 ;
  LAYER M2 ;
        RECT 12.352 10.508 12.384 10.54 ;
  LAYER M2 ;
        RECT 14.72 10.572 14.752 10.604 ;
  LAYER M2 ;
        RECT 12.352 10.636 12.384 10.668 ;
  LAYER M2 ;
        RECT 14.72 10.7 14.752 10.732 ;
  LAYER M2 ;
        RECT 12.352 10.764 12.384 10.796 ;
  LAYER M2 ;
        RECT 14.72 10.828 14.752 10.86 ;
  LAYER M2 ;
        RECT 12.352 10.892 12.384 10.924 ;
  LAYER M2 ;
        RECT 14.72 10.956 14.752 10.988 ;
  LAYER M2 ;
        RECT 12.352 11.02 12.384 11.052 ;
  LAYER M2 ;
        RECT 14.72 11.084 14.752 11.116 ;
  LAYER M2 ;
        RECT 12.352 11.148 12.384 11.18 ;
  LAYER M2 ;
        RECT 14.72 11.212 14.752 11.244 ;
  LAYER M2 ;
        RECT 12.352 11.276 12.384 11.308 ;
  LAYER M2 ;
        RECT 14.72 11.34 14.752 11.372 ;
  LAYER M2 ;
        RECT 12.352 11.404 12.384 11.436 ;
  LAYER M2 ;
        RECT 14.72 11.468 14.752 11.5 ;
  LAYER M2 ;
        RECT 12.352 11.532 12.384 11.564 ;
  LAYER M2 ;
        RECT 14.72 11.596 14.752 11.628 ;
  LAYER M2 ;
        RECT 12.352 11.66 12.384 11.692 ;
  LAYER M2 ;
        RECT 14.72 11.724 14.752 11.756 ;
  LAYER M2 ;
        RECT 12.352 11.788 12.384 11.82 ;
  LAYER M2 ;
        RECT 14.72 11.852 14.752 11.884 ;
  LAYER M2 ;
        RECT 12.352 11.916 12.384 11.948 ;
  LAYER M2 ;
        RECT 14.72 11.98 14.752 12.012 ;
  LAYER M2 ;
        RECT 12.352 12.044 12.384 12.076 ;
  LAYER M2 ;
        RECT 14.72 12.108 14.752 12.14 ;
  LAYER M2 ;
        RECT 12.352 12.172 12.384 12.204 ;
  LAYER M2 ;
        RECT 14.72 12.236 14.752 12.268 ;
  LAYER M2 ;
        RECT 12.352 12.3 12.384 12.332 ;
  LAYER M2 ;
        RECT 14.72 12.364 14.752 12.396 ;
  LAYER M2 ;
        RECT 12.352 12.428 12.384 12.46 ;
  LAYER M2 ;
        RECT 14.72 12.492 14.752 12.524 ;
  LAYER M2 ;
        RECT 12.352 12.556 12.384 12.588 ;
  LAYER M2 ;
        RECT 14.72 12.62 14.752 12.652 ;
  LAYER M2 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M1 ;
        RECT 12.352 13.404 12.384 15.912 ;
  LAYER M3 ;
        RECT 12.352 15.86 12.384 15.892 ;
  LAYER M1 ;
        RECT 12.416 13.404 12.448 15.912 ;
  LAYER M3 ;
        RECT 12.416 13.424 12.448 13.456 ;
  LAYER M1 ;
        RECT 12.48 13.404 12.512 15.912 ;
  LAYER M3 ;
        RECT 12.48 15.86 12.512 15.892 ;
  LAYER M1 ;
        RECT 12.544 13.404 12.576 15.912 ;
  LAYER M3 ;
        RECT 12.544 13.424 12.576 13.456 ;
  LAYER M1 ;
        RECT 12.608 13.404 12.64 15.912 ;
  LAYER M3 ;
        RECT 12.608 15.86 12.64 15.892 ;
  LAYER M1 ;
        RECT 12.672 13.404 12.704 15.912 ;
  LAYER M3 ;
        RECT 12.672 13.424 12.704 13.456 ;
  LAYER M1 ;
        RECT 12.736 13.404 12.768 15.912 ;
  LAYER M3 ;
        RECT 12.736 15.86 12.768 15.892 ;
  LAYER M1 ;
        RECT 12.8 13.404 12.832 15.912 ;
  LAYER M3 ;
        RECT 12.8 13.424 12.832 13.456 ;
  LAYER M1 ;
        RECT 12.864 13.404 12.896 15.912 ;
  LAYER M3 ;
        RECT 12.864 15.86 12.896 15.892 ;
  LAYER M1 ;
        RECT 12.928 13.404 12.96 15.912 ;
  LAYER M3 ;
        RECT 12.928 13.424 12.96 13.456 ;
  LAYER M1 ;
        RECT 12.992 13.404 13.024 15.912 ;
  LAYER M3 ;
        RECT 12.992 15.86 13.024 15.892 ;
  LAYER M1 ;
        RECT 13.056 13.404 13.088 15.912 ;
  LAYER M3 ;
        RECT 13.056 13.424 13.088 13.456 ;
  LAYER M1 ;
        RECT 13.12 13.404 13.152 15.912 ;
  LAYER M3 ;
        RECT 13.12 15.86 13.152 15.892 ;
  LAYER M1 ;
        RECT 13.184 13.404 13.216 15.912 ;
  LAYER M3 ;
        RECT 13.184 13.424 13.216 13.456 ;
  LAYER M1 ;
        RECT 13.248 13.404 13.28 15.912 ;
  LAYER M3 ;
        RECT 13.248 15.86 13.28 15.892 ;
  LAYER M1 ;
        RECT 13.312 13.404 13.344 15.912 ;
  LAYER M3 ;
        RECT 13.312 13.424 13.344 13.456 ;
  LAYER M1 ;
        RECT 13.376 13.404 13.408 15.912 ;
  LAYER M3 ;
        RECT 13.376 15.86 13.408 15.892 ;
  LAYER M1 ;
        RECT 13.44 13.404 13.472 15.912 ;
  LAYER M3 ;
        RECT 13.44 13.424 13.472 13.456 ;
  LAYER M1 ;
        RECT 13.504 13.404 13.536 15.912 ;
  LAYER M3 ;
        RECT 13.504 15.86 13.536 15.892 ;
  LAYER M1 ;
        RECT 13.568 13.404 13.6 15.912 ;
  LAYER M3 ;
        RECT 13.568 13.424 13.6 13.456 ;
  LAYER M1 ;
        RECT 13.632 13.404 13.664 15.912 ;
  LAYER M3 ;
        RECT 13.632 15.86 13.664 15.892 ;
  LAYER M1 ;
        RECT 13.696 13.404 13.728 15.912 ;
  LAYER M3 ;
        RECT 13.696 13.424 13.728 13.456 ;
  LAYER M1 ;
        RECT 13.76 13.404 13.792 15.912 ;
  LAYER M3 ;
        RECT 13.76 15.86 13.792 15.892 ;
  LAYER M1 ;
        RECT 13.824 13.404 13.856 15.912 ;
  LAYER M3 ;
        RECT 13.824 13.424 13.856 13.456 ;
  LAYER M1 ;
        RECT 13.888 13.404 13.92 15.912 ;
  LAYER M3 ;
        RECT 13.888 15.86 13.92 15.892 ;
  LAYER M1 ;
        RECT 13.952 13.404 13.984 15.912 ;
  LAYER M3 ;
        RECT 13.952 13.424 13.984 13.456 ;
  LAYER M1 ;
        RECT 14.016 13.404 14.048 15.912 ;
  LAYER M3 ;
        RECT 14.016 15.86 14.048 15.892 ;
  LAYER M1 ;
        RECT 14.08 13.404 14.112 15.912 ;
  LAYER M3 ;
        RECT 14.08 13.424 14.112 13.456 ;
  LAYER M1 ;
        RECT 14.144 13.404 14.176 15.912 ;
  LAYER M3 ;
        RECT 14.144 15.86 14.176 15.892 ;
  LAYER M1 ;
        RECT 14.208 13.404 14.24 15.912 ;
  LAYER M3 ;
        RECT 14.208 13.424 14.24 13.456 ;
  LAYER M1 ;
        RECT 14.272 13.404 14.304 15.912 ;
  LAYER M3 ;
        RECT 14.272 15.86 14.304 15.892 ;
  LAYER M1 ;
        RECT 14.336 13.404 14.368 15.912 ;
  LAYER M3 ;
        RECT 14.336 13.424 14.368 13.456 ;
  LAYER M1 ;
        RECT 14.4 13.404 14.432 15.912 ;
  LAYER M3 ;
        RECT 14.4 15.86 14.432 15.892 ;
  LAYER M1 ;
        RECT 14.464 13.404 14.496 15.912 ;
  LAYER M3 ;
        RECT 14.464 13.424 14.496 13.456 ;
  LAYER M1 ;
        RECT 14.528 13.404 14.56 15.912 ;
  LAYER M3 ;
        RECT 14.528 15.86 14.56 15.892 ;
  LAYER M1 ;
        RECT 14.592 13.404 14.624 15.912 ;
  LAYER M3 ;
        RECT 14.592 13.424 14.624 13.456 ;
  LAYER M1 ;
        RECT 14.656 13.404 14.688 15.912 ;
  LAYER M3 ;
        RECT 14.656 15.86 14.688 15.892 ;
  LAYER M1 ;
        RECT 14.72 13.404 14.752 15.912 ;
  LAYER M3 ;
        RECT 12.352 13.488 12.384 13.52 ;
  LAYER M2 ;
        RECT 14.72 13.552 14.752 13.584 ;
  LAYER M2 ;
        RECT 12.352 13.616 12.384 13.648 ;
  LAYER M2 ;
        RECT 14.72 13.68 14.752 13.712 ;
  LAYER M2 ;
        RECT 12.352 13.744 12.384 13.776 ;
  LAYER M2 ;
        RECT 14.72 13.808 14.752 13.84 ;
  LAYER M2 ;
        RECT 12.352 13.872 12.384 13.904 ;
  LAYER M2 ;
        RECT 14.72 13.936 14.752 13.968 ;
  LAYER M2 ;
        RECT 12.352 14 12.384 14.032 ;
  LAYER M2 ;
        RECT 14.72 14.064 14.752 14.096 ;
  LAYER M2 ;
        RECT 12.352 14.128 12.384 14.16 ;
  LAYER M2 ;
        RECT 14.72 14.192 14.752 14.224 ;
  LAYER M2 ;
        RECT 12.352 14.256 12.384 14.288 ;
  LAYER M2 ;
        RECT 14.72 14.32 14.752 14.352 ;
  LAYER M2 ;
        RECT 12.352 14.384 12.384 14.416 ;
  LAYER M2 ;
        RECT 14.72 14.448 14.752 14.48 ;
  LAYER M2 ;
        RECT 12.352 14.512 12.384 14.544 ;
  LAYER M2 ;
        RECT 14.72 14.576 14.752 14.608 ;
  LAYER M2 ;
        RECT 12.352 14.64 12.384 14.672 ;
  LAYER M2 ;
        RECT 14.72 14.704 14.752 14.736 ;
  LAYER M2 ;
        RECT 12.352 14.768 12.384 14.8 ;
  LAYER M2 ;
        RECT 14.72 14.832 14.752 14.864 ;
  LAYER M2 ;
        RECT 12.352 14.896 12.384 14.928 ;
  LAYER M2 ;
        RECT 14.72 14.96 14.752 14.992 ;
  LAYER M2 ;
        RECT 12.352 15.024 12.384 15.056 ;
  LAYER M2 ;
        RECT 14.72 15.088 14.752 15.12 ;
  LAYER M2 ;
        RECT 12.352 15.152 12.384 15.184 ;
  LAYER M2 ;
        RECT 14.72 15.216 14.752 15.248 ;
  LAYER M2 ;
        RECT 12.352 15.28 12.384 15.312 ;
  LAYER M2 ;
        RECT 14.72 15.344 14.752 15.376 ;
  LAYER M2 ;
        RECT 12.352 15.408 12.384 15.44 ;
  LAYER M2 ;
        RECT 14.72 15.472 14.752 15.504 ;
  LAYER M2 ;
        RECT 12.352 15.536 12.384 15.568 ;
  LAYER M2 ;
        RECT 14.72 15.6 14.752 15.632 ;
  LAYER M2 ;
        RECT 12.352 15.664 12.384 15.696 ;
  LAYER M2 ;
        RECT 14.72 15.728 14.752 15.76 ;
  LAYER M2 ;
        RECT 12.304 13.356 14.8 15.96 ;
  LAYER M1 ;
        RECT 15.328 0.972 15.36 3.48 ;
  LAYER M3 ;
        RECT 15.328 3.428 15.36 3.46 ;
  LAYER M1 ;
        RECT 15.392 0.972 15.424 3.48 ;
  LAYER M3 ;
        RECT 15.392 0.992 15.424 1.024 ;
  LAYER M1 ;
        RECT 15.456 0.972 15.488 3.48 ;
  LAYER M3 ;
        RECT 15.456 3.428 15.488 3.46 ;
  LAYER M1 ;
        RECT 15.52 0.972 15.552 3.48 ;
  LAYER M3 ;
        RECT 15.52 0.992 15.552 1.024 ;
  LAYER M1 ;
        RECT 15.584 0.972 15.616 3.48 ;
  LAYER M3 ;
        RECT 15.584 3.428 15.616 3.46 ;
  LAYER M1 ;
        RECT 15.648 0.972 15.68 3.48 ;
  LAYER M3 ;
        RECT 15.648 0.992 15.68 1.024 ;
  LAYER M1 ;
        RECT 15.712 0.972 15.744 3.48 ;
  LAYER M3 ;
        RECT 15.712 3.428 15.744 3.46 ;
  LAYER M1 ;
        RECT 15.776 0.972 15.808 3.48 ;
  LAYER M3 ;
        RECT 15.776 0.992 15.808 1.024 ;
  LAYER M1 ;
        RECT 15.84 0.972 15.872 3.48 ;
  LAYER M3 ;
        RECT 15.84 3.428 15.872 3.46 ;
  LAYER M1 ;
        RECT 15.904 0.972 15.936 3.48 ;
  LAYER M3 ;
        RECT 15.904 0.992 15.936 1.024 ;
  LAYER M1 ;
        RECT 15.968 0.972 16 3.48 ;
  LAYER M3 ;
        RECT 15.968 3.428 16 3.46 ;
  LAYER M1 ;
        RECT 16.032 0.972 16.064 3.48 ;
  LAYER M3 ;
        RECT 16.032 0.992 16.064 1.024 ;
  LAYER M1 ;
        RECT 16.096 0.972 16.128 3.48 ;
  LAYER M3 ;
        RECT 16.096 3.428 16.128 3.46 ;
  LAYER M1 ;
        RECT 16.16 0.972 16.192 3.48 ;
  LAYER M3 ;
        RECT 16.16 0.992 16.192 1.024 ;
  LAYER M1 ;
        RECT 16.224 0.972 16.256 3.48 ;
  LAYER M3 ;
        RECT 16.224 3.428 16.256 3.46 ;
  LAYER M1 ;
        RECT 16.288 0.972 16.32 3.48 ;
  LAYER M3 ;
        RECT 16.288 0.992 16.32 1.024 ;
  LAYER M1 ;
        RECT 16.352 0.972 16.384 3.48 ;
  LAYER M3 ;
        RECT 16.352 3.428 16.384 3.46 ;
  LAYER M1 ;
        RECT 16.416 0.972 16.448 3.48 ;
  LAYER M3 ;
        RECT 16.416 0.992 16.448 1.024 ;
  LAYER M1 ;
        RECT 16.48 0.972 16.512 3.48 ;
  LAYER M3 ;
        RECT 16.48 3.428 16.512 3.46 ;
  LAYER M1 ;
        RECT 16.544 0.972 16.576 3.48 ;
  LAYER M3 ;
        RECT 16.544 0.992 16.576 1.024 ;
  LAYER M1 ;
        RECT 16.608 0.972 16.64 3.48 ;
  LAYER M3 ;
        RECT 16.608 3.428 16.64 3.46 ;
  LAYER M1 ;
        RECT 16.672 0.972 16.704 3.48 ;
  LAYER M3 ;
        RECT 16.672 0.992 16.704 1.024 ;
  LAYER M1 ;
        RECT 16.736 0.972 16.768 3.48 ;
  LAYER M3 ;
        RECT 16.736 3.428 16.768 3.46 ;
  LAYER M1 ;
        RECT 16.8 0.972 16.832 3.48 ;
  LAYER M3 ;
        RECT 16.8 0.992 16.832 1.024 ;
  LAYER M1 ;
        RECT 16.864 0.972 16.896 3.48 ;
  LAYER M3 ;
        RECT 16.864 3.428 16.896 3.46 ;
  LAYER M1 ;
        RECT 16.928 0.972 16.96 3.48 ;
  LAYER M3 ;
        RECT 16.928 0.992 16.96 1.024 ;
  LAYER M1 ;
        RECT 16.992 0.972 17.024 3.48 ;
  LAYER M3 ;
        RECT 16.992 3.428 17.024 3.46 ;
  LAYER M1 ;
        RECT 17.056 0.972 17.088 3.48 ;
  LAYER M3 ;
        RECT 17.056 0.992 17.088 1.024 ;
  LAYER M1 ;
        RECT 17.12 0.972 17.152 3.48 ;
  LAYER M3 ;
        RECT 17.12 3.428 17.152 3.46 ;
  LAYER M1 ;
        RECT 17.184 0.972 17.216 3.48 ;
  LAYER M3 ;
        RECT 17.184 0.992 17.216 1.024 ;
  LAYER M1 ;
        RECT 17.248 0.972 17.28 3.48 ;
  LAYER M3 ;
        RECT 17.248 3.428 17.28 3.46 ;
  LAYER M1 ;
        RECT 17.312 0.972 17.344 3.48 ;
  LAYER M3 ;
        RECT 17.312 0.992 17.344 1.024 ;
  LAYER M1 ;
        RECT 17.376 0.972 17.408 3.48 ;
  LAYER M3 ;
        RECT 17.376 3.428 17.408 3.46 ;
  LAYER M1 ;
        RECT 17.44 0.972 17.472 3.48 ;
  LAYER M3 ;
        RECT 17.44 0.992 17.472 1.024 ;
  LAYER M1 ;
        RECT 17.504 0.972 17.536 3.48 ;
  LAYER M3 ;
        RECT 17.504 3.428 17.536 3.46 ;
  LAYER M1 ;
        RECT 17.568 0.972 17.6 3.48 ;
  LAYER M3 ;
        RECT 17.568 0.992 17.6 1.024 ;
  LAYER M1 ;
        RECT 17.632 0.972 17.664 3.48 ;
  LAYER M3 ;
        RECT 17.632 3.428 17.664 3.46 ;
  LAYER M1 ;
        RECT 17.696 0.972 17.728 3.48 ;
  LAYER M3 ;
        RECT 15.328 1.056 15.36 1.088 ;
  LAYER M2 ;
        RECT 17.696 1.12 17.728 1.152 ;
  LAYER M2 ;
        RECT 15.328 1.184 15.36 1.216 ;
  LAYER M2 ;
        RECT 17.696 1.248 17.728 1.28 ;
  LAYER M2 ;
        RECT 15.328 1.312 15.36 1.344 ;
  LAYER M2 ;
        RECT 17.696 1.376 17.728 1.408 ;
  LAYER M2 ;
        RECT 15.328 1.44 15.36 1.472 ;
  LAYER M2 ;
        RECT 17.696 1.504 17.728 1.536 ;
  LAYER M2 ;
        RECT 15.328 1.568 15.36 1.6 ;
  LAYER M2 ;
        RECT 17.696 1.632 17.728 1.664 ;
  LAYER M2 ;
        RECT 15.328 1.696 15.36 1.728 ;
  LAYER M2 ;
        RECT 17.696 1.76 17.728 1.792 ;
  LAYER M2 ;
        RECT 15.328 1.824 15.36 1.856 ;
  LAYER M2 ;
        RECT 17.696 1.888 17.728 1.92 ;
  LAYER M2 ;
        RECT 15.328 1.952 15.36 1.984 ;
  LAYER M2 ;
        RECT 17.696 2.016 17.728 2.048 ;
  LAYER M2 ;
        RECT 15.328 2.08 15.36 2.112 ;
  LAYER M2 ;
        RECT 17.696 2.144 17.728 2.176 ;
  LAYER M2 ;
        RECT 15.328 2.208 15.36 2.24 ;
  LAYER M2 ;
        RECT 17.696 2.272 17.728 2.304 ;
  LAYER M2 ;
        RECT 15.328 2.336 15.36 2.368 ;
  LAYER M2 ;
        RECT 17.696 2.4 17.728 2.432 ;
  LAYER M2 ;
        RECT 15.328 2.464 15.36 2.496 ;
  LAYER M2 ;
        RECT 17.696 2.528 17.728 2.56 ;
  LAYER M2 ;
        RECT 15.328 2.592 15.36 2.624 ;
  LAYER M2 ;
        RECT 17.696 2.656 17.728 2.688 ;
  LAYER M2 ;
        RECT 15.328 2.72 15.36 2.752 ;
  LAYER M2 ;
        RECT 17.696 2.784 17.728 2.816 ;
  LAYER M2 ;
        RECT 15.328 2.848 15.36 2.88 ;
  LAYER M2 ;
        RECT 17.696 2.912 17.728 2.944 ;
  LAYER M2 ;
        RECT 15.328 2.976 15.36 3.008 ;
  LAYER M2 ;
        RECT 17.696 3.04 17.728 3.072 ;
  LAYER M2 ;
        RECT 15.328 3.104 15.36 3.136 ;
  LAYER M2 ;
        RECT 17.696 3.168 17.728 3.2 ;
  LAYER M2 ;
        RECT 15.328 3.232 15.36 3.264 ;
  LAYER M2 ;
        RECT 17.696 3.296 17.728 3.328 ;
  LAYER M2 ;
        RECT 15.28 0.924 17.776 3.528 ;
  LAYER M1 ;
        RECT 15.328 4.08 15.36 6.588 ;
  LAYER M3 ;
        RECT 15.328 6.536 15.36 6.568 ;
  LAYER M1 ;
        RECT 15.392 4.08 15.424 6.588 ;
  LAYER M3 ;
        RECT 15.392 4.1 15.424 4.132 ;
  LAYER M1 ;
        RECT 15.456 4.08 15.488 6.588 ;
  LAYER M3 ;
        RECT 15.456 6.536 15.488 6.568 ;
  LAYER M1 ;
        RECT 15.52 4.08 15.552 6.588 ;
  LAYER M3 ;
        RECT 15.52 4.1 15.552 4.132 ;
  LAYER M1 ;
        RECT 15.584 4.08 15.616 6.588 ;
  LAYER M3 ;
        RECT 15.584 6.536 15.616 6.568 ;
  LAYER M1 ;
        RECT 15.648 4.08 15.68 6.588 ;
  LAYER M3 ;
        RECT 15.648 4.1 15.68 4.132 ;
  LAYER M1 ;
        RECT 15.712 4.08 15.744 6.588 ;
  LAYER M3 ;
        RECT 15.712 6.536 15.744 6.568 ;
  LAYER M1 ;
        RECT 15.776 4.08 15.808 6.588 ;
  LAYER M3 ;
        RECT 15.776 4.1 15.808 4.132 ;
  LAYER M1 ;
        RECT 15.84 4.08 15.872 6.588 ;
  LAYER M3 ;
        RECT 15.84 6.536 15.872 6.568 ;
  LAYER M1 ;
        RECT 15.904 4.08 15.936 6.588 ;
  LAYER M3 ;
        RECT 15.904 4.1 15.936 4.132 ;
  LAYER M1 ;
        RECT 15.968 4.08 16 6.588 ;
  LAYER M3 ;
        RECT 15.968 6.536 16 6.568 ;
  LAYER M1 ;
        RECT 16.032 4.08 16.064 6.588 ;
  LAYER M3 ;
        RECT 16.032 4.1 16.064 4.132 ;
  LAYER M1 ;
        RECT 16.096 4.08 16.128 6.588 ;
  LAYER M3 ;
        RECT 16.096 6.536 16.128 6.568 ;
  LAYER M1 ;
        RECT 16.16 4.08 16.192 6.588 ;
  LAYER M3 ;
        RECT 16.16 4.1 16.192 4.132 ;
  LAYER M1 ;
        RECT 16.224 4.08 16.256 6.588 ;
  LAYER M3 ;
        RECT 16.224 6.536 16.256 6.568 ;
  LAYER M1 ;
        RECT 16.288 4.08 16.32 6.588 ;
  LAYER M3 ;
        RECT 16.288 4.1 16.32 4.132 ;
  LAYER M1 ;
        RECT 16.352 4.08 16.384 6.588 ;
  LAYER M3 ;
        RECT 16.352 6.536 16.384 6.568 ;
  LAYER M1 ;
        RECT 16.416 4.08 16.448 6.588 ;
  LAYER M3 ;
        RECT 16.416 4.1 16.448 4.132 ;
  LAYER M1 ;
        RECT 16.48 4.08 16.512 6.588 ;
  LAYER M3 ;
        RECT 16.48 6.536 16.512 6.568 ;
  LAYER M1 ;
        RECT 16.544 4.08 16.576 6.588 ;
  LAYER M3 ;
        RECT 16.544 4.1 16.576 4.132 ;
  LAYER M1 ;
        RECT 16.608 4.08 16.64 6.588 ;
  LAYER M3 ;
        RECT 16.608 6.536 16.64 6.568 ;
  LAYER M1 ;
        RECT 16.672 4.08 16.704 6.588 ;
  LAYER M3 ;
        RECT 16.672 4.1 16.704 4.132 ;
  LAYER M1 ;
        RECT 16.736 4.08 16.768 6.588 ;
  LAYER M3 ;
        RECT 16.736 6.536 16.768 6.568 ;
  LAYER M1 ;
        RECT 16.8 4.08 16.832 6.588 ;
  LAYER M3 ;
        RECT 16.8 4.1 16.832 4.132 ;
  LAYER M1 ;
        RECT 16.864 4.08 16.896 6.588 ;
  LAYER M3 ;
        RECT 16.864 6.536 16.896 6.568 ;
  LAYER M1 ;
        RECT 16.928 4.08 16.96 6.588 ;
  LAYER M3 ;
        RECT 16.928 4.1 16.96 4.132 ;
  LAYER M1 ;
        RECT 16.992 4.08 17.024 6.588 ;
  LAYER M3 ;
        RECT 16.992 6.536 17.024 6.568 ;
  LAYER M1 ;
        RECT 17.056 4.08 17.088 6.588 ;
  LAYER M3 ;
        RECT 17.056 4.1 17.088 4.132 ;
  LAYER M1 ;
        RECT 17.12 4.08 17.152 6.588 ;
  LAYER M3 ;
        RECT 17.12 6.536 17.152 6.568 ;
  LAYER M1 ;
        RECT 17.184 4.08 17.216 6.588 ;
  LAYER M3 ;
        RECT 17.184 4.1 17.216 4.132 ;
  LAYER M1 ;
        RECT 17.248 4.08 17.28 6.588 ;
  LAYER M3 ;
        RECT 17.248 6.536 17.28 6.568 ;
  LAYER M1 ;
        RECT 17.312 4.08 17.344 6.588 ;
  LAYER M3 ;
        RECT 17.312 4.1 17.344 4.132 ;
  LAYER M1 ;
        RECT 17.376 4.08 17.408 6.588 ;
  LAYER M3 ;
        RECT 17.376 6.536 17.408 6.568 ;
  LAYER M1 ;
        RECT 17.44 4.08 17.472 6.588 ;
  LAYER M3 ;
        RECT 17.44 4.1 17.472 4.132 ;
  LAYER M1 ;
        RECT 17.504 4.08 17.536 6.588 ;
  LAYER M3 ;
        RECT 17.504 6.536 17.536 6.568 ;
  LAYER M1 ;
        RECT 17.568 4.08 17.6 6.588 ;
  LAYER M3 ;
        RECT 17.568 4.1 17.6 4.132 ;
  LAYER M1 ;
        RECT 17.632 4.08 17.664 6.588 ;
  LAYER M3 ;
        RECT 17.632 6.536 17.664 6.568 ;
  LAYER M1 ;
        RECT 17.696 4.08 17.728 6.588 ;
  LAYER M3 ;
        RECT 15.328 4.164 15.36 4.196 ;
  LAYER M2 ;
        RECT 17.696 4.228 17.728 4.26 ;
  LAYER M2 ;
        RECT 15.328 4.292 15.36 4.324 ;
  LAYER M2 ;
        RECT 17.696 4.356 17.728 4.388 ;
  LAYER M2 ;
        RECT 15.328 4.42 15.36 4.452 ;
  LAYER M2 ;
        RECT 17.696 4.484 17.728 4.516 ;
  LAYER M2 ;
        RECT 15.328 4.548 15.36 4.58 ;
  LAYER M2 ;
        RECT 17.696 4.612 17.728 4.644 ;
  LAYER M2 ;
        RECT 15.328 4.676 15.36 4.708 ;
  LAYER M2 ;
        RECT 17.696 4.74 17.728 4.772 ;
  LAYER M2 ;
        RECT 15.328 4.804 15.36 4.836 ;
  LAYER M2 ;
        RECT 17.696 4.868 17.728 4.9 ;
  LAYER M2 ;
        RECT 15.328 4.932 15.36 4.964 ;
  LAYER M2 ;
        RECT 17.696 4.996 17.728 5.028 ;
  LAYER M2 ;
        RECT 15.328 5.06 15.36 5.092 ;
  LAYER M2 ;
        RECT 17.696 5.124 17.728 5.156 ;
  LAYER M2 ;
        RECT 15.328 5.188 15.36 5.22 ;
  LAYER M2 ;
        RECT 17.696 5.252 17.728 5.284 ;
  LAYER M2 ;
        RECT 15.328 5.316 15.36 5.348 ;
  LAYER M2 ;
        RECT 17.696 5.38 17.728 5.412 ;
  LAYER M2 ;
        RECT 15.328 5.444 15.36 5.476 ;
  LAYER M2 ;
        RECT 17.696 5.508 17.728 5.54 ;
  LAYER M2 ;
        RECT 15.328 5.572 15.36 5.604 ;
  LAYER M2 ;
        RECT 17.696 5.636 17.728 5.668 ;
  LAYER M2 ;
        RECT 15.328 5.7 15.36 5.732 ;
  LAYER M2 ;
        RECT 17.696 5.764 17.728 5.796 ;
  LAYER M2 ;
        RECT 15.328 5.828 15.36 5.86 ;
  LAYER M2 ;
        RECT 17.696 5.892 17.728 5.924 ;
  LAYER M2 ;
        RECT 15.328 5.956 15.36 5.988 ;
  LAYER M2 ;
        RECT 17.696 6.02 17.728 6.052 ;
  LAYER M2 ;
        RECT 15.328 6.084 15.36 6.116 ;
  LAYER M2 ;
        RECT 17.696 6.148 17.728 6.18 ;
  LAYER M2 ;
        RECT 15.328 6.212 15.36 6.244 ;
  LAYER M2 ;
        RECT 17.696 6.276 17.728 6.308 ;
  LAYER M2 ;
        RECT 15.328 6.34 15.36 6.372 ;
  LAYER M2 ;
        RECT 17.696 6.404 17.728 6.436 ;
  LAYER M2 ;
        RECT 15.28 4.032 17.776 6.636 ;
  LAYER M1 ;
        RECT 15.328 7.188 15.36 9.696 ;
  LAYER M3 ;
        RECT 15.328 9.644 15.36 9.676 ;
  LAYER M1 ;
        RECT 15.392 7.188 15.424 9.696 ;
  LAYER M3 ;
        RECT 15.392 7.208 15.424 7.24 ;
  LAYER M1 ;
        RECT 15.456 7.188 15.488 9.696 ;
  LAYER M3 ;
        RECT 15.456 9.644 15.488 9.676 ;
  LAYER M1 ;
        RECT 15.52 7.188 15.552 9.696 ;
  LAYER M3 ;
        RECT 15.52 7.208 15.552 7.24 ;
  LAYER M1 ;
        RECT 15.584 7.188 15.616 9.696 ;
  LAYER M3 ;
        RECT 15.584 9.644 15.616 9.676 ;
  LAYER M1 ;
        RECT 15.648 7.188 15.68 9.696 ;
  LAYER M3 ;
        RECT 15.648 7.208 15.68 7.24 ;
  LAYER M1 ;
        RECT 15.712 7.188 15.744 9.696 ;
  LAYER M3 ;
        RECT 15.712 9.644 15.744 9.676 ;
  LAYER M1 ;
        RECT 15.776 7.188 15.808 9.696 ;
  LAYER M3 ;
        RECT 15.776 7.208 15.808 7.24 ;
  LAYER M1 ;
        RECT 15.84 7.188 15.872 9.696 ;
  LAYER M3 ;
        RECT 15.84 9.644 15.872 9.676 ;
  LAYER M1 ;
        RECT 15.904 7.188 15.936 9.696 ;
  LAYER M3 ;
        RECT 15.904 7.208 15.936 7.24 ;
  LAYER M1 ;
        RECT 15.968 7.188 16 9.696 ;
  LAYER M3 ;
        RECT 15.968 9.644 16 9.676 ;
  LAYER M1 ;
        RECT 16.032 7.188 16.064 9.696 ;
  LAYER M3 ;
        RECT 16.032 7.208 16.064 7.24 ;
  LAYER M1 ;
        RECT 16.096 7.188 16.128 9.696 ;
  LAYER M3 ;
        RECT 16.096 9.644 16.128 9.676 ;
  LAYER M1 ;
        RECT 16.16 7.188 16.192 9.696 ;
  LAYER M3 ;
        RECT 16.16 7.208 16.192 7.24 ;
  LAYER M1 ;
        RECT 16.224 7.188 16.256 9.696 ;
  LAYER M3 ;
        RECT 16.224 9.644 16.256 9.676 ;
  LAYER M1 ;
        RECT 16.288 7.188 16.32 9.696 ;
  LAYER M3 ;
        RECT 16.288 7.208 16.32 7.24 ;
  LAYER M1 ;
        RECT 16.352 7.188 16.384 9.696 ;
  LAYER M3 ;
        RECT 16.352 9.644 16.384 9.676 ;
  LAYER M1 ;
        RECT 16.416 7.188 16.448 9.696 ;
  LAYER M3 ;
        RECT 16.416 7.208 16.448 7.24 ;
  LAYER M1 ;
        RECT 16.48 7.188 16.512 9.696 ;
  LAYER M3 ;
        RECT 16.48 9.644 16.512 9.676 ;
  LAYER M1 ;
        RECT 16.544 7.188 16.576 9.696 ;
  LAYER M3 ;
        RECT 16.544 7.208 16.576 7.24 ;
  LAYER M1 ;
        RECT 16.608 7.188 16.64 9.696 ;
  LAYER M3 ;
        RECT 16.608 9.644 16.64 9.676 ;
  LAYER M1 ;
        RECT 16.672 7.188 16.704 9.696 ;
  LAYER M3 ;
        RECT 16.672 7.208 16.704 7.24 ;
  LAYER M1 ;
        RECT 16.736 7.188 16.768 9.696 ;
  LAYER M3 ;
        RECT 16.736 9.644 16.768 9.676 ;
  LAYER M1 ;
        RECT 16.8 7.188 16.832 9.696 ;
  LAYER M3 ;
        RECT 16.8 7.208 16.832 7.24 ;
  LAYER M1 ;
        RECT 16.864 7.188 16.896 9.696 ;
  LAYER M3 ;
        RECT 16.864 9.644 16.896 9.676 ;
  LAYER M1 ;
        RECT 16.928 7.188 16.96 9.696 ;
  LAYER M3 ;
        RECT 16.928 7.208 16.96 7.24 ;
  LAYER M1 ;
        RECT 16.992 7.188 17.024 9.696 ;
  LAYER M3 ;
        RECT 16.992 9.644 17.024 9.676 ;
  LAYER M1 ;
        RECT 17.056 7.188 17.088 9.696 ;
  LAYER M3 ;
        RECT 17.056 7.208 17.088 7.24 ;
  LAYER M1 ;
        RECT 17.12 7.188 17.152 9.696 ;
  LAYER M3 ;
        RECT 17.12 9.644 17.152 9.676 ;
  LAYER M1 ;
        RECT 17.184 7.188 17.216 9.696 ;
  LAYER M3 ;
        RECT 17.184 7.208 17.216 7.24 ;
  LAYER M1 ;
        RECT 17.248 7.188 17.28 9.696 ;
  LAYER M3 ;
        RECT 17.248 9.644 17.28 9.676 ;
  LAYER M1 ;
        RECT 17.312 7.188 17.344 9.696 ;
  LAYER M3 ;
        RECT 17.312 7.208 17.344 7.24 ;
  LAYER M1 ;
        RECT 17.376 7.188 17.408 9.696 ;
  LAYER M3 ;
        RECT 17.376 9.644 17.408 9.676 ;
  LAYER M1 ;
        RECT 17.44 7.188 17.472 9.696 ;
  LAYER M3 ;
        RECT 17.44 7.208 17.472 7.24 ;
  LAYER M1 ;
        RECT 17.504 7.188 17.536 9.696 ;
  LAYER M3 ;
        RECT 17.504 9.644 17.536 9.676 ;
  LAYER M1 ;
        RECT 17.568 7.188 17.6 9.696 ;
  LAYER M3 ;
        RECT 17.568 7.208 17.6 7.24 ;
  LAYER M1 ;
        RECT 17.632 7.188 17.664 9.696 ;
  LAYER M3 ;
        RECT 17.632 9.644 17.664 9.676 ;
  LAYER M1 ;
        RECT 17.696 7.188 17.728 9.696 ;
  LAYER M3 ;
        RECT 15.328 7.272 15.36 7.304 ;
  LAYER M2 ;
        RECT 17.696 7.336 17.728 7.368 ;
  LAYER M2 ;
        RECT 15.328 7.4 15.36 7.432 ;
  LAYER M2 ;
        RECT 17.696 7.464 17.728 7.496 ;
  LAYER M2 ;
        RECT 15.328 7.528 15.36 7.56 ;
  LAYER M2 ;
        RECT 17.696 7.592 17.728 7.624 ;
  LAYER M2 ;
        RECT 15.328 7.656 15.36 7.688 ;
  LAYER M2 ;
        RECT 17.696 7.72 17.728 7.752 ;
  LAYER M2 ;
        RECT 15.328 7.784 15.36 7.816 ;
  LAYER M2 ;
        RECT 17.696 7.848 17.728 7.88 ;
  LAYER M2 ;
        RECT 15.328 7.912 15.36 7.944 ;
  LAYER M2 ;
        RECT 17.696 7.976 17.728 8.008 ;
  LAYER M2 ;
        RECT 15.328 8.04 15.36 8.072 ;
  LAYER M2 ;
        RECT 17.696 8.104 17.728 8.136 ;
  LAYER M2 ;
        RECT 15.328 8.168 15.36 8.2 ;
  LAYER M2 ;
        RECT 17.696 8.232 17.728 8.264 ;
  LAYER M2 ;
        RECT 15.328 8.296 15.36 8.328 ;
  LAYER M2 ;
        RECT 17.696 8.36 17.728 8.392 ;
  LAYER M2 ;
        RECT 15.328 8.424 15.36 8.456 ;
  LAYER M2 ;
        RECT 17.696 8.488 17.728 8.52 ;
  LAYER M2 ;
        RECT 15.328 8.552 15.36 8.584 ;
  LAYER M2 ;
        RECT 17.696 8.616 17.728 8.648 ;
  LAYER M2 ;
        RECT 15.328 8.68 15.36 8.712 ;
  LAYER M2 ;
        RECT 17.696 8.744 17.728 8.776 ;
  LAYER M2 ;
        RECT 15.328 8.808 15.36 8.84 ;
  LAYER M2 ;
        RECT 17.696 8.872 17.728 8.904 ;
  LAYER M2 ;
        RECT 15.328 8.936 15.36 8.968 ;
  LAYER M2 ;
        RECT 17.696 9 17.728 9.032 ;
  LAYER M2 ;
        RECT 15.328 9.064 15.36 9.096 ;
  LAYER M2 ;
        RECT 17.696 9.128 17.728 9.16 ;
  LAYER M2 ;
        RECT 15.328 9.192 15.36 9.224 ;
  LAYER M2 ;
        RECT 17.696 9.256 17.728 9.288 ;
  LAYER M2 ;
        RECT 15.328 9.32 15.36 9.352 ;
  LAYER M2 ;
        RECT 17.696 9.384 17.728 9.416 ;
  LAYER M2 ;
        RECT 15.328 9.448 15.36 9.48 ;
  LAYER M2 ;
        RECT 17.696 9.512 17.728 9.544 ;
  LAYER M2 ;
        RECT 15.28 7.14 17.776 9.744 ;
  LAYER M1 ;
        RECT 15.328 10.296 15.36 12.804 ;
  LAYER M3 ;
        RECT 15.328 12.752 15.36 12.784 ;
  LAYER M1 ;
        RECT 15.392 10.296 15.424 12.804 ;
  LAYER M3 ;
        RECT 15.392 10.316 15.424 10.348 ;
  LAYER M1 ;
        RECT 15.456 10.296 15.488 12.804 ;
  LAYER M3 ;
        RECT 15.456 12.752 15.488 12.784 ;
  LAYER M1 ;
        RECT 15.52 10.296 15.552 12.804 ;
  LAYER M3 ;
        RECT 15.52 10.316 15.552 10.348 ;
  LAYER M1 ;
        RECT 15.584 10.296 15.616 12.804 ;
  LAYER M3 ;
        RECT 15.584 12.752 15.616 12.784 ;
  LAYER M1 ;
        RECT 15.648 10.296 15.68 12.804 ;
  LAYER M3 ;
        RECT 15.648 10.316 15.68 10.348 ;
  LAYER M1 ;
        RECT 15.712 10.296 15.744 12.804 ;
  LAYER M3 ;
        RECT 15.712 12.752 15.744 12.784 ;
  LAYER M1 ;
        RECT 15.776 10.296 15.808 12.804 ;
  LAYER M3 ;
        RECT 15.776 10.316 15.808 10.348 ;
  LAYER M1 ;
        RECT 15.84 10.296 15.872 12.804 ;
  LAYER M3 ;
        RECT 15.84 12.752 15.872 12.784 ;
  LAYER M1 ;
        RECT 15.904 10.296 15.936 12.804 ;
  LAYER M3 ;
        RECT 15.904 10.316 15.936 10.348 ;
  LAYER M1 ;
        RECT 15.968 10.296 16 12.804 ;
  LAYER M3 ;
        RECT 15.968 12.752 16 12.784 ;
  LAYER M1 ;
        RECT 16.032 10.296 16.064 12.804 ;
  LAYER M3 ;
        RECT 16.032 10.316 16.064 10.348 ;
  LAYER M1 ;
        RECT 16.096 10.296 16.128 12.804 ;
  LAYER M3 ;
        RECT 16.096 12.752 16.128 12.784 ;
  LAYER M1 ;
        RECT 16.16 10.296 16.192 12.804 ;
  LAYER M3 ;
        RECT 16.16 10.316 16.192 10.348 ;
  LAYER M1 ;
        RECT 16.224 10.296 16.256 12.804 ;
  LAYER M3 ;
        RECT 16.224 12.752 16.256 12.784 ;
  LAYER M1 ;
        RECT 16.288 10.296 16.32 12.804 ;
  LAYER M3 ;
        RECT 16.288 10.316 16.32 10.348 ;
  LAYER M1 ;
        RECT 16.352 10.296 16.384 12.804 ;
  LAYER M3 ;
        RECT 16.352 12.752 16.384 12.784 ;
  LAYER M1 ;
        RECT 16.416 10.296 16.448 12.804 ;
  LAYER M3 ;
        RECT 16.416 10.316 16.448 10.348 ;
  LAYER M1 ;
        RECT 16.48 10.296 16.512 12.804 ;
  LAYER M3 ;
        RECT 16.48 12.752 16.512 12.784 ;
  LAYER M1 ;
        RECT 16.544 10.296 16.576 12.804 ;
  LAYER M3 ;
        RECT 16.544 10.316 16.576 10.348 ;
  LAYER M1 ;
        RECT 16.608 10.296 16.64 12.804 ;
  LAYER M3 ;
        RECT 16.608 12.752 16.64 12.784 ;
  LAYER M1 ;
        RECT 16.672 10.296 16.704 12.804 ;
  LAYER M3 ;
        RECT 16.672 10.316 16.704 10.348 ;
  LAYER M1 ;
        RECT 16.736 10.296 16.768 12.804 ;
  LAYER M3 ;
        RECT 16.736 12.752 16.768 12.784 ;
  LAYER M1 ;
        RECT 16.8 10.296 16.832 12.804 ;
  LAYER M3 ;
        RECT 16.8 10.316 16.832 10.348 ;
  LAYER M1 ;
        RECT 16.864 10.296 16.896 12.804 ;
  LAYER M3 ;
        RECT 16.864 12.752 16.896 12.784 ;
  LAYER M1 ;
        RECT 16.928 10.296 16.96 12.804 ;
  LAYER M3 ;
        RECT 16.928 10.316 16.96 10.348 ;
  LAYER M1 ;
        RECT 16.992 10.296 17.024 12.804 ;
  LAYER M3 ;
        RECT 16.992 12.752 17.024 12.784 ;
  LAYER M1 ;
        RECT 17.056 10.296 17.088 12.804 ;
  LAYER M3 ;
        RECT 17.056 10.316 17.088 10.348 ;
  LAYER M1 ;
        RECT 17.12 10.296 17.152 12.804 ;
  LAYER M3 ;
        RECT 17.12 12.752 17.152 12.784 ;
  LAYER M1 ;
        RECT 17.184 10.296 17.216 12.804 ;
  LAYER M3 ;
        RECT 17.184 10.316 17.216 10.348 ;
  LAYER M1 ;
        RECT 17.248 10.296 17.28 12.804 ;
  LAYER M3 ;
        RECT 17.248 12.752 17.28 12.784 ;
  LAYER M1 ;
        RECT 17.312 10.296 17.344 12.804 ;
  LAYER M3 ;
        RECT 17.312 10.316 17.344 10.348 ;
  LAYER M1 ;
        RECT 17.376 10.296 17.408 12.804 ;
  LAYER M3 ;
        RECT 17.376 12.752 17.408 12.784 ;
  LAYER M1 ;
        RECT 17.44 10.296 17.472 12.804 ;
  LAYER M3 ;
        RECT 17.44 10.316 17.472 10.348 ;
  LAYER M1 ;
        RECT 17.504 10.296 17.536 12.804 ;
  LAYER M3 ;
        RECT 17.504 12.752 17.536 12.784 ;
  LAYER M1 ;
        RECT 17.568 10.296 17.6 12.804 ;
  LAYER M3 ;
        RECT 17.568 10.316 17.6 10.348 ;
  LAYER M1 ;
        RECT 17.632 10.296 17.664 12.804 ;
  LAYER M3 ;
        RECT 17.632 12.752 17.664 12.784 ;
  LAYER M1 ;
        RECT 17.696 10.296 17.728 12.804 ;
  LAYER M3 ;
        RECT 15.328 10.38 15.36 10.412 ;
  LAYER M2 ;
        RECT 17.696 10.444 17.728 10.476 ;
  LAYER M2 ;
        RECT 15.328 10.508 15.36 10.54 ;
  LAYER M2 ;
        RECT 17.696 10.572 17.728 10.604 ;
  LAYER M2 ;
        RECT 15.328 10.636 15.36 10.668 ;
  LAYER M2 ;
        RECT 17.696 10.7 17.728 10.732 ;
  LAYER M2 ;
        RECT 15.328 10.764 15.36 10.796 ;
  LAYER M2 ;
        RECT 17.696 10.828 17.728 10.86 ;
  LAYER M2 ;
        RECT 15.328 10.892 15.36 10.924 ;
  LAYER M2 ;
        RECT 17.696 10.956 17.728 10.988 ;
  LAYER M2 ;
        RECT 15.328 11.02 15.36 11.052 ;
  LAYER M2 ;
        RECT 17.696 11.084 17.728 11.116 ;
  LAYER M2 ;
        RECT 15.328 11.148 15.36 11.18 ;
  LAYER M2 ;
        RECT 17.696 11.212 17.728 11.244 ;
  LAYER M2 ;
        RECT 15.328 11.276 15.36 11.308 ;
  LAYER M2 ;
        RECT 17.696 11.34 17.728 11.372 ;
  LAYER M2 ;
        RECT 15.328 11.404 15.36 11.436 ;
  LAYER M2 ;
        RECT 17.696 11.468 17.728 11.5 ;
  LAYER M2 ;
        RECT 15.328 11.532 15.36 11.564 ;
  LAYER M2 ;
        RECT 17.696 11.596 17.728 11.628 ;
  LAYER M2 ;
        RECT 15.328 11.66 15.36 11.692 ;
  LAYER M2 ;
        RECT 17.696 11.724 17.728 11.756 ;
  LAYER M2 ;
        RECT 15.328 11.788 15.36 11.82 ;
  LAYER M2 ;
        RECT 17.696 11.852 17.728 11.884 ;
  LAYER M2 ;
        RECT 15.328 11.916 15.36 11.948 ;
  LAYER M2 ;
        RECT 17.696 11.98 17.728 12.012 ;
  LAYER M2 ;
        RECT 15.328 12.044 15.36 12.076 ;
  LAYER M2 ;
        RECT 17.696 12.108 17.728 12.14 ;
  LAYER M2 ;
        RECT 15.328 12.172 15.36 12.204 ;
  LAYER M2 ;
        RECT 17.696 12.236 17.728 12.268 ;
  LAYER M2 ;
        RECT 15.328 12.3 15.36 12.332 ;
  LAYER M2 ;
        RECT 17.696 12.364 17.728 12.396 ;
  LAYER M2 ;
        RECT 15.328 12.428 15.36 12.46 ;
  LAYER M2 ;
        RECT 17.696 12.492 17.728 12.524 ;
  LAYER M2 ;
        RECT 15.328 12.556 15.36 12.588 ;
  LAYER M2 ;
        RECT 17.696 12.62 17.728 12.652 ;
  LAYER M2 ;
        RECT 15.28 10.248 17.776 12.852 ;
  LAYER M1 ;
        RECT 15.328 13.404 15.36 15.912 ;
  LAYER M3 ;
        RECT 15.328 15.86 15.36 15.892 ;
  LAYER M1 ;
        RECT 15.392 13.404 15.424 15.912 ;
  LAYER M3 ;
        RECT 15.392 13.424 15.424 13.456 ;
  LAYER M1 ;
        RECT 15.456 13.404 15.488 15.912 ;
  LAYER M3 ;
        RECT 15.456 15.86 15.488 15.892 ;
  LAYER M1 ;
        RECT 15.52 13.404 15.552 15.912 ;
  LAYER M3 ;
        RECT 15.52 13.424 15.552 13.456 ;
  LAYER M1 ;
        RECT 15.584 13.404 15.616 15.912 ;
  LAYER M3 ;
        RECT 15.584 15.86 15.616 15.892 ;
  LAYER M1 ;
        RECT 15.648 13.404 15.68 15.912 ;
  LAYER M3 ;
        RECT 15.648 13.424 15.68 13.456 ;
  LAYER M1 ;
        RECT 15.712 13.404 15.744 15.912 ;
  LAYER M3 ;
        RECT 15.712 15.86 15.744 15.892 ;
  LAYER M1 ;
        RECT 15.776 13.404 15.808 15.912 ;
  LAYER M3 ;
        RECT 15.776 13.424 15.808 13.456 ;
  LAYER M1 ;
        RECT 15.84 13.404 15.872 15.912 ;
  LAYER M3 ;
        RECT 15.84 15.86 15.872 15.892 ;
  LAYER M1 ;
        RECT 15.904 13.404 15.936 15.912 ;
  LAYER M3 ;
        RECT 15.904 13.424 15.936 13.456 ;
  LAYER M1 ;
        RECT 15.968 13.404 16 15.912 ;
  LAYER M3 ;
        RECT 15.968 15.86 16 15.892 ;
  LAYER M1 ;
        RECT 16.032 13.404 16.064 15.912 ;
  LAYER M3 ;
        RECT 16.032 13.424 16.064 13.456 ;
  LAYER M1 ;
        RECT 16.096 13.404 16.128 15.912 ;
  LAYER M3 ;
        RECT 16.096 15.86 16.128 15.892 ;
  LAYER M1 ;
        RECT 16.16 13.404 16.192 15.912 ;
  LAYER M3 ;
        RECT 16.16 13.424 16.192 13.456 ;
  LAYER M1 ;
        RECT 16.224 13.404 16.256 15.912 ;
  LAYER M3 ;
        RECT 16.224 15.86 16.256 15.892 ;
  LAYER M1 ;
        RECT 16.288 13.404 16.32 15.912 ;
  LAYER M3 ;
        RECT 16.288 13.424 16.32 13.456 ;
  LAYER M1 ;
        RECT 16.352 13.404 16.384 15.912 ;
  LAYER M3 ;
        RECT 16.352 15.86 16.384 15.892 ;
  LAYER M1 ;
        RECT 16.416 13.404 16.448 15.912 ;
  LAYER M3 ;
        RECT 16.416 13.424 16.448 13.456 ;
  LAYER M1 ;
        RECT 16.48 13.404 16.512 15.912 ;
  LAYER M3 ;
        RECT 16.48 15.86 16.512 15.892 ;
  LAYER M1 ;
        RECT 16.544 13.404 16.576 15.912 ;
  LAYER M3 ;
        RECT 16.544 13.424 16.576 13.456 ;
  LAYER M1 ;
        RECT 16.608 13.404 16.64 15.912 ;
  LAYER M3 ;
        RECT 16.608 15.86 16.64 15.892 ;
  LAYER M1 ;
        RECT 16.672 13.404 16.704 15.912 ;
  LAYER M3 ;
        RECT 16.672 13.424 16.704 13.456 ;
  LAYER M1 ;
        RECT 16.736 13.404 16.768 15.912 ;
  LAYER M3 ;
        RECT 16.736 15.86 16.768 15.892 ;
  LAYER M1 ;
        RECT 16.8 13.404 16.832 15.912 ;
  LAYER M3 ;
        RECT 16.8 13.424 16.832 13.456 ;
  LAYER M1 ;
        RECT 16.864 13.404 16.896 15.912 ;
  LAYER M3 ;
        RECT 16.864 15.86 16.896 15.892 ;
  LAYER M1 ;
        RECT 16.928 13.404 16.96 15.912 ;
  LAYER M3 ;
        RECT 16.928 13.424 16.96 13.456 ;
  LAYER M1 ;
        RECT 16.992 13.404 17.024 15.912 ;
  LAYER M3 ;
        RECT 16.992 15.86 17.024 15.892 ;
  LAYER M1 ;
        RECT 17.056 13.404 17.088 15.912 ;
  LAYER M3 ;
        RECT 17.056 13.424 17.088 13.456 ;
  LAYER M1 ;
        RECT 17.12 13.404 17.152 15.912 ;
  LAYER M3 ;
        RECT 17.12 15.86 17.152 15.892 ;
  LAYER M1 ;
        RECT 17.184 13.404 17.216 15.912 ;
  LAYER M3 ;
        RECT 17.184 13.424 17.216 13.456 ;
  LAYER M1 ;
        RECT 17.248 13.404 17.28 15.912 ;
  LAYER M3 ;
        RECT 17.248 15.86 17.28 15.892 ;
  LAYER M1 ;
        RECT 17.312 13.404 17.344 15.912 ;
  LAYER M3 ;
        RECT 17.312 13.424 17.344 13.456 ;
  LAYER M1 ;
        RECT 17.376 13.404 17.408 15.912 ;
  LAYER M3 ;
        RECT 17.376 15.86 17.408 15.892 ;
  LAYER M1 ;
        RECT 17.44 13.404 17.472 15.912 ;
  LAYER M3 ;
        RECT 17.44 13.424 17.472 13.456 ;
  LAYER M1 ;
        RECT 17.504 13.404 17.536 15.912 ;
  LAYER M3 ;
        RECT 17.504 15.86 17.536 15.892 ;
  LAYER M1 ;
        RECT 17.568 13.404 17.6 15.912 ;
  LAYER M3 ;
        RECT 17.568 13.424 17.6 13.456 ;
  LAYER M1 ;
        RECT 17.632 13.404 17.664 15.912 ;
  LAYER M3 ;
        RECT 17.632 15.86 17.664 15.892 ;
  LAYER M1 ;
        RECT 17.696 13.404 17.728 15.912 ;
  LAYER M3 ;
        RECT 15.328 13.488 15.36 13.52 ;
  LAYER M2 ;
        RECT 17.696 13.552 17.728 13.584 ;
  LAYER M2 ;
        RECT 15.328 13.616 15.36 13.648 ;
  LAYER M2 ;
        RECT 17.696 13.68 17.728 13.712 ;
  LAYER M2 ;
        RECT 15.328 13.744 15.36 13.776 ;
  LAYER M2 ;
        RECT 17.696 13.808 17.728 13.84 ;
  LAYER M2 ;
        RECT 15.328 13.872 15.36 13.904 ;
  LAYER M2 ;
        RECT 17.696 13.936 17.728 13.968 ;
  LAYER M2 ;
        RECT 15.328 14 15.36 14.032 ;
  LAYER M2 ;
        RECT 17.696 14.064 17.728 14.096 ;
  LAYER M2 ;
        RECT 15.328 14.128 15.36 14.16 ;
  LAYER M2 ;
        RECT 17.696 14.192 17.728 14.224 ;
  LAYER M2 ;
        RECT 15.328 14.256 15.36 14.288 ;
  LAYER M2 ;
        RECT 17.696 14.32 17.728 14.352 ;
  LAYER M2 ;
        RECT 15.328 14.384 15.36 14.416 ;
  LAYER M2 ;
        RECT 17.696 14.448 17.728 14.48 ;
  LAYER M2 ;
        RECT 15.328 14.512 15.36 14.544 ;
  LAYER M2 ;
        RECT 17.696 14.576 17.728 14.608 ;
  LAYER M2 ;
        RECT 15.328 14.64 15.36 14.672 ;
  LAYER M2 ;
        RECT 17.696 14.704 17.728 14.736 ;
  LAYER M2 ;
        RECT 15.328 14.768 15.36 14.8 ;
  LAYER M2 ;
        RECT 17.696 14.832 17.728 14.864 ;
  LAYER M2 ;
        RECT 15.328 14.896 15.36 14.928 ;
  LAYER M2 ;
        RECT 17.696 14.96 17.728 14.992 ;
  LAYER M2 ;
        RECT 15.328 15.024 15.36 15.056 ;
  LAYER M2 ;
        RECT 17.696 15.088 17.728 15.12 ;
  LAYER M2 ;
        RECT 15.328 15.152 15.36 15.184 ;
  LAYER M2 ;
        RECT 17.696 15.216 17.728 15.248 ;
  LAYER M2 ;
        RECT 15.328 15.28 15.36 15.312 ;
  LAYER M2 ;
        RECT 17.696 15.344 17.728 15.376 ;
  LAYER M2 ;
        RECT 15.328 15.408 15.36 15.44 ;
  LAYER M2 ;
        RECT 17.696 15.472 17.728 15.504 ;
  LAYER M2 ;
        RECT 15.328 15.536 15.36 15.568 ;
  LAYER M2 ;
        RECT 17.696 15.6 17.728 15.632 ;
  LAYER M2 ;
        RECT 15.328 15.664 15.36 15.696 ;
  LAYER M2 ;
        RECT 17.696 15.728 17.728 15.76 ;
  LAYER M2 ;
        RECT 15.28 13.356 17.776 15.96 ;
  END 
END Cap_60fF_Cap_60fF
