MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 18 BY 16.884 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
      LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
      LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
      LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
      LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 8.864 0.384 8.896 0.456 ;
      LAYER M2 ;
        RECT 8.844 0.404 8.916 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
      LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
      LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
      LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
      LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
      LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
      LAYER M1 ;
        RECT 11.84 0.216 11.872 0.288 ;
      LAYER M2 ;
        RECT 11.82 0.236 11.892 0.268 ;
      LAYER M2 ;
        RECT 5.904 0.236 11.856 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.704 7.188 8.736 7.26 ;
  LAYER M2 ;
        RECT 8.684 7.208 8.756 7.24 ;
  LAYER M1 ;
        RECT 8.704 7.056 8.736 7.224 ;
  LAYER M1 ;
        RECT 8.704 7.02 8.736 7.092 ;
  LAYER M2 ;
        RECT 8.684 7.04 8.756 7.072 ;
  LAYER M2 ;
        RECT 8.72 7.04 8.88 7.072 ;
  LAYER M1 ;
        RECT 8.864 7.02 8.896 7.092 ;
  LAYER M2 ;
        RECT 8.844 7.04 8.916 7.072 ;
  LAYER M1 ;
        RECT 11.68 7.188 11.712 7.26 ;
  LAYER M2 ;
        RECT 11.66 7.208 11.732 7.24 ;
  LAYER M2 ;
        RECT 8.88 7.208 11.696 7.24 ;
  LAYER M1 ;
        RECT 8.864 7.188 8.896 7.26 ;
  LAYER M2 ;
        RECT 8.844 7.208 8.916 7.24 ;
  LAYER M1 ;
        RECT 8.704 10.296 8.736 10.368 ;
  LAYER M2 ;
        RECT 8.684 10.316 8.756 10.348 ;
  LAYER M1 ;
        RECT 8.704 10.164 8.736 10.332 ;
  LAYER M1 ;
        RECT 8.704 10.128 8.736 10.2 ;
  LAYER M2 ;
        RECT 8.684 10.148 8.756 10.18 ;
  LAYER M2 ;
        RECT 8.72 10.148 8.88 10.18 ;
  LAYER M1 ;
        RECT 8.864 10.128 8.896 10.2 ;
  LAYER M2 ;
        RECT 8.844 10.148 8.916 10.18 ;
  LAYER M1 ;
        RECT 11.68 4.08 11.712 4.152 ;
  LAYER M2 ;
        RECT 11.66 4.1 11.732 4.132 ;
  LAYER M2 ;
        RECT 8.88 4.1 11.696 4.132 ;
  LAYER M1 ;
        RECT 8.864 4.08 8.896 4.152 ;
  LAYER M2 ;
        RECT 8.844 4.1 8.916 4.132 ;
  LAYER M1 ;
        RECT 8.704 4.08 8.736 4.152 ;
  LAYER M2 ;
        RECT 8.684 4.1 8.756 4.132 ;
  LAYER M1 ;
        RECT 8.704 3.948 8.736 4.116 ;
  LAYER M1 ;
        RECT 8.704 3.912 8.736 3.984 ;
  LAYER M2 ;
        RECT 8.684 3.932 8.756 3.964 ;
  LAYER M2 ;
        RECT 8.72 3.932 8.88 3.964 ;
  LAYER M1 ;
        RECT 8.864 3.912 8.896 3.984 ;
  LAYER M2 ;
        RECT 8.844 3.932 8.916 3.964 ;
  LAYER M1 ;
        RECT 11.68 10.296 11.712 10.368 ;
  LAYER M2 ;
        RECT 11.66 10.316 11.732 10.348 ;
  LAYER M2 ;
        RECT 8.88 10.316 11.696 10.348 ;
  LAYER M1 ;
        RECT 8.864 10.296 8.896 10.368 ;
  LAYER M2 ;
        RECT 8.844 10.316 8.916 10.348 ;
  LAYER M1 ;
        RECT 8.864 0.384 8.896 0.456 ;
  LAYER M2 ;
        RECT 8.844 0.404 8.916 0.436 ;
  LAYER M1 ;
        RECT 8.864 0.42 8.896 0.672 ;
  LAYER M1 ;
        RECT 8.864 0.672 8.896 10.332 ;
  LAYER M1 ;
        RECT 5.728 7.188 5.76 7.26 ;
  LAYER M2 ;
        RECT 5.708 7.208 5.78 7.24 ;
  LAYER M1 ;
        RECT 5.728 7.056 5.76 7.224 ;
  LAYER M1 ;
        RECT 5.728 7.02 5.76 7.092 ;
  LAYER M2 ;
        RECT 5.708 7.04 5.78 7.072 ;
  LAYER M2 ;
        RECT 5.744 7.04 5.904 7.072 ;
  LAYER M1 ;
        RECT 5.888 7.02 5.92 7.092 ;
  LAYER M2 ;
        RECT 5.868 7.04 5.94 7.072 ;
  LAYER M1 ;
        RECT 5.728 10.296 5.76 10.368 ;
  LAYER M2 ;
        RECT 5.708 10.316 5.78 10.348 ;
  LAYER M1 ;
        RECT 5.728 10.164 5.76 10.332 ;
  LAYER M1 ;
        RECT 5.728 10.128 5.76 10.2 ;
  LAYER M2 ;
        RECT 5.708 10.148 5.78 10.18 ;
  LAYER M2 ;
        RECT 5.744 10.148 5.904 10.18 ;
  LAYER M1 ;
        RECT 5.888 10.128 5.92 10.2 ;
  LAYER M2 ;
        RECT 5.868 10.148 5.94 10.18 ;
  LAYER M1 ;
        RECT 5.728 4.08 5.76 4.152 ;
  LAYER M2 ;
        RECT 5.708 4.1 5.78 4.132 ;
  LAYER M1 ;
        RECT 5.728 3.948 5.76 4.116 ;
  LAYER M1 ;
        RECT 5.728 3.912 5.76 3.984 ;
  LAYER M2 ;
        RECT 5.708 3.932 5.78 3.964 ;
  LAYER M2 ;
        RECT 5.744 3.932 5.904 3.964 ;
  LAYER M1 ;
        RECT 5.888 3.912 5.92 3.984 ;
  LAYER M2 ;
        RECT 5.868 3.932 5.94 3.964 ;
  LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
  LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
  LAYER M1 ;
        RECT 5.888 0.252 5.92 0.672 ;
  LAYER M1 ;
        RECT 5.888 0.672 5.92 10.164 ;
  LAYER M1 ;
        RECT 14.656 7.188 14.688 7.26 ;
  LAYER M2 ;
        RECT 14.636 7.208 14.708 7.24 ;
  LAYER M2 ;
        RECT 11.856 7.208 14.672 7.24 ;
  LAYER M1 ;
        RECT 11.84 7.188 11.872 7.26 ;
  LAYER M2 ;
        RECT 11.82 7.208 11.892 7.24 ;
  LAYER M1 ;
        RECT 14.656 4.08 14.688 4.152 ;
  LAYER M2 ;
        RECT 14.636 4.1 14.708 4.132 ;
  LAYER M2 ;
        RECT 11.856 4.1 14.672 4.132 ;
  LAYER M1 ;
        RECT 11.84 4.08 11.872 4.152 ;
  LAYER M2 ;
        RECT 11.82 4.1 11.892 4.132 ;
  LAYER M1 ;
        RECT 14.656 10.296 14.688 10.368 ;
  LAYER M2 ;
        RECT 14.636 10.316 14.708 10.348 ;
  LAYER M2 ;
        RECT 11.856 10.316 14.672 10.348 ;
  LAYER M1 ;
        RECT 11.84 10.296 11.872 10.368 ;
  LAYER M2 ;
        RECT 11.82 10.316 11.892 10.348 ;
  LAYER M1 ;
        RECT 11.84 0.216 11.872 0.288 ;
  LAYER M2 ;
        RECT 11.82 0.236 11.892 0.268 ;
  LAYER M1 ;
        RECT 11.84 0.252 11.872 0.672 ;
  LAYER M1 ;
        RECT 11.84 0.672 11.872 10.332 ;
  LAYER M2 ;
        RECT 5.904 0.236 11.856 0.268 ;
  LAYER M1 ;
        RECT 2.752 0.972 2.784 1.044 ;
  LAYER M2 ;
        RECT 2.732 0.992 2.804 1.024 ;
  LAYER M1 ;
        RECT 2.752 0.84 2.784 1.008 ;
  LAYER M1 ;
        RECT 2.752 0.804 2.784 0.876 ;
  LAYER M2 ;
        RECT 2.732 0.824 2.804 0.856 ;
  LAYER M2 ;
        RECT 2.768 0.824 2.928 0.856 ;
  LAYER M1 ;
        RECT 2.912 0.804 2.944 0.876 ;
  LAYER M2 ;
        RECT 2.892 0.824 2.964 0.856 ;
  LAYER M1 ;
        RECT 2.752 4.08 2.784 4.152 ;
  LAYER M2 ;
        RECT 2.732 4.1 2.804 4.132 ;
  LAYER M1 ;
        RECT 2.752 3.948 2.784 4.116 ;
  LAYER M1 ;
        RECT 2.752 3.912 2.784 3.984 ;
  LAYER M2 ;
        RECT 2.732 3.932 2.804 3.964 ;
  LAYER M2 ;
        RECT 2.768 3.932 2.928 3.964 ;
  LAYER M1 ;
        RECT 2.912 3.912 2.944 3.984 ;
  LAYER M2 ;
        RECT 2.892 3.932 2.964 3.964 ;
  LAYER M1 ;
        RECT 2.752 7.188 2.784 7.26 ;
  LAYER M2 ;
        RECT 2.732 7.208 2.804 7.24 ;
  LAYER M1 ;
        RECT 2.752 7.056 2.784 7.224 ;
  LAYER M1 ;
        RECT 2.752 7.02 2.784 7.092 ;
  LAYER M2 ;
        RECT 2.732 7.04 2.804 7.072 ;
  LAYER M2 ;
        RECT 2.768 7.04 2.928 7.072 ;
  LAYER M1 ;
        RECT 2.912 7.02 2.944 7.092 ;
  LAYER M2 ;
        RECT 2.892 7.04 2.964 7.072 ;
  LAYER M1 ;
        RECT 2.752 10.296 2.784 10.368 ;
  LAYER M2 ;
        RECT 2.732 10.316 2.804 10.348 ;
  LAYER M1 ;
        RECT 2.752 10.164 2.784 10.332 ;
  LAYER M1 ;
        RECT 2.752 10.128 2.784 10.2 ;
  LAYER M2 ;
        RECT 2.732 10.148 2.804 10.18 ;
  LAYER M2 ;
        RECT 2.768 10.148 2.928 10.18 ;
  LAYER M1 ;
        RECT 2.912 10.128 2.944 10.2 ;
  LAYER M2 ;
        RECT 2.892 10.148 2.964 10.18 ;
  LAYER M1 ;
        RECT 2.752 13.404 2.784 13.476 ;
  LAYER M2 ;
        RECT 2.732 13.424 2.804 13.456 ;
  LAYER M1 ;
        RECT 2.752 13.272 2.784 13.44 ;
  LAYER M1 ;
        RECT 2.752 13.236 2.784 13.308 ;
  LAYER M2 ;
        RECT 2.732 13.256 2.804 13.288 ;
  LAYER M2 ;
        RECT 2.768 13.256 2.928 13.288 ;
  LAYER M1 ;
        RECT 2.912 13.236 2.944 13.308 ;
  LAYER M2 ;
        RECT 2.892 13.256 2.964 13.288 ;
  LAYER M1 ;
        RECT 5.728 0.972 5.76 1.044 ;
  LAYER M2 ;
        RECT 5.708 0.992 5.78 1.024 ;
  LAYER M2 ;
        RECT 2.928 0.992 5.744 1.024 ;
  LAYER M1 ;
        RECT 2.912 0.972 2.944 1.044 ;
  LAYER M2 ;
        RECT 2.892 0.992 2.964 1.024 ;
  LAYER M1 ;
        RECT 5.728 13.404 5.76 13.476 ;
  LAYER M2 ;
        RECT 5.708 13.424 5.78 13.456 ;
  LAYER M2 ;
        RECT 2.928 13.424 5.744 13.456 ;
  LAYER M1 ;
        RECT 2.912 13.404 2.944 13.476 ;
  LAYER M2 ;
        RECT 2.892 13.424 2.964 13.456 ;
  LAYER M1 ;
        RECT 2.912 0.048 2.944 0.12 ;
  LAYER M2 ;
        RECT 2.892 0.068 2.964 0.1 ;
  LAYER M1 ;
        RECT 2.912 0.084 2.944 0.672 ;
  LAYER M1 ;
        RECT 2.912 0.672 2.944 13.44 ;
  LAYER M1 ;
        RECT 14.656 0.972 14.688 1.044 ;
  LAYER M2 ;
        RECT 14.636 0.992 14.708 1.024 ;
  LAYER M1 ;
        RECT 14.656 0.84 14.688 1.008 ;
  LAYER M1 ;
        RECT 14.656 0.804 14.688 0.876 ;
  LAYER M2 ;
        RECT 14.636 0.824 14.708 0.856 ;
  LAYER M2 ;
        RECT 14.672 0.824 14.832 0.856 ;
  LAYER M1 ;
        RECT 14.816 0.804 14.848 0.876 ;
  LAYER M2 ;
        RECT 14.796 0.824 14.868 0.856 ;
  LAYER M1 ;
        RECT 14.656 13.404 14.688 13.476 ;
  LAYER M2 ;
        RECT 14.636 13.424 14.708 13.456 ;
  LAYER M1 ;
        RECT 14.656 13.272 14.688 13.44 ;
  LAYER M1 ;
        RECT 14.656 13.236 14.688 13.308 ;
  LAYER M2 ;
        RECT 14.636 13.256 14.708 13.288 ;
  LAYER M2 ;
        RECT 14.672 13.256 14.832 13.288 ;
  LAYER M1 ;
        RECT 14.816 13.236 14.848 13.308 ;
  LAYER M2 ;
        RECT 14.796 13.256 14.868 13.288 ;
  LAYER M1 ;
        RECT 17.632 0.972 17.664 1.044 ;
  LAYER M2 ;
        RECT 17.612 0.992 17.684 1.024 ;
  LAYER M2 ;
        RECT 14.832 0.992 17.648 1.024 ;
  LAYER M1 ;
        RECT 14.816 0.972 14.848 1.044 ;
  LAYER M2 ;
        RECT 14.796 0.992 14.868 1.024 ;
  LAYER M1 ;
        RECT 17.632 4.08 17.664 4.152 ;
  LAYER M2 ;
        RECT 17.612 4.1 17.684 4.132 ;
  LAYER M2 ;
        RECT 14.832 4.1 17.648 4.132 ;
  LAYER M1 ;
        RECT 14.816 4.08 14.848 4.152 ;
  LAYER M2 ;
        RECT 14.796 4.1 14.868 4.132 ;
  LAYER M1 ;
        RECT 17.632 7.188 17.664 7.26 ;
  LAYER M2 ;
        RECT 17.612 7.208 17.684 7.24 ;
  LAYER M2 ;
        RECT 14.832 7.208 17.648 7.24 ;
  LAYER M1 ;
        RECT 14.816 7.188 14.848 7.26 ;
  LAYER M2 ;
        RECT 14.796 7.208 14.868 7.24 ;
  LAYER M1 ;
        RECT 17.632 10.296 17.664 10.368 ;
  LAYER M2 ;
        RECT 17.612 10.316 17.684 10.348 ;
  LAYER M2 ;
        RECT 14.832 10.316 17.648 10.348 ;
  LAYER M1 ;
        RECT 14.816 10.296 14.848 10.368 ;
  LAYER M2 ;
        RECT 14.796 10.316 14.868 10.348 ;
  LAYER M1 ;
        RECT 17.632 13.404 17.664 13.476 ;
  LAYER M2 ;
        RECT 17.612 13.424 17.684 13.456 ;
  LAYER M2 ;
        RECT 14.832 13.424 17.648 13.456 ;
  LAYER M1 ;
        RECT 14.816 13.404 14.848 13.476 ;
  LAYER M2 ;
        RECT 14.796 13.424 14.868 13.456 ;
  LAYER M1 ;
        RECT 14.816 0.048 14.848 0.12 ;
  LAYER M2 ;
        RECT 14.796 0.068 14.868 0.1 ;
  LAYER M1 ;
        RECT 14.816 0.084 14.848 0.672 ;
  LAYER M1 ;
        RECT 14.816 0.672 14.848 13.44 ;
  LAYER M2 ;
        RECT 2.928 0.068 14.832 0.1 ;
  LAYER M1 ;
        RECT 8.704 13.404 8.736 13.476 ;
  LAYER M2 ;
        RECT 8.684 13.424 8.756 13.456 ;
  LAYER M2 ;
        RECT 5.744 13.424 8.72 13.456 ;
  LAYER M1 ;
        RECT 5.728 13.404 5.76 13.476 ;
  LAYER M2 ;
        RECT 5.708 13.424 5.78 13.456 ;
  LAYER M1 ;
        RECT 11.68 13.404 11.712 13.476 ;
  LAYER M2 ;
        RECT 11.66 13.424 11.732 13.456 ;
  LAYER M2 ;
        RECT 8.72 13.424 11.696 13.456 ;
  LAYER M1 ;
        RECT 8.704 13.404 8.736 13.476 ;
  LAYER M2 ;
        RECT 8.684 13.424 8.756 13.456 ;
  LAYER M1 ;
        RECT 11.68 0.972 11.712 1.044 ;
  LAYER M2 ;
        RECT 11.66 0.992 11.732 1.024 ;
  LAYER M2 ;
        RECT 11.696 0.992 14.672 1.024 ;
  LAYER M1 ;
        RECT 14.656 0.972 14.688 1.044 ;
  LAYER M2 ;
        RECT 14.636 0.992 14.708 1.024 ;
  LAYER M1 ;
        RECT 8.704 0.972 8.736 1.044 ;
  LAYER M2 ;
        RECT 8.684 0.992 8.756 1.024 ;
  LAYER M2 ;
        RECT 8.72 0.992 11.696 1.024 ;
  LAYER M1 ;
        RECT 11.68 0.972 11.712 1.044 ;
  LAYER M2 ;
        RECT 11.66 0.992 11.732 1.024 ;
  LAYER M1 ;
        RECT 6.336 9.624 6.368 9.696 ;
  LAYER M2 ;
        RECT 6.316 9.644 6.388 9.676 ;
  LAYER M2 ;
        RECT 6.192 9.644 6.352 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 6.336 12.732 6.368 12.804 ;
  LAYER M2 ;
        RECT 6.316 12.752 6.388 12.784 ;
  LAYER M2 ;
        RECT 6.192 12.752 6.352 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 6.336 6.516 6.368 6.588 ;
  LAYER M2 ;
        RECT 6.316 6.536 6.388 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.352 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
  LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
  LAYER M1 ;
        RECT 6.176 16.212 6.208 16.464 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 16.212 ;
  LAYER M1 ;
        RECT 9.312 9.624 9.344 9.696 ;
  LAYER M2 ;
        RECT 9.292 9.644 9.364 9.676 ;
  LAYER M1 ;
        RECT 9.312 9.66 9.344 9.828 ;
  LAYER M1 ;
        RECT 9.312 9.792 9.344 9.864 ;
  LAYER M2 ;
        RECT 9.292 9.812 9.364 9.844 ;
  LAYER M2 ;
        RECT 9.328 9.812 12.144 9.844 ;
  LAYER M1 ;
        RECT 12.128 9.792 12.16 9.864 ;
  LAYER M2 ;
        RECT 12.108 9.812 12.18 9.844 ;
  LAYER M1 ;
        RECT 9.312 6.516 9.344 6.588 ;
  LAYER M2 ;
        RECT 9.292 6.536 9.364 6.568 ;
  LAYER M1 ;
        RECT 9.312 6.552 9.344 6.72 ;
  LAYER M1 ;
        RECT 9.312 6.684 9.344 6.756 ;
  LAYER M2 ;
        RECT 9.292 6.704 9.364 6.736 ;
  LAYER M2 ;
        RECT 9.328 6.704 12.144 6.736 ;
  LAYER M1 ;
        RECT 12.128 6.684 12.16 6.756 ;
  LAYER M2 ;
        RECT 12.108 6.704 12.18 6.736 ;
  LAYER M1 ;
        RECT 9.312 12.732 9.344 12.804 ;
  LAYER M2 ;
        RECT 9.292 12.752 9.364 12.784 ;
  LAYER M1 ;
        RECT 9.312 12.768 9.344 12.936 ;
  LAYER M1 ;
        RECT 9.312 12.9 9.344 12.972 ;
  LAYER M2 ;
        RECT 9.292 12.92 9.364 12.952 ;
  LAYER M2 ;
        RECT 9.328 12.92 12.144 12.952 ;
  LAYER M1 ;
        RECT 12.128 12.9 12.16 12.972 ;
  LAYER M2 ;
        RECT 12.108 12.92 12.18 12.952 ;
  LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
  LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
  LAYER M1 ;
        RECT 12.128 16.212 12.16 16.464 ;
  LAYER M1 ;
        RECT 12.128 6.72 12.16 16.212 ;
  LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
  LAYER M1 ;
        RECT 3.36 9.624 3.392 9.696 ;
  LAYER M2 ;
        RECT 3.34 9.644 3.412 9.676 ;
  LAYER M2 ;
        RECT 3.216 9.644 3.376 9.676 ;
  LAYER M1 ;
        RECT 3.2 9.624 3.232 9.696 ;
  LAYER M2 ;
        RECT 3.18 9.644 3.252 9.676 ;
  LAYER M1 ;
        RECT 3.36 12.732 3.392 12.804 ;
  LAYER M2 ;
        RECT 3.34 12.752 3.412 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.376 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.36 6.516 3.392 6.588 ;
  LAYER M2 ;
        RECT 3.34 6.536 3.412 6.568 ;
  LAYER M2 ;
        RECT 3.216 6.536 3.376 6.568 ;
  LAYER M1 ;
        RECT 3.2 6.516 3.232 6.588 ;
  LAYER M2 ;
        RECT 3.18 6.536 3.252 6.568 ;
  LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
  LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
  LAYER M1 ;
        RECT 3.2 16.212 3.232 16.632 ;
  LAYER M1 ;
        RECT 3.2 6.552 3.232 16.212 ;
  LAYER M1 ;
        RECT 12.288 9.624 12.32 9.696 ;
  LAYER M2 ;
        RECT 12.268 9.644 12.34 9.676 ;
  LAYER M1 ;
        RECT 12.288 9.66 12.32 9.828 ;
  LAYER M1 ;
        RECT 12.288 9.792 12.32 9.864 ;
  LAYER M2 ;
        RECT 12.268 9.812 12.34 9.844 ;
  LAYER M2 ;
        RECT 12.304 9.812 15.12 9.844 ;
  LAYER M1 ;
        RECT 15.104 9.792 15.136 9.864 ;
  LAYER M2 ;
        RECT 15.084 9.812 15.156 9.844 ;
  LAYER M1 ;
        RECT 12.288 6.516 12.32 6.588 ;
  LAYER M2 ;
        RECT 12.268 6.536 12.34 6.568 ;
  LAYER M1 ;
        RECT 12.288 6.552 12.32 6.72 ;
  LAYER M1 ;
        RECT 12.288 6.684 12.32 6.756 ;
  LAYER M2 ;
        RECT 12.268 6.704 12.34 6.736 ;
  LAYER M2 ;
        RECT 12.304 6.704 15.12 6.736 ;
  LAYER M1 ;
        RECT 15.104 6.684 15.136 6.756 ;
  LAYER M2 ;
        RECT 15.084 6.704 15.156 6.736 ;
  LAYER M1 ;
        RECT 12.288 12.732 12.32 12.804 ;
  LAYER M2 ;
        RECT 12.268 12.752 12.34 12.784 ;
  LAYER M1 ;
        RECT 12.288 12.768 12.32 12.936 ;
  LAYER M1 ;
        RECT 12.288 12.9 12.32 12.972 ;
  LAYER M2 ;
        RECT 12.268 12.92 12.34 12.952 ;
  LAYER M2 ;
        RECT 12.304 12.92 15.12 12.952 ;
  LAYER M1 ;
        RECT 15.104 12.9 15.136 12.972 ;
  LAYER M2 ;
        RECT 15.084 12.92 15.156 12.952 ;
  LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
  LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
  LAYER M1 ;
        RECT 15.104 16.212 15.136 16.632 ;
  LAYER M1 ;
        RECT 15.104 6.72 15.136 16.212 ;
  LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
  LAYER M1 ;
        RECT 0.384 3.408 0.416 3.48 ;
  LAYER M2 ;
        RECT 0.364 3.428 0.436 3.46 ;
  LAYER M2 ;
        RECT 0.08 3.428 0.4 3.46 ;
  LAYER M1 ;
        RECT 0.064 3.408 0.096 3.48 ;
  LAYER M2 ;
        RECT 0.044 3.428 0.116 3.46 ;
  LAYER M1 ;
        RECT 0.384 6.516 0.416 6.588 ;
  LAYER M2 ;
        RECT 0.364 6.536 0.436 6.568 ;
  LAYER M2 ;
        RECT 0.08 6.536 0.4 6.568 ;
  LAYER M1 ;
        RECT 0.064 6.516 0.096 6.588 ;
  LAYER M2 ;
        RECT 0.044 6.536 0.116 6.568 ;
  LAYER M1 ;
        RECT 0.384 9.624 0.416 9.696 ;
  LAYER M2 ;
        RECT 0.364 9.644 0.436 9.676 ;
  LAYER M2 ;
        RECT 0.08 9.644 0.4 9.676 ;
  LAYER M1 ;
        RECT 0.064 9.624 0.096 9.696 ;
  LAYER M2 ;
        RECT 0.044 9.644 0.116 9.676 ;
  LAYER M1 ;
        RECT 0.384 12.732 0.416 12.804 ;
  LAYER M2 ;
        RECT 0.364 12.752 0.436 12.784 ;
  LAYER M2 ;
        RECT 0.08 12.752 0.4 12.784 ;
  LAYER M1 ;
        RECT 0.064 12.732 0.096 12.804 ;
  LAYER M2 ;
        RECT 0.044 12.752 0.116 12.784 ;
  LAYER M1 ;
        RECT 0.384 15.84 0.416 15.912 ;
  LAYER M2 ;
        RECT 0.364 15.86 0.436 15.892 ;
  LAYER M2 ;
        RECT 0.08 15.86 0.4 15.892 ;
  LAYER M1 ;
        RECT 0.064 15.84 0.096 15.912 ;
  LAYER M2 ;
        RECT 0.044 15.86 0.116 15.892 ;
  LAYER M1 ;
        RECT 0.064 16.764 0.096 16.836 ;
  LAYER M2 ;
        RECT 0.044 16.784 0.116 16.816 ;
  LAYER M1 ;
        RECT 0.064 16.212 0.096 16.8 ;
  LAYER M1 ;
        RECT 0.064 3.444 0.096 16.212 ;
  LAYER M1 ;
        RECT 15.264 3.408 15.296 3.48 ;
  LAYER M2 ;
        RECT 15.244 3.428 15.316 3.46 ;
  LAYER M1 ;
        RECT 15.264 3.444 15.296 3.612 ;
  LAYER M1 ;
        RECT 15.264 3.576 15.296 3.648 ;
  LAYER M2 ;
        RECT 15.244 3.596 15.316 3.628 ;
  LAYER M2 ;
        RECT 15.28 3.596 17.936 3.628 ;
  LAYER M1 ;
        RECT 17.92 3.576 17.952 3.648 ;
  LAYER M2 ;
        RECT 17.9 3.596 17.972 3.628 ;
  LAYER M1 ;
        RECT 15.264 6.516 15.296 6.588 ;
  LAYER M2 ;
        RECT 15.244 6.536 15.316 6.568 ;
  LAYER M1 ;
        RECT 15.264 6.552 15.296 6.72 ;
  LAYER M1 ;
        RECT 15.264 6.684 15.296 6.756 ;
  LAYER M2 ;
        RECT 15.244 6.704 15.316 6.736 ;
  LAYER M2 ;
        RECT 15.28 6.704 17.936 6.736 ;
  LAYER M1 ;
        RECT 17.92 6.684 17.952 6.756 ;
  LAYER M2 ;
        RECT 17.9 6.704 17.972 6.736 ;
  LAYER M1 ;
        RECT 15.264 9.624 15.296 9.696 ;
  LAYER M2 ;
        RECT 15.244 9.644 15.316 9.676 ;
  LAYER M1 ;
        RECT 15.264 9.66 15.296 9.828 ;
  LAYER M1 ;
        RECT 15.264 9.792 15.296 9.864 ;
  LAYER M2 ;
        RECT 15.244 9.812 15.316 9.844 ;
  LAYER M2 ;
        RECT 15.28 9.812 17.936 9.844 ;
  LAYER M1 ;
        RECT 17.92 9.792 17.952 9.864 ;
  LAYER M2 ;
        RECT 17.9 9.812 17.972 9.844 ;
  LAYER M1 ;
        RECT 15.264 12.732 15.296 12.804 ;
  LAYER M2 ;
        RECT 15.244 12.752 15.316 12.784 ;
  LAYER M1 ;
        RECT 15.264 12.768 15.296 12.936 ;
  LAYER M1 ;
        RECT 15.264 12.9 15.296 12.972 ;
  LAYER M2 ;
        RECT 15.244 12.92 15.316 12.952 ;
  LAYER M2 ;
        RECT 15.28 12.92 17.936 12.952 ;
  LAYER M1 ;
        RECT 17.92 12.9 17.952 12.972 ;
  LAYER M2 ;
        RECT 17.9 12.92 17.972 12.952 ;
  LAYER M1 ;
        RECT 15.264 15.84 15.296 15.912 ;
  LAYER M2 ;
        RECT 15.244 15.86 15.316 15.892 ;
  LAYER M1 ;
        RECT 15.264 15.876 15.296 16.044 ;
  LAYER M1 ;
        RECT 15.264 16.008 15.296 16.08 ;
  LAYER M2 ;
        RECT 15.244 16.028 15.316 16.06 ;
  LAYER M2 ;
        RECT 15.28 16.028 17.936 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.008 17.952 16.08 ;
  LAYER M2 ;
        RECT 17.9 16.028 17.972 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.764 17.952 16.836 ;
  LAYER M2 ;
        RECT 17.9 16.784 17.972 16.816 ;
  LAYER M1 ;
        RECT 17.92 16.212 17.952 16.8 ;
  LAYER M1 ;
        RECT 17.92 3.612 17.952 16.212 ;
  LAYER M2 ;
        RECT 0.08 16.784 17.936 16.816 ;
  LAYER M1 ;
        RECT 3.36 3.408 3.392 3.48 ;
  LAYER M2 ;
        RECT 3.34 3.428 3.412 3.46 ;
  LAYER M2 ;
        RECT 0.4 3.428 3.376 3.46 ;
  LAYER M1 ;
        RECT 0.384 3.408 0.416 3.48 ;
  LAYER M2 ;
        RECT 0.364 3.428 0.436 3.46 ;
  LAYER M1 ;
        RECT 3.36 15.84 3.392 15.912 ;
  LAYER M2 ;
        RECT 3.34 15.86 3.412 15.892 ;
  LAYER M2 ;
        RECT 0.4 15.86 3.376 15.892 ;
  LAYER M1 ;
        RECT 0.384 15.84 0.416 15.912 ;
  LAYER M2 ;
        RECT 0.364 15.86 0.436 15.892 ;
  LAYER M1 ;
        RECT 6.336 15.84 6.368 15.912 ;
  LAYER M2 ;
        RECT 6.316 15.86 6.388 15.892 ;
  LAYER M2 ;
        RECT 3.376 15.86 6.352 15.892 ;
  LAYER M1 ;
        RECT 3.36 15.84 3.392 15.912 ;
  LAYER M2 ;
        RECT 3.34 15.86 3.412 15.892 ;
  LAYER M1 ;
        RECT 9.312 15.84 9.344 15.912 ;
  LAYER M2 ;
        RECT 9.292 15.86 9.364 15.892 ;
  LAYER M2 ;
        RECT 6.352 15.86 9.328 15.892 ;
  LAYER M1 ;
        RECT 6.336 15.84 6.368 15.912 ;
  LAYER M2 ;
        RECT 6.316 15.86 6.388 15.892 ;
  LAYER M1 ;
        RECT 12.288 15.84 12.32 15.912 ;
  LAYER M2 ;
        RECT 12.268 15.86 12.34 15.892 ;
  LAYER M2 ;
        RECT 9.328 15.86 12.304 15.892 ;
  LAYER M1 ;
        RECT 9.312 15.84 9.344 15.912 ;
  LAYER M2 ;
        RECT 9.292 15.86 9.364 15.892 ;
  LAYER M1 ;
        RECT 12.288 3.408 12.32 3.48 ;
  LAYER M2 ;
        RECT 12.268 3.428 12.34 3.46 ;
  LAYER M2 ;
        RECT 12.304 3.428 15.28 3.46 ;
  LAYER M1 ;
        RECT 15.264 3.408 15.296 3.48 ;
  LAYER M2 ;
        RECT 15.244 3.428 15.316 3.46 ;
  LAYER M1 ;
        RECT 9.312 3.408 9.344 3.48 ;
  LAYER M2 ;
        RECT 9.292 3.428 9.364 3.46 ;
  LAYER M2 ;
        RECT 9.328 3.428 12.304 3.46 ;
  LAYER M1 ;
        RECT 12.288 3.408 12.32 3.48 ;
  LAYER M2 ;
        RECT 12.268 3.428 12.34 3.46 ;
  LAYER M1 ;
        RECT 6.336 3.408 6.368 3.48 ;
  LAYER M2 ;
        RECT 6.316 3.428 6.388 3.46 ;
  LAYER M2 ;
        RECT 6.352 3.428 9.328 3.46 ;
  LAYER M1 ;
        RECT 9.312 3.408 9.344 3.48 ;
  LAYER M2 ;
        RECT 9.292 3.428 9.364 3.46 ;
  LAYER M1 ;
        RECT 0.336 0.924 2.832 3.528 ;
  LAYER M3 ;
        RECT 0.336 0.924 2.832 3.528 ;
  LAYER M2 ;
        RECT 0.336 0.924 2.832 3.528 ;
  LAYER M1 ;
        RECT 0.336 4.032 2.832 6.636 ;
  LAYER M3 ;
        RECT 0.336 4.032 2.832 6.636 ;
  LAYER M2 ;
        RECT 0.336 4.032 2.832 6.636 ;
  LAYER M1 ;
        RECT 0.336 7.14 2.832 9.744 ;
  LAYER M3 ;
        RECT 0.336 7.14 2.832 9.744 ;
  LAYER M2 ;
        RECT 0.336 7.14 2.832 9.744 ;
  LAYER M1 ;
        RECT 0.336 10.248 2.832 12.852 ;
  LAYER M3 ;
        RECT 0.336 10.248 2.832 12.852 ;
  LAYER M2 ;
        RECT 0.336 10.248 2.832 12.852 ;
  LAYER M1 ;
        RECT 0.336 13.356 2.832 15.96 ;
  LAYER M3 ;
        RECT 0.336 13.356 2.832 15.96 ;
  LAYER M2 ;
        RECT 0.336 13.356 2.832 15.96 ;
  LAYER M1 ;
        RECT 3.312 0.924 5.808 3.528 ;
  LAYER M3 ;
        RECT 3.312 0.924 5.808 3.528 ;
  LAYER M2 ;
        RECT 3.312 0.924 5.808 3.528 ;
  LAYER M1 ;
        RECT 3.312 4.032 5.808 6.636 ;
  LAYER M3 ;
        RECT 3.312 4.032 5.808 6.636 ;
  LAYER M2 ;
        RECT 3.312 4.032 5.808 6.636 ;
  LAYER M1 ;
        RECT 3.312 7.14 5.808 9.744 ;
  LAYER M3 ;
        RECT 3.312 7.14 5.808 9.744 ;
  LAYER M2 ;
        RECT 3.312 7.14 5.808 9.744 ;
  LAYER M1 ;
        RECT 3.312 10.248 5.808 12.852 ;
  LAYER M3 ;
        RECT 3.312 10.248 5.808 12.852 ;
  LAYER M2 ;
        RECT 3.312 10.248 5.808 12.852 ;
  LAYER M1 ;
        RECT 3.312 13.356 5.808 15.96 ;
  LAYER M3 ;
        RECT 3.312 13.356 5.808 15.96 ;
  LAYER M2 ;
        RECT 3.312 13.356 5.808 15.96 ;
  LAYER M1 ;
        RECT 6.288 0.924 8.784 3.528 ;
  LAYER M3 ;
        RECT 6.288 0.924 8.784 3.528 ;
  LAYER M2 ;
        RECT 6.288 0.924 8.784 3.528 ;
  LAYER M1 ;
        RECT 6.288 4.032 8.784 6.636 ;
  LAYER M3 ;
        RECT 6.288 4.032 8.784 6.636 ;
  LAYER M2 ;
        RECT 6.288 4.032 8.784 6.636 ;
  LAYER M1 ;
        RECT 6.288 7.14 8.784 9.744 ;
  LAYER M3 ;
        RECT 6.288 7.14 8.784 9.744 ;
  LAYER M2 ;
        RECT 6.288 7.14 8.784 9.744 ;
  LAYER M1 ;
        RECT 6.288 10.248 8.784 12.852 ;
  LAYER M3 ;
        RECT 6.288 10.248 8.784 12.852 ;
  LAYER M2 ;
        RECT 6.288 10.248 8.784 12.852 ;
  LAYER M1 ;
        RECT 6.288 13.356 8.784 15.96 ;
  LAYER M3 ;
        RECT 6.288 13.356 8.784 15.96 ;
  LAYER M2 ;
        RECT 6.288 13.356 8.784 15.96 ;
  LAYER M1 ;
        RECT 9.264 0.924 11.76 3.528 ;
  LAYER M3 ;
        RECT 9.264 0.924 11.76 3.528 ;
  LAYER M2 ;
        RECT 9.264 0.924 11.76 3.528 ;
  LAYER M1 ;
        RECT 9.264 4.032 11.76 6.636 ;
  LAYER M3 ;
        RECT 9.264 4.032 11.76 6.636 ;
  LAYER M2 ;
        RECT 9.264 4.032 11.76 6.636 ;
  LAYER M1 ;
        RECT 9.264 7.14 11.76 9.744 ;
  LAYER M3 ;
        RECT 9.264 7.14 11.76 9.744 ;
  LAYER M2 ;
        RECT 9.264 7.14 11.76 9.744 ;
  LAYER M1 ;
        RECT 9.264 10.248 11.76 12.852 ;
  LAYER M3 ;
        RECT 9.264 10.248 11.76 12.852 ;
  LAYER M2 ;
        RECT 9.264 10.248 11.76 12.852 ;
  LAYER M1 ;
        RECT 9.264 13.356 11.76 15.96 ;
  LAYER M3 ;
        RECT 9.264 13.356 11.76 15.96 ;
  LAYER M2 ;
        RECT 9.264 13.356 11.76 15.96 ;
  LAYER M1 ;
        RECT 12.24 0.924 14.736 3.528 ;
  LAYER M3 ;
        RECT 12.24 0.924 14.736 3.528 ;
  LAYER M2 ;
        RECT 12.24 0.924 14.736 3.528 ;
  LAYER M1 ;
        RECT 12.24 4.032 14.736 6.636 ;
  LAYER M3 ;
        RECT 12.24 4.032 14.736 6.636 ;
  LAYER M2 ;
        RECT 12.24 4.032 14.736 6.636 ;
  LAYER M1 ;
        RECT 12.24 7.14 14.736 9.744 ;
  LAYER M3 ;
        RECT 12.24 7.14 14.736 9.744 ;
  LAYER M2 ;
        RECT 12.24 7.14 14.736 9.744 ;
  LAYER M1 ;
        RECT 12.24 10.248 14.736 12.852 ;
  LAYER M3 ;
        RECT 12.24 10.248 14.736 12.852 ;
  LAYER M2 ;
        RECT 12.24 10.248 14.736 12.852 ;
  LAYER M1 ;
        RECT 12.24 13.356 14.736 15.96 ;
  LAYER M3 ;
        RECT 12.24 13.356 14.736 15.96 ;
  LAYER M2 ;
        RECT 12.24 13.356 14.736 15.96 ;
  LAYER M1 ;
        RECT 15.216 0.924 17.712 3.528 ;
  LAYER M3 ;
        RECT 15.216 0.924 17.712 3.528 ;
  LAYER M2 ;
        RECT 15.216 0.924 17.712 3.528 ;
  LAYER M1 ;
        RECT 15.216 4.032 17.712 6.636 ;
  LAYER M3 ;
        RECT 15.216 4.032 17.712 6.636 ;
  LAYER M2 ;
        RECT 15.216 4.032 17.712 6.636 ;
  LAYER M1 ;
        RECT 15.216 7.14 17.712 9.744 ;
  LAYER M3 ;
        RECT 15.216 7.14 17.712 9.744 ;
  LAYER M2 ;
        RECT 15.216 7.14 17.712 9.744 ;
  LAYER M1 ;
        RECT 15.216 10.248 17.712 12.852 ;
  LAYER M3 ;
        RECT 15.216 10.248 17.712 12.852 ;
  LAYER M2 ;
        RECT 15.216 10.248 17.712 12.852 ;
  LAYER M1 ;
        RECT 15.216 13.356 17.712 15.96 ;
  LAYER M3 ;
        RECT 15.216 13.356 17.712 15.96 ;
  LAYER M2 ;
        RECT 15.216 13.356 17.712 15.96 ;
  END 
END Cap_60fF_Cap_60fF
