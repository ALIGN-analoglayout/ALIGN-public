VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RES_w1u_l14u
  UNITS 
    DATABASE MICRONS UNITS 1 ;
  END UNITS 

  ORIGIN 0 0 ;
  FOREIGN RES_w1u_l14u 0 0 ;
  SIZE 14.54 BY 1.3 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0 0.15 0.32 1.15 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.22 0.15 14.54 1.15 ;
    END
  END MINUS
END RES_w1u_l14u

