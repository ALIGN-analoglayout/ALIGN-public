MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 18 BY 16.884 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
      LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
      LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
      LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
      LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
      LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
      LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
      LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
      LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
      LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
      LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
      LAYER M2 ;
        RECT 6.032 0.236 11.984 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M1 ;
        RECT 8.768 7.056 8.8 7.224 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M2 ;
        RECT 8.784 7.04 9.008 7.072 ;
  LAYER M1 ;
        RECT 8.992 7.02 9.024 7.092 ;
  LAYER M2 ;
        RECT 8.972 7.04 9.044 7.072 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M2 ;
        RECT 9.008 7.208 11.76 7.24 ;
  LAYER M1 ;
        RECT 8.992 7.188 9.024 7.26 ;
  LAYER M2 ;
        RECT 8.972 7.208 9.044 7.24 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.164 8.8 10.332 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M2 ;
        RECT 8.784 10.148 9.008 10.18 ;
  LAYER M1 ;
        RECT 8.992 10.128 9.024 10.2 ;
  LAYER M2 ;
        RECT 8.972 10.148 9.044 10.18 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M2 ;
        RECT 9.008 4.1 11.76 4.132 ;
  LAYER M1 ;
        RECT 8.992 4.08 9.024 4.152 ;
  LAYER M2 ;
        RECT 8.972 4.1 9.044 4.132 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M1 ;
        RECT 8.768 3.948 8.8 4.116 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 8.784 3.932 9.008 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M2 ;
        RECT 9.008 10.316 11.76 10.348 ;
  LAYER M1 ;
        RECT 8.992 10.296 9.024 10.368 ;
  LAYER M2 ;
        RECT 8.972 10.316 9.044 10.348 ;
  LAYER M1 ;
        RECT 8.992 0.384 9.024 0.456 ;
  LAYER M2 ;
        RECT 8.972 0.404 9.044 0.436 ;
  LAYER M1 ;
        RECT 8.992 0.42 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 10.332 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M1 ;
        RECT 5.792 7.056 5.824 7.224 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M2 ;
        RECT 5.808 7.04 6.032 7.072 ;
  LAYER M1 ;
        RECT 6.016 7.02 6.048 7.092 ;
  LAYER M2 ;
        RECT 5.996 7.04 6.068 7.072 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.164 5.824 10.332 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M1 ;
        RECT 5.792 3.948 5.824 4.116 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M2 ;
        RECT 5.808 3.932 6.032 3.964 ;
  LAYER M1 ;
        RECT 6.016 3.912 6.048 3.984 ;
  LAYER M2 ;
        RECT 5.996 3.932 6.068 3.964 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 10.164 ;
  LAYER M1 ;
        RECT 14.72 7.188 14.752 7.26 ;
  LAYER M2 ;
        RECT 14.7 7.208 14.772 7.24 ;
  LAYER M2 ;
        RECT 11.984 7.208 14.736 7.24 ;
  LAYER M1 ;
        RECT 11.968 7.188 12 7.26 ;
  LAYER M2 ;
        RECT 11.948 7.208 12.02 7.24 ;
  LAYER M1 ;
        RECT 14.72 4.08 14.752 4.152 ;
  LAYER M2 ;
        RECT 14.7 4.1 14.772 4.132 ;
  LAYER M2 ;
        RECT 11.984 4.1 14.736 4.132 ;
  LAYER M1 ;
        RECT 11.968 4.08 12 4.152 ;
  LAYER M2 ;
        RECT 11.948 4.1 12.02 4.132 ;
  LAYER M1 ;
        RECT 14.72 10.296 14.752 10.368 ;
  LAYER M2 ;
        RECT 14.7 10.316 14.772 10.348 ;
  LAYER M2 ;
        RECT 11.984 10.316 14.736 10.348 ;
  LAYER M1 ;
        RECT 11.968 10.296 12 10.368 ;
  LAYER M2 ;
        RECT 11.948 10.316 12.02 10.348 ;
  LAYER M1 ;
        RECT 11.968 0.216 12 0.288 ;
  LAYER M2 ;
        RECT 11.948 0.236 12.02 0.268 ;
  LAYER M1 ;
        RECT 11.968 0.252 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 10.332 ;
  LAYER M2 ;
        RECT 6.032 0.236 11.984 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.84 2.848 1.008 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M2 ;
        RECT 2.832 0.824 3.056 0.856 ;
  LAYER M1 ;
        RECT 3.04 0.804 3.072 0.876 ;
  LAYER M2 ;
        RECT 3.02 0.824 3.092 0.856 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M1 ;
        RECT 2.816 3.948 2.848 4.116 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M2 ;
        RECT 2.832 3.932 3.056 3.964 ;
  LAYER M1 ;
        RECT 3.04 3.912 3.072 3.984 ;
  LAYER M2 ;
        RECT 3.02 3.932 3.092 3.964 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M1 ;
        RECT 2.816 7.056 2.848 7.224 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M2 ;
        RECT 2.832 7.04 3.056 7.072 ;
  LAYER M1 ;
        RECT 3.04 7.02 3.072 7.092 ;
  LAYER M2 ;
        RECT 3.02 7.04 3.092 7.072 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M1 ;
        RECT 2.816 10.164 2.848 10.332 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M2 ;
        RECT 2.832 10.148 3.056 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M1 ;
        RECT 2.816 13.272 2.848 13.44 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 13.308 ;
  LAYER M2 ;
        RECT 2.796 13.256 2.868 13.288 ;
  LAYER M2 ;
        RECT 2.832 13.256 3.056 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 3.056 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 3.04 0.972 3.072 1.044 ;
  LAYER M2 ;
        RECT 3.02 0.992 3.092 1.024 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M2 ;
        RECT 3.056 13.424 5.808 13.456 ;
  LAYER M1 ;
        RECT 3.04 13.404 3.072 13.476 ;
  LAYER M2 ;
        RECT 3.02 13.424 3.092 13.456 ;
  LAYER M1 ;
        RECT 3.04 0.048 3.072 0.12 ;
  LAYER M2 ;
        RECT 3.02 0.068 3.092 0.1 ;
  LAYER M1 ;
        RECT 3.04 0.084 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 13.44 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.84 14.752 1.008 ;
  LAYER M1 ;
        RECT 14.72 0.804 14.752 0.876 ;
  LAYER M2 ;
        RECT 14.7 0.824 14.772 0.856 ;
  LAYER M2 ;
        RECT 14.736 0.824 14.96 0.856 ;
  LAYER M1 ;
        RECT 14.944 0.804 14.976 0.876 ;
  LAYER M2 ;
        RECT 14.924 0.824 14.996 0.856 ;
  LAYER M1 ;
        RECT 14.72 13.404 14.752 13.476 ;
  LAYER M2 ;
        RECT 14.7 13.424 14.772 13.456 ;
  LAYER M1 ;
        RECT 14.72 13.272 14.752 13.44 ;
  LAYER M1 ;
        RECT 14.72 13.236 14.752 13.308 ;
  LAYER M2 ;
        RECT 14.7 13.256 14.772 13.288 ;
  LAYER M2 ;
        RECT 14.736 13.256 14.96 13.288 ;
  LAYER M1 ;
        RECT 14.944 13.236 14.976 13.308 ;
  LAYER M2 ;
        RECT 14.924 13.256 14.996 13.288 ;
  LAYER M1 ;
        RECT 17.696 0.972 17.728 1.044 ;
  LAYER M2 ;
        RECT 17.676 0.992 17.748 1.024 ;
  LAYER M2 ;
        RECT 14.96 0.992 17.712 1.024 ;
  LAYER M1 ;
        RECT 14.944 0.972 14.976 1.044 ;
  LAYER M2 ;
        RECT 14.924 0.992 14.996 1.024 ;
  LAYER M1 ;
        RECT 17.696 4.08 17.728 4.152 ;
  LAYER M2 ;
        RECT 17.676 4.1 17.748 4.132 ;
  LAYER M2 ;
        RECT 14.96 4.1 17.712 4.132 ;
  LAYER M1 ;
        RECT 14.944 4.08 14.976 4.152 ;
  LAYER M2 ;
        RECT 14.924 4.1 14.996 4.132 ;
  LAYER M1 ;
        RECT 17.696 7.188 17.728 7.26 ;
  LAYER M2 ;
        RECT 17.676 7.208 17.748 7.24 ;
  LAYER M2 ;
        RECT 14.96 7.208 17.712 7.24 ;
  LAYER M1 ;
        RECT 14.944 7.188 14.976 7.26 ;
  LAYER M2 ;
        RECT 14.924 7.208 14.996 7.24 ;
  LAYER M1 ;
        RECT 17.696 10.296 17.728 10.368 ;
  LAYER M2 ;
        RECT 17.676 10.316 17.748 10.348 ;
  LAYER M2 ;
        RECT 14.96 10.316 17.712 10.348 ;
  LAYER M1 ;
        RECT 14.944 10.296 14.976 10.368 ;
  LAYER M2 ;
        RECT 14.924 10.316 14.996 10.348 ;
  LAYER M1 ;
        RECT 17.696 13.404 17.728 13.476 ;
  LAYER M2 ;
        RECT 17.676 13.424 17.748 13.456 ;
  LAYER M2 ;
        RECT 14.96 13.424 17.712 13.456 ;
  LAYER M1 ;
        RECT 14.944 13.404 14.976 13.476 ;
  LAYER M2 ;
        RECT 14.924 13.424 14.996 13.456 ;
  LAYER M1 ;
        RECT 14.944 0.048 14.976 0.12 ;
  LAYER M2 ;
        RECT 14.924 0.068 14.996 0.1 ;
  LAYER M1 ;
        RECT 14.944 0.084 14.976 0.672 ;
  LAYER M1 ;
        RECT 14.944 0.672 14.976 13.44 ;
  LAYER M2 ;
        RECT 3.056 0.068 14.96 0.1 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M2 ;
        RECT 5.808 13.424 8.784 13.456 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 13.476 ;
  LAYER M2 ;
        RECT 11.724 13.424 11.796 13.456 ;
  LAYER M2 ;
        RECT 8.784 13.424 11.76 13.456 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M2 ;
        RECT 11.76 0.992 14.736 1.024 ;
  LAYER M1 ;
        RECT 14.72 0.972 14.752 1.044 ;
  LAYER M2 ;
        RECT 14.7 0.992 14.772 1.024 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M2 ;
        RECT 6.192 9.644 6.416 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 6.192 12.752 6.416 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.416 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 6.176 16.428 6.208 16.5 ;
  LAYER M2 ;
        RECT 6.156 16.448 6.228 16.48 ;
  LAYER M1 ;
        RECT 6.176 16.212 6.208 16.464 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 16.212 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M1 ;
        RECT 9.376 9.66 9.408 9.828 ;
  LAYER M1 ;
        RECT 9.376 9.792 9.408 9.864 ;
  LAYER M2 ;
        RECT 9.356 9.812 9.428 9.844 ;
  LAYER M2 ;
        RECT 9.392 9.812 12.144 9.844 ;
  LAYER M1 ;
        RECT 12.128 9.792 12.16 9.864 ;
  LAYER M2 ;
        RECT 12.108 9.812 12.18 9.844 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.376 6.552 9.408 6.72 ;
  LAYER M1 ;
        RECT 9.376 6.684 9.408 6.756 ;
  LAYER M2 ;
        RECT 9.356 6.704 9.428 6.736 ;
  LAYER M2 ;
        RECT 9.392 6.704 12.144 6.736 ;
  LAYER M1 ;
        RECT 12.128 6.684 12.16 6.756 ;
  LAYER M2 ;
        RECT 12.108 6.704 12.18 6.736 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M1 ;
        RECT 9.376 12.768 9.408 12.936 ;
  LAYER M1 ;
        RECT 9.376 12.9 9.408 12.972 ;
  LAYER M2 ;
        RECT 9.356 12.92 9.428 12.952 ;
  LAYER M2 ;
        RECT 9.392 12.92 12.144 12.952 ;
  LAYER M1 ;
        RECT 12.128 12.9 12.16 12.972 ;
  LAYER M2 ;
        RECT 12.108 12.92 12.18 12.952 ;
  LAYER M1 ;
        RECT 12.128 16.428 12.16 16.5 ;
  LAYER M2 ;
        RECT 12.108 16.448 12.18 16.48 ;
  LAYER M1 ;
        RECT 12.128 16.212 12.16 16.464 ;
  LAYER M1 ;
        RECT 12.128 6.72 12.16 16.212 ;
  LAYER M2 ;
        RECT 6.192 16.448 12.144 16.48 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.216 9.644 3.44 9.676 ;
  LAYER M1 ;
        RECT 3.2 9.624 3.232 9.696 ;
  LAYER M2 ;
        RECT 3.18 9.644 3.252 9.676 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 3.216 6.536 3.44 6.568 ;
  LAYER M1 ;
        RECT 3.2 6.516 3.232 6.588 ;
  LAYER M2 ;
        RECT 3.18 6.536 3.252 6.568 ;
  LAYER M1 ;
        RECT 3.2 16.596 3.232 16.668 ;
  LAYER M2 ;
        RECT 3.18 16.616 3.252 16.648 ;
  LAYER M1 ;
        RECT 3.2 16.212 3.232 16.632 ;
  LAYER M1 ;
        RECT 3.2 6.552 3.232 16.212 ;
  LAYER M1 ;
        RECT 12.352 9.624 12.384 9.696 ;
  LAYER M2 ;
        RECT 12.332 9.644 12.404 9.676 ;
  LAYER M1 ;
        RECT 12.352 9.66 12.384 9.828 ;
  LAYER M1 ;
        RECT 12.352 9.792 12.384 9.864 ;
  LAYER M2 ;
        RECT 12.332 9.812 12.404 9.844 ;
  LAYER M2 ;
        RECT 12.368 9.812 15.12 9.844 ;
  LAYER M1 ;
        RECT 15.104 9.792 15.136 9.864 ;
  LAYER M2 ;
        RECT 15.084 9.812 15.156 9.844 ;
  LAYER M1 ;
        RECT 12.352 6.516 12.384 6.588 ;
  LAYER M2 ;
        RECT 12.332 6.536 12.404 6.568 ;
  LAYER M1 ;
        RECT 12.352 6.552 12.384 6.72 ;
  LAYER M1 ;
        RECT 12.352 6.684 12.384 6.756 ;
  LAYER M2 ;
        RECT 12.332 6.704 12.404 6.736 ;
  LAYER M2 ;
        RECT 12.368 6.704 15.12 6.736 ;
  LAYER M1 ;
        RECT 15.104 6.684 15.136 6.756 ;
  LAYER M2 ;
        RECT 15.084 6.704 15.156 6.736 ;
  LAYER M1 ;
        RECT 12.352 12.732 12.384 12.804 ;
  LAYER M2 ;
        RECT 12.332 12.752 12.404 12.784 ;
  LAYER M1 ;
        RECT 12.352 12.768 12.384 12.936 ;
  LAYER M1 ;
        RECT 12.352 12.9 12.384 12.972 ;
  LAYER M2 ;
        RECT 12.332 12.92 12.404 12.952 ;
  LAYER M2 ;
        RECT 12.368 12.92 15.12 12.952 ;
  LAYER M1 ;
        RECT 15.104 12.9 15.136 12.972 ;
  LAYER M2 ;
        RECT 15.084 12.92 15.156 12.952 ;
  LAYER M1 ;
        RECT 15.104 16.596 15.136 16.668 ;
  LAYER M2 ;
        RECT 15.084 16.616 15.156 16.648 ;
  LAYER M1 ;
        RECT 15.104 16.212 15.136 16.632 ;
  LAYER M1 ;
        RECT 15.104 6.72 15.136 16.212 ;
  LAYER M2 ;
        RECT 3.216 16.616 15.12 16.648 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.08 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.064 3.408 0.096 3.48 ;
  LAYER M2 ;
        RECT 0.044 3.428 0.116 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.08 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.064 6.516 0.096 6.588 ;
  LAYER M2 ;
        RECT 0.044 6.536 0.116 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.08 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.064 9.624 0.096 9.696 ;
  LAYER M2 ;
        RECT 0.044 9.644 0.116 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.08 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.064 12.732 0.096 12.804 ;
  LAYER M2 ;
        RECT 0.044 12.752 0.116 12.784 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M2 ;
        RECT 0.08 15.86 0.464 15.892 ;
  LAYER M1 ;
        RECT 0.064 15.84 0.096 15.912 ;
  LAYER M2 ;
        RECT 0.044 15.86 0.116 15.892 ;
  LAYER M1 ;
        RECT 0.064 16.764 0.096 16.836 ;
  LAYER M2 ;
        RECT 0.044 16.784 0.116 16.816 ;
  LAYER M1 ;
        RECT 0.064 16.212 0.096 16.8 ;
  LAYER M1 ;
        RECT 0.064 3.444 0.096 16.212 ;
  LAYER M1 ;
        RECT 15.328 3.408 15.36 3.48 ;
  LAYER M2 ;
        RECT 15.308 3.428 15.38 3.46 ;
  LAYER M1 ;
        RECT 15.328 3.444 15.36 3.612 ;
  LAYER M1 ;
        RECT 15.328 3.576 15.36 3.648 ;
  LAYER M2 ;
        RECT 15.308 3.596 15.38 3.628 ;
  LAYER M2 ;
        RECT 15.344 3.596 17.936 3.628 ;
  LAYER M1 ;
        RECT 17.92 3.576 17.952 3.648 ;
  LAYER M2 ;
        RECT 17.9 3.596 17.972 3.628 ;
  LAYER M1 ;
        RECT 15.328 6.516 15.36 6.588 ;
  LAYER M2 ;
        RECT 15.308 6.536 15.38 6.568 ;
  LAYER M1 ;
        RECT 15.328 6.552 15.36 6.72 ;
  LAYER M1 ;
        RECT 15.328 6.684 15.36 6.756 ;
  LAYER M2 ;
        RECT 15.308 6.704 15.38 6.736 ;
  LAYER M2 ;
        RECT 15.344 6.704 17.936 6.736 ;
  LAYER M1 ;
        RECT 17.92 6.684 17.952 6.756 ;
  LAYER M2 ;
        RECT 17.9 6.704 17.972 6.736 ;
  LAYER M1 ;
        RECT 15.328 9.624 15.36 9.696 ;
  LAYER M2 ;
        RECT 15.308 9.644 15.38 9.676 ;
  LAYER M1 ;
        RECT 15.328 9.66 15.36 9.828 ;
  LAYER M1 ;
        RECT 15.328 9.792 15.36 9.864 ;
  LAYER M2 ;
        RECT 15.308 9.812 15.38 9.844 ;
  LAYER M2 ;
        RECT 15.344 9.812 17.936 9.844 ;
  LAYER M1 ;
        RECT 17.92 9.792 17.952 9.864 ;
  LAYER M2 ;
        RECT 17.9 9.812 17.972 9.844 ;
  LAYER M1 ;
        RECT 15.328 12.732 15.36 12.804 ;
  LAYER M2 ;
        RECT 15.308 12.752 15.38 12.784 ;
  LAYER M1 ;
        RECT 15.328 12.768 15.36 12.936 ;
  LAYER M1 ;
        RECT 15.328 12.9 15.36 12.972 ;
  LAYER M2 ;
        RECT 15.308 12.92 15.38 12.952 ;
  LAYER M2 ;
        RECT 15.344 12.92 17.936 12.952 ;
  LAYER M1 ;
        RECT 17.92 12.9 17.952 12.972 ;
  LAYER M2 ;
        RECT 17.9 12.92 17.972 12.952 ;
  LAYER M1 ;
        RECT 15.328 15.84 15.36 15.912 ;
  LAYER M2 ;
        RECT 15.308 15.86 15.38 15.892 ;
  LAYER M1 ;
        RECT 15.328 15.876 15.36 16.044 ;
  LAYER M1 ;
        RECT 15.328 16.008 15.36 16.08 ;
  LAYER M2 ;
        RECT 15.308 16.028 15.38 16.06 ;
  LAYER M2 ;
        RECT 15.344 16.028 17.936 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.008 17.952 16.08 ;
  LAYER M2 ;
        RECT 17.9 16.028 17.972 16.06 ;
  LAYER M1 ;
        RECT 17.92 16.764 17.952 16.836 ;
  LAYER M2 ;
        RECT 17.9 16.784 17.972 16.816 ;
  LAYER M1 ;
        RECT 17.92 16.212 17.952 16.8 ;
  LAYER M1 ;
        RECT 17.92 3.612 17.952 16.212 ;
  LAYER M2 ;
        RECT 0.08 16.784 17.936 16.816 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 0.464 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M2 ;
        RECT 3.44 15.86 6.416 15.892 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M2 ;
        RECT 6.416 15.86 9.392 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M1 ;
        RECT 12.352 15.84 12.384 15.912 ;
  LAYER M2 ;
        RECT 12.332 15.86 12.404 15.892 ;
  LAYER M2 ;
        RECT 9.392 15.86 12.368 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M2 ;
        RECT 12.368 3.428 15.344 3.46 ;
  LAYER M1 ;
        RECT 15.328 3.408 15.36 3.48 ;
  LAYER M2 ;
        RECT 15.308 3.428 15.38 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M2 ;
        RECT 9.392 3.428 12.368 3.46 ;
  LAYER M1 ;
        RECT 12.352 3.408 12.384 3.48 ;
  LAYER M2 ;
        RECT 12.332 3.428 12.404 3.46 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M3 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M3 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M3 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M3 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M2 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M1 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M3 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M3 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M3 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M3 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M3 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M2 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M1 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M3 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M3 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M3 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M3 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M3 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M2 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M1 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M3 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M3 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M3 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M3 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M3 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M2 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M1 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M3 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M2 ;
        RECT 12.304 0.924 14.8 3.528 ;
  LAYER M1 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M3 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M2 ;
        RECT 12.304 4.032 14.8 6.636 ;
  LAYER M1 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M3 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M2 ;
        RECT 12.304 7.14 14.8 9.744 ;
  LAYER M1 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M3 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M2 ;
        RECT 12.304 10.248 14.8 12.852 ;
  LAYER M1 ;
        RECT 12.304 13.356 14.8 15.96 ;
  LAYER M3 ;
        RECT 12.304 13.356 14.8 15.96 ;
  LAYER M2 ;
        RECT 12.304 13.356 14.8 15.96 ;
  LAYER M1 ;
        RECT 15.28 0.924 17.776 3.528 ;
  LAYER M3 ;
        RECT 15.28 0.924 17.776 3.528 ;
  LAYER M2 ;
        RECT 15.28 0.924 17.776 3.528 ;
  LAYER M1 ;
        RECT 15.28 4.032 17.776 6.636 ;
  LAYER M3 ;
        RECT 15.28 4.032 17.776 6.636 ;
  LAYER M2 ;
        RECT 15.28 4.032 17.776 6.636 ;
  LAYER M1 ;
        RECT 15.28 7.14 17.776 9.744 ;
  LAYER M3 ;
        RECT 15.28 7.14 17.776 9.744 ;
  LAYER M2 ;
        RECT 15.28 7.14 17.776 9.744 ;
  LAYER M1 ;
        RECT 15.28 10.248 17.776 12.852 ;
  LAYER M3 ;
        RECT 15.28 10.248 17.776 12.852 ;
  LAYER M2 ;
        RECT 15.28 10.248 17.776 12.852 ;
  LAYER M1 ;
        RECT 15.28 13.356 17.776 15.96 ;
  LAYER M3 ;
        RECT 15.28 13.356 17.776 15.96 ;
  LAYER M2 ;
        RECT 15.28 13.356 17.776 15.96 ;
  END 
END Cap_60fF_Cap_60fF
