.model plplvt pmos w=1 l=1 nfin=1 nf=1 m=1
.subckt powertrain vcc vg vout
mmp0 vout vg vcc vcc plplvt w=180n l=40n nfin=4 nf=8 m=20
.ends
