
.subckt Sanitized_CK_Divider8 PRESET VDD VSS CKIN COMPEN QPHASE OUTPHASE INPHASE
XI14 PRESET VDD VSS net039 INVD2LVT
XI51<18> VDD VSS DCAP8LVT
XI51<17> VDD VSS DCAP8LVT
XI51<16> VDD VSS DCAP8LVT
XI51<15> VDD VSS DCAP8LVT
XI51<14> VDD VSS DCAP8LVT
XI51<13> VDD VSS DCAP8LVT
XI51<12> VDD VSS DCAP8LVT
XI51<11> VDD VSS DCAP8LVT
XI51<10> VDD VSS DCAP8LVT
XI51<9> VDD VSS DCAP8LVT
XI51<8> VDD VSS DCAP8LVT
XI51<7> VDD VSS DCAP8LVT
XI51<6> VDD VSS DCAP8LVT
XI51<5> VDD VSS DCAP8LVT
XI51<4> VDD VSS DCAP8LVT
XI51<3> VDD VSS DCAP8LVT
XI51<2> VDD VSS DCAP8LVT
XI51<1> VDD VSS DCAP8LVT
XI51<0> VDD VSS DCAP8LVT
XI50 PRESET VDD VSS net048 INVD1LVT
XI6 CKIN VDD VSS net45 CKBD1LVT
XI139 net048 net015 VDD VSS COMPEN AN2D1LVT
XI5 net45 VDD VSS net49 CKND1LVT
XI8 net039 net011 net48 net015 net48 VDD VSS DFCND1LVT
XI7 net039 net018 net50 net076 net50 VDD VSS DFCND1LVT
XI43 net076 VDD VSS net059 CKND3LVT
XI39 net48 VDD VSS net063 CKND3LVT
XI37 net015 VDD VSS net064 CKND3LVT
XI42 net059 VDD VSS QPHASE CKND8LVT
XI38 net063 VDD VSS OUTPHASE CKND8LVT
XI20 net064 VDD VSS INPHASE CKND8LVT
XI29 net039 net49 net016 net016 VDD VSS DFCND1LVT_schematic
XI28 net039 net016 net018 net018 VDD VSS DFCND1LVT_schematic
XI27 net039 net45 net040 net040 VDD VSS DFCND1LVT_schematic
XI26 net039 net040 net011 net011 VDD VSS DFCND1LVT_schematic
.ends Sanitized_CK_Divider8

.subckt INVD2LVT I VDD VSS ZN
xMMU1_0_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_0_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD2LVT

.subckt Switch_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=2
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=2
.ends Switch_NMOS_n12_X1_Y1

.subckt Switch_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=2
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=2
.ends Switch_PMOS_n12_X1_Y1

.subckt DCAP8LVT VDD VSS
xMMI4 VSS net9 VSS Dcap_NMOS_n12_X1_Y1
xMM_u2 net11 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI3 VDD net11 VDD Dcap_PMOS_n12_X1_Y1
xMM_u1 net9 net11 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DCAP8LVT

.subckt Dcap_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_NMOS_n12_X1_Y1

.subckt Dcap_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_PMOS_n12_X1_Y1

.subckt INVD1LVT I VDD VSS ZN
xMMU1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD1LVT

.subckt INV_LVT zn i SN SP
xxm0 zn i SN SN Switch_NMOS_n12_X1_Y1
xxm1 zn i SP SP Switch_PMOS_n12_X1_Y1
.ends INV_LVT

.subckt stage2_inv G1 SN G2 SP
MM0_MM2 D SN SP G1 INV_LVT
MM1_MM3 G2 SN SP D INV_LVT
.ends stage2_inv

.subckt CKBD1LVT I VDD VSS Z
MMU23_MM_u15_MMU21_MM_u3 VSS I VDD Z stage2_inv
.ends CKBD1LVT

.subckt AN2D1LVT A1 A2 VDD VSS Z
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u4 net17 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net17 VSS Switch_NMOS_n12_X1_Y1
.ends AN2D1LVT

.subckt CKND1LVT I VDD VSS ZN
xMM_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u1 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKND1LVT

.subckt tgate D GA S GB
xM0 D GA S BN Switch_NMOS_n12_X1_Y1
xM1 D GB S BP Switch_PMOS_n12_X1_Y1
.ends tgate

.subckt DFCND1LVT CDN CP D Q QN VDD VSS
xMMI4 net53 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u3 net95 net79 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net81 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net25 D net53 VSS Switch_NMOS_n12_X1_Y1
xMMI49 net20 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net17 net81 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 Q net95 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u4 net9 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net25 net67 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI43 net72 net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net25 D net104 VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 Q net95 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI44 net72 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net81 net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u1 net95 net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI45 net25 net5 net72 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net104 net67 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u2 net95 CDN VDD VDD Switch_PMOS_n12_X1_Y1
MMI32_M_u2_MMI22_M_u2_MMI32_M_u3_MMI22_M_u3 VSS CP VDD net67 stage2_inv
MMI29_M_u2_MMI14_M_u2_MMI29_M_u3_MMI14_M_u3 VSS net95 VDD QN stage2_inv
MMI15_MMI16 net67 net79 net5 net81 tgate
MMI18_MMI17 net5 net79 net67 net33 tgate
.ends DFCND1LVT

.subckt CKND3LVT I VDD VSS ZN
xMM_u1_0 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u1_1 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_1 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
.ends CKND3LVT

.subckt CKND8LVT I VDD VSS ZN
xMM_u1_1 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
.ends CKND8LVT

.subckt DFCND1LVT_schematic CDN CP D QN VDD VSS
xMMI4 net53 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u3 net95 net79 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net81 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net25 D net53 VSS Switch_NMOS_n12_X1_Y1
xMMI49 net20 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net17 net81 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 net036 net95 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u4 net9 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net25 net67 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI43 net72 net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net25 D net104 VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 net036 net95 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI44 net72 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net81 net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u1 net95 net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI45 net25 net5 net72 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net104 net67 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u2 net95 CDN VDD VDD Switch_PMOS_n12_X1_Y1
MMI32_M_u2_MMI22_M_u2_MMI32_M_u3_MMI22_M_u3 VSS CP VDD net67 stage2_inv
MMI29_M_u2_MMI14_M_u2_MMI29_M_u3_MMI14_M_u3 VSS net95 VDD QN stage2_inv
MMI15_MMI16 net67 net79 net5 net81 tgate
MMI18_MMI17 net5 net79 net67 net33 tgate
.ends DFCND1LVT_schematic
