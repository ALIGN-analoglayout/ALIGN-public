MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 9.92 BY 33.684 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.584 33.228 3.616 33.3 ;
      LAYER M2 ;
        RECT 3.564 33.248 3.636 33.28 ;
      LAYER M1 ;
        RECT 6.784 33.228 6.816 33.3 ;
      LAYER M2 ;
        RECT 6.764 33.248 6.836 33.28 ;
      LAYER M2 ;
        RECT 3.6 33.248 6.8 33.28 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.264 0.384 3.296 0.456 ;
      LAYER M2 ;
        RECT 3.244 0.404 3.316 0.436 ;
      LAYER M1 ;
        RECT 6.464 0.384 6.496 0.456 ;
      LAYER M2 ;
        RECT 6.444 0.404 6.516 0.436 ;
      LAYER M2 ;
        RECT 3.28 0.404 6.48 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.744 33.396 3.776 33.468 ;
      LAYER M2 ;
        RECT 3.724 33.416 3.796 33.448 ;
      LAYER M1 ;
        RECT 6.944 33.396 6.976 33.468 ;
      LAYER M2 ;
        RECT 6.924 33.416 6.996 33.448 ;
      LAYER M2 ;
        RECT 3.76 33.416 6.96 33.448 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.424 0.216 3.456 0.288 ;
      LAYER M2 ;
        RECT 3.404 0.236 3.476 0.268 ;
      LAYER M1 ;
        RECT 6.624 0.216 6.656 0.288 ;
      LAYER M2 ;
        RECT 6.604 0.236 6.676 0.268 ;
      LAYER M2 ;
        RECT 3.44 0.236 6.64 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.304 15.588 6.336 15.66 ;
  LAYER M2 ;
        RECT 6.284 15.608 6.356 15.64 ;
  LAYER M2 ;
        RECT 3.28 15.608 6.32 15.64 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M1 ;
        RECT 6.304 3.828 6.336 3.9 ;
  LAYER M2 ;
        RECT 6.284 3.848 6.356 3.88 ;
  LAYER M2 ;
        RECT 3.28 3.848 6.32 3.88 ;
  LAYER M1 ;
        RECT 3.264 3.828 3.296 3.9 ;
  LAYER M2 ;
        RECT 3.244 3.848 3.316 3.88 ;
  LAYER M1 ;
        RECT 6.304 27.348 6.336 27.42 ;
  LAYER M2 ;
        RECT 6.284 27.368 6.356 27.4 ;
  LAYER M2 ;
        RECT 3.28 27.368 6.32 27.4 ;
  LAYER M1 ;
        RECT 3.264 27.348 3.296 27.42 ;
  LAYER M2 ;
        RECT 3.244 27.368 3.316 27.4 ;
  LAYER M1 ;
        RECT 3.264 0.384 3.296 0.456 ;
  LAYER M2 ;
        RECT 3.244 0.404 3.316 0.436 ;
  LAYER M1 ;
        RECT 3.264 0.42 3.296 0.588 ;
  LAYER M1 ;
        RECT 3.264 0.588 3.296 27.384 ;
  LAYER M1 ;
        RECT 6.304 15.588 6.336 15.66 ;
  LAYER M2 ;
        RECT 6.284 15.608 6.356 15.64 ;
  LAYER M1 ;
        RECT 6.304 15.456 6.336 15.624 ;
  LAYER M1 ;
        RECT 6.304 15.42 6.336 15.492 ;
  LAYER M2 ;
        RECT 6.284 15.44 6.356 15.472 ;
  LAYER M2 ;
        RECT 6.32 15.44 6.48 15.472 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 15.492 ;
  LAYER M2 ;
        RECT 6.444 15.44 6.516 15.472 ;
  LAYER M1 ;
        RECT 6.304 3.828 6.336 3.9 ;
  LAYER M2 ;
        RECT 6.284 3.848 6.356 3.88 ;
  LAYER M1 ;
        RECT 6.304 3.696 6.336 3.864 ;
  LAYER M1 ;
        RECT 6.304 3.66 6.336 3.732 ;
  LAYER M2 ;
        RECT 6.284 3.68 6.356 3.712 ;
  LAYER M2 ;
        RECT 6.32 3.68 6.48 3.712 ;
  LAYER M1 ;
        RECT 6.464 3.66 6.496 3.732 ;
  LAYER M2 ;
        RECT 6.444 3.68 6.516 3.712 ;
  LAYER M1 ;
        RECT 6.304 27.348 6.336 27.42 ;
  LAYER M2 ;
        RECT 6.284 27.368 6.356 27.4 ;
  LAYER M1 ;
        RECT 6.304 27.216 6.336 27.384 ;
  LAYER M1 ;
        RECT 6.304 27.18 6.336 27.252 ;
  LAYER M2 ;
        RECT 6.284 27.2 6.356 27.232 ;
  LAYER M2 ;
        RECT 6.32 27.2 6.48 27.232 ;
  LAYER M1 ;
        RECT 6.464 27.18 6.496 27.252 ;
  LAYER M2 ;
        RECT 6.444 27.2 6.516 27.232 ;
  LAYER M1 ;
        RECT 6.464 0.384 6.496 0.456 ;
  LAYER M2 ;
        RECT 6.444 0.404 6.516 0.436 ;
  LAYER M1 ;
        RECT 6.464 0.42 6.496 0.588 ;
  LAYER M1 ;
        RECT 6.464 0.588 6.496 27.216 ;
  LAYER M2 ;
        RECT 3.28 0.404 6.48 0.436 ;
  LAYER M1 ;
        RECT 6.304 12.648 6.336 12.72 ;
  LAYER M2 ;
        RECT 6.284 12.668 6.356 12.7 ;
  LAYER M2 ;
        RECT 3.44 12.668 6.32 12.7 ;
  LAYER M1 ;
        RECT 3.424 12.648 3.456 12.72 ;
  LAYER M2 ;
        RECT 3.404 12.668 3.476 12.7 ;
  LAYER M1 ;
        RECT 6.304 18.528 6.336 18.6 ;
  LAYER M2 ;
        RECT 6.284 18.548 6.356 18.58 ;
  LAYER M2 ;
        RECT 3.44 18.548 6.32 18.58 ;
  LAYER M1 ;
        RECT 3.424 18.528 3.456 18.6 ;
  LAYER M2 ;
        RECT 3.404 18.548 3.476 18.58 ;
  LAYER M1 ;
        RECT 6.304 9.708 6.336 9.78 ;
  LAYER M2 ;
        RECT 6.284 9.728 6.356 9.76 ;
  LAYER M2 ;
        RECT 3.44 9.728 6.32 9.76 ;
  LAYER M1 ;
        RECT 3.424 9.708 3.456 9.78 ;
  LAYER M2 ;
        RECT 3.404 9.728 3.476 9.76 ;
  LAYER M1 ;
        RECT 6.304 21.468 6.336 21.54 ;
  LAYER M2 ;
        RECT 6.284 21.488 6.356 21.52 ;
  LAYER M2 ;
        RECT 3.44 21.488 6.32 21.52 ;
  LAYER M1 ;
        RECT 3.424 21.468 3.456 21.54 ;
  LAYER M2 ;
        RECT 3.404 21.488 3.476 21.52 ;
  LAYER M1 ;
        RECT 6.304 6.768 6.336 6.84 ;
  LAYER M2 ;
        RECT 6.284 6.788 6.356 6.82 ;
  LAYER M2 ;
        RECT 3.44 6.788 6.32 6.82 ;
  LAYER M1 ;
        RECT 3.424 6.768 3.456 6.84 ;
  LAYER M2 ;
        RECT 3.404 6.788 3.476 6.82 ;
  LAYER M1 ;
        RECT 6.304 24.408 6.336 24.48 ;
  LAYER M2 ;
        RECT 6.284 24.428 6.356 24.46 ;
  LAYER M2 ;
        RECT 3.44 24.428 6.32 24.46 ;
  LAYER M1 ;
        RECT 3.424 24.408 3.456 24.48 ;
  LAYER M2 ;
        RECT 3.404 24.428 3.476 24.46 ;
  LAYER M1 ;
        RECT 3.424 0.216 3.456 0.288 ;
  LAYER M2 ;
        RECT 3.404 0.236 3.476 0.268 ;
  LAYER M1 ;
        RECT 3.424 0.252 3.456 0.588 ;
  LAYER M1 ;
        RECT 3.424 0.588 3.456 24.444 ;
  LAYER M1 ;
        RECT 6.304 12.648 6.336 12.72 ;
  LAYER M2 ;
        RECT 6.284 12.668 6.356 12.7 ;
  LAYER M1 ;
        RECT 6.304 12.516 6.336 12.684 ;
  LAYER M1 ;
        RECT 6.304 12.48 6.336 12.552 ;
  LAYER M2 ;
        RECT 6.284 12.5 6.356 12.532 ;
  LAYER M2 ;
        RECT 6.32 12.5 6.64 12.532 ;
  LAYER M1 ;
        RECT 6.624 12.48 6.656 12.552 ;
  LAYER M2 ;
        RECT 6.604 12.5 6.676 12.532 ;
  LAYER M1 ;
        RECT 6.304 18.528 6.336 18.6 ;
  LAYER M2 ;
        RECT 6.284 18.548 6.356 18.58 ;
  LAYER M1 ;
        RECT 6.304 18.396 6.336 18.564 ;
  LAYER M1 ;
        RECT 6.304 18.36 6.336 18.432 ;
  LAYER M2 ;
        RECT 6.284 18.38 6.356 18.412 ;
  LAYER M2 ;
        RECT 6.32 18.38 6.64 18.412 ;
  LAYER M1 ;
        RECT 6.624 18.36 6.656 18.432 ;
  LAYER M2 ;
        RECT 6.604 18.38 6.676 18.412 ;
  LAYER M1 ;
        RECT 6.304 9.708 6.336 9.78 ;
  LAYER M2 ;
        RECT 6.284 9.728 6.356 9.76 ;
  LAYER M1 ;
        RECT 6.304 9.576 6.336 9.744 ;
  LAYER M1 ;
        RECT 6.304 9.54 6.336 9.612 ;
  LAYER M2 ;
        RECT 6.284 9.56 6.356 9.592 ;
  LAYER M2 ;
        RECT 6.32 9.56 6.64 9.592 ;
  LAYER M1 ;
        RECT 6.624 9.54 6.656 9.612 ;
  LAYER M2 ;
        RECT 6.604 9.56 6.676 9.592 ;
  LAYER M1 ;
        RECT 6.304 21.468 6.336 21.54 ;
  LAYER M2 ;
        RECT 6.284 21.488 6.356 21.52 ;
  LAYER M1 ;
        RECT 6.304 21.336 6.336 21.504 ;
  LAYER M1 ;
        RECT 6.304 21.3 6.336 21.372 ;
  LAYER M2 ;
        RECT 6.284 21.32 6.356 21.352 ;
  LAYER M2 ;
        RECT 6.32 21.32 6.64 21.352 ;
  LAYER M1 ;
        RECT 6.624 21.3 6.656 21.372 ;
  LAYER M2 ;
        RECT 6.604 21.32 6.676 21.352 ;
  LAYER M1 ;
        RECT 6.304 6.768 6.336 6.84 ;
  LAYER M2 ;
        RECT 6.284 6.788 6.356 6.82 ;
  LAYER M1 ;
        RECT 6.304 6.636 6.336 6.804 ;
  LAYER M1 ;
        RECT 6.304 6.6 6.336 6.672 ;
  LAYER M2 ;
        RECT 6.284 6.62 6.356 6.652 ;
  LAYER M2 ;
        RECT 6.32 6.62 6.64 6.652 ;
  LAYER M1 ;
        RECT 6.624 6.6 6.656 6.672 ;
  LAYER M2 ;
        RECT 6.604 6.62 6.676 6.652 ;
  LAYER M1 ;
        RECT 6.304 24.408 6.336 24.48 ;
  LAYER M2 ;
        RECT 6.284 24.428 6.356 24.46 ;
  LAYER M1 ;
        RECT 6.304 24.276 6.336 24.444 ;
  LAYER M1 ;
        RECT 6.304 24.24 6.336 24.312 ;
  LAYER M2 ;
        RECT 6.284 24.26 6.356 24.292 ;
  LAYER M2 ;
        RECT 6.32 24.26 6.64 24.292 ;
  LAYER M1 ;
        RECT 6.624 24.24 6.656 24.312 ;
  LAYER M2 ;
        RECT 6.604 24.26 6.676 24.292 ;
  LAYER M1 ;
        RECT 6.624 0.216 6.656 0.288 ;
  LAYER M2 ;
        RECT 6.604 0.236 6.676 0.268 ;
  LAYER M1 ;
        RECT 6.624 0.252 6.656 0.588 ;
  LAYER M1 ;
        RECT 6.624 0.588 6.656 24.276 ;
  LAYER M2 ;
        RECT 3.44 0.236 6.64 0.268 ;
  LAYER M1 ;
        RECT 3.104 0.888 3.136 0.96 ;
  LAYER M2 ;
        RECT 3.084 0.908 3.156 0.94 ;
  LAYER M2 ;
        RECT 0.08 0.908 3.12 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 3.104 3.828 3.136 3.9 ;
  LAYER M2 ;
        RECT 3.084 3.848 3.156 3.88 ;
  LAYER M2 ;
        RECT 0.08 3.848 3.12 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 3.104 6.768 3.136 6.84 ;
  LAYER M2 ;
        RECT 3.084 6.788 3.156 6.82 ;
  LAYER M2 ;
        RECT 0.08 6.788 3.12 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 3.104 9.708 3.136 9.78 ;
  LAYER M2 ;
        RECT 3.084 9.728 3.156 9.76 ;
  LAYER M2 ;
        RECT 0.08 9.728 3.12 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 3.104 12.648 3.136 12.72 ;
  LAYER M2 ;
        RECT 3.084 12.668 3.156 12.7 ;
  LAYER M2 ;
        RECT 0.08 12.668 3.12 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 3.104 15.588 3.136 15.66 ;
  LAYER M2 ;
        RECT 3.084 15.608 3.156 15.64 ;
  LAYER M2 ;
        RECT 0.08 15.608 3.12 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 3.104 18.528 3.136 18.6 ;
  LAYER M2 ;
        RECT 3.084 18.548 3.156 18.58 ;
  LAYER M2 ;
        RECT 0.08 18.548 3.12 18.58 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M1 ;
        RECT 3.104 21.468 3.136 21.54 ;
  LAYER M2 ;
        RECT 3.084 21.488 3.156 21.52 ;
  LAYER M2 ;
        RECT 0.08 21.488 3.12 21.52 ;
  LAYER M1 ;
        RECT 0.064 21.468 0.096 21.54 ;
  LAYER M2 ;
        RECT 0.044 21.488 0.116 21.52 ;
  LAYER M1 ;
        RECT 3.104 24.408 3.136 24.48 ;
  LAYER M2 ;
        RECT 3.084 24.428 3.156 24.46 ;
  LAYER M2 ;
        RECT 0.08 24.428 3.12 24.46 ;
  LAYER M1 ;
        RECT 0.064 24.408 0.096 24.48 ;
  LAYER M2 ;
        RECT 0.044 24.428 0.116 24.46 ;
  LAYER M1 ;
        RECT 3.104 27.348 3.136 27.42 ;
  LAYER M2 ;
        RECT 3.084 27.368 3.156 27.4 ;
  LAYER M2 ;
        RECT 0.08 27.368 3.12 27.4 ;
  LAYER M1 ;
        RECT 0.064 27.348 0.096 27.42 ;
  LAYER M2 ;
        RECT 0.044 27.368 0.116 27.4 ;
  LAYER M1 ;
        RECT 3.104 30.288 3.136 30.36 ;
  LAYER M2 ;
        RECT 3.084 30.308 3.156 30.34 ;
  LAYER M2 ;
        RECT 0.08 30.308 3.12 30.34 ;
  LAYER M1 ;
        RECT 0.064 30.288 0.096 30.36 ;
  LAYER M2 ;
        RECT 0.044 30.308 0.116 30.34 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.588 ;
  LAYER M1 ;
        RECT 0.064 0.588 0.096 30.324 ;
  LAYER M1 ;
        RECT 9.504 0.888 9.536 0.96 ;
  LAYER M2 ;
        RECT 9.484 0.908 9.556 0.94 ;
  LAYER M1 ;
        RECT 9.504 0.756 9.536 0.924 ;
  LAYER M1 ;
        RECT 9.504 0.72 9.536 0.792 ;
  LAYER M2 ;
        RECT 9.484 0.74 9.556 0.772 ;
  LAYER M2 ;
        RECT 9.52 0.74 9.68 0.772 ;
  LAYER M1 ;
        RECT 9.664 0.72 9.696 0.792 ;
  LAYER M2 ;
        RECT 9.644 0.74 9.716 0.772 ;
  LAYER M1 ;
        RECT 9.504 3.828 9.536 3.9 ;
  LAYER M2 ;
        RECT 9.484 3.848 9.556 3.88 ;
  LAYER M1 ;
        RECT 9.504 3.696 9.536 3.864 ;
  LAYER M1 ;
        RECT 9.504 3.66 9.536 3.732 ;
  LAYER M2 ;
        RECT 9.484 3.68 9.556 3.712 ;
  LAYER M2 ;
        RECT 9.52 3.68 9.68 3.712 ;
  LAYER M1 ;
        RECT 9.664 3.66 9.696 3.732 ;
  LAYER M2 ;
        RECT 9.644 3.68 9.716 3.712 ;
  LAYER M1 ;
        RECT 9.504 6.768 9.536 6.84 ;
  LAYER M2 ;
        RECT 9.484 6.788 9.556 6.82 ;
  LAYER M1 ;
        RECT 9.504 6.636 9.536 6.804 ;
  LAYER M1 ;
        RECT 9.504 6.6 9.536 6.672 ;
  LAYER M2 ;
        RECT 9.484 6.62 9.556 6.652 ;
  LAYER M2 ;
        RECT 9.52 6.62 9.68 6.652 ;
  LAYER M1 ;
        RECT 9.664 6.6 9.696 6.672 ;
  LAYER M2 ;
        RECT 9.644 6.62 9.716 6.652 ;
  LAYER M1 ;
        RECT 9.504 9.708 9.536 9.78 ;
  LAYER M2 ;
        RECT 9.484 9.728 9.556 9.76 ;
  LAYER M1 ;
        RECT 9.504 9.576 9.536 9.744 ;
  LAYER M1 ;
        RECT 9.504 9.54 9.536 9.612 ;
  LAYER M2 ;
        RECT 9.484 9.56 9.556 9.592 ;
  LAYER M2 ;
        RECT 9.52 9.56 9.68 9.592 ;
  LAYER M1 ;
        RECT 9.664 9.54 9.696 9.612 ;
  LAYER M2 ;
        RECT 9.644 9.56 9.716 9.592 ;
  LAYER M1 ;
        RECT 9.504 12.648 9.536 12.72 ;
  LAYER M2 ;
        RECT 9.484 12.668 9.556 12.7 ;
  LAYER M1 ;
        RECT 9.504 12.516 9.536 12.684 ;
  LAYER M1 ;
        RECT 9.504 12.48 9.536 12.552 ;
  LAYER M2 ;
        RECT 9.484 12.5 9.556 12.532 ;
  LAYER M2 ;
        RECT 9.52 12.5 9.68 12.532 ;
  LAYER M1 ;
        RECT 9.664 12.48 9.696 12.552 ;
  LAYER M2 ;
        RECT 9.644 12.5 9.716 12.532 ;
  LAYER M1 ;
        RECT 9.504 15.588 9.536 15.66 ;
  LAYER M2 ;
        RECT 9.484 15.608 9.556 15.64 ;
  LAYER M1 ;
        RECT 9.504 15.456 9.536 15.624 ;
  LAYER M1 ;
        RECT 9.504 15.42 9.536 15.492 ;
  LAYER M2 ;
        RECT 9.484 15.44 9.556 15.472 ;
  LAYER M2 ;
        RECT 9.52 15.44 9.68 15.472 ;
  LAYER M1 ;
        RECT 9.664 15.42 9.696 15.492 ;
  LAYER M2 ;
        RECT 9.644 15.44 9.716 15.472 ;
  LAYER M1 ;
        RECT 9.504 18.528 9.536 18.6 ;
  LAYER M2 ;
        RECT 9.484 18.548 9.556 18.58 ;
  LAYER M1 ;
        RECT 9.504 18.396 9.536 18.564 ;
  LAYER M1 ;
        RECT 9.504 18.36 9.536 18.432 ;
  LAYER M2 ;
        RECT 9.484 18.38 9.556 18.412 ;
  LAYER M2 ;
        RECT 9.52 18.38 9.68 18.412 ;
  LAYER M1 ;
        RECT 9.664 18.36 9.696 18.432 ;
  LAYER M2 ;
        RECT 9.644 18.38 9.716 18.412 ;
  LAYER M1 ;
        RECT 9.504 21.468 9.536 21.54 ;
  LAYER M2 ;
        RECT 9.484 21.488 9.556 21.52 ;
  LAYER M1 ;
        RECT 9.504 21.336 9.536 21.504 ;
  LAYER M1 ;
        RECT 9.504 21.3 9.536 21.372 ;
  LAYER M2 ;
        RECT 9.484 21.32 9.556 21.352 ;
  LAYER M2 ;
        RECT 9.52 21.32 9.68 21.352 ;
  LAYER M1 ;
        RECT 9.664 21.3 9.696 21.372 ;
  LAYER M2 ;
        RECT 9.644 21.32 9.716 21.352 ;
  LAYER M1 ;
        RECT 9.504 24.408 9.536 24.48 ;
  LAYER M2 ;
        RECT 9.484 24.428 9.556 24.46 ;
  LAYER M1 ;
        RECT 9.504 24.276 9.536 24.444 ;
  LAYER M1 ;
        RECT 9.504 24.24 9.536 24.312 ;
  LAYER M2 ;
        RECT 9.484 24.26 9.556 24.292 ;
  LAYER M2 ;
        RECT 9.52 24.26 9.68 24.292 ;
  LAYER M1 ;
        RECT 9.664 24.24 9.696 24.312 ;
  LAYER M2 ;
        RECT 9.644 24.26 9.716 24.292 ;
  LAYER M1 ;
        RECT 9.504 27.348 9.536 27.42 ;
  LAYER M2 ;
        RECT 9.484 27.368 9.556 27.4 ;
  LAYER M1 ;
        RECT 9.504 27.216 9.536 27.384 ;
  LAYER M1 ;
        RECT 9.504 27.18 9.536 27.252 ;
  LAYER M2 ;
        RECT 9.484 27.2 9.556 27.232 ;
  LAYER M2 ;
        RECT 9.52 27.2 9.68 27.232 ;
  LAYER M1 ;
        RECT 9.664 27.18 9.696 27.252 ;
  LAYER M2 ;
        RECT 9.644 27.2 9.716 27.232 ;
  LAYER M1 ;
        RECT 9.504 30.288 9.536 30.36 ;
  LAYER M2 ;
        RECT 9.484 30.308 9.556 30.34 ;
  LAYER M1 ;
        RECT 9.504 30.156 9.536 30.324 ;
  LAYER M1 ;
        RECT 9.504 30.12 9.536 30.192 ;
  LAYER M2 ;
        RECT 9.484 30.14 9.556 30.172 ;
  LAYER M2 ;
        RECT 9.52 30.14 9.68 30.172 ;
  LAYER M1 ;
        RECT 9.664 30.12 9.696 30.192 ;
  LAYER M2 ;
        RECT 9.644 30.14 9.716 30.172 ;
  LAYER M1 ;
        RECT 9.664 0.048 9.696 0.12 ;
  LAYER M2 ;
        RECT 9.644 0.068 9.716 0.1 ;
  LAYER M1 ;
        RECT 9.664 0.084 9.696 0.588 ;
  LAYER M1 ;
        RECT 9.664 0.588 9.696 30.156 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.68 0.1 ;
  LAYER M1 ;
        RECT 6.304 0.888 6.336 0.96 ;
  LAYER M2 ;
        RECT 6.284 0.908 6.356 0.94 ;
  LAYER M2 ;
        RECT 3.12 0.908 6.32 0.94 ;
  LAYER M1 ;
        RECT 3.104 0.888 3.136 0.96 ;
  LAYER M2 ;
        RECT 3.084 0.908 3.156 0.94 ;
  LAYER M1 ;
        RECT 6.304 30.288 6.336 30.36 ;
  LAYER M2 ;
        RECT 6.284 30.308 6.356 30.34 ;
  LAYER M2 ;
        RECT 3.12 30.308 6.32 30.34 ;
  LAYER M1 ;
        RECT 3.104 30.288 3.136 30.36 ;
  LAYER M2 ;
        RECT 3.084 30.308 3.156 30.34 ;
  LAYER M1 ;
        RECT 3.904 18.024 3.936 18.096 ;
  LAYER M2 ;
        RECT 3.884 18.044 3.956 18.076 ;
  LAYER M2 ;
        RECT 3.6 18.044 3.92 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M1 ;
        RECT 3.904 6.264 3.936 6.336 ;
  LAYER M2 ;
        RECT 3.884 6.284 3.956 6.316 ;
  LAYER M2 ;
        RECT 3.6 6.284 3.92 6.316 ;
  LAYER M1 ;
        RECT 3.584 6.264 3.616 6.336 ;
  LAYER M2 ;
        RECT 3.564 6.284 3.636 6.316 ;
  LAYER M1 ;
        RECT 3.904 29.784 3.936 29.856 ;
  LAYER M2 ;
        RECT 3.884 29.804 3.956 29.836 ;
  LAYER M2 ;
        RECT 3.6 29.804 3.92 29.836 ;
  LAYER M1 ;
        RECT 3.584 29.784 3.616 29.856 ;
  LAYER M2 ;
        RECT 3.564 29.804 3.636 29.836 ;
  LAYER M1 ;
        RECT 3.584 33.228 3.616 33.3 ;
  LAYER M2 ;
        RECT 3.564 33.248 3.636 33.28 ;
  LAYER M1 ;
        RECT 3.584 33.096 3.616 33.264 ;
  LAYER M1 ;
        RECT 3.584 6.3 3.616 33.096 ;
  LAYER M1 ;
        RECT 3.904 18.024 3.936 18.096 ;
  LAYER M2 ;
        RECT 3.884 18.044 3.956 18.076 ;
  LAYER M1 ;
        RECT 3.904 18.06 3.936 18.228 ;
  LAYER M1 ;
        RECT 3.904 18.192 3.936 18.264 ;
  LAYER M2 ;
        RECT 3.884 18.212 3.956 18.244 ;
  LAYER M2 ;
        RECT 3.92 18.212 6.8 18.244 ;
  LAYER M1 ;
        RECT 6.784 18.192 6.816 18.264 ;
  LAYER M2 ;
        RECT 6.764 18.212 6.836 18.244 ;
  LAYER M1 ;
        RECT 3.904 6.264 3.936 6.336 ;
  LAYER M2 ;
        RECT 3.884 6.284 3.956 6.316 ;
  LAYER M1 ;
        RECT 3.904 6.3 3.936 6.468 ;
  LAYER M1 ;
        RECT 3.904 6.432 3.936 6.504 ;
  LAYER M2 ;
        RECT 3.884 6.452 3.956 6.484 ;
  LAYER M2 ;
        RECT 3.92 6.452 6.8 6.484 ;
  LAYER M1 ;
        RECT 6.784 6.432 6.816 6.504 ;
  LAYER M2 ;
        RECT 6.764 6.452 6.836 6.484 ;
  LAYER M1 ;
        RECT 3.904 29.784 3.936 29.856 ;
  LAYER M2 ;
        RECT 3.884 29.804 3.956 29.836 ;
  LAYER M1 ;
        RECT 3.904 29.82 3.936 29.988 ;
  LAYER M1 ;
        RECT 3.904 29.952 3.936 30.024 ;
  LAYER M2 ;
        RECT 3.884 29.972 3.956 30.004 ;
  LAYER M2 ;
        RECT 3.92 29.972 6.8 30.004 ;
  LAYER M1 ;
        RECT 6.784 29.952 6.816 30.024 ;
  LAYER M2 ;
        RECT 6.764 29.972 6.836 30.004 ;
  LAYER M1 ;
        RECT 6.784 33.228 6.816 33.3 ;
  LAYER M2 ;
        RECT 6.764 33.248 6.836 33.28 ;
  LAYER M1 ;
        RECT 6.784 33.096 6.816 33.264 ;
  LAYER M1 ;
        RECT 6.784 6.468 6.816 33.096 ;
  LAYER M2 ;
        RECT 3.6 33.248 6.8 33.28 ;
  LAYER M1 ;
        RECT 3.904 15.084 3.936 15.156 ;
  LAYER M2 ;
        RECT 3.884 15.104 3.956 15.136 ;
  LAYER M2 ;
        RECT 3.76 15.104 3.92 15.136 ;
  LAYER M1 ;
        RECT 3.744 15.084 3.776 15.156 ;
  LAYER M2 ;
        RECT 3.724 15.104 3.796 15.136 ;
  LAYER M1 ;
        RECT 3.904 20.964 3.936 21.036 ;
  LAYER M2 ;
        RECT 3.884 20.984 3.956 21.016 ;
  LAYER M2 ;
        RECT 3.76 20.984 3.92 21.016 ;
  LAYER M1 ;
        RECT 3.744 20.964 3.776 21.036 ;
  LAYER M2 ;
        RECT 3.724 20.984 3.796 21.016 ;
  LAYER M1 ;
        RECT 3.904 12.144 3.936 12.216 ;
  LAYER M2 ;
        RECT 3.884 12.164 3.956 12.196 ;
  LAYER M2 ;
        RECT 3.76 12.164 3.92 12.196 ;
  LAYER M1 ;
        RECT 3.744 12.144 3.776 12.216 ;
  LAYER M2 ;
        RECT 3.724 12.164 3.796 12.196 ;
  LAYER M1 ;
        RECT 3.904 23.904 3.936 23.976 ;
  LAYER M2 ;
        RECT 3.884 23.924 3.956 23.956 ;
  LAYER M2 ;
        RECT 3.76 23.924 3.92 23.956 ;
  LAYER M1 ;
        RECT 3.744 23.904 3.776 23.976 ;
  LAYER M2 ;
        RECT 3.724 23.924 3.796 23.956 ;
  LAYER M1 ;
        RECT 3.904 9.204 3.936 9.276 ;
  LAYER M2 ;
        RECT 3.884 9.224 3.956 9.256 ;
  LAYER M2 ;
        RECT 3.76 9.224 3.92 9.256 ;
  LAYER M1 ;
        RECT 3.744 9.204 3.776 9.276 ;
  LAYER M2 ;
        RECT 3.724 9.224 3.796 9.256 ;
  LAYER M1 ;
        RECT 3.904 26.844 3.936 26.916 ;
  LAYER M2 ;
        RECT 3.884 26.864 3.956 26.896 ;
  LAYER M2 ;
        RECT 3.76 26.864 3.92 26.896 ;
  LAYER M1 ;
        RECT 3.744 26.844 3.776 26.916 ;
  LAYER M2 ;
        RECT 3.724 26.864 3.796 26.896 ;
  LAYER M1 ;
        RECT 3.744 33.396 3.776 33.468 ;
  LAYER M2 ;
        RECT 3.724 33.416 3.796 33.448 ;
  LAYER M1 ;
        RECT 3.744 33.096 3.776 33.432 ;
  LAYER M1 ;
        RECT 3.744 9.24 3.776 33.096 ;
  LAYER M1 ;
        RECT 3.904 15.084 3.936 15.156 ;
  LAYER M2 ;
        RECT 3.884 15.104 3.956 15.136 ;
  LAYER M1 ;
        RECT 3.904 15.12 3.936 15.288 ;
  LAYER M1 ;
        RECT 3.904 15.252 3.936 15.324 ;
  LAYER M2 ;
        RECT 3.884 15.272 3.956 15.304 ;
  LAYER M2 ;
        RECT 3.92 15.272 6.96 15.304 ;
  LAYER M1 ;
        RECT 6.944 15.252 6.976 15.324 ;
  LAYER M2 ;
        RECT 6.924 15.272 6.996 15.304 ;
  LAYER M1 ;
        RECT 3.904 20.964 3.936 21.036 ;
  LAYER M2 ;
        RECT 3.884 20.984 3.956 21.016 ;
  LAYER M1 ;
        RECT 3.904 21 3.936 21.168 ;
  LAYER M1 ;
        RECT 3.904 21.132 3.936 21.204 ;
  LAYER M2 ;
        RECT 3.884 21.152 3.956 21.184 ;
  LAYER M2 ;
        RECT 3.92 21.152 6.96 21.184 ;
  LAYER M1 ;
        RECT 6.944 21.132 6.976 21.204 ;
  LAYER M2 ;
        RECT 6.924 21.152 6.996 21.184 ;
  LAYER M1 ;
        RECT 3.904 12.144 3.936 12.216 ;
  LAYER M2 ;
        RECT 3.884 12.164 3.956 12.196 ;
  LAYER M1 ;
        RECT 3.904 12.18 3.936 12.348 ;
  LAYER M1 ;
        RECT 3.904 12.312 3.936 12.384 ;
  LAYER M2 ;
        RECT 3.884 12.332 3.956 12.364 ;
  LAYER M2 ;
        RECT 3.92 12.332 6.96 12.364 ;
  LAYER M1 ;
        RECT 6.944 12.312 6.976 12.384 ;
  LAYER M2 ;
        RECT 6.924 12.332 6.996 12.364 ;
  LAYER M1 ;
        RECT 3.904 23.904 3.936 23.976 ;
  LAYER M2 ;
        RECT 3.884 23.924 3.956 23.956 ;
  LAYER M1 ;
        RECT 3.904 23.94 3.936 24.108 ;
  LAYER M1 ;
        RECT 3.904 24.072 3.936 24.144 ;
  LAYER M2 ;
        RECT 3.884 24.092 3.956 24.124 ;
  LAYER M2 ;
        RECT 3.92 24.092 6.96 24.124 ;
  LAYER M1 ;
        RECT 6.944 24.072 6.976 24.144 ;
  LAYER M2 ;
        RECT 6.924 24.092 6.996 24.124 ;
  LAYER M1 ;
        RECT 3.904 9.204 3.936 9.276 ;
  LAYER M2 ;
        RECT 3.884 9.224 3.956 9.256 ;
  LAYER M1 ;
        RECT 3.904 9.24 3.936 9.408 ;
  LAYER M1 ;
        RECT 3.904 9.372 3.936 9.444 ;
  LAYER M2 ;
        RECT 3.884 9.392 3.956 9.424 ;
  LAYER M2 ;
        RECT 3.92 9.392 6.96 9.424 ;
  LAYER M1 ;
        RECT 6.944 9.372 6.976 9.444 ;
  LAYER M2 ;
        RECT 6.924 9.392 6.996 9.424 ;
  LAYER M1 ;
        RECT 3.904 26.844 3.936 26.916 ;
  LAYER M2 ;
        RECT 3.884 26.864 3.956 26.896 ;
  LAYER M1 ;
        RECT 3.904 26.88 3.936 27.048 ;
  LAYER M1 ;
        RECT 3.904 27.012 3.936 27.084 ;
  LAYER M2 ;
        RECT 3.884 27.032 3.956 27.064 ;
  LAYER M2 ;
        RECT 3.92 27.032 6.96 27.064 ;
  LAYER M1 ;
        RECT 6.944 27.012 6.976 27.084 ;
  LAYER M2 ;
        RECT 6.924 27.032 6.996 27.064 ;
  LAYER M1 ;
        RECT 6.944 33.396 6.976 33.468 ;
  LAYER M2 ;
        RECT 6.924 33.416 6.996 33.448 ;
  LAYER M1 ;
        RECT 6.944 33.096 6.976 33.432 ;
  LAYER M1 ;
        RECT 6.944 9.408 6.976 33.096 ;
  LAYER M2 ;
        RECT 3.76 33.416 6.96 33.448 ;
  LAYER M1 ;
        RECT 0.704 3.324 0.736 3.396 ;
  LAYER M2 ;
        RECT 0.684 3.344 0.756 3.376 ;
  LAYER M2 ;
        RECT 0.24 3.344 0.72 3.376 ;
  LAYER M1 ;
        RECT 0.224 3.324 0.256 3.396 ;
  LAYER M2 ;
        RECT 0.204 3.344 0.276 3.376 ;
  LAYER M1 ;
        RECT 0.704 6.264 0.736 6.336 ;
  LAYER M2 ;
        RECT 0.684 6.284 0.756 6.316 ;
  LAYER M2 ;
        RECT 0.24 6.284 0.72 6.316 ;
  LAYER M1 ;
        RECT 0.224 6.264 0.256 6.336 ;
  LAYER M2 ;
        RECT 0.204 6.284 0.276 6.316 ;
  LAYER M1 ;
        RECT 0.704 9.204 0.736 9.276 ;
  LAYER M2 ;
        RECT 0.684 9.224 0.756 9.256 ;
  LAYER M2 ;
        RECT 0.24 9.224 0.72 9.256 ;
  LAYER M1 ;
        RECT 0.224 9.204 0.256 9.276 ;
  LAYER M2 ;
        RECT 0.204 9.224 0.276 9.256 ;
  LAYER M1 ;
        RECT 0.704 12.144 0.736 12.216 ;
  LAYER M2 ;
        RECT 0.684 12.164 0.756 12.196 ;
  LAYER M2 ;
        RECT 0.24 12.164 0.72 12.196 ;
  LAYER M1 ;
        RECT 0.224 12.144 0.256 12.216 ;
  LAYER M2 ;
        RECT 0.204 12.164 0.276 12.196 ;
  LAYER M1 ;
        RECT 0.704 15.084 0.736 15.156 ;
  LAYER M2 ;
        RECT 0.684 15.104 0.756 15.136 ;
  LAYER M2 ;
        RECT 0.24 15.104 0.72 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.084 0.256 15.156 ;
  LAYER M2 ;
        RECT 0.204 15.104 0.276 15.136 ;
  LAYER M1 ;
        RECT 0.704 18.024 0.736 18.096 ;
  LAYER M2 ;
        RECT 0.684 18.044 0.756 18.076 ;
  LAYER M2 ;
        RECT 0.24 18.044 0.72 18.076 ;
  LAYER M1 ;
        RECT 0.224 18.024 0.256 18.096 ;
  LAYER M2 ;
        RECT 0.204 18.044 0.276 18.076 ;
  LAYER M1 ;
        RECT 0.704 20.964 0.736 21.036 ;
  LAYER M2 ;
        RECT 0.684 20.984 0.756 21.016 ;
  LAYER M2 ;
        RECT 0.24 20.984 0.72 21.016 ;
  LAYER M1 ;
        RECT 0.224 20.964 0.256 21.036 ;
  LAYER M2 ;
        RECT 0.204 20.984 0.276 21.016 ;
  LAYER M1 ;
        RECT 0.704 23.904 0.736 23.976 ;
  LAYER M2 ;
        RECT 0.684 23.924 0.756 23.956 ;
  LAYER M2 ;
        RECT 0.24 23.924 0.72 23.956 ;
  LAYER M1 ;
        RECT 0.224 23.904 0.256 23.976 ;
  LAYER M2 ;
        RECT 0.204 23.924 0.276 23.956 ;
  LAYER M1 ;
        RECT 0.704 26.844 0.736 26.916 ;
  LAYER M2 ;
        RECT 0.684 26.864 0.756 26.896 ;
  LAYER M2 ;
        RECT 0.24 26.864 0.72 26.896 ;
  LAYER M1 ;
        RECT 0.224 26.844 0.256 26.916 ;
  LAYER M2 ;
        RECT 0.204 26.864 0.276 26.896 ;
  LAYER M1 ;
        RECT 0.704 29.784 0.736 29.856 ;
  LAYER M2 ;
        RECT 0.684 29.804 0.756 29.836 ;
  LAYER M2 ;
        RECT 0.24 29.804 0.72 29.836 ;
  LAYER M1 ;
        RECT 0.224 29.784 0.256 29.856 ;
  LAYER M2 ;
        RECT 0.204 29.804 0.276 29.836 ;
  LAYER M1 ;
        RECT 0.704 32.724 0.736 32.796 ;
  LAYER M2 ;
        RECT 0.684 32.744 0.756 32.776 ;
  LAYER M2 ;
        RECT 0.24 32.744 0.72 32.776 ;
  LAYER M1 ;
        RECT 0.224 32.724 0.256 32.796 ;
  LAYER M2 ;
        RECT 0.204 32.744 0.276 32.776 ;
  LAYER M1 ;
        RECT 0.224 33.564 0.256 33.636 ;
  LAYER M2 ;
        RECT 0.204 33.584 0.276 33.616 ;
  LAYER M1 ;
        RECT 0.224 33.096 0.256 33.6 ;
  LAYER M1 ;
        RECT 0.224 3.36 0.256 33.096 ;
  LAYER M1 ;
        RECT 7.104 3.324 7.136 3.396 ;
  LAYER M2 ;
        RECT 7.084 3.344 7.156 3.376 ;
  LAYER M1 ;
        RECT 7.104 3.36 7.136 3.528 ;
  LAYER M1 ;
        RECT 7.104 3.492 7.136 3.564 ;
  LAYER M2 ;
        RECT 7.084 3.512 7.156 3.544 ;
  LAYER M2 ;
        RECT 7.12 3.512 9.84 3.544 ;
  LAYER M1 ;
        RECT 9.824 3.492 9.856 3.564 ;
  LAYER M2 ;
        RECT 9.804 3.512 9.876 3.544 ;
  LAYER M1 ;
        RECT 7.104 6.264 7.136 6.336 ;
  LAYER M2 ;
        RECT 7.084 6.284 7.156 6.316 ;
  LAYER M1 ;
        RECT 7.104 6.3 7.136 6.468 ;
  LAYER M1 ;
        RECT 7.104 6.432 7.136 6.504 ;
  LAYER M2 ;
        RECT 7.084 6.452 7.156 6.484 ;
  LAYER M2 ;
        RECT 7.12 6.452 9.84 6.484 ;
  LAYER M1 ;
        RECT 9.824 6.432 9.856 6.504 ;
  LAYER M2 ;
        RECT 9.804 6.452 9.876 6.484 ;
  LAYER M1 ;
        RECT 7.104 9.204 7.136 9.276 ;
  LAYER M2 ;
        RECT 7.084 9.224 7.156 9.256 ;
  LAYER M1 ;
        RECT 7.104 9.24 7.136 9.408 ;
  LAYER M1 ;
        RECT 7.104 9.372 7.136 9.444 ;
  LAYER M2 ;
        RECT 7.084 9.392 7.156 9.424 ;
  LAYER M2 ;
        RECT 7.12 9.392 9.84 9.424 ;
  LAYER M1 ;
        RECT 9.824 9.372 9.856 9.444 ;
  LAYER M2 ;
        RECT 9.804 9.392 9.876 9.424 ;
  LAYER M1 ;
        RECT 7.104 12.144 7.136 12.216 ;
  LAYER M2 ;
        RECT 7.084 12.164 7.156 12.196 ;
  LAYER M1 ;
        RECT 7.104 12.18 7.136 12.348 ;
  LAYER M1 ;
        RECT 7.104 12.312 7.136 12.384 ;
  LAYER M2 ;
        RECT 7.084 12.332 7.156 12.364 ;
  LAYER M2 ;
        RECT 7.12 12.332 9.84 12.364 ;
  LAYER M1 ;
        RECT 9.824 12.312 9.856 12.384 ;
  LAYER M2 ;
        RECT 9.804 12.332 9.876 12.364 ;
  LAYER M1 ;
        RECT 7.104 15.084 7.136 15.156 ;
  LAYER M2 ;
        RECT 7.084 15.104 7.156 15.136 ;
  LAYER M1 ;
        RECT 7.104 15.12 7.136 15.288 ;
  LAYER M1 ;
        RECT 7.104 15.252 7.136 15.324 ;
  LAYER M2 ;
        RECT 7.084 15.272 7.156 15.304 ;
  LAYER M2 ;
        RECT 7.12 15.272 9.84 15.304 ;
  LAYER M1 ;
        RECT 9.824 15.252 9.856 15.324 ;
  LAYER M2 ;
        RECT 9.804 15.272 9.876 15.304 ;
  LAYER M1 ;
        RECT 7.104 18.024 7.136 18.096 ;
  LAYER M2 ;
        RECT 7.084 18.044 7.156 18.076 ;
  LAYER M1 ;
        RECT 7.104 18.06 7.136 18.228 ;
  LAYER M1 ;
        RECT 7.104 18.192 7.136 18.264 ;
  LAYER M2 ;
        RECT 7.084 18.212 7.156 18.244 ;
  LAYER M2 ;
        RECT 7.12 18.212 9.84 18.244 ;
  LAYER M1 ;
        RECT 9.824 18.192 9.856 18.264 ;
  LAYER M2 ;
        RECT 9.804 18.212 9.876 18.244 ;
  LAYER M1 ;
        RECT 7.104 20.964 7.136 21.036 ;
  LAYER M2 ;
        RECT 7.084 20.984 7.156 21.016 ;
  LAYER M1 ;
        RECT 7.104 21 7.136 21.168 ;
  LAYER M1 ;
        RECT 7.104 21.132 7.136 21.204 ;
  LAYER M2 ;
        RECT 7.084 21.152 7.156 21.184 ;
  LAYER M2 ;
        RECT 7.12 21.152 9.84 21.184 ;
  LAYER M1 ;
        RECT 9.824 21.132 9.856 21.204 ;
  LAYER M2 ;
        RECT 9.804 21.152 9.876 21.184 ;
  LAYER M1 ;
        RECT 7.104 23.904 7.136 23.976 ;
  LAYER M2 ;
        RECT 7.084 23.924 7.156 23.956 ;
  LAYER M1 ;
        RECT 7.104 23.94 7.136 24.108 ;
  LAYER M1 ;
        RECT 7.104 24.072 7.136 24.144 ;
  LAYER M2 ;
        RECT 7.084 24.092 7.156 24.124 ;
  LAYER M2 ;
        RECT 7.12 24.092 9.84 24.124 ;
  LAYER M1 ;
        RECT 9.824 24.072 9.856 24.144 ;
  LAYER M2 ;
        RECT 9.804 24.092 9.876 24.124 ;
  LAYER M1 ;
        RECT 7.104 26.844 7.136 26.916 ;
  LAYER M2 ;
        RECT 7.084 26.864 7.156 26.896 ;
  LAYER M1 ;
        RECT 7.104 26.88 7.136 27.048 ;
  LAYER M1 ;
        RECT 7.104 27.012 7.136 27.084 ;
  LAYER M2 ;
        RECT 7.084 27.032 7.156 27.064 ;
  LAYER M2 ;
        RECT 7.12 27.032 9.84 27.064 ;
  LAYER M1 ;
        RECT 9.824 27.012 9.856 27.084 ;
  LAYER M2 ;
        RECT 9.804 27.032 9.876 27.064 ;
  LAYER M1 ;
        RECT 7.104 29.784 7.136 29.856 ;
  LAYER M2 ;
        RECT 7.084 29.804 7.156 29.836 ;
  LAYER M1 ;
        RECT 7.104 29.82 7.136 29.988 ;
  LAYER M1 ;
        RECT 7.104 29.952 7.136 30.024 ;
  LAYER M2 ;
        RECT 7.084 29.972 7.156 30.004 ;
  LAYER M2 ;
        RECT 7.12 29.972 9.84 30.004 ;
  LAYER M1 ;
        RECT 9.824 29.952 9.856 30.024 ;
  LAYER M2 ;
        RECT 9.804 29.972 9.876 30.004 ;
  LAYER M1 ;
        RECT 7.104 32.724 7.136 32.796 ;
  LAYER M2 ;
        RECT 7.084 32.744 7.156 32.776 ;
  LAYER M1 ;
        RECT 7.104 32.76 7.136 32.928 ;
  LAYER M1 ;
        RECT 7.104 32.892 7.136 32.964 ;
  LAYER M2 ;
        RECT 7.084 32.912 7.156 32.944 ;
  LAYER M2 ;
        RECT 7.12 32.912 9.84 32.944 ;
  LAYER M1 ;
        RECT 9.824 32.892 9.856 32.964 ;
  LAYER M2 ;
        RECT 9.804 32.912 9.876 32.944 ;
  LAYER M1 ;
        RECT 9.824 33.564 9.856 33.636 ;
  LAYER M2 ;
        RECT 9.804 33.584 9.876 33.616 ;
  LAYER M1 ;
        RECT 9.824 33.096 9.856 33.6 ;
  LAYER M1 ;
        RECT 9.824 3.528 9.856 33.096 ;
  LAYER M2 ;
        RECT 0.24 33.584 9.84 33.616 ;
  LAYER M1 ;
        RECT 3.904 3.324 3.936 3.396 ;
  LAYER M2 ;
        RECT 3.884 3.344 3.956 3.376 ;
  LAYER M2 ;
        RECT 0.72 3.344 3.92 3.376 ;
  LAYER M1 ;
        RECT 0.704 3.324 0.736 3.396 ;
  LAYER M2 ;
        RECT 0.684 3.344 0.756 3.376 ;
  LAYER M1 ;
        RECT 3.904 32.724 3.936 32.796 ;
  LAYER M2 ;
        RECT 3.884 32.744 3.956 32.776 ;
  LAYER M2 ;
        RECT 0.72 32.744 3.92 32.776 ;
  LAYER M1 ;
        RECT 0.704 32.724 0.736 32.796 ;
  LAYER M2 ;
        RECT 0.684 32.744 0.756 32.776 ;
  LAYER M1 ;
        RECT 0.72 0.924 3.12 3.36 ;
  LAYER M2 ;
        RECT 0.72 0.924 3.12 3.36 ;
  LAYER M3 ;
        RECT 0.72 0.924 3.12 3.36 ;
  LAYER M1 ;
        RECT 0.72 3.864 3.12 6.3 ;
  LAYER M2 ;
        RECT 0.72 3.864 3.12 6.3 ;
  LAYER M3 ;
        RECT 0.72 3.864 3.12 6.3 ;
  LAYER M1 ;
        RECT 0.72 6.804 3.12 9.24 ;
  LAYER M2 ;
        RECT 0.72 6.804 3.12 9.24 ;
  LAYER M3 ;
        RECT 0.72 6.804 3.12 9.24 ;
  LAYER M1 ;
        RECT 0.72 9.744 3.12 12.18 ;
  LAYER M2 ;
        RECT 0.72 9.744 3.12 12.18 ;
  LAYER M3 ;
        RECT 0.72 9.744 3.12 12.18 ;
  LAYER M1 ;
        RECT 0.72 12.684 3.12 15.12 ;
  LAYER M2 ;
        RECT 0.72 12.684 3.12 15.12 ;
  LAYER M3 ;
        RECT 0.72 12.684 3.12 15.12 ;
  LAYER M1 ;
        RECT 0.72 15.624 3.12 18.06 ;
  LAYER M2 ;
        RECT 0.72 15.624 3.12 18.06 ;
  LAYER M3 ;
        RECT 0.72 15.624 3.12 18.06 ;
  LAYER M1 ;
        RECT 0.72 18.564 3.12 21 ;
  LAYER M2 ;
        RECT 0.72 18.564 3.12 21 ;
  LAYER M3 ;
        RECT 0.72 18.564 3.12 21 ;
  LAYER M1 ;
        RECT 0.72 21.504 3.12 23.94 ;
  LAYER M2 ;
        RECT 0.72 21.504 3.12 23.94 ;
  LAYER M3 ;
        RECT 0.72 21.504 3.12 23.94 ;
  LAYER M1 ;
        RECT 0.72 24.444 3.12 26.88 ;
  LAYER M2 ;
        RECT 0.72 24.444 3.12 26.88 ;
  LAYER M3 ;
        RECT 0.72 24.444 3.12 26.88 ;
  LAYER M1 ;
        RECT 0.72 27.384 3.12 29.82 ;
  LAYER M2 ;
        RECT 0.72 27.384 3.12 29.82 ;
  LAYER M3 ;
        RECT 0.72 27.384 3.12 29.82 ;
  LAYER M1 ;
        RECT 0.72 30.324 3.12 32.76 ;
  LAYER M2 ;
        RECT 0.72 30.324 3.12 32.76 ;
  LAYER M3 ;
        RECT 0.72 30.324 3.12 32.76 ;
  LAYER M1 ;
        RECT 3.92 0.924 6.32 3.36 ;
  LAYER M2 ;
        RECT 3.92 0.924 6.32 3.36 ;
  LAYER M3 ;
        RECT 3.92 0.924 6.32 3.36 ;
  LAYER M1 ;
        RECT 3.92 3.864 6.32 6.3 ;
  LAYER M2 ;
        RECT 3.92 3.864 6.32 6.3 ;
  LAYER M3 ;
        RECT 3.92 3.864 6.32 6.3 ;
  LAYER M1 ;
        RECT 3.92 6.804 6.32 9.24 ;
  LAYER M2 ;
        RECT 3.92 6.804 6.32 9.24 ;
  LAYER M3 ;
        RECT 3.92 6.804 6.32 9.24 ;
  LAYER M1 ;
        RECT 3.92 9.744 6.32 12.18 ;
  LAYER M2 ;
        RECT 3.92 9.744 6.32 12.18 ;
  LAYER M3 ;
        RECT 3.92 9.744 6.32 12.18 ;
  LAYER M1 ;
        RECT 3.92 12.684 6.32 15.12 ;
  LAYER M2 ;
        RECT 3.92 12.684 6.32 15.12 ;
  LAYER M3 ;
        RECT 3.92 12.684 6.32 15.12 ;
  LAYER M1 ;
        RECT 3.92 15.624 6.32 18.06 ;
  LAYER M2 ;
        RECT 3.92 15.624 6.32 18.06 ;
  LAYER M3 ;
        RECT 3.92 15.624 6.32 18.06 ;
  LAYER M1 ;
        RECT 3.92 18.564 6.32 21 ;
  LAYER M2 ;
        RECT 3.92 18.564 6.32 21 ;
  LAYER M3 ;
        RECT 3.92 18.564 6.32 21 ;
  LAYER M1 ;
        RECT 3.92 21.504 6.32 23.94 ;
  LAYER M2 ;
        RECT 3.92 21.504 6.32 23.94 ;
  LAYER M3 ;
        RECT 3.92 21.504 6.32 23.94 ;
  LAYER M1 ;
        RECT 3.92 24.444 6.32 26.88 ;
  LAYER M2 ;
        RECT 3.92 24.444 6.32 26.88 ;
  LAYER M3 ;
        RECT 3.92 24.444 6.32 26.88 ;
  LAYER M1 ;
        RECT 3.92 27.384 6.32 29.82 ;
  LAYER M2 ;
        RECT 3.92 27.384 6.32 29.82 ;
  LAYER M3 ;
        RECT 3.92 27.384 6.32 29.82 ;
  LAYER M1 ;
        RECT 3.92 30.324 6.32 32.76 ;
  LAYER M2 ;
        RECT 3.92 30.324 6.32 32.76 ;
  LAYER M3 ;
        RECT 3.92 30.324 6.32 32.76 ;
  LAYER M1 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M2 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M3 ;
        RECT 7.12 0.924 9.52 3.36 ;
  LAYER M1 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M2 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M3 ;
        RECT 7.12 3.864 9.52 6.3 ;
  LAYER M1 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M2 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M3 ;
        RECT 7.12 6.804 9.52 9.24 ;
  LAYER M1 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M2 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M3 ;
        RECT 7.12 9.744 9.52 12.18 ;
  LAYER M1 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M2 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M3 ;
        RECT 7.12 12.684 9.52 15.12 ;
  LAYER M1 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M2 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M3 ;
        RECT 7.12 15.624 9.52 18.06 ;
  LAYER M1 ;
        RECT 7.12 18.564 9.52 21 ;
  LAYER M2 ;
        RECT 7.12 18.564 9.52 21 ;
  LAYER M3 ;
        RECT 7.12 18.564 9.52 21 ;
  LAYER M1 ;
        RECT 7.12 21.504 9.52 23.94 ;
  LAYER M2 ;
        RECT 7.12 21.504 9.52 23.94 ;
  LAYER M3 ;
        RECT 7.12 21.504 9.52 23.94 ;
  LAYER M1 ;
        RECT 7.12 24.444 9.52 26.88 ;
  LAYER M2 ;
        RECT 7.12 24.444 9.52 26.88 ;
  LAYER M3 ;
        RECT 7.12 24.444 9.52 26.88 ;
  LAYER M1 ;
        RECT 7.12 27.384 9.52 29.82 ;
  LAYER M2 ;
        RECT 7.12 27.384 9.52 29.82 ;
  LAYER M3 ;
        RECT 7.12 27.384 9.52 29.82 ;
  LAYER M1 ;
        RECT 7.12 30.324 9.52 32.76 ;
  LAYER M2 ;
        RECT 7.12 30.324 9.52 32.76 ;
  LAYER M3 ;
        RECT 7.12 30.324 9.52 32.76 ;
  END 
END Cap_30fF_Cap_60fF
