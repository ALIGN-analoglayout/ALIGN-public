MACRO switched_capacitor_combination
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_combination 0 0 ;
  SIZE 15.52 BY 29.904 ;
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.46 0.384 10.5 0.708 ;
      LAYER M3 ;
        RECT 10.22 0.384 10.26 0.708 ;
      LAYER M2 ;
        RECT 9.564 0.488 9.796 0.52 ;
      LAYER M2 ;
        RECT 7.724 0.488 7.956 0.52 ;
      LAYER M3 ;
        RECT 10.22 0.252 10.26 0.504 ;
      LAYER M2 ;
        RECT 9.76 0.236 10.24 0.268 ;
      LAYER M3 ;
        RECT 9.74 0.252 9.78 0.504 ;
      LAYER M2 ;
        RECT 9.66 0.488 9.86 0.52 ;
      LAYER M2 ;
        RECT 7.92 0.488 9.6 0.52 ;
    END
  END phi2
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.62 0.552 10.66 0.876 ;
      LAYER M3 ;
        RECT 10.38 0.552 10.42 0.876 ;
      LAYER M2 ;
        RECT 9.644 0.656 9.876 0.688 ;
      LAYER M2 ;
        RECT 7.644 0.656 7.876 0.688 ;
      LAYER M3 ;
        RECT 10.38 0.42 10.42 0.672 ;
      LAYER M4 ;
        RECT 10.08 0.4 10.4 0.44 ;
      LAYER M3 ;
        RECT 10.06 0.42 10.1 0.672 ;
      LAYER M2 ;
        RECT 9.84 0.656 10.08 0.688 ;
      LAYER M2 ;
        RECT 7.76 0.656 9.68 0.688 ;
    END
  END agnd
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.38 17.436 0.42 17.76 ;
      LAYER M3 ;
        RECT 0.14 17.436 0.18 17.76 ;
      LAYER M2 ;
        RECT 9.084 0.572 9.316 0.604 ;
      LAYER M2 ;
        RECT 8.204 0.572 8.436 0.604 ;
      LAYER M3 ;
        RECT 0.38 10.416 0.42 17.472 ;
      LAYER M2 ;
        RECT 0.4 10.4 6.64 10.432 ;
      LAYER M3 ;
        RECT 6.62 8.4 6.66 10.416 ;
      LAYER M4 ;
        RECT 6.64 8.38 8.208 8.42 ;
      LAYER M5 ;
        RECT 8.176 0.588 8.24 8.4 ;
      LAYER M4 ;
        RECT 8.208 0.568 8.64 0.608 ;
      LAYER M3 ;
        RECT 8.62 0.483 8.66 0.693 ;
      LAYER M2 ;
        RECT 8.4 0.572 8.64 0.604 ;
      LAYER M2 ;
        RECT 8.64 0.572 9.12 0.604 ;
    END
  END phi1
  PIN Vin
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.54 17.604 0.58 17.928 ;
      LAYER M3 ;
        RECT 0.3 17.604 0.34 17.928 ;
    END
  END Vin
  PIN Vin_ota
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.164 0.74 9.396 0.772 ;
      LAYER M1 ;
        RECT 3.664 16.764 3.696 16.836 ;
      LAYER M2 ;
        RECT 3.644 16.784 3.716 16.816 ;
      LAYER M1 ;
        RECT 12.304 16.764 12.336 16.836 ;
      LAYER M2 ;
        RECT 12.284 16.784 12.356 16.816 ;
      LAYER M2 ;
        RECT 3.68 16.784 12.32 16.816 ;
      LAYER M2 ;
        RECT 8.96 0.74 9.2 0.772 ;
      LAYER M3 ;
        RECT 8.94 0.756 8.98 1.764 ;
      LAYER M4 ;
        RECT 8.64 1.744 8.96 1.784 ;
      LAYER M5 ;
        RECT 8.608 1.764 8.672 16.548 ;
      LAYER M4 ;
        RECT 8.57 16.528 8.71 16.568 ;
      LAYER M3 ;
        RECT 8.62 16.548 8.66 16.8 ;
      LAYER M2 ;
        RECT 8.54 16.784 8.74 16.816 ;
    END
  END Vin_ota
  PIN Voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.124 0.74 8.356 0.772 ;
      LAYER M1 ;
        RECT 3.824 1.224 3.856 1.296 ;
      LAYER M2 ;
        RECT 3.804 1.244 3.876 1.276 ;
      LAYER M1 ;
        RECT 12.464 1.224 12.496 1.296 ;
      LAYER M2 ;
        RECT 12.444 1.244 12.516 1.276 ;
      LAYER M2 ;
        RECT 3.84 1.244 12.48 1.276 ;
      LAYER M2 ;
        RECT 8.22 0.74 8.42 0.772 ;
      LAYER M3 ;
        RECT 8.3 0.756 8.34 1.26 ;
      LAYER M2 ;
        RECT 8.22 1.244 8.42 1.276 ;
    END
  END Voutn
  OBS 
  LAYER M1 ;
        RECT 9.344 29.616 9.376 29.688 ;
  LAYER M2 ;
        RECT 9.324 29.636 9.396 29.668 ;
  LAYER M1 ;
        RECT 6.464 29.616 6.496 29.688 ;
  LAYER M2 ;
        RECT 6.444 29.636 6.516 29.668 ;
  LAYER M2 ;
        RECT 6.48 29.636 9.36 29.668 ;
  LAYER M2 ;
        RECT 9.004 0.824 9.716 0.856 ;
  LAYER M1 ;
        RECT 6.544 16.596 6.576 16.668 ;
  LAYER M2 ;
        RECT 6.524 16.616 6.596 16.648 ;
  LAYER M1 ;
        RECT 9.424 16.596 9.456 16.668 ;
  LAYER M2 ;
        RECT 9.404 16.616 9.476 16.648 ;
  LAYER M2 ;
        RECT 6.56 16.616 9.44 16.648 ;
  LAYER M2 ;
        RECT 7.1 29.636 7.3 29.668 ;
  LAYER M3 ;
        RECT 7.18 29.4 7.22 29.652 ;
  LAYER M4 ;
        RECT 7.13 29.38 7.27 29.42 ;
  LAYER M5 ;
        RECT 7.168 16.884 7.232 29.4 ;
  LAYER M4 ;
        RECT 7.13 16.864 7.27 16.904 ;
  LAYER M3 ;
        RECT 7.18 16.632 7.22 16.884 ;
  LAYER M2 ;
        RECT 7.1 16.616 7.3 16.648 ;
  LAYER M2 ;
        RECT 9.26 16.616 9.46 16.648 ;
  LAYER M3 ;
        RECT 9.34 1.512 9.38 16.632 ;
  LAYER M4 ;
        RECT 9.29 1.492 9.43 1.532 ;
  LAYER M5 ;
        RECT 9.328 1.344 9.392 1.512 ;
  LAYER M4 ;
        RECT 9.29 1.324 9.43 1.364 ;
  LAYER M3 ;
        RECT 9.34 0.84 9.38 1.344 ;
  LAYER M2 ;
        RECT 9.26 0.824 9.46 0.856 ;
  LAYER M1 ;
        RECT 9.504 17.352 9.536 17.424 ;
  LAYER M2 ;
        RECT 9.484 17.372 9.556 17.404 ;
  LAYER M1 ;
        RECT 6.624 17.352 6.656 17.424 ;
  LAYER M2 ;
        RECT 6.604 17.372 6.676 17.404 ;
  LAYER M2 ;
        RECT 6.64 17.372 9.52 17.404 ;
  LAYER M3 ;
        RECT 10.54 0.468 10.58 0.792 ;
  LAYER M3 ;
        RECT 10.3 0.468 10.34 0.792 ;
  LAYER M3 ;
        RECT 0.46 17.52 0.5 17.844 ;
  LAYER M3 ;
        RECT 0.22 17.52 0.26 17.844 ;
  LAYER M2 ;
        RECT 0.64 17.372 6.64 17.404 ;
  LAYER M3 ;
        RECT 0.62 17.283 0.66 17.493 ;
  LAYER M4 ;
        RECT 0.48 17.368 0.64 17.408 ;
  LAYER M3 ;
        RECT 0.46 17.388 0.5 17.64 ;
  LAYER M2 ;
        RECT 9.42 17.372 9.62 17.404 ;
  LAYER M3 ;
        RECT 9.5 0.756 9.54 17.388 ;
  LAYER M4 ;
        RECT 9.52 0.736 10.32 0.776 ;
  LAYER M3 ;
        RECT 10.3 0.651 10.34 0.861 ;
  LAYER M2 ;
        RECT 7.804 0.824 8.516 0.856 ;
  LAYER M1 ;
        RECT 6.704 1.392 6.736 1.464 ;
  LAYER M2 ;
        RECT 6.684 1.412 6.756 1.444 ;
  LAYER M1 ;
        RECT 9.584 1.392 9.616 1.464 ;
  LAYER M2 ;
        RECT 9.564 1.412 9.636 1.444 ;
  LAYER M2 ;
        RECT 6.72 1.412 9.6 1.444 ;
  LAYER M2 ;
        RECT 7.98 0.824 8.18 0.856 ;
  LAYER M3 ;
        RECT 8.06 0.84 8.1 1.344 ;
  LAYER M4 ;
        RECT 7.92 1.324 8.08 1.364 ;
  LAYER M5 ;
        RECT 7.888 1.336 7.952 1.436 ;
  LAYER M4 ;
        RECT 7.85 1.408 7.99 1.448 ;
  LAYER M3 ;
        RECT 7.9 1.323 7.94 1.533 ;
  LAYER M2 ;
        RECT 7.82 1.412 8.02 1.444 ;
  LAYER M1 ;
        RECT 6.784 20.796 6.816 20.868 ;
  LAYER M2 ;
        RECT 6.764 20.816 6.836 20.848 ;
  LAYER M2 ;
        RECT 6.8 20.816 9.52 20.848 ;
  LAYER M1 ;
        RECT 9.504 20.796 9.536 20.868 ;
  LAYER M2 ;
        RECT 9.484 20.816 9.556 20.848 ;
  LAYER M1 ;
        RECT 6.784 23.736 6.816 23.808 ;
  LAYER M2 ;
        RECT 6.764 23.756 6.836 23.788 ;
  LAYER M2 ;
        RECT 6.8 23.756 9.52 23.788 ;
  LAYER M1 ;
        RECT 9.504 23.736 9.536 23.808 ;
  LAYER M2 ;
        RECT 9.484 23.756 9.556 23.788 ;
  LAYER M1 ;
        RECT 9.664 20.796 9.696 20.868 ;
  LAYER M2 ;
        RECT 9.644 20.816 9.716 20.848 ;
  LAYER M1 ;
        RECT 9.664 20.664 9.696 20.832 ;
  LAYER M1 ;
        RECT 9.664 20.628 9.696 20.7 ;
  LAYER M2 ;
        RECT 9.644 20.648 9.716 20.68 ;
  LAYER M2 ;
        RECT 9.52 20.648 9.68 20.68 ;
  LAYER M1 ;
        RECT 9.504 20.628 9.536 20.7 ;
  LAYER M2 ;
        RECT 9.484 20.648 9.556 20.68 ;
  LAYER M1 ;
        RECT 9.664 23.736 9.696 23.808 ;
  LAYER M2 ;
        RECT 9.644 23.756 9.716 23.788 ;
  LAYER M1 ;
        RECT 9.664 23.604 9.696 23.772 ;
  LAYER M1 ;
        RECT 9.664 23.568 9.696 23.64 ;
  LAYER M2 ;
        RECT 9.644 23.588 9.716 23.62 ;
  LAYER M2 ;
        RECT 9.52 23.588 9.68 23.62 ;
  LAYER M1 ;
        RECT 9.504 23.568 9.536 23.64 ;
  LAYER M2 ;
        RECT 9.484 23.588 9.556 23.62 ;
  LAYER M1 ;
        RECT 9.504 17.352 9.536 17.424 ;
  LAYER M2 ;
        RECT 9.484 17.372 9.556 17.404 ;
  LAYER M1 ;
        RECT 9.504 17.388 9.536 17.556 ;
  LAYER M1 ;
        RECT 9.504 17.556 9.536 23.772 ;
  LAYER M1 ;
        RECT 3.904 23.736 3.936 23.808 ;
  LAYER M2 ;
        RECT 3.884 23.756 3.956 23.788 ;
  LAYER M2 ;
        RECT 3.92 23.756 6.64 23.788 ;
  LAYER M1 ;
        RECT 6.624 23.736 6.656 23.808 ;
  LAYER M2 ;
        RECT 6.604 23.756 6.676 23.788 ;
  LAYER M1 ;
        RECT 3.904 20.796 3.936 20.868 ;
  LAYER M2 ;
        RECT 3.884 20.816 3.956 20.848 ;
  LAYER M2 ;
        RECT 3.92 20.816 6.64 20.848 ;
  LAYER M1 ;
        RECT 6.624 20.796 6.656 20.868 ;
  LAYER M2 ;
        RECT 6.604 20.816 6.676 20.848 ;
  LAYER M1 ;
        RECT 6.624 17.352 6.656 17.424 ;
  LAYER M2 ;
        RECT 6.604 17.372 6.676 17.404 ;
  LAYER M1 ;
        RECT 6.624 17.388 6.656 17.556 ;
  LAYER M1 ;
        RECT 6.624 17.556 6.656 23.772 ;
  LAYER M2 ;
        RECT 6.64 17.372 9.52 17.404 ;
  LAYER M1 ;
        RECT 12.544 17.856 12.576 17.928 ;
  LAYER M2 ;
        RECT 12.524 17.876 12.596 17.908 ;
  LAYER M1 ;
        RECT 12.544 17.724 12.576 17.892 ;
  LAYER M1 ;
        RECT 12.544 17.688 12.576 17.76 ;
  LAYER M2 ;
        RECT 12.524 17.708 12.596 17.74 ;
  LAYER M2 ;
        RECT 12.4 17.708 12.56 17.74 ;
  LAYER M1 ;
        RECT 12.384 17.688 12.416 17.76 ;
  LAYER M2 ;
        RECT 12.364 17.708 12.436 17.74 ;
  LAYER M1 ;
        RECT 12.544 20.796 12.576 20.868 ;
  LAYER M2 ;
        RECT 12.524 20.816 12.596 20.848 ;
  LAYER M1 ;
        RECT 12.544 20.664 12.576 20.832 ;
  LAYER M1 ;
        RECT 12.544 20.628 12.576 20.7 ;
  LAYER M2 ;
        RECT 12.524 20.648 12.596 20.68 ;
  LAYER M2 ;
        RECT 12.4 20.648 12.56 20.68 ;
  LAYER M1 ;
        RECT 12.384 20.628 12.416 20.7 ;
  LAYER M2 ;
        RECT 12.364 20.648 12.436 20.68 ;
  LAYER M1 ;
        RECT 12.544 23.736 12.576 23.808 ;
  LAYER M2 ;
        RECT 12.524 23.756 12.596 23.788 ;
  LAYER M1 ;
        RECT 12.544 23.604 12.576 23.772 ;
  LAYER M1 ;
        RECT 12.544 23.568 12.576 23.64 ;
  LAYER M2 ;
        RECT 12.524 23.588 12.596 23.62 ;
  LAYER M2 ;
        RECT 12.4 23.588 12.56 23.62 ;
  LAYER M1 ;
        RECT 12.384 23.568 12.416 23.64 ;
  LAYER M2 ;
        RECT 12.364 23.588 12.436 23.62 ;
  LAYER M1 ;
        RECT 12.544 26.676 12.576 26.748 ;
  LAYER M2 ;
        RECT 12.524 26.696 12.596 26.728 ;
  LAYER M1 ;
        RECT 12.544 26.544 12.576 26.712 ;
  LAYER M1 ;
        RECT 12.544 26.508 12.576 26.58 ;
  LAYER M2 ;
        RECT 12.524 26.528 12.596 26.56 ;
  LAYER M2 ;
        RECT 12.4 26.528 12.56 26.56 ;
  LAYER M1 ;
        RECT 12.384 26.508 12.416 26.58 ;
  LAYER M2 ;
        RECT 12.364 26.528 12.436 26.56 ;
  LAYER M1 ;
        RECT 9.664 17.856 9.696 17.928 ;
  LAYER M2 ;
        RECT 9.644 17.876 9.716 17.908 ;
  LAYER M2 ;
        RECT 9.68 17.876 12.4 17.908 ;
  LAYER M1 ;
        RECT 12.384 17.856 12.416 17.928 ;
  LAYER M2 ;
        RECT 12.364 17.876 12.436 17.908 ;
  LAYER M1 ;
        RECT 9.664 26.676 9.696 26.748 ;
  LAYER M2 ;
        RECT 9.644 26.696 9.716 26.728 ;
  LAYER M2 ;
        RECT 9.68 26.696 12.4 26.728 ;
  LAYER M1 ;
        RECT 12.384 26.676 12.416 26.748 ;
  LAYER M2 ;
        RECT 12.364 26.696 12.436 26.728 ;
  LAYER M1 ;
        RECT 12.384 17.184 12.416 17.256 ;
  LAYER M2 ;
        RECT 12.364 17.204 12.436 17.236 ;
  LAYER M1 ;
        RECT 12.384 17.22 12.416 17.556 ;
  LAYER M1 ;
        RECT 12.384 17.556 12.416 26.712 ;
  LAYER M1 ;
        RECT 3.904 17.856 3.936 17.928 ;
  LAYER M2 ;
        RECT 3.884 17.876 3.956 17.908 ;
  LAYER M1 ;
        RECT 3.904 17.724 3.936 17.892 ;
  LAYER M1 ;
        RECT 3.904 17.688 3.936 17.76 ;
  LAYER M2 ;
        RECT 3.884 17.708 3.956 17.74 ;
  LAYER M2 ;
        RECT 3.76 17.708 3.92 17.74 ;
  LAYER M1 ;
        RECT 3.744 17.688 3.776 17.76 ;
  LAYER M2 ;
        RECT 3.724 17.708 3.796 17.74 ;
  LAYER M1 ;
        RECT 3.904 26.676 3.936 26.748 ;
  LAYER M2 ;
        RECT 3.884 26.696 3.956 26.728 ;
  LAYER M1 ;
        RECT 3.904 26.544 3.936 26.712 ;
  LAYER M1 ;
        RECT 3.904 26.508 3.936 26.58 ;
  LAYER M2 ;
        RECT 3.884 26.528 3.956 26.56 ;
  LAYER M2 ;
        RECT 3.76 26.528 3.92 26.56 ;
  LAYER M1 ;
        RECT 3.744 26.508 3.776 26.58 ;
  LAYER M2 ;
        RECT 3.724 26.528 3.796 26.56 ;
  LAYER M1 ;
        RECT 1.024 17.856 1.056 17.928 ;
  LAYER M2 ;
        RECT 1.004 17.876 1.076 17.908 ;
  LAYER M2 ;
        RECT 1.04 17.876 3.76 17.908 ;
  LAYER M1 ;
        RECT 3.744 17.856 3.776 17.928 ;
  LAYER M2 ;
        RECT 3.724 17.876 3.796 17.908 ;
  LAYER M1 ;
        RECT 1.024 20.796 1.056 20.868 ;
  LAYER M2 ;
        RECT 1.004 20.816 1.076 20.848 ;
  LAYER M2 ;
        RECT 1.04 20.816 3.76 20.848 ;
  LAYER M1 ;
        RECT 3.744 20.796 3.776 20.868 ;
  LAYER M2 ;
        RECT 3.724 20.816 3.796 20.848 ;
  LAYER M1 ;
        RECT 1.024 23.736 1.056 23.808 ;
  LAYER M2 ;
        RECT 1.004 23.756 1.076 23.788 ;
  LAYER M2 ;
        RECT 1.04 23.756 3.76 23.788 ;
  LAYER M1 ;
        RECT 3.744 23.736 3.776 23.808 ;
  LAYER M2 ;
        RECT 3.724 23.756 3.796 23.788 ;
  LAYER M1 ;
        RECT 1.024 26.676 1.056 26.748 ;
  LAYER M2 ;
        RECT 1.004 26.696 1.076 26.728 ;
  LAYER M2 ;
        RECT 1.04 26.696 3.76 26.728 ;
  LAYER M1 ;
        RECT 3.744 26.676 3.776 26.748 ;
  LAYER M2 ;
        RECT 3.724 26.696 3.796 26.728 ;
  LAYER M1 ;
        RECT 3.744 17.184 3.776 17.256 ;
  LAYER M2 ;
        RECT 3.724 17.204 3.796 17.236 ;
  LAYER M1 ;
        RECT 3.744 17.22 3.776 17.556 ;
  LAYER M1 ;
        RECT 3.744 17.556 3.776 26.712 ;
  LAYER M2 ;
        RECT 3.76 17.204 12.4 17.236 ;
  LAYER M1 ;
        RECT 6.784 26.676 6.816 26.748 ;
  LAYER M2 ;
        RECT 6.764 26.696 6.836 26.728 ;
  LAYER M2 ;
        RECT 6.8 26.696 9.68 26.728 ;
  LAYER M1 ;
        RECT 9.664 26.676 9.696 26.748 ;
  LAYER M2 ;
        RECT 9.644 26.696 9.716 26.728 ;
  LAYER M1 ;
        RECT 6.784 17.856 6.816 17.928 ;
  LAYER M2 ;
        RECT 6.764 17.876 6.836 17.908 ;
  LAYER M2 ;
        RECT 3.92 17.876 6.8 17.908 ;
  LAYER M1 ;
        RECT 3.904 17.856 3.936 17.928 ;
  LAYER M2 ;
        RECT 3.884 17.876 3.956 17.908 ;
  LAYER M1 ;
        RECT 9.184 23.232 9.216 23.304 ;
  LAYER M2 ;
        RECT 9.164 23.252 9.236 23.284 ;
  LAYER M2 ;
        RECT 9.2 23.252 9.36 23.284 ;
  LAYER M1 ;
        RECT 9.344 23.232 9.376 23.304 ;
  LAYER M2 ;
        RECT 9.324 23.252 9.396 23.284 ;
  LAYER M1 ;
        RECT 9.184 26.172 9.216 26.244 ;
  LAYER M2 ;
        RECT 9.164 26.192 9.236 26.224 ;
  LAYER M2 ;
        RECT 9.2 26.192 9.36 26.224 ;
  LAYER M1 ;
        RECT 9.344 26.172 9.376 26.244 ;
  LAYER M2 ;
        RECT 9.324 26.192 9.396 26.224 ;
  LAYER M1 ;
        RECT 12.064 23.232 12.096 23.304 ;
  LAYER M2 ;
        RECT 12.044 23.252 12.116 23.284 ;
  LAYER M1 ;
        RECT 12.064 23.268 12.096 23.436 ;
  LAYER M1 ;
        RECT 12.064 23.4 12.096 23.472 ;
  LAYER M2 ;
        RECT 12.044 23.42 12.116 23.452 ;
  LAYER M2 ;
        RECT 9.36 23.42 12.08 23.452 ;
  LAYER M1 ;
        RECT 9.344 23.4 9.376 23.472 ;
  LAYER M2 ;
        RECT 9.324 23.42 9.396 23.452 ;
  LAYER M1 ;
        RECT 12.064 26.172 12.096 26.244 ;
  LAYER M2 ;
        RECT 12.044 26.192 12.116 26.224 ;
  LAYER M1 ;
        RECT 12.064 26.208 12.096 26.376 ;
  LAYER M1 ;
        RECT 12.064 26.34 12.096 26.412 ;
  LAYER M2 ;
        RECT 12.044 26.36 12.116 26.392 ;
  LAYER M2 ;
        RECT 9.36 26.36 12.08 26.392 ;
  LAYER M1 ;
        RECT 9.344 26.34 9.376 26.412 ;
  LAYER M2 ;
        RECT 9.324 26.36 9.396 26.392 ;
  LAYER M1 ;
        RECT 9.344 29.616 9.376 29.688 ;
  LAYER M2 ;
        RECT 9.324 29.636 9.396 29.668 ;
  LAYER M1 ;
        RECT 9.344 29.484 9.376 29.652 ;
  LAYER M1 ;
        RECT 9.344 23.268 9.376 29.484 ;
  LAYER M1 ;
        RECT 6.304 26.172 6.336 26.244 ;
  LAYER M2 ;
        RECT 6.284 26.192 6.356 26.224 ;
  LAYER M2 ;
        RECT 6.32 26.192 6.48 26.224 ;
  LAYER M1 ;
        RECT 6.464 26.172 6.496 26.244 ;
  LAYER M2 ;
        RECT 6.444 26.192 6.516 26.224 ;
  LAYER M1 ;
        RECT 6.304 23.232 6.336 23.304 ;
  LAYER M2 ;
        RECT 6.284 23.252 6.356 23.284 ;
  LAYER M2 ;
        RECT 6.32 23.252 6.48 23.284 ;
  LAYER M1 ;
        RECT 6.464 23.232 6.496 23.304 ;
  LAYER M2 ;
        RECT 6.444 23.252 6.516 23.284 ;
  LAYER M1 ;
        RECT 6.464 29.616 6.496 29.688 ;
  LAYER M2 ;
        RECT 6.444 29.636 6.516 29.668 ;
  LAYER M1 ;
        RECT 6.464 29.484 6.496 29.652 ;
  LAYER M1 ;
        RECT 6.464 23.268 6.496 29.484 ;
  LAYER M2 ;
        RECT 6.48 29.636 9.36 29.668 ;
  LAYER M1 ;
        RECT 14.944 20.292 14.976 20.364 ;
  LAYER M2 ;
        RECT 14.924 20.312 14.996 20.344 ;
  LAYER M2 ;
        RECT 14.96 20.312 15.28 20.344 ;
  LAYER M1 ;
        RECT 15.264 20.292 15.296 20.364 ;
  LAYER M2 ;
        RECT 15.244 20.312 15.316 20.344 ;
  LAYER M1 ;
        RECT 14.944 23.232 14.976 23.304 ;
  LAYER M2 ;
        RECT 14.924 23.252 14.996 23.284 ;
  LAYER M2 ;
        RECT 14.96 23.252 15.28 23.284 ;
  LAYER M1 ;
        RECT 15.264 23.232 15.296 23.304 ;
  LAYER M2 ;
        RECT 15.244 23.252 15.316 23.284 ;
  LAYER M1 ;
        RECT 14.944 26.172 14.976 26.244 ;
  LAYER M2 ;
        RECT 14.924 26.192 14.996 26.224 ;
  LAYER M2 ;
        RECT 14.96 26.192 15.28 26.224 ;
  LAYER M1 ;
        RECT 15.264 26.172 15.296 26.244 ;
  LAYER M2 ;
        RECT 15.244 26.192 15.316 26.224 ;
  LAYER M1 ;
        RECT 14.944 29.112 14.976 29.184 ;
  LAYER M2 ;
        RECT 14.924 29.132 14.996 29.164 ;
  LAYER M2 ;
        RECT 14.96 29.132 15.28 29.164 ;
  LAYER M1 ;
        RECT 15.264 29.112 15.296 29.184 ;
  LAYER M2 ;
        RECT 15.244 29.132 15.316 29.164 ;
  LAYER M1 ;
        RECT 15.264 29.784 15.296 29.856 ;
  LAYER M2 ;
        RECT 15.244 29.804 15.316 29.836 ;
  LAYER M1 ;
        RECT 15.264 29.484 15.296 29.82 ;
  LAYER M1 ;
        RECT 15.264 20.328 15.296 29.484 ;
  LAYER M1 ;
        RECT 3.424 20.292 3.456 20.364 ;
  LAYER M2 ;
        RECT 3.404 20.312 3.476 20.344 ;
  LAYER M1 ;
        RECT 3.424 20.328 3.456 20.496 ;
  LAYER M1 ;
        RECT 3.424 20.46 3.456 20.532 ;
  LAYER M2 ;
        RECT 3.404 20.48 3.476 20.512 ;
  LAYER M2 ;
        RECT 0.88 20.48 3.44 20.512 ;
  LAYER M1 ;
        RECT 0.864 20.46 0.896 20.532 ;
  LAYER M2 ;
        RECT 0.844 20.48 0.916 20.512 ;
  LAYER M1 ;
        RECT 3.424 23.232 3.456 23.304 ;
  LAYER M2 ;
        RECT 3.404 23.252 3.476 23.284 ;
  LAYER M1 ;
        RECT 3.424 23.268 3.456 23.436 ;
  LAYER M1 ;
        RECT 3.424 23.4 3.456 23.472 ;
  LAYER M2 ;
        RECT 3.404 23.42 3.476 23.452 ;
  LAYER M2 ;
        RECT 0.88 23.42 3.44 23.452 ;
  LAYER M1 ;
        RECT 0.864 23.4 0.896 23.472 ;
  LAYER M2 ;
        RECT 0.844 23.42 0.916 23.452 ;
  LAYER M1 ;
        RECT 3.424 26.172 3.456 26.244 ;
  LAYER M2 ;
        RECT 3.404 26.192 3.476 26.224 ;
  LAYER M1 ;
        RECT 3.424 26.208 3.456 26.376 ;
  LAYER M1 ;
        RECT 3.424 26.34 3.456 26.412 ;
  LAYER M2 ;
        RECT 3.404 26.36 3.476 26.392 ;
  LAYER M2 ;
        RECT 0.88 26.36 3.44 26.392 ;
  LAYER M1 ;
        RECT 0.864 26.34 0.896 26.412 ;
  LAYER M2 ;
        RECT 0.844 26.36 0.916 26.392 ;
  LAYER M1 ;
        RECT 3.424 29.112 3.456 29.184 ;
  LAYER M2 ;
        RECT 3.404 29.132 3.476 29.164 ;
  LAYER M1 ;
        RECT 3.424 29.148 3.456 29.316 ;
  LAYER M1 ;
        RECT 3.424 29.28 3.456 29.352 ;
  LAYER M2 ;
        RECT 3.404 29.3 3.476 29.332 ;
  LAYER M2 ;
        RECT 0.88 29.3 3.44 29.332 ;
  LAYER M1 ;
        RECT 0.864 29.28 0.896 29.352 ;
  LAYER M2 ;
        RECT 0.844 29.3 0.916 29.332 ;
  LAYER M1 ;
        RECT 0.864 29.784 0.896 29.856 ;
  LAYER M2 ;
        RECT 0.844 29.804 0.916 29.836 ;
  LAYER M1 ;
        RECT 0.864 29.484 0.896 29.82 ;
  LAYER M1 ;
        RECT 0.864 20.496 0.896 29.484 ;
  LAYER M2 ;
        RECT 0.88 29.804 15.28 29.836 ;
  LAYER M1 ;
        RECT 12.064 20.292 12.096 20.364 ;
  LAYER M2 ;
        RECT 12.044 20.312 12.116 20.344 ;
  LAYER M2 ;
        RECT 12.08 20.312 14.96 20.344 ;
  LAYER M1 ;
        RECT 14.944 20.292 14.976 20.364 ;
  LAYER M2 ;
        RECT 14.924 20.312 14.996 20.344 ;
  LAYER M1 ;
        RECT 12.064 29.112 12.096 29.184 ;
  LAYER M2 ;
        RECT 12.044 29.132 12.116 29.164 ;
  LAYER M2 ;
        RECT 12.08 29.132 14.96 29.164 ;
  LAYER M1 ;
        RECT 14.944 29.112 14.976 29.184 ;
  LAYER M2 ;
        RECT 14.924 29.132 14.996 29.164 ;
  LAYER M1 ;
        RECT 9.184 29.112 9.216 29.184 ;
  LAYER M2 ;
        RECT 9.164 29.132 9.236 29.164 ;
  LAYER M2 ;
        RECT 9.2 29.132 12.08 29.164 ;
  LAYER M1 ;
        RECT 12.064 29.112 12.096 29.184 ;
  LAYER M2 ;
        RECT 12.044 29.132 12.116 29.164 ;
  LAYER M1 ;
        RECT 6.304 29.112 6.336 29.184 ;
  LAYER M2 ;
        RECT 6.284 29.132 6.356 29.164 ;
  LAYER M2 ;
        RECT 6.32 29.132 9.2 29.164 ;
  LAYER M1 ;
        RECT 9.184 29.112 9.216 29.184 ;
  LAYER M2 ;
        RECT 9.164 29.132 9.236 29.164 ;
  LAYER M1 ;
        RECT 6.304 20.292 6.336 20.364 ;
  LAYER M2 ;
        RECT 6.284 20.312 6.356 20.344 ;
  LAYER M2 ;
        RECT 3.44 20.312 6.32 20.344 ;
  LAYER M1 ;
        RECT 3.424 20.292 3.456 20.364 ;
  LAYER M2 ;
        RECT 3.404 20.312 3.476 20.344 ;
  LAYER M1 ;
        RECT 9.184 20.292 9.216 20.364 ;
  LAYER M2 ;
        RECT 9.164 20.312 9.236 20.344 ;
  LAYER M2 ;
        RECT 6.32 20.312 9.2 20.344 ;
  LAYER M1 ;
        RECT 6.304 20.292 6.336 20.364 ;
  LAYER M2 ;
        RECT 6.284 20.312 6.356 20.344 ;
  LAYER M1 ;
        RECT 12.56 17.892 14.96 20.328 ;
  LAYER M2 ;
        RECT 12.56 17.892 14.96 20.328 ;
  LAYER M3 ;
        RECT 12.56 17.892 14.96 20.328 ;
  LAYER M1 ;
        RECT 12.56 20.832 14.96 23.268 ;
  LAYER M2 ;
        RECT 12.56 20.832 14.96 23.268 ;
  LAYER M3 ;
        RECT 12.56 20.832 14.96 23.268 ;
  LAYER M1 ;
        RECT 12.56 23.772 14.96 26.208 ;
  LAYER M2 ;
        RECT 12.56 23.772 14.96 26.208 ;
  LAYER M3 ;
        RECT 12.56 23.772 14.96 26.208 ;
  LAYER M1 ;
        RECT 12.56 26.712 14.96 29.148 ;
  LAYER M2 ;
        RECT 12.56 26.712 14.96 29.148 ;
  LAYER M3 ;
        RECT 12.56 26.712 14.96 29.148 ;
  LAYER M1 ;
        RECT 9.68 17.892 12.08 20.328 ;
  LAYER M2 ;
        RECT 9.68 17.892 12.08 20.328 ;
  LAYER M3 ;
        RECT 9.68 17.892 12.08 20.328 ;
  LAYER M1 ;
        RECT 9.68 20.832 12.08 23.268 ;
  LAYER M2 ;
        RECT 9.68 20.832 12.08 23.268 ;
  LAYER M3 ;
        RECT 9.68 20.832 12.08 23.268 ;
  LAYER M1 ;
        RECT 9.68 23.772 12.08 26.208 ;
  LAYER M2 ;
        RECT 9.68 23.772 12.08 26.208 ;
  LAYER M3 ;
        RECT 9.68 23.772 12.08 26.208 ;
  LAYER M1 ;
        RECT 9.68 26.712 12.08 29.148 ;
  LAYER M2 ;
        RECT 9.68 26.712 12.08 29.148 ;
  LAYER M3 ;
        RECT 9.68 26.712 12.08 29.148 ;
  LAYER M1 ;
        RECT 6.8 17.892 9.2 20.328 ;
  LAYER M2 ;
        RECT 6.8 17.892 9.2 20.328 ;
  LAYER M3 ;
        RECT 6.8 17.892 9.2 20.328 ;
  LAYER M1 ;
        RECT 6.8 20.832 9.2 23.268 ;
  LAYER M2 ;
        RECT 6.8 20.832 9.2 23.268 ;
  LAYER M3 ;
        RECT 6.8 20.832 9.2 23.268 ;
  LAYER M1 ;
        RECT 6.8 23.772 9.2 26.208 ;
  LAYER M2 ;
        RECT 6.8 23.772 9.2 26.208 ;
  LAYER M3 ;
        RECT 6.8 23.772 9.2 26.208 ;
  LAYER M1 ;
        RECT 6.8 26.712 9.2 29.148 ;
  LAYER M2 ;
        RECT 6.8 26.712 9.2 29.148 ;
  LAYER M3 ;
        RECT 6.8 26.712 9.2 29.148 ;
  LAYER M1 ;
        RECT 3.92 17.892 6.32 20.328 ;
  LAYER M2 ;
        RECT 3.92 17.892 6.32 20.328 ;
  LAYER M3 ;
        RECT 3.92 17.892 6.32 20.328 ;
  LAYER M1 ;
        RECT 3.92 20.832 6.32 23.268 ;
  LAYER M2 ;
        RECT 3.92 20.832 6.32 23.268 ;
  LAYER M3 ;
        RECT 3.92 20.832 6.32 23.268 ;
  LAYER M1 ;
        RECT 3.92 23.772 6.32 26.208 ;
  LAYER M2 ;
        RECT 3.92 23.772 6.32 26.208 ;
  LAYER M3 ;
        RECT 3.92 23.772 6.32 26.208 ;
  LAYER M1 ;
        RECT 3.92 26.712 6.32 29.148 ;
  LAYER M2 ;
        RECT 3.92 26.712 6.32 29.148 ;
  LAYER M3 ;
        RECT 3.92 26.712 6.32 29.148 ;
  LAYER M1 ;
        RECT 1.04 17.892 3.44 20.328 ;
  LAYER M2 ;
        RECT 1.04 17.892 3.44 20.328 ;
  LAYER M3 ;
        RECT 1.04 17.892 3.44 20.328 ;
  LAYER M1 ;
        RECT 1.04 20.832 3.44 23.268 ;
  LAYER M2 ;
        RECT 1.04 20.832 3.44 23.268 ;
  LAYER M3 ;
        RECT 1.04 20.832 3.44 23.268 ;
  LAYER M1 ;
        RECT 1.04 23.772 3.44 26.208 ;
  LAYER M2 ;
        RECT 1.04 23.772 3.44 26.208 ;
  LAYER M3 ;
        RECT 1.04 23.772 3.44 26.208 ;
  LAYER M1 ;
        RECT 1.04 26.712 3.44 29.148 ;
  LAYER M2 ;
        RECT 1.04 26.712 3.44 29.148 ;
  LAYER M3 ;
        RECT 1.04 26.712 3.44 29.148 ;
  LAYER M1 ;
        RECT 10.464 0.216 10.496 0.876 ;
  LAYER M1 ;
        RECT 10.544 0.216 10.576 0.876 ;
  LAYER M1 ;
        RECT 10.384 0.216 10.416 0.876 ;
  LAYER M2 ;
        RECT 10.364 0.824 10.676 0.856 ;
  LAYER M2 ;
        RECT 10.364 0.572 10.676 0.604 ;
  LAYER M2 ;
        RECT 10.284 0.74 10.596 0.772 ;
  LAYER M2 ;
        RECT 10.284 0.488 10.596 0.52 ;
  LAYER M2 ;
        RECT 10.204 0.656 10.596 0.688 ;
  LAYER M2 ;
        RECT 10.204 0.404 10.596 0.436 ;
  LAYER M1 ;
        RECT 0.384 17.268 0.416 17.928 ;
  LAYER M1 ;
        RECT 0.464 17.268 0.496 17.928 ;
  LAYER M1 ;
        RECT 0.304 17.268 0.336 17.928 ;
  LAYER M2 ;
        RECT 0.284 17.876 0.596 17.908 ;
  LAYER M2 ;
        RECT 0.284 17.624 0.596 17.656 ;
  LAYER M2 ;
        RECT 0.204 17.792 0.516 17.824 ;
  LAYER M2 ;
        RECT 0.204 17.54 0.516 17.572 ;
  LAYER M2 ;
        RECT 0.124 17.708 0.516 17.74 ;
  LAYER M2 ;
        RECT 0.124 17.456 0.516 17.488 ;
  LAYER M1 ;
        RECT 9.104 0.216 9.136 0.876 ;
  LAYER M1 ;
        RECT 9.024 0.216 9.056 0.876 ;
  LAYER M1 ;
        RECT 9.184 0.216 9.216 0.876 ;
  LAYER M1 ;
        RECT 9.744 0.216 9.776 0.876 ;
  LAYER M1 ;
        RECT 9.664 0.216 9.696 0.876 ;
  LAYER M1 ;
        RECT 9.824 0.216 9.856 0.876 ;
  LAYER M1 ;
        RECT 8.384 0.216 8.416 0.876 ;
  LAYER M1 ;
        RECT 8.464 0.216 8.496 0.876 ;
  LAYER M1 ;
        RECT 8.304 0.216 8.336 0.876 ;
  LAYER M1 ;
        RECT 7.744 0.216 7.776 0.876 ;
  LAYER M1 ;
        RECT 7.824 0.216 7.856 0.876 ;
  LAYER M1 ;
        RECT 7.664 0.216 7.696 0.876 ;
  LAYER M1 ;
        RECT 9.264 10.212 9.296 10.284 ;
  LAYER M2 ;
        RECT 9.244 10.232 9.316 10.264 ;
  LAYER M2 ;
        RECT 6.56 10.232 9.28 10.264 ;
  LAYER M1 ;
        RECT 6.544 10.212 6.576 10.284 ;
  LAYER M2 ;
        RECT 6.524 10.232 6.596 10.264 ;
  LAYER M1 ;
        RECT 6.384 7.272 6.416 7.344 ;
  LAYER M2 ;
        RECT 6.364 7.292 6.436 7.324 ;
  LAYER M1 ;
        RECT 6.384 7.308 6.416 7.476 ;
  LAYER M1 ;
        RECT 6.384 7.44 6.416 7.512 ;
  LAYER M2 ;
        RECT 6.364 7.46 6.436 7.492 ;
  LAYER M2 ;
        RECT 6.4 7.46 6.56 7.492 ;
  LAYER M1 ;
        RECT 6.544 7.44 6.576 7.512 ;
  LAYER M2 ;
        RECT 6.524 7.46 6.596 7.492 ;
  LAYER M1 ;
        RECT 6.544 16.596 6.576 16.668 ;
  LAYER M2 ;
        RECT 6.524 16.616 6.596 16.648 ;
  LAYER M1 ;
        RECT 6.544 16.464 6.576 16.632 ;
  LAYER M1 ;
        RECT 6.544 7.476 6.576 16.464 ;
  LAYER M1 ;
        RECT 12.144 13.152 12.176 13.224 ;
  LAYER M2 ;
        RECT 12.124 13.172 12.196 13.204 ;
  LAYER M2 ;
        RECT 9.44 13.172 12.16 13.204 ;
  LAYER M1 ;
        RECT 9.424 13.152 9.456 13.224 ;
  LAYER M2 ;
        RECT 9.404 13.172 9.476 13.204 ;
  LAYER M1 ;
        RECT 9.424 16.596 9.456 16.668 ;
  LAYER M2 ;
        RECT 9.404 16.616 9.476 16.648 ;
  LAYER M1 ;
        RECT 9.424 16.464 9.456 16.632 ;
  LAYER M1 ;
        RECT 9.424 13.188 9.456 16.464 ;
  LAYER M2 ;
        RECT 6.56 16.616 9.44 16.648 ;
  LAYER M1 ;
        RECT 6.384 10.212 6.416 10.284 ;
  LAYER M2 ;
        RECT 6.364 10.232 6.436 10.264 ;
  LAYER M2 ;
        RECT 3.68 10.232 6.4 10.264 ;
  LAYER M1 ;
        RECT 3.664 10.212 3.696 10.284 ;
  LAYER M2 ;
        RECT 3.644 10.232 3.716 10.264 ;
  LAYER M1 ;
        RECT 6.384 13.152 6.416 13.224 ;
  LAYER M2 ;
        RECT 6.364 13.172 6.436 13.204 ;
  LAYER M2 ;
        RECT 3.68 13.172 6.4 13.204 ;
  LAYER M1 ;
        RECT 3.664 13.152 3.696 13.224 ;
  LAYER M2 ;
        RECT 3.644 13.172 3.716 13.204 ;
  LAYER M1 ;
        RECT 3.664 16.764 3.696 16.836 ;
  LAYER M2 ;
        RECT 3.644 16.784 3.716 16.816 ;
  LAYER M1 ;
        RECT 3.664 16.464 3.696 16.8 ;
  LAYER M1 ;
        RECT 3.664 10.248 3.696 16.464 ;
  LAYER M1 ;
        RECT 12.144 10.212 12.176 10.284 ;
  LAYER M2 ;
        RECT 12.124 10.232 12.196 10.264 ;
  LAYER M1 ;
        RECT 12.144 10.248 12.176 10.416 ;
  LAYER M1 ;
        RECT 12.144 10.38 12.176 10.452 ;
  LAYER M2 ;
        RECT 12.124 10.4 12.196 10.432 ;
  LAYER M2 ;
        RECT 12.16 10.4 12.32 10.432 ;
  LAYER M1 ;
        RECT 12.304 10.38 12.336 10.452 ;
  LAYER M2 ;
        RECT 12.284 10.4 12.356 10.432 ;
  LAYER M1 ;
        RECT 12.144 7.272 12.176 7.344 ;
  LAYER M2 ;
        RECT 12.124 7.292 12.196 7.324 ;
  LAYER M1 ;
        RECT 12.144 7.308 12.176 7.476 ;
  LAYER M1 ;
        RECT 12.144 7.44 12.176 7.512 ;
  LAYER M2 ;
        RECT 12.124 7.46 12.196 7.492 ;
  LAYER M2 ;
        RECT 12.16 7.46 12.32 7.492 ;
  LAYER M1 ;
        RECT 12.304 7.44 12.336 7.512 ;
  LAYER M2 ;
        RECT 12.284 7.46 12.356 7.492 ;
  LAYER M1 ;
        RECT 12.304 16.764 12.336 16.836 ;
  LAYER M2 ;
        RECT 12.284 16.784 12.356 16.816 ;
  LAYER M1 ;
        RECT 12.304 16.464 12.336 16.8 ;
  LAYER M1 ;
        RECT 12.304 7.476 12.336 16.464 ;
  LAYER M2 ;
        RECT 3.68 16.784 12.32 16.816 ;
  LAYER M1 ;
        RECT 9.264 13.152 9.296 13.224 ;
  LAYER M2 ;
        RECT 9.244 13.172 9.316 13.204 ;
  LAYER M2 ;
        RECT 6.4 13.172 9.28 13.204 ;
  LAYER M1 ;
        RECT 6.384 13.152 6.416 13.224 ;
  LAYER M2 ;
        RECT 6.364 13.172 6.436 13.204 ;
  LAYER M1 ;
        RECT 9.264 7.272 9.296 7.344 ;
  LAYER M2 ;
        RECT 9.244 7.292 9.316 7.324 ;
  LAYER M2 ;
        RECT 9.28 7.292 12.16 7.324 ;
  LAYER M1 ;
        RECT 12.144 7.272 12.176 7.344 ;
  LAYER M2 ;
        RECT 12.124 7.292 12.196 7.324 ;
  LAYER M1 ;
        RECT 3.504 16.092 3.536 16.164 ;
  LAYER M2 ;
        RECT 3.484 16.112 3.556 16.144 ;
  LAYER M2 ;
        RECT 0.8 16.112 3.52 16.144 ;
  LAYER M1 ;
        RECT 0.784 16.092 0.816 16.164 ;
  LAYER M2 ;
        RECT 0.764 16.112 0.836 16.144 ;
  LAYER M1 ;
        RECT 3.504 13.152 3.536 13.224 ;
  LAYER M2 ;
        RECT 3.484 13.172 3.556 13.204 ;
  LAYER M2 ;
        RECT 0.8 13.172 3.52 13.204 ;
  LAYER M1 ;
        RECT 0.784 13.152 0.816 13.224 ;
  LAYER M2 ;
        RECT 0.764 13.172 0.836 13.204 ;
  LAYER M1 ;
        RECT 3.504 10.212 3.536 10.284 ;
  LAYER M2 ;
        RECT 3.484 10.232 3.556 10.264 ;
  LAYER M2 ;
        RECT 0.8 10.232 3.52 10.264 ;
  LAYER M1 ;
        RECT 0.784 10.212 0.816 10.284 ;
  LAYER M2 ;
        RECT 0.764 10.232 0.836 10.264 ;
  LAYER M1 ;
        RECT 3.504 7.272 3.536 7.344 ;
  LAYER M2 ;
        RECT 3.484 7.292 3.556 7.324 ;
  LAYER M2 ;
        RECT 0.8 7.292 3.52 7.324 ;
  LAYER M1 ;
        RECT 0.784 7.272 0.816 7.344 ;
  LAYER M2 ;
        RECT 0.764 7.292 0.836 7.324 ;
  LAYER M1 ;
        RECT 3.504 4.332 3.536 4.404 ;
  LAYER M2 ;
        RECT 3.484 4.352 3.556 4.384 ;
  LAYER M2 ;
        RECT 0.8 4.352 3.52 4.384 ;
  LAYER M1 ;
        RECT 0.784 4.332 0.816 4.404 ;
  LAYER M2 ;
        RECT 0.764 4.352 0.836 4.384 ;
  LAYER M1 ;
        RECT 0.784 16.932 0.816 17.004 ;
  LAYER M2 ;
        RECT 0.764 16.952 0.836 16.984 ;
  LAYER M1 ;
        RECT 0.784 16.464 0.816 16.968 ;
  LAYER M1 ;
        RECT 0.784 4.368 0.816 16.464 ;
  LAYER M1 ;
        RECT 15.024 16.092 15.056 16.164 ;
  LAYER M2 ;
        RECT 15.004 16.112 15.076 16.144 ;
  LAYER M1 ;
        RECT 15.024 16.128 15.056 16.296 ;
  LAYER M1 ;
        RECT 15.024 16.26 15.056 16.332 ;
  LAYER M2 ;
        RECT 15.004 16.28 15.076 16.312 ;
  LAYER M2 ;
        RECT 15.04 16.28 15.2 16.312 ;
  LAYER M1 ;
        RECT 15.184 16.26 15.216 16.332 ;
  LAYER M2 ;
        RECT 15.164 16.28 15.236 16.312 ;
  LAYER M1 ;
        RECT 15.024 13.152 15.056 13.224 ;
  LAYER M2 ;
        RECT 15.004 13.172 15.076 13.204 ;
  LAYER M1 ;
        RECT 15.024 13.188 15.056 13.356 ;
  LAYER M1 ;
        RECT 15.024 13.32 15.056 13.392 ;
  LAYER M2 ;
        RECT 15.004 13.34 15.076 13.372 ;
  LAYER M2 ;
        RECT 15.04 13.34 15.2 13.372 ;
  LAYER M1 ;
        RECT 15.184 13.32 15.216 13.392 ;
  LAYER M2 ;
        RECT 15.164 13.34 15.236 13.372 ;
  LAYER M1 ;
        RECT 15.024 10.212 15.056 10.284 ;
  LAYER M2 ;
        RECT 15.004 10.232 15.076 10.264 ;
  LAYER M1 ;
        RECT 15.024 10.248 15.056 10.416 ;
  LAYER M1 ;
        RECT 15.024 10.38 15.056 10.452 ;
  LAYER M2 ;
        RECT 15.004 10.4 15.076 10.432 ;
  LAYER M2 ;
        RECT 15.04 10.4 15.2 10.432 ;
  LAYER M1 ;
        RECT 15.184 10.38 15.216 10.452 ;
  LAYER M2 ;
        RECT 15.164 10.4 15.236 10.432 ;
  LAYER M1 ;
        RECT 15.024 7.272 15.056 7.344 ;
  LAYER M2 ;
        RECT 15.004 7.292 15.076 7.324 ;
  LAYER M1 ;
        RECT 15.024 7.308 15.056 7.476 ;
  LAYER M1 ;
        RECT 15.024 7.44 15.056 7.512 ;
  LAYER M2 ;
        RECT 15.004 7.46 15.076 7.492 ;
  LAYER M2 ;
        RECT 15.04 7.46 15.2 7.492 ;
  LAYER M1 ;
        RECT 15.184 7.44 15.216 7.512 ;
  LAYER M2 ;
        RECT 15.164 7.46 15.236 7.492 ;
  LAYER M1 ;
        RECT 15.024 4.332 15.056 4.404 ;
  LAYER M2 ;
        RECT 15.004 4.352 15.076 4.384 ;
  LAYER M1 ;
        RECT 15.024 4.368 15.056 4.536 ;
  LAYER M1 ;
        RECT 15.024 4.5 15.056 4.572 ;
  LAYER M2 ;
        RECT 15.004 4.52 15.076 4.552 ;
  LAYER M2 ;
        RECT 15.04 4.52 15.2 4.552 ;
  LAYER M1 ;
        RECT 15.184 4.5 15.216 4.572 ;
  LAYER M2 ;
        RECT 15.164 4.52 15.236 4.552 ;
  LAYER M1 ;
        RECT 15.184 16.932 15.216 17.004 ;
  LAYER M2 ;
        RECT 15.164 16.952 15.236 16.984 ;
  LAYER M1 ;
        RECT 15.184 16.464 15.216 16.968 ;
  LAYER M1 ;
        RECT 15.184 4.536 15.216 16.464 ;
  LAYER M2 ;
        RECT 0.8 16.952 15.2 16.984 ;
  LAYER M1 ;
        RECT 6.384 16.092 6.416 16.164 ;
  LAYER M2 ;
        RECT 6.364 16.112 6.436 16.144 ;
  LAYER M2 ;
        RECT 3.52 16.112 6.4 16.144 ;
  LAYER M1 ;
        RECT 3.504 16.092 3.536 16.164 ;
  LAYER M2 ;
        RECT 3.484 16.112 3.556 16.144 ;
  LAYER M1 ;
        RECT 6.384 4.332 6.416 4.404 ;
  LAYER M2 ;
        RECT 6.364 4.352 6.436 4.384 ;
  LAYER M2 ;
        RECT 3.52 4.352 6.4 4.384 ;
  LAYER M1 ;
        RECT 3.504 4.332 3.536 4.404 ;
  LAYER M2 ;
        RECT 3.484 4.352 3.556 4.384 ;
  LAYER M1 ;
        RECT 9.264 4.332 9.296 4.404 ;
  LAYER M2 ;
        RECT 9.244 4.352 9.316 4.384 ;
  LAYER M2 ;
        RECT 6.4 4.352 9.28 4.384 ;
  LAYER M1 ;
        RECT 6.384 4.332 6.416 4.404 ;
  LAYER M2 ;
        RECT 6.364 4.352 6.436 4.384 ;
  LAYER M1 ;
        RECT 12.144 4.332 12.176 4.404 ;
  LAYER M2 ;
        RECT 12.124 4.352 12.196 4.384 ;
  LAYER M2 ;
        RECT 9.28 4.352 12.16 4.384 ;
  LAYER M1 ;
        RECT 9.264 4.332 9.296 4.404 ;
  LAYER M2 ;
        RECT 9.244 4.352 9.316 4.384 ;
  LAYER M1 ;
        RECT 12.144 16.092 12.176 16.164 ;
  LAYER M2 ;
        RECT 12.124 16.112 12.196 16.144 ;
  LAYER M2 ;
        RECT 12.16 16.112 15.04 16.144 ;
  LAYER M1 ;
        RECT 15.024 16.092 15.056 16.164 ;
  LAYER M2 ;
        RECT 15.004 16.112 15.076 16.144 ;
  LAYER M1 ;
        RECT 9.264 16.092 9.296 16.164 ;
  LAYER M2 ;
        RECT 9.244 16.112 9.316 16.144 ;
  LAYER M2 ;
        RECT 9.28 16.112 12.16 16.144 ;
  LAYER M1 ;
        RECT 12.144 16.092 12.176 16.164 ;
  LAYER M2 ;
        RECT 12.124 16.112 12.196 16.144 ;
  LAYER M1 ;
        RECT 6.864 7.776 6.896 7.848 ;
  LAYER M2 ;
        RECT 6.844 7.796 6.916 7.828 ;
  LAYER M2 ;
        RECT 6.72 7.796 6.88 7.828 ;
  LAYER M1 ;
        RECT 6.704 7.776 6.736 7.848 ;
  LAYER M2 ;
        RECT 6.684 7.796 6.756 7.828 ;
  LAYER M1 ;
        RECT 3.984 4.836 4.016 4.908 ;
  LAYER M2 ;
        RECT 3.964 4.856 4.036 4.888 ;
  LAYER M1 ;
        RECT 3.984 4.704 4.016 4.872 ;
  LAYER M1 ;
        RECT 3.984 4.668 4.016 4.74 ;
  LAYER M2 ;
        RECT 3.964 4.688 4.036 4.72 ;
  LAYER M2 ;
        RECT 4 4.688 6.72 4.72 ;
  LAYER M1 ;
        RECT 6.704 4.668 6.736 4.74 ;
  LAYER M2 ;
        RECT 6.684 4.688 6.756 4.72 ;
  LAYER M1 ;
        RECT 6.704 1.392 6.736 1.464 ;
  LAYER M2 ;
        RECT 6.684 1.412 6.756 1.444 ;
  LAYER M1 ;
        RECT 6.704 1.428 6.736 1.596 ;
  LAYER M1 ;
        RECT 6.704 1.596 6.736 7.812 ;
  LAYER M1 ;
        RECT 9.744 10.716 9.776 10.788 ;
  LAYER M2 ;
        RECT 9.724 10.736 9.796 10.768 ;
  LAYER M2 ;
        RECT 9.6 10.736 9.76 10.768 ;
  LAYER M1 ;
        RECT 9.584 10.716 9.616 10.788 ;
  LAYER M2 ;
        RECT 9.564 10.736 9.636 10.768 ;
  LAYER M1 ;
        RECT 9.584 1.392 9.616 1.464 ;
  LAYER M2 ;
        RECT 9.564 1.412 9.636 1.444 ;
  LAYER M1 ;
        RECT 9.584 1.428 9.616 1.596 ;
  LAYER M1 ;
        RECT 9.584 1.596 9.616 10.752 ;
  LAYER M2 ;
        RECT 6.72 1.412 9.6 1.444 ;
  LAYER M1 ;
        RECT 3.984 7.776 4.016 7.848 ;
  LAYER M2 ;
        RECT 3.964 7.796 4.036 7.828 ;
  LAYER M2 ;
        RECT 3.84 7.796 4 7.828 ;
  LAYER M1 ;
        RECT 3.824 7.776 3.856 7.848 ;
  LAYER M2 ;
        RECT 3.804 7.796 3.876 7.828 ;
  LAYER M1 ;
        RECT 3.984 10.716 4.016 10.788 ;
  LAYER M2 ;
        RECT 3.964 10.736 4.036 10.768 ;
  LAYER M2 ;
        RECT 3.84 10.736 4 10.768 ;
  LAYER M1 ;
        RECT 3.824 10.716 3.856 10.788 ;
  LAYER M2 ;
        RECT 3.804 10.736 3.876 10.768 ;
  LAYER M1 ;
        RECT 3.824 1.224 3.856 1.296 ;
  LAYER M2 ;
        RECT 3.804 1.244 3.876 1.276 ;
  LAYER M1 ;
        RECT 3.824 1.26 3.856 1.596 ;
  LAYER M1 ;
        RECT 3.824 1.596 3.856 10.752 ;
  LAYER M1 ;
        RECT 9.744 7.776 9.776 7.848 ;
  LAYER M2 ;
        RECT 9.724 7.796 9.796 7.828 ;
  LAYER M1 ;
        RECT 9.744 7.644 9.776 7.812 ;
  LAYER M1 ;
        RECT 9.744 7.608 9.776 7.68 ;
  LAYER M2 ;
        RECT 9.724 7.628 9.796 7.66 ;
  LAYER M2 ;
        RECT 9.76 7.628 12.48 7.66 ;
  LAYER M1 ;
        RECT 12.464 7.608 12.496 7.68 ;
  LAYER M2 ;
        RECT 12.444 7.628 12.516 7.66 ;
  LAYER M1 ;
        RECT 9.744 4.836 9.776 4.908 ;
  LAYER M2 ;
        RECT 9.724 4.856 9.796 4.888 ;
  LAYER M1 ;
        RECT 9.744 4.704 9.776 4.872 ;
  LAYER M1 ;
        RECT 9.744 4.668 9.776 4.74 ;
  LAYER M2 ;
        RECT 9.724 4.688 9.796 4.72 ;
  LAYER M2 ;
        RECT 9.76 4.688 12.48 4.72 ;
  LAYER M1 ;
        RECT 12.464 4.668 12.496 4.74 ;
  LAYER M2 ;
        RECT 12.444 4.688 12.516 4.72 ;
  LAYER M1 ;
        RECT 12.464 1.224 12.496 1.296 ;
  LAYER M2 ;
        RECT 12.444 1.244 12.516 1.276 ;
  LAYER M1 ;
        RECT 12.464 1.26 12.496 1.596 ;
  LAYER M1 ;
        RECT 12.464 1.596 12.496 7.644 ;
  LAYER M2 ;
        RECT 3.84 1.244 12.48 1.276 ;
  LAYER M1 ;
        RECT 6.864 10.716 6.896 10.788 ;
  LAYER M2 ;
        RECT 6.844 10.736 6.916 10.768 ;
  LAYER M2 ;
        RECT 4 10.736 6.88 10.768 ;
  LAYER M1 ;
        RECT 3.984 10.716 4.016 10.788 ;
  LAYER M2 ;
        RECT 3.964 10.736 4.036 10.768 ;
  LAYER M1 ;
        RECT 6.864 4.836 6.896 4.908 ;
  LAYER M2 ;
        RECT 6.844 4.856 6.916 4.888 ;
  LAYER M2 ;
        RECT 6.88 4.856 9.76 4.888 ;
  LAYER M1 ;
        RECT 9.744 4.836 9.776 4.908 ;
  LAYER M2 ;
        RECT 9.724 4.856 9.796 4.888 ;
  LAYER M1 ;
        RECT 1.104 13.656 1.136 13.728 ;
  LAYER M2 ;
        RECT 1.084 13.676 1.156 13.708 ;
  LAYER M2 ;
        RECT 0.96 13.676 1.12 13.708 ;
  LAYER M1 ;
        RECT 0.944 13.656 0.976 13.728 ;
  LAYER M2 ;
        RECT 0.924 13.676 0.996 13.708 ;
  LAYER M1 ;
        RECT 1.104 10.716 1.136 10.788 ;
  LAYER M2 ;
        RECT 1.084 10.736 1.156 10.768 ;
  LAYER M2 ;
        RECT 0.96 10.736 1.12 10.768 ;
  LAYER M1 ;
        RECT 0.944 10.716 0.976 10.788 ;
  LAYER M2 ;
        RECT 0.924 10.736 0.996 10.768 ;
  LAYER M1 ;
        RECT 1.104 7.776 1.136 7.848 ;
  LAYER M2 ;
        RECT 1.084 7.796 1.156 7.828 ;
  LAYER M2 ;
        RECT 0.96 7.796 1.12 7.828 ;
  LAYER M1 ;
        RECT 0.944 7.776 0.976 7.848 ;
  LAYER M2 ;
        RECT 0.924 7.796 0.996 7.828 ;
  LAYER M1 ;
        RECT 1.104 4.836 1.136 4.908 ;
  LAYER M2 ;
        RECT 1.084 4.856 1.156 4.888 ;
  LAYER M2 ;
        RECT 0.96 4.856 1.12 4.888 ;
  LAYER M1 ;
        RECT 0.944 4.836 0.976 4.908 ;
  LAYER M2 ;
        RECT 0.924 4.856 0.996 4.888 ;
  LAYER M1 ;
        RECT 1.104 1.896 1.136 1.968 ;
  LAYER M2 ;
        RECT 1.084 1.916 1.156 1.948 ;
  LAYER M2 ;
        RECT 0.96 1.916 1.12 1.948 ;
  LAYER M1 ;
        RECT 0.944 1.896 0.976 1.968 ;
  LAYER M2 ;
        RECT 0.924 1.916 0.996 1.948 ;
  LAYER M1 ;
        RECT 0.944 1.056 0.976 1.128 ;
  LAYER M2 ;
        RECT 0.924 1.076 0.996 1.108 ;
  LAYER M1 ;
        RECT 0.944 1.092 0.976 1.596 ;
  LAYER M1 ;
        RECT 0.944 1.596 0.976 13.692 ;
  LAYER M1 ;
        RECT 12.624 13.656 12.656 13.728 ;
  LAYER M2 ;
        RECT 12.604 13.676 12.676 13.708 ;
  LAYER M1 ;
        RECT 12.624 13.524 12.656 13.692 ;
  LAYER M1 ;
        RECT 12.624 13.488 12.656 13.56 ;
  LAYER M2 ;
        RECT 12.604 13.508 12.676 13.54 ;
  LAYER M2 ;
        RECT 12.64 13.508 15.36 13.54 ;
  LAYER M1 ;
        RECT 15.344 13.488 15.376 13.56 ;
  LAYER M2 ;
        RECT 15.324 13.508 15.396 13.54 ;
  LAYER M1 ;
        RECT 12.624 10.716 12.656 10.788 ;
  LAYER M2 ;
        RECT 12.604 10.736 12.676 10.768 ;
  LAYER M1 ;
        RECT 12.624 10.584 12.656 10.752 ;
  LAYER M1 ;
        RECT 12.624 10.548 12.656 10.62 ;
  LAYER M2 ;
        RECT 12.604 10.568 12.676 10.6 ;
  LAYER M2 ;
        RECT 12.64 10.568 15.36 10.6 ;
  LAYER M1 ;
        RECT 15.344 10.548 15.376 10.62 ;
  LAYER M2 ;
        RECT 15.324 10.568 15.396 10.6 ;
  LAYER M1 ;
        RECT 12.624 7.776 12.656 7.848 ;
  LAYER M2 ;
        RECT 12.604 7.796 12.676 7.828 ;
  LAYER M1 ;
        RECT 12.624 7.644 12.656 7.812 ;
  LAYER M1 ;
        RECT 12.624 7.608 12.656 7.68 ;
  LAYER M2 ;
        RECT 12.604 7.628 12.676 7.66 ;
  LAYER M2 ;
        RECT 12.64 7.628 15.36 7.66 ;
  LAYER M1 ;
        RECT 15.344 7.608 15.376 7.68 ;
  LAYER M2 ;
        RECT 15.324 7.628 15.396 7.66 ;
  LAYER M1 ;
        RECT 12.624 4.836 12.656 4.908 ;
  LAYER M2 ;
        RECT 12.604 4.856 12.676 4.888 ;
  LAYER M1 ;
        RECT 12.624 4.704 12.656 4.872 ;
  LAYER M1 ;
        RECT 12.624 4.668 12.656 4.74 ;
  LAYER M2 ;
        RECT 12.604 4.688 12.676 4.72 ;
  LAYER M2 ;
        RECT 12.64 4.688 15.36 4.72 ;
  LAYER M1 ;
        RECT 15.344 4.668 15.376 4.74 ;
  LAYER M2 ;
        RECT 15.324 4.688 15.396 4.72 ;
  LAYER M1 ;
        RECT 12.624 1.896 12.656 1.968 ;
  LAYER M2 ;
        RECT 12.604 1.916 12.676 1.948 ;
  LAYER M1 ;
        RECT 12.624 1.764 12.656 1.932 ;
  LAYER M1 ;
        RECT 12.624 1.728 12.656 1.8 ;
  LAYER M2 ;
        RECT 12.604 1.748 12.676 1.78 ;
  LAYER M2 ;
        RECT 12.64 1.748 15.36 1.78 ;
  LAYER M1 ;
        RECT 15.344 1.728 15.376 1.8 ;
  LAYER M2 ;
        RECT 15.324 1.748 15.396 1.78 ;
  LAYER M1 ;
        RECT 15.344 1.056 15.376 1.128 ;
  LAYER M2 ;
        RECT 15.324 1.076 15.396 1.108 ;
  LAYER M1 ;
        RECT 15.344 1.092 15.376 1.596 ;
  LAYER M1 ;
        RECT 15.344 1.596 15.376 13.524 ;
  LAYER M2 ;
        RECT 0.96 1.076 15.36 1.108 ;
  LAYER M1 ;
        RECT 3.984 13.656 4.016 13.728 ;
  LAYER M2 ;
        RECT 3.964 13.676 4.036 13.708 ;
  LAYER M2 ;
        RECT 1.12 13.676 4 13.708 ;
  LAYER M1 ;
        RECT 1.104 13.656 1.136 13.728 ;
  LAYER M2 ;
        RECT 1.084 13.676 1.156 13.708 ;
  LAYER M1 ;
        RECT 3.984 1.896 4.016 1.968 ;
  LAYER M2 ;
        RECT 3.964 1.916 4.036 1.948 ;
  LAYER M2 ;
        RECT 1.12 1.916 4 1.948 ;
  LAYER M1 ;
        RECT 1.104 1.896 1.136 1.968 ;
  LAYER M2 ;
        RECT 1.084 1.916 1.156 1.948 ;
  LAYER M1 ;
        RECT 6.864 1.896 6.896 1.968 ;
  LAYER M2 ;
        RECT 6.844 1.916 6.916 1.948 ;
  LAYER M2 ;
        RECT 4 1.916 6.88 1.948 ;
  LAYER M1 ;
        RECT 3.984 1.896 4.016 1.968 ;
  LAYER M2 ;
        RECT 3.964 1.916 4.036 1.948 ;
  LAYER M1 ;
        RECT 9.744 1.896 9.776 1.968 ;
  LAYER M2 ;
        RECT 9.724 1.916 9.796 1.948 ;
  LAYER M2 ;
        RECT 6.88 1.916 9.76 1.948 ;
  LAYER M1 ;
        RECT 6.864 1.896 6.896 1.968 ;
  LAYER M2 ;
        RECT 6.844 1.916 6.916 1.948 ;
  LAYER M1 ;
        RECT 9.744 13.656 9.776 13.728 ;
  LAYER M2 ;
        RECT 9.724 13.676 9.796 13.708 ;
  LAYER M2 ;
        RECT 9.76 13.676 12.64 13.708 ;
  LAYER M1 ;
        RECT 12.624 13.656 12.656 13.728 ;
  LAYER M2 ;
        RECT 12.604 13.676 12.676 13.708 ;
  LAYER M1 ;
        RECT 6.864 13.656 6.896 13.728 ;
  LAYER M2 ;
        RECT 6.844 13.676 6.916 13.708 ;
  LAYER M2 ;
        RECT 6.88 13.676 9.76 13.708 ;
  LAYER M1 ;
        RECT 9.744 13.656 9.776 13.728 ;
  LAYER M2 ;
        RECT 9.724 13.676 9.796 13.708 ;
  LAYER M1 ;
        RECT 1.12 13.692 3.52 16.128 ;
  LAYER M2 ;
        RECT 1.12 13.692 3.52 16.128 ;
  LAYER M3 ;
        RECT 1.12 13.692 3.52 16.128 ;
  LAYER M1 ;
        RECT 1.12 10.752 3.52 13.188 ;
  LAYER M2 ;
        RECT 1.12 10.752 3.52 13.188 ;
  LAYER M3 ;
        RECT 1.12 10.752 3.52 13.188 ;
  LAYER M1 ;
        RECT 1.12 7.812 3.52 10.248 ;
  LAYER M2 ;
        RECT 1.12 7.812 3.52 10.248 ;
  LAYER M3 ;
        RECT 1.12 7.812 3.52 10.248 ;
  LAYER M1 ;
        RECT 1.12 4.872 3.52 7.308 ;
  LAYER M2 ;
        RECT 1.12 4.872 3.52 7.308 ;
  LAYER M3 ;
        RECT 1.12 4.872 3.52 7.308 ;
  LAYER M1 ;
        RECT 1.12 1.932 3.52 4.368 ;
  LAYER M2 ;
        RECT 1.12 1.932 3.52 4.368 ;
  LAYER M3 ;
        RECT 1.12 1.932 3.52 4.368 ;
  LAYER M1 ;
        RECT 4 13.692 6.4 16.128 ;
  LAYER M2 ;
        RECT 4 13.692 6.4 16.128 ;
  LAYER M3 ;
        RECT 4 13.692 6.4 16.128 ;
  LAYER M1 ;
        RECT 4 10.752 6.4 13.188 ;
  LAYER M2 ;
        RECT 4 10.752 6.4 13.188 ;
  LAYER M3 ;
        RECT 4 10.752 6.4 13.188 ;
  LAYER M1 ;
        RECT 4 7.812 6.4 10.248 ;
  LAYER M2 ;
        RECT 4 7.812 6.4 10.248 ;
  LAYER M3 ;
        RECT 4 7.812 6.4 10.248 ;
  LAYER M1 ;
        RECT 4 4.872 6.4 7.308 ;
  LAYER M2 ;
        RECT 4 4.872 6.4 7.308 ;
  LAYER M3 ;
        RECT 4 4.872 6.4 7.308 ;
  LAYER M1 ;
        RECT 4 1.932 6.4 4.368 ;
  LAYER M2 ;
        RECT 4 1.932 6.4 4.368 ;
  LAYER M3 ;
        RECT 4 1.932 6.4 4.368 ;
  LAYER M1 ;
        RECT 6.88 13.692 9.28 16.128 ;
  LAYER M2 ;
        RECT 6.88 13.692 9.28 16.128 ;
  LAYER M3 ;
        RECT 6.88 13.692 9.28 16.128 ;
  LAYER M1 ;
        RECT 6.88 10.752 9.28 13.188 ;
  LAYER M2 ;
        RECT 6.88 10.752 9.28 13.188 ;
  LAYER M3 ;
        RECT 6.88 10.752 9.28 13.188 ;
  LAYER M1 ;
        RECT 6.88 7.812 9.28 10.248 ;
  LAYER M2 ;
        RECT 6.88 7.812 9.28 10.248 ;
  LAYER M3 ;
        RECT 6.88 7.812 9.28 10.248 ;
  LAYER M1 ;
        RECT 6.88 4.872 9.28 7.308 ;
  LAYER M2 ;
        RECT 6.88 4.872 9.28 7.308 ;
  LAYER M3 ;
        RECT 6.88 4.872 9.28 7.308 ;
  LAYER M1 ;
        RECT 6.88 1.932 9.28 4.368 ;
  LAYER M2 ;
        RECT 6.88 1.932 9.28 4.368 ;
  LAYER M3 ;
        RECT 6.88 1.932 9.28 4.368 ;
  LAYER M1 ;
        RECT 9.76 13.692 12.16 16.128 ;
  LAYER M2 ;
        RECT 9.76 13.692 12.16 16.128 ;
  LAYER M3 ;
        RECT 9.76 13.692 12.16 16.128 ;
  LAYER M1 ;
        RECT 9.76 10.752 12.16 13.188 ;
  LAYER M2 ;
        RECT 9.76 10.752 12.16 13.188 ;
  LAYER M3 ;
        RECT 9.76 10.752 12.16 13.188 ;
  LAYER M1 ;
        RECT 9.76 7.812 12.16 10.248 ;
  LAYER M2 ;
        RECT 9.76 7.812 12.16 10.248 ;
  LAYER M3 ;
        RECT 9.76 7.812 12.16 10.248 ;
  LAYER M1 ;
        RECT 9.76 4.872 12.16 7.308 ;
  LAYER M2 ;
        RECT 9.76 4.872 12.16 7.308 ;
  LAYER M3 ;
        RECT 9.76 4.872 12.16 7.308 ;
  LAYER M1 ;
        RECT 9.76 1.932 12.16 4.368 ;
  LAYER M2 ;
        RECT 9.76 1.932 12.16 4.368 ;
  LAYER M3 ;
        RECT 9.76 1.932 12.16 4.368 ;
  LAYER M1 ;
        RECT 12.64 13.692 15.04 16.128 ;
  LAYER M2 ;
        RECT 12.64 13.692 15.04 16.128 ;
  LAYER M3 ;
        RECT 12.64 13.692 15.04 16.128 ;
  LAYER M1 ;
        RECT 12.64 10.752 15.04 13.188 ;
  LAYER M2 ;
        RECT 12.64 10.752 15.04 13.188 ;
  LAYER M3 ;
        RECT 12.64 10.752 15.04 13.188 ;
  LAYER M1 ;
        RECT 12.64 7.812 15.04 10.248 ;
  LAYER M2 ;
        RECT 12.64 7.812 15.04 10.248 ;
  LAYER M3 ;
        RECT 12.64 7.812 15.04 10.248 ;
  LAYER M1 ;
        RECT 12.64 4.872 15.04 7.308 ;
  LAYER M2 ;
        RECT 12.64 4.872 15.04 7.308 ;
  LAYER M3 ;
        RECT 12.64 4.872 15.04 7.308 ;
  LAYER M1 ;
        RECT 12.64 1.932 15.04 4.368 ;
  LAYER M2 ;
        RECT 12.64 1.932 15.04 4.368 ;
  LAYER M3 ;
        RECT 12.64 1.932 15.04 4.368 ;
  END 
END switched_capacitor_combination
