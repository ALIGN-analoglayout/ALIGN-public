module testcase_EA_placer ( 0, 1 ); 
input 0, 1;

CMC_PMOS_S_n12_X1_Y1 m1 ( .G(0) );
CMC_PMOS_S_n12_X1_Y1 m2 ( .G(1) );
CMC_PMOS_S_n12_X1_Y1 m2 ( .G(1) );

endmodule
