MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 2.5600 BY 1.7640 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
      LAYER M2 ;
        RECT 0.2040 0.9500 2.1960 0.9820 ;
    END
  END S
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4460 1.6360 0.4780 ;
      LAYER M2 ;
        RECT 0.2840 1.2860 2.2760 1.3180 ;
    END
  END GB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 2.2760 0.3940 ;
      LAYER M2 ;
        RECT 0.9240 1.2020 1.6360 1.2340 ;
    END
  END GA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
      LAYER M2 ;
        RECT 1.0040 1.0340 1.7160 1.0660 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
      LAYER M2 ;
        RECT 0.3640 1.1180 2.3560 1.1500 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 0.1620 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER M3 ;
      RECT 1.0200 0.1740 1.0600 0.2460 ;
    LAYER V2 ;
      RECT 1.0200 0.1940 1.0600 0.2260 ;
    LAYER V2 ;
      RECT 1.0200 0.1940 1.0600 0.2260 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER M3 ;
      RECT 1.3400 0.2580 1.3800 0.3300 ;
    LAYER V2 ;
      RECT 1.3400 0.2780 1.3800 0.3100 ;
    LAYER V2 ;
      RECT 1.3400 0.2780 1.3800 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER M3 ;
      RECT 1.1000 0.3420 1.1400 0.4140 ;
    LAYER V2 ;
      RECT 1.1000 0.3620 1.1400 0.3940 ;
    LAYER V2 ;
      RECT 1.1000 0.3620 1.1400 0.3940 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 2.2240 0.3620 2.2560 0.3940 ;
    LAYER M3 ;
      RECT 1.2600 0.4260 1.3000 0.4980 ;
    LAYER V2 ;
      RECT 1.2600 0.4460 1.3000 0.4780 ;
    LAYER V2 ;
      RECT 1.2600 0.4460 1.3000 0.4780 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
    LAYER M1 ;
      RECT 0.3040 0.9300 0.3360 1.5900 ;
    LAYER M1 ;
      RECT 2.2240 0.9300 2.2560 1.5900 ;
    LAYER M1 ;
      RECT 0.9440 0.9300 0.9760 1.5900 ;
    LAYER M1 ;
      RECT 1.5840 0.9300 1.6160 1.5900 ;
    LAYER M1 ;
      RECT 0.2240 0.9300 0.2560 1.5900 ;
    LAYER V0 ;
      RECT 0.2240 1.1180 0.2560 1.1500 ;
    LAYER V0 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V0 ;
      RECT 0.2240 1.3700 0.2560 1.4020 ;
    LAYER M1 ;
      RECT 2.1440 0.9300 2.1760 1.5900 ;
    LAYER V0 ;
      RECT 2.1440 1.1180 2.1760 1.1500 ;
    LAYER V0 ;
      RECT 2.1440 1.2440 2.1760 1.2760 ;
    LAYER V0 ;
      RECT 2.1440 1.3700 2.1760 1.4020 ;
    LAYER M1 ;
      RECT 0.8640 0.9300 0.8960 1.5900 ;
    LAYER V0 ;
      RECT 0.8640 1.1180 0.8960 1.1500 ;
    LAYER V0 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V0 ;
      RECT 0.8640 1.3700 0.8960 1.4020 ;
    LAYER M1 ;
      RECT 1.5040 0.9300 1.5360 1.5900 ;
    LAYER V0 ;
      RECT 1.5040 1.1180 1.5360 1.1500 ;
    LAYER V0 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V0 ;
      RECT 1.5040 1.3700 1.5360 1.4020 ;
    LAYER M1 ;
      RECT 0.3840 0.9300 0.4160 1.5900 ;
    LAYER V0 ;
      RECT 0.3840 1.1180 0.4160 1.1500 ;
    LAYER V0 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V0 ;
      RECT 0.3840 1.3700 0.4160 1.4020 ;
    LAYER M1 ;
      RECT 2.3040 0.9300 2.3360 1.5900 ;
    LAYER V0 ;
      RECT 2.3040 1.1180 2.3360 1.1500 ;
    LAYER V0 ;
      RECT 2.3040 1.2440 2.3360 1.2760 ;
    LAYER V0 ;
      RECT 2.3040 1.3700 2.3360 1.4020 ;
    LAYER M1 ;
      RECT 1.0240 0.9300 1.0560 1.5900 ;
    LAYER V0 ;
      RECT 1.0240 1.1180 1.0560 1.1500 ;
    LAYER V0 ;
      RECT 1.0240 1.2440 1.0560 1.2760 ;
    LAYER V0 ;
      RECT 1.0240 1.3700 1.0560 1.4020 ;
    LAYER M1 ;
      RECT 1.6640 0.9300 1.6960 1.5900 ;
    LAYER V0 ;
      RECT 1.6640 1.1180 1.6960 1.1500 ;
    LAYER V0 ;
      RECT 1.6640 1.2440 1.6960 1.2760 ;
    LAYER V0 ;
      RECT 1.6640 1.3700 1.6960 1.4020 ;
    LAYER M3 ;
      RECT 1.1800 0.0900 1.2200 1.0020 ;
    LAYER V2 ;
      RECT 1.1800 0.1100 1.2200 0.1420 ;
    LAYER V2 ;
      RECT 1.1800 0.9500 1.2200 0.9820 ;
    LAYER V1 ;
      RECT 0.2240 0.9500 0.2560 0.9820 ;
    LAYER V1 ;
      RECT 2.1440 0.9500 2.1760 0.9820 ;
    LAYER V1 ;
      RECT 0.8640 0.9500 0.8960 0.9820 ;
    LAYER V1 ;
      RECT 1.5040 0.9500 1.5360 0.9820 ;
    LAYER M3 ;
      RECT 1.0200 0.1740 1.0600 1.0860 ;
    LAYER V2 ;
      RECT 1.0200 0.1940 1.0600 0.2260 ;
    LAYER V2 ;
      RECT 1.0200 1.0340 1.0600 1.0660 ;
    LAYER V1 ;
      RECT 1.0240 1.0340 1.0560 1.0660 ;
    LAYER V1 ;
      RECT 1.6640 1.0340 1.6960 1.0660 ;
    LAYER M3 ;
      RECT 1.3400 0.2580 1.3800 1.1700 ;
    LAYER V2 ;
      RECT 1.3400 0.2780 1.3800 0.3100 ;
    LAYER V2 ;
      RECT 1.3400 1.1180 1.3800 1.1500 ;
    LAYER V1 ;
      RECT 0.3840 1.1180 0.4160 1.1500 ;
    LAYER V1 ;
      RECT 2.3040 1.1180 2.3360 1.1500 ;
    LAYER M3 ;
      RECT 1.1000 0.3420 1.1400 1.2540 ;
    LAYER V2 ;
      RECT 1.1000 0.3620 1.1400 0.3940 ;
    LAYER V2 ;
      RECT 1.1000 1.2020 1.1400 1.2340 ;
    LAYER V1 ;
      RECT 0.9440 1.2020 0.9760 1.2340 ;
    LAYER V1 ;
      RECT 1.5840 1.2020 1.6160 1.2340 ;
    LAYER M3 ;
      RECT 1.2600 0.4260 1.3000 1.3380 ;
    LAYER V2 ;
      RECT 1.2600 0.4460 1.3000 0.4780 ;
    LAYER V2 ;
      RECT 1.2600 1.2860 1.3000 1.3180 ;
    LAYER V1 ;
      RECT 0.3040 1.2860 0.3360 1.3180 ;
    LAYER V1 ;
      RECT 2.2240 1.2860 2.2560 1.3180 ;
  END
END test
