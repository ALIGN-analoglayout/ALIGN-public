MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 10.32 BY 26.208 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.808 25.752 3.84 25.824 ;
      LAYER M2 ;
        RECT 3.788 25.772 3.86 25.804 ;
      LAYER M1 ;
        RECT 7.104 25.752 7.136 25.824 ;
      LAYER M2 ;
        RECT 7.084 25.772 7.156 25.804 ;
      LAYER M2 ;
        RECT 3.824 25.772 7.12 25.804 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
      LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
      LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
      LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
      LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.968 25.92 4 25.992 ;
      LAYER M2 ;
        RECT 3.948 25.94 4.02 25.972 ;
      LAYER M1 ;
        RECT 7.264 25.92 7.296 25.992 ;
      LAYER M2 ;
        RECT 7.244 25.94 7.316 25.972 ;
      LAYER M2 ;
        RECT 3.984 25.94 7.28 25.972 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
      LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
      LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
      LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
      LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.496 13.404 6.528 13.476 ;
  LAYER M2 ;
        RECT 6.476 13.424 6.548 13.456 ;
  LAYER M2 ;
        RECT 3.376 13.424 6.512 13.456 ;
  LAYER M1 ;
        RECT 3.36 13.404 3.392 13.476 ;
  LAYER M2 ;
        RECT 3.34 13.424 3.412 13.456 ;
  LAYER M1 ;
        RECT 6.496 7.188 6.528 7.26 ;
  LAYER M2 ;
        RECT 6.476 7.208 6.548 7.24 ;
  LAYER M2 ;
        RECT 3.376 7.208 6.512 7.24 ;
  LAYER M1 ;
        RECT 3.36 7.188 3.392 7.26 ;
  LAYER M2 ;
        RECT 3.34 7.208 3.412 7.24 ;
  LAYER M1 ;
        RECT 6.496 16.512 6.528 16.584 ;
  LAYER M2 ;
        RECT 6.476 16.532 6.548 16.564 ;
  LAYER M2 ;
        RECT 3.376 16.532 6.512 16.564 ;
  LAYER M1 ;
        RECT 3.36 16.512 3.392 16.584 ;
  LAYER M2 ;
        RECT 3.34 16.532 3.412 16.564 ;
  LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
  LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
  LAYER M1 ;
        RECT 3.36 0.42 3.392 0.672 ;
  LAYER M1 ;
        RECT 3.36 0.672 3.392 16.548 ;
  LAYER M1 ;
        RECT 6.496 13.404 6.528 13.476 ;
  LAYER M2 ;
        RECT 6.476 13.424 6.548 13.456 ;
  LAYER M1 ;
        RECT 6.496 13.272 6.528 13.44 ;
  LAYER M1 ;
        RECT 6.496 13.236 6.528 13.308 ;
  LAYER M2 ;
        RECT 6.476 13.256 6.548 13.288 ;
  LAYER M2 ;
        RECT 6.512 13.256 6.672 13.288 ;
  LAYER M1 ;
        RECT 6.656 13.236 6.688 13.308 ;
  LAYER M2 ;
        RECT 6.636 13.256 6.708 13.288 ;
  LAYER M1 ;
        RECT 6.496 7.188 6.528 7.26 ;
  LAYER M2 ;
        RECT 6.476 7.208 6.548 7.24 ;
  LAYER M1 ;
        RECT 6.496 7.056 6.528 7.224 ;
  LAYER M1 ;
        RECT 6.496 7.02 6.528 7.092 ;
  LAYER M2 ;
        RECT 6.476 7.04 6.548 7.072 ;
  LAYER M2 ;
        RECT 6.512 7.04 6.672 7.072 ;
  LAYER M1 ;
        RECT 6.656 7.02 6.688 7.092 ;
  LAYER M2 ;
        RECT 6.636 7.04 6.708 7.072 ;
  LAYER M1 ;
        RECT 6.496 16.512 6.528 16.584 ;
  LAYER M2 ;
        RECT 6.476 16.532 6.548 16.564 ;
  LAYER M1 ;
        RECT 6.496 16.38 6.528 16.548 ;
  LAYER M1 ;
        RECT 6.496 16.344 6.528 16.416 ;
  LAYER M2 ;
        RECT 6.476 16.364 6.548 16.396 ;
  LAYER M2 ;
        RECT 6.512 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 16.416 ;
  LAYER M2 ;
        RECT 6.636 16.364 6.708 16.396 ;
  LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
  LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
  LAYER M1 ;
        RECT 6.656 0.42 6.688 0.672 ;
  LAYER M1 ;
        RECT 6.656 0.672 6.688 16.38 ;
  LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
  LAYER M1 ;
        RECT 6.496 10.296 6.528 10.368 ;
  LAYER M2 ;
        RECT 6.476 10.316 6.548 10.348 ;
  LAYER M2 ;
        RECT 3.536 10.316 6.512 10.348 ;
  LAYER M1 ;
        RECT 3.52 10.296 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.5 10.316 3.572 10.348 ;
  LAYER M1 ;
        RECT 6.496 4.08 6.528 4.152 ;
  LAYER M2 ;
        RECT 6.476 4.1 6.548 4.132 ;
  LAYER M2 ;
        RECT 3.536 4.1 6.512 4.132 ;
  LAYER M1 ;
        RECT 3.52 4.08 3.552 4.152 ;
  LAYER M2 ;
        RECT 3.5 4.1 3.572 4.132 ;
  LAYER M1 ;
        RECT 6.496 19.62 6.528 19.692 ;
  LAYER M2 ;
        RECT 6.476 19.64 6.548 19.672 ;
  LAYER M2 ;
        RECT 3.536 19.64 6.512 19.672 ;
  LAYER M1 ;
        RECT 3.52 19.62 3.552 19.692 ;
  LAYER M2 ;
        RECT 3.5 19.64 3.572 19.672 ;
  LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
  LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
  LAYER M1 ;
        RECT 3.52 0.252 3.552 0.672 ;
  LAYER M1 ;
        RECT 3.52 0.672 3.552 19.656 ;
  LAYER M1 ;
        RECT 6.496 10.296 6.528 10.368 ;
  LAYER M2 ;
        RECT 6.476 10.316 6.548 10.348 ;
  LAYER M1 ;
        RECT 6.496 10.164 6.528 10.332 ;
  LAYER M1 ;
        RECT 6.496 10.128 6.528 10.2 ;
  LAYER M2 ;
        RECT 6.476 10.148 6.548 10.18 ;
  LAYER M2 ;
        RECT 6.512 10.148 6.832 10.18 ;
  LAYER M1 ;
        RECT 6.816 10.128 6.848 10.2 ;
  LAYER M2 ;
        RECT 6.796 10.148 6.868 10.18 ;
  LAYER M1 ;
        RECT 6.496 4.08 6.528 4.152 ;
  LAYER M2 ;
        RECT 6.476 4.1 6.548 4.132 ;
  LAYER M1 ;
        RECT 6.496 3.948 6.528 4.116 ;
  LAYER M1 ;
        RECT 6.496 3.912 6.528 3.984 ;
  LAYER M2 ;
        RECT 6.476 3.932 6.548 3.964 ;
  LAYER M2 ;
        RECT 6.512 3.932 6.832 3.964 ;
  LAYER M1 ;
        RECT 6.816 3.912 6.848 3.984 ;
  LAYER M2 ;
        RECT 6.796 3.932 6.868 3.964 ;
  LAYER M1 ;
        RECT 6.496 19.62 6.528 19.692 ;
  LAYER M2 ;
        RECT 6.476 19.64 6.548 19.672 ;
  LAYER M1 ;
        RECT 6.496 19.488 6.528 19.656 ;
  LAYER M1 ;
        RECT 6.496 19.452 6.528 19.524 ;
  LAYER M2 ;
        RECT 6.476 19.472 6.548 19.504 ;
  LAYER M2 ;
        RECT 6.512 19.472 6.832 19.504 ;
  LAYER M1 ;
        RECT 6.816 19.452 6.848 19.524 ;
  LAYER M2 ;
        RECT 6.796 19.472 6.868 19.504 ;
  LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
  LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
  LAYER M1 ;
        RECT 6.816 0.252 6.848 0.672 ;
  LAYER M1 ;
        RECT 6.816 0.672 6.848 19.488 ;
  LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
  LAYER M1 ;
        RECT 3.2 0.972 3.232 1.044 ;
  LAYER M2 ;
        RECT 3.18 0.992 3.252 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 3.216 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 3.2 4.08 3.232 4.152 ;
  LAYER M2 ;
        RECT 3.18 4.1 3.252 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 3.216 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 3.2 7.188 3.232 7.26 ;
  LAYER M2 ;
        RECT 3.18 7.208 3.252 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 3.216 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 3.2 10.296 3.232 10.368 ;
  LAYER M2 ;
        RECT 3.18 10.316 3.252 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 3.216 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 3.2 13.404 3.232 13.476 ;
  LAYER M2 ;
        RECT 3.18 13.424 3.252 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 3.216 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 3.2 16.512 3.232 16.584 ;
  LAYER M2 ;
        RECT 3.18 16.532 3.252 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 3.216 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 3.2 19.62 3.232 19.692 ;
  LAYER M2 ;
        RECT 3.18 19.64 3.252 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 3.216 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 3.2 22.728 3.232 22.8 ;
  LAYER M2 ;
        RECT 3.18 22.748 3.252 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 3.216 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 22.764 ;
  LAYER M1 ;
        RECT 9.792 0.972 9.824 1.044 ;
  LAYER M2 ;
        RECT 9.772 0.992 9.844 1.024 ;
  LAYER M1 ;
        RECT 9.792 0.84 9.824 1.008 ;
  LAYER M1 ;
        RECT 9.792 0.804 9.824 0.876 ;
  LAYER M2 ;
        RECT 9.772 0.824 9.844 0.856 ;
  LAYER M2 ;
        RECT 9.808 0.824 9.968 0.856 ;
  LAYER M1 ;
        RECT 9.952 0.804 9.984 0.876 ;
  LAYER M2 ;
        RECT 9.932 0.824 10.004 0.856 ;
  LAYER M1 ;
        RECT 9.792 4.08 9.824 4.152 ;
  LAYER M2 ;
        RECT 9.772 4.1 9.844 4.132 ;
  LAYER M1 ;
        RECT 9.792 3.948 9.824 4.116 ;
  LAYER M1 ;
        RECT 9.792 3.912 9.824 3.984 ;
  LAYER M2 ;
        RECT 9.772 3.932 9.844 3.964 ;
  LAYER M2 ;
        RECT 9.808 3.932 9.968 3.964 ;
  LAYER M1 ;
        RECT 9.952 3.912 9.984 3.984 ;
  LAYER M2 ;
        RECT 9.932 3.932 10.004 3.964 ;
  LAYER M1 ;
        RECT 9.792 7.188 9.824 7.26 ;
  LAYER M2 ;
        RECT 9.772 7.208 9.844 7.24 ;
  LAYER M1 ;
        RECT 9.792 7.056 9.824 7.224 ;
  LAYER M1 ;
        RECT 9.792 7.02 9.824 7.092 ;
  LAYER M2 ;
        RECT 9.772 7.04 9.844 7.072 ;
  LAYER M2 ;
        RECT 9.808 7.04 9.968 7.072 ;
  LAYER M1 ;
        RECT 9.952 7.02 9.984 7.092 ;
  LAYER M2 ;
        RECT 9.932 7.04 10.004 7.072 ;
  LAYER M1 ;
        RECT 9.792 10.296 9.824 10.368 ;
  LAYER M2 ;
        RECT 9.772 10.316 9.844 10.348 ;
  LAYER M1 ;
        RECT 9.792 10.164 9.824 10.332 ;
  LAYER M1 ;
        RECT 9.792 10.128 9.824 10.2 ;
  LAYER M2 ;
        RECT 9.772 10.148 9.844 10.18 ;
  LAYER M2 ;
        RECT 9.808 10.148 9.968 10.18 ;
  LAYER M1 ;
        RECT 9.952 10.128 9.984 10.2 ;
  LAYER M2 ;
        RECT 9.932 10.148 10.004 10.18 ;
  LAYER M1 ;
        RECT 9.792 13.404 9.824 13.476 ;
  LAYER M2 ;
        RECT 9.772 13.424 9.844 13.456 ;
  LAYER M1 ;
        RECT 9.792 13.272 9.824 13.44 ;
  LAYER M1 ;
        RECT 9.792 13.236 9.824 13.308 ;
  LAYER M2 ;
        RECT 9.772 13.256 9.844 13.288 ;
  LAYER M2 ;
        RECT 9.808 13.256 9.968 13.288 ;
  LAYER M1 ;
        RECT 9.952 13.236 9.984 13.308 ;
  LAYER M2 ;
        RECT 9.932 13.256 10.004 13.288 ;
  LAYER M1 ;
        RECT 9.792 16.512 9.824 16.584 ;
  LAYER M2 ;
        RECT 9.772 16.532 9.844 16.564 ;
  LAYER M1 ;
        RECT 9.792 16.38 9.824 16.548 ;
  LAYER M1 ;
        RECT 9.792 16.344 9.824 16.416 ;
  LAYER M2 ;
        RECT 9.772 16.364 9.844 16.396 ;
  LAYER M2 ;
        RECT 9.808 16.364 9.968 16.396 ;
  LAYER M1 ;
        RECT 9.952 16.344 9.984 16.416 ;
  LAYER M2 ;
        RECT 9.932 16.364 10.004 16.396 ;
  LAYER M1 ;
        RECT 9.792 19.62 9.824 19.692 ;
  LAYER M2 ;
        RECT 9.772 19.64 9.844 19.672 ;
  LAYER M1 ;
        RECT 9.792 19.488 9.824 19.656 ;
  LAYER M1 ;
        RECT 9.792 19.452 9.824 19.524 ;
  LAYER M2 ;
        RECT 9.772 19.472 9.844 19.504 ;
  LAYER M2 ;
        RECT 9.808 19.472 9.968 19.504 ;
  LAYER M1 ;
        RECT 9.952 19.452 9.984 19.524 ;
  LAYER M2 ;
        RECT 9.932 19.472 10.004 19.504 ;
  LAYER M1 ;
        RECT 9.792 22.728 9.824 22.8 ;
  LAYER M2 ;
        RECT 9.772 22.748 9.844 22.78 ;
  LAYER M1 ;
        RECT 9.792 22.596 9.824 22.764 ;
  LAYER M1 ;
        RECT 9.792 22.56 9.824 22.632 ;
  LAYER M2 ;
        RECT 9.772 22.58 9.844 22.612 ;
  LAYER M2 ;
        RECT 9.808 22.58 9.968 22.612 ;
  LAYER M1 ;
        RECT 9.952 22.56 9.984 22.632 ;
  LAYER M2 ;
        RECT 9.932 22.58 10.004 22.612 ;
  LAYER M1 ;
        RECT 9.952 0.048 9.984 0.12 ;
  LAYER M2 ;
        RECT 9.932 0.068 10.004 0.1 ;
  LAYER M1 ;
        RECT 9.952 0.084 9.984 0.672 ;
  LAYER M1 ;
        RECT 9.952 0.672 9.984 22.596 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.968 0.1 ;
  LAYER M1 ;
        RECT 6.496 0.972 6.528 1.044 ;
  LAYER M2 ;
        RECT 6.476 0.992 6.548 1.024 ;
  LAYER M2 ;
        RECT 3.216 0.992 6.512 1.024 ;
  LAYER M1 ;
        RECT 3.2 0.972 3.232 1.044 ;
  LAYER M2 ;
        RECT 3.18 0.992 3.252 1.024 ;
  LAYER M1 ;
        RECT 6.496 22.728 6.528 22.8 ;
  LAYER M2 ;
        RECT 6.476 22.748 6.548 22.78 ;
  LAYER M2 ;
        RECT 3.216 22.748 6.512 22.78 ;
  LAYER M1 ;
        RECT 3.2 22.728 3.232 22.8 ;
  LAYER M2 ;
        RECT 3.18 22.748 3.252 22.78 ;
  LAYER M1 ;
        RECT 4.128 15.84 4.16 15.912 ;
  LAYER M2 ;
        RECT 4.108 15.86 4.18 15.892 ;
  LAYER M2 ;
        RECT 3.824 15.86 4.144 15.892 ;
  LAYER M1 ;
        RECT 3.808 15.84 3.84 15.912 ;
  LAYER M2 ;
        RECT 3.788 15.86 3.86 15.892 ;
  LAYER M1 ;
        RECT 4.128 9.624 4.16 9.696 ;
  LAYER M2 ;
        RECT 4.108 9.644 4.18 9.676 ;
  LAYER M2 ;
        RECT 3.824 9.644 4.144 9.676 ;
  LAYER M1 ;
        RECT 3.808 9.624 3.84 9.696 ;
  LAYER M2 ;
        RECT 3.788 9.644 3.86 9.676 ;
  LAYER M1 ;
        RECT 4.128 18.948 4.16 19.02 ;
  LAYER M2 ;
        RECT 4.108 18.968 4.18 19 ;
  LAYER M2 ;
        RECT 3.824 18.968 4.144 19 ;
  LAYER M1 ;
        RECT 3.808 18.948 3.84 19.02 ;
  LAYER M2 ;
        RECT 3.788 18.968 3.86 19 ;
  LAYER M1 ;
        RECT 3.808 25.752 3.84 25.824 ;
  LAYER M2 ;
        RECT 3.788 25.772 3.86 25.804 ;
  LAYER M1 ;
        RECT 3.808 25.536 3.84 25.788 ;
  LAYER M1 ;
        RECT 3.808 9.66 3.84 25.536 ;
  LAYER M1 ;
        RECT 4.128 15.84 4.16 15.912 ;
  LAYER M2 ;
        RECT 4.108 15.86 4.18 15.892 ;
  LAYER M1 ;
        RECT 4.128 15.876 4.16 16.044 ;
  LAYER M1 ;
        RECT 4.128 16.008 4.16 16.08 ;
  LAYER M2 ;
        RECT 4.108 16.028 4.18 16.06 ;
  LAYER M2 ;
        RECT 4.144 16.028 7.12 16.06 ;
  LAYER M1 ;
        RECT 7.104 16.008 7.136 16.08 ;
  LAYER M2 ;
        RECT 7.084 16.028 7.156 16.06 ;
  LAYER M1 ;
        RECT 4.128 9.624 4.16 9.696 ;
  LAYER M2 ;
        RECT 4.108 9.644 4.18 9.676 ;
  LAYER M1 ;
        RECT 4.128 9.66 4.16 9.828 ;
  LAYER M1 ;
        RECT 4.128 9.792 4.16 9.864 ;
  LAYER M2 ;
        RECT 4.108 9.812 4.18 9.844 ;
  LAYER M2 ;
        RECT 4.144 9.812 7.12 9.844 ;
  LAYER M1 ;
        RECT 7.104 9.792 7.136 9.864 ;
  LAYER M2 ;
        RECT 7.084 9.812 7.156 9.844 ;
  LAYER M1 ;
        RECT 4.128 18.948 4.16 19.02 ;
  LAYER M2 ;
        RECT 4.108 18.968 4.18 19 ;
  LAYER M1 ;
        RECT 4.128 18.984 4.16 19.152 ;
  LAYER M1 ;
        RECT 4.128 19.116 4.16 19.188 ;
  LAYER M2 ;
        RECT 4.108 19.136 4.18 19.168 ;
  LAYER M2 ;
        RECT 4.144 19.136 7.12 19.168 ;
  LAYER M1 ;
        RECT 7.104 19.116 7.136 19.188 ;
  LAYER M2 ;
        RECT 7.084 19.136 7.156 19.168 ;
  LAYER M1 ;
        RECT 7.104 25.752 7.136 25.824 ;
  LAYER M2 ;
        RECT 7.084 25.772 7.156 25.804 ;
  LAYER M1 ;
        RECT 7.104 25.536 7.136 25.788 ;
  LAYER M1 ;
        RECT 7.104 9.828 7.136 25.536 ;
  LAYER M2 ;
        RECT 3.824 25.772 7.12 25.804 ;
  LAYER M1 ;
        RECT 4.128 12.732 4.16 12.804 ;
  LAYER M2 ;
        RECT 4.108 12.752 4.18 12.784 ;
  LAYER M2 ;
        RECT 3.984 12.752 4.144 12.784 ;
  LAYER M1 ;
        RECT 3.968 12.732 4 12.804 ;
  LAYER M2 ;
        RECT 3.948 12.752 4.02 12.784 ;
  LAYER M1 ;
        RECT 4.128 6.516 4.16 6.588 ;
  LAYER M2 ;
        RECT 4.108 6.536 4.18 6.568 ;
  LAYER M2 ;
        RECT 3.984 6.536 4.144 6.568 ;
  LAYER M1 ;
        RECT 3.968 6.516 4 6.588 ;
  LAYER M2 ;
        RECT 3.948 6.536 4.02 6.568 ;
  LAYER M1 ;
        RECT 4.128 22.056 4.16 22.128 ;
  LAYER M2 ;
        RECT 4.108 22.076 4.18 22.108 ;
  LAYER M2 ;
        RECT 3.984 22.076 4.144 22.108 ;
  LAYER M1 ;
        RECT 3.968 22.056 4 22.128 ;
  LAYER M2 ;
        RECT 3.948 22.076 4.02 22.108 ;
  LAYER M1 ;
        RECT 3.968 25.92 4 25.992 ;
  LAYER M2 ;
        RECT 3.948 25.94 4.02 25.972 ;
  LAYER M1 ;
        RECT 3.968 25.536 4 25.956 ;
  LAYER M1 ;
        RECT 3.968 6.552 4 25.536 ;
  LAYER M1 ;
        RECT 4.128 12.732 4.16 12.804 ;
  LAYER M2 ;
        RECT 4.108 12.752 4.18 12.784 ;
  LAYER M1 ;
        RECT 4.128 12.768 4.16 12.936 ;
  LAYER M1 ;
        RECT 4.128 12.9 4.16 12.972 ;
  LAYER M2 ;
        RECT 4.108 12.92 4.18 12.952 ;
  LAYER M2 ;
        RECT 4.144 12.92 7.28 12.952 ;
  LAYER M1 ;
        RECT 7.264 12.9 7.296 12.972 ;
  LAYER M2 ;
        RECT 7.244 12.92 7.316 12.952 ;
  LAYER M1 ;
        RECT 4.128 6.516 4.16 6.588 ;
  LAYER M2 ;
        RECT 4.108 6.536 4.18 6.568 ;
  LAYER M1 ;
        RECT 4.128 6.552 4.16 6.72 ;
  LAYER M1 ;
        RECT 4.128 6.684 4.16 6.756 ;
  LAYER M2 ;
        RECT 4.108 6.704 4.18 6.736 ;
  LAYER M2 ;
        RECT 4.144 6.704 7.28 6.736 ;
  LAYER M1 ;
        RECT 7.264 6.684 7.296 6.756 ;
  LAYER M2 ;
        RECT 7.244 6.704 7.316 6.736 ;
  LAYER M1 ;
        RECT 4.128 22.056 4.16 22.128 ;
  LAYER M2 ;
        RECT 4.108 22.076 4.18 22.108 ;
  LAYER M1 ;
        RECT 4.128 22.092 4.16 22.26 ;
  LAYER M1 ;
        RECT 4.128 22.224 4.16 22.296 ;
  LAYER M2 ;
        RECT 4.108 22.244 4.18 22.276 ;
  LAYER M2 ;
        RECT 4.144 22.244 7.28 22.276 ;
  LAYER M1 ;
        RECT 7.264 22.224 7.296 22.296 ;
  LAYER M2 ;
        RECT 7.244 22.244 7.316 22.276 ;
  LAYER M1 ;
        RECT 7.264 25.92 7.296 25.992 ;
  LAYER M2 ;
        RECT 7.244 25.94 7.316 25.972 ;
  LAYER M1 ;
        RECT 7.264 25.536 7.296 25.956 ;
  LAYER M1 ;
        RECT 7.264 6.72 7.296 25.536 ;
  LAYER M2 ;
        RECT 3.984 25.94 7.28 25.972 ;
  LAYER M1 ;
        RECT 0.832 3.408 0.864 3.48 ;
  LAYER M2 ;
        RECT 0.812 3.428 0.884 3.46 ;
  LAYER M2 ;
        RECT 0.368 3.428 0.848 3.46 ;
  LAYER M1 ;
        RECT 0.352 3.408 0.384 3.48 ;
  LAYER M2 ;
        RECT 0.332 3.428 0.404 3.46 ;
  LAYER M1 ;
        RECT 0.832 6.516 0.864 6.588 ;
  LAYER M2 ;
        RECT 0.812 6.536 0.884 6.568 ;
  LAYER M2 ;
        RECT 0.368 6.536 0.848 6.568 ;
  LAYER M1 ;
        RECT 0.352 6.516 0.384 6.588 ;
  LAYER M2 ;
        RECT 0.332 6.536 0.404 6.568 ;
  LAYER M1 ;
        RECT 0.832 9.624 0.864 9.696 ;
  LAYER M2 ;
        RECT 0.812 9.644 0.884 9.676 ;
  LAYER M2 ;
        RECT 0.368 9.644 0.848 9.676 ;
  LAYER M1 ;
        RECT 0.352 9.624 0.384 9.696 ;
  LAYER M2 ;
        RECT 0.332 9.644 0.404 9.676 ;
  LAYER M1 ;
        RECT 0.832 12.732 0.864 12.804 ;
  LAYER M2 ;
        RECT 0.812 12.752 0.884 12.784 ;
  LAYER M2 ;
        RECT 0.368 12.752 0.848 12.784 ;
  LAYER M1 ;
        RECT 0.352 12.732 0.384 12.804 ;
  LAYER M2 ;
        RECT 0.332 12.752 0.404 12.784 ;
  LAYER M1 ;
        RECT 0.832 15.84 0.864 15.912 ;
  LAYER M2 ;
        RECT 0.812 15.86 0.884 15.892 ;
  LAYER M2 ;
        RECT 0.368 15.86 0.848 15.892 ;
  LAYER M1 ;
        RECT 0.352 15.84 0.384 15.912 ;
  LAYER M2 ;
        RECT 0.332 15.86 0.404 15.892 ;
  LAYER M1 ;
        RECT 0.832 18.948 0.864 19.02 ;
  LAYER M2 ;
        RECT 0.812 18.968 0.884 19 ;
  LAYER M2 ;
        RECT 0.368 18.968 0.848 19 ;
  LAYER M1 ;
        RECT 0.352 18.948 0.384 19.02 ;
  LAYER M2 ;
        RECT 0.332 18.968 0.404 19 ;
  LAYER M1 ;
        RECT 0.832 22.056 0.864 22.128 ;
  LAYER M2 ;
        RECT 0.812 22.076 0.884 22.108 ;
  LAYER M2 ;
        RECT 0.368 22.076 0.848 22.108 ;
  LAYER M1 ;
        RECT 0.352 22.056 0.384 22.128 ;
  LAYER M2 ;
        RECT 0.332 22.076 0.404 22.108 ;
  LAYER M1 ;
        RECT 0.832 25.164 0.864 25.236 ;
  LAYER M2 ;
        RECT 0.812 25.184 0.884 25.216 ;
  LAYER M2 ;
        RECT 0.368 25.184 0.848 25.216 ;
  LAYER M1 ;
        RECT 0.352 25.164 0.384 25.236 ;
  LAYER M2 ;
        RECT 0.332 25.184 0.404 25.216 ;
  LAYER M1 ;
        RECT 0.352 26.088 0.384 26.16 ;
  LAYER M2 ;
        RECT 0.332 26.108 0.404 26.14 ;
  LAYER M1 ;
        RECT 0.352 25.536 0.384 26.124 ;
  LAYER M1 ;
        RECT 0.352 3.444 0.384 25.536 ;
  LAYER M1 ;
        RECT 7.424 3.408 7.456 3.48 ;
  LAYER M2 ;
        RECT 7.404 3.428 7.476 3.46 ;
  LAYER M1 ;
        RECT 7.424 3.444 7.456 3.612 ;
  LAYER M1 ;
        RECT 7.424 3.576 7.456 3.648 ;
  LAYER M2 ;
        RECT 7.404 3.596 7.476 3.628 ;
  LAYER M2 ;
        RECT 7.44 3.596 10.256 3.628 ;
  LAYER M1 ;
        RECT 10.24 3.576 10.272 3.648 ;
  LAYER M2 ;
        RECT 10.22 3.596 10.292 3.628 ;
  LAYER M1 ;
        RECT 7.424 6.516 7.456 6.588 ;
  LAYER M2 ;
        RECT 7.404 6.536 7.476 6.568 ;
  LAYER M1 ;
        RECT 7.424 6.552 7.456 6.72 ;
  LAYER M1 ;
        RECT 7.424 6.684 7.456 6.756 ;
  LAYER M2 ;
        RECT 7.404 6.704 7.476 6.736 ;
  LAYER M2 ;
        RECT 7.44 6.704 10.256 6.736 ;
  LAYER M1 ;
        RECT 10.24 6.684 10.272 6.756 ;
  LAYER M2 ;
        RECT 10.22 6.704 10.292 6.736 ;
  LAYER M1 ;
        RECT 7.424 9.624 7.456 9.696 ;
  LAYER M2 ;
        RECT 7.404 9.644 7.476 9.676 ;
  LAYER M1 ;
        RECT 7.424 9.66 7.456 9.828 ;
  LAYER M1 ;
        RECT 7.424 9.792 7.456 9.864 ;
  LAYER M2 ;
        RECT 7.404 9.812 7.476 9.844 ;
  LAYER M2 ;
        RECT 7.44 9.812 10.256 9.844 ;
  LAYER M1 ;
        RECT 10.24 9.792 10.272 9.864 ;
  LAYER M2 ;
        RECT 10.22 9.812 10.292 9.844 ;
  LAYER M1 ;
        RECT 7.424 12.732 7.456 12.804 ;
  LAYER M2 ;
        RECT 7.404 12.752 7.476 12.784 ;
  LAYER M1 ;
        RECT 7.424 12.768 7.456 12.936 ;
  LAYER M1 ;
        RECT 7.424 12.9 7.456 12.972 ;
  LAYER M2 ;
        RECT 7.404 12.92 7.476 12.952 ;
  LAYER M2 ;
        RECT 7.44 12.92 10.256 12.952 ;
  LAYER M1 ;
        RECT 10.24 12.9 10.272 12.972 ;
  LAYER M2 ;
        RECT 10.22 12.92 10.292 12.952 ;
  LAYER M1 ;
        RECT 7.424 15.84 7.456 15.912 ;
  LAYER M2 ;
        RECT 7.404 15.86 7.476 15.892 ;
  LAYER M1 ;
        RECT 7.424 15.876 7.456 16.044 ;
  LAYER M1 ;
        RECT 7.424 16.008 7.456 16.08 ;
  LAYER M2 ;
        RECT 7.404 16.028 7.476 16.06 ;
  LAYER M2 ;
        RECT 7.44 16.028 10.256 16.06 ;
  LAYER M1 ;
        RECT 10.24 16.008 10.272 16.08 ;
  LAYER M2 ;
        RECT 10.22 16.028 10.292 16.06 ;
  LAYER M1 ;
        RECT 7.424 18.948 7.456 19.02 ;
  LAYER M2 ;
        RECT 7.404 18.968 7.476 19 ;
  LAYER M1 ;
        RECT 7.424 18.984 7.456 19.152 ;
  LAYER M1 ;
        RECT 7.424 19.116 7.456 19.188 ;
  LAYER M2 ;
        RECT 7.404 19.136 7.476 19.168 ;
  LAYER M2 ;
        RECT 7.44 19.136 10.256 19.168 ;
  LAYER M1 ;
        RECT 10.24 19.116 10.272 19.188 ;
  LAYER M2 ;
        RECT 10.22 19.136 10.292 19.168 ;
  LAYER M1 ;
        RECT 7.424 22.056 7.456 22.128 ;
  LAYER M2 ;
        RECT 7.404 22.076 7.476 22.108 ;
  LAYER M1 ;
        RECT 7.424 22.092 7.456 22.26 ;
  LAYER M1 ;
        RECT 7.424 22.224 7.456 22.296 ;
  LAYER M2 ;
        RECT 7.404 22.244 7.476 22.276 ;
  LAYER M2 ;
        RECT 7.44 22.244 10.256 22.276 ;
  LAYER M1 ;
        RECT 10.24 22.224 10.272 22.296 ;
  LAYER M2 ;
        RECT 10.22 22.244 10.292 22.276 ;
  LAYER M1 ;
        RECT 7.424 25.164 7.456 25.236 ;
  LAYER M2 ;
        RECT 7.404 25.184 7.476 25.216 ;
  LAYER M1 ;
        RECT 7.424 25.2 7.456 25.368 ;
  LAYER M1 ;
        RECT 7.424 25.332 7.456 25.404 ;
  LAYER M2 ;
        RECT 7.404 25.352 7.476 25.384 ;
  LAYER M2 ;
        RECT 7.44 25.352 10.256 25.384 ;
  LAYER M1 ;
        RECT 10.24 25.332 10.272 25.404 ;
  LAYER M2 ;
        RECT 10.22 25.352 10.292 25.384 ;
  LAYER M1 ;
        RECT 10.24 26.088 10.272 26.16 ;
  LAYER M2 ;
        RECT 10.22 26.108 10.292 26.14 ;
  LAYER M1 ;
        RECT 10.24 25.536 10.272 26.124 ;
  LAYER M1 ;
        RECT 10.24 3.612 10.272 25.536 ;
  LAYER M2 ;
        RECT 0.368 26.108 10.256 26.14 ;
  LAYER M1 ;
        RECT 4.128 3.408 4.16 3.48 ;
  LAYER M2 ;
        RECT 4.108 3.428 4.18 3.46 ;
  LAYER M2 ;
        RECT 0.848 3.428 4.144 3.46 ;
  LAYER M1 ;
        RECT 0.832 3.408 0.864 3.48 ;
  LAYER M2 ;
        RECT 0.812 3.428 0.884 3.46 ;
  LAYER M1 ;
        RECT 4.128 25.164 4.16 25.236 ;
  LAYER M2 ;
        RECT 4.108 25.184 4.18 25.216 ;
  LAYER M2 ;
        RECT 0.848 25.184 4.144 25.216 ;
  LAYER M1 ;
        RECT 0.832 25.164 0.864 25.236 ;
  LAYER M2 ;
        RECT 0.812 25.184 0.884 25.216 ;
  LAYER M1 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M3 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M2 ;
        RECT 0.784 0.924 3.28 3.528 ;
  LAYER M1 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M3 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M2 ;
        RECT 0.784 4.032 3.28 6.636 ;
  LAYER M1 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M3 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M2 ;
        RECT 0.784 7.14 3.28 9.744 ;
  LAYER M1 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M3 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M2 ;
        RECT 0.784 10.248 3.28 12.852 ;
  LAYER M1 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M3 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M2 ;
        RECT 0.784 13.356 3.28 15.96 ;
  LAYER M1 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M3 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M2 ;
        RECT 0.784 16.464 3.28 19.068 ;
  LAYER M1 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M3 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M2 ;
        RECT 0.784 19.572 3.28 22.176 ;
  LAYER M1 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M3 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M2 ;
        RECT 0.784 22.68 3.28 25.284 ;
  LAYER M1 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M3 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M2 ;
        RECT 4.08 0.924 6.576 3.528 ;
  LAYER M1 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M3 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M2 ;
        RECT 4.08 4.032 6.576 6.636 ;
  LAYER M1 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M3 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M2 ;
        RECT 4.08 7.14 6.576 9.744 ;
  LAYER M1 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M3 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M2 ;
        RECT 4.08 10.248 6.576 12.852 ;
  LAYER M1 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M3 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M2 ;
        RECT 4.08 13.356 6.576 15.96 ;
  LAYER M1 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M3 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M2 ;
        RECT 4.08 16.464 6.576 19.068 ;
  LAYER M1 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M3 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M2 ;
        RECT 4.08 19.572 6.576 22.176 ;
  LAYER M1 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M3 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M2 ;
        RECT 4.08 22.68 6.576 25.284 ;
  LAYER M1 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M3 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M2 ;
        RECT 7.376 0.924 9.872 3.528 ;
  LAYER M1 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M3 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M2 ;
        RECT 7.376 4.032 9.872 6.636 ;
  LAYER M1 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M3 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M2 ;
        RECT 7.376 7.14 9.872 9.744 ;
  LAYER M1 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M3 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M2 ;
        RECT 7.376 10.248 9.872 12.852 ;
  LAYER M1 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M3 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M2 ;
        RECT 7.376 13.356 9.872 15.96 ;
  LAYER M1 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M3 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M2 ;
        RECT 7.376 16.464 9.872 19.068 ;
  LAYER M1 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M3 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M2 ;
        RECT 7.376 19.572 9.872 22.176 ;
  LAYER M1 ;
        RECT 7.376 22.68 9.872 25.284 ;
  LAYER M3 ;
        RECT 7.376 22.68 9.872 25.284 ;
  LAYER M2 ;
        RECT 7.376 22.68 9.872 25.284 ;
  END 
END Cap_30fF_Cap_30fF
