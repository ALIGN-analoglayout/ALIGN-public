MACRO __json_dp_nmos_cand
  ORIGIN 0 0 ;
  FOREIGN __json_dp_nmos_cand 0 0 ;
  SIZE 256000.0000 BY 168000.0000 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20400.0000 6800.0000 235600.0000 10000.0000 ;
      LAYER M2 ;
        RECT 20400.0000 90800.0000 235600.0000 94000.0000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36400.0000 15200.0000 219600.0000 18400.0000 ;
      LAYER M2 ;
        RECT 100400.0000 99200.0000 155600.0000 102400.0000 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100400.0000 23600.0000 155600.0000 26800.0000 ;
      LAYER M2 ;
        RECT 36400.0000 107600.0000 219600.0000 110800.0000 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28400.0000 32000.0000 227600.0000 35200.0000 ;
      LAYER M2 ;
        RECT 92400.0000 116000.0000 163600.0000 119200.0000 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92400.0000 40400.0000 163600.0000 43600.0000 ;
      LAYER M2 ;
        RECT 28400.0000 124400.0000 227600.0000 127600.0000 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 30400.0000 4800.0000 33600.0000 70800.0000 ;
    LAYER M1 ;
      RECT 222400.0000 4800.0000 225600.0000 70800.0000 ;
    LAYER M1 ;
      RECT 94400.0000 4800.0000 97600.0000 70800.0000 ;
    LAYER M1 ;
      RECT 158400.0000 4800.0000 161600.0000 70800.0000 ;
    LAYER M1 ;
      RECT 22400.0000 4800.0000 25600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 22400.0000 23600.0000 25600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 22400.0000 36200.0000 25600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 22400.0000 48800.0000 25600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 230400.0000 4800.0000 233600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 230400.0000 23600.0000 233600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 230400.0000 36200.0000 233600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 230400.0000 48800.0000 233600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 86400.0000 4800.0000 89600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 86400.0000 23600.0000 89600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 86400.0000 36200.0000 89600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 86400.0000 48800.0000 89600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 166400.0000 4800.0000 169600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 166400.0000 23600.0000 169600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 166400.0000 36200.0000 169600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 166400.0000 48800.0000 169600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 38400.0000 4800.0000 41600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 38400.0000 23600.0000 41600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 38400.0000 36200.0000 41600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 38400.0000 48800.0000 41600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 214400.0000 4800.0000 217600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 214400.0000 23600.0000 217600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 214400.0000 36200.0000 217600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 214400.0000 48800.0000 217600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 102400.0000 4800.0000 105600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 102400.0000 23600.0000 105600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 102400.0000 36200.0000 105600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 102400.0000 48800.0000 105600.0000 52000.0000 ;
    LAYER M1 ;
      RECT 150400.0000 4800.0000 153600.0000 70800.0000 ;
    LAYER V0 ;
      RECT 150400.0000 23600.0000 153600.0000 26800.0000 ;
    LAYER V0 ;
      RECT 150400.0000 36200.0000 153600.0000 39400.0000 ;
    LAYER V0 ;
      RECT 150400.0000 48800.0000 153600.0000 52000.0000 ;
    LAYER M3 ;
      RECT 126000.0000 4800.0000 130000.0000 12000.0000 ;
    LAYER V2 ;
      RECT 126000.0000 6800.0000 130000.0000 10000.0000 ;
    LAYER V2 ;
      RECT 126000.0000 6800.0000 130000.0000 10000.0000 ;
    LAYER V1 ;
      RECT 22400.0000 6800.0000 25600.0000 10000.0000 ;
    LAYER V1 ;
      RECT 230400.0000 6800.0000 233600.0000 10000.0000 ;
    LAYER V1 ;
      RECT 86400.0000 6800.0000 89600.0000 10000.0000 ;
    LAYER V1 ;
      RECT 166400.0000 6800.0000 169600.0000 10000.0000 ;
    LAYER M3 ;
      RECT 118000.0000 13200.0000 122000.0000 20400.0000 ;
    LAYER V2 ;
      RECT 118000.0000 15200.0000 122000.0000 18400.0000 ;
    LAYER V2 ;
      RECT 118000.0000 15200.0000 122000.0000 18400.0000 ;
    LAYER V1 ;
      RECT 38400.0000 15200.0000 41600.0000 18400.0000 ;
    LAYER V1 ;
      RECT 214400.0000 15200.0000 217600.0000 18400.0000 ;
    LAYER M3 ;
      RECT 134000.0000 21600.0000 138000.0000 28800.0000 ;
    LAYER V2 ;
      RECT 134000.0000 23600.0000 138000.0000 26800.0000 ;
    LAYER V2 ;
      RECT 134000.0000 23600.0000 138000.0000 26800.0000 ;
    LAYER V1 ;
      RECT 102400.0000 23600.0000 105600.0000 26800.0000 ;
    LAYER V1 ;
      RECT 150400.0000 23600.0000 153600.0000 26800.0000 ;
    LAYER M3 ;
      RECT 110000.0000 30000.0000 114000.0000 37200.0000 ;
    LAYER V2 ;
      RECT 110000.0000 32000.0000 114000.0000 35200.0000 ;
    LAYER V2 ;
      RECT 110000.0000 32000.0000 114000.0000 35200.0000 ;
    LAYER V1 ;
      RECT 30400.0000 32000.0000 33600.0000 35200.0000 ;
    LAYER V1 ;
      RECT 222400.0000 32000.0000 225600.0000 35200.0000 ;
    LAYER M3 ;
      RECT 142000.0000 38400.0000 146000.0000 45600.0000 ;
    LAYER V2 ;
      RECT 142000.0000 40400.0000 146000.0000 43600.0000 ;
    LAYER V2 ;
      RECT 142000.0000 40400.0000 146000.0000 43600.0000 ;
    LAYER V1 ;
      RECT 94400.0000 40400.0000 97600.0000 43600.0000 ;
    LAYER V1 ;
      RECT 158400.0000 40400.0000 161600.0000 43600.0000 ;
    LAYER M1 ;
      RECT 30400.0000 88800.0000 33600.0000 154800.0000 ;
    LAYER M1 ;
      RECT 222400.0000 88800.0000 225600.0000 154800.0000 ;
    LAYER M1 ;
      RECT 94400.0000 88800.0000 97600.0000 154800.0000 ;
    LAYER M1 ;
      RECT 158400.0000 88800.0000 161600.0000 154800.0000 ;
    LAYER M1 ;
      RECT 22400.0000 88800.0000 25600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 22400.0000 107600.0000 25600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 22400.0000 120200.0000 25600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 22400.0000 132800.0000 25600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 230400.0000 88800.0000 233600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 230400.0000 107600.0000 233600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 230400.0000 120200.0000 233600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 230400.0000 132800.0000 233600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 86400.0000 88800.0000 89600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 86400.0000 107600.0000 89600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 86400.0000 120200.0000 89600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 86400.0000 132800.0000 89600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 166400.0000 88800.0000 169600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 166400.0000 107600.0000 169600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 166400.0000 120200.0000 169600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 166400.0000 132800.0000 169600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 38400.0000 88800.0000 41600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 38400.0000 107600.0000 41600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 38400.0000 120200.0000 41600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 38400.0000 132800.0000 41600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 214400.0000 88800.0000 217600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 214400.0000 107600.0000 217600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 214400.0000 120200.0000 217600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 214400.0000 132800.0000 217600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 102400.0000 88800.0000 105600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 102400.0000 107600.0000 105600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 102400.0000 120200.0000 105600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 102400.0000 132800.0000 105600.0000 136000.0000 ;
    LAYER M1 ;
      RECT 150400.0000 88800.0000 153600.0000 154800.0000 ;
    LAYER V0 ;
      RECT 150400.0000 107600.0000 153600.0000 110800.0000 ;
    LAYER V0 ;
      RECT 150400.0000 120200.0000 153600.0000 123400.0000 ;
    LAYER V0 ;
      RECT 150400.0000 132800.0000 153600.0000 136000.0000 ;
    LAYER M3 ;
      RECT 126000.0000 4800.0000 130000.0000 96000.0000 ;
    LAYER V2 ;
      RECT 126000.0000 6800.0000 130000.0000 10000.0000 ;
    LAYER V2 ;
      RECT 126000.0000 90800.0000 130000.0000 94000.0000 ;
    LAYER V1 ;
      RECT 22400.0000 90800.0000 25600.0000 94000.0000 ;
    LAYER V1 ;
      RECT 230400.0000 90800.0000 233600.0000 94000.0000 ;
    LAYER V1 ;
      RECT 86400.0000 90800.0000 89600.0000 94000.0000 ;
    LAYER V1 ;
      RECT 166400.0000 90800.0000 169600.0000 94000.0000 ;
    LAYER M3 ;
      RECT 118000.0000 13200.0000 122000.0000 104400.0000 ;
    LAYER V2 ;
      RECT 118000.0000 15200.0000 122000.0000 18400.0000 ;
    LAYER V2 ;
      RECT 118000.0000 99200.0000 122000.0000 102400.0000 ;
    LAYER V1 ;
      RECT 102400.0000 99200.0000 105600.0000 102400.0000 ;
    LAYER V1 ;
      RECT 150400.0000 99200.0000 153600.0000 102400.0000 ;
    LAYER M3 ;
      RECT 134000.0000 21600.0000 138000.0000 112800.0000 ;
    LAYER V2 ;
      RECT 134000.0000 23600.0000 138000.0000 26800.0000 ;
    LAYER V2 ;
      RECT 134000.0000 107600.0000 138000.0000 110800.0000 ;
    LAYER V1 ;
      RECT 38400.0000 107600.0000 41600.0000 110800.0000 ;
    LAYER V1 ;
      RECT 214400.0000 107600.0000 217600.0000 110800.0000 ;
    LAYER M3 ;
      RECT 110000.0000 30000.0000 114000.0000 121200.0000 ;
    LAYER V2 ;
      RECT 110000.0000 32000.0000 114000.0000 35200.0000 ;
    LAYER V2 ;
      RECT 110000.0000 116000.0000 114000.0000 119200.0000 ;
    LAYER V1 ;
      RECT 94400.0000 116000.0000 97600.0000 119200.0000 ;
    LAYER V1 ;
      RECT 158400.0000 116000.0000 161600.0000 119200.0000 ;
    LAYER M3 ;
      RECT 142000.0000 38400.0000 146000.0000 129600.0000 ;
    LAYER V2 ;
      RECT 142000.0000 40400.0000 146000.0000 43600.0000 ;
    LAYER V2 ;
      RECT 142000.0000 124400.0000 146000.0000 127600.0000 ;
    LAYER V1 ;
      RECT 30400.0000 124400.0000 33600.0000 127600.0000 ;
    LAYER V1 ;
      RECT 222400.0000 124400.0000 225600.0000 127600.0000 ;
  END
END __json_dp_nmos_cand
