MACRO CMC_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.8360 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 3.4760 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 3.6360 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 3.5560 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
  END
END CMC_NMOS_n12_X3_Y1
MACRO CMC_PMOS_S_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.4560 ;
      LAYER M3 ;
        RECT 0.7000 0.0480 0.7400 0.4560 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.5400 ;
      LAYER M3 ;
        RECT 0.7800 0.1320 0.8200 0.5400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.2160 0.5800 0.6240 ;
      LAYER M3 ;
        RECT 0.8600 0.2160 0.9000 0.6240 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.3000 0.6600 0.7080 ;
      LAYER M3 ;
        RECT 0.9400 0.3000 0.9800 0.7080 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 0.9160 0.4360 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4880 0.8360 0.5200 ;
    LAYER M2 ;
      RECT 0.5240 0.2360 1.0760 0.2680 ;
    LAYER M2 ;
      RECT 0.5240 0.5720 1.0760 0.6040 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 0.9960 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.6560 0.9960 0.6880 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END CMC_PMOS_S_n12_X1_Y1
MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 1.5560 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 2.2760 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
  END
END CMC_PMOS_n12_X2_Y1
MACRO CMFB_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMFB_NMOS_n12_X3_Y1 0 0 ;
  SIZE 5.1200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.3000 0.0480 2.3400 0.4560 ;
      LAYER M3 ;
        RECT 2.6200 0.0480 2.6600 0.4560 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.3800 0.1320 2.4200 0.5400 ;
      LAYER M3 ;
        RECT 2.7000 0.1320 2.7400 0.5400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.4600 0.2160 2.5000 0.6240 ;
      LAYER M3 ;
        RECT 2.7800 0.2160 2.8200 0.6240 ;
    END
  END DB
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.5400 0.3000 2.5800 0.7080 ;
      LAYER M3 ;
        RECT 2.8600 0.3000 2.9000 0.7080 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M1 ;
      RECT 4.1440 0.0480 4.1760 0.7080 ;
    LAYER M1 ;
      RECT 4.0640 0.0480 4.0960 0.7080 ;
    LAYER M1 ;
      RECT 4.2240 0.0480 4.2560 0.7080 ;
    LAYER M1 ;
      RECT 4.7840 0.0480 4.8160 0.7080 ;
    LAYER M1 ;
      RECT 4.7040 0.0480 4.7360 0.7080 ;
    LAYER M1 ;
      RECT 4.8640 0.0480 4.8960 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 4.7560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 4.7560 0.4360 ;
    LAYER M2 ;
      RECT 2.2040 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 2.2040 0.4880 2.9960 0.5200 ;
    LAYER M2 ;
      RECT 0.3640 0.2360 4.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.3640 0.5720 4.9160 0.6040 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 4.8360 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.6560 4.8360 0.6880 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
    LAYER pc ;
      RECT 4.1110 0.0680 4.2090 0.1000 ;
    LAYER pc ;
      RECT 4.7510 0.0680 4.8490 0.1000 ;
  END
END CMFB_NMOS_n12_X3_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.0480 0.5800 0.2880 ;
      LAYER M3 ;
        RECT 0.7000 0.0480 0.7400 0.2880 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.1320 0.6600 0.3720 ;
      LAYER M3 ;
        RECT 0.7800 0.1320 0.8200 0.3720 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 1.0760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 1.0760 0.3520 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DP_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 0.5960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.0760 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 0.5160 0.3520 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7640 0.4040 0.9960 0.4360 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END DP_NMOS_n12_X1_Y1
MACRO DP_NMOS_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X3_Y2 0 0 ;
  SIZE 3.8400 BY 1.6800 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.7400 0.0480 1.7800 0.9600 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.8200 0.1320 1.8600 1.0440 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9000 0.2160 1.9400 1.1280 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9800 0.3000 2.0200 1.2120 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.0600 0.3840 2.1000 1.2960 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.8880 3.5360 1.5480 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.4240 0.8880 3.4560 1.5480 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.8880 3.6160 1.5480 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 3.4760 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 1.0040 0.2360 3.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 2.9160 0.3520 ;
    LAYER M2 ;
      RECT 0.9240 0.4040 3.5560 0.4360 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 3.4760 0.9400 ;
    LAYER M2 ;
      RECT 1.0040 0.9920 3.6360 1.0240 ;
    LAYER M2 ;
      RECT 0.3640 1.0760 2.9960 1.1080 ;
    LAYER M2 ;
      RECT 0.9240 1.1600 3.5560 1.1920 ;
    LAYER M2 ;
      RECT 0.2840 1.2440 2.9160 1.2760 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 2.1910 0.0680 2.2890 0.1000 ;
    LAYER pc ;
      RECT 2.8310 0.0680 2.9290 0.1000 ;
    LAYER pc ;
      RECT 3.4710 0.0680 3.5690 0.1000 ;
    LAYER pc ;
      RECT 0.2710 0.9080 0.3690 0.9400 ;
    LAYER pc ;
      RECT 0.9110 0.9080 1.0090 0.9400 ;
    LAYER pc ;
      RECT 1.5510 0.9080 1.6490 0.9400 ;
    LAYER pc ;
      RECT 2.1910 0.9080 2.2890 0.9400 ;
    LAYER pc ;
      RECT 2.8310 0.9080 2.9290 0.9400 ;
    LAYER pc ;
      RECT 3.4710 0.9080 3.5690 0.9400 ;
  END
END DP_NMOS_n12_X3_Y2
MACRO Switch_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 0.3720 ;
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.4560 ;
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 0.5400 ;
      LAYER M3 ;
        RECT 0.5400 0.2160 0.5800 0.5400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 0.3200 0.4360 0.3520 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 0.5160 0.4360 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.5960 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.4880 0.5960 0.5200 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
  END
END Switch_NMOS_n12_X1_Y1
MACRO Switch_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y1 0 0 ;
  SIZE 1.9200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.0480 0.8200 0.3720 ;
      LAYER M3 ;
        RECT 1.0200 0.0480 1.0600 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8600 0.1320 0.9000 0.4560 ;
      LAYER M3 ;
        RECT 1.1000 0.1320 1.1400 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9400 0.2160 0.9800 0.5400 ;
      LAYER M3 ;
        RECT 1.1800 0.2160 1.2200 0.5400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 1.5560 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 1.7160 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 1.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 1.6360 0.5200 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
  END
END Switch_NMOS_n12_X3_Y1
MACRO Switch_NMOS_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y2 0 0 ;
  SIZE 1.9200 BY 1.6800 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.0480 0.8200 1.2120 ;
      LAYER M3 ;
        RECT 1.0200 0.0480 1.0600 1.2120 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8600 0.1320 0.9000 1.2960 ;
      LAYER M3 ;
        RECT 1.1000 0.1320 1.1400 1.2960 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9400 0.2160 0.9800 1.3800 ;
      LAYER M3 ;
        RECT 1.1800 0.2160 1.2200 1.3800 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 1.5560 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 1.7160 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 1.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 1.6360 0.5200 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 1.5560 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.1600 1.5560 1.1920 ;
    LAYER M2 ;
      RECT 0.3640 0.9920 1.7160 1.0240 ;
    LAYER M2 ;
      RECT 0.3640 1.2440 1.7160 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.0760 1.6360 1.1080 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 1.6360 1.3600 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
    LAYER pc ;
      RECT 1.5510 0.0680 1.6490 0.1000 ;
    LAYER pc ;
      RECT 0.2710 0.9080 0.3690 0.9400 ;
    LAYER pc ;
      RECT 0.9110 0.9080 1.0090 0.9400 ;
    LAYER pc ;
      RECT 1.5510 0.9080 1.6490 0.9400 ;
  END
END Switch_NMOS_n12_X3_Y2
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 0.3720 ;
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.4560 ;
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 0.5400 ;
      LAYER M3 ;
        RECT 0.5400 0.2160 0.5800 0.5400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 0.3200 0.4360 0.3520 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 0.5160 0.4360 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.5960 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.4880 0.5960 0.5200 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 0.3720 ;
      LAYER M3 ;
        RECT 0.7000 0.0480 0.7400 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 0.4560 ;
      LAYER M3 ;
        RECT 0.7800 0.1320 0.8200 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.2160 0.6600 0.5400 ;
      LAYER M3 ;
        RECT 0.8600 0.2160 0.9000 0.5400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 0.9160 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.0760 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 1.0760 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.9960 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 0.9960 0.5200 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END Switch_PMOS_n12_X2_Y1
MACRO cap_12f
  ORIGIN 0 0 ;
  FOREIGN cap_12f 0 0 ;
  SIZE 2.4000 BY 2.4360 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 -0.0160 2.4360 0.0160 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0360 2.4200 2.4360 2.4520 ;
    END
  END MINUS
  OBS
    LAYER boundary ;
      RECT 0.0000 0.0000 2.4000 2.4360 ;
    LAYER M1 ;
      RECT -0.0160 -0.0360 0.0160 2.4720 ;
    LAYER M1 ;
      RECT 0.0480 -0.0360 0.0800 2.4720 ;
    LAYER M1 ;
      RECT 0.1120 -0.0360 0.1440 2.4720 ;
    LAYER M1 ;
      RECT 0.1760 -0.0360 0.2080 2.4720 ;
    LAYER M1 ;
      RECT 0.2400 -0.0360 0.2720 2.4720 ;
    LAYER M1 ;
      RECT 0.3040 -0.0360 0.3360 2.4720 ;
    LAYER M1 ;
      RECT 0.3680 -0.0360 0.4000 2.4720 ;
    LAYER M1 ;
      RECT 0.4320 -0.0360 0.4640 2.4720 ;
    LAYER M1 ;
      RECT 0.4960 -0.0360 0.5280 2.4720 ;
    LAYER M1 ;
      RECT 0.5600 -0.0360 0.5920 2.4720 ;
    LAYER M1 ;
      RECT 0.6240 -0.0360 0.6560 2.4720 ;
    LAYER M1 ;
      RECT 0.6880 -0.0360 0.7200 2.4720 ;
    LAYER M1 ;
      RECT 0.7520 -0.0360 0.7840 2.4720 ;
    LAYER M1 ;
      RECT 0.8160 -0.0360 0.8480 2.4720 ;
    LAYER M1 ;
      RECT 0.8800 -0.0360 0.9120 2.4720 ;
    LAYER M1 ;
      RECT 0.9440 -0.0360 0.9760 2.4720 ;
    LAYER M1 ;
      RECT 1.0080 -0.0360 1.0400 2.4720 ;
    LAYER M1 ;
      RECT 1.0720 -0.0360 1.1040 2.4720 ;
    LAYER M1 ;
      RECT 1.1360 -0.0360 1.1680 2.4720 ;
    LAYER M1 ;
      RECT 1.2000 -0.0360 1.2320 2.4720 ;
    LAYER M1 ;
      RECT 1.2640 -0.0360 1.2960 2.4720 ;
    LAYER M1 ;
      RECT 1.3280 -0.0360 1.3600 2.4720 ;
    LAYER M1 ;
      RECT 1.3920 -0.0360 1.4240 2.4720 ;
    LAYER M1 ;
      RECT 1.4560 -0.0360 1.4880 2.4720 ;
    LAYER M1 ;
      RECT 1.5200 -0.0360 1.5520 2.4720 ;
    LAYER M1 ;
      RECT 1.5840 -0.0360 1.6160 2.4720 ;
    LAYER M1 ;
      RECT 1.6480 -0.0360 1.6800 2.4720 ;
    LAYER M1 ;
      RECT 1.7120 -0.0360 1.7440 2.4720 ;
    LAYER M1 ;
      RECT 1.7760 -0.0360 1.8080 2.4720 ;
    LAYER M1 ;
      RECT 1.8400 -0.0360 1.8720 2.4720 ;
    LAYER M1 ;
      RECT 1.9040 -0.0360 1.9360 2.4720 ;
    LAYER M1 ;
      RECT 1.9680 -0.0360 2.0000 2.4720 ;
    LAYER M1 ;
      RECT 2.0320 -0.0360 2.0640 2.4720 ;
    LAYER M1 ;
      RECT 2.0960 -0.0360 2.1280 2.4720 ;
    LAYER M1 ;
      RECT 2.1600 -0.0360 2.1920 2.4720 ;
    LAYER M1 ;
      RECT 2.2240 -0.0360 2.2560 2.4720 ;
    LAYER M1 ;
      RECT 2.2880 -0.0360 2.3200 2.4720 ;
    LAYER M1 ;
      RECT 2.3840 -0.0360 2.4160 2.4720 ;
    LAYER M2 ;
      RECT -0.0360 0.0480 2.4360 0.0800 ;
    LAYER M2 ;
      RECT -0.0360 0.1120 2.4360 0.1440 ;
    LAYER M2 ;
      RECT -0.0360 0.1760 2.4360 0.2080 ;
    LAYER M2 ;
      RECT -0.0360 0.2400 2.4360 0.2720 ;
    LAYER M2 ;
      RECT -0.0360 0.3040 2.4360 0.3360 ;
    LAYER M2 ;
      RECT -0.0360 0.3680 2.4360 0.4000 ;
    LAYER M2 ;
      RECT -0.0360 0.4320 2.4360 0.4640 ;
    LAYER M2 ;
      RECT -0.0360 0.4960 2.4360 0.5280 ;
    LAYER M2 ;
      RECT -0.0360 0.5600 2.4360 0.5920 ;
    LAYER M2 ;
      RECT -0.0360 0.6240 2.4360 0.6560 ;
    LAYER M2 ;
      RECT -0.0360 0.6880 2.4360 0.7200 ;
    LAYER M2 ;
      RECT -0.0360 0.7520 2.4360 0.7840 ;
    LAYER M2 ;
      RECT -0.0360 0.8160 2.4360 0.8480 ;
    LAYER M2 ;
      RECT -0.0360 0.8800 2.4360 0.9120 ;
    LAYER M2 ;
      RECT -0.0360 0.9440 2.4360 0.9760 ;
    LAYER M2 ;
      RECT -0.0360 1.0080 2.4360 1.0400 ;
    LAYER M2 ;
      RECT -0.0360 1.0720 2.4360 1.1040 ;
    LAYER M2 ;
      RECT -0.0360 1.1360 2.4360 1.1680 ;
    LAYER M2 ;
      RECT -0.0360 1.2000 2.4360 1.2320 ;
    LAYER M2 ;
      RECT -0.0360 1.2640 2.4360 1.2960 ;
    LAYER M2 ;
      RECT -0.0360 1.3280 2.4360 1.3600 ;
    LAYER M2 ;
      RECT -0.0360 1.3920 2.4360 1.4240 ;
    LAYER M2 ;
      RECT -0.0360 1.4560 2.4360 1.4880 ;
    LAYER M2 ;
      RECT -0.0360 1.5200 2.4360 1.5520 ;
    LAYER M2 ;
      RECT -0.0360 1.5840 2.4360 1.6160 ;
    LAYER M2 ;
      RECT -0.0360 1.6480 2.4360 1.6800 ;
    LAYER M2 ;
      RECT -0.0360 1.7120 2.4360 1.7440 ;
    LAYER M2 ;
      RECT -0.0360 1.7760 2.4360 1.8080 ;
    LAYER M2 ;
      RECT -0.0360 1.8400 2.4360 1.8720 ;
    LAYER M2 ;
      RECT -0.0360 1.9040 2.4360 1.9360 ;
    LAYER M2 ;
      RECT -0.0360 1.9680 2.4360 2.0000 ;
    LAYER M2 ;
      RECT -0.0360 2.0320 2.4360 2.0640 ;
    LAYER M2 ;
      RECT -0.0360 2.0960 2.4360 2.1280 ;
    LAYER M2 ;
      RECT -0.0360 2.1600 2.4360 2.1920 ;
    LAYER M2 ;
      RECT -0.0360 2.2240 2.4360 2.2560 ;
    LAYER M2 ;
      RECT -0.0360 2.2880 2.4360 2.3200 ;
    LAYER M3 ;
      RECT -0.0160 -0.0360 0.0160 2.4720 ;
    LAYER M3 ;
      RECT 0.0480 -0.0360 0.0800 2.4720 ;
    LAYER M3 ;
      RECT 0.1120 -0.0360 0.1440 2.4720 ;
    LAYER M3 ;
      RECT 0.1760 -0.0360 0.2080 2.4720 ;
    LAYER M3 ;
      RECT 0.2400 -0.0360 0.2720 2.4720 ;
    LAYER M3 ;
      RECT 0.3040 -0.0360 0.3360 2.4720 ;
    LAYER M3 ;
      RECT 0.3680 -0.0360 0.4000 2.4720 ;
    LAYER M3 ;
      RECT 0.4320 -0.0360 0.4640 2.4720 ;
    LAYER M3 ;
      RECT 0.4960 -0.0360 0.5280 2.4720 ;
    LAYER M3 ;
      RECT 0.5600 -0.0360 0.5920 2.4720 ;
    LAYER M3 ;
      RECT 0.6240 -0.0360 0.6560 2.4720 ;
    LAYER M3 ;
      RECT 0.6880 -0.0360 0.7200 2.4720 ;
    LAYER M3 ;
      RECT 0.7520 -0.0360 0.7840 2.4720 ;
    LAYER M3 ;
      RECT 0.8160 -0.0360 0.8480 2.4720 ;
    LAYER M3 ;
      RECT 0.8800 -0.0360 0.9120 2.4720 ;
    LAYER M3 ;
      RECT 0.9440 -0.0360 0.9760 2.4720 ;
    LAYER M3 ;
      RECT 1.0080 -0.0360 1.0400 2.4720 ;
    LAYER M3 ;
      RECT 1.0720 -0.0360 1.1040 2.4720 ;
    LAYER M3 ;
      RECT 1.1360 -0.0360 1.1680 2.4720 ;
    LAYER M3 ;
      RECT 1.2000 -0.0360 1.2320 2.4720 ;
    LAYER M3 ;
      RECT 1.2640 -0.0360 1.2960 2.4720 ;
    LAYER M3 ;
      RECT 1.3280 -0.0360 1.3600 2.4720 ;
    LAYER M3 ;
      RECT 1.3920 -0.0360 1.4240 2.4720 ;
    LAYER M3 ;
      RECT 1.4560 -0.0360 1.4880 2.4720 ;
    LAYER M3 ;
      RECT 1.5200 -0.0360 1.5520 2.4720 ;
    LAYER M3 ;
      RECT 1.5840 -0.0360 1.6160 2.4720 ;
    LAYER M3 ;
      RECT 1.6480 -0.0360 1.6800 2.4720 ;
    LAYER M3 ;
      RECT 1.7120 -0.0360 1.7440 2.4720 ;
    LAYER M3 ;
      RECT 1.7760 -0.0360 1.8080 2.4720 ;
    LAYER M3 ;
      RECT 1.8400 -0.0360 1.8720 2.4720 ;
    LAYER M3 ;
      RECT 1.9040 -0.0360 1.9360 2.4720 ;
    LAYER M3 ;
      RECT 1.9680 -0.0360 2.0000 2.4720 ;
    LAYER M3 ;
      RECT 2.0320 -0.0360 2.0640 2.4720 ;
    LAYER M3 ;
      RECT 2.0960 -0.0360 2.1280 2.4720 ;
    LAYER M3 ;
      RECT 2.1600 -0.0360 2.1920 2.4720 ;
    LAYER M3 ;
      RECT 2.2240 -0.0360 2.2560 2.4720 ;
    LAYER M3 ;
      RECT 2.2880 -0.0360 2.3200 2.4720 ;
    LAYER M3 ;
      RECT 2.3840 -0.0360 2.4160 2.4720 ;
  END
END cap_12f
