MACRO CMC_S_NMOS_B_nfin10_n12_X1_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN CMC_S_NMOS_B_nfin10_n12_X1_Y1_RVT 0 0 ;
  SIZE 1.2800 BY 1.8480 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.4360 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.5160 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.0760 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.7640 0.3200 0.9960 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.9960 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 0.9960 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
  END
END CMC_S_NMOS_B_nfin10_n12_X1_Y1_RVT
MACRO DP_NMOS_B_nfin75_n12_X7_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin75_n12_X7_Y1_RVT 0 0 ;
  SIZE 2.7200 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.5160 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 2.2760 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 2.4360 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 2.2760 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.9920 2.4360 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 2.4360 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 0.7920 ;
    LAYER M1 ;
      RECT 1.2640 0.8880 1.2960 1.1280 ;
    LAYER M1 ;
      RECT 1.2640 1.3920 1.2960 1.6320 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.0480 1.4560 0.7920 ;
    LAYER M1 ;
      RECT 1.4240 0.8880 1.4560 1.1280 ;
    LAYER M1 ;
      RECT 1.4240 1.3920 1.4560 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.3920 1.6160 1.6320 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.0480 1.7760 0.7920 ;
    LAYER M1 ;
      RECT 1.7440 0.8880 1.7760 1.1280 ;
    LAYER M1 ;
      RECT 1.7440 1.3920 1.7760 1.6320 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 0.7920 ;
    LAYER M1 ;
      RECT 1.9040 0.8880 1.9360 1.1280 ;
    LAYER M1 ;
      RECT 1.9040 1.3920 1.9360 1.6320 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.0480 2.0960 0.7920 ;
    LAYER M1 ;
      RECT 2.0640 0.8880 2.0960 1.1280 ;
    LAYER M1 ;
      RECT 2.0640 1.3920 2.0960 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.3920 2.2560 1.6320 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.0480 2.4160 0.7920 ;
    LAYER M1 ;
      RECT 2.3840 0.8880 2.4160 1.1280 ;
    LAYER M1 ;
      RECT 2.3840 1.3920 2.4160 1.6320 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.3440 0.0680 1.3760 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.9840 0.0680 2.0160 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 1.2640 0.1520 1.2960 0.1840 ;
    LAYER V1 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V1 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V1 ;
      RECT 1.5840 0.1520 1.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V1 ;
      RECT 1.9040 0.1520 1.9360 0.1840 ;
    LAYER V1 ;
      RECT 1.9040 0.9080 1.9360 0.9400 ;
    LAYER V1 ;
      RECT 1.9040 1.4960 1.9360 1.5280 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9920 0.8160 1.0240 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V1 ;
      RECT 1.4240 0.2360 1.4560 0.2680 ;
    LAYER V1 ;
      RECT 1.4240 0.9920 1.4560 1.0240 ;
    LAYER V1 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V1 ;
      RECT 1.7440 0.2360 1.7760 0.2680 ;
    LAYER V1 ;
      RECT 1.7440 0.9920 1.7760 1.0240 ;
    LAYER V1 ;
      RECT 1.7440 1.4960 1.7760 1.5280 ;
    LAYER V1 ;
      RECT 2.0640 0.2360 2.0960 0.2680 ;
    LAYER V1 ;
      RECT 2.0640 0.9920 2.0960 1.0240 ;
    LAYER V1 ;
      RECT 2.0640 1.4960 2.0960 1.5280 ;
    LAYER V1 ;
      RECT 2.3840 0.2360 2.4160 0.2680 ;
    LAYER V1 ;
      RECT 2.3840 0.9920 2.4160 1.0240 ;
    LAYER V1 ;
      RECT 2.3840 1.4960 2.4160 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.4040 1.2960 0.4360 ;
    LAYER V0 ;
      RECT 1.2640 0.5300 1.2960 0.5620 ;
    LAYER V0 ;
      RECT 1.2640 0.6560 1.2960 0.6880 ;
    LAYER V0 ;
      RECT 1.2640 0.9080 1.2960 0.9400 ;
    LAYER V0 ;
      RECT 1.2640 1.4960 1.2960 1.5280 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.4040 1.4560 0.4360 ;
    LAYER V0 ;
      RECT 1.4240 0.5300 1.4560 0.5620 ;
    LAYER V0 ;
      RECT 1.4240 0.6560 1.4560 0.6880 ;
    LAYER V0 ;
      RECT 1.4240 0.9080 1.4560 0.9400 ;
    LAYER V0 ;
      RECT 1.4240 1.4960 1.4560 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.4040 1.7760 0.4360 ;
    LAYER V0 ;
      RECT 1.7440 0.5300 1.7760 0.5620 ;
    LAYER V0 ;
      RECT 1.7440 0.6560 1.7760 0.6880 ;
    LAYER V0 ;
      RECT 1.7440 0.9080 1.7760 0.9400 ;
    LAYER V0 ;
      RECT 1.7440 1.4960 1.7760 1.5280 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.4040 1.9360 0.4360 ;
    LAYER V0 ;
      RECT 1.9040 0.5300 1.9360 0.5620 ;
    LAYER V0 ;
      RECT 1.9040 0.6560 1.9360 0.6880 ;
    LAYER V0 ;
      RECT 1.9040 0.9080 1.9360 0.9400 ;
    LAYER V0 ;
      RECT 1.9040 1.4960 1.9360 1.5280 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.4040 2.0960 0.4360 ;
    LAYER V0 ;
      RECT 2.0640 0.5300 2.0960 0.5620 ;
    LAYER V0 ;
      RECT 2.0640 0.6560 2.0960 0.6880 ;
    LAYER V0 ;
      RECT 2.0640 0.9080 2.0960 0.9400 ;
    LAYER V0 ;
      RECT 2.0640 1.4960 2.0960 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.4040 2.4160 0.4360 ;
    LAYER V0 ;
      RECT 2.3840 0.5300 2.4160 0.5620 ;
    LAYER V0 ;
      RECT 2.3840 0.6560 2.4160 0.6880 ;
    LAYER V0 ;
      RECT 2.3840 0.9080 2.4160 0.9400 ;
    LAYER V0 ;
      RECT 2.3840 1.4960 2.4160 1.5280 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
  END
END DP_NMOS_B_nfin75_n12_X7_Y1_RVT
MACRO CMC_S_PMOS_B_nfin15_n12_X2_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN CMC_S_PMOS_B_nfin15_n12_X2_Y1_RVT 0 0 ;
  SIZE 2.5600 BY 1.8480 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 2.2760 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.3200 1.6360 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 2.2760 0.9400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 2.2760 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7920 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.1280 ;
    LAYER M1 ;
      RECT 1.5840 1.3920 1.6160 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7920 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.1280 ;
    LAYER M1 ;
      RECT 2.2240 1.3920 2.2560 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V1 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.3200 1.6160 0.3520 ;
    LAYER V1 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V1 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V0 ;
      RECT 1.5840 0.5300 1.6160 0.5620 ;
    LAYER V0 ;
      RECT 1.5840 0.6560 1.6160 0.6880 ;
    LAYER V0 ;
      RECT 1.5840 0.9080 1.6160 0.9400 ;
    LAYER V0 ;
      RECT 1.5840 1.4960 1.6160 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V0 ;
      RECT 2.2240 0.5300 2.2560 0.5620 ;
    LAYER V0 ;
      RECT 2.2240 0.6560 2.2560 0.6880 ;
    LAYER V0 ;
      RECT 2.2240 0.9080 2.2560 0.9400 ;
    LAYER V0 ;
      RECT 2.2240 1.4960 2.2560 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
  END
END CMC_S_PMOS_B_nfin15_n12_X2_Y1_RVT
MACRO CMC_PMOS_nfin15_nf2_n12_X3_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_nfin15_nf2_n12_X3_Y1_RVT 0 0 ;
  SIZE 1.4400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 1.1560 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 1.1560 0.9400 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M2 ;
      RECT 0.2840 1.4960 1.1560 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
  END
END CMC_PMOS_nfin15_nf2_n12_X3_Y1_RVT
MACRO SCM_NMOS_nfin15_nf2_n12_X3_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin15_nf2_n12_X3_Y1_RVT 0 0 ;
  SIZE 1.4400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 1.1560 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M2 ;
      RECT 0.2840 1.4960 1.1560 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.2360 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 1.1560 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.9960 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.5440 0.1520 0.5760 0.1840 ;
    LAYER V2 ;
      RECT 0.5440 0.9080 0.5760 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
  END
END SCM_NMOS_nfin15_nf2_n12_X3_Y1_RVT
MACRO guard_ring
  ORIGIN 0 0 ;
  FOREIGN guard_ring 0 0 ;
  SIZE 1.4400 BY 1.4280 ;
  PIN Body
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3440 0.3360 1.0960 1.0920 ;
    END
  END Body
  OBS
    LAYER V0 ;
      RECT 0.3840 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 1.0560 0.5200 ;
    LAYER V0 ;
      RECT 0.3840 0.5720 1.0560 0.6040 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.7400 1.0560 0.7720 ;
    LAYER V0 ;
      RECT 0.3840 0.8240 1.0560 0.8560 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 0.9920 1.0560 1.0240 ;
  END
END guard_ring