MACRO switched_capacitor_filter
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_filter 0 0 ;
  SIZE 46.08 BY 37.8 ;
  PIN id
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.184 -0.016 23.216 0.016 ;
      LAYER M3 ;
        RECT 23.18 0.3 23.22 0.708 ;
      LAYER M3 ;
        RECT 22.86 0.3 22.9 0.708 ;
      LAYER M3 ;
        RECT 23.18 0.316 23.22 0.356 ;
      LAYER M4 ;
        RECT 23.04 0.316 23.2 0.356 ;
      LAYER M5 ;
        RECT 23.008 0 23.072 0.336 ;
      LAYER M4 ;
        RECT 23.04 -0.02 23.2 0.02 ;
      LAYER M3 ;
        RECT 23.18 -0.02 23.22 0.02 ;
      LAYER M2 ;
        RECT 23.184 -0.016 23.216 0.016 ;
    END
  END id
  PIN voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.344 37.784 15.376 37.816 ;
      LAYER M2 ;
        RECT 22.124 4.436 23.956 4.468 ;
      LAYER M2 ;
        RECT 21.964 3.008 24.596 3.04 ;
      LAYER M2 ;
        RECT 22.544 4.436 22.576 4.468 ;
      LAYER M3 ;
        RECT 22.54 3.192 22.58 4.452 ;
      LAYER M4 ;
        RECT 22.54 3.172 22.58 3.212 ;
      LAYER M5 ;
        RECT 22.528 3.024 22.592 3.192 ;
      LAYER M4 ;
        RECT 22.54 3.004 22.58 3.044 ;
      LAYER M3 ;
        RECT 22.54 3.004 22.58 3.044 ;
      LAYER M2 ;
        RECT 22.544 3.008 22.576 3.04 ;
      LAYER M2 ;
        RECT 7.244 0.824 7.476 0.856 ;
      LAYER M1 ;
        RECT 11.744 1.308 11.776 1.38 ;
      LAYER M2 ;
        RECT 11.724 1.328 11.796 1.36 ;
      LAYER M1 ;
        RECT 3.104 1.308 3.136 1.38 ;
      LAYER M2 ;
        RECT 3.084 1.328 3.156 1.36 ;
      LAYER M2 ;
        RECT 3.12 1.328 11.76 1.36 ;
      LAYER M2 ;
        RECT 7.424 0.824 7.456 0.856 ;
      LAYER M3 ;
        RECT 7.42 0.84 7.46 1.344 ;
      LAYER M2 ;
        RECT 7.424 1.328 7.456 1.36 ;
      LAYER M1 ;
        RECT 21.504 37.344 21.536 37.416 ;
      LAYER M2 ;
        RECT 21.484 37.364 21.556 37.396 ;
      LAYER M1 ;
        RECT 24.384 37.344 24.416 37.416 ;
      LAYER M2 ;
        RECT 24.364 37.364 24.436 37.396 ;
      LAYER M2 ;
        RECT 21.52 37.364 24.4 37.396 ;
      LAYER M2 ;
        RECT 21.04 3.008 22 3.04 ;
      LAYER M3 ;
        RECT 21.02 3.004 21.06 3.044 ;
      LAYER M4 ;
        RECT 20.88 3.004 21.04 3.044 ;
      LAYER M5 ;
        RECT 20.848 3.024 20.912 3.36 ;
      LAYER M4 ;
        RECT 12.816 3.34 20.88 3.38 ;
      LAYER M5 ;
        RECT 12.784 1.596 12.848 3.36 ;
      LAYER M4 ;
        RECT 12.24 1.576 12.816 1.616 ;
      LAYER M3 ;
        RECT 12.22 1.344 12.26 1.596 ;
      LAYER M2 ;
        RECT 11.76 1.328 12.24 1.36 ;
      LAYER M2 ;
        RECT 23.744 4.436 23.776 4.468 ;
      LAYER M3 ;
        RECT 23.74 4.452 23.78 4.956 ;
      LAYER M4 ;
        RECT 23.76 4.936 25.632 4.976 ;
      LAYER M5 ;
        RECT 25.6 4.956 25.664 37.38 ;
      LAYER M4 ;
        RECT 25.2 37.36 25.632 37.4 ;
      LAYER M3 ;
        RECT 25.18 37.36 25.22 37.4 ;
      LAYER M2 ;
        RECT 24.72 37.364 25.2 37.396 ;
      LAYER M3 ;
        RECT 24.7 37.36 24.74 37.4 ;
      LAYER M4 ;
        RECT 24.4 37.36 24.72 37.4 ;
      LAYER M3 ;
        RECT 24.38 37.36 24.42 37.4 ;
      LAYER M2 ;
        RECT 24.384 37.364 24.416 37.396 ;
      LAYER M2 ;
        RECT 20.08 37.364 21.52 37.396 ;
      LAYER M3 ;
        RECT 20.06 36.372 20.1 37.38 ;
      LAYER M4 ;
        RECT 19.296 36.352 20.08 36.392 ;
      LAYER M5 ;
        RECT 19.264 35.28 19.328 36.372 ;
      LAYER M6 ;
        RECT 15.84 35.248 19.296 35.312 ;
      LAYER M5 ;
        RECT 15.808 35.28 15.872 37.548 ;
      LAYER M4 ;
        RECT 15.82 37.528 15.86 37.568 ;
      LAYER M3 ;
        RECT 15.82 37.528 15.86 37.568 ;
      LAYER M2 ;
        RECT 15.36 37.532 15.84 37.564 ;
      LAYER M3 ;
        RECT 15.34 37.548 15.38 37.8 ;
      LAYER M2 ;
        RECT 15.344 37.784 15.376 37.816 ;
    END
  END voutn
  PIN voutp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 30.704 37.784 30.736 37.816 ;
      LAYER M2 ;
        RECT 22.764 4.268 23.316 4.3 ;
      LAYER M2 ;
        RECT 21.324 3.176 23.956 3.208 ;
      LAYER M2 ;
        RECT 23.264 4.268 23.296 4.3 ;
      LAYER M3 ;
        RECT 23.26 4.032 23.3 4.284 ;
      LAYER M4 ;
        RECT 23.26 4.012 23.3 4.052 ;
      LAYER M5 ;
        RECT 23.248 3.696 23.312 4.032 ;
      LAYER M4 ;
        RECT 23.26 3.676 23.3 3.716 ;
      LAYER M3 ;
        RECT 23.26 3.192 23.3 3.696 ;
      LAYER M2 ;
        RECT 23.264 3.176 23.296 3.208 ;
      LAYER M2 ;
        RECT 38.604 0.824 38.836 0.856 ;
      LAYER M1 ;
        RECT 34.304 1.308 34.336 1.38 ;
      LAYER M2 ;
        RECT 34.284 1.328 34.356 1.36 ;
      LAYER M1 ;
        RECT 42.944 1.308 42.976 1.38 ;
      LAYER M2 ;
        RECT 42.924 1.328 42.996 1.36 ;
      LAYER M2 ;
        RECT 34.32 1.328 42.96 1.36 ;
      LAYER M2 ;
        RECT 38.624 0.824 38.656 0.856 ;
      LAYER M3 ;
        RECT 38.62 0.84 38.66 1.344 ;
      LAYER M2 ;
        RECT 38.624 1.328 38.656 1.36 ;
      LAYER M1 ;
        RECT 18.624 37.512 18.656 37.584 ;
      LAYER M2 ;
        RECT 18.604 37.532 18.676 37.564 ;
      LAYER M1 ;
        RECT 27.264 37.512 27.296 37.584 ;
      LAYER M2 ;
        RECT 27.244 37.532 27.316 37.564 ;
      LAYER M2 ;
        RECT 18.64 37.532 27.28 37.564 ;
      LAYER M2 ;
        RECT 23.92 3.176 25.36 3.208 ;
      LAYER M3 ;
        RECT 25.34 3.172 25.38 3.212 ;
      LAYER M4 ;
        RECT 25.36 3.172 25.488 3.212 ;
      LAYER M5 ;
        RECT 25.456 3.192 25.52 3.36 ;
      LAYER M4 ;
        RECT 25.488 3.34 33.552 3.38 ;
      LAYER M5 ;
        RECT 33.52 1.596 33.584 3.36 ;
      LAYER M4 ;
        RECT 33.552 1.576 34.32 1.616 ;
      LAYER M3 ;
        RECT 34.3 1.344 34.34 1.596 ;
      LAYER M2 ;
        RECT 34.304 1.328 34.336 1.36 ;
      LAYER M4 ;
        RECT 25.9 3.34 25.94 3.38 ;
      LAYER M3 ;
        RECT 25.9 3.36 25.94 5.628 ;
      LAYER M4 ;
        RECT 25.9 5.608 25.94 5.648 ;
      LAYER M5 ;
        RECT 25.888 5.628 25.952 37.548 ;
      LAYER M4 ;
        RECT 25.9 37.528 25.94 37.568 ;
      LAYER M3 ;
        RECT 25.9 37.528 25.94 37.568 ;
      LAYER M2 ;
        RECT 25.904 37.532 25.936 37.564 ;
      LAYER M2 ;
        RECT 27.28 37.532 30.4 37.564 ;
      LAYER M3 ;
        RECT 30.38 37.548 30.42 37.8 ;
      LAYER M4 ;
        RECT 30.4 37.78 30.72 37.82 ;
      LAYER M3 ;
        RECT 30.7 37.78 30.74 37.82 ;
      LAYER M2 ;
        RECT 30.704 37.784 30.736 37.816 ;
    END
  END voutp
  PIN vss
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.344 -0.016 23.376 0.016 ;
      LAYER M3 ;
        RECT 23.26 0.216 23.3 0.624 ;
      LAYER M3 ;
        RECT 22.94 0.216 22.98 0.624 ;
      LAYER M1 ;
        RECT 21.664 19.2 21.696 19.272 ;
      LAYER M2 ;
        RECT 21.644 19.22 21.716 19.252 ;
      LAYER M1 ;
        RECT 24.544 19.2 24.576 19.272 ;
      LAYER M2 ;
        RECT 24.524 19.22 24.596 19.252 ;
      LAYER M2 ;
        RECT 21.68 19.22 24.56 19.252 ;
      LAYER M1 ;
        RECT 18.784 19.032 18.816 19.104 ;
      LAYER M2 ;
        RECT 18.764 19.052 18.836 19.084 ;
      LAYER M1 ;
        RECT 27.424 19.032 27.456 19.104 ;
      LAYER M2 ;
        RECT 27.404 19.052 27.476 19.084 ;
      LAYER M2 ;
        RECT 18.8 19.052 27.44 19.084 ;
      LAYER M3 ;
        RECT 23.26 0.232 23.3 0.272 ;
      LAYER M4 ;
        RECT 23.28 0.232 23.6 0.272 ;
      LAYER M3 ;
        RECT 23.58 0 23.62 0.252 ;
      LAYER M2 ;
        RECT 23.36 -0.016 23.6 0.016 ;
      LAYER M3 ;
        RECT 23.26 0.588 23.3 1.344 ;
      LAYER M2 ;
        RECT 23.28 1.328 25.68 1.36 ;
      LAYER M3 ;
        RECT 25.66 1.344 25.7 19.236 ;
      LAYER M2 ;
        RECT 24.48 19.22 25.68 19.252 ;
      LAYER M3 ;
        RECT 25.66 19.048 25.7 19.088 ;
      LAYER M2 ;
        RECT 25.664 19.052 25.696 19.084 ;
    END
  END vss
  PIN vinn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.024 -0.016 15.056 0.016 ;
      LAYER M3 ;
        RECT 15.02 17.688 15.06 18.012 ;
      LAYER M3 ;
        RECT 15.26 17.688 15.3 18.012 ;
      LAYER M1 ;
        RECT 27.424 18.444 27.456 18.516 ;
      LAYER M2 ;
        RECT 27.404 18.464 27.476 18.496 ;
      LAYER M1 ;
        RECT 18.784 18.444 18.816 18.516 ;
      LAYER M2 ;
        RECT 18.764 18.464 18.836 18.496 ;
      LAYER M2 ;
        RECT 18.8 18.464 27.44 18.496 ;
      LAYER M3 ;
        RECT 15.26 17.976 15.3 18.48 ;
      LAYER M2 ;
        RECT 15.28 18.464 18.88 18.496 ;
      LAYER M3 ;
        RECT 15.02 16.968 15.06 17.724 ;
      LAYER M4 ;
        RECT 14.4 16.948 15.04 16.988 ;
      LAYER M5 ;
        RECT 14.368 0 14.432 16.968 ;
      LAYER M4 ;
        RECT 14.4 -0.02 15.04 0.02 ;
      LAYER M3 ;
        RECT 15.02 -0.02 15.06 0.02 ;
      LAYER M2 ;
        RECT 15.024 -0.016 15.056 0.016 ;
    END
  END vinn
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.344 -0.016 15.376 0.016 ;
      LAYER M3 ;
        RECT 4.94 0.636 4.98 0.96 ;
      LAYER M3 ;
        RECT 5.18 0.636 5.22 0.96 ;
      LAYER M2 ;
        RECT 5.724 0.74 5.956 0.772 ;
      LAYER M2 ;
        RECT 7.724 0.74 7.956 0.772 ;
      LAYER M3 ;
        RECT 5.18 0.736 5.22 0.776 ;
      LAYER M4 ;
        RECT 5.2 0.736 5.52 0.776 ;
      LAYER M3 ;
        RECT 5.5 0.736 5.54 0.776 ;
      LAYER M2 ;
        RECT 5.52 0.74 5.76 0.772 ;
      LAYER M2 ;
        RECT 5.92 0.74 7.84 0.772 ;
      LAYER M3 ;
        RECT 41.1 0.636 41.14 0.96 ;
      LAYER M3 ;
        RECT 40.86 0.636 40.9 0.96 ;
      LAYER M2 ;
        RECT 40.124 0.74 40.356 0.772 ;
      LAYER M2 ;
        RECT 38.124 0.74 38.356 0.772 ;
      LAYER M3 ;
        RECT 40.86 0.736 40.9 0.776 ;
      LAYER M4 ;
        RECT 40.56 0.736 40.88 0.776 ;
      LAYER M3 ;
        RECT 40.54 0.736 40.58 0.776 ;
      LAYER M2 ;
        RECT 40.32 0.74 40.56 0.772 ;
      LAYER M2 ;
        RECT 38.24 0.74 40.16 0.772 ;
      LAYER M2 ;
        RECT 7.904 0.74 7.936 0.772 ;
      LAYER M3 ;
        RECT 7.9 0.736 7.94 0.776 ;
      LAYER M4 ;
        RECT 7.9 0.736 7.94 0.776 ;
      LAYER M5 ;
        RECT 7.888 0.756 7.952 1.68 ;
      LAYER M4 ;
        RECT 7.92 1.66 14.256 1.7 ;
      LAYER M5 ;
        RECT 14.224 0.756 14.288 1.68 ;
      LAYER M4 ;
        RECT 14.256 0.736 15.36 0.776 ;
      LAYER M3 ;
        RECT 15.34 0 15.38 0.756 ;
      LAYER M2 ;
        RECT 15.344 -0.016 15.376 0.016 ;
      LAYER M5 ;
        RECT 14.224 1.596 14.288 5.04 ;
      LAYER M4 ;
        RECT 14.256 5.02 17.568 5.06 ;
      LAYER M5 ;
        RECT 17.536 5.04 17.6 6.72 ;
      LAYER M4 ;
        RECT 17.568 6.7 38.16 6.74 ;
      LAYER M5 ;
        RECT 38.128 0.756 38.192 6.72 ;
      LAYER M4 ;
        RECT 38.14 0.736 38.18 0.776 ;
      LAYER M3 ;
        RECT 38.14 0.736 38.18 0.776 ;
      LAYER M2 ;
        RECT 38.144 0.74 38.176 0.772 ;
    END
  END agnd
  PIN vinp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.024 -0.016 31.056 0.016 ;
      LAYER M3 ;
        RECT 31.02 17.688 31.06 18.012 ;
      LAYER M3 ;
        RECT 30.78 17.688 30.82 18.012 ;
      LAYER M1 ;
        RECT 24.544 18.276 24.576 18.348 ;
      LAYER M2 ;
        RECT 24.524 18.296 24.596 18.328 ;
      LAYER M1 ;
        RECT 21.664 18.276 21.696 18.348 ;
      LAYER M2 ;
        RECT 21.644 18.296 21.716 18.328 ;
      LAYER M2 ;
        RECT 21.68 18.296 24.56 18.328 ;
      LAYER M3 ;
        RECT 30.78 17.976 30.82 18.48 ;
      LAYER M2 ;
        RECT 27.68 18.464 30.8 18.496 ;
      LAYER M3 ;
        RECT 27.66 18.46 27.7 18.5 ;
      LAYER M4 ;
        RECT 25.2 18.46 27.68 18.5 ;
      LAYER M5 ;
        RECT 25.168 18.312 25.232 18.48 ;
      LAYER M4 ;
        RECT 25.18 18.292 25.22 18.332 ;
      LAYER M3 ;
        RECT 25.18 18.292 25.22 18.332 ;
      LAYER M2 ;
        RECT 24.48 18.296 25.2 18.328 ;
      LAYER M3 ;
        RECT 31.02 17.872 31.06 17.912 ;
      LAYER M4 ;
        RECT 31.04 17.872 31.36 17.912 ;
      LAYER M3 ;
        RECT 31.34 16.884 31.38 17.892 ;
      LAYER M2 ;
        RECT 31.36 16.868 32.08 16.9 ;
      LAYER M3 ;
        RECT 32.06 0 32.1 16.884 ;
      LAYER M4 ;
        RECT 31.28 -0.02 32.08 0.02 ;
      LAYER M3 ;
        RECT 31.26 -0.02 31.3 0.02 ;
      LAYER M2 ;
        RECT 31.04 -0.016 31.28 0.016 ;
    END
  END vinp
  OBS 
  LAYER M2 ;
        RECT 21.404 3.26 24.676 3.292 ;
  LAYER M3 ;
        RECT 23.02 0.468 23.06 0.876 ;
  LAYER M3 ;
        RECT 22.7 0.468 22.74 0.876 ;
  LAYER M3 ;
        RECT 23.02 5.004 23.06 5.412 ;
  LAYER M3 ;
        RECT 22.7 5.004 22.74 5.412 ;
  LAYER M2 ;
        RECT 22.044 4.184 24.036 4.216 ;
  LAYER M3 ;
        RECT 23.26 4.752 23.3 5.16 ;
  LAYER M3 ;
        RECT 22.94 4.752 22.98 5.16 ;
  LAYER M3 ;
        RECT 23.1 1.56 23.14 2.472 ;
  LAYER M2 ;
        RECT 39.644 0.824 39.876 0.856 ;
  LAYER M1 ;
        RECT 34.144 16.848 34.176 16.92 ;
  LAYER M2 ;
        RECT 34.124 16.868 34.196 16.9 ;
  LAYER M1 ;
        RECT 42.784 16.848 42.816 16.92 ;
  LAYER M2 ;
        RECT 42.764 16.868 42.836 16.9 ;
  LAYER M2 ;
        RECT 34.16 16.868 42.8 16.9 ;
  LAYER M2 ;
        RECT 39.44 0.824 39.68 0.856 ;
  LAYER M3 ;
        RECT 39.42 0.84 39.46 16.212 ;
  LAYER M4 ;
        RECT 39.12 16.192 39.44 16.232 ;
  LAYER M5 ;
        RECT 39.088 16.212 39.152 16.632 ;
  LAYER M4 ;
        RECT 39.1 16.612 39.14 16.652 ;
  LAYER M3 ;
        RECT 39.1 16.632 39.14 16.884 ;
  LAYER M2 ;
        RECT 39.104 16.868 39.136 16.9 ;
  LAYER M1 ;
        RECT 27.264 5.844 27.296 5.916 ;
  LAYER M2 ;
        RECT 27.244 5.864 27.316 5.896 ;
  LAYER M1 ;
        RECT 18.624 5.844 18.656 5.916 ;
  LAYER M2 ;
        RECT 18.604 5.864 18.676 5.896 ;
  LAYER M2 ;
        RECT 18.64 5.864 27.28 5.896 ;
  LAYER M3 ;
        RECT 23.1 2.248 23.14 2.288 ;
  LAYER M4 ;
        RECT 23.12 2.248 23.28 2.288 ;
  LAYER M3 ;
        RECT 23.26 2.248 23.3 2.288 ;
  LAYER M2 ;
        RECT 23.28 2.252 24 2.284 ;
  LAYER M3 ;
        RECT 23.98 2.268 24.02 5.04 ;
  LAYER M2 ;
        RECT 24 5.024 28.8 5.056 ;
  LAYER M3 ;
        RECT 28.78 5.02 28.82 5.06 ;
  LAYER M4 ;
        RECT 28.8 5.02 39.44 5.06 ;
  LAYER M3 ;
        RECT 39.42 5.02 39.46 5.06 ;
  LAYER M3 ;
        RECT 23.98 4.872 24.02 5.88 ;
  LAYER M2 ;
        RECT 23.984 5.864 24.016 5.896 ;
  LAYER M3 ;
        RECT 23.18 1.476 23.22 2.388 ;
  LAYER M2 ;
        RECT 6.204 0.824 6.436 0.856 ;
  LAYER M1 ;
        RECT 11.904 16.848 11.936 16.92 ;
  LAYER M2 ;
        RECT 11.884 16.868 11.956 16.9 ;
  LAYER M1 ;
        RECT 3.264 16.848 3.296 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.868 3.316 16.9 ;
  LAYER M2 ;
        RECT 3.28 16.868 11.92 16.9 ;
  LAYER M2 ;
        RECT 6.4 0.824 6.64 0.856 ;
  LAYER M3 ;
        RECT 6.62 0.84 6.66 16.212 ;
  LAYER M4 ;
        RECT 6.64 16.192 6.96 16.232 ;
  LAYER M5 ;
        RECT 6.928 16.212 6.992 16.632 ;
  LAYER M4 ;
        RECT 6.94 16.612 6.98 16.652 ;
  LAYER M3 ;
        RECT 6.94 16.632 6.98 16.884 ;
  LAYER M2 ;
        RECT 6.944 16.868 6.976 16.9 ;
  LAYER M1 ;
        RECT 24.384 6.012 24.416 6.084 ;
  LAYER M2 ;
        RECT 24.364 6.032 24.436 6.064 ;
  LAYER M1 ;
        RECT 21.504 6.012 21.536 6.084 ;
  LAYER M2 ;
        RECT 21.484 6.032 21.556 6.064 ;
  LAYER M2 ;
        RECT 21.52 6.032 24.4 6.064 ;
  LAYER M3 ;
        RECT 23.18 2.352 23.22 2.856 ;
  LAYER M2 ;
        RECT 20.8 2.84 23.2 2.872 ;
  LAYER M3 ;
        RECT 20.78 2.856 20.82 5.124 ;
  LAYER M4 ;
        RECT 6.64 5.104 20.8 5.144 ;
  LAYER M3 ;
        RECT 6.62 5.104 6.66 5.144 ;
  LAYER M3 ;
        RECT 20.78 5.04 20.82 6.048 ;
  LAYER M2 ;
        RECT 20.8 6.032 21.52 6.064 ;
  LAYER M3 ;
        RECT 15.18 17.52 15.22 17.844 ;
  LAYER M3 ;
        RECT 15.42 17.52 15.46 17.844 ;
  LAYER M2 ;
        RECT 6.284 0.656 6.516 0.688 ;
  LAYER M2 ;
        RECT 7.164 0.656 7.396 0.688 ;
  LAYER M3 ;
        RECT 15.18 10.5 15.22 17.556 ;
  LAYER M2 ;
        RECT 7.28 10.484 15.2 10.516 ;
  LAYER M3 ;
        RECT 7.26 0.672 7.3 10.5 ;
  LAYER M2 ;
        RECT 7.264 0.656 7.296 0.688 ;
  LAYER M2 ;
        RECT 6.48 0.656 7.2 0.688 ;
  LAYER M3 ;
        RECT 30.86 17.52 30.9 17.844 ;
  LAYER M3 ;
        RECT 30.62 17.52 30.66 17.844 ;
  LAYER M2 ;
        RECT 39.564 0.656 39.796 0.688 ;
  LAYER M2 ;
        RECT 38.684 0.656 38.916 0.688 ;
  LAYER M3 ;
        RECT 30.86 10.5 30.9 17.556 ;
  LAYER M2 ;
        RECT 30.88 10.484 38.8 10.516 ;
  LAYER M3 ;
        RECT 38.78 0.672 38.82 10.5 ;
  LAYER M2 ;
        RECT 38.784 0.656 38.816 0.688 ;
  LAYER M2 ;
        RECT 38.88 0.656 39.6 0.688 ;
  LAYER M3 ;
        RECT 15.18 11.992 15.22 12.032 ;
  LAYER M4 ;
        RECT 15.2 11.992 15.52 12.032 ;
  LAYER M3 ;
        RECT 15.5 11.992 15.54 12.032 ;
  LAYER M2 ;
        RECT 15.52 11.996 30.88 12.028 ;
  LAYER M3 ;
        RECT 30.86 11.992 30.9 12.032 ;
  LAYER M3 ;
        RECT 5.1 0.468 5.14 0.792 ;
  LAYER M3 ;
        RECT 5.34 0.468 5.38 0.792 ;
  LAYER M2 ;
        RECT 5.804 0.572 6.036 0.604 ;
  LAYER M2 ;
        RECT 7.644 0.572 7.876 0.604 ;
  LAYER M3 ;
        RECT 5.1 0.568 5.14 0.608 ;
  LAYER M4 ;
        RECT 5.12 0.568 5.6 0.608 ;
  LAYER M3 ;
        RECT 5.58 0.568 5.62 0.608 ;
  LAYER M2 ;
        RECT 5.6 0.572 5.84 0.604 ;
  LAYER M2 ;
        RECT 6 0.572 7.68 0.604 ;
  LAYER M3 ;
        RECT 40.94 0.468 40.98 0.792 ;
  LAYER M3 ;
        RECT 40.7 0.468 40.74 0.792 ;
  LAYER M2 ;
        RECT 40.044 0.572 40.276 0.604 ;
  LAYER M2 ;
        RECT 38.204 0.572 38.436 0.604 ;
  LAYER M3 ;
        RECT 40.94 0.568 40.98 0.608 ;
  LAYER M4 ;
        RECT 40.48 0.568 40.96 0.608 ;
  LAYER M3 ;
        RECT 40.46 0.568 40.5 0.608 ;
  LAYER M2 ;
        RECT 40.24 0.572 40.48 0.604 ;
  LAYER M2 ;
        RECT 38.4 0.572 40.08 0.604 ;
  LAYER M2 ;
        RECT 7.84 0.572 20.32 0.604 ;
  LAYER M3 ;
        RECT 20.3 0.568 20.34 0.608 ;
  LAYER M4 ;
        RECT 20.32 0.568 38.24 0.608 ;
  LAYER M3 ;
        RECT 38.22 0.568 38.26 0.608 ;
  LAYER M2 ;
        RECT 38.224 0.572 38.256 0.604 ;
  LAYER M3 ;
        RECT 23.18 4.836 23.22 5.244 ;
  LAYER M3 ;
        RECT 22.86 4.836 22.9 5.244 ;
  LAYER M2 ;
        RECT 22.604 4.352 23.476 4.384 ;
  LAYER M3 ;
        RECT 22.86 4.368 22.9 4.872 ;
  LAYER M2 ;
        RECT 22.864 4.352 22.896 4.384 ;
  LAYER M3 ;
        RECT 23.1 4.92 23.14 5.328 ;
  LAYER M3 ;
        RECT 22.78 4.92 22.82 5.328 ;
  LAYER M2 ;
        RECT 21.964 4.52 24.116 4.552 ;
  LAYER M3 ;
        RECT 22.78 4.536 22.82 5.04 ;
  LAYER M2 ;
        RECT 22.784 4.52 22.816 4.552 ;
  LAYER M3 ;
        RECT 22.94 1.728 22.98 2.64 ;
  LAYER M2 ;
        RECT 21.484 3.092 24.116 3.124 ;
  LAYER M3 ;
        RECT 22.94 2.604 22.98 3.108 ;
  LAYER M2 ;
        RECT 22.944 3.092 22.976 3.124 ;
  LAYER M3 ;
        RECT 22.86 1.812 22.9 2.724 ;
  LAYER M3 ;
        RECT 23.1 0.384 23.14 0.792 ;
  LAYER M3 ;
        RECT 22.78 0.384 22.82 0.792 ;
  LAYER M3 ;
        RECT 22.86 0.924 22.9 1.932 ;
  LAYER M2 ;
        RECT 22.88 0.908 23.12 0.94 ;
  LAYER M3 ;
        RECT 23.1 0.672 23.14 0.924 ;
  LAYER M3 ;
        RECT 23.02 1.644 23.06 2.556 ;
  LAYER M2 ;
        RECT 22.124 2.924 24.756 2.956 ;
  LAYER M3 ;
        RECT 23.02 2.436 23.06 2.94 ;
  LAYER M2 ;
        RECT 23.024 2.924 23.056 2.956 ;
  LAYER M1 ;
        RECT 23.344 4.752 23.376 5.412 ;
  LAYER M1 ;
        RECT 23.424 4.752 23.456 5.412 ;
  LAYER M1 ;
        RECT 23.264 4.752 23.296 5.412 ;
  LAYER M1 ;
        RECT 22.704 4.752 22.736 5.412 ;
  LAYER M1 ;
        RECT 22.784 4.752 22.816 5.412 ;
  LAYER M1 ;
        RECT 22.624 4.752 22.656 5.412 ;
  LAYER M2 ;
        RECT 22.764 4.772 23.476 4.804 ;
  LAYER M2 ;
        RECT 22.764 5.108 23.476 5.14 ;
  LAYER M2 ;
        RECT 22.844 4.856 23.316 4.888 ;
  LAYER M2 ;
        RECT 22.844 5.192 23.316 5.224 ;
  LAYER M2 ;
        RECT 22.604 4.94 23.156 4.972 ;
  LAYER M2 ;
        RECT 22.604 5.276 23.156 5.308 ;
  LAYER M2 ;
        RECT 22.684 5.024 23.396 5.056 ;
  LAYER M2 ;
        RECT 22.684 5.36 23.396 5.392 ;
  LAYER M1 ;
        RECT 21.424 2.064 21.456 2.724 ;
  LAYER M1 ;
        RECT 21.424 1.224 21.456 1.884 ;
  LAYER M1 ;
        RECT 21.344 2.064 21.376 2.724 ;
  LAYER M1 ;
        RECT 21.344 1.224 21.376 1.884 ;
  LAYER M1 ;
        RECT 21.504 2.064 21.536 2.724 ;
  LAYER M1 ;
        RECT 21.504 1.224 21.536 1.884 ;
  LAYER M1 ;
        RECT 22.064 2.064 22.096 2.724 ;
  LAYER M1 ;
        RECT 22.064 1.224 22.096 1.884 ;
  LAYER M1 ;
        RECT 21.984 2.064 22.016 2.724 ;
  LAYER M1 ;
        RECT 21.984 1.224 22.016 1.884 ;
  LAYER M1 ;
        RECT 22.144 2.064 22.176 2.724 ;
  LAYER M1 ;
        RECT 22.144 1.224 22.176 1.884 ;
  LAYER M1 ;
        RECT 22.704 2.064 22.736 2.724 ;
  LAYER M1 ;
        RECT 22.704 1.224 22.736 1.884 ;
  LAYER M1 ;
        RECT 22.624 2.064 22.656 2.724 ;
  LAYER M1 ;
        RECT 22.624 1.224 22.656 1.884 ;
  LAYER M1 ;
        RECT 22.784 2.064 22.816 2.724 ;
  LAYER M1 ;
        RECT 22.784 1.224 22.816 1.884 ;
  LAYER M1 ;
        RECT 23.344 2.064 23.376 2.724 ;
  LAYER M1 ;
        RECT 23.344 1.224 23.376 1.884 ;
  LAYER M1 ;
        RECT 23.264 2.064 23.296 2.724 ;
  LAYER M1 ;
        RECT 23.264 1.224 23.296 1.884 ;
  LAYER M1 ;
        RECT 23.424 2.064 23.456 2.724 ;
  LAYER M1 ;
        RECT 23.424 1.224 23.456 1.884 ;
  LAYER M1 ;
        RECT 23.984 2.064 24.016 2.724 ;
  LAYER M1 ;
        RECT 23.984 1.224 24.016 1.884 ;
  LAYER M1 ;
        RECT 23.904 2.064 23.936 2.724 ;
  LAYER M1 ;
        RECT 23.904 1.224 23.936 1.884 ;
  LAYER M1 ;
        RECT 24.064 2.064 24.096 2.724 ;
  LAYER M1 ;
        RECT 24.064 1.224 24.096 1.884 ;
  LAYER M1 ;
        RECT 24.624 2.064 24.656 2.724 ;
  LAYER M1 ;
        RECT 24.624 1.224 24.656 1.884 ;
  LAYER M1 ;
        RECT 24.544 2.064 24.576 2.724 ;
  LAYER M1 ;
        RECT 24.544 1.224 24.576 1.884 ;
  LAYER M1 ;
        RECT 24.704 2.064 24.736 2.724 ;
  LAYER M1 ;
        RECT 24.704 1.224 24.736 1.884 ;
  LAYER M2 ;
        RECT 21.324 2.672 24.596 2.704 ;
  LAYER M2 ;
        RECT 21.484 2.588 24.116 2.62 ;
  LAYER M2 ;
        RECT 22.124 2.504 24.756 2.536 ;
  LAYER M2 ;
        RECT 21.404 2.42 24.036 2.452 ;
  LAYER M2 ;
        RECT 22.044 2.336 24.676 2.368 ;
  LAYER M2 ;
        RECT 21.324 1.832 24.596 1.864 ;
  LAYER M2 ;
        RECT 22.124 1.748 24.756 1.78 ;
  LAYER M2 ;
        RECT 21.484 1.664 24.116 1.696 ;
  LAYER M2 ;
        RECT 22.044 1.58 24.676 1.612 ;
  LAYER M2 ;
        RECT 21.404 1.496 24.036 1.528 ;
  LAYER M1 ;
        RECT 25.264 0.216 25.296 0.876 ;
  LAYER M1 ;
        RECT 25.344 0.216 25.376 0.876 ;
  LAYER M1 ;
        RECT 25.184 0.216 25.216 0.876 ;
  LAYER M1 ;
        RECT 24.624 0.216 24.656 0.876 ;
  LAYER M1 ;
        RECT 24.704 0.216 24.736 0.876 ;
  LAYER M1 ;
        RECT 24.544 0.216 24.576 0.876 ;
  LAYER M1 ;
        RECT 23.984 0.216 24.016 0.876 ;
  LAYER M1 ;
        RECT 24.064 0.216 24.096 0.876 ;
  LAYER M1 ;
        RECT 23.904 0.216 23.936 0.876 ;
  LAYER M1 ;
        RECT 23.344 0.216 23.376 0.876 ;
  LAYER M1 ;
        RECT 23.424 0.216 23.456 0.876 ;
  LAYER M1 ;
        RECT 23.264 0.216 23.296 0.876 ;
  LAYER M1 ;
        RECT 22.704 0.216 22.736 0.876 ;
  LAYER M1 ;
        RECT 22.784 0.216 22.816 0.876 ;
  LAYER M1 ;
        RECT 22.624 0.216 22.656 0.876 ;
  LAYER M1 ;
        RECT 22.064 0.216 22.096 0.876 ;
  LAYER M1 ;
        RECT 22.144 0.216 22.176 0.876 ;
  LAYER M1 ;
        RECT 21.984 0.216 22.016 0.876 ;
  LAYER M1 ;
        RECT 21.424 0.216 21.456 0.876 ;
  LAYER M1 ;
        RECT 21.504 0.216 21.536 0.876 ;
  LAYER M1 ;
        RECT 21.344 0.216 21.376 0.876 ;
  LAYER M1 ;
        RECT 20.784 0.216 20.816 0.876 ;
  LAYER M1 ;
        RECT 20.864 0.216 20.896 0.876 ;
  LAYER M1 ;
        RECT 20.704 0.216 20.736 0.876 ;
  LAYER M2 ;
        RECT 20.844 0.236 25.396 0.268 ;
  LAYER M2 ;
        RECT 20.844 0.572 25.396 0.604 ;
  LAYER M2 ;
        RECT 22.604 0.32 23.396 0.352 ;
  LAYER M2 ;
        RECT 22.604 0.656 23.396 0.688 ;
  LAYER M2 ;
        RECT 20.684 0.404 25.236 0.436 ;
  LAYER M2 ;
        RECT 20.684 0.74 25.236 0.772 ;
  LAYER M2 ;
        RECT 20.764 0.488 25.316 0.52 ;
  LAYER M2 ;
        RECT 20.764 0.824 25.316 0.856 ;
  LAYER M1 ;
        RECT 22.064 3.912 22.096 4.572 ;
  LAYER M1 ;
        RECT 21.984 3.912 22.016 4.572 ;
  LAYER M1 ;
        RECT 22.144 3.912 22.176 4.572 ;
  LAYER M1 ;
        RECT 22.704 3.912 22.736 4.572 ;
  LAYER M1 ;
        RECT 22.624 3.912 22.656 4.572 ;
  LAYER M1 ;
        RECT 22.784 3.912 22.816 4.572 ;
  LAYER M1 ;
        RECT 23.344 3.912 23.376 4.572 ;
  LAYER M1 ;
        RECT 23.424 3.912 23.456 4.572 ;
  LAYER M1 ;
        RECT 23.264 3.912 23.296 4.572 ;
  LAYER M1 ;
        RECT 23.984 3.912 24.016 4.572 ;
  LAYER M1 ;
        RECT 24.064 3.912 24.096 4.572 ;
  LAYER M1 ;
        RECT 23.904 3.912 23.936 4.572 ;
  LAYER M1 ;
        RECT 24.624 2.904 24.656 3.564 ;
  LAYER M1 ;
        RECT 24.704 2.904 24.736 3.564 ;
  LAYER M1 ;
        RECT 24.544 2.904 24.576 3.564 ;
  LAYER M1 ;
        RECT 23.984 2.904 24.016 3.564 ;
  LAYER M1 ;
        RECT 24.064 2.904 24.096 3.564 ;
  LAYER M1 ;
        RECT 23.904 2.904 23.936 3.564 ;
  LAYER M1 ;
        RECT 23.344 2.904 23.376 3.564 ;
  LAYER M1 ;
        RECT 23.424 2.904 23.456 3.564 ;
  LAYER M1 ;
        RECT 23.264 2.904 23.296 3.564 ;
  LAYER M1 ;
        RECT 22.704 2.904 22.736 3.564 ;
  LAYER M1 ;
        RECT 22.784 2.904 22.816 3.564 ;
  LAYER M1 ;
        RECT 22.624 2.904 22.656 3.564 ;
  LAYER M1 ;
        RECT 22.064 2.904 22.096 3.564 ;
  LAYER M1 ;
        RECT 22.144 2.904 22.176 3.564 ;
  LAYER M1 ;
        RECT 21.984 2.904 22.016 3.564 ;
  LAYER M1 ;
        RECT 21.424 2.904 21.456 3.564 ;
  LAYER M1 ;
        RECT 21.504 2.904 21.536 3.564 ;
  LAYER M1 ;
        RECT 21.344 2.904 21.376 3.564 ;
  LAYER M1 ;
        RECT 6.224 29.7 6.256 29.772 ;
  LAYER M2 ;
        RECT 6.204 29.72 6.276 29.752 ;
  LAYER M1 ;
        RECT 9.104 29.7 9.136 29.772 ;
  LAYER M2 ;
        RECT 9.084 29.72 9.156 29.752 ;
  LAYER M2 ;
        RECT 6.24 29.72 9.12 29.752 ;
  LAYER M2 ;
        RECT 5.884 0.908 6.596 0.94 ;
  LAYER M1 ;
        RECT 9.024 16.68 9.056 16.752 ;
  LAYER M2 ;
        RECT 9.004 16.7 9.076 16.732 ;
  LAYER M1 ;
        RECT 6.144 16.68 6.176 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.7 6.196 16.732 ;
  LAYER M2 ;
        RECT 6.16 16.7 9.04 16.732 ;
  LAYER M2 ;
        RECT 8.384 29.72 8.416 29.752 ;
  LAYER M3 ;
        RECT 8.38 29.484 8.42 29.736 ;
  LAYER M4 ;
        RECT 8.38 29.464 8.42 29.504 ;
  LAYER M5 ;
        RECT 8.368 16.968 8.432 29.484 ;
  LAYER M4 ;
        RECT 8.38 16.948 8.42 16.988 ;
  LAYER M3 ;
        RECT 8.38 16.716 8.42 16.968 ;
  LAYER M2 ;
        RECT 8.384 16.7 8.416 16.732 ;
  LAYER M2 ;
        RECT 6.224 16.7 6.256 16.732 ;
  LAYER M3 ;
        RECT 6.22 1.596 6.26 16.716 ;
  LAYER M4 ;
        RECT 6.22 1.576 6.26 1.616 ;
  LAYER M5 ;
        RECT 6.208 1.428 6.272 1.596 ;
  LAYER M4 ;
        RECT 6.22 1.408 6.26 1.448 ;
  LAYER M3 ;
        RECT 6.22 0.924 6.26 1.428 ;
  LAYER M2 ;
        RECT 6.224 0.908 6.256 0.94 ;
  LAYER M1 ;
        RECT 6.064 17.436 6.096 17.508 ;
  LAYER M2 ;
        RECT 6.044 17.456 6.116 17.488 ;
  LAYER M1 ;
        RECT 8.944 17.436 8.976 17.508 ;
  LAYER M2 ;
        RECT 8.924 17.456 8.996 17.488 ;
  LAYER M2 ;
        RECT 6.08 17.456 8.96 17.488 ;
  LAYER M3 ;
        RECT 5.02 0.552 5.06 0.876 ;
  LAYER M3 ;
        RECT 5.26 0.552 5.3 0.876 ;
  LAYER M3 ;
        RECT 15.1 17.604 15.14 17.928 ;
  LAYER M3 ;
        RECT 15.34 17.604 15.38 17.928 ;
  LAYER M2 ;
        RECT 8.88 17.456 15.12 17.488 ;
  LAYER M3 ;
        RECT 15.1 17.472 15.14 17.724 ;
  LAYER M2 ;
        RECT 6.064 17.456 6.096 17.488 ;
  LAYER M3 ;
        RECT 6.06 0.84 6.1 17.472 ;
  LAYER M4 ;
        RECT 5.28 0.82 6.08 0.86 ;
  LAYER M3 ;
        RECT 5.26 0.82 5.3 0.86 ;
  LAYER M2 ;
        RECT 7.084 0.908 7.796 0.94 ;
  LAYER M1 ;
        RECT 8.864 1.476 8.896 1.548 ;
  LAYER M2 ;
        RECT 8.844 1.496 8.916 1.528 ;
  LAYER M1 ;
        RECT 5.984 1.476 6.016 1.548 ;
  LAYER M2 ;
        RECT 5.964 1.496 6.036 1.528 ;
  LAYER M2 ;
        RECT 6 1.496 8.88 1.528 ;
  LAYER M2 ;
        RECT 7.664 0.908 7.696 0.94 ;
  LAYER M3 ;
        RECT 7.66 0.924 7.7 1.428 ;
  LAYER M4 ;
        RECT 7.66 1.408 7.7 1.448 ;
  LAYER M5 ;
        RECT 7.648 1.428 7.712 1.512 ;
  LAYER M4 ;
        RECT 7.66 1.492 7.7 1.532 ;
  LAYER M3 ;
        RECT 7.66 1.492 7.7 1.532 ;
  LAYER M2 ;
        RECT 7.664 1.496 7.696 1.528 ;
  LAYER M1 ;
        RECT 6.384 20.88 6.416 20.952 ;
  LAYER M2 ;
        RECT 6.364 20.9 6.436 20.932 ;
  LAYER M2 ;
        RECT 6.08 20.9 6.4 20.932 ;
  LAYER M1 ;
        RECT 6.064 20.88 6.096 20.952 ;
  LAYER M2 ;
        RECT 6.044 20.9 6.116 20.932 ;
  LAYER M1 ;
        RECT 6.384 23.82 6.416 23.892 ;
  LAYER M2 ;
        RECT 6.364 23.84 6.436 23.872 ;
  LAYER M2 ;
        RECT 6.08 23.84 6.4 23.872 ;
  LAYER M1 ;
        RECT 6.064 23.82 6.096 23.892 ;
  LAYER M2 ;
        RECT 6.044 23.84 6.116 23.872 ;
  LAYER M1 ;
        RECT 3.504 20.88 3.536 20.952 ;
  LAYER M2 ;
        RECT 3.484 20.9 3.556 20.932 ;
  LAYER M1 ;
        RECT 3.504 20.748 3.536 20.916 ;
  LAYER M1 ;
        RECT 3.504 20.712 3.536 20.784 ;
  LAYER M2 ;
        RECT 3.484 20.732 3.556 20.764 ;
  LAYER M2 ;
        RECT 3.52 20.732 6.08 20.764 ;
  LAYER M1 ;
        RECT 6.064 20.712 6.096 20.784 ;
  LAYER M2 ;
        RECT 6.044 20.732 6.116 20.764 ;
  LAYER M1 ;
        RECT 3.504 23.82 3.536 23.892 ;
  LAYER M2 ;
        RECT 3.484 23.84 3.556 23.872 ;
  LAYER M1 ;
        RECT 3.504 23.688 3.536 23.856 ;
  LAYER M1 ;
        RECT 3.504 23.652 3.536 23.724 ;
  LAYER M2 ;
        RECT 3.484 23.672 3.556 23.704 ;
  LAYER M2 ;
        RECT 3.52 23.672 6.08 23.704 ;
  LAYER M1 ;
        RECT 6.064 23.652 6.096 23.724 ;
  LAYER M2 ;
        RECT 6.044 23.672 6.116 23.704 ;
  LAYER M1 ;
        RECT 6.064 17.436 6.096 17.508 ;
  LAYER M2 ;
        RECT 6.044 17.456 6.116 17.488 ;
  LAYER M1 ;
        RECT 6.064 17.472 6.096 17.64 ;
  LAYER M1 ;
        RECT 6.064 17.64 6.096 23.856 ;
  LAYER M1 ;
        RECT 9.264 23.82 9.296 23.892 ;
  LAYER M2 ;
        RECT 9.244 23.84 9.316 23.872 ;
  LAYER M2 ;
        RECT 8.96 23.84 9.28 23.872 ;
  LAYER M1 ;
        RECT 8.944 23.82 8.976 23.892 ;
  LAYER M2 ;
        RECT 8.924 23.84 8.996 23.872 ;
  LAYER M1 ;
        RECT 9.264 20.88 9.296 20.952 ;
  LAYER M2 ;
        RECT 9.244 20.9 9.316 20.932 ;
  LAYER M2 ;
        RECT 8.96 20.9 9.28 20.932 ;
  LAYER M1 ;
        RECT 8.944 20.88 8.976 20.952 ;
  LAYER M2 ;
        RECT 8.924 20.9 8.996 20.932 ;
  LAYER M1 ;
        RECT 8.944 17.436 8.976 17.508 ;
  LAYER M2 ;
        RECT 8.924 17.456 8.996 17.488 ;
  LAYER M1 ;
        RECT 8.944 17.472 8.976 17.64 ;
  LAYER M1 ;
        RECT 8.944 17.64 8.976 23.856 ;
  LAYER M2 ;
        RECT 6.08 17.456 8.96 17.488 ;
  LAYER M1 ;
        RECT 0.624 17.94 0.656 18.012 ;
  LAYER M2 ;
        RECT 0.604 17.96 0.676 17.992 ;
  LAYER M1 ;
        RECT 0.624 17.808 0.656 17.976 ;
  LAYER M1 ;
        RECT 0.624 17.772 0.656 17.844 ;
  LAYER M2 ;
        RECT 0.604 17.792 0.676 17.824 ;
  LAYER M2 ;
        RECT 0.64 17.792 3.2 17.824 ;
  LAYER M1 ;
        RECT 3.184 17.772 3.216 17.844 ;
  LAYER M2 ;
        RECT 3.164 17.792 3.236 17.824 ;
  LAYER M1 ;
        RECT 0.624 20.88 0.656 20.952 ;
  LAYER M2 ;
        RECT 0.604 20.9 0.676 20.932 ;
  LAYER M1 ;
        RECT 0.624 20.748 0.656 20.916 ;
  LAYER M1 ;
        RECT 0.624 20.712 0.656 20.784 ;
  LAYER M2 ;
        RECT 0.604 20.732 0.676 20.764 ;
  LAYER M2 ;
        RECT 0.64 20.732 3.2 20.764 ;
  LAYER M1 ;
        RECT 3.184 20.712 3.216 20.784 ;
  LAYER M2 ;
        RECT 3.164 20.732 3.236 20.764 ;
  LAYER M1 ;
        RECT 0.624 23.82 0.656 23.892 ;
  LAYER M2 ;
        RECT 0.604 23.84 0.676 23.872 ;
  LAYER M1 ;
        RECT 0.624 23.688 0.656 23.856 ;
  LAYER M1 ;
        RECT 0.624 23.652 0.656 23.724 ;
  LAYER M2 ;
        RECT 0.604 23.672 0.676 23.704 ;
  LAYER M2 ;
        RECT 0.64 23.672 3.2 23.704 ;
  LAYER M1 ;
        RECT 3.184 23.652 3.216 23.724 ;
  LAYER M2 ;
        RECT 3.164 23.672 3.236 23.704 ;
  LAYER M1 ;
        RECT 0.624 26.76 0.656 26.832 ;
  LAYER M2 ;
        RECT 0.604 26.78 0.676 26.812 ;
  LAYER M1 ;
        RECT 0.624 26.628 0.656 26.796 ;
  LAYER M1 ;
        RECT 0.624 26.592 0.656 26.664 ;
  LAYER M2 ;
        RECT 0.604 26.612 0.676 26.644 ;
  LAYER M2 ;
        RECT 0.64 26.612 3.2 26.644 ;
  LAYER M1 ;
        RECT 3.184 26.592 3.216 26.664 ;
  LAYER M2 ;
        RECT 3.164 26.612 3.236 26.644 ;
  LAYER M1 ;
        RECT 3.504 17.94 3.536 18.012 ;
  LAYER M2 ;
        RECT 3.484 17.96 3.556 17.992 ;
  LAYER M2 ;
        RECT 3.2 17.96 3.52 17.992 ;
  LAYER M1 ;
        RECT 3.184 17.94 3.216 18.012 ;
  LAYER M2 ;
        RECT 3.164 17.96 3.236 17.992 ;
  LAYER M1 ;
        RECT 3.504 26.76 3.536 26.832 ;
  LAYER M2 ;
        RECT 3.484 26.78 3.556 26.812 ;
  LAYER M2 ;
        RECT 3.2 26.78 3.52 26.812 ;
  LAYER M1 ;
        RECT 3.184 26.76 3.216 26.832 ;
  LAYER M2 ;
        RECT 3.164 26.78 3.236 26.812 ;
  LAYER M1 ;
        RECT 3.184 17.268 3.216 17.34 ;
  LAYER M2 ;
        RECT 3.164 17.288 3.236 17.32 ;
  LAYER M1 ;
        RECT 3.184 17.304 3.216 17.64 ;
  LAYER M1 ;
        RECT 3.184 17.64 3.216 26.796 ;
  LAYER M1 ;
        RECT 9.264 17.94 9.296 18.012 ;
  LAYER M2 ;
        RECT 9.244 17.96 9.316 17.992 ;
  LAYER M1 ;
        RECT 9.264 17.808 9.296 17.976 ;
  LAYER M1 ;
        RECT 9.264 17.772 9.296 17.844 ;
  LAYER M2 ;
        RECT 9.244 17.792 9.316 17.824 ;
  LAYER M2 ;
        RECT 9.28 17.792 11.84 17.824 ;
  LAYER M1 ;
        RECT 11.824 17.772 11.856 17.844 ;
  LAYER M2 ;
        RECT 11.804 17.792 11.876 17.824 ;
  LAYER M1 ;
        RECT 9.264 26.76 9.296 26.832 ;
  LAYER M2 ;
        RECT 9.244 26.78 9.316 26.812 ;
  LAYER M1 ;
        RECT 9.264 26.628 9.296 26.796 ;
  LAYER M1 ;
        RECT 9.264 26.592 9.296 26.664 ;
  LAYER M2 ;
        RECT 9.244 26.612 9.316 26.644 ;
  LAYER M2 ;
        RECT 9.28 26.612 11.84 26.644 ;
  LAYER M1 ;
        RECT 11.824 26.592 11.856 26.664 ;
  LAYER M2 ;
        RECT 11.804 26.612 11.876 26.644 ;
  LAYER M1 ;
        RECT 12.144 17.94 12.176 18.012 ;
  LAYER M2 ;
        RECT 12.124 17.96 12.196 17.992 ;
  LAYER M2 ;
        RECT 11.84 17.96 12.16 17.992 ;
  LAYER M1 ;
        RECT 11.824 17.94 11.856 18.012 ;
  LAYER M2 ;
        RECT 11.804 17.96 11.876 17.992 ;
  LAYER M1 ;
        RECT 12.144 20.88 12.176 20.952 ;
  LAYER M2 ;
        RECT 12.124 20.9 12.196 20.932 ;
  LAYER M2 ;
        RECT 11.84 20.9 12.16 20.932 ;
  LAYER M1 ;
        RECT 11.824 20.88 11.856 20.952 ;
  LAYER M2 ;
        RECT 11.804 20.9 11.876 20.932 ;
  LAYER M1 ;
        RECT 12.144 23.82 12.176 23.892 ;
  LAYER M2 ;
        RECT 12.124 23.84 12.196 23.872 ;
  LAYER M2 ;
        RECT 11.84 23.84 12.16 23.872 ;
  LAYER M1 ;
        RECT 11.824 23.82 11.856 23.892 ;
  LAYER M2 ;
        RECT 11.804 23.84 11.876 23.872 ;
  LAYER M1 ;
        RECT 12.144 26.76 12.176 26.832 ;
  LAYER M2 ;
        RECT 12.124 26.78 12.196 26.812 ;
  LAYER M2 ;
        RECT 11.84 26.78 12.16 26.812 ;
  LAYER M1 ;
        RECT 11.824 26.76 11.856 26.832 ;
  LAYER M2 ;
        RECT 11.804 26.78 11.876 26.812 ;
  LAYER M1 ;
        RECT 11.824 17.268 11.856 17.34 ;
  LAYER M2 ;
        RECT 11.804 17.288 11.876 17.32 ;
  LAYER M1 ;
        RECT 11.824 17.304 11.856 17.64 ;
  LAYER M1 ;
        RECT 11.824 17.64 11.856 26.796 ;
  LAYER M2 ;
        RECT 3.2 17.288 11.84 17.32 ;
  LAYER M1 ;
        RECT 6.384 26.76 6.416 26.832 ;
  LAYER M2 ;
        RECT 6.364 26.78 6.436 26.812 ;
  LAYER M2 ;
        RECT 3.52 26.78 6.4 26.812 ;
  LAYER M1 ;
        RECT 3.504 26.76 3.536 26.832 ;
  LAYER M2 ;
        RECT 3.484 26.78 3.556 26.812 ;
  LAYER M1 ;
        RECT 6.384 17.94 6.416 18.012 ;
  LAYER M2 ;
        RECT 6.364 17.96 6.436 17.992 ;
  LAYER M2 ;
        RECT 6.4 17.96 9.28 17.992 ;
  LAYER M1 ;
        RECT 9.264 17.94 9.296 18.012 ;
  LAYER M2 ;
        RECT 9.244 17.96 9.316 17.992 ;
  LAYER M1 ;
        RECT 8.784 23.316 8.816 23.388 ;
  LAYER M2 ;
        RECT 8.764 23.336 8.836 23.368 ;
  LAYER M2 ;
        RECT 6.24 23.336 8.8 23.368 ;
  LAYER M1 ;
        RECT 6.224 23.316 6.256 23.388 ;
  LAYER M2 ;
        RECT 6.204 23.336 6.276 23.368 ;
  LAYER M1 ;
        RECT 8.784 26.256 8.816 26.328 ;
  LAYER M2 ;
        RECT 8.764 26.276 8.836 26.308 ;
  LAYER M2 ;
        RECT 6.24 26.276 8.8 26.308 ;
  LAYER M1 ;
        RECT 6.224 26.256 6.256 26.328 ;
  LAYER M2 ;
        RECT 6.204 26.276 6.276 26.308 ;
  LAYER M1 ;
        RECT 5.904 23.316 5.936 23.388 ;
  LAYER M2 ;
        RECT 5.884 23.336 5.956 23.368 ;
  LAYER M1 ;
        RECT 5.904 23.352 5.936 23.52 ;
  LAYER M1 ;
        RECT 5.904 23.484 5.936 23.556 ;
  LAYER M2 ;
        RECT 5.884 23.504 5.956 23.536 ;
  LAYER M2 ;
        RECT 5.92 23.504 6.24 23.536 ;
  LAYER M1 ;
        RECT 6.224 23.484 6.256 23.556 ;
  LAYER M2 ;
        RECT 6.204 23.504 6.276 23.536 ;
  LAYER M1 ;
        RECT 5.904 26.256 5.936 26.328 ;
  LAYER M2 ;
        RECT 5.884 26.276 5.956 26.308 ;
  LAYER M1 ;
        RECT 5.904 26.292 5.936 26.46 ;
  LAYER M1 ;
        RECT 5.904 26.424 5.936 26.496 ;
  LAYER M2 ;
        RECT 5.884 26.444 5.956 26.476 ;
  LAYER M2 ;
        RECT 5.92 26.444 6.24 26.476 ;
  LAYER M1 ;
        RECT 6.224 26.424 6.256 26.496 ;
  LAYER M2 ;
        RECT 6.204 26.444 6.276 26.476 ;
  LAYER M1 ;
        RECT 6.224 29.7 6.256 29.772 ;
  LAYER M2 ;
        RECT 6.204 29.72 6.276 29.752 ;
  LAYER M1 ;
        RECT 6.224 29.568 6.256 29.736 ;
  LAYER M1 ;
        RECT 6.224 23.352 6.256 29.568 ;
  LAYER M1 ;
        RECT 11.664 26.256 11.696 26.328 ;
  LAYER M2 ;
        RECT 11.644 26.276 11.716 26.308 ;
  LAYER M2 ;
        RECT 9.12 26.276 11.68 26.308 ;
  LAYER M1 ;
        RECT 9.104 26.256 9.136 26.328 ;
  LAYER M2 ;
        RECT 9.084 26.276 9.156 26.308 ;
  LAYER M1 ;
        RECT 11.664 23.316 11.696 23.388 ;
  LAYER M2 ;
        RECT 11.644 23.336 11.716 23.368 ;
  LAYER M2 ;
        RECT 9.12 23.336 11.68 23.368 ;
  LAYER M1 ;
        RECT 9.104 23.316 9.136 23.388 ;
  LAYER M2 ;
        RECT 9.084 23.336 9.156 23.368 ;
  LAYER M1 ;
        RECT 9.104 29.7 9.136 29.772 ;
  LAYER M2 ;
        RECT 9.084 29.72 9.156 29.752 ;
  LAYER M1 ;
        RECT 9.104 29.568 9.136 29.736 ;
  LAYER M1 ;
        RECT 9.104 23.352 9.136 29.568 ;
  LAYER M2 ;
        RECT 6.24 29.72 9.12 29.752 ;
  LAYER M1 ;
        RECT 3.024 20.376 3.056 20.448 ;
  LAYER M2 ;
        RECT 3.004 20.396 3.076 20.428 ;
  LAYER M2 ;
        RECT 0.32 20.396 3.04 20.428 ;
  LAYER M1 ;
        RECT 0.304 20.376 0.336 20.448 ;
  LAYER M2 ;
        RECT 0.284 20.396 0.356 20.428 ;
  LAYER M1 ;
        RECT 3.024 23.316 3.056 23.388 ;
  LAYER M2 ;
        RECT 3.004 23.336 3.076 23.368 ;
  LAYER M2 ;
        RECT 0.32 23.336 3.04 23.368 ;
  LAYER M1 ;
        RECT 0.304 23.316 0.336 23.388 ;
  LAYER M2 ;
        RECT 0.284 23.336 0.356 23.368 ;
  LAYER M1 ;
        RECT 3.024 26.256 3.056 26.328 ;
  LAYER M2 ;
        RECT 3.004 26.276 3.076 26.308 ;
  LAYER M2 ;
        RECT 0.32 26.276 3.04 26.308 ;
  LAYER M1 ;
        RECT 0.304 26.256 0.336 26.328 ;
  LAYER M2 ;
        RECT 0.284 26.276 0.356 26.308 ;
  LAYER M1 ;
        RECT 3.024 29.196 3.056 29.268 ;
  LAYER M2 ;
        RECT 3.004 29.216 3.076 29.248 ;
  LAYER M2 ;
        RECT 0.32 29.216 3.04 29.248 ;
  LAYER M1 ;
        RECT 0.304 29.196 0.336 29.268 ;
  LAYER M2 ;
        RECT 0.284 29.216 0.356 29.248 ;
  LAYER M1 ;
        RECT 0.304 29.868 0.336 29.94 ;
  LAYER M2 ;
        RECT 0.284 29.888 0.356 29.92 ;
  LAYER M1 ;
        RECT 0.304 29.568 0.336 29.904 ;
  LAYER M1 ;
        RECT 0.304 20.412 0.336 29.568 ;
  LAYER M1 ;
        RECT 14.544 20.376 14.576 20.448 ;
  LAYER M2 ;
        RECT 14.524 20.396 14.596 20.428 ;
  LAYER M1 ;
        RECT 14.544 20.412 14.576 20.58 ;
  LAYER M1 ;
        RECT 14.544 20.544 14.576 20.616 ;
  LAYER M2 ;
        RECT 14.524 20.564 14.596 20.596 ;
  LAYER M2 ;
        RECT 14.56 20.564 14.72 20.596 ;
  LAYER M1 ;
        RECT 14.704 20.544 14.736 20.616 ;
  LAYER M2 ;
        RECT 14.684 20.564 14.756 20.596 ;
  LAYER M1 ;
        RECT 14.544 23.316 14.576 23.388 ;
  LAYER M2 ;
        RECT 14.524 23.336 14.596 23.368 ;
  LAYER M1 ;
        RECT 14.544 23.352 14.576 23.52 ;
  LAYER M1 ;
        RECT 14.544 23.484 14.576 23.556 ;
  LAYER M2 ;
        RECT 14.524 23.504 14.596 23.536 ;
  LAYER M2 ;
        RECT 14.56 23.504 14.72 23.536 ;
  LAYER M1 ;
        RECT 14.704 23.484 14.736 23.556 ;
  LAYER M2 ;
        RECT 14.684 23.504 14.756 23.536 ;
  LAYER M1 ;
        RECT 14.544 26.256 14.576 26.328 ;
  LAYER M2 ;
        RECT 14.524 26.276 14.596 26.308 ;
  LAYER M1 ;
        RECT 14.544 26.292 14.576 26.46 ;
  LAYER M1 ;
        RECT 14.544 26.424 14.576 26.496 ;
  LAYER M2 ;
        RECT 14.524 26.444 14.596 26.476 ;
  LAYER M2 ;
        RECT 14.56 26.444 14.72 26.476 ;
  LAYER M1 ;
        RECT 14.704 26.424 14.736 26.496 ;
  LAYER M2 ;
        RECT 14.684 26.444 14.756 26.476 ;
  LAYER M1 ;
        RECT 14.544 29.196 14.576 29.268 ;
  LAYER M2 ;
        RECT 14.524 29.216 14.596 29.248 ;
  LAYER M1 ;
        RECT 14.544 29.232 14.576 29.4 ;
  LAYER M1 ;
        RECT 14.544 29.364 14.576 29.436 ;
  LAYER M2 ;
        RECT 14.524 29.384 14.596 29.416 ;
  LAYER M2 ;
        RECT 14.56 29.384 14.72 29.416 ;
  LAYER M1 ;
        RECT 14.704 29.364 14.736 29.436 ;
  LAYER M2 ;
        RECT 14.684 29.384 14.756 29.416 ;
  LAYER M1 ;
        RECT 14.704 29.868 14.736 29.94 ;
  LAYER M2 ;
        RECT 14.684 29.888 14.756 29.92 ;
  LAYER M1 ;
        RECT 14.704 29.568 14.736 29.904 ;
  LAYER M1 ;
        RECT 14.704 20.58 14.736 29.568 ;
  LAYER M2 ;
        RECT 0.32 29.888 14.72 29.92 ;
  LAYER M1 ;
        RECT 5.904 20.376 5.936 20.448 ;
  LAYER M2 ;
        RECT 5.884 20.396 5.956 20.428 ;
  LAYER M2 ;
        RECT 3.04 20.396 5.92 20.428 ;
  LAYER M1 ;
        RECT 3.024 20.376 3.056 20.448 ;
  LAYER M2 ;
        RECT 3.004 20.396 3.076 20.428 ;
  LAYER M1 ;
        RECT 5.904 29.196 5.936 29.268 ;
  LAYER M2 ;
        RECT 5.884 29.216 5.956 29.248 ;
  LAYER M2 ;
        RECT 3.04 29.216 5.92 29.248 ;
  LAYER M1 ;
        RECT 3.024 29.196 3.056 29.268 ;
  LAYER M2 ;
        RECT 3.004 29.216 3.076 29.248 ;
  LAYER M1 ;
        RECT 8.784 29.196 8.816 29.268 ;
  LAYER M2 ;
        RECT 8.764 29.216 8.836 29.248 ;
  LAYER M2 ;
        RECT 5.92 29.216 8.8 29.248 ;
  LAYER M1 ;
        RECT 5.904 29.196 5.936 29.268 ;
  LAYER M2 ;
        RECT 5.884 29.216 5.956 29.248 ;
  LAYER M1 ;
        RECT 11.664 29.196 11.696 29.268 ;
  LAYER M2 ;
        RECT 11.644 29.216 11.716 29.248 ;
  LAYER M2 ;
        RECT 8.8 29.216 11.68 29.248 ;
  LAYER M1 ;
        RECT 8.784 29.196 8.816 29.268 ;
  LAYER M2 ;
        RECT 8.764 29.216 8.836 29.248 ;
  LAYER M1 ;
        RECT 11.664 20.376 11.696 20.448 ;
  LAYER M2 ;
        RECT 11.644 20.396 11.716 20.428 ;
  LAYER M2 ;
        RECT 11.68 20.396 14.56 20.428 ;
  LAYER M1 ;
        RECT 14.544 20.376 14.576 20.448 ;
  LAYER M2 ;
        RECT 14.524 20.396 14.596 20.428 ;
  LAYER M1 ;
        RECT 8.784 20.376 8.816 20.448 ;
  LAYER M2 ;
        RECT 8.764 20.396 8.836 20.428 ;
  LAYER M2 ;
        RECT 8.8 20.396 11.68 20.428 ;
  LAYER M1 ;
        RECT 11.664 20.376 11.696 20.448 ;
  LAYER M2 ;
        RECT 11.644 20.396 11.716 20.428 ;
  LAYER M1 ;
        RECT 0.624 17.94 0.656 20.448 ;
  LAYER M1 ;
        RECT 0.688 17.94 0.72 20.448 ;
  LAYER M1 ;
        RECT 0.752 17.94 0.784 20.448 ;
  LAYER M1 ;
        RECT 0.816 17.94 0.848 20.448 ;
  LAYER M1 ;
        RECT 0.88 17.94 0.912 20.448 ;
  LAYER M1 ;
        RECT 0.944 17.94 0.976 20.448 ;
  LAYER M1 ;
        RECT 1.008 17.94 1.04 20.448 ;
  LAYER M1 ;
        RECT 1.072 17.94 1.104 20.448 ;
  LAYER M1 ;
        RECT 1.136 17.94 1.168 20.448 ;
  LAYER M1 ;
        RECT 1.2 17.94 1.232 20.448 ;
  LAYER M1 ;
        RECT 1.264 17.94 1.296 20.448 ;
  LAYER M1 ;
        RECT 1.328 17.94 1.36 20.448 ;
  LAYER M1 ;
        RECT 1.392 17.94 1.424 20.448 ;
  LAYER M1 ;
        RECT 1.456 17.94 1.488 20.448 ;
  LAYER M1 ;
        RECT 1.52 17.94 1.552 20.448 ;
  LAYER M1 ;
        RECT 1.584 17.94 1.616 20.448 ;
  LAYER M1 ;
        RECT 1.648 17.94 1.68 20.448 ;
  LAYER M1 ;
        RECT 1.712 17.94 1.744 20.448 ;
  LAYER M1 ;
        RECT 1.776 17.94 1.808 20.448 ;
  LAYER M1 ;
        RECT 1.84 17.94 1.872 20.448 ;
  LAYER M1 ;
        RECT 1.904 17.94 1.936 20.448 ;
  LAYER M1 ;
        RECT 1.968 17.94 2 20.448 ;
  LAYER M1 ;
        RECT 2.032 17.94 2.064 20.448 ;
  LAYER M1 ;
        RECT 2.096 17.94 2.128 20.448 ;
  LAYER M1 ;
        RECT 2.16 17.94 2.192 20.448 ;
  LAYER M1 ;
        RECT 2.224 17.94 2.256 20.448 ;
  LAYER M1 ;
        RECT 2.288 17.94 2.32 20.448 ;
  LAYER M1 ;
        RECT 2.352 17.94 2.384 20.448 ;
  LAYER M1 ;
        RECT 2.416 17.94 2.448 20.448 ;
  LAYER M1 ;
        RECT 2.48 17.94 2.512 20.448 ;
  LAYER M1 ;
        RECT 2.544 17.94 2.576 20.448 ;
  LAYER M1 ;
        RECT 2.608 17.94 2.64 20.448 ;
  LAYER M1 ;
        RECT 2.672 17.94 2.704 20.448 ;
  LAYER M1 ;
        RECT 2.736 17.94 2.768 20.448 ;
  LAYER M1 ;
        RECT 2.8 17.94 2.832 20.448 ;
  LAYER M1 ;
        RECT 2.864 17.94 2.896 20.448 ;
  LAYER M1 ;
        RECT 2.928 17.94 2.96 20.448 ;
  LAYER M2 ;
        RECT 0.604 18.024 3.076 18.056 ;
  LAYER M2 ;
        RECT 0.604 18.088 3.076 18.12 ;
  LAYER M2 ;
        RECT 0.604 18.152 3.076 18.184 ;
  LAYER M2 ;
        RECT 0.604 18.216 3.076 18.248 ;
  LAYER M2 ;
        RECT 0.604 18.28 3.076 18.312 ;
  LAYER M2 ;
        RECT 0.604 18.344 3.076 18.376 ;
  LAYER M2 ;
        RECT 0.604 18.408 3.076 18.44 ;
  LAYER M2 ;
        RECT 0.604 18.472 3.076 18.504 ;
  LAYER M2 ;
        RECT 0.604 18.536 3.076 18.568 ;
  LAYER M2 ;
        RECT 0.604 18.6 3.076 18.632 ;
  LAYER M2 ;
        RECT 0.604 18.664 3.076 18.696 ;
  LAYER M2 ;
        RECT 0.604 18.728 3.076 18.76 ;
  LAYER M2 ;
        RECT 0.604 18.792 3.076 18.824 ;
  LAYER M2 ;
        RECT 0.604 18.856 3.076 18.888 ;
  LAYER M2 ;
        RECT 0.604 18.92 3.076 18.952 ;
  LAYER M2 ;
        RECT 0.604 18.984 3.076 19.016 ;
  LAYER M2 ;
        RECT 0.604 19.048 3.076 19.08 ;
  LAYER M2 ;
        RECT 0.604 19.112 3.076 19.144 ;
  LAYER M2 ;
        RECT 0.604 19.176 3.076 19.208 ;
  LAYER M2 ;
        RECT 0.604 19.24 3.076 19.272 ;
  LAYER M2 ;
        RECT 0.604 19.304 3.076 19.336 ;
  LAYER M2 ;
        RECT 0.604 19.368 3.076 19.4 ;
  LAYER M2 ;
        RECT 0.604 19.432 3.076 19.464 ;
  LAYER M2 ;
        RECT 0.604 19.496 3.076 19.528 ;
  LAYER M2 ;
        RECT 0.604 19.56 3.076 19.592 ;
  LAYER M2 ;
        RECT 0.604 19.624 3.076 19.656 ;
  LAYER M2 ;
        RECT 0.604 19.688 3.076 19.72 ;
  LAYER M2 ;
        RECT 0.604 19.752 3.076 19.784 ;
  LAYER M2 ;
        RECT 0.604 19.816 3.076 19.848 ;
  LAYER M2 ;
        RECT 0.604 19.88 3.076 19.912 ;
  LAYER M2 ;
        RECT 0.604 19.944 3.076 19.976 ;
  LAYER M2 ;
        RECT 0.604 20.008 3.076 20.04 ;
  LAYER M2 ;
        RECT 0.604 20.072 3.076 20.104 ;
  LAYER M2 ;
        RECT 0.604 20.136 3.076 20.168 ;
  LAYER M2 ;
        RECT 0.604 20.2 3.076 20.232 ;
  LAYER M2 ;
        RECT 0.604 20.264 3.076 20.296 ;
  LAYER M3 ;
        RECT 0.624 17.94 0.656 20.448 ;
  LAYER M3 ;
        RECT 0.688 17.94 0.72 20.448 ;
  LAYER M3 ;
        RECT 0.752 17.94 0.784 20.448 ;
  LAYER M3 ;
        RECT 0.816 17.94 0.848 20.448 ;
  LAYER M3 ;
        RECT 0.88 17.94 0.912 20.448 ;
  LAYER M3 ;
        RECT 0.944 17.94 0.976 20.448 ;
  LAYER M3 ;
        RECT 1.008 17.94 1.04 20.448 ;
  LAYER M3 ;
        RECT 1.072 17.94 1.104 20.448 ;
  LAYER M3 ;
        RECT 1.136 17.94 1.168 20.448 ;
  LAYER M3 ;
        RECT 1.2 17.94 1.232 20.448 ;
  LAYER M3 ;
        RECT 1.264 17.94 1.296 20.448 ;
  LAYER M3 ;
        RECT 1.328 17.94 1.36 20.448 ;
  LAYER M3 ;
        RECT 1.392 17.94 1.424 20.448 ;
  LAYER M3 ;
        RECT 1.456 17.94 1.488 20.448 ;
  LAYER M3 ;
        RECT 1.52 17.94 1.552 20.448 ;
  LAYER M3 ;
        RECT 1.584 17.94 1.616 20.448 ;
  LAYER M3 ;
        RECT 1.648 17.94 1.68 20.448 ;
  LAYER M3 ;
        RECT 1.712 17.94 1.744 20.448 ;
  LAYER M3 ;
        RECT 1.776 17.94 1.808 20.448 ;
  LAYER M3 ;
        RECT 1.84 17.94 1.872 20.448 ;
  LAYER M3 ;
        RECT 1.904 17.94 1.936 20.448 ;
  LAYER M3 ;
        RECT 1.968 17.94 2 20.448 ;
  LAYER M3 ;
        RECT 2.032 17.94 2.064 20.448 ;
  LAYER M3 ;
        RECT 2.096 17.94 2.128 20.448 ;
  LAYER M3 ;
        RECT 2.16 17.94 2.192 20.448 ;
  LAYER M3 ;
        RECT 2.224 17.94 2.256 20.448 ;
  LAYER M3 ;
        RECT 2.288 17.94 2.32 20.448 ;
  LAYER M3 ;
        RECT 2.352 17.94 2.384 20.448 ;
  LAYER M3 ;
        RECT 2.416 17.94 2.448 20.448 ;
  LAYER M3 ;
        RECT 2.48 17.94 2.512 20.448 ;
  LAYER M3 ;
        RECT 2.544 17.94 2.576 20.448 ;
  LAYER M3 ;
        RECT 2.608 17.94 2.64 20.448 ;
  LAYER M3 ;
        RECT 2.672 17.94 2.704 20.448 ;
  LAYER M3 ;
        RECT 2.736 17.94 2.768 20.448 ;
  LAYER M3 ;
        RECT 2.8 17.94 2.832 20.448 ;
  LAYER M3 ;
        RECT 2.864 17.94 2.896 20.448 ;
  LAYER M3 ;
        RECT 2.928 17.94 2.96 20.448 ;
  LAYER M3 ;
        RECT 3.024 17.94 3.056 20.448 ;
  LAYER M1 ;
        RECT 0.639 17.976 0.641 20.412 ;
  LAYER M1 ;
        RECT 0.719 17.976 0.721 20.412 ;
  LAYER M1 ;
        RECT 0.799 17.976 0.801 20.412 ;
  LAYER M1 ;
        RECT 0.879 17.976 0.881 20.412 ;
  LAYER M1 ;
        RECT 0.959 17.976 0.961 20.412 ;
  LAYER M1 ;
        RECT 1.039 17.976 1.041 20.412 ;
  LAYER M1 ;
        RECT 1.119 17.976 1.121 20.412 ;
  LAYER M1 ;
        RECT 1.199 17.976 1.201 20.412 ;
  LAYER M1 ;
        RECT 1.279 17.976 1.281 20.412 ;
  LAYER M1 ;
        RECT 1.359 17.976 1.361 20.412 ;
  LAYER M1 ;
        RECT 1.439 17.976 1.441 20.412 ;
  LAYER M1 ;
        RECT 1.519 17.976 1.521 20.412 ;
  LAYER M1 ;
        RECT 1.599 17.976 1.601 20.412 ;
  LAYER M1 ;
        RECT 1.679 17.976 1.681 20.412 ;
  LAYER M1 ;
        RECT 1.759 17.976 1.761 20.412 ;
  LAYER M1 ;
        RECT 1.839 17.976 1.841 20.412 ;
  LAYER M1 ;
        RECT 1.919 17.976 1.921 20.412 ;
  LAYER M1 ;
        RECT 1.999 17.976 2.001 20.412 ;
  LAYER M1 ;
        RECT 2.079 17.976 2.081 20.412 ;
  LAYER M1 ;
        RECT 2.159 17.976 2.161 20.412 ;
  LAYER M1 ;
        RECT 2.239 17.976 2.241 20.412 ;
  LAYER M1 ;
        RECT 2.319 17.976 2.321 20.412 ;
  LAYER M1 ;
        RECT 2.399 17.976 2.401 20.412 ;
  LAYER M1 ;
        RECT 2.479 17.976 2.481 20.412 ;
  LAYER M1 ;
        RECT 2.559 17.976 2.561 20.412 ;
  LAYER M1 ;
        RECT 2.639 17.976 2.641 20.412 ;
  LAYER M1 ;
        RECT 2.719 17.976 2.721 20.412 ;
  LAYER M1 ;
        RECT 2.799 17.976 2.801 20.412 ;
  LAYER M1 ;
        RECT 2.879 17.976 2.881 20.412 ;
  LAYER M1 ;
        RECT 2.959 17.976 2.961 20.412 ;
  LAYER M2 ;
        RECT 0.64 17.975 3.04 17.977 ;
  LAYER M2 ;
        RECT 0.64 18.059 3.04 18.061 ;
  LAYER M2 ;
        RECT 0.64 18.143 3.04 18.145 ;
  LAYER M2 ;
        RECT 0.64 18.227 3.04 18.229 ;
  LAYER M2 ;
        RECT 0.64 18.311 3.04 18.313 ;
  LAYER M2 ;
        RECT 0.64 18.395 3.04 18.397 ;
  LAYER M2 ;
        RECT 0.64 18.479 3.04 18.481 ;
  LAYER M2 ;
        RECT 0.64 18.563 3.04 18.565 ;
  LAYER M2 ;
        RECT 0.64 18.647 3.04 18.649 ;
  LAYER M2 ;
        RECT 0.64 18.731 3.04 18.733 ;
  LAYER M2 ;
        RECT 0.64 18.815 3.04 18.817 ;
  LAYER M2 ;
        RECT 0.64 18.899 3.04 18.901 ;
  LAYER M2 ;
        RECT 0.64 18.9825 3.04 18.9845 ;
  LAYER M2 ;
        RECT 0.64 19.067 3.04 19.069 ;
  LAYER M2 ;
        RECT 0.64 19.151 3.04 19.153 ;
  LAYER M2 ;
        RECT 0.64 19.235 3.04 19.237 ;
  LAYER M2 ;
        RECT 0.64 19.319 3.04 19.321 ;
  LAYER M2 ;
        RECT 0.64 19.403 3.04 19.405 ;
  LAYER M2 ;
        RECT 0.64 19.487 3.04 19.489 ;
  LAYER M2 ;
        RECT 0.64 19.571 3.04 19.573 ;
  LAYER M2 ;
        RECT 0.64 19.655 3.04 19.657 ;
  LAYER M2 ;
        RECT 0.64 19.739 3.04 19.741 ;
  LAYER M2 ;
        RECT 0.64 19.823 3.04 19.825 ;
  LAYER M2 ;
        RECT 0.64 19.907 3.04 19.909 ;
  LAYER M2 ;
        RECT 0.64 19.991 3.04 19.993 ;
  LAYER M2 ;
        RECT 0.64 20.075 3.04 20.077 ;
  LAYER M2 ;
        RECT 0.64 20.159 3.04 20.161 ;
  LAYER M2 ;
        RECT 0.64 20.243 3.04 20.245 ;
  LAYER M2 ;
        RECT 0.64 20.327 3.04 20.329 ;
  LAYER M1 ;
        RECT 0.624 20.88 0.656 23.388 ;
  LAYER M1 ;
        RECT 0.688 20.88 0.72 23.388 ;
  LAYER M1 ;
        RECT 0.752 20.88 0.784 23.388 ;
  LAYER M1 ;
        RECT 0.816 20.88 0.848 23.388 ;
  LAYER M1 ;
        RECT 0.88 20.88 0.912 23.388 ;
  LAYER M1 ;
        RECT 0.944 20.88 0.976 23.388 ;
  LAYER M1 ;
        RECT 1.008 20.88 1.04 23.388 ;
  LAYER M1 ;
        RECT 1.072 20.88 1.104 23.388 ;
  LAYER M1 ;
        RECT 1.136 20.88 1.168 23.388 ;
  LAYER M1 ;
        RECT 1.2 20.88 1.232 23.388 ;
  LAYER M1 ;
        RECT 1.264 20.88 1.296 23.388 ;
  LAYER M1 ;
        RECT 1.328 20.88 1.36 23.388 ;
  LAYER M1 ;
        RECT 1.392 20.88 1.424 23.388 ;
  LAYER M1 ;
        RECT 1.456 20.88 1.488 23.388 ;
  LAYER M1 ;
        RECT 1.52 20.88 1.552 23.388 ;
  LAYER M1 ;
        RECT 1.584 20.88 1.616 23.388 ;
  LAYER M1 ;
        RECT 1.648 20.88 1.68 23.388 ;
  LAYER M1 ;
        RECT 1.712 20.88 1.744 23.388 ;
  LAYER M1 ;
        RECT 1.776 20.88 1.808 23.388 ;
  LAYER M1 ;
        RECT 1.84 20.88 1.872 23.388 ;
  LAYER M1 ;
        RECT 1.904 20.88 1.936 23.388 ;
  LAYER M1 ;
        RECT 1.968 20.88 2 23.388 ;
  LAYER M1 ;
        RECT 2.032 20.88 2.064 23.388 ;
  LAYER M1 ;
        RECT 2.096 20.88 2.128 23.388 ;
  LAYER M1 ;
        RECT 2.16 20.88 2.192 23.388 ;
  LAYER M1 ;
        RECT 2.224 20.88 2.256 23.388 ;
  LAYER M1 ;
        RECT 2.288 20.88 2.32 23.388 ;
  LAYER M1 ;
        RECT 2.352 20.88 2.384 23.388 ;
  LAYER M1 ;
        RECT 2.416 20.88 2.448 23.388 ;
  LAYER M1 ;
        RECT 2.48 20.88 2.512 23.388 ;
  LAYER M1 ;
        RECT 2.544 20.88 2.576 23.388 ;
  LAYER M1 ;
        RECT 2.608 20.88 2.64 23.388 ;
  LAYER M1 ;
        RECT 2.672 20.88 2.704 23.388 ;
  LAYER M1 ;
        RECT 2.736 20.88 2.768 23.388 ;
  LAYER M1 ;
        RECT 2.8 20.88 2.832 23.388 ;
  LAYER M1 ;
        RECT 2.864 20.88 2.896 23.388 ;
  LAYER M1 ;
        RECT 2.928 20.88 2.96 23.388 ;
  LAYER M2 ;
        RECT 0.604 20.964 3.076 20.996 ;
  LAYER M2 ;
        RECT 0.604 21.028 3.076 21.06 ;
  LAYER M2 ;
        RECT 0.604 21.092 3.076 21.124 ;
  LAYER M2 ;
        RECT 0.604 21.156 3.076 21.188 ;
  LAYER M2 ;
        RECT 0.604 21.22 3.076 21.252 ;
  LAYER M2 ;
        RECT 0.604 21.284 3.076 21.316 ;
  LAYER M2 ;
        RECT 0.604 21.348 3.076 21.38 ;
  LAYER M2 ;
        RECT 0.604 21.412 3.076 21.444 ;
  LAYER M2 ;
        RECT 0.604 21.476 3.076 21.508 ;
  LAYER M2 ;
        RECT 0.604 21.54 3.076 21.572 ;
  LAYER M2 ;
        RECT 0.604 21.604 3.076 21.636 ;
  LAYER M2 ;
        RECT 0.604 21.668 3.076 21.7 ;
  LAYER M2 ;
        RECT 0.604 21.732 3.076 21.764 ;
  LAYER M2 ;
        RECT 0.604 21.796 3.076 21.828 ;
  LAYER M2 ;
        RECT 0.604 21.86 3.076 21.892 ;
  LAYER M2 ;
        RECT 0.604 21.924 3.076 21.956 ;
  LAYER M2 ;
        RECT 0.604 21.988 3.076 22.02 ;
  LAYER M2 ;
        RECT 0.604 22.052 3.076 22.084 ;
  LAYER M2 ;
        RECT 0.604 22.116 3.076 22.148 ;
  LAYER M2 ;
        RECT 0.604 22.18 3.076 22.212 ;
  LAYER M2 ;
        RECT 0.604 22.244 3.076 22.276 ;
  LAYER M2 ;
        RECT 0.604 22.308 3.076 22.34 ;
  LAYER M2 ;
        RECT 0.604 22.372 3.076 22.404 ;
  LAYER M2 ;
        RECT 0.604 22.436 3.076 22.468 ;
  LAYER M2 ;
        RECT 0.604 22.5 3.076 22.532 ;
  LAYER M2 ;
        RECT 0.604 22.564 3.076 22.596 ;
  LAYER M2 ;
        RECT 0.604 22.628 3.076 22.66 ;
  LAYER M2 ;
        RECT 0.604 22.692 3.076 22.724 ;
  LAYER M2 ;
        RECT 0.604 22.756 3.076 22.788 ;
  LAYER M2 ;
        RECT 0.604 22.82 3.076 22.852 ;
  LAYER M2 ;
        RECT 0.604 22.884 3.076 22.916 ;
  LAYER M2 ;
        RECT 0.604 22.948 3.076 22.98 ;
  LAYER M2 ;
        RECT 0.604 23.012 3.076 23.044 ;
  LAYER M2 ;
        RECT 0.604 23.076 3.076 23.108 ;
  LAYER M2 ;
        RECT 0.604 23.14 3.076 23.172 ;
  LAYER M2 ;
        RECT 0.604 23.204 3.076 23.236 ;
  LAYER M3 ;
        RECT 0.624 20.88 0.656 23.388 ;
  LAYER M3 ;
        RECT 0.688 20.88 0.72 23.388 ;
  LAYER M3 ;
        RECT 0.752 20.88 0.784 23.388 ;
  LAYER M3 ;
        RECT 0.816 20.88 0.848 23.388 ;
  LAYER M3 ;
        RECT 0.88 20.88 0.912 23.388 ;
  LAYER M3 ;
        RECT 0.944 20.88 0.976 23.388 ;
  LAYER M3 ;
        RECT 1.008 20.88 1.04 23.388 ;
  LAYER M3 ;
        RECT 1.072 20.88 1.104 23.388 ;
  LAYER M3 ;
        RECT 1.136 20.88 1.168 23.388 ;
  LAYER M3 ;
        RECT 1.2 20.88 1.232 23.388 ;
  LAYER M3 ;
        RECT 1.264 20.88 1.296 23.388 ;
  LAYER M3 ;
        RECT 1.328 20.88 1.36 23.388 ;
  LAYER M3 ;
        RECT 1.392 20.88 1.424 23.388 ;
  LAYER M3 ;
        RECT 1.456 20.88 1.488 23.388 ;
  LAYER M3 ;
        RECT 1.52 20.88 1.552 23.388 ;
  LAYER M3 ;
        RECT 1.584 20.88 1.616 23.388 ;
  LAYER M3 ;
        RECT 1.648 20.88 1.68 23.388 ;
  LAYER M3 ;
        RECT 1.712 20.88 1.744 23.388 ;
  LAYER M3 ;
        RECT 1.776 20.88 1.808 23.388 ;
  LAYER M3 ;
        RECT 1.84 20.88 1.872 23.388 ;
  LAYER M3 ;
        RECT 1.904 20.88 1.936 23.388 ;
  LAYER M3 ;
        RECT 1.968 20.88 2 23.388 ;
  LAYER M3 ;
        RECT 2.032 20.88 2.064 23.388 ;
  LAYER M3 ;
        RECT 2.096 20.88 2.128 23.388 ;
  LAYER M3 ;
        RECT 2.16 20.88 2.192 23.388 ;
  LAYER M3 ;
        RECT 2.224 20.88 2.256 23.388 ;
  LAYER M3 ;
        RECT 2.288 20.88 2.32 23.388 ;
  LAYER M3 ;
        RECT 2.352 20.88 2.384 23.388 ;
  LAYER M3 ;
        RECT 2.416 20.88 2.448 23.388 ;
  LAYER M3 ;
        RECT 2.48 20.88 2.512 23.388 ;
  LAYER M3 ;
        RECT 2.544 20.88 2.576 23.388 ;
  LAYER M3 ;
        RECT 2.608 20.88 2.64 23.388 ;
  LAYER M3 ;
        RECT 2.672 20.88 2.704 23.388 ;
  LAYER M3 ;
        RECT 2.736 20.88 2.768 23.388 ;
  LAYER M3 ;
        RECT 2.8 20.88 2.832 23.388 ;
  LAYER M3 ;
        RECT 2.864 20.88 2.896 23.388 ;
  LAYER M3 ;
        RECT 2.928 20.88 2.96 23.388 ;
  LAYER M3 ;
        RECT 3.024 20.88 3.056 23.388 ;
  LAYER M1 ;
        RECT 0.639 20.916 0.641 23.352 ;
  LAYER M1 ;
        RECT 0.719 20.916 0.721 23.352 ;
  LAYER M1 ;
        RECT 0.799 20.916 0.801 23.352 ;
  LAYER M1 ;
        RECT 0.879 20.916 0.881 23.352 ;
  LAYER M1 ;
        RECT 0.959 20.916 0.961 23.352 ;
  LAYER M1 ;
        RECT 1.039 20.916 1.041 23.352 ;
  LAYER M1 ;
        RECT 1.119 20.916 1.121 23.352 ;
  LAYER M1 ;
        RECT 1.199 20.916 1.201 23.352 ;
  LAYER M1 ;
        RECT 1.279 20.916 1.281 23.352 ;
  LAYER M1 ;
        RECT 1.359 20.916 1.361 23.352 ;
  LAYER M1 ;
        RECT 1.439 20.916 1.441 23.352 ;
  LAYER M1 ;
        RECT 1.519 20.916 1.521 23.352 ;
  LAYER M1 ;
        RECT 1.599 20.916 1.601 23.352 ;
  LAYER M1 ;
        RECT 1.679 20.916 1.681 23.352 ;
  LAYER M1 ;
        RECT 1.759 20.916 1.761 23.352 ;
  LAYER M1 ;
        RECT 1.839 20.916 1.841 23.352 ;
  LAYER M1 ;
        RECT 1.919 20.916 1.921 23.352 ;
  LAYER M1 ;
        RECT 1.999 20.916 2.001 23.352 ;
  LAYER M1 ;
        RECT 2.079 20.916 2.081 23.352 ;
  LAYER M1 ;
        RECT 2.159 20.916 2.161 23.352 ;
  LAYER M1 ;
        RECT 2.239 20.916 2.241 23.352 ;
  LAYER M1 ;
        RECT 2.319 20.916 2.321 23.352 ;
  LAYER M1 ;
        RECT 2.399 20.916 2.401 23.352 ;
  LAYER M1 ;
        RECT 2.479 20.916 2.481 23.352 ;
  LAYER M1 ;
        RECT 2.559 20.916 2.561 23.352 ;
  LAYER M1 ;
        RECT 2.639 20.916 2.641 23.352 ;
  LAYER M1 ;
        RECT 2.719 20.916 2.721 23.352 ;
  LAYER M1 ;
        RECT 2.799 20.916 2.801 23.352 ;
  LAYER M1 ;
        RECT 2.879 20.916 2.881 23.352 ;
  LAYER M1 ;
        RECT 2.959 20.916 2.961 23.352 ;
  LAYER M2 ;
        RECT 0.64 20.915 3.04 20.917 ;
  LAYER M2 ;
        RECT 0.64 20.999 3.04 21.001 ;
  LAYER M2 ;
        RECT 0.64 21.083 3.04 21.085 ;
  LAYER M2 ;
        RECT 0.64 21.167 3.04 21.169 ;
  LAYER M2 ;
        RECT 0.64 21.251 3.04 21.253 ;
  LAYER M2 ;
        RECT 0.64 21.335 3.04 21.337 ;
  LAYER M2 ;
        RECT 0.64 21.419 3.04 21.421 ;
  LAYER M2 ;
        RECT 0.64 21.503 3.04 21.505 ;
  LAYER M2 ;
        RECT 0.64 21.587 3.04 21.589 ;
  LAYER M2 ;
        RECT 0.64 21.671 3.04 21.673 ;
  LAYER M2 ;
        RECT 0.64 21.755 3.04 21.757 ;
  LAYER M2 ;
        RECT 0.64 21.839 3.04 21.841 ;
  LAYER M2 ;
        RECT 0.64 21.9225 3.04 21.9245 ;
  LAYER M2 ;
        RECT 0.64 22.007 3.04 22.009 ;
  LAYER M2 ;
        RECT 0.64 22.091 3.04 22.093 ;
  LAYER M2 ;
        RECT 0.64 22.175 3.04 22.177 ;
  LAYER M2 ;
        RECT 0.64 22.259 3.04 22.261 ;
  LAYER M2 ;
        RECT 0.64 22.343 3.04 22.345 ;
  LAYER M2 ;
        RECT 0.64 22.427 3.04 22.429 ;
  LAYER M2 ;
        RECT 0.64 22.511 3.04 22.513 ;
  LAYER M2 ;
        RECT 0.64 22.595 3.04 22.597 ;
  LAYER M2 ;
        RECT 0.64 22.679 3.04 22.681 ;
  LAYER M2 ;
        RECT 0.64 22.763 3.04 22.765 ;
  LAYER M2 ;
        RECT 0.64 22.847 3.04 22.849 ;
  LAYER M2 ;
        RECT 0.64 22.931 3.04 22.933 ;
  LAYER M2 ;
        RECT 0.64 23.015 3.04 23.017 ;
  LAYER M2 ;
        RECT 0.64 23.099 3.04 23.101 ;
  LAYER M2 ;
        RECT 0.64 23.183 3.04 23.185 ;
  LAYER M2 ;
        RECT 0.64 23.267 3.04 23.269 ;
  LAYER M1 ;
        RECT 0.624 23.82 0.656 26.328 ;
  LAYER M1 ;
        RECT 0.688 23.82 0.72 26.328 ;
  LAYER M1 ;
        RECT 0.752 23.82 0.784 26.328 ;
  LAYER M1 ;
        RECT 0.816 23.82 0.848 26.328 ;
  LAYER M1 ;
        RECT 0.88 23.82 0.912 26.328 ;
  LAYER M1 ;
        RECT 0.944 23.82 0.976 26.328 ;
  LAYER M1 ;
        RECT 1.008 23.82 1.04 26.328 ;
  LAYER M1 ;
        RECT 1.072 23.82 1.104 26.328 ;
  LAYER M1 ;
        RECT 1.136 23.82 1.168 26.328 ;
  LAYER M1 ;
        RECT 1.2 23.82 1.232 26.328 ;
  LAYER M1 ;
        RECT 1.264 23.82 1.296 26.328 ;
  LAYER M1 ;
        RECT 1.328 23.82 1.36 26.328 ;
  LAYER M1 ;
        RECT 1.392 23.82 1.424 26.328 ;
  LAYER M1 ;
        RECT 1.456 23.82 1.488 26.328 ;
  LAYER M1 ;
        RECT 1.52 23.82 1.552 26.328 ;
  LAYER M1 ;
        RECT 1.584 23.82 1.616 26.328 ;
  LAYER M1 ;
        RECT 1.648 23.82 1.68 26.328 ;
  LAYER M1 ;
        RECT 1.712 23.82 1.744 26.328 ;
  LAYER M1 ;
        RECT 1.776 23.82 1.808 26.328 ;
  LAYER M1 ;
        RECT 1.84 23.82 1.872 26.328 ;
  LAYER M1 ;
        RECT 1.904 23.82 1.936 26.328 ;
  LAYER M1 ;
        RECT 1.968 23.82 2 26.328 ;
  LAYER M1 ;
        RECT 2.032 23.82 2.064 26.328 ;
  LAYER M1 ;
        RECT 2.096 23.82 2.128 26.328 ;
  LAYER M1 ;
        RECT 2.16 23.82 2.192 26.328 ;
  LAYER M1 ;
        RECT 2.224 23.82 2.256 26.328 ;
  LAYER M1 ;
        RECT 2.288 23.82 2.32 26.328 ;
  LAYER M1 ;
        RECT 2.352 23.82 2.384 26.328 ;
  LAYER M1 ;
        RECT 2.416 23.82 2.448 26.328 ;
  LAYER M1 ;
        RECT 2.48 23.82 2.512 26.328 ;
  LAYER M1 ;
        RECT 2.544 23.82 2.576 26.328 ;
  LAYER M1 ;
        RECT 2.608 23.82 2.64 26.328 ;
  LAYER M1 ;
        RECT 2.672 23.82 2.704 26.328 ;
  LAYER M1 ;
        RECT 2.736 23.82 2.768 26.328 ;
  LAYER M1 ;
        RECT 2.8 23.82 2.832 26.328 ;
  LAYER M1 ;
        RECT 2.864 23.82 2.896 26.328 ;
  LAYER M1 ;
        RECT 2.928 23.82 2.96 26.328 ;
  LAYER M2 ;
        RECT 0.604 23.904 3.076 23.936 ;
  LAYER M2 ;
        RECT 0.604 23.968 3.076 24 ;
  LAYER M2 ;
        RECT 0.604 24.032 3.076 24.064 ;
  LAYER M2 ;
        RECT 0.604 24.096 3.076 24.128 ;
  LAYER M2 ;
        RECT 0.604 24.16 3.076 24.192 ;
  LAYER M2 ;
        RECT 0.604 24.224 3.076 24.256 ;
  LAYER M2 ;
        RECT 0.604 24.288 3.076 24.32 ;
  LAYER M2 ;
        RECT 0.604 24.352 3.076 24.384 ;
  LAYER M2 ;
        RECT 0.604 24.416 3.076 24.448 ;
  LAYER M2 ;
        RECT 0.604 24.48 3.076 24.512 ;
  LAYER M2 ;
        RECT 0.604 24.544 3.076 24.576 ;
  LAYER M2 ;
        RECT 0.604 24.608 3.076 24.64 ;
  LAYER M2 ;
        RECT 0.604 24.672 3.076 24.704 ;
  LAYER M2 ;
        RECT 0.604 24.736 3.076 24.768 ;
  LAYER M2 ;
        RECT 0.604 24.8 3.076 24.832 ;
  LAYER M2 ;
        RECT 0.604 24.864 3.076 24.896 ;
  LAYER M2 ;
        RECT 0.604 24.928 3.076 24.96 ;
  LAYER M2 ;
        RECT 0.604 24.992 3.076 25.024 ;
  LAYER M2 ;
        RECT 0.604 25.056 3.076 25.088 ;
  LAYER M2 ;
        RECT 0.604 25.12 3.076 25.152 ;
  LAYER M2 ;
        RECT 0.604 25.184 3.076 25.216 ;
  LAYER M2 ;
        RECT 0.604 25.248 3.076 25.28 ;
  LAYER M2 ;
        RECT 0.604 25.312 3.076 25.344 ;
  LAYER M2 ;
        RECT 0.604 25.376 3.076 25.408 ;
  LAYER M2 ;
        RECT 0.604 25.44 3.076 25.472 ;
  LAYER M2 ;
        RECT 0.604 25.504 3.076 25.536 ;
  LAYER M2 ;
        RECT 0.604 25.568 3.076 25.6 ;
  LAYER M2 ;
        RECT 0.604 25.632 3.076 25.664 ;
  LAYER M2 ;
        RECT 0.604 25.696 3.076 25.728 ;
  LAYER M2 ;
        RECT 0.604 25.76 3.076 25.792 ;
  LAYER M2 ;
        RECT 0.604 25.824 3.076 25.856 ;
  LAYER M2 ;
        RECT 0.604 25.888 3.076 25.92 ;
  LAYER M2 ;
        RECT 0.604 25.952 3.076 25.984 ;
  LAYER M2 ;
        RECT 0.604 26.016 3.076 26.048 ;
  LAYER M2 ;
        RECT 0.604 26.08 3.076 26.112 ;
  LAYER M2 ;
        RECT 0.604 26.144 3.076 26.176 ;
  LAYER M3 ;
        RECT 0.624 23.82 0.656 26.328 ;
  LAYER M3 ;
        RECT 0.688 23.82 0.72 26.328 ;
  LAYER M3 ;
        RECT 0.752 23.82 0.784 26.328 ;
  LAYER M3 ;
        RECT 0.816 23.82 0.848 26.328 ;
  LAYER M3 ;
        RECT 0.88 23.82 0.912 26.328 ;
  LAYER M3 ;
        RECT 0.944 23.82 0.976 26.328 ;
  LAYER M3 ;
        RECT 1.008 23.82 1.04 26.328 ;
  LAYER M3 ;
        RECT 1.072 23.82 1.104 26.328 ;
  LAYER M3 ;
        RECT 1.136 23.82 1.168 26.328 ;
  LAYER M3 ;
        RECT 1.2 23.82 1.232 26.328 ;
  LAYER M3 ;
        RECT 1.264 23.82 1.296 26.328 ;
  LAYER M3 ;
        RECT 1.328 23.82 1.36 26.328 ;
  LAYER M3 ;
        RECT 1.392 23.82 1.424 26.328 ;
  LAYER M3 ;
        RECT 1.456 23.82 1.488 26.328 ;
  LAYER M3 ;
        RECT 1.52 23.82 1.552 26.328 ;
  LAYER M3 ;
        RECT 1.584 23.82 1.616 26.328 ;
  LAYER M3 ;
        RECT 1.648 23.82 1.68 26.328 ;
  LAYER M3 ;
        RECT 1.712 23.82 1.744 26.328 ;
  LAYER M3 ;
        RECT 1.776 23.82 1.808 26.328 ;
  LAYER M3 ;
        RECT 1.84 23.82 1.872 26.328 ;
  LAYER M3 ;
        RECT 1.904 23.82 1.936 26.328 ;
  LAYER M3 ;
        RECT 1.968 23.82 2 26.328 ;
  LAYER M3 ;
        RECT 2.032 23.82 2.064 26.328 ;
  LAYER M3 ;
        RECT 2.096 23.82 2.128 26.328 ;
  LAYER M3 ;
        RECT 2.16 23.82 2.192 26.328 ;
  LAYER M3 ;
        RECT 2.224 23.82 2.256 26.328 ;
  LAYER M3 ;
        RECT 2.288 23.82 2.32 26.328 ;
  LAYER M3 ;
        RECT 2.352 23.82 2.384 26.328 ;
  LAYER M3 ;
        RECT 2.416 23.82 2.448 26.328 ;
  LAYER M3 ;
        RECT 2.48 23.82 2.512 26.328 ;
  LAYER M3 ;
        RECT 2.544 23.82 2.576 26.328 ;
  LAYER M3 ;
        RECT 2.608 23.82 2.64 26.328 ;
  LAYER M3 ;
        RECT 2.672 23.82 2.704 26.328 ;
  LAYER M3 ;
        RECT 2.736 23.82 2.768 26.328 ;
  LAYER M3 ;
        RECT 2.8 23.82 2.832 26.328 ;
  LAYER M3 ;
        RECT 2.864 23.82 2.896 26.328 ;
  LAYER M3 ;
        RECT 2.928 23.82 2.96 26.328 ;
  LAYER M3 ;
        RECT 3.024 23.82 3.056 26.328 ;
  LAYER M1 ;
        RECT 0.639 23.856 0.641 26.292 ;
  LAYER M1 ;
        RECT 0.719 23.856 0.721 26.292 ;
  LAYER M1 ;
        RECT 0.799 23.856 0.801 26.292 ;
  LAYER M1 ;
        RECT 0.879 23.856 0.881 26.292 ;
  LAYER M1 ;
        RECT 0.959 23.856 0.961 26.292 ;
  LAYER M1 ;
        RECT 1.039 23.856 1.041 26.292 ;
  LAYER M1 ;
        RECT 1.119 23.856 1.121 26.292 ;
  LAYER M1 ;
        RECT 1.199 23.856 1.201 26.292 ;
  LAYER M1 ;
        RECT 1.279 23.856 1.281 26.292 ;
  LAYER M1 ;
        RECT 1.359 23.856 1.361 26.292 ;
  LAYER M1 ;
        RECT 1.439 23.856 1.441 26.292 ;
  LAYER M1 ;
        RECT 1.519 23.856 1.521 26.292 ;
  LAYER M1 ;
        RECT 1.599 23.856 1.601 26.292 ;
  LAYER M1 ;
        RECT 1.679 23.856 1.681 26.292 ;
  LAYER M1 ;
        RECT 1.759 23.856 1.761 26.292 ;
  LAYER M1 ;
        RECT 1.839 23.856 1.841 26.292 ;
  LAYER M1 ;
        RECT 1.919 23.856 1.921 26.292 ;
  LAYER M1 ;
        RECT 1.999 23.856 2.001 26.292 ;
  LAYER M1 ;
        RECT 2.079 23.856 2.081 26.292 ;
  LAYER M1 ;
        RECT 2.159 23.856 2.161 26.292 ;
  LAYER M1 ;
        RECT 2.239 23.856 2.241 26.292 ;
  LAYER M1 ;
        RECT 2.319 23.856 2.321 26.292 ;
  LAYER M1 ;
        RECT 2.399 23.856 2.401 26.292 ;
  LAYER M1 ;
        RECT 2.479 23.856 2.481 26.292 ;
  LAYER M1 ;
        RECT 2.559 23.856 2.561 26.292 ;
  LAYER M1 ;
        RECT 2.639 23.856 2.641 26.292 ;
  LAYER M1 ;
        RECT 2.719 23.856 2.721 26.292 ;
  LAYER M1 ;
        RECT 2.799 23.856 2.801 26.292 ;
  LAYER M1 ;
        RECT 2.879 23.856 2.881 26.292 ;
  LAYER M1 ;
        RECT 2.959 23.856 2.961 26.292 ;
  LAYER M2 ;
        RECT 0.64 23.855 3.04 23.857 ;
  LAYER M2 ;
        RECT 0.64 23.939 3.04 23.941 ;
  LAYER M2 ;
        RECT 0.64 24.023 3.04 24.025 ;
  LAYER M2 ;
        RECT 0.64 24.107 3.04 24.109 ;
  LAYER M2 ;
        RECT 0.64 24.191 3.04 24.193 ;
  LAYER M2 ;
        RECT 0.64 24.275 3.04 24.277 ;
  LAYER M2 ;
        RECT 0.64 24.359 3.04 24.361 ;
  LAYER M2 ;
        RECT 0.64 24.443 3.04 24.445 ;
  LAYER M2 ;
        RECT 0.64 24.527 3.04 24.529 ;
  LAYER M2 ;
        RECT 0.64 24.611 3.04 24.613 ;
  LAYER M2 ;
        RECT 0.64 24.695 3.04 24.697 ;
  LAYER M2 ;
        RECT 0.64 24.779 3.04 24.781 ;
  LAYER M2 ;
        RECT 0.64 24.8625 3.04 24.8645 ;
  LAYER M2 ;
        RECT 0.64 24.947 3.04 24.949 ;
  LAYER M2 ;
        RECT 0.64 25.031 3.04 25.033 ;
  LAYER M2 ;
        RECT 0.64 25.115 3.04 25.117 ;
  LAYER M2 ;
        RECT 0.64 25.199 3.04 25.201 ;
  LAYER M2 ;
        RECT 0.64 25.283 3.04 25.285 ;
  LAYER M2 ;
        RECT 0.64 25.367 3.04 25.369 ;
  LAYER M2 ;
        RECT 0.64 25.451 3.04 25.453 ;
  LAYER M2 ;
        RECT 0.64 25.535 3.04 25.537 ;
  LAYER M2 ;
        RECT 0.64 25.619 3.04 25.621 ;
  LAYER M2 ;
        RECT 0.64 25.703 3.04 25.705 ;
  LAYER M2 ;
        RECT 0.64 25.787 3.04 25.789 ;
  LAYER M2 ;
        RECT 0.64 25.871 3.04 25.873 ;
  LAYER M2 ;
        RECT 0.64 25.955 3.04 25.957 ;
  LAYER M2 ;
        RECT 0.64 26.039 3.04 26.041 ;
  LAYER M2 ;
        RECT 0.64 26.123 3.04 26.125 ;
  LAYER M2 ;
        RECT 0.64 26.207 3.04 26.209 ;
  LAYER M1 ;
        RECT 0.624 26.76 0.656 29.268 ;
  LAYER M1 ;
        RECT 0.688 26.76 0.72 29.268 ;
  LAYER M1 ;
        RECT 0.752 26.76 0.784 29.268 ;
  LAYER M1 ;
        RECT 0.816 26.76 0.848 29.268 ;
  LAYER M1 ;
        RECT 0.88 26.76 0.912 29.268 ;
  LAYER M1 ;
        RECT 0.944 26.76 0.976 29.268 ;
  LAYER M1 ;
        RECT 1.008 26.76 1.04 29.268 ;
  LAYER M1 ;
        RECT 1.072 26.76 1.104 29.268 ;
  LAYER M1 ;
        RECT 1.136 26.76 1.168 29.268 ;
  LAYER M1 ;
        RECT 1.2 26.76 1.232 29.268 ;
  LAYER M1 ;
        RECT 1.264 26.76 1.296 29.268 ;
  LAYER M1 ;
        RECT 1.328 26.76 1.36 29.268 ;
  LAYER M1 ;
        RECT 1.392 26.76 1.424 29.268 ;
  LAYER M1 ;
        RECT 1.456 26.76 1.488 29.268 ;
  LAYER M1 ;
        RECT 1.52 26.76 1.552 29.268 ;
  LAYER M1 ;
        RECT 1.584 26.76 1.616 29.268 ;
  LAYER M1 ;
        RECT 1.648 26.76 1.68 29.268 ;
  LAYER M1 ;
        RECT 1.712 26.76 1.744 29.268 ;
  LAYER M1 ;
        RECT 1.776 26.76 1.808 29.268 ;
  LAYER M1 ;
        RECT 1.84 26.76 1.872 29.268 ;
  LAYER M1 ;
        RECT 1.904 26.76 1.936 29.268 ;
  LAYER M1 ;
        RECT 1.968 26.76 2 29.268 ;
  LAYER M1 ;
        RECT 2.032 26.76 2.064 29.268 ;
  LAYER M1 ;
        RECT 2.096 26.76 2.128 29.268 ;
  LAYER M1 ;
        RECT 2.16 26.76 2.192 29.268 ;
  LAYER M1 ;
        RECT 2.224 26.76 2.256 29.268 ;
  LAYER M1 ;
        RECT 2.288 26.76 2.32 29.268 ;
  LAYER M1 ;
        RECT 2.352 26.76 2.384 29.268 ;
  LAYER M1 ;
        RECT 2.416 26.76 2.448 29.268 ;
  LAYER M1 ;
        RECT 2.48 26.76 2.512 29.268 ;
  LAYER M1 ;
        RECT 2.544 26.76 2.576 29.268 ;
  LAYER M1 ;
        RECT 2.608 26.76 2.64 29.268 ;
  LAYER M1 ;
        RECT 2.672 26.76 2.704 29.268 ;
  LAYER M1 ;
        RECT 2.736 26.76 2.768 29.268 ;
  LAYER M1 ;
        RECT 2.8 26.76 2.832 29.268 ;
  LAYER M1 ;
        RECT 2.864 26.76 2.896 29.268 ;
  LAYER M1 ;
        RECT 2.928 26.76 2.96 29.268 ;
  LAYER M2 ;
        RECT 0.604 26.844 3.076 26.876 ;
  LAYER M2 ;
        RECT 0.604 26.908 3.076 26.94 ;
  LAYER M2 ;
        RECT 0.604 26.972 3.076 27.004 ;
  LAYER M2 ;
        RECT 0.604 27.036 3.076 27.068 ;
  LAYER M2 ;
        RECT 0.604 27.1 3.076 27.132 ;
  LAYER M2 ;
        RECT 0.604 27.164 3.076 27.196 ;
  LAYER M2 ;
        RECT 0.604 27.228 3.076 27.26 ;
  LAYER M2 ;
        RECT 0.604 27.292 3.076 27.324 ;
  LAYER M2 ;
        RECT 0.604 27.356 3.076 27.388 ;
  LAYER M2 ;
        RECT 0.604 27.42 3.076 27.452 ;
  LAYER M2 ;
        RECT 0.604 27.484 3.076 27.516 ;
  LAYER M2 ;
        RECT 0.604 27.548 3.076 27.58 ;
  LAYER M2 ;
        RECT 0.604 27.612 3.076 27.644 ;
  LAYER M2 ;
        RECT 0.604 27.676 3.076 27.708 ;
  LAYER M2 ;
        RECT 0.604 27.74 3.076 27.772 ;
  LAYER M2 ;
        RECT 0.604 27.804 3.076 27.836 ;
  LAYER M2 ;
        RECT 0.604 27.868 3.076 27.9 ;
  LAYER M2 ;
        RECT 0.604 27.932 3.076 27.964 ;
  LAYER M2 ;
        RECT 0.604 27.996 3.076 28.028 ;
  LAYER M2 ;
        RECT 0.604 28.06 3.076 28.092 ;
  LAYER M2 ;
        RECT 0.604 28.124 3.076 28.156 ;
  LAYER M2 ;
        RECT 0.604 28.188 3.076 28.22 ;
  LAYER M2 ;
        RECT 0.604 28.252 3.076 28.284 ;
  LAYER M2 ;
        RECT 0.604 28.316 3.076 28.348 ;
  LAYER M2 ;
        RECT 0.604 28.38 3.076 28.412 ;
  LAYER M2 ;
        RECT 0.604 28.444 3.076 28.476 ;
  LAYER M2 ;
        RECT 0.604 28.508 3.076 28.54 ;
  LAYER M2 ;
        RECT 0.604 28.572 3.076 28.604 ;
  LAYER M2 ;
        RECT 0.604 28.636 3.076 28.668 ;
  LAYER M2 ;
        RECT 0.604 28.7 3.076 28.732 ;
  LAYER M2 ;
        RECT 0.604 28.764 3.076 28.796 ;
  LAYER M2 ;
        RECT 0.604 28.828 3.076 28.86 ;
  LAYER M2 ;
        RECT 0.604 28.892 3.076 28.924 ;
  LAYER M2 ;
        RECT 0.604 28.956 3.076 28.988 ;
  LAYER M2 ;
        RECT 0.604 29.02 3.076 29.052 ;
  LAYER M2 ;
        RECT 0.604 29.084 3.076 29.116 ;
  LAYER M3 ;
        RECT 0.624 26.76 0.656 29.268 ;
  LAYER M3 ;
        RECT 0.688 26.76 0.72 29.268 ;
  LAYER M3 ;
        RECT 0.752 26.76 0.784 29.268 ;
  LAYER M3 ;
        RECT 0.816 26.76 0.848 29.268 ;
  LAYER M3 ;
        RECT 0.88 26.76 0.912 29.268 ;
  LAYER M3 ;
        RECT 0.944 26.76 0.976 29.268 ;
  LAYER M3 ;
        RECT 1.008 26.76 1.04 29.268 ;
  LAYER M3 ;
        RECT 1.072 26.76 1.104 29.268 ;
  LAYER M3 ;
        RECT 1.136 26.76 1.168 29.268 ;
  LAYER M3 ;
        RECT 1.2 26.76 1.232 29.268 ;
  LAYER M3 ;
        RECT 1.264 26.76 1.296 29.268 ;
  LAYER M3 ;
        RECT 1.328 26.76 1.36 29.268 ;
  LAYER M3 ;
        RECT 1.392 26.76 1.424 29.268 ;
  LAYER M3 ;
        RECT 1.456 26.76 1.488 29.268 ;
  LAYER M3 ;
        RECT 1.52 26.76 1.552 29.268 ;
  LAYER M3 ;
        RECT 1.584 26.76 1.616 29.268 ;
  LAYER M3 ;
        RECT 1.648 26.76 1.68 29.268 ;
  LAYER M3 ;
        RECT 1.712 26.76 1.744 29.268 ;
  LAYER M3 ;
        RECT 1.776 26.76 1.808 29.268 ;
  LAYER M3 ;
        RECT 1.84 26.76 1.872 29.268 ;
  LAYER M3 ;
        RECT 1.904 26.76 1.936 29.268 ;
  LAYER M3 ;
        RECT 1.968 26.76 2 29.268 ;
  LAYER M3 ;
        RECT 2.032 26.76 2.064 29.268 ;
  LAYER M3 ;
        RECT 2.096 26.76 2.128 29.268 ;
  LAYER M3 ;
        RECT 2.16 26.76 2.192 29.268 ;
  LAYER M3 ;
        RECT 2.224 26.76 2.256 29.268 ;
  LAYER M3 ;
        RECT 2.288 26.76 2.32 29.268 ;
  LAYER M3 ;
        RECT 2.352 26.76 2.384 29.268 ;
  LAYER M3 ;
        RECT 2.416 26.76 2.448 29.268 ;
  LAYER M3 ;
        RECT 2.48 26.76 2.512 29.268 ;
  LAYER M3 ;
        RECT 2.544 26.76 2.576 29.268 ;
  LAYER M3 ;
        RECT 2.608 26.76 2.64 29.268 ;
  LAYER M3 ;
        RECT 2.672 26.76 2.704 29.268 ;
  LAYER M3 ;
        RECT 2.736 26.76 2.768 29.268 ;
  LAYER M3 ;
        RECT 2.8 26.76 2.832 29.268 ;
  LAYER M3 ;
        RECT 2.864 26.76 2.896 29.268 ;
  LAYER M3 ;
        RECT 2.928 26.76 2.96 29.268 ;
  LAYER M3 ;
        RECT 3.024 26.76 3.056 29.268 ;
  LAYER M1 ;
        RECT 0.639 26.796 0.641 29.232 ;
  LAYER M1 ;
        RECT 0.719 26.796 0.721 29.232 ;
  LAYER M1 ;
        RECT 0.799 26.796 0.801 29.232 ;
  LAYER M1 ;
        RECT 0.879 26.796 0.881 29.232 ;
  LAYER M1 ;
        RECT 0.959 26.796 0.961 29.232 ;
  LAYER M1 ;
        RECT 1.039 26.796 1.041 29.232 ;
  LAYER M1 ;
        RECT 1.119 26.796 1.121 29.232 ;
  LAYER M1 ;
        RECT 1.199 26.796 1.201 29.232 ;
  LAYER M1 ;
        RECT 1.279 26.796 1.281 29.232 ;
  LAYER M1 ;
        RECT 1.359 26.796 1.361 29.232 ;
  LAYER M1 ;
        RECT 1.439 26.796 1.441 29.232 ;
  LAYER M1 ;
        RECT 1.519 26.796 1.521 29.232 ;
  LAYER M1 ;
        RECT 1.599 26.796 1.601 29.232 ;
  LAYER M1 ;
        RECT 1.679 26.796 1.681 29.232 ;
  LAYER M1 ;
        RECT 1.759 26.796 1.761 29.232 ;
  LAYER M1 ;
        RECT 1.839 26.796 1.841 29.232 ;
  LAYER M1 ;
        RECT 1.919 26.796 1.921 29.232 ;
  LAYER M1 ;
        RECT 1.999 26.796 2.001 29.232 ;
  LAYER M1 ;
        RECT 2.079 26.796 2.081 29.232 ;
  LAYER M1 ;
        RECT 2.159 26.796 2.161 29.232 ;
  LAYER M1 ;
        RECT 2.239 26.796 2.241 29.232 ;
  LAYER M1 ;
        RECT 2.319 26.796 2.321 29.232 ;
  LAYER M1 ;
        RECT 2.399 26.796 2.401 29.232 ;
  LAYER M1 ;
        RECT 2.479 26.796 2.481 29.232 ;
  LAYER M1 ;
        RECT 2.559 26.796 2.561 29.232 ;
  LAYER M1 ;
        RECT 2.639 26.796 2.641 29.232 ;
  LAYER M1 ;
        RECT 2.719 26.796 2.721 29.232 ;
  LAYER M1 ;
        RECT 2.799 26.796 2.801 29.232 ;
  LAYER M1 ;
        RECT 2.879 26.796 2.881 29.232 ;
  LAYER M1 ;
        RECT 2.959 26.796 2.961 29.232 ;
  LAYER M2 ;
        RECT 0.64 26.795 3.04 26.797 ;
  LAYER M2 ;
        RECT 0.64 26.879 3.04 26.881 ;
  LAYER M2 ;
        RECT 0.64 26.963 3.04 26.965 ;
  LAYER M2 ;
        RECT 0.64 27.047 3.04 27.049 ;
  LAYER M2 ;
        RECT 0.64 27.131 3.04 27.133 ;
  LAYER M2 ;
        RECT 0.64 27.215 3.04 27.217 ;
  LAYER M2 ;
        RECT 0.64 27.299 3.04 27.301 ;
  LAYER M2 ;
        RECT 0.64 27.383 3.04 27.385 ;
  LAYER M2 ;
        RECT 0.64 27.467 3.04 27.469 ;
  LAYER M2 ;
        RECT 0.64 27.551 3.04 27.553 ;
  LAYER M2 ;
        RECT 0.64 27.635 3.04 27.637 ;
  LAYER M2 ;
        RECT 0.64 27.719 3.04 27.721 ;
  LAYER M2 ;
        RECT 0.64 27.8025 3.04 27.8045 ;
  LAYER M2 ;
        RECT 0.64 27.887 3.04 27.889 ;
  LAYER M2 ;
        RECT 0.64 27.971 3.04 27.973 ;
  LAYER M2 ;
        RECT 0.64 28.055 3.04 28.057 ;
  LAYER M2 ;
        RECT 0.64 28.139 3.04 28.141 ;
  LAYER M2 ;
        RECT 0.64 28.223 3.04 28.225 ;
  LAYER M2 ;
        RECT 0.64 28.307 3.04 28.309 ;
  LAYER M2 ;
        RECT 0.64 28.391 3.04 28.393 ;
  LAYER M2 ;
        RECT 0.64 28.475 3.04 28.477 ;
  LAYER M2 ;
        RECT 0.64 28.559 3.04 28.561 ;
  LAYER M2 ;
        RECT 0.64 28.643 3.04 28.645 ;
  LAYER M2 ;
        RECT 0.64 28.727 3.04 28.729 ;
  LAYER M2 ;
        RECT 0.64 28.811 3.04 28.813 ;
  LAYER M2 ;
        RECT 0.64 28.895 3.04 28.897 ;
  LAYER M2 ;
        RECT 0.64 28.979 3.04 28.981 ;
  LAYER M2 ;
        RECT 0.64 29.063 3.04 29.065 ;
  LAYER M2 ;
        RECT 0.64 29.147 3.04 29.149 ;
  LAYER M1 ;
        RECT 3.504 17.94 3.536 20.448 ;
  LAYER M1 ;
        RECT 3.568 17.94 3.6 20.448 ;
  LAYER M1 ;
        RECT 3.632 17.94 3.664 20.448 ;
  LAYER M1 ;
        RECT 3.696 17.94 3.728 20.448 ;
  LAYER M1 ;
        RECT 3.76 17.94 3.792 20.448 ;
  LAYER M1 ;
        RECT 3.824 17.94 3.856 20.448 ;
  LAYER M1 ;
        RECT 3.888 17.94 3.92 20.448 ;
  LAYER M1 ;
        RECT 3.952 17.94 3.984 20.448 ;
  LAYER M1 ;
        RECT 4.016 17.94 4.048 20.448 ;
  LAYER M1 ;
        RECT 4.08 17.94 4.112 20.448 ;
  LAYER M1 ;
        RECT 4.144 17.94 4.176 20.448 ;
  LAYER M1 ;
        RECT 4.208 17.94 4.24 20.448 ;
  LAYER M1 ;
        RECT 4.272 17.94 4.304 20.448 ;
  LAYER M1 ;
        RECT 4.336 17.94 4.368 20.448 ;
  LAYER M1 ;
        RECT 4.4 17.94 4.432 20.448 ;
  LAYER M1 ;
        RECT 4.464 17.94 4.496 20.448 ;
  LAYER M1 ;
        RECT 4.528 17.94 4.56 20.448 ;
  LAYER M1 ;
        RECT 4.592 17.94 4.624 20.448 ;
  LAYER M1 ;
        RECT 4.656 17.94 4.688 20.448 ;
  LAYER M1 ;
        RECT 4.72 17.94 4.752 20.448 ;
  LAYER M1 ;
        RECT 4.784 17.94 4.816 20.448 ;
  LAYER M1 ;
        RECT 4.848 17.94 4.88 20.448 ;
  LAYER M1 ;
        RECT 4.912 17.94 4.944 20.448 ;
  LAYER M1 ;
        RECT 4.976 17.94 5.008 20.448 ;
  LAYER M1 ;
        RECT 5.04 17.94 5.072 20.448 ;
  LAYER M1 ;
        RECT 5.104 17.94 5.136 20.448 ;
  LAYER M1 ;
        RECT 5.168 17.94 5.2 20.448 ;
  LAYER M1 ;
        RECT 5.232 17.94 5.264 20.448 ;
  LAYER M1 ;
        RECT 5.296 17.94 5.328 20.448 ;
  LAYER M1 ;
        RECT 5.36 17.94 5.392 20.448 ;
  LAYER M1 ;
        RECT 5.424 17.94 5.456 20.448 ;
  LAYER M1 ;
        RECT 5.488 17.94 5.52 20.448 ;
  LAYER M1 ;
        RECT 5.552 17.94 5.584 20.448 ;
  LAYER M1 ;
        RECT 5.616 17.94 5.648 20.448 ;
  LAYER M1 ;
        RECT 5.68 17.94 5.712 20.448 ;
  LAYER M1 ;
        RECT 5.744 17.94 5.776 20.448 ;
  LAYER M1 ;
        RECT 5.808 17.94 5.84 20.448 ;
  LAYER M2 ;
        RECT 3.484 18.024 5.956 18.056 ;
  LAYER M2 ;
        RECT 3.484 18.088 5.956 18.12 ;
  LAYER M2 ;
        RECT 3.484 18.152 5.956 18.184 ;
  LAYER M2 ;
        RECT 3.484 18.216 5.956 18.248 ;
  LAYER M2 ;
        RECT 3.484 18.28 5.956 18.312 ;
  LAYER M2 ;
        RECT 3.484 18.344 5.956 18.376 ;
  LAYER M2 ;
        RECT 3.484 18.408 5.956 18.44 ;
  LAYER M2 ;
        RECT 3.484 18.472 5.956 18.504 ;
  LAYER M2 ;
        RECT 3.484 18.536 5.956 18.568 ;
  LAYER M2 ;
        RECT 3.484 18.6 5.956 18.632 ;
  LAYER M2 ;
        RECT 3.484 18.664 5.956 18.696 ;
  LAYER M2 ;
        RECT 3.484 18.728 5.956 18.76 ;
  LAYER M2 ;
        RECT 3.484 18.792 5.956 18.824 ;
  LAYER M2 ;
        RECT 3.484 18.856 5.956 18.888 ;
  LAYER M2 ;
        RECT 3.484 18.92 5.956 18.952 ;
  LAYER M2 ;
        RECT 3.484 18.984 5.956 19.016 ;
  LAYER M2 ;
        RECT 3.484 19.048 5.956 19.08 ;
  LAYER M2 ;
        RECT 3.484 19.112 5.956 19.144 ;
  LAYER M2 ;
        RECT 3.484 19.176 5.956 19.208 ;
  LAYER M2 ;
        RECT 3.484 19.24 5.956 19.272 ;
  LAYER M2 ;
        RECT 3.484 19.304 5.956 19.336 ;
  LAYER M2 ;
        RECT 3.484 19.368 5.956 19.4 ;
  LAYER M2 ;
        RECT 3.484 19.432 5.956 19.464 ;
  LAYER M2 ;
        RECT 3.484 19.496 5.956 19.528 ;
  LAYER M2 ;
        RECT 3.484 19.56 5.956 19.592 ;
  LAYER M2 ;
        RECT 3.484 19.624 5.956 19.656 ;
  LAYER M2 ;
        RECT 3.484 19.688 5.956 19.72 ;
  LAYER M2 ;
        RECT 3.484 19.752 5.956 19.784 ;
  LAYER M2 ;
        RECT 3.484 19.816 5.956 19.848 ;
  LAYER M2 ;
        RECT 3.484 19.88 5.956 19.912 ;
  LAYER M2 ;
        RECT 3.484 19.944 5.956 19.976 ;
  LAYER M2 ;
        RECT 3.484 20.008 5.956 20.04 ;
  LAYER M2 ;
        RECT 3.484 20.072 5.956 20.104 ;
  LAYER M2 ;
        RECT 3.484 20.136 5.956 20.168 ;
  LAYER M2 ;
        RECT 3.484 20.2 5.956 20.232 ;
  LAYER M2 ;
        RECT 3.484 20.264 5.956 20.296 ;
  LAYER M3 ;
        RECT 3.504 17.94 3.536 20.448 ;
  LAYER M3 ;
        RECT 3.568 17.94 3.6 20.448 ;
  LAYER M3 ;
        RECT 3.632 17.94 3.664 20.448 ;
  LAYER M3 ;
        RECT 3.696 17.94 3.728 20.448 ;
  LAYER M3 ;
        RECT 3.76 17.94 3.792 20.448 ;
  LAYER M3 ;
        RECT 3.824 17.94 3.856 20.448 ;
  LAYER M3 ;
        RECT 3.888 17.94 3.92 20.448 ;
  LAYER M3 ;
        RECT 3.952 17.94 3.984 20.448 ;
  LAYER M3 ;
        RECT 4.016 17.94 4.048 20.448 ;
  LAYER M3 ;
        RECT 4.08 17.94 4.112 20.448 ;
  LAYER M3 ;
        RECT 4.144 17.94 4.176 20.448 ;
  LAYER M3 ;
        RECT 4.208 17.94 4.24 20.448 ;
  LAYER M3 ;
        RECT 4.272 17.94 4.304 20.448 ;
  LAYER M3 ;
        RECT 4.336 17.94 4.368 20.448 ;
  LAYER M3 ;
        RECT 4.4 17.94 4.432 20.448 ;
  LAYER M3 ;
        RECT 4.464 17.94 4.496 20.448 ;
  LAYER M3 ;
        RECT 4.528 17.94 4.56 20.448 ;
  LAYER M3 ;
        RECT 4.592 17.94 4.624 20.448 ;
  LAYER M3 ;
        RECT 4.656 17.94 4.688 20.448 ;
  LAYER M3 ;
        RECT 4.72 17.94 4.752 20.448 ;
  LAYER M3 ;
        RECT 4.784 17.94 4.816 20.448 ;
  LAYER M3 ;
        RECT 4.848 17.94 4.88 20.448 ;
  LAYER M3 ;
        RECT 4.912 17.94 4.944 20.448 ;
  LAYER M3 ;
        RECT 4.976 17.94 5.008 20.448 ;
  LAYER M3 ;
        RECT 5.04 17.94 5.072 20.448 ;
  LAYER M3 ;
        RECT 5.104 17.94 5.136 20.448 ;
  LAYER M3 ;
        RECT 5.168 17.94 5.2 20.448 ;
  LAYER M3 ;
        RECT 5.232 17.94 5.264 20.448 ;
  LAYER M3 ;
        RECT 5.296 17.94 5.328 20.448 ;
  LAYER M3 ;
        RECT 5.36 17.94 5.392 20.448 ;
  LAYER M3 ;
        RECT 5.424 17.94 5.456 20.448 ;
  LAYER M3 ;
        RECT 5.488 17.94 5.52 20.448 ;
  LAYER M3 ;
        RECT 5.552 17.94 5.584 20.448 ;
  LAYER M3 ;
        RECT 5.616 17.94 5.648 20.448 ;
  LAYER M3 ;
        RECT 5.68 17.94 5.712 20.448 ;
  LAYER M3 ;
        RECT 5.744 17.94 5.776 20.448 ;
  LAYER M3 ;
        RECT 5.808 17.94 5.84 20.448 ;
  LAYER M3 ;
        RECT 5.904 17.94 5.936 20.448 ;
  LAYER M1 ;
        RECT 3.519 17.976 3.521 20.412 ;
  LAYER M1 ;
        RECT 3.599 17.976 3.601 20.412 ;
  LAYER M1 ;
        RECT 3.679 17.976 3.681 20.412 ;
  LAYER M1 ;
        RECT 3.759 17.976 3.761 20.412 ;
  LAYER M1 ;
        RECT 3.839 17.976 3.841 20.412 ;
  LAYER M1 ;
        RECT 3.919 17.976 3.921 20.412 ;
  LAYER M1 ;
        RECT 3.999 17.976 4.001 20.412 ;
  LAYER M1 ;
        RECT 4.079 17.976 4.081 20.412 ;
  LAYER M1 ;
        RECT 4.159 17.976 4.161 20.412 ;
  LAYER M1 ;
        RECT 4.239 17.976 4.241 20.412 ;
  LAYER M1 ;
        RECT 4.319 17.976 4.321 20.412 ;
  LAYER M1 ;
        RECT 4.399 17.976 4.401 20.412 ;
  LAYER M1 ;
        RECT 4.479 17.976 4.481 20.412 ;
  LAYER M1 ;
        RECT 4.559 17.976 4.561 20.412 ;
  LAYER M1 ;
        RECT 4.639 17.976 4.641 20.412 ;
  LAYER M1 ;
        RECT 4.719 17.976 4.721 20.412 ;
  LAYER M1 ;
        RECT 4.799 17.976 4.801 20.412 ;
  LAYER M1 ;
        RECT 4.879 17.976 4.881 20.412 ;
  LAYER M1 ;
        RECT 4.959 17.976 4.961 20.412 ;
  LAYER M1 ;
        RECT 5.039 17.976 5.041 20.412 ;
  LAYER M1 ;
        RECT 5.119 17.976 5.121 20.412 ;
  LAYER M1 ;
        RECT 5.199 17.976 5.201 20.412 ;
  LAYER M1 ;
        RECT 5.279 17.976 5.281 20.412 ;
  LAYER M1 ;
        RECT 5.359 17.976 5.361 20.412 ;
  LAYER M1 ;
        RECT 5.439 17.976 5.441 20.412 ;
  LAYER M1 ;
        RECT 5.519 17.976 5.521 20.412 ;
  LAYER M1 ;
        RECT 5.599 17.976 5.601 20.412 ;
  LAYER M1 ;
        RECT 5.679 17.976 5.681 20.412 ;
  LAYER M1 ;
        RECT 5.759 17.976 5.761 20.412 ;
  LAYER M1 ;
        RECT 5.839 17.976 5.841 20.412 ;
  LAYER M2 ;
        RECT 3.52 17.975 5.92 17.977 ;
  LAYER M2 ;
        RECT 3.52 18.059 5.92 18.061 ;
  LAYER M2 ;
        RECT 3.52 18.143 5.92 18.145 ;
  LAYER M2 ;
        RECT 3.52 18.227 5.92 18.229 ;
  LAYER M2 ;
        RECT 3.52 18.311 5.92 18.313 ;
  LAYER M2 ;
        RECT 3.52 18.395 5.92 18.397 ;
  LAYER M2 ;
        RECT 3.52 18.479 5.92 18.481 ;
  LAYER M2 ;
        RECT 3.52 18.563 5.92 18.565 ;
  LAYER M2 ;
        RECT 3.52 18.647 5.92 18.649 ;
  LAYER M2 ;
        RECT 3.52 18.731 5.92 18.733 ;
  LAYER M2 ;
        RECT 3.52 18.815 5.92 18.817 ;
  LAYER M2 ;
        RECT 3.52 18.899 5.92 18.901 ;
  LAYER M2 ;
        RECT 3.52 18.9825 5.92 18.9845 ;
  LAYER M2 ;
        RECT 3.52 19.067 5.92 19.069 ;
  LAYER M2 ;
        RECT 3.52 19.151 5.92 19.153 ;
  LAYER M2 ;
        RECT 3.52 19.235 5.92 19.237 ;
  LAYER M2 ;
        RECT 3.52 19.319 5.92 19.321 ;
  LAYER M2 ;
        RECT 3.52 19.403 5.92 19.405 ;
  LAYER M2 ;
        RECT 3.52 19.487 5.92 19.489 ;
  LAYER M2 ;
        RECT 3.52 19.571 5.92 19.573 ;
  LAYER M2 ;
        RECT 3.52 19.655 5.92 19.657 ;
  LAYER M2 ;
        RECT 3.52 19.739 5.92 19.741 ;
  LAYER M2 ;
        RECT 3.52 19.823 5.92 19.825 ;
  LAYER M2 ;
        RECT 3.52 19.907 5.92 19.909 ;
  LAYER M2 ;
        RECT 3.52 19.991 5.92 19.993 ;
  LAYER M2 ;
        RECT 3.52 20.075 5.92 20.077 ;
  LAYER M2 ;
        RECT 3.52 20.159 5.92 20.161 ;
  LAYER M2 ;
        RECT 3.52 20.243 5.92 20.245 ;
  LAYER M2 ;
        RECT 3.52 20.327 5.92 20.329 ;
  LAYER M1 ;
        RECT 3.504 20.88 3.536 23.388 ;
  LAYER M1 ;
        RECT 3.568 20.88 3.6 23.388 ;
  LAYER M1 ;
        RECT 3.632 20.88 3.664 23.388 ;
  LAYER M1 ;
        RECT 3.696 20.88 3.728 23.388 ;
  LAYER M1 ;
        RECT 3.76 20.88 3.792 23.388 ;
  LAYER M1 ;
        RECT 3.824 20.88 3.856 23.388 ;
  LAYER M1 ;
        RECT 3.888 20.88 3.92 23.388 ;
  LAYER M1 ;
        RECT 3.952 20.88 3.984 23.388 ;
  LAYER M1 ;
        RECT 4.016 20.88 4.048 23.388 ;
  LAYER M1 ;
        RECT 4.08 20.88 4.112 23.388 ;
  LAYER M1 ;
        RECT 4.144 20.88 4.176 23.388 ;
  LAYER M1 ;
        RECT 4.208 20.88 4.24 23.388 ;
  LAYER M1 ;
        RECT 4.272 20.88 4.304 23.388 ;
  LAYER M1 ;
        RECT 4.336 20.88 4.368 23.388 ;
  LAYER M1 ;
        RECT 4.4 20.88 4.432 23.388 ;
  LAYER M1 ;
        RECT 4.464 20.88 4.496 23.388 ;
  LAYER M1 ;
        RECT 4.528 20.88 4.56 23.388 ;
  LAYER M1 ;
        RECT 4.592 20.88 4.624 23.388 ;
  LAYER M1 ;
        RECT 4.656 20.88 4.688 23.388 ;
  LAYER M1 ;
        RECT 4.72 20.88 4.752 23.388 ;
  LAYER M1 ;
        RECT 4.784 20.88 4.816 23.388 ;
  LAYER M1 ;
        RECT 4.848 20.88 4.88 23.388 ;
  LAYER M1 ;
        RECT 4.912 20.88 4.944 23.388 ;
  LAYER M1 ;
        RECT 4.976 20.88 5.008 23.388 ;
  LAYER M1 ;
        RECT 5.04 20.88 5.072 23.388 ;
  LAYER M1 ;
        RECT 5.104 20.88 5.136 23.388 ;
  LAYER M1 ;
        RECT 5.168 20.88 5.2 23.388 ;
  LAYER M1 ;
        RECT 5.232 20.88 5.264 23.388 ;
  LAYER M1 ;
        RECT 5.296 20.88 5.328 23.388 ;
  LAYER M1 ;
        RECT 5.36 20.88 5.392 23.388 ;
  LAYER M1 ;
        RECT 5.424 20.88 5.456 23.388 ;
  LAYER M1 ;
        RECT 5.488 20.88 5.52 23.388 ;
  LAYER M1 ;
        RECT 5.552 20.88 5.584 23.388 ;
  LAYER M1 ;
        RECT 5.616 20.88 5.648 23.388 ;
  LAYER M1 ;
        RECT 5.68 20.88 5.712 23.388 ;
  LAYER M1 ;
        RECT 5.744 20.88 5.776 23.388 ;
  LAYER M1 ;
        RECT 5.808 20.88 5.84 23.388 ;
  LAYER M2 ;
        RECT 3.484 20.964 5.956 20.996 ;
  LAYER M2 ;
        RECT 3.484 21.028 5.956 21.06 ;
  LAYER M2 ;
        RECT 3.484 21.092 5.956 21.124 ;
  LAYER M2 ;
        RECT 3.484 21.156 5.956 21.188 ;
  LAYER M2 ;
        RECT 3.484 21.22 5.956 21.252 ;
  LAYER M2 ;
        RECT 3.484 21.284 5.956 21.316 ;
  LAYER M2 ;
        RECT 3.484 21.348 5.956 21.38 ;
  LAYER M2 ;
        RECT 3.484 21.412 5.956 21.444 ;
  LAYER M2 ;
        RECT 3.484 21.476 5.956 21.508 ;
  LAYER M2 ;
        RECT 3.484 21.54 5.956 21.572 ;
  LAYER M2 ;
        RECT 3.484 21.604 5.956 21.636 ;
  LAYER M2 ;
        RECT 3.484 21.668 5.956 21.7 ;
  LAYER M2 ;
        RECT 3.484 21.732 5.956 21.764 ;
  LAYER M2 ;
        RECT 3.484 21.796 5.956 21.828 ;
  LAYER M2 ;
        RECT 3.484 21.86 5.956 21.892 ;
  LAYER M2 ;
        RECT 3.484 21.924 5.956 21.956 ;
  LAYER M2 ;
        RECT 3.484 21.988 5.956 22.02 ;
  LAYER M2 ;
        RECT 3.484 22.052 5.956 22.084 ;
  LAYER M2 ;
        RECT 3.484 22.116 5.956 22.148 ;
  LAYER M2 ;
        RECT 3.484 22.18 5.956 22.212 ;
  LAYER M2 ;
        RECT 3.484 22.244 5.956 22.276 ;
  LAYER M2 ;
        RECT 3.484 22.308 5.956 22.34 ;
  LAYER M2 ;
        RECT 3.484 22.372 5.956 22.404 ;
  LAYER M2 ;
        RECT 3.484 22.436 5.956 22.468 ;
  LAYER M2 ;
        RECT 3.484 22.5 5.956 22.532 ;
  LAYER M2 ;
        RECT 3.484 22.564 5.956 22.596 ;
  LAYER M2 ;
        RECT 3.484 22.628 5.956 22.66 ;
  LAYER M2 ;
        RECT 3.484 22.692 5.956 22.724 ;
  LAYER M2 ;
        RECT 3.484 22.756 5.956 22.788 ;
  LAYER M2 ;
        RECT 3.484 22.82 5.956 22.852 ;
  LAYER M2 ;
        RECT 3.484 22.884 5.956 22.916 ;
  LAYER M2 ;
        RECT 3.484 22.948 5.956 22.98 ;
  LAYER M2 ;
        RECT 3.484 23.012 5.956 23.044 ;
  LAYER M2 ;
        RECT 3.484 23.076 5.956 23.108 ;
  LAYER M2 ;
        RECT 3.484 23.14 5.956 23.172 ;
  LAYER M2 ;
        RECT 3.484 23.204 5.956 23.236 ;
  LAYER M3 ;
        RECT 3.504 20.88 3.536 23.388 ;
  LAYER M3 ;
        RECT 3.568 20.88 3.6 23.388 ;
  LAYER M3 ;
        RECT 3.632 20.88 3.664 23.388 ;
  LAYER M3 ;
        RECT 3.696 20.88 3.728 23.388 ;
  LAYER M3 ;
        RECT 3.76 20.88 3.792 23.388 ;
  LAYER M3 ;
        RECT 3.824 20.88 3.856 23.388 ;
  LAYER M3 ;
        RECT 3.888 20.88 3.92 23.388 ;
  LAYER M3 ;
        RECT 3.952 20.88 3.984 23.388 ;
  LAYER M3 ;
        RECT 4.016 20.88 4.048 23.388 ;
  LAYER M3 ;
        RECT 4.08 20.88 4.112 23.388 ;
  LAYER M3 ;
        RECT 4.144 20.88 4.176 23.388 ;
  LAYER M3 ;
        RECT 4.208 20.88 4.24 23.388 ;
  LAYER M3 ;
        RECT 4.272 20.88 4.304 23.388 ;
  LAYER M3 ;
        RECT 4.336 20.88 4.368 23.388 ;
  LAYER M3 ;
        RECT 4.4 20.88 4.432 23.388 ;
  LAYER M3 ;
        RECT 4.464 20.88 4.496 23.388 ;
  LAYER M3 ;
        RECT 4.528 20.88 4.56 23.388 ;
  LAYER M3 ;
        RECT 4.592 20.88 4.624 23.388 ;
  LAYER M3 ;
        RECT 4.656 20.88 4.688 23.388 ;
  LAYER M3 ;
        RECT 4.72 20.88 4.752 23.388 ;
  LAYER M3 ;
        RECT 4.784 20.88 4.816 23.388 ;
  LAYER M3 ;
        RECT 4.848 20.88 4.88 23.388 ;
  LAYER M3 ;
        RECT 4.912 20.88 4.944 23.388 ;
  LAYER M3 ;
        RECT 4.976 20.88 5.008 23.388 ;
  LAYER M3 ;
        RECT 5.04 20.88 5.072 23.388 ;
  LAYER M3 ;
        RECT 5.104 20.88 5.136 23.388 ;
  LAYER M3 ;
        RECT 5.168 20.88 5.2 23.388 ;
  LAYER M3 ;
        RECT 5.232 20.88 5.264 23.388 ;
  LAYER M3 ;
        RECT 5.296 20.88 5.328 23.388 ;
  LAYER M3 ;
        RECT 5.36 20.88 5.392 23.388 ;
  LAYER M3 ;
        RECT 5.424 20.88 5.456 23.388 ;
  LAYER M3 ;
        RECT 5.488 20.88 5.52 23.388 ;
  LAYER M3 ;
        RECT 5.552 20.88 5.584 23.388 ;
  LAYER M3 ;
        RECT 5.616 20.88 5.648 23.388 ;
  LAYER M3 ;
        RECT 5.68 20.88 5.712 23.388 ;
  LAYER M3 ;
        RECT 5.744 20.88 5.776 23.388 ;
  LAYER M3 ;
        RECT 5.808 20.88 5.84 23.388 ;
  LAYER M3 ;
        RECT 5.904 20.88 5.936 23.388 ;
  LAYER M1 ;
        RECT 3.519 20.916 3.521 23.352 ;
  LAYER M1 ;
        RECT 3.599 20.916 3.601 23.352 ;
  LAYER M1 ;
        RECT 3.679 20.916 3.681 23.352 ;
  LAYER M1 ;
        RECT 3.759 20.916 3.761 23.352 ;
  LAYER M1 ;
        RECT 3.839 20.916 3.841 23.352 ;
  LAYER M1 ;
        RECT 3.919 20.916 3.921 23.352 ;
  LAYER M1 ;
        RECT 3.999 20.916 4.001 23.352 ;
  LAYER M1 ;
        RECT 4.079 20.916 4.081 23.352 ;
  LAYER M1 ;
        RECT 4.159 20.916 4.161 23.352 ;
  LAYER M1 ;
        RECT 4.239 20.916 4.241 23.352 ;
  LAYER M1 ;
        RECT 4.319 20.916 4.321 23.352 ;
  LAYER M1 ;
        RECT 4.399 20.916 4.401 23.352 ;
  LAYER M1 ;
        RECT 4.479 20.916 4.481 23.352 ;
  LAYER M1 ;
        RECT 4.559 20.916 4.561 23.352 ;
  LAYER M1 ;
        RECT 4.639 20.916 4.641 23.352 ;
  LAYER M1 ;
        RECT 4.719 20.916 4.721 23.352 ;
  LAYER M1 ;
        RECT 4.799 20.916 4.801 23.352 ;
  LAYER M1 ;
        RECT 4.879 20.916 4.881 23.352 ;
  LAYER M1 ;
        RECT 4.959 20.916 4.961 23.352 ;
  LAYER M1 ;
        RECT 5.039 20.916 5.041 23.352 ;
  LAYER M1 ;
        RECT 5.119 20.916 5.121 23.352 ;
  LAYER M1 ;
        RECT 5.199 20.916 5.201 23.352 ;
  LAYER M1 ;
        RECT 5.279 20.916 5.281 23.352 ;
  LAYER M1 ;
        RECT 5.359 20.916 5.361 23.352 ;
  LAYER M1 ;
        RECT 5.439 20.916 5.441 23.352 ;
  LAYER M1 ;
        RECT 5.519 20.916 5.521 23.352 ;
  LAYER M1 ;
        RECT 5.599 20.916 5.601 23.352 ;
  LAYER M1 ;
        RECT 5.679 20.916 5.681 23.352 ;
  LAYER M1 ;
        RECT 5.759 20.916 5.761 23.352 ;
  LAYER M1 ;
        RECT 5.839 20.916 5.841 23.352 ;
  LAYER M2 ;
        RECT 3.52 20.915 5.92 20.917 ;
  LAYER M2 ;
        RECT 3.52 20.999 5.92 21.001 ;
  LAYER M2 ;
        RECT 3.52 21.083 5.92 21.085 ;
  LAYER M2 ;
        RECT 3.52 21.167 5.92 21.169 ;
  LAYER M2 ;
        RECT 3.52 21.251 5.92 21.253 ;
  LAYER M2 ;
        RECT 3.52 21.335 5.92 21.337 ;
  LAYER M2 ;
        RECT 3.52 21.419 5.92 21.421 ;
  LAYER M2 ;
        RECT 3.52 21.503 5.92 21.505 ;
  LAYER M2 ;
        RECT 3.52 21.587 5.92 21.589 ;
  LAYER M2 ;
        RECT 3.52 21.671 5.92 21.673 ;
  LAYER M2 ;
        RECT 3.52 21.755 5.92 21.757 ;
  LAYER M2 ;
        RECT 3.52 21.839 5.92 21.841 ;
  LAYER M2 ;
        RECT 3.52 21.9225 5.92 21.9245 ;
  LAYER M2 ;
        RECT 3.52 22.007 5.92 22.009 ;
  LAYER M2 ;
        RECT 3.52 22.091 5.92 22.093 ;
  LAYER M2 ;
        RECT 3.52 22.175 5.92 22.177 ;
  LAYER M2 ;
        RECT 3.52 22.259 5.92 22.261 ;
  LAYER M2 ;
        RECT 3.52 22.343 5.92 22.345 ;
  LAYER M2 ;
        RECT 3.52 22.427 5.92 22.429 ;
  LAYER M2 ;
        RECT 3.52 22.511 5.92 22.513 ;
  LAYER M2 ;
        RECT 3.52 22.595 5.92 22.597 ;
  LAYER M2 ;
        RECT 3.52 22.679 5.92 22.681 ;
  LAYER M2 ;
        RECT 3.52 22.763 5.92 22.765 ;
  LAYER M2 ;
        RECT 3.52 22.847 5.92 22.849 ;
  LAYER M2 ;
        RECT 3.52 22.931 5.92 22.933 ;
  LAYER M2 ;
        RECT 3.52 23.015 5.92 23.017 ;
  LAYER M2 ;
        RECT 3.52 23.099 5.92 23.101 ;
  LAYER M2 ;
        RECT 3.52 23.183 5.92 23.185 ;
  LAYER M2 ;
        RECT 3.52 23.267 5.92 23.269 ;
  LAYER M1 ;
        RECT 3.504 23.82 3.536 26.328 ;
  LAYER M1 ;
        RECT 3.568 23.82 3.6 26.328 ;
  LAYER M1 ;
        RECT 3.632 23.82 3.664 26.328 ;
  LAYER M1 ;
        RECT 3.696 23.82 3.728 26.328 ;
  LAYER M1 ;
        RECT 3.76 23.82 3.792 26.328 ;
  LAYER M1 ;
        RECT 3.824 23.82 3.856 26.328 ;
  LAYER M1 ;
        RECT 3.888 23.82 3.92 26.328 ;
  LAYER M1 ;
        RECT 3.952 23.82 3.984 26.328 ;
  LAYER M1 ;
        RECT 4.016 23.82 4.048 26.328 ;
  LAYER M1 ;
        RECT 4.08 23.82 4.112 26.328 ;
  LAYER M1 ;
        RECT 4.144 23.82 4.176 26.328 ;
  LAYER M1 ;
        RECT 4.208 23.82 4.24 26.328 ;
  LAYER M1 ;
        RECT 4.272 23.82 4.304 26.328 ;
  LAYER M1 ;
        RECT 4.336 23.82 4.368 26.328 ;
  LAYER M1 ;
        RECT 4.4 23.82 4.432 26.328 ;
  LAYER M1 ;
        RECT 4.464 23.82 4.496 26.328 ;
  LAYER M1 ;
        RECT 4.528 23.82 4.56 26.328 ;
  LAYER M1 ;
        RECT 4.592 23.82 4.624 26.328 ;
  LAYER M1 ;
        RECT 4.656 23.82 4.688 26.328 ;
  LAYER M1 ;
        RECT 4.72 23.82 4.752 26.328 ;
  LAYER M1 ;
        RECT 4.784 23.82 4.816 26.328 ;
  LAYER M1 ;
        RECT 4.848 23.82 4.88 26.328 ;
  LAYER M1 ;
        RECT 4.912 23.82 4.944 26.328 ;
  LAYER M1 ;
        RECT 4.976 23.82 5.008 26.328 ;
  LAYER M1 ;
        RECT 5.04 23.82 5.072 26.328 ;
  LAYER M1 ;
        RECT 5.104 23.82 5.136 26.328 ;
  LAYER M1 ;
        RECT 5.168 23.82 5.2 26.328 ;
  LAYER M1 ;
        RECT 5.232 23.82 5.264 26.328 ;
  LAYER M1 ;
        RECT 5.296 23.82 5.328 26.328 ;
  LAYER M1 ;
        RECT 5.36 23.82 5.392 26.328 ;
  LAYER M1 ;
        RECT 5.424 23.82 5.456 26.328 ;
  LAYER M1 ;
        RECT 5.488 23.82 5.52 26.328 ;
  LAYER M1 ;
        RECT 5.552 23.82 5.584 26.328 ;
  LAYER M1 ;
        RECT 5.616 23.82 5.648 26.328 ;
  LAYER M1 ;
        RECT 5.68 23.82 5.712 26.328 ;
  LAYER M1 ;
        RECT 5.744 23.82 5.776 26.328 ;
  LAYER M1 ;
        RECT 5.808 23.82 5.84 26.328 ;
  LAYER M2 ;
        RECT 3.484 23.904 5.956 23.936 ;
  LAYER M2 ;
        RECT 3.484 23.968 5.956 24 ;
  LAYER M2 ;
        RECT 3.484 24.032 5.956 24.064 ;
  LAYER M2 ;
        RECT 3.484 24.096 5.956 24.128 ;
  LAYER M2 ;
        RECT 3.484 24.16 5.956 24.192 ;
  LAYER M2 ;
        RECT 3.484 24.224 5.956 24.256 ;
  LAYER M2 ;
        RECT 3.484 24.288 5.956 24.32 ;
  LAYER M2 ;
        RECT 3.484 24.352 5.956 24.384 ;
  LAYER M2 ;
        RECT 3.484 24.416 5.956 24.448 ;
  LAYER M2 ;
        RECT 3.484 24.48 5.956 24.512 ;
  LAYER M2 ;
        RECT 3.484 24.544 5.956 24.576 ;
  LAYER M2 ;
        RECT 3.484 24.608 5.956 24.64 ;
  LAYER M2 ;
        RECT 3.484 24.672 5.956 24.704 ;
  LAYER M2 ;
        RECT 3.484 24.736 5.956 24.768 ;
  LAYER M2 ;
        RECT 3.484 24.8 5.956 24.832 ;
  LAYER M2 ;
        RECT 3.484 24.864 5.956 24.896 ;
  LAYER M2 ;
        RECT 3.484 24.928 5.956 24.96 ;
  LAYER M2 ;
        RECT 3.484 24.992 5.956 25.024 ;
  LAYER M2 ;
        RECT 3.484 25.056 5.956 25.088 ;
  LAYER M2 ;
        RECT 3.484 25.12 5.956 25.152 ;
  LAYER M2 ;
        RECT 3.484 25.184 5.956 25.216 ;
  LAYER M2 ;
        RECT 3.484 25.248 5.956 25.28 ;
  LAYER M2 ;
        RECT 3.484 25.312 5.956 25.344 ;
  LAYER M2 ;
        RECT 3.484 25.376 5.956 25.408 ;
  LAYER M2 ;
        RECT 3.484 25.44 5.956 25.472 ;
  LAYER M2 ;
        RECT 3.484 25.504 5.956 25.536 ;
  LAYER M2 ;
        RECT 3.484 25.568 5.956 25.6 ;
  LAYER M2 ;
        RECT 3.484 25.632 5.956 25.664 ;
  LAYER M2 ;
        RECT 3.484 25.696 5.956 25.728 ;
  LAYER M2 ;
        RECT 3.484 25.76 5.956 25.792 ;
  LAYER M2 ;
        RECT 3.484 25.824 5.956 25.856 ;
  LAYER M2 ;
        RECT 3.484 25.888 5.956 25.92 ;
  LAYER M2 ;
        RECT 3.484 25.952 5.956 25.984 ;
  LAYER M2 ;
        RECT 3.484 26.016 5.956 26.048 ;
  LAYER M2 ;
        RECT 3.484 26.08 5.956 26.112 ;
  LAYER M2 ;
        RECT 3.484 26.144 5.956 26.176 ;
  LAYER M3 ;
        RECT 3.504 23.82 3.536 26.328 ;
  LAYER M3 ;
        RECT 3.568 23.82 3.6 26.328 ;
  LAYER M3 ;
        RECT 3.632 23.82 3.664 26.328 ;
  LAYER M3 ;
        RECT 3.696 23.82 3.728 26.328 ;
  LAYER M3 ;
        RECT 3.76 23.82 3.792 26.328 ;
  LAYER M3 ;
        RECT 3.824 23.82 3.856 26.328 ;
  LAYER M3 ;
        RECT 3.888 23.82 3.92 26.328 ;
  LAYER M3 ;
        RECT 3.952 23.82 3.984 26.328 ;
  LAYER M3 ;
        RECT 4.016 23.82 4.048 26.328 ;
  LAYER M3 ;
        RECT 4.08 23.82 4.112 26.328 ;
  LAYER M3 ;
        RECT 4.144 23.82 4.176 26.328 ;
  LAYER M3 ;
        RECT 4.208 23.82 4.24 26.328 ;
  LAYER M3 ;
        RECT 4.272 23.82 4.304 26.328 ;
  LAYER M3 ;
        RECT 4.336 23.82 4.368 26.328 ;
  LAYER M3 ;
        RECT 4.4 23.82 4.432 26.328 ;
  LAYER M3 ;
        RECT 4.464 23.82 4.496 26.328 ;
  LAYER M3 ;
        RECT 4.528 23.82 4.56 26.328 ;
  LAYER M3 ;
        RECT 4.592 23.82 4.624 26.328 ;
  LAYER M3 ;
        RECT 4.656 23.82 4.688 26.328 ;
  LAYER M3 ;
        RECT 4.72 23.82 4.752 26.328 ;
  LAYER M3 ;
        RECT 4.784 23.82 4.816 26.328 ;
  LAYER M3 ;
        RECT 4.848 23.82 4.88 26.328 ;
  LAYER M3 ;
        RECT 4.912 23.82 4.944 26.328 ;
  LAYER M3 ;
        RECT 4.976 23.82 5.008 26.328 ;
  LAYER M3 ;
        RECT 5.04 23.82 5.072 26.328 ;
  LAYER M3 ;
        RECT 5.104 23.82 5.136 26.328 ;
  LAYER M3 ;
        RECT 5.168 23.82 5.2 26.328 ;
  LAYER M3 ;
        RECT 5.232 23.82 5.264 26.328 ;
  LAYER M3 ;
        RECT 5.296 23.82 5.328 26.328 ;
  LAYER M3 ;
        RECT 5.36 23.82 5.392 26.328 ;
  LAYER M3 ;
        RECT 5.424 23.82 5.456 26.328 ;
  LAYER M3 ;
        RECT 5.488 23.82 5.52 26.328 ;
  LAYER M3 ;
        RECT 5.552 23.82 5.584 26.328 ;
  LAYER M3 ;
        RECT 5.616 23.82 5.648 26.328 ;
  LAYER M3 ;
        RECT 5.68 23.82 5.712 26.328 ;
  LAYER M3 ;
        RECT 5.744 23.82 5.776 26.328 ;
  LAYER M3 ;
        RECT 5.808 23.82 5.84 26.328 ;
  LAYER M3 ;
        RECT 5.904 23.82 5.936 26.328 ;
  LAYER M1 ;
        RECT 3.519 23.856 3.521 26.292 ;
  LAYER M1 ;
        RECT 3.599 23.856 3.601 26.292 ;
  LAYER M1 ;
        RECT 3.679 23.856 3.681 26.292 ;
  LAYER M1 ;
        RECT 3.759 23.856 3.761 26.292 ;
  LAYER M1 ;
        RECT 3.839 23.856 3.841 26.292 ;
  LAYER M1 ;
        RECT 3.919 23.856 3.921 26.292 ;
  LAYER M1 ;
        RECT 3.999 23.856 4.001 26.292 ;
  LAYER M1 ;
        RECT 4.079 23.856 4.081 26.292 ;
  LAYER M1 ;
        RECT 4.159 23.856 4.161 26.292 ;
  LAYER M1 ;
        RECT 4.239 23.856 4.241 26.292 ;
  LAYER M1 ;
        RECT 4.319 23.856 4.321 26.292 ;
  LAYER M1 ;
        RECT 4.399 23.856 4.401 26.292 ;
  LAYER M1 ;
        RECT 4.479 23.856 4.481 26.292 ;
  LAYER M1 ;
        RECT 4.559 23.856 4.561 26.292 ;
  LAYER M1 ;
        RECT 4.639 23.856 4.641 26.292 ;
  LAYER M1 ;
        RECT 4.719 23.856 4.721 26.292 ;
  LAYER M1 ;
        RECT 4.799 23.856 4.801 26.292 ;
  LAYER M1 ;
        RECT 4.879 23.856 4.881 26.292 ;
  LAYER M1 ;
        RECT 4.959 23.856 4.961 26.292 ;
  LAYER M1 ;
        RECT 5.039 23.856 5.041 26.292 ;
  LAYER M1 ;
        RECT 5.119 23.856 5.121 26.292 ;
  LAYER M1 ;
        RECT 5.199 23.856 5.201 26.292 ;
  LAYER M1 ;
        RECT 5.279 23.856 5.281 26.292 ;
  LAYER M1 ;
        RECT 5.359 23.856 5.361 26.292 ;
  LAYER M1 ;
        RECT 5.439 23.856 5.441 26.292 ;
  LAYER M1 ;
        RECT 5.519 23.856 5.521 26.292 ;
  LAYER M1 ;
        RECT 5.599 23.856 5.601 26.292 ;
  LAYER M1 ;
        RECT 5.679 23.856 5.681 26.292 ;
  LAYER M1 ;
        RECT 5.759 23.856 5.761 26.292 ;
  LAYER M1 ;
        RECT 5.839 23.856 5.841 26.292 ;
  LAYER M2 ;
        RECT 3.52 23.855 5.92 23.857 ;
  LAYER M2 ;
        RECT 3.52 23.939 5.92 23.941 ;
  LAYER M2 ;
        RECT 3.52 24.023 5.92 24.025 ;
  LAYER M2 ;
        RECT 3.52 24.107 5.92 24.109 ;
  LAYER M2 ;
        RECT 3.52 24.191 5.92 24.193 ;
  LAYER M2 ;
        RECT 3.52 24.275 5.92 24.277 ;
  LAYER M2 ;
        RECT 3.52 24.359 5.92 24.361 ;
  LAYER M2 ;
        RECT 3.52 24.443 5.92 24.445 ;
  LAYER M2 ;
        RECT 3.52 24.527 5.92 24.529 ;
  LAYER M2 ;
        RECT 3.52 24.611 5.92 24.613 ;
  LAYER M2 ;
        RECT 3.52 24.695 5.92 24.697 ;
  LAYER M2 ;
        RECT 3.52 24.779 5.92 24.781 ;
  LAYER M2 ;
        RECT 3.52 24.8625 5.92 24.8645 ;
  LAYER M2 ;
        RECT 3.52 24.947 5.92 24.949 ;
  LAYER M2 ;
        RECT 3.52 25.031 5.92 25.033 ;
  LAYER M2 ;
        RECT 3.52 25.115 5.92 25.117 ;
  LAYER M2 ;
        RECT 3.52 25.199 5.92 25.201 ;
  LAYER M2 ;
        RECT 3.52 25.283 5.92 25.285 ;
  LAYER M2 ;
        RECT 3.52 25.367 5.92 25.369 ;
  LAYER M2 ;
        RECT 3.52 25.451 5.92 25.453 ;
  LAYER M2 ;
        RECT 3.52 25.535 5.92 25.537 ;
  LAYER M2 ;
        RECT 3.52 25.619 5.92 25.621 ;
  LAYER M2 ;
        RECT 3.52 25.703 5.92 25.705 ;
  LAYER M2 ;
        RECT 3.52 25.787 5.92 25.789 ;
  LAYER M2 ;
        RECT 3.52 25.871 5.92 25.873 ;
  LAYER M2 ;
        RECT 3.52 25.955 5.92 25.957 ;
  LAYER M2 ;
        RECT 3.52 26.039 5.92 26.041 ;
  LAYER M2 ;
        RECT 3.52 26.123 5.92 26.125 ;
  LAYER M2 ;
        RECT 3.52 26.207 5.92 26.209 ;
  LAYER M1 ;
        RECT 3.504 26.76 3.536 29.268 ;
  LAYER M1 ;
        RECT 3.568 26.76 3.6 29.268 ;
  LAYER M1 ;
        RECT 3.632 26.76 3.664 29.268 ;
  LAYER M1 ;
        RECT 3.696 26.76 3.728 29.268 ;
  LAYER M1 ;
        RECT 3.76 26.76 3.792 29.268 ;
  LAYER M1 ;
        RECT 3.824 26.76 3.856 29.268 ;
  LAYER M1 ;
        RECT 3.888 26.76 3.92 29.268 ;
  LAYER M1 ;
        RECT 3.952 26.76 3.984 29.268 ;
  LAYER M1 ;
        RECT 4.016 26.76 4.048 29.268 ;
  LAYER M1 ;
        RECT 4.08 26.76 4.112 29.268 ;
  LAYER M1 ;
        RECT 4.144 26.76 4.176 29.268 ;
  LAYER M1 ;
        RECT 4.208 26.76 4.24 29.268 ;
  LAYER M1 ;
        RECT 4.272 26.76 4.304 29.268 ;
  LAYER M1 ;
        RECT 4.336 26.76 4.368 29.268 ;
  LAYER M1 ;
        RECT 4.4 26.76 4.432 29.268 ;
  LAYER M1 ;
        RECT 4.464 26.76 4.496 29.268 ;
  LAYER M1 ;
        RECT 4.528 26.76 4.56 29.268 ;
  LAYER M1 ;
        RECT 4.592 26.76 4.624 29.268 ;
  LAYER M1 ;
        RECT 4.656 26.76 4.688 29.268 ;
  LAYER M1 ;
        RECT 4.72 26.76 4.752 29.268 ;
  LAYER M1 ;
        RECT 4.784 26.76 4.816 29.268 ;
  LAYER M1 ;
        RECT 4.848 26.76 4.88 29.268 ;
  LAYER M1 ;
        RECT 4.912 26.76 4.944 29.268 ;
  LAYER M1 ;
        RECT 4.976 26.76 5.008 29.268 ;
  LAYER M1 ;
        RECT 5.04 26.76 5.072 29.268 ;
  LAYER M1 ;
        RECT 5.104 26.76 5.136 29.268 ;
  LAYER M1 ;
        RECT 5.168 26.76 5.2 29.268 ;
  LAYER M1 ;
        RECT 5.232 26.76 5.264 29.268 ;
  LAYER M1 ;
        RECT 5.296 26.76 5.328 29.268 ;
  LAYER M1 ;
        RECT 5.36 26.76 5.392 29.268 ;
  LAYER M1 ;
        RECT 5.424 26.76 5.456 29.268 ;
  LAYER M1 ;
        RECT 5.488 26.76 5.52 29.268 ;
  LAYER M1 ;
        RECT 5.552 26.76 5.584 29.268 ;
  LAYER M1 ;
        RECT 5.616 26.76 5.648 29.268 ;
  LAYER M1 ;
        RECT 5.68 26.76 5.712 29.268 ;
  LAYER M1 ;
        RECT 5.744 26.76 5.776 29.268 ;
  LAYER M1 ;
        RECT 5.808 26.76 5.84 29.268 ;
  LAYER M2 ;
        RECT 3.484 26.844 5.956 26.876 ;
  LAYER M2 ;
        RECT 3.484 26.908 5.956 26.94 ;
  LAYER M2 ;
        RECT 3.484 26.972 5.956 27.004 ;
  LAYER M2 ;
        RECT 3.484 27.036 5.956 27.068 ;
  LAYER M2 ;
        RECT 3.484 27.1 5.956 27.132 ;
  LAYER M2 ;
        RECT 3.484 27.164 5.956 27.196 ;
  LAYER M2 ;
        RECT 3.484 27.228 5.956 27.26 ;
  LAYER M2 ;
        RECT 3.484 27.292 5.956 27.324 ;
  LAYER M2 ;
        RECT 3.484 27.356 5.956 27.388 ;
  LAYER M2 ;
        RECT 3.484 27.42 5.956 27.452 ;
  LAYER M2 ;
        RECT 3.484 27.484 5.956 27.516 ;
  LAYER M2 ;
        RECT 3.484 27.548 5.956 27.58 ;
  LAYER M2 ;
        RECT 3.484 27.612 5.956 27.644 ;
  LAYER M2 ;
        RECT 3.484 27.676 5.956 27.708 ;
  LAYER M2 ;
        RECT 3.484 27.74 5.956 27.772 ;
  LAYER M2 ;
        RECT 3.484 27.804 5.956 27.836 ;
  LAYER M2 ;
        RECT 3.484 27.868 5.956 27.9 ;
  LAYER M2 ;
        RECT 3.484 27.932 5.956 27.964 ;
  LAYER M2 ;
        RECT 3.484 27.996 5.956 28.028 ;
  LAYER M2 ;
        RECT 3.484 28.06 5.956 28.092 ;
  LAYER M2 ;
        RECT 3.484 28.124 5.956 28.156 ;
  LAYER M2 ;
        RECT 3.484 28.188 5.956 28.22 ;
  LAYER M2 ;
        RECT 3.484 28.252 5.956 28.284 ;
  LAYER M2 ;
        RECT 3.484 28.316 5.956 28.348 ;
  LAYER M2 ;
        RECT 3.484 28.38 5.956 28.412 ;
  LAYER M2 ;
        RECT 3.484 28.444 5.956 28.476 ;
  LAYER M2 ;
        RECT 3.484 28.508 5.956 28.54 ;
  LAYER M2 ;
        RECT 3.484 28.572 5.956 28.604 ;
  LAYER M2 ;
        RECT 3.484 28.636 5.956 28.668 ;
  LAYER M2 ;
        RECT 3.484 28.7 5.956 28.732 ;
  LAYER M2 ;
        RECT 3.484 28.764 5.956 28.796 ;
  LAYER M2 ;
        RECT 3.484 28.828 5.956 28.86 ;
  LAYER M2 ;
        RECT 3.484 28.892 5.956 28.924 ;
  LAYER M2 ;
        RECT 3.484 28.956 5.956 28.988 ;
  LAYER M2 ;
        RECT 3.484 29.02 5.956 29.052 ;
  LAYER M2 ;
        RECT 3.484 29.084 5.956 29.116 ;
  LAYER M3 ;
        RECT 3.504 26.76 3.536 29.268 ;
  LAYER M3 ;
        RECT 3.568 26.76 3.6 29.268 ;
  LAYER M3 ;
        RECT 3.632 26.76 3.664 29.268 ;
  LAYER M3 ;
        RECT 3.696 26.76 3.728 29.268 ;
  LAYER M3 ;
        RECT 3.76 26.76 3.792 29.268 ;
  LAYER M3 ;
        RECT 3.824 26.76 3.856 29.268 ;
  LAYER M3 ;
        RECT 3.888 26.76 3.92 29.268 ;
  LAYER M3 ;
        RECT 3.952 26.76 3.984 29.268 ;
  LAYER M3 ;
        RECT 4.016 26.76 4.048 29.268 ;
  LAYER M3 ;
        RECT 4.08 26.76 4.112 29.268 ;
  LAYER M3 ;
        RECT 4.144 26.76 4.176 29.268 ;
  LAYER M3 ;
        RECT 4.208 26.76 4.24 29.268 ;
  LAYER M3 ;
        RECT 4.272 26.76 4.304 29.268 ;
  LAYER M3 ;
        RECT 4.336 26.76 4.368 29.268 ;
  LAYER M3 ;
        RECT 4.4 26.76 4.432 29.268 ;
  LAYER M3 ;
        RECT 4.464 26.76 4.496 29.268 ;
  LAYER M3 ;
        RECT 4.528 26.76 4.56 29.268 ;
  LAYER M3 ;
        RECT 4.592 26.76 4.624 29.268 ;
  LAYER M3 ;
        RECT 4.656 26.76 4.688 29.268 ;
  LAYER M3 ;
        RECT 4.72 26.76 4.752 29.268 ;
  LAYER M3 ;
        RECT 4.784 26.76 4.816 29.268 ;
  LAYER M3 ;
        RECT 4.848 26.76 4.88 29.268 ;
  LAYER M3 ;
        RECT 4.912 26.76 4.944 29.268 ;
  LAYER M3 ;
        RECT 4.976 26.76 5.008 29.268 ;
  LAYER M3 ;
        RECT 5.04 26.76 5.072 29.268 ;
  LAYER M3 ;
        RECT 5.104 26.76 5.136 29.268 ;
  LAYER M3 ;
        RECT 5.168 26.76 5.2 29.268 ;
  LAYER M3 ;
        RECT 5.232 26.76 5.264 29.268 ;
  LAYER M3 ;
        RECT 5.296 26.76 5.328 29.268 ;
  LAYER M3 ;
        RECT 5.36 26.76 5.392 29.268 ;
  LAYER M3 ;
        RECT 5.424 26.76 5.456 29.268 ;
  LAYER M3 ;
        RECT 5.488 26.76 5.52 29.268 ;
  LAYER M3 ;
        RECT 5.552 26.76 5.584 29.268 ;
  LAYER M3 ;
        RECT 5.616 26.76 5.648 29.268 ;
  LAYER M3 ;
        RECT 5.68 26.76 5.712 29.268 ;
  LAYER M3 ;
        RECT 5.744 26.76 5.776 29.268 ;
  LAYER M3 ;
        RECT 5.808 26.76 5.84 29.268 ;
  LAYER M3 ;
        RECT 5.904 26.76 5.936 29.268 ;
  LAYER M1 ;
        RECT 3.519 26.796 3.521 29.232 ;
  LAYER M1 ;
        RECT 3.599 26.796 3.601 29.232 ;
  LAYER M1 ;
        RECT 3.679 26.796 3.681 29.232 ;
  LAYER M1 ;
        RECT 3.759 26.796 3.761 29.232 ;
  LAYER M1 ;
        RECT 3.839 26.796 3.841 29.232 ;
  LAYER M1 ;
        RECT 3.919 26.796 3.921 29.232 ;
  LAYER M1 ;
        RECT 3.999 26.796 4.001 29.232 ;
  LAYER M1 ;
        RECT 4.079 26.796 4.081 29.232 ;
  LAYER M1 ;
        RECT 4.159 26.796 4.161 29.232 ;
  LAYER M1 ;
        RECT 4.239 26.796 4.241 29.232 ;
  LAYER M1 ;
        RECT 4.319 26.796 4.321 29.232 ;
  LAYER M1 ;
        RECT 4.399 26.796 4.401 29.232 ;
  LAYER M1 ;
        RECT 4.479 26.796 4.481 29.232 ;
  LAYER M1 ;
        RECT 4.559 26.796 4.561 29.232 ;
  LAYER M1 ;
        RECT 4.639 26.796 4.641 29.232 ;
  LAYER M1 ;
        RECT 4.719 26.796 4.721 29.232 ;
  LAYER M1 ;
        RECT 4.799 26.796 4.801 29.232 ;
  LAYER M1 ;
        RECT 4.879 26.796 4.881 29.232 ;
  LAYER M1 ;
        RECT 4.959 26.796 4.961 29.232 ;
  LAYER M1 ;
        RECT 5.039 26.796 5.041 29.232 ;
  LAYER M1 ;
        RECT 5.119 26.796 5.121 29.232 ;
  LAYER M1 ;
        RECT 5.199 26.796 5.201 29.232 ;
  LAYER M1 ;
        RECT 5.279 26.796 5.281 29.232 ;
  LAYER M1 ;
        RECT 5.359 26.796 5.361 29.232 ;
  LAYER M1 ;
        RECT 5.439 26.796 5.441 29.232 ;
  LAYER M1 ;
        RECT 5.519 26.796 5.521 29.232 ;
  LAYER M1 ;
        RECT 5.599 26.796 5.601 29.232 ;
  LAYER M1 ;
        RECT 5.679 26.796 5.681 29.232 ;
  LAYER M1 ;
        RECT 5.759 26.796 5.761 29.232 ;
  LAYER M1 ;
        RECT 5.839 26.796 5.841 29.232 ;
  LAYER M2 ;
        RECT 3.52 26.795 5.92 26.797 ;
  LAYER M2 ;
        RECT 3.52 26.879 5.92 26.881 ;
  LAYER M2 ;
        RECT 3.52 26.963 5.92 26.965 ;
  LAYER M2 ;
        RECT 3.52 27.047 5.92 27.049 ;
  LAYER M2 ;
        RECT 3.52 27.131 5.92 27.133 ;
  LAYER M2 ;
        RECT 3.52 27.215 5.92 27.217 ;
  LAYER M2 ;
        RECT 3.52 27.299 5.92 27.301 ;
  LAYER M2 ;
        RECT 3.52 27.383 5.92 27.385 ;
  LAYER M2 ;
        RECT 3.52 27.467 5.92 27.469 ;
  LAYER M2 ;
        RECT 3.52 27.551 5.92 27.553 ;
  LAYER M2 ;
        RECT 3.52 27.635 5.92 27.637 ;
  LAYER M2 ;
        RECT 3.52 27.719 5.92 27.721 ;
  LAYER M2 ;
        RECT 3.52 27.8025 5.92 27.8045 ;
  LAYER M2 ;
        RECT 3.52 27.887 5.92 27.889 ;
  LAYER M2 ;
        RECT 3.52 27.971 5.92 27.973 ;
  LAYER M2 ;
        RECT 3.52 28.055 5.92 28.057 ;
  LAYER M2 ;
        RECT 3.52 28.139 5.92 28.141 ;
  LAYER M2 ;
        RECT 3.52 28.223 5.92 28.225 ;
  LAYER M2 ;
        RECT 3.52 28.307 5.92 28.309 ;
  LAYER M2 ;
        RECT 3.52 28.391 5.92 28.393 ;
  LAYER M2 ;
        RECT 3.52 28.475 5.92 28.477 ;
  LAYER M2 ;
        RECT 3.52 28.559 5.92 28.561 ;
  LAYER M2 ;
        RECT 3.52 28.643 5.92 28.645 ;
  LAYER M2 ;
        RECT 3.52 28.727 5.92 28.729 ;
  LAYER M2 ;
        RECT 3.52 28.811 5.92 28.813 ;
  LAYER M2 ;
        RECT 3.52 28.895 5.92 28.897 ;
  LAYER M2 ;
        RECT 3.52 28.979 5.92 28.981 ;
  LAYER M2 ;
        RECT 3.52 29.063 5.92 29.065 ;
  LAYER M2 ;
        RECT 3.52 29.147 5.92 29.149 ;
  LAYER M1 ;
        RECT 6.384 17.94 6.416 20.448 ;
  LAYER M1 ;
        RECT 6.448 17.94 6.48 20.448 ;
  LAYER M1 ;
        RECT 6.512 17.94 6.544 20.448 ;
  LAYER M1 ;
        RECT 6.576 17.94 6.608 20.448 ;
  LAYER M1 ;
        RECT 6.64 17.94 6.672 20.448 ;
  LAYER M1 ;
        RECT 6.704 17.94 6.736 20.448 ;
  LAYER M1 ;
        RECT 6.768 17.94 6.8 20.448 ;
  LAYER M1 ;
        RECT 6.832 17.94 6.864 20.448 ;
  LAYER M1 ;
        RECT 6.896 17.94 6.928 20.448 ;
  LAYER M1 ;
        RECT 6.96 17.94 6.992 20.448 ;
  LAYER M1 ;
        RECT 7.024 17.94 7.056 20.448 ;
  LAYER M1 ;
        RECT 7.088 17.94 7.12 20.448 ;
  LAYER M1 ;
        RECT 7.152 17.94 7.184 20.448 ;
  LAYER M1 ;
        RECT 7.216 17.94 7.248 20.448 ;
  LAYER M1 ;
        RECT 7.28 17.94 7.312 20.448 ;
  LAYER M1 ;
        RECT 7.344 17.94 7.376 20.448 ;
  LAYER M1 ;
        RECT 7.408 17.94 7.44 20.448 ;
  LAYER M1 ;
        RECT 7.472 17.94 7.504 20.448 ;
  LAYER M1 ;
        RECT 7.536 17.94 7.568 20.448 ;
  LAYER M1 ;
        RECT 7.6 17.94 7.632 20.448 ;
  LAYER M1 ;
        RECT 7.664 17.94 7.696 20.448 ;
  LAYER M1 ;
        RECT 7.728 17.94 7.76 20.448 ;
  LAYER M1 ;
        RECT 7.792 17.94 7.824 20.448 ;
  LAYER M1 ;
        RECT 7.856 17.94 7.888 20.448 ;
  LAYER M1 ;
        RECT 7.92 17.94 7.952 20.448 ;
  LAYER M1 ;
        RECT 7.984 17.94 8.016 20.448 ;
  LAYER M1 ;
        RECT 8.048 17.94 8.08 20.448 ;
  LAYER M1 ;
        RECT 8.112 17.94 8.144 20.448 ;
  LAYER M1 ;
        RECT 8.176 17.94 8.208 20.448 ;
  LAYER M1 ;
        RECT 8.24 17.94 8.272 20.448 ;
  LAYER M1 ;
        RECT 8.304 17.94 8.336 20.448 ;
  LAYER M1 ;
        RECT 8.368 17.94 8.4 20.448 ;
  LAYER M1 ;
        RECT 8.432 17.94 8.464 20.448 ;
  LAYER M1 ;
        RECT 8.496 17.94 8.528 20.448 ;
  LAYER M1 ;
        RECT 8.56 17.94 8.592 20.448 ;
  LAYER M1 ;
        RECT 8.624 17.94 8.656 20.448 ;
  LAYER M1 ;
        RECT 8.688 17.94 8.72 20.448 ;
  LAYER M2 ;
        RECT 6.364 18.024 8.836 18.056 ;
  LAYER M2 ;
        RECT 6.364 18.088 8.836 18.12 ;
  LAYER M2 ;
        RECT 6.364 18.152 8.836 18.184 ;
  LAYER M2 ;
        RECT 6.364 18.216 8.836 18.248 ;
  LAYER M2 ;
        RECT 6.364 18.28 8.836 18.312 ;
  LAYER M2 ;
        RECT 6.364 18.344 8.836 18.376 ;
  LAYER M2 ;
        RECT 6.364 18.408 8.836 18.44 ;
  LAYER M2 ;
        RECT 6.364 18.472 8.836 18.504 ;
  LAYER M2 ;
        RECT 6.364 18.536 8.836 18.568 ;
  LAYER M2 ;
        RECT 6.364 18.6 8.836 18.632 ;
  LAYER M2 ;
        RECT 6.364 18.664 8.836 18.696 ;
  LAYER M2 ;
        RECT 6.364 18.728 8.836 18.76 ;
  LAYER M2 ;
        RECT 6.364 18.792 8.836 18.824 ;
  LAYER M2 ;
        RECT 6.364 18.856 8.836 18.888 ;
  LAYER M2 ;
        RECT 6.364 18.92 8.836 18.952 ;
  LAYER M2 ;
        RECT 6.364 18.984 8.836 19.016 ;
  LAYER M2 ;
        RECT 6.364 19.048 8.836 19.08 ;
  LAYER M2 ;
        RECT 6.364 19.112 8.836 19.144 ;
  LAYER M2 ;
        RECT 6.364 19.176 8.836 19.208 ;
  LAYER M2 ;
        RECT 6.364 19.24 8.836 19.272 ;
  LAYER M2 ;
        RECT 6.364 19.304 8.836 19.336 ;
  LAYER M2 ;
        RECT 6.364 19.368 8.836 19.4 ;
  LAYER M2 ;
        RECT 6.364 19.432 8.836 19.464 ;
  LAYER M2 ;
        RECT 6.364 19.496 8.836 19.528 ;
  LAYER M2 ;
        RECT 6.364 19.56 8.836 19.592 ;
  LAYER M2 ;
        RECT 6.364 19.624 8.836 19.656 ;
  LAYER M2 ;
        RECT 6.364 19.688 8.836 19.72 ;
  LAYER M2 ;
        RECT 6.364 19.752 8.836 19.784 ;
  LAYER M2 ;
        RECT 6.364 19.816 8.836 19.848 ;
  LAYER M2 ;
        RECT 6.364 19.88 8.836 19.912 ;
  LAYER M2 ;
        RECT 6.364 19.944 8.836 19.976 ;
  LAYER M2 ;
        RECT 6.364 20.008 8.836 20.04 ;
  LAYER M2 ;
        RECT 6.364 20.072 8.836 20.104 ;
  LAYER M2 ;
        RECT 6.364 20.136 8.836 20.168 ;
  LAYER M2 ;
        RECT 6.364 20.2 8.836 20.232 ;
  LAYER M2 ;
        RECT 6.364 20.264 8.836 20.296 ;
  LAYER M3 ;
        RECT 6.384 17.94 6.416 20.448 ;
  LAYER M3 ;
        RECT 6.448 17.94 6.48 20.448 ;
  LAYER M3 ;
        RECT 6.512 17.94 6.544 20.448 ;
  LAYER M3 ;
        RECT 6.576 17.94 6.608 20.448 ;
  LAYER M3 ;
        RECT 6.64 17.94 6.672 20.448 ;
  LAYER M3 ;
        RECT 6.704 17.94 6.736 20.448 ;
  LAYER M3 ;
        RECT 6.768 17.94 6.8 20.448 ;
  LAYER M3 ;
        RECT 6.832 17.94 6.864 20.448 ;
  LAYER M3 ;
        RECT 6.896 17.94 6.928 20.448 ;
  LAYER M3 ;
        RECT 6.96 17.94 6.992 20.448 ;
  LAYER M3 ;
        RECT 7.024 17.94 7.056 20.448 ;
  LAYER M3 ;
        RECT 7.088 17.94 7.12 20.448 ;
  LAYER M3 ;
        RECT 7.152 17.94 7.184 20.448 ;
  LAYER M3 ;
        RECT 7.216 17.94 7.248 20.448 ;
  LAYER M3 ;
        RECT 7.28 17.94 7.312 20.448 ;
  LAYER M3 ;
        RECT 7.344 17.94 7.376 20.448 ;
  LAYER M3 ;
        RECT 7.408 17.94 7.44 20.448 ;
  LAYER M3 ;
        RECT 7.472 17.94 7.504 20.448 ;
  LAYER M3 ;
        RECT 7.536 17.94 7.568 20.448 ;
  LAYER M3 ;
        RECT 7.6 17.94 7.632 20.448 ;
  LAYER M3 ;
        RECT 7.664 17.94 7.696 20.448 ;
  LAYER M3 ;
        RECT 7.728 17.94 7.76 20.448 ;
  LAYER M3 ;
        RECT 7.792 17.94 7.824 20.448 ;
  LAYER M3 ;
        RECT 7.856 17.94 7.888 20.448 ;
  LAYER M3 ;
        RECT 7.92 17.94 7.952 20.448 ;
  LAYER M3 ;
        RECT 7.984 17.94 8.016 20.448 ;
  LAYER M3 ;
        RECT 8.048 17.94 8.08 20.448 ;
  LAYER M3 ;
        RECT 8.112 17.94 8.144 20.448 ;
  LAYER M3 ;
        RECT 8.176 17.94 8.208 20.448 ;
  LAYER M3 ;
        RECT 8.24 17.94 8.272 20.448 ;
  LAYER M3 ;
        RECT 8.304 17.94 8.336 20.448 ;
  LAYER M3 ;
        RECT 8.368 17.94 8.4 20.448 ;
  LAYER M3 ;
        RECT 8.432 17.94 8.464 20.448 ;
  LAYER M3 ;
        RECT 8.496 17.94 8.528 20.448 ;
  LAYER M3 ;
        RECT 8.56 17.94 8.592 20.448 ;
  LAYER M3 ;
        RECT 8.624 17.94 8.656 20.448 ;
  LAYER M3 ;
        RECT 8.688 17.94 8.72 20.448 ;
  LAYER M3 ;
        RECT 8.784 17.94 8.816 20.448 ;
  LAYER M1 ;
        RECT 6.399 17.976 6.401 20.412 ;
  LAYER M1 ;
        RECT 6.479 17.976 6.481 20.412 ;
  LAYER M1 ;
        RECT 6.559 17.976 6.561 20.412 ;
  LAYER M1 ;
        RECT 6.639 17.976 6.641 20.412 ;
  LAYER M1 ;
        RECT 6.719 17.976 6.721 20.412 ;
  LAYER M1 ;
        RECT 6.799 17.976 6.801 20.412 ;
  LAYER M1 ;
        RECT 6.879 17.976 6.881 20.412 ;
  LAYER M1 ;
        RECT 6.959 17.976 6.961 20.412 ;
  LAYER M1 ;
        RECT 7.039 17.976 7.041 20.412 ;
  LAYER M1 ;
        RECT 7.119 17.976 7.121 20.412 ;
  LAYER M1 ;
        RECT 7.199 17.976 7.201 20.412 ;
  LAYER M1 ;
        RECT 7.279 17.976 7.281 20.412 ;
  LAYER M1 ;
        RECT 7.359 17.976 7.361 20.412 ;
  LAYER M1 ;
        RECT 7.439 17.976 7.441 20.412 ;
  LAYER M1 ;
        RECT 7.519 17.976 7.521 20.412 ;
  LAYER M1 ;
        RECT 7.599 17.976 7.601 20.412 ;
  LAYER M1 ;
        RECT 7.679 17.976 7.681 20.412 ;
  LAYER M1 ;
        RECT 7.759 17.976 7.761 20.412 ;
  LAYER M1 ;
        RECT 7.839 17.976 7.841 20.412 ;
  LAYER M1 ;
        RECT 7.919 17.976 7.921 20.412 ;
  LAYER M1 ;
        RECT 7.999 17.976 8.001 20.412 ;
  LAYER M1 ;
        RECT 8.079 17.976 8.081 20.412 ;
  LAYER M1 ;
        RECT 8.159 17.976 8.161 20.412 ;
  LAYER M1 ;
        RECT 8.239 17.976 8.241 20.412 ;
  LAYER M1 ;
        RECT 8.319 17.976 8.321 20.412 ;
  LAYER M1 ;
        RECT 8.399 17.976 8.401 20.412 ;
  LAYER M1 ;
        RECT 8.479 17.976 8.481 20.412 ;
  LAYER M1 ;
        RECT 8.559 17.976 8.561 20.412 ;
  LAYER M1 ;
        RECT 8.639 17.976 8.641 20.412 ;
  LAYER M1 ;
        RECT 8.719 17.976 8.721 20.412 ;
  LAYER M2 ;
        RECT 6.4 17.975 8.8 17.977 ;
  LAYER M2 ;
        RECT 6.4 18.059 8.8 18.061 ;
  LAYER M2 ;
        RECT 6.4 18.143 8.8 18.145 ;
  LAYER M2 ;
        RECT 6.4 18.227 8.8 18.229 ;
  LAYER M2 ;
        RECT 6.4 18.311 8.8 18.313 ;
  LAYER M2 ;
        RECT 6.4 18.395 8.8 18.397 ;
  LAYER M2 ;
        RECT 6.4 18.479 8.8 18.481 ;
  LAYER M2 ;
        RECT 6.4 18.563 8.8 18.565 ;
  LAYER M2 ;
        RECT 6.4 18.647 8.8 18.649 ;
  LAYER M2 ;
        RECT 6.4 18.731 8.8 18.733 ;
  LAYER M2 ;
        RECT 6.4 18.815 8.8 18.817 ;
  LAYER M2 ;
        RECT 6.4 18.899 8.8 18.901 ;
  LAYER M2 ;
        RECT 6.4 18.9825 8.8 18.9845 ;
  LAYER M2 ;
        RECT 6.4 19.067 8.8 19.069 ;
  LAYER M2 ;
        RECT 6.4 19.151 8.8 19.153 ;
  LAYER M2 ;
        RECT 6.4 19.235 8.8 19.237 ;
  LAYER M2 ;
        RECT 6.4 19.319 8.8 19.321 ;
  LAYER M2 ;
        RECT 6.4 19.403 8.8 19.405 ;
  LAYER M2 ;
        RECT 6.4 19.487 8.8 19.489 ;
  LAYER M2 ;
        RECT 6.4 19.571 8.8 19.573 ;
  LAYER M2 ;
        RECT 6.4 19.655 8.8 19.657 ;
  LAYER M2 ;
        RECT 6.4 19.739 8.8 19.741 ;
  LAYER M2 ;
        RECT 6.4 19.823 8.8 19.825 ;
  LAYER M2 ;
        RECT 6.4 19.907 8.8 19.909 ;
  LAYER M2 ;
        RECT 6.4 19.991 8.8 19.993 ;
  LAYER M2 ;
        RECT 6.4 20.075 8.8 20.077 ;
  LAYER M2 ;
        RECT 6.4 20.159 8.8 20.161 ;
  LAYER M2 ;
        RECT 6.4 20.243 8.8 20.245 ;
  LAYER M2 ;
        RECT 6.4 20.327 8.8 20.329 ;
  LAYER M1 ;
        RECT 6.384 20.88 6.416 23.388 ;
  LAYER M1 ;
        RECT 6.448 20.88 6.48 23.388 ;
  LAYER M1 ;
        RECT 6.512 20.88 6.544 23.388 ;
  LAYER M1 ;
        RECT 6.576 20.88 6.608 23.388 ;
  LAYER M1 ;
        RECT 6.64 20.88 6.672 23.388 ;
  LAYER M1 ;
        RECT 6.704 20.88 6.736 23.388 ;
  LAYER M1 ;
        RECT 6.768 20.88 6.8 23.388 ;
  LAYER M1 ;
        RECT 6.832 20.88 6.864 23.388 ;
  LAYER M1 ;
        RECT 6.896 20.88 6.928 23.388 ;
  LAYER M1 ;
        RECT 6.96 20.88 6.992 23.388 ;
  LAYER M1 ;
        RECT 7.024 20.88 7.056 23.388 ;
  LAYER M1 ;
        RECT 7.088 20.88 7.12 23.388 ;
  LAYER M1 ;
        RECT 7.152 20.88 7.184 23.388 ;
  LAYER M1 ;
        RECT 7.216 20.88 7.248 23.388 ;
  LAYER M1 ;
        RECT 7.28 20.88 7.312 23.388 ;
  LAYER M1 ;
        RECT 7.344 20.88 7.376 23.388 ;
  LAYER M1 ;
        RECT 7.408 20.88 7.44 23.388 ;
  LAYER M1 ;
        RECT 7.472 20.88 7.504 23.388 ;
  LAYER M1 ;
        RECT 7.536 20.88 7.568 23.388 ;
  LAYER M1 ;
        RECT 7.6 20.88 7.632 23.388 ;
  LAYER M1 ;
        RECT 7.664 20.88 7.696 23.388 ;
  LAYER M1 ;
        RECT 7.728 20.88 7.76 23.388 ;
  LAYER M1 ;
        RECT 7.792 20.88 7.824 23.388 ;
  LAYER M1 ;
        RECT 7.856 20.88 7.888 23.388 ;
  LAYER M1 ;
        RECT 7.92 20.88 7.952 23.388 ;
  LAYER M1 ;
        RECT 7.984 20.88 8.016 23.388 ;
  LAYER M1 ;
        RECT 8.048 20.88 8.08 23.388 ;
  LAYER M1 ;
        RECT 8.112 20.88 8.144 23.388 ;
  LAYER M1 ;
        RECT 8.176 20.88 8.208 23.388 ;
  LAYER M1 ;
        RECT 8.24 20.88 8.272 23.388 ;
  LAYER M1 ;
        RECT 8.304 20.88 8.336 23.388 ;
  LAYER M1 ;
        RECT 8.368 20.88 8.4 23.388 ;
  LAYER M1 ;
        RECT 8.432 20.88 8.464 23.388 ;
  LAYER M1 ;
        RECT 8.496 20.88 8.528 23.388 ;
  LAYER M1 ;
        RECT 8.56 20.88 8.592 23.388 ;
  LAYER M1 ;
        RECT 8.624 20.88 8.656 23.388 ;
  LAYER M1 ;
        RECT 8.688 20.88 8.72 23.388 ;
  LAYER M2 ;
        RECT 6.364 20.964 8.836 20.996 ;
  LAYER M2 ;
        RECT 6.364 21.028 8.836 21.06 ;
  LAYER M2 ;
        RECT 6.364 21.092 8.836 21.124 ;
  LAYER M2 ;
        RECT 6.364 21.156 8.836 21.188 ;
  LAYER M2 ;
        RECT 6.364 21.22 8.836 21.252 ;
  LAYER M2 ;
        RECT 6.364 21.284 8.836 21.316 ;
  LAYER M2 ;
        RECT 6.364 21.348 8.836 21.38 ;
  LAYER M2 ;
        RECT 6.364 21.412 8.836 21.444 ;
  LAYER M2 ;
        RECT 6.364 21.476 8.836 21.508 ;
  LAYER M2 ;
        RECT 6.364 21.54 8.836 21.572 ;
  LAYER M2 ;
        RECT 6.364 21.604 8.836 21.636 ;
  LAYER M2 ;
        RECT 6.364 21.668 8.836 21.7 ;
  LAYER M2 ;
        RECT 6.364 21.732 8.836 21.764 ;
  LAYER M2 ;
        RECT 6.364 21.796 8.836 21.828 ;
  LAYER M2 ;
        RECT 6.364 21.86 8.836 21.892 ;
  LAYER M2 ;
        RECT 6.364 21.924 8.836 21.956 ;
  LAYER M2 ;
        RECT 6.364 21.988 8.836 22.02 ;
  LAYER M2 ;
        RECT 6.364 22.052 8.836 22.084 ;
  LAYER M2 ;
        RECT 6.364 22.116 8.836 22.148 ;
  LAYER M2 ;
        RECT 6.364 22.18 8.836 22.212 ;
  LAYER M2 ;
        RECT 6.364 22.244 8.836 22.276 ;
  LAYER M2 ;
        RECT 6.364 22.308 8.836 22.34 ;
  LAYER M2 ;
        RECT 6.364 22.372 8.836 22.404 ;
  LAYER M2 ;
        RECT 6.364 22.436 8.836 22.468 ;
  LAYER M2 ;
        RECT 6.364 22.5 8.836 22.532 ;
  LAYER M2 ;
        RECT 6.364 22.564 8.836 22.596 ;
  LAYER M2 ;
        RECT 6.364 22.628 8.836 22.66 ;
  LAYER M2 ;
        RECT 6.364 22.692 8.836 22.724 ;
  LAYER M2 ;
        RECT 6.364 22.756 8.836 22.788 ;
  LAYER M2 ;
        RECT 6.364 22.82 8.836 22.852 ;
  LAYER M2 ;
        RECT 6.364 22.884 8.836 22.916 ;
  LAYER M2 ;
        RECT 6.364 22.948 8.836 22.98 ;
  LAYER M2 ;
        RECT 6.364 23.012 8.836 23.044 ;
  LAYER M2 ;
        RECT 6.364 23.076 8.836 23.108 ;
  LAYER M2 ;
        RECT 6.364 23.14 8.836 23.172 ;
  LAYER M2 ;
        RECT 6.364 23.204 8.836 23.236 ;
  LAYER M3 ;
        RECT 6.384 20.88 6.416 23.388 ;
  LAYER M3 ;
        RECT 6.448 20.88 6.48 23.388 ;
  LAYER M3 ;
        RECT 6.512 20.88 6.544 23.388 ;
  LAYER M3 ;
        RECT 6.576 20.88 6.608 23.388 ;
  LAYER M3 ;
        RECT 6.64 20.88 6.672 23.388 ;
  LAYER M3 ;
        RECT 6.704 20.88 6.736 23.388 ;
  LAYER M3 ;
        RECT 6.768 20.88 6.8 23.388 ;
  LAYER M3 ;
        RECT 6.832 20.88 6.864 23.388 ;
  LAYER M3 ;
        RECT 6.896 20.88 6.928 23.388 ;
  LAYER M3 ;
        RECT 6.96 20.88 6.992 23.388 ;
  LAYER M3 ;
        RECT 7.024 20.88 7.056 23.388 ;
  LAYER M3 ;
        RECT 7.088 20.88 7.12 23.388 ;
  LAYER M3 ;
        RECT 7.152 20.88 7.184 23.388 ;
  LAYER M3 ;
        RECT 7.216 20.88 7.248 23.388 ;
  LAYER M3 ;
        RECT 7.28 20.88 7.312 23.388 ;
  LAYER M3 ;
        RECT 7.344 20.88 7.376 23.388 ;
  LAYER M3 ;
        RECT 7.408 20.88 7.44 23.388 ;
  LAYER M3 ;
        RECT 7.472 20.88 7.504 23.388 ;
  LAYER M3 ;
        RECT 7.536 20.88 7.568 23.388 ;
  LAYER M3 ;
        RECT 7.6 20.88 7.632 23.388 ;
  LAYER M3 ;
        RECT 7.664 20.88 7.696 23.388 ;
  LAYER M3 ;
        RECT 7.728 20.88 7.76 23.388 ;
  LAYER M3 ;
        RECT 7.792 20.88 7.824 23.388 ;
  LAYER M3 ;
        RECT 7.856 20.88 7.888 23.388 ;
  LAYER M3 ;
        RECT 7.92 20.88 7.952 23.388 ;
  LAYER M3 ;
        RECT 7.984 20.88 8.016 23.388 ;
  LAYER M3 ;
        RECT 8.048 20.88 8.08 23.388 ;
  LAYER M3 ;
        RECT 8.112 20.88 8.144 23.388 ;
  LAYER M3 ;
        RECT 8.176 20.88 8.208 23.388 ;
  LAYER M3 ;
        RECT 8.24 20.88 8.272 23.388 ;
  LAYER M3 ;
        RECT 8.304 20.88 8.336 23.388 ;
  LAYER M3 ;
        RECT 8.368 20.88 8.4 23.388 ;
  LAYER M3 ;
        RECT 8.432 20.88 8.464 23.388 ;
  LAYER M3 ;
        RECT 8.496 20.88 8.528 23.388 ;
  LAYER M3 ;
        RECT 8.56 20.88 8.592 23.388 ;
  LAYER M3 ;
        RECT 8.624 20.88 8.656 23.388 ;
  LAYER M3 ;
        RECT 8.688 20.88 8.72 23.388 ;
  LAYER M3 ;
        RECT 8.784 20.88 8.816 23.388 ;
  LAYER M1 ;
        RECT 6.399 20.916 6.401 23.352 ;
  LAYER M1 ;
        RECT 6.479 20.916 6.481 23.352 ;
  LAYER M1 ;
        RECT 6.559 20.916 6.561 23.352 ;
  LAYER M1 ;
        RECT 6.639 20.916 6.641 23.352 ;
  LAYER M1 ;
        RECT 6.719 20.916 6.721 23.352 ;
  LAYER M1 ;
        RECT 6.799 20.916 6.801 23.352 ;
  LAYER M1 ;
        RECT 6.879 20.916 6.881 23.352 ;
  LAYER M1 ;
        RECT 6.959 20.916 6.961 23.352 ;
  LAYER M1 ;
        RECT 7.039 20.916 7.041 23.352 ;
  LAYER M1 ;
        RECT 7.119 20.916 7.121 23.352 ;
  LAYER M1 ;
        RECT 7.199 20.916 7.201 23.352 ;
  LAYER M1 ;
        RECT 7.279 20.916 7.281 23.352 ;
  LAYER M1 ;
        RECT 7.359 20.916 7.361 23.352 ;
  LAYER M1 ;
        RECT 7.439 20.916 7.441 23.352 ;
  LAYER M1 ;
        RECT 7.519 20.916 7.521 23.352 ;
  LAYER M1 ;
        RECT 7.599 20.916 7.601 23.352 ;
  LAYER M1 ;
        RECT 7.679 20.916 7.681 23.352 ;
  LAYER M1 ;
        RECT 7.759 20.916 7.761 23.352 ;
  LAYER M1 ;
        RECT 7.839 20.916 7.841 23.352 ;
  LAYER M1 ;
        RECT 7.919 20.916 7.921 23.352 ;
  LAYER M1 ;
        RECT 7.999 20.916 8.001 23.352 ;
  LAYER M1 ;
        RECT 8.079 20.916 8.081 23.352 ;
  LAYER M1 ;
        RECT 8.159 20.916 8.161 23.352 ;
  LAYER M1 ;
        RECT 8.239 20.916 8.241 23.352 ;
  LAYER M1 ;
        RECT 8.319 20.916 8.321 23.352 ;
  LAYER M1 ;
        RECT 8.399 20.916 8.401 23.352 ;
  LAYER M1 ;
        RECT 8.479 20.916 8.481 23.352 ;
  LAYER M1 ;
        RECT 8.559 20.916 8.561 23.352 ;
  LAYER M1 ;
        RECT 8.639 20.916 8.641 23.352 ;
  LAYER M1 ;
        RECT 8.719 20.916 8.721 23.352 ;
  LAYER M2 ;
        RECT 6.4 20.915 8.8 20.917 ;
  LAYER M2 ;
        RECT 6.4 20.999 8.8 21.001 ;
  LAYER M2 ;
        RECT 6.4 21.083 8.8 21.085 ;
  LAYER M2 ;
        RECT 6.4 21.167 8.8 21.169 ;
  LAYER M2 ;
        RECT 6.4 21.251 8.8 21.253 ;
  LAYER M2 ;
        RECT 6.4 21.335 8.8 21.337 ;
  LAYER M2 ;
        RECT 6.4 21.419 8.8 21.421 ;
  LAYER M2 ;
        RECT 6.4 21.503 8.8 21.505 ;
  LAYER M2 ;
        RECT 6.4 21.587 8.8 21.589 ;
  LAYER M2 ;
        RECT 6.4 21.671 8.8 21.673 ;
  LAYER M2 ;
        RECT 6.4 21.755 8.8 21.757 ;
  LAYER M2 ;
        RECT 6.4 21.839 8.8 21.841 ;
  LAYER M2 ;
        RECT 6.4 21.9225 8.8 21.9245 ;
  LAYER M2 ;
        RECT 6.4 22.007 8.8 22.009 ;
  LAYER M2 ;
        RECT 6.4 22.091 8.8 22.093 ;
  LAYER M2 ;
        RECT 6.4 22.175 8.8 22.177 ;
  LAYER M2 ;
        RECT 6.4 22.259 8.8 22.261 ;
  LAYER M2 ;
        RECT 6.4 22.343 8.8 22.345 ;
  LAYER M2 ;
        RECT 6.4 22.427 8.8 22.429 ;
  LAYER M2 ;
        RECT 6.4 22.511 8.8 22.513 ;
  LAYER M2 ;
        RECT 6.4 22.595 8.8 22.597 ;
  LAYER M2 ;
        RECT 6.4 22.679 8.8 22.681 ;
  LAYER M2 ;
        RECT 6.4 22.763 8.8 22.765 ;
  LAYER M2 ;
        RECT 6.4 22.847 8.8 22.849 ;
  LAYER M2 ;
        RECT 6.4 22.931 8.8 22.933 ;
  LAYER M2 ;
        RECT 6.4 23.015 8.8 23.017 ;
  LAYER M2 ;
        RECT 6.4 23.099 8.8 23.101 ;
  LAYER M2 ;
        RECT 6.4 23.183 8.8 23.185 ;
  LAYER M2 ;
        RECT 6.4 23.267 8.8 23.269 ;
  LAYER M1 ;
        RECT 6.384 23.82 6.416 26.328 ;
  LAYER M1 ;
        RECT 6.448 23.82 6.48 26.328 ;
  LAYER M1 ;
        RECT 6.512 23.82 6.544 26.328 ;
  LAYER M1 ;
        RECT 6.576 23.82 6.608 26.328 ;
  LAYER M1 ;
        RECT 6.64 23.82 6.672 26.328 ;
  LAYER M1 ;
        RECT 6.704 23.82 6.736 26.328 ;
  LAYER M1 ;
        RECT 6.768 23.82 6.8 26.328 ;
  LAYER M1 ;
        RECT 6.832 23.82 6.864 26.328 ;
  LAYER M1 ;
        RECT 6.896 23.82 6.928 26.328 ;
  LAYER M1 ;
        RECT 6.96 23.82 6.992 26.328 ;
  LAYER M1 ;
        RECT 7.024 23.82 7.056 26.328 ;
  LAYER M1 ;
        RECT 7.088 23.82 7.12 26.328 ;
  LAYER M1 ;
        RECT 7.152 23.82 7.184 26.328 ;
  LAYER M1 ;
        RECT 7.216 23.82 7.248 26.328 ;
  LAYER M1 ;
        RECT 7.28 23.82 7.312 26.328 ;
  LAYER M1 ;
        RECT 7.344 23.82 7.376 26.328 ;
  LAYER M1 ;
        RECT 7.408 23.82 7.44 26.328 ;
  LAYER M1 ;
        RECT 7.472 23.82 7.504 26.328 ;
  LAYER M1 ;
        RECT 7.536 23.82 7.568 26.328 ;
  LAYER M1 ;
        RECT 7.6 23.82 7.632 26.328 ;
  LAYER M1 ;
        RECT 7.664 23.82 7.696 26.328 ;
  LAYER M1 ;
        RECT 7.728 23.82 7.76 26.328 ;
  LAYER M1 ;
        RECT 7.792 23.82 7.824 26.328 ;
  LAYER M1 ;
        RECT 7.856 23.82 7.888 26.328 ;
  LAYER M1 ;
        RECT 7.92 23.82 7.952 26.328 ;
  LAYER M1 ;
        RECT 7.984 23.82 8.016 26.328 ;
  LAYER M1 ;
        RECT 8.048 23.82 8.08 26.328 ;
  LAYER M1 ;
        RECT 8.112 23.82 8.144 26.328 ;
  LAYER M1 ;
        RECT 8.176 23.82 8.208 26.328 ;
  LAYER M1 ;
        RECT 8.24 23.82 8.272 26.328 ;
  LAYER M1 ;
        RECT 8.304 23.82 8.336 26.328 ;
  LAYER M1 ;
        RECT 8.368 23.82 8.4 26.328 ;
  LAYER M1 ;
        RECT 8.432 23.82 8.464 26.328 ;
  LAYER M1 ;
        RECT 8.496 23.82 8.528 26.328 ;
  LAYER M1 ;
        RECT 8.56 23.82 8.592 26.328 ;
  LAYER M1 ;
        RECT 8.624 23.82 8.656 26.328 ;
  LAYER M1 ;
        RECT 8.688 23.82 8.72 26.328 ;
  LAYER M2 ;
        RECT 6.364 23.904 8.836 23.936 ;
  LAYER M2 ;
        RECT 6.364 23.968 8.836 24 ;
  LAYER M2 ;
        RECT 6.364 24.032 8.836 24.064 ;
  LAYER M2 ;
        RECT 6.364 24.096 8.836 24.128 ;
  LAYER M2 ;
        RECT 6.364 24.16 8.836 24.192 ;
  LAYER M2 ;
        RECT 6.364 24.224 8.836 24.256 ;
  LAYER M2 ;
        RECT 6.364 24.288 8.836 24.32 ;
  LAYER M2 ;
        RECT 6.364 24.352 8.836 24.384 ;
  LAYER M2 ;
        RECT 6.364 24.416 8.836 24.448 ;
  LAYER M2 ;
        RECT 6.364 24.48 8.836 24.512 ;
  LAYER M2 ;
        RECT 6.364 24.544 8.836 24.576 ;
  LAYER M2 ;
        RECT 6.364 24.608 8.836 24.64 ;
  LAYER M2 ;
        RECT 6.364 24.672 8.836 24.704 ;
  LAYER M2 ;
        RECT 6.364 24.736 8.836 24.768 ;
  LAYER M2 ;
        RECT 6.364 24.8 8.836 24.832 ;
  LAYER M2 ;
        RECT 6.364 24.864 8.836 24.896 ;
  LAYER M2 ;
        RECT 6.364 24.928 8.836 24.96 ;
  LAYER M2 ;
        RECT 6.364 24.992 8.836 25.024 ;
  LAYER M2 ;
        RECT 6.364 25.056 8.836 25.088 ;
  LAYER M2 ;
        RECT 6.364 25.12 8.836 25.152 ;
  LAYER M2 ;
        RECT 6.364 25.184 8.836 25.216 ;
  LAYER M2 ;
        RECT 6.364 25.248 8.836 25.28 ;
  LAYER M2 ;
        RECT 6.364 25.312 8.836 25.344 ;
  LAYER M2 ;
        RECT 6.364 25.376 8.836 25.408 ;
  LAYER M2 ;
        RECT 6.364 25.44 8.836 25.472 ;
  LAYER M2 ;
        RECT 6.364 25.504 8.836 25.536 ;
  LAYER M2 ;
        RECT 6.364 25.568 8.836 25.6 ;
  LAYER M2 ;
        RECT 6.364 25.632 8.836 25.664 ;
  LAYER M2 ;
        RECT 6.364 25.696 8.836 25.728 ;
  LAYER M2 ;
        RECT 6.364 25.76 8.836 25.792 ;
  LAYER M2 ;
        RECT 6.364 25.824 8.836 25.856 ;
  LAYER M2 ;
        RECT 6.364 25.888 8.836 25.92 ;
  LAYER M2 ;
        RECT 6.364 25.952 8.836 25.984 ;
  LAYER M2 ;
        RECT 6.364 26.016 8.836 26.048 ;
  LAYER M2 ;
        RECT 6.364 26.08 8.836 26.112 ;
  LAYER M2 ;
        RECT 6.364 26.144 8.836 26.176 ;
  LAYER M3 ;
        RECT 6.384 23.82 6.416 26.328 ;
  LAYER M3 ;
        RECT 6.448 23.82 6.48 26.328 ;
  LAYER M3 ;
        RECT 6.512 23.82 6.544 26.328 ;
  LAYER M3 ;
        RECT 6.576 23.82 6.608 26.328 ;
  LAYER M3 ;
        RECT 6.64 23.82 6.672 26.328 ;
  LAYER M3 ;
        RECT 6.704 23.82 6.736 26.328 ;
  LAYER M3 ;
        RECT 6.768 23.82 6.8 26.328 ;
  LAYER M3 ;
        RECT 6.832 23.82 6.864 26.328 ;
  LAYER M3 ;
        RECT 6.896 23.82 6.928 26.328 ;
  LAYER M3 ;
        RECT 6.96 23.82 6.992 26.328 ;
  LAYER M3 ;
        RECT 7.024 23.82 7.056 26.328 ;
  LAYER M3 ;
        RECT 7.088 23.82 7.12 26.328 ;
  LAYER M3 ;
        RECT 7.152 23.82 7.184 26.328 ;
  LAYER M3 ;
        RECT 7.216 23.82 7.248 26.328 ;
  LAYER M3 ;
        RECT 7.28 23.82 7.312 26.328 ;
  LAYER M3 ;
        RECT 7.344 23.82 7.376 26.328 ;
  LAYER M3 ;
        RECT 7.408 23.82 7.44 26.328 ;
  LAYER M3 ;
        RECT 7.472 23.82 7.504 26.328 ;
  LAYER M3 ;
        RECT 7.536 23.82 7.568 26.328 ;
  LAYER M3 ;
        RECT 7.6 23.82 7.632 26.328 ;
  LAYER M3 ;
        RECT 7.664 23.82 7.696 26.328 ;
  LAYER M3 ;
        RECT 7.728 23.82 7.76 26.328 ;
  LAYER M3 ;
        RECT 7.792 23.82 7.824 26.328 ;
  LAYER M3 ;
        RECT 7.856 23.82 7.888 26.328 ;
  LAYER M3 ;
        RECT 7.92 23.82 7.952 26.328 ;
  LAYER M3 ;
        RECT 7.984 23.82 8.016 26.328 ;
  LAYER M3 ;
        RECT 8.048 23.82 8.08 26.328 ;
  LAYER M3 ;
        RECT 8.112 23.82 8.144 26.328 ;
  LAYER M3 ;
        RECT 8.176 23.82 8.208 26.328 ;
  LAYER M3 ;
        RECT 8.24 23.82 8.272 26.328 ;
  LAYER M3 ;
        RECT 8.304 23.82 8.336 26.328 ;
  LAYER M3 ;
        RECT 8.368 23.82 8.4 26.328 ;
  LAYER M3 ;
        RECT 8.432 23.82 8.464 26.328 ;
  LAYER M3 ;
        RECT 8.496 23.82 8.528 26.328 ;
  LAYER M3 ;
        RECT 8.56 23.82 8.592 26.328 ;
  LAYER M3 ;
        RECT 8.624 23.82 8.656 26.328 ;
  LAYER M3 ;
        RECT 8.688 23.82 8.72 26.328 ;
  LAYER M3 ;
        RECT 8.784 23.82 8.816 26.328 ;
  LAYER M1 ;
        RECT 6.399 23.856 6.401 26.292 ;
  LAYER M1 ;
        RECT 6.479 23.856 6.481 26.292 ;
  LAYER M1 ;
        RECT 6.559 23.856 6.561 26.292 ;
  LAYER M1 ;
        RECT 6.639 23.856 6.641 26.292 ;
  LAYER M1 ;
        RECT 6.719 23.856 6.721 26.292 ;
  LAYER M1 ;
        RECT 6.799 23.856 6.801 26.292 ;
  LAYER M1 ;
        RECT 6.879 23.856 6.881 26.292 ;
  LAYER M1 ;
        RECT 6.959 23.856 6.961 26.292 ;
  LAYER M1 ;
        RECT 7.039 23.856 7.041 26.292 ;
  LAYER M1 ;
        RECT 7.119 23.856 7.121 26.292 ;
  LAYER M1 ;
        RECT 7.199 23.856 7.201 26.292 ;
  LAYER M1 ;
        RECT 7.279 23.856 7.281 26.292 ;
  LAYER M1 ;
        RECT 7.359 23.856 7.361 26.292 ;
  LAYER M1 ;
        RECT 7.439 23.856 7.441 26.292 ;
  LAYER M1 ;
        RECT 7.519 23.856 7.521 26.292 ;
  LAYER M1 ;
        RECT 7.599 23.856 7.601 26.292 ;
  LAYER M1 ;
        RECT 7.679 23.856 7.681 26.292 ;
  LAYER M1 ;
        RECT 7.759 23.856 7.761 26.292 ;
  LAYER M1 ;
        RECT 7.839 23.856 7.841 26.292 ;
  LAYER M1 ;
        RECT 7.919 23.856 7.921 26.292 ;
  LAYER M1 ;
        RECT 7.999 23.856 8.001 26.292 ;
  LAYER M1 ;
        RECT 8.079 23.856 8.081 26.292 ;
  LAYER M1 ;
        RECT 8.159 23.856 8.161 26.292 ;
  LAYER M1 ;
        RECT 8.239 23.856 8.241 26.292 ;
  LAYER M1 ;
        RECT 8.319 23.856 8.321 26.292 ;
  LAYER M1 ;
        RECT 8.399 23.856 8.401 26.292 ;
  LAYER M1 ;
        RECT 8.479 23.856 8.481 26.292 ;
  LAYER M1 ;
        RECT 8.559 23.856 8.561 26.292 ;
  LAYER M1 ;
        RECT 8.639 23.856 8.641 26.292 ;
  LAYER M1 ;
        RECT 8.719 23.856 8.721 26.292 ;
  LAYER M2 ;
        RECT 6.4 23.855 8.8 23.857 ;
  LAYER M2 ;
        RECT 6.4 23.939 8.8 23.941 ;
  LAYER M2 ;
        RECT 6.4 24.023 8.8 24.025 ;
  LAYER M2 ;
        RECT 6.4 24.107 8.8 24.109 ;
  LAYER M2 ;
        RECT 6.4 24.191 8.8 24.193 ;
  LAYER M2 ;
        RECT 6.4 24.275 8.8 24.277 ;
  LAYER M2 ;
        RECT 6.4 24.359 8.8 24.361 ;
  LAYER M2 ;
        RECT 6.4 24.443 8.8 24.445 ;
  LAYER M2 ;
        RECT 6.4 24.527 8.8 24.529 ;
  LAYER M2 ;
        RECT 6.4 24.611 8.8 24.613 ;
  LAYER M2 ;
        RECT 6.4 24.695 8.8 24.697 ;
  LAYER M2 ;
        RECT 6.4 24.779 8.8 24.781 ;
  LAYER M2 ;
        RECT 6.4 24.8625 8.8 24.8645 ;
  LAYER M2 ;
        RECT 6.4 24.947 8.8 24.949 ;
  LAYER M2 ;
        RECT 6.4 25.031 8.8 25.033 ;
  LAYER M2 ;
        RECT 6.4 25.115 8.8 25.117 ;
  LAYER M2 ;
        RECT 6.4 25.199 8.8 25.201 ;
  LAYER M2 ;
        RECT 6.4 25.283 8.8 25.285 ;
  LAYER M2 ;
        RECT 6.4 25.367 8.8 25.369 ;
  LAYER M2 ;
        RECT 6.4 25.451 8.8 25.453 ;
  LAYER M2 ;
        RECT 6.4 25.535 8.8 25.537 ;
  LAYER M2 ;
        RECT 6.4 25.619 8.8 25.621 ;
  LAYER M2 ;
        RECT 6.4 25.703 8.8 25.705 ;
  LAYER M2 ;
        RECT 6.4 25.787 8.8 25.789 ;
  LAYER M2 ;
        RECT 6.4 25.871 8.8 25.873 ;
  LAYER M2 ;
        RECT 6.4 25.955 8.8 25.957 ;
  LAYER M2 ;
        RECT 6.4 26.039 8.8 26.041 ;
  LAYER M2 ;
        RECT 6.4 26.123 8.8 26.125 ;
  LAYER M2 ;
        RECT 6.4 26.207 8.8 26.209 ;
  LAYER M1 ;
        RECT 6.384 26.76 6.416 29.268 ;
  LAYER M1 ;
        RECT 6.448 26.76 6.48 29.268 ;
  LAYER M1 ;
        RECT 6.512 26.76 6.544 29.268 ;
  LAYER M1 ;
        RECT 6.576 26.76 6.608 29.268 ;
  LAYER M1 ;
        RECT 6.64 26.76 6.672 29.268 ;
  LAYER M1 ;
        RECT 6.704 26.76 6.736 29.268 ;
  LAYER M1 ;
        RECT 6.768 26.76 6.8 29.268 ;
  LAYER M1 ;
        RECT 6.832 26.76 6.864 29.268 ;
  LAYER M1 ;
        RECT 6.896 26.76 6.928 29.268 ;
  LAYER M1 ;
        RECT 6.96 26.76 6.992 29.268 ;
  LAYER M1 ;
        RECT 7.024 26.76 7.056 29.268 ;
  LAYER M1 ;
        RECT 7.088 26.76 7.12 29.268 ;
  LAYER M1 ;
        RECT 7.152 26.76 7.184 29.268 ;
  LAYER M1 ;
        RECT 7.216 26.76 7.248 29.268 ;
  LAYER M1 ;
        RECT 7.28 26.76 7.312 29.268 ;
  LAYER M1 ;
        RECT 7.344 26.76 7.376 29.268 ;
  LAYER M1 ;
        RECT 7.408 26.76 7.44 29.268 ;
  LAYER M1 ;
        RECT 7.472 26.76 7.504 29.268 ;
  LAYER M1 ;
        RECT 7.536 26.76 7.568 29.268 ;
  LAYER M1 ;
        RECT 7.6 26.76 7.632 29.268 ;
  LAYER M1 ;
        RECT 7.664 26.76 7.696 29.268 ;
  LAYER M1 ;
        RECT 7.728 26.76 7.76 29.268 ;
  LAYER M1 ;
        RECT 7.792 26.76 7.824 29.268 ;
  LAYER M1 ;
        RECT 7.856 26.76 7.888 29.268 ;
  LAYER M1 ;
        RECT 7.92 26.76 7.952 29.268 ;
  LAYER M1 ;
        RECT 7.984 26.76 8.016 29.268 ;
  LAYER M1 ;
        RECT 8.048 26.76 8.08 29.268 ;
  LAYER M1 ;
        RECT 8.112 26.76 8.144 29.268 ;
  LAYER M1 ;
        RECT 8.176 26.76 8.208 29.268 ;
  LAYER M1 ;
        RECT 8.24 26.76 8.272 29.268 ;
  LAYER M1 ;
        RECT 8.304 26.76 8.336 29.268 ;
  LAYER M1 ;
        RECT 8.368 26.76 8.4 29.268 ;
  LAYER M1 ;
        RECT 8.432 26.76 8.464 29.268 ;
  LAYER M1 ;
        RECT 8.496 26.76 8.528 29.268 ;
  LAYER M1 ;
        RECT 8.56 26.76 8.592 29.268 ;
  LAYER M1 ;
        RECT 8.624 26.76 8.656 29.268 ;
  LAYER M1 ;
        RECT 8.688 26.76 8.72 29.268 ;
  LAYER M2 ;
        RECT 6.364 26.844 8.836 26.876 ;
  LAYER M2 ;
        RECT 6.364 26.908 8.836 26.94 ;
  LAYER M2 ;
        RECT 6.364 26.972 8.836 27.004 ;
  LAYER M2 ;
        RECT 6.364 27.036 8.836 27.068 ;
  LAYER M2 ;
        RECT 6.364 27.1 8.836 27.132 ;
  LAYER M2 ;
        RECT 6.364 27.164 8.836 27.196 ;
  LAYER M2 ;
        RECT 6.364 27.228 8.836 27.26 ;
  LAYER M2 ;
        RECT 6.364 27.292 8.836 27.324 ;
  LAYER M2 ;
        RECT 6.364 27.356 8.836 27.388 ;
  LAYER M2 ;
        RECT 6.364 27.42 8.836 27.452 ;
  LAYER M2 ;
        RECT 6.364 27.484 8.836 27.516 ;
  LAYER M2 ;
        RECT 6.364 27.548 8.836 27.58 ;
  LAYER M2 ;
        RECT 6.364 27.612 8.836 27.644 ;
  LAYER M2 ;
        RECT 6.364 27.676 8.836 27.708 ;
  LAYER M2 ;
        RECT 6.364 27.74 8.836 27.772 ;
  LAYER M2 ;
        RECT 6.364 27.804 8.836 27.836 ;
  LAYER M2 ;
        RECT 6.364 27.868 8.836 27.9 ;
  LAYER M2 ;
        RECT 6.364 27.932 8.836 27.964 ;
  LAYER M2 ;
        RECT 6.364 27.996 8.836 28.028 ;
  LAYER M2 ;
        RECT 6.364 28.06 8.836 28.092 ;
  LAYER M2 ;
        RECT 6.364 28.124 8.836 28.156 ;
  LAYER M2 ;
        RECT 6.364 28.188 8.836 28.22 ;
  LAYER M2 ;
        RECT 6.364 28.252 8.836 28.284 ;
  LAYER M2 ;
        RECT 6.364 28.316 8.836 28.348 ;
  LAYER M2 ;
        RECT 6.364 28.38 8.836 28.412 ;
  LAYER M2 ;
        RECT 6.364 28.444 8.836 28.476 ;
  LAYER M2 ;
        RECT 6.364 28.508 8.836 28.54 ;
  LAYER M2 ;
        RECT 6.364 28.572 8.836 28.604 ;
  LAYER M2 ;
        RECT 6.364 28.636 8.836 28.668 ;
  LAYER M2 ;
        RECT 6.364 28.7 8.836 28.732 ;
  LAYER M2 ;
        RECT 6.364 28.764 8.836 28.796 ;
  LAYER M2 ;
        RECT 6.364 28.828 8.836 28.86 ;
  LAYER M2 ;
        RECT 6.364 28.892 8.836 28.924 ;
  LAYER M2 ;
        RECT 6.364 28.956 8.836 28.988 ;
  LAYER M2 ;
        RECT 6.364 29.02 8.836 29.052 ;
  LAYER M2 ;
        RECT 6.364 29.084 8.836 29.116 ;
  LAYER M3 ;
        RECT 6.384 26.76 6.416 29.268 ;
  LAYER M3 ;
        RECT 6.448 26.76 6.48 29.268 ;
  LAYER M3 ;
        RECT 6.512 26.76 6.544 29.268 ;
  LAYER M3 ;
        RECT 6.576 26.76 6.608 29.268 ;
  LAYER M3 ;
        RECT 6.64 26.76 6.672 29.268 ;
  LAYER M3 ;
        RECT 6.704 26.76 6.736 29.268 ;
  LAYER M3 ;
        RECT 6.768 26.76 6.8 29.268 ;
  LAYER M3 ;
        RECT 6.832 26.76 6.864 29.268 ;
  LAYER M3 ;
        RECT 6.896 26.76 6.928 29.268 ;
  LAYER M3 ;
        RECT 6.96 26.76 6.992 29.268 ;
  LAYER M3 ;
        RECT 7.024 26.76 7.056 29.268 ;
  LAYER M3 ;
        RECT 7.088 26.76 7.12 29.268 ;
  LAYER M3 ;
        RECT 7.152 26.76 7.184 29.268 ;
  LAYER M3 ;
        RECT 7.216 26.76 7.248 29.268 ;
  LAYER M3 ;
        RECT 7.28 26.76 7.312 29.268 ;
  LAYER M3 ;
        RECT 7.344 26.76 7.376 29.268 ;
  LAYER M3 ;
        RECT 7.408 26.76 7.44 29.268 ;
  LAYER M3 ;
        RECT 7.472 26.76 7.504 29.268 ;
  LAYER M3 ;
        RECT 7.536 26.76 7.568 29.268 ;
  LAYER M3 ;
        RECT 7.6 26.76 7.632 29.268 ;
  LAYER M3 ;
        RECT 7.664 26.76 7.696 29.268 ;
  LAYER M3 ;
        RECT 7.728 26.76 7.76 29.268 ;
  LAYER M3 ;
        RECT 7.792 26.76 7.824 29.268 ;
  LAYER M3 ;
        RECT 7.856 26.76 7.888 29.268 ;
  LAYER M3 ;
        RECT 7.92 26.76 7.952 29.268 ;
  LAYER M3 ;
        RECT 7.984 26.76 8.016 29.268 ;
  LAYER M3 ;
        RECT 8.048 26.76 8.08 29.268 ;
  LAYER M3 ;
        RECT 8.112 26.76 8.144 29.268 ;
  LAYER M3 ;
        RECT 8.176 26.76 8.208 29.268 ;
  LAYER M3 ;
        RECT 8.24 26.76 8.272 29.268 ;
  LAYER M3 ;
        RECT 8.304 26.76 8.336 29.268 ;
  LAYER M3 ;
        RECT 8.368 26.76 8.4 29.268 ;
  LAYER M3 ;
        RECT 8.432 26.76 8.464 29.268 ;
  LAYER M3 ;
        RECT 8.496 26.76 8.528 29.268 ;
  LAYER M3 ;
        RECT 8.56 26.76 8.592 29.268 ;
  LAYER M3 ;
        RECT 8.624 26.76 8.656 29.268 ;
  LAYER M3 ;
        RECT 8.688 26.76 8.72 29.268 ;
  LAYER M3 ;
        RECT 8.784 26.76 8.816 29.268 ;
  LAYER M1 ;
        RECT 6.399 26.796 6.401 29.232 ;
  LAYER M1 ;
        RECT 6.479 26.796 6.481 29.232 ;
  LAYER M1 ;
        RECT 6.559 26.796 6.561 29.232 ;
  LAYER M1 ;
        RECT 6.639 26.796 6.641 29.232 ;
  LAYER M1 ;
        RECT 6.719 26.796 6.721 29.232 ;
  LAYER M1 ;
        RECT 6.799 26.796 6.801 29.232 ;
  LAYER M1 ;
        RECT 6.879 26.796 6.881 29.232 ;
  LAYER M1 ;
        RECT 6.959 26.796 6.961 29.232 ;
  LAYER M1 ;
        RECT 7.039 26.796 7.041 29.232 ;
  LAYER M1 ;
        RECT 7.119 26.796 7.121 29.232 ;
  LAYER M1 ;
        RECT 7.199 26.796 7.201 29.232 ;
  LAYER M1 ;
        RECT 7.279 26.796 7.281 29.232 ;
  LAYER M1 ;
        RECT 7.359 26.796 7.361 29.232 ;
  LAYER M1 ;
        RECT 7.439 26.796 7.441 29.232 ;
  LAYER M1 ;
        RECT 7.519 26.796 7.521 29.232 ;
  LAYER M1 ;
        RECT 7.599 26.796 7.601 29.232 ;
  LAYER M1 ;
        RECT 7.679 26.796 7.681 29.232 ;
  LAYER M1 ;
        RECT 7.759 26.796 7.761 29.232 ;
  LAYER M1 ;
        RECT 7.839 26.796 7.841 29.232 ;
  LAYER M1 ;
        RECT 7.919 26.796 7.921 29.232 ;
  LAYER M1 ;
        RECT 7.999 26.796 8.001 29.232 ;
  LAYER M1 ;
        RECT 8.079 26.796 8.081 29.232 ;
  LAYER M1 ;
        RECT 8.159 26.796 8.161 29.232 ;
  LAYER M1 ;
        RECT 8.239 26.796 8.241 29.232 ;
  LAYER M1 ;
        RECT 8.319 26.796 8.321 29.232 ;
  LAYER M1 ;
        RECT 8.399 26.796 8.401 29.232 ;
  LAYER M1 ;
        RECT 8.479 26.796 8.481 29.232 ;
  LAYER M1 ;
        RECT 8.559 26.796 8.561 29.232 ;
  LAYER M1 ;
        RECT 8.639 26.796 8.641 29.232 ;
  LAYER M1 ;
        RECT 8.719 26.796 8.721 29.232 ;
  LAYER M2 ;
        RECT 6.4 26.795 8.8 26.797 ;
  LAYER M2 ;
        RECT 6.4 26.879 8.8 26.881 ;
  LAYER M2 ;
        RECT 6.4 26.963 8.8 26.965 ;
  LAYER M2 ;
        RECT 6.4 27.047 8.8 27.049 ;
  LAYER M2 ;
        RECT 6.4 27.131 8.8 27.133 ;
  LAYER M2 ;
        RECT 6.4 27.215 8.8 27.217 ;
  LAYER M2 ;
        RECT 6.4 27.299 8.8 27.301 ;
  LAYER M2 ;
        RECT 6.4 27.383 8.8 27.385 ;
  LAYER M2 ;
        RECT 6.4 27.467 8.8 27.469 ;
  LAYER M2 ;
        RECT 6.4 27.551 8.8 27.553 ;
  LAYER M2 ;
        RECT 6.4 27.635 8.8 27.637 ;
  LAYER M2 ;
        RECT 6.4 27.719 8.8 27.721 ;
  LAYER M2 ;
        RECT 6.4 27.8025 8.8 27.8045 ;
  LAYER M2 ;
        RECT 6.4 27.887 8.8 27.889 ;
  LAYER M2 ;
        RECT 6.4 27.971 8.8 27.973 ;
  LAYER M2 ;
        RECT 6.4 28.055 8.8 28.057 ;
  LAYER M2 ;
        RECT 6.4 28.139 8.8 28.141 ;
  LAYER M2 ;
        RECT 6.4 28.223 8.8 28.225 ;
  LAYER M2 ;
        RECT 6.4 28.307 8.8 28.309 ;
  LAYER M2 ;
        RECT 6.4 28.391 8.8 28.393 ;
  LAYER M2 ;
        RECT 6.4 28.475 8.8 28.477 ;
  LAYER M2 ;
        RECT 6.4 28.559 8.8 28.561 ;
  LAYER M2 ;
        RECT 6.4 28.643 8.8 28.645 ;
  LAYER M2 ;
        RECT 6.4 28.727 8.8 28.729 ;
  LAYER M2 ;
        RECT 6.4 28.811 8.8 28.813 ;
  LAYER M2 ;
        RECT 6.4 28.895 8.8 28.897 ;
  LAYER M2 ;
        RECT 6.4 28.979 8.8 28.981 ;
  LAYER M2 ;
        RECT 6.4 29.063 8.8 29.065 ;
  LAYER M2 ;
        RECT 6.4 29.147 8.8 29.149 ;
  LAYER M1 ;
        RECT 9.264 17.94 9.296 20.448 ;
  LAYER M1 ;
        RECT 9.328 17.94 9.36 20.448 ;
  LAYER M1 ;
        RECT 9.392 17.94 9.424 20.448 ;
  LAYER M1 ;
        RECT 9.456 17.94 9.488 20.448 ;
  LAYER M1 ;
        RECT 9.52 17.94 9.552 20.448 ;
  LAYER M1 ;
        RECT 9.584 17.94 9.616 20.448 ;
  LAYER M1 ;
        RECT 9.648 17.94 9.68 20.448 ;
  LAYER M1 ;
        RECT 9.712 17.94 9.744 20.448 ;
  LAYER M1 ;
        RECT 9.776 17.94 9.808 20.448 ;
  LAYER M1 ;
        RECT 9.84 17.94 9.872 20.448 ;
  LAYER M1 ;
        RECT 9.904 17.94 9.936 20.448 ;
  LAYER M1 ;
        RECT 9.968 17.94 10 20.448 ;
  LAYER M1 ;
        RECT 10.032 17.94 10.064 20.448 ;
  LAYER M1 ;
        RECT 10.096 17.94 10.128 20.448 ;
  LAYER M1 ;
        RECT 10.16 17.94 10.192 20.448 ;
  LAYER M1 ;
        RECT 10.224 17.94 10.256 20.448 ;
  LAYER M1 ;
        RECT 10.288 17.94 10.32 20.448 ;
  LAYER M1 ;
        RECT 10.352 17.94 10.384 20.448 ;
  LAYER M1 ;
        RECT 10.416 17.94 10.448 20.448 ;
  LAYER M1 ;
        RECT 10.48 17.94 10.512 20.448 ;
  LAYER M1 ;
        RECT 10.544 17.94 10.576 20.448 ;
  LAYER M1 ;
        RECT 10.608 17.94 10.64 20.448 ;
  LAYER M1 ;
        RECT 10.672 17.94 10.704 20.448 ;
  LAYER M1 ;
        RECT 10.736 17.94 10.768 20.448 ;
  LAYER M1 ;
        RECT 10.8 17.94 10.832 20.448 ;
  LAYER M1 ;
        RECT 10.864 17.94 10.896 20.448 ;
  LAYER M1 ;
        RECT 10.928 17.94 10.96 20.448 ;
  LAYER M1 ;
        RECT 10.992 17.94 11.024 20.448 ;
  LAYER M1 ;
        RECT 11.056 17.94 11.088 20.448 ;
  LAYER M1 ;
        RECT 11.12 17.94 11.152 20.448 ;
  LAYER M1 ;
        RECT 11.184 17.94 11.216 20.448 ;
  LAYER M1 ;
        RECT 11.248 17.94 11.28 20.448 ;
  LAYER M1 ;
        RECT 11.312 17.94 11.344 20.448 ;
  LAYER M1 ;
        RECT 11.376 17.94 11.408 20.448 ;
  LAYER M1 ;
        RECT 11.44 17.94 11.472 20.448 ;
  LAYER M1 ;
        RECT 11.504 17.94 11.536 20.448 ;
  LAYER M1 ;
        RECT 11.568 17.94 11.6 20.448 ;
  LAYER M2 ;
        RECT 9.244 18.024 11.716 18.056 ;
  LAYER M2 ;
        RECT 9.244 18.088 11.716 18.12 ;
  LAYER M2 ;
        RECT 9.244 18.152 11.716 18.184 ;
  LAYER M2 ;
        RECT 9.244 18.216 11.716 18.248 ;
  LAYER M2 ;
        RECT 9.244 18.28 11.716 18.312 ;
  LAYER M2 ;
        RECT 9.244 18.344 11.716 18.376 ;
  LAYER M2 ;
        RECT 9.244 18.408 11.716 18.44 ;
  LAYER M2 ;
        RECT 9.244 18.472 11.716 18.504 ;
  LAYER M2 ;
        RECT 9.244 18.536 11.716 18.568 ;
  LAYER M2 ;
        RECT 9.244 18.6 11.716 18.632 ;
  LAYER M2 ;
        RECT 9.244 18.664 11.716 18.696 ;
  LAYER M2 ;
        RECT 9.244 18.728 11.716 18.76 ;
  LAYER M2 ;
        RECT 9.244 18.792 11.716 18.824 ;
  LAYER M2 ;
        RECT 9.244 18.856 11.716 18.888 ;
  LAYER M2 ;
        RECT 9.244 18.92 11.716 18.952 ;
  LAYER M2 ;
        RECT 9.244 18.984 11.716 19.016 ;
  LAYER M2 ;
        RECT 9.244 19.048 11.716 19.08 ;
  LAYER M2 ;
        RECT 9.244 19.112 11.716 19.144 ;
  LAYER M2 ;
        RECT 9.244 19.176 11.716 19.208 ;
  LAYER M2 ;
        RECT 9.244 19.24 11.716 19.272 ;
  LAYER M2 ;
        RECT 9.244 19.304 11.716 19.336 ;
  LAYER M2 ;
        RECT 9.244 19.368 11.716 19.4 ;
  LAYER M2 ;
        RECT 9.244 19.432 11.716 19.464 ;
  LAYER M2 ;
        RECT 9.244 19.496 11.716 19.528 ;
  LAYER M2 ;
        RECT 9.244 19.56 11.716 19.592 ;
  LAYER M2 ;
        RECT 9.244 19.624 11.716 19.656 ;
  LAYER M2 ;
        RECT 9.244 19.688 11.716 19.72 ;
  LAYER M2 ;
        RECT 9.244 19.752 11.716 19.784 ;
  LAYER M2 ;
        RECT 9.244 19.816 11.716 19.848 ;
  LAYER M2 ;
        RECT 9.244 19.88 11.716 19.912 ;
  LAYER M2 ;
        RECT 9.244 19.944 11.716 19.976 ;
  LAYER M2 ;
        RECT 9.244 20.008 11.716 20.04 ;
  LAYER M2 ;
        RECT 9.244 20.072 11.716 20.104 ;
  LAYER M2 ;
        RECT 9.244 20.136 11.716 20.168 ;
  LAYER M2 ;
        RECT 9.244 20.2 11.716 20.232 ;
  LAYER M2 ;
        RECT 9.244 20.264 11.716 20.296 ;
  LAYER M3 ;
        RECT 9.264 17.94 9.296 20.448 ;
  LAYER M3 ;
        RECT 9.328 17.94 9.36 20.448 ;
  LAYER M3 ;
        RECT 9.392 17.94 9.424 20.448 ;
  LAYER M3 ;
        RECT 9.456 17.94 9.488 20.448 ;
  LAYER M3 ;
        RECT 9.52 17.94 9.552 20.448 ;
  LAYER M3 ;
        RECT 9.584 17.94 9.616 20.448 ;
  LAYER M3 ;
        RECT 9.648 17.94 9.68 20.448 ;
  LAYER M3 ;
        RECT 9.712 17.94 9.744 20.448 ;
  LAYER M3 ;
        RECT 9.776 17.94 9.808 20.448 ;
  LAYER M3 ;
        RECT 9.84 17.94 9.872 20.448 ;
  LAYER M3 ;
        RECT 9.904 17.94 9.936 20.448 ;
  LAYER M3 ;
        RECT 9.968 17.94 10 20.448 ;
  LAYER M3 ;
        RECT 10.032 17.94 10.064 20.448 ;
  LAYER M3 ;
        RECT 10.096 17.94 10.128 20.448 ;
  LAYER M3 ;
        RECT 10.16 17.94 10.192 20.448 ;
  LAYER M3 ;
        RECT 10.224 17.94 10.256 20.448 ;
  LAYER M3 ;
        RECT 10.288 17.94 10.32 20.448 ;
  LAYER M3 ;
        RECT 10.352 17.94 10.384 20.448 ;
  LAYER M3 ;
        RECT 10.416 17.94 10.448 20.448 ;
  LAYER M3 ;
        RECT 10.48 17.94 10.512 20.448 ;
  LAYER M3 ;
        RECT 10.544 17.94 10.576 20.448 ;
  LAYER M3 ;
        RECT 10.608 17.94 10.64 20.448 ;
  LAYER M3 ;
        RECT 10.672 17.94 10.704 20.448 ;
  LAYER M3 ;
        RECT 10.736 17.94 10.768 20.448 ;
  LAYER M3 ;
        RECT 10.8 17.94 10.832 20.448 ;
  LAYER M3 ;
        RECT 10.864 17.94 10.896 20.448 ;
  LAYER M3 ;
        RECT 10.928 17.94 10.96 20.448 ;
  LAYER M3 ;
        RECT 10.992 17.94 11.024 20.448 ;
  LAYER M3 ;
        RECT 11.056 17.94 11.088 20.448 ;
  LAYER M3 ;
        RECT 11.12 17.94 11.152 20.448 ;
  LAYER M3 ;
        RECT 11.184 17.94 11.216 20.448 ;
  LAYER M3 ;
        RECT 11.248 17.94 11.28 20.448 ;
  LAYER M3 ;
        RECT 11.312 17.94 11.344 20.448 ;
  LAYER M3 ;
        RECT 11.376 17.94 11.408 20.448 ;
  LAYER M3 ;
        RECT 11.44 17.94 11.472 20.448 ;
  LAYER M3 ;
        RECT 11.504 17.94 11.536 20.448 ;
  LAYER M3 ;
        RECT 11.568 17.94 11.6 20.448 ;
  LAYER M3 ;
        RECT 11.664 17.94 11.696 20.448 ;
  LAYER M1 ;
        RECT 9.279 17.976 9.281 20.412 ;
  LAYER M1 ;
        RECT 9.359 17.976 9.361 20.412 ;
  LAYER M1 ;
        RECT 9.439 17.976 9.441 20.412 ;
  LAYER M1 ;
        RECT 9.519 17.976 9.521 20.412 ;
  LAYER M1 ;
        RECT 9.599 17.976 9.601 20.412 ;
  LAYER M1 ;
        RECT 9.679 17.976 9.681 20.412 ;
  LAYER M1 ;
        RECT 9.759 17.976 9.761 20.412 ;
  LAYER M1 ;
        RECT 9.839 17.976 9.841 20.412 ;
  LAYER M1 ;
        RECT 9.919 17.976 9.921 20.412 ;
  LAYER M1 ;
        RECT 9.999 17.976 10.001 20.412 ;
  LAYER M1 ;
        RECT 10.079 17.976 10.081 20.412 ;
  LAYER M1 ;
        RECT 10.159 17.976 10.161 20.412 ;
  LAYER M1 ;
        RECT 10.239 17.976 10.241 20.412 ;
  LAYER M1 ;
        RECT 10.319 17.976 10.321 20.412 ;
  LAYER M1 ;
        RECT 10.399 17.976 10.401 20.412 ;
  LAYER M1 ;
        RECT 10.479 17.976 10.481 20.412 ;
  LAYER M1 ;
        RECT 10.559 17.976 10.561 20.412 ;
  LAYER M1 ;
        RECT 10.639 17.976 10.641 20.412 ;
  LAYER M1 ;
        RECT 10.719 17.976 10.721 20.412 ;
  LAYER M1 ;
        RECT 10.799 17.976 10.801 20.412 ;
  LAYER M1 ;
        RECT 10.879 17.976 10.881 20.412 ;
  LAYER M1 ;
        RECT 10.959 17.976 10.961 20.412 ;
  LAYER M1 ;
        RECT 11.039 17.976 11.041 20.412 ;
  LAYER M1 ;
        RECT 11.119 17.976 11.121 20.412 ;
  LAYER M1 ;
        RECT 11.199 17.976 11.201 20.412 ;
  LAYER M1 ;
        RECT 11.279 17.976 11.281 20.412 ;
  LAYER M1 ;
        RECT 11.359 17.976 11.361 20.412 ;
  LAYER M1 ;
        RECT 11.439 17.976 11.441 20.412 ;
  LAYER M1 ;
        RECT 11.519 17.976 11.521 20.412 ;
  LAYER M1 ;
        RECT 11.599 17.976 11.601 20.412 ;
  LAYER M2 ;
        RECT 9.28 17.975 11.68 17.977 ;
  LAYER M2 ;
        RECT 9.28 18.059 11.68 18.061 ;
  LAYER M2 ;
        RECT 9.28 18.143 11.68 18.145 ;
  LAYER M2 ;
        RECT 9.28 18.227 11.68 18.229 ;
  LAYER M2 ;
        RECT 9.28 18.311 11.68 18.313 ;
  LAYER M2 ;
        RECT 9.28 18.395 11.68 18.397 ;
  LAYER M2 ;
        RECT 9.28 18.479 11.68 18.481 ;
  LAYER M2 ;
        RECT 9.28 18.563 11.68 18.565 ;
  LAYER M2 ;
        RECT 9.28 18.647 11.68 18.649 ;
  LAYER M2 ;
        RECT 9.28 18.731 11.68 18.733 ;
  LAYER M2 ;
        RECT 9.28 18.815 11.68 18.817 ;
  LAYER M2 ;
        RECT 9.28 18.899 11.68 18.901 ;
  LAYER M2 ;
        RECT 9.28 18.9825 11.68 18.9845 ;
  LAYER M2 ;
        RECT 9.28 19.067 11.68 19.069 ;
  LAYER M2 ;
        RECT 9.28 19.151 11.68 19.153 ;
  LAYER M2 ;
        RECT 9.28 19.235 11.68 19.237 ;
  LAYER M2 ;
        RECT 9.28 19.319 11.68 19.321 ;
  LAYER M2 ;
        RECT 9.28 19.403 11.68 19.405 ;
  LAYER M2 ;
        RECT 9.28 19.487 11.68 19.489 ;
  LAYER M2 ;
        RECT 9.28 19.571 11.68 19.573 ;
  LAYER M2 ;
        RECT 9.28 19.655 11.68 19.657 ;
  LAYER M2 ;
        RECT 9.28 19.739 11.68 19.741 ;
  LAYER M2 ;
        RECT 9.28 19.823 11.68 19.825 ;
  LAYER M2 ;
        RECT 9.28 19.907 11.68 19.909 ;
  LAYER M2 ;
        RECT 9.28 19.991 11.68 19.993 ;
  LAYER M2 ;
        RECT 9.28 20.075 11.68 20.077 ;
  LAYER M2 ;
        RECT 9.28 20.159 11.68 20.161 ;
  LAYER M2 ;
        RECT 9.28 20.243 11.68 20.245 ;
  LAYER M2 ;
        RECT 9.28 20.327 11.68 20.329 ;
  LAYER M1 ;
        RECT 9.264 20.88 9.296 23.388 ;
  LAYER M1 ;
        RECT 9.328 20.88 9.36 23.388 ;
  LAYER M1 ;
        RECT 9.392 20.88 9.424 23.388 ;
  LAYER M1 ;
        RECT 9.456 20.88 9.488 23.388 ;
  LAYER M1 ;
        RECT 9.52 20.88 9.552 23.388 ;
  LAYER M1 ;
        RECT 9.584 20.88 9.616 23.388 ;
  LAYER M1 ;
        RECT 9.648 20.88 9.68 23.388 ;
  LAYER M1 ;
        RECT 9.712 20.88 9.744 23.388 ;
  LAYER M1 ;
        RECT 9.776 20.88 9.808 23.388 ;
  LAYER M1 ;
        RECT 9.84 20.88 9.872 23.388 ;
  LAYER M1 ;
        RECT 9.904 20.88 9.936 23.388 ;
  LAYER M1 ;
        RECT 9.968 20.88 10 23.388 ;
  LAYER M1 ;
        RECT 10.032 20.88 10.064 23.388 ;
  LAYER M1 ;
        RECT 10.096 20.88 10.128 23.388 ;
  LAYER M1 ;
        RECT 10.16 20.88 10.192 23.388 ;
  LAYER M1 ;
        RECT 10.224 20.88 10.256 23.388 ;
  LAYER M1 ;
        RECT 10.288 20.88 10.32 23.388 ;
  LAYER M1 ;
        RECT 10.352 20.88 10.384 23.388 ;
  LAYER M1 ;
        RECT 10.416 20.88 10.448 23.388 ;
  LAYER M1 ;
        RECT 10.48 20.88 10.512 23.388 ;
  LAYER M1 ;
        RECT 10.544 20.88 10.576 23.388 ;
  LAYER M1 ;
        RECT 10.608 20.88 10.64 23.388 ;
  LAYER M1 ;
        RECT 10.672 20.88 10.704 23.388 ;
  LAYER M1 ;
        RECT 10.736 20.88 10.768 23.388 ;
  LAYER M1 ;
        RECT 10.8 20.88 10.832 23.388 ;
  LAYER M1 ;
        RECT 10.864 20.88 10.896 23.388 ;
  LAYER M1 ;
        RECT 10.928 20.88 10.96 23.388 ;
  LAYER M1 ;
        RECT 10.992 20.88 11.024 23.388 ;
  LAYER M1 ;
        RECT 11.056 20.88 11.088 23.388 ;
  LAYER M1 ;
        RECT 11.12 20.88 11.152 23.388 ;
  LAYER M1 ;
        RECT 11.184 20.88 11.216 23.388 ;
  LAYER M1 ;
        RECT 11.248 20.88 11.28 23.388 ;
  LAYER M1 ;
        RECT 11.312 20.88 11.344 23.388 ;
  LAYER M1 ;
        RECT 11.376 20.88 11.408 23.388 ;
  LAYER M1 ;
        RECT 11.44 20.88 11.472 23.388 ;
  LAYER M1 ;
        RECT 11.504 20.88 11.536 23.388 ;
  LAYER M1 ;
        RECT 11.568 20.88 11.6 23.388 ;
  LAYER M2 ;
        RECT 9.244 20.964 11.716 20.996 ;
  LAYER M2 ;
        RECT 9.244 21.028 11.716 21.06 ;
  LAYER M2 ;
        RECT 9.244 21.092 11.716 21.124 ;
  LAYER M2 ;
        RECT 9.244 21.156 11.716 21.188 ;
  LAYER M2 ;
        RECT 9.244 21.22 11.716 21.252 ;
  LAYER M2 ;
        RECT 9.244 21.284 11.716 21.316 ;
  LAYER M2 ;
        RECT 9.244 21.348 11.716 21.38 ;
  LAYER M2 ;
        RECT 9.244 21.412 11.716 21.444 ;
  LAYER M2 ;
        RECT 9.244 21.476 11.716 21.508 ;
  LAYER M2 ;
        RECT 9.244 21.54 11.716 21.572 ;
  LAYER M2 ;
        RECT 9.244 21.604 11.716 21.636 ;
  LAYER M2 ;
        RECT 9.244 21.668 11.716 21.7 ;
  LAYER M2 ;
        RECT 9.244 21.732 11.716 21.764 ;
  LAYER M2 ;
        RECT 9.244 21.796 11.716 21.828 ;
  LAYER M2 ;
        RECT 9.244 21.86 11.716 21.892 ;
  LAYER M2 ;
        RECT 9.244 21.924 11.716 21.956 ;
  LAYER M2 ;
        RECT 9.244 21.988 11.716 22.02 ;
  LAYER M2 ;
        RECT 9.244 22.052 11.716 22.084 ;
  LAYER M2 ;
        RECT 9.244 22.116 11.716 22.148 ;
  LAYER M2 ;
        RECT 9.244 22.18 11.716 22.212 ;
  LAYER M2 ;
        RECT 9.244 22.244 11.716 22.276 ;
  LAYER M2 ;
        RECT 9.244 22.308 11.716 22.34 ;
  LAYER M2 ;
        RECT 9.244 22.372 11.716 22.404 ;
  LAYER M2 ;
        RECT 9.244 22.436 11.716 22.468 ;
  LAYER M2 ;
        RECT 9.244 22.5 11.716 22.532 ;
  LAYER M2 ;
        RECT 9.244 22.564 11.716 22.596 ;
  LAYER M2 ;
        RECT 9.244 22.628 11.716 22.66 ;
  LAYER M2 ;
        RECT 9.244 22.692 11.716 22.724 ;
  LAYER M2 ;
        RECT 9.244 22.756 11.716 22.788 ;
  LAYER M2 ;
        RECT 9.244 22.82 11.716 22.852 ;
  LAYER M2 ;
        RECT 9.244 22.884 11.716 22.916 ;
  LAYER M2 ;
        RECT 9.244 22.948 11.716 22.98 ;
  LAYER M2 ;
        RECT 9.244 23.012 11.716 23.044 ;
  LAYER M2 ;
        RECT 9.244 23.076 11.716 23.108 ;
  LAYER M2 ;
        RECT 9.244 23.14 11.716 23.172 ;
  LAYER M2 ;
        RECT 9.244 23.204 11.716 23.236 ;
  LAYER M3 ;
        RECT 9.264 20.88 9.296 23.388 ;
  LAYER M3 ;
        RECT 9.328 20.88 9.36 23.388 ;
  LAYER M3 ;
        RECT 9.392 20.88 9.424 23.388 ;
  LAYER M3 ;
        RECT 9.456 20.88 9.488 23.388 ;
  LAYER M3 ;
        RECT 9.52 20.88 9.552 23.388 ;
  LAYER M3 ;
        RECT 9.584 20.88 9.616 23.388 ;
  LAYER M3 ;
        RECT 9.648 20.88 9.68 23.388 ;
  LAYER M3 ;
        RECT 9.712 20.88 9.744 23.388 ;
  LAYER M3 ;
        RECT 9.776 20.88 9.808 23.388 ;
  LAYER M3 ;
        RECT 9.84 20.88 9.872 23.388 ;
  LAYER M3 ;
        RECT 9.904 20.88 9.936 23.388 ;
  LAYER M3 ;
        RECT 9.968 20.88 10 23.388 ;
  LAYER M3 ;
        RECT 10.032 20.88 10.064 23.388 ;
  LAYER M3 ;
        RECT 10.096 20.88 10.128 23.388 ;
  LAYER M3 ;
        RECT 10.16 20.88 10.192 23.388 ;
  LAYER M3 ;
        RECT 10.224 20.88 10.256 23.388 ;
  LAYER M3 ;
        RECT 10.288 20.88 10.32 23.388 ;
  LAYER M3 ;
        RECT 10.352 20.88 10.384 23.388 ;
  LAYER M3 ;
        RECT 10.416 20.88 10.448 23.388 ;
  LAYER M3 ;
        RECT 10.48 20.88 10.512 23.388 ;
  LAYER M3 ;
        RECT 10.544 20.88 10.576 23.388 ;
  LAYER M3 ;
        RECT 10.608 20.88 10.64 23.388 ;
  LAYER M3 ;
        RECT 10.672 20.88 10.704 23.388 ;
  LAYER M3 ;
        RECT 10.736 20.88 10.768 23.388 ;
  LAYER M3 ;
        RECT 10.8 20.88 10.832 23.388 ;
  LAYER M3 ;
        RECT 10.864 20.88 10.896 23.388 ;
  LAYER M3 ;
        RECT 10.928 20.88 10.96 23.388 ;
  LAYER M3 ;
        RECT 10.992 20.88 11.024 23.388 ;
  LAYER M3 ;
        RECT 11.056 20.88 11.088 23.388 ;
  LAYER M3 ;
        RECT 11.12 20.88 11.152 23.388 ;
  LAYER M3 ;
        RECT 11.184 20.88 11.216 23.388 ;
  LAYER M3 ;
        RECT 11.248 20.88 11.28 23.388 ;
  LAYER M3 ;
        RECT 11.312 20.88 11.344 23.388 ;
  LAYER M3 ;
        RECT 11.376 20.88 11.408 23.388 ;
  LAYER M3 ;
        RECT 11.44 20.88 11.472 23.388 ;
  LAYER M3 ;
        RECT 11.504 20.88 11.536 23.388 ;
  LAYER M3 ;
        RECT 11.568 20.88 11.6 23.388 ;
  LAYER M3 ;
        RECT 11.664 20.88 11.696 23.388 ;
  LAYER M1 ;
        RECT 9.279 20.916 9.281 23.352 ;
  LAYER M1 ;
        RECT 9.359 20.916 9.361 23.352 ;
  LAYER M1 ;
        RECT 9.439 20.916 9.441 23.352 ;
  LAYER M1 ;
        RECT 9.519 20.916 9.521 23.352 ;
  LAYER M1 ;
        RECT 9.599 20.916 9.601 23.352 ;
  LAYER M1 ;
        RECT 9.679 20.916 9.681 23.352 ;
  LAYER M1 ;
        RECT 9.759 20.916 9.761 23.352 ;
  LAYER M1 ;
        RECT 9.839 20.916 9.841 23.352 ;
  LAYER M1 ;
        RECT 9.919 20.916 9.921 23.352 ;
  LAYER M1 ;
        RECT 9.999 20.916 10.001 23.352 ;
  LAYER M1 ;
        RECT 10.079 20.916 10.081 23.352 ;
  LAYER M1 ;
        RECT 10.159 20.916 10.161 23.352 ;
  LAYER M1 ;
        RECT 10.239 20.916 10.241 23.352 ;
  LAYER M1 ;
        RECT 10.319 20.916 10.321 23.352 ;
  LAYER M1 ;
        RECT 10.399 20.916 10.401 23.352 ;
  LAYER M1 ;
        RECT 10.479 20.916 10.481 23.352 ;
  LAYER M1 ;
        RECT 10.559 20.916 10.561 23.352 ;
  LAYER M1 ;
        RECT 10.639 20.916 10.641 23.352 ;
  LAYER M1 ;
        RECT 10.719 20.916 10.721 23.352 ;
  LAYER M1 ;
        RECT 10.799 20.916 10.801 23.352 ;
  LAYER M1 ;
        RECT 10.879 20.916 10.881 23.352 ;
  LAYER M1 ;
        RECT 10.959 20.916 10.961 23.352 ;
  LAYER M1 ;
        RECT 11.039 20.916 11.041 23.352 ;
  LAYER M1 ;
        RECT 11.119 20.916 11.121 23.352 ;
  LAYER M1 ;
        RECT 11.199 20.916 11.201 23.352 ;
  LAYER M1 ;
        RECT 11.279 20.916 11.281 23.352 ;
  LAYER M1 ;
        RECT 11.359 20.916 11.361 23.352 ;
  LAYER M1 ;
        RECT 11.439 20.916 11.441 23.352 ;
  LAYER M1 ;
        RECT 11.519 20.916 11.521 23.352 ;
  LAYER M1 ;
        RECT 11.599 20.916 11.601 23.352 ;
  LAYER M2 ;
        RECT 9.28 20.915 11.68 20.917 ;
  LAYER M2 ;
        RECT 9.28 20.999 11.68 21.001 ;
  LAYER M2 ;
        RECT 9.28 21.083 11.68 21.085 ;
  LAYER M2 ;
        RECT 9.28 21.167 11.68 21.169 ;
  LAYER M2 ;
        RECT 9.28 21.251 11.68 21.253 ;
  LAYER M2 ;
        RECT 9.28 21.335 11.68 21.337 ;
  LAYER M2 ;
        RECT 9.28 21.419 11.68 21.421 ;
  LAYER M2 ;
        RECT 9.28 21.503 11.68 21.505 ;
  LAYER M2 ;
        RECT 9.28 21.587 11.68 21.589 ;
  LAYER M2 ;
        RECT 9.28 21.671 11.68 21.673 ;
  LAYER M2 ;
        RECT 9.28 21.755 11.68 21.757 ;
  LAYER M2 ;
        RECT 9.28 21.839 11.68 21.841 ;
  LAYER M2 ;
        RECT 9.28 21.9225 11.68 21.9245 ;
  LAYER M2 ;
        RECT 9.28 22.007 11.68 22.009 ;
  LAYER M2 ;
        RECT 9.28 22.091 11.68 22.093 ;
  LAYER M2 ;
        RECT 9.28 22.175 11.68 22.177 ;
  LAYER M2 ;
        RECT 9.28 22.259 11.68 22.261 ;
  LAYER M2 ;
        RECT 9.28 22.343 11.68 22.345 ;
  LAYER M2 ;
        RECT 9.28 22.427 11.68 22.429 ;
  LAYER M2 ;
        RECT 9.28 22.511 11.68 22.513 ;
  LAYER M2 ;
        RECT 9.28 22.595 11.68 22.597 ;
  LAYER M2 ;
        RECT 9.28 22.679 11.68 22.681 ;
  LAYER M2 ;
        RECT 9.28 22.763 11.68 22.765 ;
  LAYER M2 ;
        RECT 9.28 22.847 11.68 22.849 ;
  LAYER M2 ;
        RECT 9.28 22.931 11.68 22.933 ;
  LAYER M2 ;
        RECT 9.28 23.015 11.68 23.017 ;
  LAYER M2 ;
        RECT 9.28 23.099 11.68 23.101 ;
  LAYER M2 ;
        RECT 9.28 23.183 11.68 23.185 ;
  LAYER M2 ;
        RECT 9.28 23.267 11.68 23.269 ;
  LAYER M1 ;
        RECT 9.264 23.82 9.296 26.328 ;
  LAYER M1 ;
        RECT 9.328 23.82 9.36 26.328 ;
  LAYER M1 ;
        RECT 9.392 23.82 9.424 26.328 ;
  LAYER M1 ;
        RECT 9.456 23.82 9.488 26.328 ;
  LAYER M1 ;
        RECT 9.52 23.82 9.552 26.328 ;
  LAYER M1 ;
        RECT 9.584 23.82 9.616 26.328 ;
  LAYER M1 ;
        RECT 9.648 23.82 9.68 26.328 ;
  LAYER M1 ;
        RECT 9.712 23.82 9.744 26.328 ;
  LAYER M1 ;
        RECT 9.776 23.82 9.808 26.328 ;
  LAYER M1 ;
        RECT 9.84 23.82 9.872 26.328 ;
  LAYER M1 ;
        RECT 9.904 23.82 9.936 26.328 ;
  LAYER M1 ;
        RECT 9.968 23.82 10 26.328 ;
  LAYER M1 ;
        RECT 10.032 23.82 10.064 26.328 ;
  LAYER M1 ;
        RECT 10.096 23.82 10.128 26.328 ;
  LAYER M1 ;
        RECT 10.16 23.82 10.192 26.328 ;
  LAYER M1 ;
        RECT 10.224 23.82 10.256 26.328 ;
  LAYER M1 ;
        RECT 10.288 23.82 10.32 26.328 ;
  LAYER M1 ;
        RECT 10.352 23.82 10.384 26.328 ;
  LAYER M1 ;
        RECT 10.416 23.82 10.448 26.328 ;
  LAYER M1 ;
        RECT 10.48 23.82 10.512 26.328 ;
  LAYER M1 ;
        RECT 10.544 23.82 10.576 26.328 ;
  LAYER M1 ;
        RECT 10.608 23.82 10.64 26.328 ;
  LAYER M1 ;
        RECT 10.672 23.82 10.704 26.328 ;
  LAYER M1 ;
        RECT 10.736 23.82 10.768 26.328 ;
  LAYER M1 ;
        RECT 10.8 23.82 10.832 26.328 ;
  LAYER M1 ;
        RECT 10.864 23.82 10.896 26.328 ;
  LAYER M1 ;
        RECT 10.928 23.82 10.96 26.328 ;
  LAYER M1 ;
        RECT 10.992 23.82 11.024 26.328 ;
  LAYER M1 ;
        RECT 11.056 23.82 11.088 26.328 ;
  LAYER M1 ;
        RECT 11.12 23.82 11.152 26.328 ;
  LAYER M1 ;
        RECT 11.184 23.82 11.216 26.328 ;
  LAYER M1 ;
        RECT 11.248 23.82 11.28 26.328 ;
  LAYER M1 ;
        RECT 11.312 23.82 11.344 26.328 ;
  LAYER M1 ;
        RECT 11.376 23.82 11.408 26.328 ;
  LAYER M1 ;
        RECT 11.44 23.82 11.472 26.328 ;
  LAYER M1 ;
        RECT 11.504 23.82 11.536 26.328 ;
  LAYER M1 ;
        RECT 11.568 23.82 11.6 26.328 ;
  LAYER M2 ;
        RECT 9.244 23.904 11.716 23.936 ;
  LAYER M2 ;
        RECT 9.244 23.968 11.716 24 ;
  LAYER M2 ;
        RECT 9.244 24.032 11.716 24.064 ;
  LAYER M2 ;
        RECT 9.244 24.096 11.716 24.128 ;
  LAYER M2 ;
        RECT 9.244 24.16 11.716 24.192 ;
  LAYER M2 ;
        RECT 9.244 24.224 11.716 24.256 ;
  LAYER M2 ;
        RECT 9.244 24.288 11.716 24.32 ;
  LAYER M2 ;
        RECT 9.244 24.352 11.716 24.384 ;
  LAYER M2 ;
        RECT 9.244 24.416 11.716 24.448 ;
  LAYER M2 ;
        RECT 9.244 24.48 11.716 24.512 ;
  LAYER M2 ;
        RECT 9.244 24.544 11.716 24.576 ;
  LAYER M2 ;
        RECT 9.244 24.608 11.716 24.64 ;
  LAYER M2 ;
        RECT 9.244 24.672 11.716 24.704 ;
  LAYER M2 ;
        RECT 9.244 24.736 11.716 24.768 ;
  LAYER M2 ;
        RECT 9.244 24.8 11.716 24.832 ;
  LAYER M2 ;
        RECT 9.244 24.864 11.716 24.896 ;
  LAYER M2 ;
        RECT 9.244 24.928 11.716 24.96 ;
  LAYER M2 ;
        RECT 9.244 24.992 11.716 25.024 ;
  LAYER M2 ;
        RECT 9.244 25.056 11.716 25.088 ;
  LAYER M2 ;
        RECT 9.244 25.12 11.716 25.152 ;
  LAYER M2 ;
        RECT 9.244 25.184 11.716 25.216 ;
  LAYER M2 ;
        RECT 9.244 25.248 11.716 25.28 ;
  LAYER M2 ;
        RECT 9.244 25.312 11.716 25.344 ;
  LAYER M2 ;
        RECT 9.244 25.376 11.716 25.408 ;
  LAYER M2 ;
        RECT 9.244 25.44 11.716 25.472 ;
  LAYER M2 ;
        RECT 9.244 25.504 11.716 25.536 ;
  LAYER M2 ;
        RECT 9.244 25.568 11.716 25.6 ;
  LAYER M2 ;
        RECT 9.244 25.632 11.716 25.664 ;
  LAYER M2 ;
        RECT 9.244 25.696 11.716 25.728 ;
  LAYER M2 ;
        RECT 9.244 25.76 11.716 25.792 ;
  LAYER M2 ;
        RECT 9.244 25.824 11.716 25.856 ;
  LAYER M2 ;
        RECT 9.244 25.888 11.716 25.92 ;
  LAYER M2 ;
        RECT 9.244 25.952 11.716 25.984 ;
  LAYER M2 ;
        RECT 9.244 26.016 11.716 26.048 ;
  LAYER M2 ;
        RECT 9.244 26.08 11.716 26.112 ;
  LAYER M2 ;
        RECT 9.244 26.144 11.716 26.176 ;
  LAYER M3 ;
        RECT 9.264 23.82 9.296 26.328 ;
  LAYER M3 ;
        RECT 9.328 23.82 9.36 26.328 ;
  LAYER M3 ;
        RECT 9.392 23.82 9.424 26.328 ;
  LAYER M3 ;
        RECT 9.456 23.82 9.488 26.328 ;
  LAYER M3 ;
        RECT 9.52 23.82 9.552 26.328 ;
  LAYER M3 ;
        RECT 9.584 23.82 9.616 26.328 ;
  LAYER M3 ;
        RECT 9.648 23.82 9.68 26.328 ;
  LAYER M3 ;
        RECT 9.712 23.82 9.744 26.328 ;
  LAYER M3 ;
        RECT 9.776 23.82 9.808 26.328 ;
  LAYER M3 ;
        RECT 9.84 23.82 9.872 26.328 ;
  LAYER M3 ;
        RECT 9.904 23.82 9.936 26.328 ;
  LAYER M3 ;
        RECT 9.968 23.82 10 26.328 ;
  LAYER M3 ;
        RECT 10.032 23.82 10.064 26.328 ;
  LAYER M3 ;
        RECT 10.096 23.82 10.128 26.328 ;
  LAYER M3 ;
        RECT 10.16 23.82 10.192 26.328 ;
  LAYER M3 ;
        RECT 10.224 23.82 10.256 26.328 ;
  LAYER M3 ;
        RECT 10.288 23.82 10.32 26.328 ;
  LAYER M3 ;
        RECT 10.352 23.82 10.384 26.328 ;
  LAYER M3 ;
        RECT 10.416 23.82 10.448 26.328 ;
  LAYER M3 ;
        RECT 10.48 23.82 10.512 26.328 ;
  LAYER M3 ;
        RECT 10.544 23.82 10.576 26.328 ;
  LAYER M3 ;
        RECT 10.608 23.82 10.64 26.328 ;
  LAYER M3 ;
        RECT 10.672 23.82 10.704 26.328 ;
  LAYER M3 ;
        RECT 10.736 23.82 10.768 26.328 ;
  LAYER M3 ;
        RECT 10.8 23.82 10.832 26.328 ;
  LAYER M3 ;
        RECT 10.864 23.82 10.896 26.328 ;
  LAYER M3 ;
        RECT 10.928 23.82 10.96 26.328 ;
  LAYER M3 ;
        RECT 10.992 23.82 11.024 26.328 ;
  LAYER M3 ;
        RECT 11.056 23.82 11.088 26.328 ;
  LAYER M3 ;
        RECT 11.12 23.82 11.152 26.328 ;
  LAYER M3 ;
        RECT 11.184 23.82 11.216 26.328 ;
  LAYER M3 ;
        RECT 11.248 23.82 11.28 26.328 ;
  LAYER M3 ;
        RECT 11.312 23.82 11.344 26.328 ;
  LAYER M3 ;
        RECT 11.376 23.82 11.408 26.328 ;
  LAYER M3 ;
        RECT 11.44 23.82 11.472 26.328 ;
  LAYER M3 ;
        RECT 11.504 23.82 11.536 26.328 ;
  LAYER M3 ;
        RECT 11.568 23.82 11.6 26.328 ;
  LAYER M3 ;
        RECT 11.664 23.82 11.696 26.328 ;
  LAYER M1 ;
        RECT 9.279 23.856 9.281 26.292 ;
  LAYER M1 ;
        RECT 9.359 23.856 9.361 26.292 ;
  LAYER M1 ;
        RECT 9.439 23.856 9.441 26.292 ;
  LAYER M1 ;
        RECT 9.519 23.856 9.521 26.292 ;
  LAYER M1 ;
        RECT 9.599 23.856 9.601 26.292 ;
  LAYER M1 ;
        RECT 9.679 23.856 9.681 26.292 ;
  LAYER M1 ;
        RECT 9.759 23.856 9.761 26.292 ;
  LAYER M1 ;
        RECT 9.839 23.856 9.841 26.292 ;
  LAYER M1 ;
        RECT 9.919 23.856 9.921 26.292 ;
  LAYER M1 ;
        RECT 9.999 23.856 10.001 26.292 ;
  LAYER M1 ;
        RECT 10.079 23.856 10.081 26.292 ;
  LAYER M1 ;
        RECT 10.159 23.856 10.161 26.292 ;
  LAYER M1 ;
        RECT 10.239 23.856 10.241 26.292 ;
  LAYER M1 ;
        RECT 10.319 23.856 10.321 26.292 ;
  LAYER M1 ;
        RECT 10.399 23.856 10.401 26.292 ;
  LAYER M1 ;
        RECT 10.479 23.856 10.481 26.292 ;
  LAYER M1 ;
        RECT 10.559 23.856 10.561 26.292 ;
  LAYER M1 ;
        RECT 10.639 23.856 10.641 26.292 ;
  LAYER M1 ;
        RECT 10.719 23.856 10.721 26.292 ;
  LAYER M1 ;
        RECT 10.799 23.856 10.801 26.292 ;
  LAYER M1 ;
        RECT 10.879 23.856 10.881 26.292 ;
  LAYER M1 ;
        RECT 10.959 23.856 10.961 26.292 ;
  LAYER M1 ;
        RECT 11.039 23.856 11.041 26.292 ;
  LAYER M1 ;
        RECT 11.119 23.856 11.121 26.292 ;
  LAYER M1 ;
        RECT 11.199 23.856 11.201 26.292 ;
  LAYER M1 ;
        RECT 11.279 23.856 11.281 26.292 ;
  LAYER M1 ;
        RECT 11.359 23.856 11.361 26.292 ;
  LAYER M1 ;
        RECT 11.439 23.856 11.441 26.292 ;
  LAYER M1 ;
        RECT 11.519 23.856 11.521 26.292 ;
  LAYER M1 ;
        RECT 11.599 23.856 11.601 26.292 ;
  LAYER M2 ;
        RECT 9.28 23.855 11.68 23.857 ;
  LAYER M2 ;
        RECT 9.28 23.939 11.68 23.941 ;
  LAYER M2 ;
        RECT 9.28 24.023 11.68 24.025 ;
  LAYER M2 ;
        RECT 9.28 24.107 11.68 24.109 ;
  LAYER M2 ;
        RECT 9.28 24.191 11.68 24.193 ;
  LAYER M2 ;
        RECT 9.28 24.275 11.68 24.277 ;
  LAYER M2 ;
        RECT 9.28 24.359 11.68 24.361 ;
  LAYER M2 ;
        RECT 9.28 24.443 11.68 24.445 ;
  LAYER M2 ;
        RECT 9.28 24.527 11.68 24.529 ;
  LAYER M2 ;
        RECT 9.28 24.611 11.68 24.613 ;
  LAYER M2 ;
        RECT 9.28 24.695 11.68 24.697 ;
  LAYER M2 ;
        RECT 9.28 24.779 11.68 24.781 ;
  LAYER M2 ;
        RECT 9.28 24.8625 11.68 24.8645 ;
  LAYER M2 ;
        RECT 9.28 24.947 11.68 24.949 ;
  LAYER M2 ;
        RECT 9.28 25.031 11.68 25.033 ;
  LAYER M2 ;
        RECT 9.28 25.115 11.68 25.117 ;
  LAYER M2 ;
        RECT 9.28 25.199 11.68 25.201 ;
  LAYER M2 ;
        RECT 9.28 25.283 11.68 25.285 ;
  LAYER M2 ;
        RECT 9.28 25.367 11.68 25.369 ;
  LAYER M2 ;
        RECT 9.28 25.451 11.68 25.453 ;
  LAYER M2 ;
        RECT 9.28 25.535 11.68 25.537 ;
  LAYER M2 ;
        RECT 9.28 25.619 11.68 25.621 ;
  LAYER M2 ;
        RECT 9.28 25.703 11.68 25.705 ;
  LAYER M2 ;
        RECT 9.28 25.787 11.68 25.789 ;
  LAYER M2 ;
        RECT 9.28 25.871 11.68 25.873 ;
  LAYER M2 ;
        RECT 9.28 25.955 11.68 25.957 ;
  LAYER M2 ;
        RECT 9.28 26.039 11.68 26.041 ;
  LAYER M2 ;
        RECT 9.28 26.123 11.68 26.125 ;
  LAYER M2 ;
        RECT 9.28 26.207 11.68 26.209 ;
  LAYER M1 ;
        RECT 9.264 26.76 9.296 29.268 ;
  LAYER M1 ;
        RECT 9.328 26.76 9.36 29.268 ;
  LAYER M1 ;
        RECT 9.392 26.76 9.424 29.268 ;
  LAYER M1 ;
        RECT 9.456 26.76 9.488 29.268 ;
  LAYER M1 ;
        RECT 9.52 26.76 9.552 29.268 ;
  LAYER M1 ;
        RECT 9.584 26.76 9.616 29.268 ;
  LAYER M1 ;
        RECT 9.648 26.76 9.68 29.268 ;
  LAYER M1 ;
        RECT 9.712 26.76 9.744 29.268 ;
  LAYER M1 ;
        RECT 9.776 26.76 9.808 29.268 ;
  LAYER M1 ;
        RECT 9.84 26.76 9.872 29.268 ;
  LAYER M1 ;
        RECT 9.904 26.76 9.936 29.268 ;
  LAYER M1 ;
        RECT 9.968 26.76 10 29.268 ;
  LAYER M1 ;
        RECT 10.032 26.76 10.064 29.268 ;
  LAYER M1 ;
        RECT 10.096 26.76 10.128 29.268 ;
  LAYER M1 ;
        RECT 10.16 26.76 10.192 29.268 ;
  LAYER M1 ;
        RECT 10.224 26.76 10.256 29.268 ;
  LAYER M1 ;
        RECT 10.288 26.76 10.32 29.268 ;
  LAYER M1 ;
        RECT 10.352 26.76 10.384 29.268 ;
  LAYER M1 ;
        RECT 10.416 26.76 10.448 29.268 ;
  LAYER M1 ;
        RECT 10.48 26.76 10.512 29.268 ;
  LAYER M1 ;
        RECT 10.544 26.76 10.576 29.268 ;
  LAYER M1 ;
        RECT 10.608 26.76 10.64 29.268 ;
  LAYER M1 ;
        RECT 10.672 26.76 10.704 29.268 ;
  LAYER M1 ;
        RECT 10.736 26.76 10.768 29.268 ;
  LAYER M1 ;
        RECT 10.8 26.76 10.832 29.268 ;
  LAYER M1 ;
        RECT 10.864 26.76 10.896 29.268 ;
  LAYER M1 ;
        RECT 10.928 26.76 10.96 29.268 ;
  LAYER M1 ;
        RECT 10.992 26.76 11.024 29.268 ;
  LAYER M1 ;
        RECT 11.056 26.76 11.088 29.268 ;
  LAYER M1 ;
        RECT 11.12 26.76 11.152 29.268 ;
  LAYER M1 ;
        RECT 11.184 26.76 11.216 29.268 ;
  LAYER M1 ;
        RECT 11.248 26.76 11.28 29.268 ;
  LAYER M1 ;
        RECT 11.312 26.76 11.344 29.268 ;
  LAYER M1 ;
        RECT 11.376 26.76 11.408 29.268 ;
  LAYER M1 ;
        RECT 11.44 26.76 11.472 29.268 ;
  LAYER M1 ;
        RECT 11.504 26.76 11.536 29.268 ;
  LAYER M1 ;
        RECT 11.568 26.76 11.6 29.268 ;
  LAYER M2 ;
        RECT 9.244 26.844 11.716 26.876 ;
  LAYER M2 ;
        RECT 9.244 26.908 11.716 26.94 ;
  LAYER M2 ;
        RECT 9.244 26.972 11.716 27.004 ;
  LAYER M2 ;
        RECT 9.244 27.036 11.716 27.068 ;
  LAYER M2 ;
        RECT 9.244 27.1 11.716 27.132 ;
  LAYER M2 ;
        RECT 9.244 27.164 11.716 27.196 ;
  LAYER M2 ;
        RECT 9.244 27.228 11.716 27.26 ;
  LAYER M2 ;
        RECT 9.244 27.292 11.716 27.324 ;
  LAYER M2 ;
        RECT 9.244 27.356 11.716 27.388 ;
  LAYER M2 ;
        RECT 9.244 27.42 11.716 27.452 ;
  LAYER M2 ;
        RECT 9.244 27.484 11.716 27.516 ;
  LAYER M2 ;
        RECT 9.244 27.548 11.716 27.58 ;
  LAYER M2 ;
        RECT 9.244 27.612 11.716 27.644 ;
  LAYER M2 ;
        RECT 9.244 27.676 11.716 27.708 ;
  LAYER M2 ;
        RECT 9.244 27.74 11.716 27.772 ;
  LAYER M2 ;
        RECT 9.244 27.804 11.716 27.836 ;
  LAYER M2 ;
        RECT 9.244 27.868 11.716 27.9 ;
  LAYER M2 ;
        RECT 9.244 27.932 11.716 27.964 ;
  LAYER M2 ;
        RECT 9.244 27.996 11.716 28.028 ;
  LAYER M2 ;
        RECT 9.244 28.06 11.716 28.092 ;
  LAYER M2 ;
        RECT 9.244 28.124 11.716 28.156 ;
  LAYER M2 ;
        RECT 9.244 28.188 11.716 28.22 ;
  LAYER M2 ;
        RECT 9.244 28.252 11.716 28.284 ;
  LAYER M2 ;
        RECT 9.244 28.316 11.716 28.348 ;
  LAYER M2 ;
        RECT 9.244 28.38 11.716 28.412 ;
  LAYER M2 ;
        RECT 9.244 28.444 11.716 28.476 ;
  LAYER M2 ;
        RECT 9.244 28.508 11.716 28.54 ;
  LAYER M2 ;
        RECT 9.244 28.572 11.716 28.604 ;
  LAYER M2 ;
        RECT 9.244 28.636 11.716 28.668 ;
  LAYER M2 ;
        RECT 9.244 28.7 11.716 28.732 ;
  LAYER M2 ;
        RECT 9.244 28.764 11.716 28.796 ;
  LAYER M2 ;
        RECT 9.244 28.828 11.716 28.86 ;
  LAYER M2 ;
        RECT 9.244 28.892 11.716 28.924 ;
  LAYER M2 ;
        RECT 9.244 28.956 11.716 28.988 ;
  LAYER M2 ;
        RECT 9.244 29.02 11.716 29.052 ;
  LAYER M2 ;
        RECT 9.244 29.084 11.716 29.116 ;
  LAYER M3 ;
        RECT 9.264 26.76 9.296 29.268 ;
  LAYER M3 ;
        RECT 9.328 26.76 9.36 29.268 ;
  LAYER M3 ;
        RECT 9.392 26.76 9.424 29.268 ;
  LAYER M3 ;
        RECT 9.456 26.76 9.488 29.268 ;
  LAYER M3 ;
        RECT 9.52 26.76 9.552 29.268 ;
  LAYER M3 ;
        RECT 9.584 26.76 9.616 29.268 ;
  LAYER M3 ;
        RECT 9.648 26.76 9.68 29.268 ;
  LAYER M3 ;
        RECT 9.712 26.76 9.744 29.268 ;
  LAYER M3 ;
        RECT 9.776 26.76 9.808 29.268 ;
  LAYER M3 ;
        RECT 9.84 26.76 9.872 29.268 ;
  LAYER M3 ;
        RECT 9.904 26.76 9.936 29.268 ;
  LAYER M3 ;
        RECT 9.968 26.76 10 29.268 ;
  LAYER M3 ;
        RECT 10.032 26.76 10.064 29.268 ;
  LAYER M3 ;
        RECT 10.096 26.76 10.128 29.268 ;
  LAYER M3 ;
        RECT 10.16 26.76 10.192 29.268 ;
  LAYER M3 ;
        RECT 10.224 26.76 10.256 29.268 ;
  LAYER M3 ;
        RECT 10.288 26.76 10.32 29.268 ;
  LAYER M3 ;
        RECT 10.352 26.76 10.384 29.268 ;
  LAYER M3 ;
        RECT 10.416 26.76 10.448 29.268 ;
  LAYER M3 ;
        RECT 10.48 26.76 10.512 29.268 ;
  LAYER M3 ;
        RECT 10.544 26.76 10.576 29.268 ;
  LAYER M3 ;
        RECT 10.608 26.76 10.64 29.268 ;
  LAYER M3 ;
        RECT 10.672 26.76 10.704 29.268 ;
  LAYER M3 ;
        RECT 10.736 26.76 10.768 29.268 ;
  LAYER M3 ;
        RECT 10.8 26.76 10.832 29.268 ;
  LAYER M3 ;
        RECT 10.864 26.76 10.896 29.268 ;
  LAYER M3 ;
        RECT 10.928 26.76 10.96 29.268 ;
  LAYER M3 ;
        RECT 10.992 26.76 11.024 29.268 ;
  LAYER M3 ;
        RECT 11.056 26.76 11.088 29.268 ;
  LAYER M3 ;
        RECT 11.12 26.76 11.152 29.268 ;
  LAYER M3 ;
        RECT 11.184 26.76 11.216 29.268 ;
  LAYER M3 ;
        RECT 11.248 26.76 11.28 29.268 ;
  LAYER M3 ;
        RECT 11.312 26.76 11.344 29.268 ;
  LAYER M3 ;
        RECT 11.376 26.76 11.408 29.268 ;
  LAYER M3 ;
        RECT 11.44 26.76 11.472 29.268 ;
  LAYER M3 ;
        RECT 11.504 26.76 11.536 29.268 ;
  LAYER M3 ;
        RECT 11.568 26.76 11.6 29.268 ;
  LAYER M3 ;
        RECT 11.664 26.76 11.696 29.268 ;
  LAYER M1 ;
        RECT 9.279 26.796 9.281 29.232 ;
  LAYER M1 ;
        RECT 9.359 26.796 9.361 29.232 ;
  LAYER M1 ;
        RECT 9.439 26.796 9.441 29.232 ;
  LAYER M1 ;
        RECT 9.519 26.796 9.521 29.232 ;
  LAYER M1 ;
        RECT 9.599 26.796 9.601 29.232 ;
  LAYER M1 ;
        RECT 9.679 26.796 9.681 29.232 ;
  LAYER M1 ;
        RECT 9.759 26.796 9.761 29.232 ;
  LAYER M1 ;
        RECT 9.839 26.796 9.841 29.232 ;
  LAYER M1 ;
        RECT 9.919 26.796 9.921 29.232 ;
  LAYER M1 ;
        RECT 9.999 26.796 10.001 29.232 ;
  LAYER M1 ;
        RECT 10.079 26.796 10.081 29.232 ;
  LAYER M1 ;
        RECT 10.159 26.796 10.161 29.232 ;
  LAYER M1 ;
        RECT 10.239 26.796 10.241 29.232 ;
  LAYER M1 ;
        RECT 10.319 26.796 10.321 29.232 ;
  LAYER M1 ;
        RECT 10.399 26.796 10.401 29.232 ;
  LAYER M1 ;
        RECT 10.479 26.796 10.481 29.232 ;
  LAYER M1 ;
        RECT 10.559 26.796 10.561 29.232 ;
  LAYER M1 ;
        RECT 10.639 26.796 10.641 29.232 ;
  LAYER M1 ;
        RECT 10.719 26.796 10.721 29.232 ;
  LAYER M1 ;
        RECT 10.799 26.796 10.801 29.232 ;
  LAYER M1 ;
        RECT 10.879 26.796 10.881 29.232 ;
  LAYER M1 ;
        RECT 10.959 26.796 10.961 29.232 ;
  LAYER M1 ;
        RECT 11.039 26.796 11.041 29.232 ;
  LAYER M1 ;
        RECT 11.119 26.796 11.121 29.232 ;
  LAYER M1 ;
        RECT 11.199 26.796 11.201 29.232 ;
  LAYER M1 ;
        RECT 11.279 26.796 11.281 29.232 ;
  LAYER M1 ;
        RECT 11.359 26.796 11.361 29.232 ;
  LAYER M1 ;
        RECT 11.439 26.796 11.441 29.232 ;
  LAYER M1 ;
        RECT 11.519 26.796 11.521 29.232 ;
  LAYER M1 ;
        RECT 11.599 26.796 11.601 29.232 ;
  LAYER M2 ;
        RECT 9.28 26.795 11.68 26.797 ;
  LAYER M2 ;
        RECT 9.28 26.879 11.68 26.881 ;
  LAYER M2 ;
        RECT 9.28 26.963 11.68 26.965 ;
  LAYER M2 ;
        RECT 9.28 27.047 11.68 27.049 ;
  LAYER M2 ;
        RECT 9.28 27.131 11.68 27.133 ;
  LAYER M2 ;
        RECT 9.28 27.215 11.68 27.217 ;
  LAYER M2 ;
        RECT 9.28 27.299 11.68 27.301 ;
  LAYER M2 ;
        RECT 9.28 27.383 11.68 27.385 ;
  LAYER M2 ;
        RECT 9.28 27.467 11.68 27.469 ;
  LAYER M2 ;
        RECT 9.28 27.551 11.68 27.553 ;
  LAYER M2 ;
        RECT 9.28 27.635 11.68 27.637 ;
  LAYER M2 ;
        RECT 9.28 27.719 11.68 27.721 ;
  LAYER M2 ;
        RECT 9.28 27.8025 11.68 27.8045 ;
  LAYER M2 ;
        RECT 9.28 27.887 11.68 27.889 ;
  LAYER M2 ;
        RECT 9.28 27.971 11.68 27.973 ;
  LAYER M2 ;
        RECT 9.28 28.055 11.68 28.057 ;
  LAYER M2 ;
        RECT 9.28 28.139 11.68 28.141 ;
  LAYER M2 ;
        RECT 9.28 28.223 11.68 28.225 ;
  LAYER M2 ;
        RECT 9.28 28.307 11.68 28.309 ;
  LAYER M2 ;
        RECT 9.28 28.391 11.68 28.393 ;
  LAYER M2 ;
        RECT 9.28 28.475 11.68 28.477 ;
  LAYER M2 ;
        RECT 9.28 28.559 11.68 28.561 ;
  LAYER M2 ;
        RECT 9.28 28.643 11.68 28.645 ;
  LAYER M2 ;
        RECT 9.28 28.727 11.68 28.729 ;
  LAYER M2 ;
        RECT 9.28 28.811 11.68 28.813 ;
  LAYER M2 ;
        RECT 9.28 28.895 11.68 28.897 ;
  LAYER M2 ;
        RECT 9.28 28.979 11.68 28.981 ;
  LAYER M2 ;
        RECT 9.28 29.063 11.68 29.065 ;
  LAYER M2 ;
        RECT 9.28 29.147 11.68 29.149 ;
  LAYER M1 ;
        RECT 12.144 17.94 12.176 20.448 ;
  LAYER M1 ;
        RECT 12.208 17.94 12.24 20.448 ;
  LAYER M1 ;
        RECT 12.272 17.94 12.304 20.448 ;
  LAYER M1 ;
        RECT 12.336 17.94 12.368 20.448 ;
  LAYER M1 ;
        RECT 12.4 17.94 12.432 20.448 ;
  LAYER M1 ;
        RECT 12.464 17.94 12.496 20.448 ;
  LAYER M1 ;
        RECT 12.528 17.94 12.56 20.448 ;
  LAYER M1 ;
        RECT 12.592 17.94 12.624 20.448 ;
  LAYER M1 ;
        RECT 12.656 17.94 12.688 20.448 ;
  LAYER M1 ;
        RECT 12.72 17.94 12.752 20.448 ;
  LAYER M1 ;
        RECT 12.784 17.94 12.816 20.448 ;
  LAYER M1 ;
        RECT 12.848 17.94 12.88 20.448 ;
  LAYER M1 ;
        RECT 12.912 17.94 12.944 20.448 ;
  LAYER M1 ;
        RECT 12.976 17.94 13.008 20.448 ;
  LAYER M1 ;
        RECT 13.04 17.94 13.072 20.448 ;
  LAYER M1 ;
        RECT 13.104 17.94 13.136 20.448 ;
  LAYER M1 ;
        RECT 13.168 17.94 13.2 20.448 ;
  LAYER M1 ;
        RECT 13.232 17.94 13.264 20.448 ;
  LAYER M1 ;
        RECT 13.296 17.94 13.328 20.448 ;
  LAYER M1 ;
        RECT 13.36 17.94 13.392 20.448 ;
  LAYER M1 ;
        RECT 13.424 17.94 13.456 20.448 ;
  LAYER M1 ;
        RECT 13.488 17.94 13.52 20.448 ;
  LAYER M1 ;
        RECT 13.552 17.94 13.584 20.448 ;
  LAYER M1 ;
        RECT 13.616 17.94 13.648 20.448 ;
  LAYER M1 ;
        RECT 13.68 17.94 13.712 20.448 ;
  LAYER M1 ;
        RECT 13.744 17.94 13.776 20.448 ;
  LAYER M1 ;
        RECT 13.808 17.94 13.84 20.448 ;
  LAYER M1 ;
        RECT 13.872 17.94 13.904 20.448 ;
  LAYER M1 ;
        RECT 13.936 17.94 13.968 20.448 ;
  LAYER M1 ;
        RECT 14 17.94 14.032 20.448 ;
  LAYER M1 ;
        RECT 14.064 17.94 14.096 20.448 ;
  LAYER M1 ;
        RECT 14.128 17.94 14.16 20.448 ;
  LAYER M1 ;
        RECT 14.192 17.94 14.224 20.448 ;
  LAYER M1 ;
        RECT 14.256 17.94 14.288 20.448 ;
  LAYER M1 ;
        RECT 14.32 17.94 14.352 20.448 ;
  LAYER M1 ;
        RECT 14.384 17.94 14.416 20.448 ;
  LAYER M1 ;
        RECT 14.448 17.94 14.48 20.448 ;
  LAYER M2 ;
        RECT 12.124 18.024 14.596 18.056 ;
  LAYER M2 ;
        RECT 12.124 18.088 14.596 18.12 ;
  LAYER M2 ;
        RECT 12.124 18.152 14.596 18.184 ;
  LAYER M2 ;
        RECT 12.124 18.216 14.596 18.248 ;
  LAYER M2 ;
        RECT 12.124 18.28 14.596 18.312 ;
  LAYER M2 ;
        RECT 12.124 18.344 14.596 18.376 ;
  LAYER M2 ;
        RECT 12.124 18.408 14.596 18.44 ;
  LAYER M2 ;
        RECT 12.124 18.472 14.596 18.504 ;
  LAYER M2 ;
        RECT 12.124 18.536 14.596 18.568 ;
  LAYER M2 ;
        RECT 12.124 18.6 14.596 18.632 ;
  LAYER M2 ;
        RECT 12.124 18.664 14.596 18.696 ;
  LAYER M2 ;
        RECT 12.124 18.728 14.596 18.76 ;
  LAYER M2 ;
        RECT 12.124 18.792 14.596 18.824 ;
  LAYER M2 ;
        RECT 12.124 18.856 14.596 18.888 ;
  LAYER M2 ;
        RECT 12.124 18.92 14.596 18.952 ;
  LAYER M2 ;
        RECT 12.124 18.984 14.596 19.016 ;
  LAYER M2 ;
        RECT 12.124 19.048 14.596 19.08 ;
  LAYER M2 ;
        RECT 12.124 19.112 14.596 19.144 ;
  LAYER M2 ;
        RECT 12.124 19.176 14.596 19.208 ;
  LAYER M2 ;
        RECT 12.124 19.24 14.596 19.272 ;
  LAYER M2 ;
        RECT 12.124 19.304 14.596 19.336 ;
  LAYER M2 ;
        RECT 12.124 19.368 14.596 19.4 ;
  LAYER M2 ;
        RECT 12.124 19.432 14.596 19.464 ;
  LAYER M2 ;
        RECT 12.124 19.496 14.596 19.528 ;
  LAYER M2 ;
        RECT 12.124 19.56 14.596 19.592 ;
  LAYER M2 ;
        RECT 12.124 19.624 14.596 19.656 ;
  LAYER M2 ;
        RECT 12.124 19.688 14.596 19.72 ;
  LAYER M2 ;
        RECT 12.124 19.752 14.596 19.784 ;
  LAYER M2 ;
        RECT 12.124 19.816 14.596 19.848 ;
  LAYER M2 ;
        RECT 12.124 19.88 14.596 19.912 ;
  LAYER M2 ;
        RECT 12.124 19.944 14.596 19.976 ;
  LAYER M2 ;
        RECT 12.124 20.008 14.596 20.04 ;
  LAYER M2 ;
        RECT 12.124 20.072 14.596 20.104 ;
  LAYER M2 ;
        RECT 12.124 20.136 14.596 20.168 ;
  LAYER M2 ;
        RECT 12.124 20.2 14.596 20.232 ;
  LAYER M2 ;
        RECT 12.124 20.264 14.596 20.296 ;
  LAYER M3 ;
        RECT 12.144 17.94 12.176 20.448 ;
  LAYER M3 ;
        RECT 12.208 17.94 12.24 20.448 ;
  LAYER M3 ;
        RECT 12.272 17.94 12.304 20.448 ;
  LAYER M3 ;
        RECT 12.336 17.94 12.368 20.448 ;
  LAYER M3 ;
        RECT 12.4 17.94 12.432 20.448 ;
  LAYER M3 ;
        RECT 12.464 17.94 12.496 20.448 ;
  LAYER M3 ;
        RECT 12.528 17.94 12.56 20.448 ;
  LAYER M3 ;
        RECT 12.592 17.94 12.624 20.448 ;
  LAYER M3 ;
        RECT 12.656 17.94 12.688 20.448 ;
  LAYER M3 ;
        RECT 12.72 17.94 12.752 20.448 ;
  LAYER M3 ;
        RECT 12.784 17.94 12.816 20.448 ;
  LAYER M3 ;
        RECT 12.848 17.94 12.88 20.448 ;
  LAYER M3 ;
        RECT 12.912 17.94 12.944 20.448 ;
  LAYER M3 ;
        RECT 12.976 17.94 13.008 20.448 ;
  LAYER M3 ;
        RECT 13.04 17.94 13.072 20.448 ;
  LAYER M3 ;
        RECT 13.104 17.94 13.136 20.448 ;
  LAYER M3 ;
        RECT 13.168 17.94 13.2 20.448 ;
  LAYER M3 ;
        RECT 13.232 17.94 13.264 20.448 ;
  LAYER M3 ;
        RECT 13.296 17.94 13.328 20.448 ;
  LAYER M3 ;
        RECT 13.36 17.94 13.392 20.448 ;
  LAYER M3 ;
        RECT 13.424 17.94 13.456 20.448 ;
  LAYER M3 ;
        RECT 13.488 17.94 13.52 20.448 ;
  LAYER M3 ;
        RECT 13.552 17.94 13.584 20.448 ;
  LAYER M3 ;
        RECT 13.616 17.94 13.648 20.448 ;
  LAYER M3 ;
        RECT 13.68 17.94 13.712 20.448 ;
  LAYER M3 ;
        RECT 13.744 17.94 13.776 20.448 ;
  LAYER M3 ;
        RECT 13.808 17.94 13.84 20.448 ;
  LAYER M3 ;
        RECT 13.872 17.94 13.904 20.448 ;
  LAYER M3 ;
        RECT 13.936 17.94 13.968 20.448 ;
  LAYER M3 ;
        RECT 14 17.94 14.032 20.448 ;
  LAYER M3 ;
        RECT 14.064 17.94 14.096 20.448 ;
  LAYER M3 ;
        RECT 14.128 17.94 14.16 20.448 ;
  LAYER M3 ;
        RECT 14.192 17.94 14.224 20.448 ;
  LAYER M3 ;
        RECT 14.256 17.94 14.288 20.448 ;
  LAYER M3 ;
        RECT 14.32 17.94 14.352 20.448 ;
  LAYER M3 ;
        RECT 14.384 17.94 14.416 20.448 ;
  LAYER M3 ;
        RECT 14.448 17.94 14.48 20.448 ;
  LAYER M3 ;
        RECT 14.544 17.94 14.576 20.448 ;
  LAYER M1 ;
        RECT 12.159 17.976 12.161 20.412 ;
  LAYER M1 ;
        RECT 12.239 17.976 12.241 20.412 ;
  LAYER M1 ;
        RECT 12.319 17.976 12.321 20.412 ;
  LAYER M1 ;
        RECT 12.399 17.976 12.401 20.412 ;
  LAYER M1 ;
        RECT 12.479 17.976 12.481 20.412 ;
  LAYER M1 ;
        RECT 12.559 17.976 12.561 20.412 ;
  LAYER M1 ;
        RECT 12.639 17.976 12.641 20.412 ;
  LAYER M1 ;
        RECT 12.719 17.976 12.721 20.412 ;
  LAYER M1 ;
        RECT 12.799 17.976 12.801 20.412 ;
  LAYER M1 ;
        RECT 12.879 17.976 12.881 20.412 ;
  LAYER M1 ;
        RECT 12.959 17.976 12.961 20.412 ;
  LAYER M1 ;
        RECT 13.039 17.976 13.041 20.412 ;
  LAYER M1 ;
        RECT 13.119 17.976 13.121 20.412 ;
  LAYER M1 ;
        RECT 13.199 17.976 13.201 20.412 ;
  LAYER M1 ;
        RECT 13.279 17.976 13.281 20.412 ;
  LAYER M1 ;
        RECT 13.359 17.976 13.361 20.412 ;
  LAYER M1 ;
        RECT 13.439 17.976 13.441 20.412 ;
  LAYER M1 ;
        RECT 13.519 17.976 13.521 20.412 ;
  LAYER M1 ;
        RECT 13.599 17.976 13.601 20.412 ;
  LAYER M1 ;
        RECT 13.679 17.976 13.681 20.412 ;
  LAYER M1 ;
        RECT 13.759 17.976 13.761 20.412 ;
  LAYER M1 ;
        RECT 13.839 17.976 13.841 20.412 ;
  LAYER M1 ;
        RECT 13.919 17.976 13.921 20.412 ;
  LAYER M1 ;
        RECT 13.999 17.976 14.001 20.412 ;
  LAYER M1 ;
        RECT 14.079 17.976 14.081 20.412 ;
  LAYER M1 ;
        RECT 14.159 17.976 14.161 20.412 ;
  LAYER M1 ;
        RECT 14.239 17.976 14.241 20.412 ;
  LAYER M1 ;
        RECT 14.319 17.976 14.321 20.412 ;
  LAYER M1 ;
        RECT 14.399 17.976 14.401 20.412 ;
  LAYER M1 ;
        RECT 14.479 17.976 14.481 20.412 ;
  LAYER M2 ;
        RECT 12.16 17.975 14.56 17.977 ;
  LAYER M2 ;
        RECT 12.16 18.059 14.56 18.061 ;
  LAYER M2 ;
        RECT 12.16 18.143 14.56 18.145 ;
  LAYER M2 ;
        RECT 12.16 18.227 14.56 18.229 ;
  LAYER M2 ;
        RECT 12.16 18.311 14.56 18.313 ;
  LAYER M2 ;
        RECT 12.16 18.395 14.56 18.397 ;
  LAYER M2 ;
        RECT 12.16 18.479 14.56 18.481 ;
  LAYER M2 ;
        RECT 12.16 18.563 14.56 18.565 ;
  LAYER M2 ;
        RECT 12.16 18.647 14.56 18.649 ;
  LAYER M2 ;
        RECT 12.16 18.731 14.56 18.733 ;
  LAYER M2 ;
        RECT 12.16 18.815 14.56 18.817 ;
  LAYER M2 ;
        RECT 12.16 18.899 14.56 18.901 ;
  LAYER M2 ;
        RECT 12.16 18.9825 14.56 18.9845 ;
  LAYER M2 ;
        RECT 12.16 19.067 14.56 19.069 ;
  LAYER M2 ;
        RECT 12.16 19.151 14.56 19.153 ;
  LAYER M2 ;
        RECT 12.16 19.235 14.56 19.237 ;
  LAYER M2 ;
        RECT 12.16 19.319 14.56 19.321 ;
  LAYER M2 ;
        RECT 12.16 19.403 14.56 19.405 ;
  LAYER M2 ;
        RECT 12.16 19.487 14.56 19.489 ;
  LAYER M2 ;
        RECT 12.16 19.571 14.56 19.573 ;
  LAYER M2 ;
        RECT 12.16 19.655 14.56 19.657 ;
  LAYER M2 ;
        RECT 12.16 19.739 14.56 19.741 ;
  LAYER M2 ;
        RECT 12.16 19.823 14.56 19.825 ;
  LAYER M2 ;
        RECT 12.16 19.907 14.56 19.909 ;
  LAYER M2 ;
        RECT 12.16 19.991 14.56 19.993 ;
  LAYER M2 ;
        RECT 12.16 20.075 14.56 20.077 ;
  LAYER M2 ;
        RECT 12.16 20.159 14.56 20.161 ;
  LAYER M2 ;
        RECT 12.16 20.243 14.56 20.245 ;
  LAYER M2 ;
        RECT 12.16 20.327 14.56 20.329 ;
  LAYER M1 ;
        RECT 12.144 20.88 12.176 23.388 ;
  LAYER M1 ;
        RECT 12.208 20.88 12.24 23.388 ;
  LAYER M1 ;
        RECT 12.272 20.88 12.304 23.388 ;
  LAYER M1 ;
        RECT 12.336 20.88 12.368 23.388 ;
  LAYER M1 ;
        RECT 12.4 20.88 12.432 23.388 ;
  LAYER M1 ;
        RECT 12.464 20.88 12.496 23.388 ;
  LAYER M1 ;
        RECT 12.528 20.88 12.56 23.388 ;
  LAYER M1 ;
        RECT 12.592 20.88 12.624 23.388 ;
  LAYER M1 ;
        RECT 12.656 20.88 12.688 23.388 ;
  LAYER M1 ;
        RECT 12.72 20.88 12.752 23.388 ;
  LAYER M1 ;
        RECT 12.784 20.88 12.816 23.388 ;
  LAYER M1 ;
        RECT 12.848 20.88 12.88 23.388 ;
  LAYER M1 ;
        RECT 12.912 20.88 12.944 23.388 ;
  LAYER M1 ;
        RECT 12.976 20.88 13.008 23.388 ;
  LAYER M1 ;
        RECT 13.04 20.88 13.072 23.388 ;
  LAYER M1 ;
        RECT 13.104 20.88 13.136 23.388 ;
  LAYER M1 ;
        RECT 13.168 20.88 13.2 23.388 ;
  LAYER M1 ;
        RECT 13.232 20.88 13.264 23.388 ;
  LAYER M1 ;
        RECT 13.296 20.88 13.328 23.388 ;
  LAYER M1 ;
        RECT 13.36 20.88 13.392 23.388 ;
  LAYER M1 ;
        RECT 13.424 20.88 13.456 23.388 ;
  LAYER M1 ;
        RECT 13.488 20.88 13.52 23.388 ;
  LAYER M1 ;
        RECT 13.552 20.88 13.584 23.388 ;
  LAYER M1 ;
        RECT 13.616 20.88 13.648 23.388 ;
  LAYER M1 ;
        RECT 13.68 20.88 13.712 23.388 ;
  LAYER M1 ;
        RECT 13.744 20.88 13.776 23.388 ;
  LAYER M1 ;
        RECT 13.808 20.88 13.84 23.388 ;
  LAYER M1 ;
        RECT 13.872 20.88 13.904 23.388 ;
  LAYER M1 ;
        RECT 13.936 20.88 13.968 23.388 ;
  LAYER M1 ;
        RECT 14 20.88 14.032 23.388 ;
  LAYER M1 ;
        RECT 14.064 20.88 14.096 23.388 ;
  LAYER M1 ;
        RECT 14.128 20.88 14.16 23.388 ;
  LAYER M1 ;
        RECT 14.192 20.88 14.224 23.388 ;
  LAYER M1 ;
        RECT 14.256 20.88 14.288 23.388 ;
  LAYER M1 ;
        RECT 14.32 20.88 14.352 23.388 ;
  LAYER M1 ;
        RECT 14.384 20.88 14.416 23.388 ;
  LAYER M1 ;
        RECT 14.448 20.88 14.48 23.388 ;
  LAYER M2 ;
        RECT 12.124 20.964 14.596 20.996 ;
  LAYER M2 ;
        RECT 12.124 21.028 14.596 21.06 ;
  LAYER M2 ;
        RECT 12.124 21.092 14.596 21.124 ;
  LAYER M2 ;
        RECT 12.124 21.156 14.596 21.188 ;
  LAYER M2 ;
        RECT 12.124 21.22 14.596 21.252 ;
  LAYER M2 ;
        RECT 12.124 21.284 14.596 21.316 ;
  LAYER M2 ;
        RECT 12.124 21.348 14.596 21.38 ;
  LAYER M2 ;
        RECT 12.124 21.412 14.596 21.444 ;
  LAYER M2 ;
        RECT 12.124 21.476 14.596 21.508 ;
  LAYER M2 ;
        RECT 12.124 21.54 14.596 21.572 ;
  LAYER M2 ;
        RECT 12.124 21.604 14.596 21.636 ;
  LAYER M2 ;
        RECT 12.124 21.668 14.596 21.7 ;
  LAYER M2 ;
        RECT 12.124 21.732 14.596 21.764 ;
  LAYER M2 ;
        RECT 12.124 21.796 14.596 21.828 ;
  LAYER M2 ;
        RECT 12.124 21.86 14.596 21.892 ;
  LAYER M2 ;
        RECT 12.124 21.924 14.596 21.956 ;
  LAYER M2 ;
        RECT 12.124 21.988 14.596 22.02 ;
  LAYER M2 ;
        RECT 12.124 22.052 14.596 22.084 ;
  LAYER M2 ;
        RECT 12.124 22.116 14.596 22.148 ;
  LAYER M2 ;
        RECT 12.124 22.18 14.596 22.212 ;
  LAYER M2 ;
        RECT 12.124 22.244 14.596 22.276 ;
  LAYER M2 ;
        RECT 12.124 22.308 14.596 22.34 ;
  LAYER M2 ;
        RECT 12.124 22.372 14.596 22.404 ;
  LAYER M2 ;
        RECT 12.124 22.436 14.596 22.468 ;
  LAYER M2 ;
        RECT 12.124 22.5 14.596 22.532 ;
  LAYER M2 ;
        RECT 12.124 22.564 14.596 22.596 ;
  LAYER M2 ;
        RECT 12.124 22.628 14.596 22.66 ;
  LAYER M2 ;
        RECT 12.124 22.692 14.596 22.724 ;
  LAYER M2 ;
        RECT 12.124 22.756 14.596 22.788 ;
  LAYER M2 ;
        RECT 12.124 22.82 14.596 22.852 ;
  LAYER M2 ;
        RECT 12.124 22.884 14.596 22.916 ;
  LAYER M2 ;
        RECT 12.124 22.948 14.596 22.98 ;
  LAYER M2 ;
        RECT 12.124 23.012 14.596 23.044 ;
  LAYER M2 ;
        RECT 12.124 23.076 14.596 23.108 ;
  LAYER M2 ;
        RECT 12.124 23.14 14.596 23.172 ;
  LAYER M2 ;
        RECT 12.124 23.204 14.596 23.236 ;
  LAYER M3 ;
        RECT 12.144 20.88 12.176 23.388 ;
  LAYER M3 ;
        RECT 12.208 20.88 12.24 23.388 ;
  LAYER M3 ;
        RECT 12.272 20.88 12.304 23.388 ;
  LAYER M3 ;
        RECT 12.336 20.88 12.368 23.388 ;
  LAYER M3 ;
        RECT 12.4 20.88 12.432 23.388 ;
  LAYER M3 ;
        RECT 12.464 20.88 12.496 23.388 ;
  LAYER M3 ;
        RECT 12.528 20.88 12.56 23.388 ;
  LAYER M3 ;
        RECT 12.592 20.88 12.624 23.388 ;
  LAYER M3 ;
        RECT 12.656 20.88 12.688 23.388 ;
  LAYER M3 ;
        RECT 12.72 20.88 12.752 23.388 ;
  LAYER M3 ;
        RECT 12.784 20.88 12.816 23.388 ;
  LAYER M3 ;
        RECT 12.848 20.88 12.88 23.388 ;
  LAYER M3 ;
        RECT 12.912 20.88 12.944 23.388 ;
  LAYER M3 ;
        RECT 12.976 20.88 13.008 23.388 ;
  LAYER M3 ;
        RECT 13.04 20.88 13.072 23.388 ;
  LAYER M3 ;
        RECT 13.104 20.88 13.136 23.388 ;
  LAYER M3 ;
        RECT 13.168 20.88 13.2 23.388 ;
  LAYER M3 ;
        RECT 13.232 20.88 13.264 23.388 ;
  LAYER M3 ;
        RECT 13.296 20.88 13.328 23.388 ;
  LAYER M3 ;
        RECT 13.36 20.88 13.392 23.388 ;
  LAYER M3 ;
        RECT 13.424 20.88 13.456 23.388 ;
  LAYER M3 ;
        RECT 13.488 20.88 13.52 23.388 ;
  LAYER M3 ;
        RECT 13.552 20.88 13.584 23.388 ;
  LAYER M3 ;
        RECT 13.616 20.88 13.648 23.388 ;
  LAYER M3 ;
        RECT 13.68 20.88 13.712 23.388 ;
  LAYER M3 ;
        RECT 13.744 20.88 13.776 23.388 ;
  LAYER M3 ;
        RECT 13.808 20.88 13.84 23.388 ;
  LAYER M3 ;
        RECT 13.872 20.88 13.904 23.388 ;
  LAYER M3 ;
        RECT 13.936 20.88 13.968 23.388 ;
  LAYER M3 ;
        RECT 14 20.88 14.032 23.388 ;
  LAYER M3 ;
        RECT 14.064 20.88 14.096 23.388 ;
  LAYER M3 ;
        RECT 14.128 20.88 14.16 23.388 ;
  LAYER M3 ;
        RECT 14.192 20.88 14.224 23.388 ;
  LAYER M3 ;
        RECT 14.256 20.88 14.288 23.388 ;
  LAYER M3 ;
        RECT 14.32 20.88 14.352 23.388 ;
  LAYER M3 ;
        RECT 14.384 20.88 14.416 23.388 ;
  LAYER M3 ;
        RECT 14.448 20.88 14.48 23.388 ;
  LAYER M3 ;
        RECT 14.544 20.88 14.576 23.388 ;
  LAYER M1 ;
        RECT 12.159 20.916 12.161 23.352 ;
  LAYER M1 ;
        RECT 12.239 20.916 12.241 23.352 ;
  LAYER M1 ;
        RECT 12.319 20.916 12.321 23.352 ;
  LAYER M1 ;
        RECT 12.399 20.916 12.401 23.352 ;
  LAYER M1 ;
        RECT 12.479 20.916 12.481 23.352 ;
  LAYER M1 ;
        RECT 12.559 20.916 12.561 23.352 ;
  LAYER M1 ;
        RECT 12.639 20.916 12.641 23.352 ;
  LAYER M1 ;
        RECT 12.719 20.916 12.721 23.352 ;
  LAYER M1 ;
        RECT 12.799 20.916 12.801 23.352 ;
  LAYER M1 ;
        RECT 12.879 20.916 12.881 23.352 ;
  LAYER M1 ;
        RECT 12.959 20.916 12.961 23.352 ;
  LAYER M1 ;
        RECT 13.039 20.916 13.041 23.352 ;
  LAYER M1 ;
        RECT 13.119 20.916 13.121 23.352 ;
  LAYER M1 ;
        RECT 13.199 20.916 13.201 23.352 ;
  LAYER M1 ;
        RECT 13.279 20.916 13.281 23.352 ;
  LAYER M1 ;
        RECT 13.359 20.916 13.361 23.352 ;
  LAYER M1 ;
        RECT 13.439 20.916 13.441 23.352 ;
  LAYER M1 ;
        RECT 13.519 20.916 13.521 23.352 ;
  LAYER M1 ;
        RECT 13.599 20.916 13.601 23.352 ;
  LAYER M1 ;
        RECT 13.679 20.916 13.681 23.352 ;
  LAYER M1 ;
        RECT 13.759 20.916 13.761 23.352 ;
  LAYER M1 ;
        RECT 13.839 20.916 13.841 23.352 ;
  LAYER M1 ;
        RECT 13.919 20.916 13.921 23.352 ;
  LAYER M1 ;
        RECT 13.999 20.916 14.001 23.352 ;
  LAYER M1 ;
        RECT 14.079 20.916 14.081 23.352 ;
  LAYER M1 ;
        RECT 14.159 20.916 14.161 23.352 ;
  LAYER M1 ;
        RECT 14.239 20.916 14.241 23.352 ;
  LAYER M1 ;
        RECT 14.319 20.916 14.321 23.352 ;
  LAYER M1 ;
        RECT 14.399 20.916 14.401 23.352 ;
  LAYER M1 ;
        RECT 14.479 20.916 14.481 23.352 ;
  LAYER M2 ;
        RECT 12.16 20.915 14.56 20.917 ;
  LAYER M2 ;
        RECT 12.16 20.999 14.56 21.001 ;
  LAYER M2 ;
        RECT 12.16 21.083 14.56 21.085 ;
  LAYER M2 ;
        RECT 12.16 21.167 14.56 21.169 ;
  LAYER M2 ;
        RECT 12.16 21.251 14.56 21.253 ;
  LAYER M2 ;
        RECT 12.16 21.335 14.56 21.337 ;
  LAYER M2 ;
        RECT 12.16 21.419 14.56 21.421 ;
  LAYER M2 ;
        RECT 12.16 21.503 14.56 21.505 ;
  LAYER M2 ;
        RECT 12.16 21.587 14.56 21.589 ;
  LAYER M2 ;
        RECT 12.16 21.671 14.56 21.673 ;
  LAYER M2 ;
        RECT 12.16 21.755 14.56 21.757 ;
  LAYER M2 ;
        RECT 12.16 21.839 14.56 21.841 ;
  LAYER M2 ;
        RECT 12.16 21.9225 14.56 21.9245 ;
  LAYER M2 ;
        RECT 12.16 22.007 14.56 22.009 ;
  LAYER M2 ;
        RECT 12.16 22.091 14.56 22.093 ;
  LAYER M2 ;
        RECT 12.16 22.175 14.56 22.177 ;
  LAYER M2 ;
        RECT 12.16 22.259 14.56 22.261 ;
  LAYER M2 ;
        RECT 12.16 22.343 14.56 22.345 ;
  LAYER M2 ;
        RECT 12.16 22.427 14.56 22.429 ;
  LAYER M2 ;
        RECT 12.16 22.511 14.56 22.513 ;
  LAYER M2 ;
        RECT 12.16 22.595 14.56 22.597 ;
  LAYER M2 ;
        RECT 12.16 22.679 14.56 22.681 ;
  LAYER M2 ;
        RECT 12.16 22.763 14.56 22.765 ;
  LAYER M2 ;
        RECT 12.16 22.847 14.56 22.849 ;
  LAYER M2 ;
        RECT 12.16 22.931 14.56 22.933 ;
  LAYER M2 ;
        RECT 12.16 23.015 14.56 23.017 ;
  LAYER M2 ;
        RECT 12.16 23.099 14.56 23.101 ;
  LAYER M2 ;
        RECT 12.16 23.183 14.56 23.185 ;
  LAYER M2 ;
        RECT 12.16 23.267 14.56 23.269 ;
  LAYER M1 ;
        RECT 12.144 23.82 12.176 26.328 ;
  LAYER M1 ;
        RECT 12.208 23.82 12.24 26.328 ;
  LAYER M1 ;
        RECT 12.272 23.82 12.304 26.328 ;
  LAYER M1 ;
        RECT 12.336 23.82 12.368 26.328 ;
  LAYER M1 ;
        RECT 12.4 23.82 12.432 26.328 ;
  LAYER M1 ;
        RECT 12.464 23.82 12.496 26.328 ;
  LAYER M1 ;
        RECT 12.528 23.82 12.56 26.328 ;
  LAYER M1 ;
        RECT 12.592 23.82 12.624 26.328 ;
  LAYER M1 ;
        RECT 12.656 23.82 12.688 26.328 ;
  LAYER M1 ;
        RECT 12.72 23.82 12.752 26.328 ;
  LAYER M1 ;
        RECT 12.784 23.82 12.816 26.328 ;
  LAYER M1 ;
        RECT 12.848 23.82 12.88 26.328 ;
  LAYER M1 ;
        RECT 12.912 23.82 12.944 26.328 ;
  LAYER M1 ;
        RECT 12.976 23.82 13.008 26.328 ;
  LAYER M1 ;
        RECT 13.04 23.82 13.072 26.328 ;
  LAYER M1 ;
        RECT 13.104 23.82 13.136 26.328 ;
  LAYER M1 ;
        RECT 13.168 23.82 13.2 26.328 ;
  LAYER M1 ;
        RECT 13.232 23.82 13.264 26.328 ;
  LAYER M1 ;
        RECT 13.296 23.82 13.328 26.328 ;
  LAYER M1 ;
        RECT 13.36 23.82 13.392 26.328 ;
  LAYER M1 ;
        RECT 13.424 23.82 13.456 26.328 ;
  LAYER M1 ;
        RECT 13.488 23.82 13.52 26.328 ;
  LAYER M1 ;
        RECT 13.552 23.82 13.584 26.328 ;
  LAYER M1 ;
        RECT 13.616 23.82 13.648 26.328 ;
  LAYER M1 ;
        RECT 13.68 23.82 13.712 26.328 ;
  LAYER M1 ;
        RECT 13.744 23.82 13.776 26.328 ;
  LAYER M1 ;
        RECT 13.808 23.82 13.84 26.328 ;
  LAYER M1 ;
        RECT 13.872 23.82 13.904 26.328 ;
  LAYER M1 ;
        RECT 13.936 23.82 13.968 26.328 ;
  LAYER M1 ;
        RECT 14 23.82 14.032 26.328 ;
  LAYER M1 ;
        RECT 14.064 23.82 14.096 26.328 ;
  LAYER M1 ;
        RECT 14.128 23.82 14.16 26.328 ;
  LAYER M1 ;
        RECT 14.192 23.82 14.224 26.328 ;
  LAYER M1 ;
        RECT 14.256 23.82 14.288 26.328 ;
  LAYER M1 ;
        RECT 14.32 23.82 14.352 26.328 ;
  LAYER M1 ;
        RECT 14.384 23.82 14.416 26.328 ;
  LAYER M1 ;
        RECT 14.448 23.82 14.48 26.328 ;
  LAYER M2 ;
        RECT 12.124 23.904 14.596 23.936 ;
  LAYER M2 ;
        RECT 12.124 23.968 14.596 24 ;
  LAYER M2 ;
        RECT 12.124 24.032 14.596 24.064 ;
  LAYER M2 ;
        RECT 12.124 24.096 14.596 24.128 ;
  LAYER M2 ;
        RECT 12.124 24.16 14.596 24.192 ;
  LAYER M2 ;
        RECT 12.124 24.224 14.596 24.256 ;
  LAYER M2 ;
        RECT 12.124 24.288 14.596 24.32 ;
  LAYER M2 ;
        RECT 12.124 24.352 14.596 24.384 ;
  LAYER M2 ;
        RECT 12.124 24.416 14.596 24.448 ;
  LAYER M2 ;
        RECT 12.124 24.48 14.596 24.512 ;
  LAYER M2 ;
        RECT 12.124 24.544 14.596 24.576 ;
  LAYER M2 ;
        RECT 12.124 24.608 14.596 24.64 ;
  LAYER M2 ;
        RECT 12.124 24.672 14.596 24.704 ;
  LAYER M2 ;
        RECT 12.124 24.736 14.596 24.768 ;
  LAYER M2 ;
        RECT 12.124 24.8 14.596 24.832 ;
  LAYER M2 ;
        RECT 12.124 24.864 14.596 24.896 ;
  LAYER M2 ;
        RECT 12.124 24.928 14.596 24.96 ;
  LAYER M2 ;
        RECT 12.124 24.992 14.596 25.024 ;
  LAYER M2 ;
        RECT 12.124 25.056 14.596 25.088 ;
  LAYER M2 ;
        RECT 12.124 25.12 14.596 25.152 ;
  LAYER M2 ;
        RECT 12.124 25.184 14.596 25.216 ;
  LAYER M2 ;
        RECT 12.124 25.248 14.596 25.28 ;
  LAYER M2 ;
        RECT 12.124 25.312 14.596 25.344 ;
  LAYER M2 ;
        RECT 12.124 25.376 14.596 25.408 ;
  LAYER M2 ;
        RECT 12.124 25.44 14.596 25.472 ;
  LAYER M2 ;
        RECT 12.124 25.504 14.596 25.536 ;
  LAYER M2 ;
        RECT 12.124 25.568 14.596 25.6 ;
  LAYER M2 ;
        RECT 12.124 25.632 14.596 25.664 ;
  LAYER M2 ;
        RECT 12.124 25.696 14.596 25.728 ;
  LAYER M2 ;
        RECT 12.124 25.76 14.596 25.792 ;
  LAYER M2 ;
        RECT 12.124 25.824 14.596 25.856 ;
  LAYER M2 ;
        RECT 12.124 25.888 14.596 25.92 ;
  LAYER M2 ;
        RECT 12.124 25.952 14.596 25.984 ;
  LAYER M2 ;
        RECT 12.124 26.016 14.596 26.048 ;
  LAYER M2 ;
        RECT 12.124 26.08 14.596 26.112 ;
  LAYER M2 ;
        RECT 12.124 26.144 14.596 26.176 ;
  LAYER M3 ;
        RECT 12.144 23.82 12.176 26.328 ;
  LAYER M3 ;
        RECT 12.208 23.82 12.24 26.328 ;
  LAYER M3 ;
        RECT 12.272 23.82 12.304 26.328 ;
  LAYER M3 ;
        RECT 12.336 23.82 12.368 26.328 ;
  LAYER M3 ;
        RECT 12.4 23.82 12.432 26.328 ;
  LAYER M3 ;
        RECT 12.464 23.82 12.496 26.328 ;
  LAYER M3 ;
        RECT 12.528 23.82 12.56 26.328 ;
  LAYER M3 ;
        RECT 12.592 23.82 12.624 26.328 ;
  LAYER M3 ;
        RECT 12.656 23.82 12.688 26.328 ;
  LAYER M3 ;
        RECT 12.72 23.82 12.752 26.328 ;
  LAYER M3 ;
        RECT 12.784 23.82 12.816 26.328 ;
  LAYER M3 ;
        RECT 12.848 23.82 12.88 26.328 ;
  LAYER M3 ;
        RECT 12.912 23.82 12.944 26.328 ;
  LAYER M3 ;
        RECT 12.976 23.82 13.008 26.328 ;
  LAYER M3 ;
        RECT 13.04 23.82 13.072 26.328 ;
  LAYER M3 ;
        RECT 13.104 23.82 13.136 26.328 ;
  LAYER M3 ;
        RECT 13.168 23.82 13.2 26.328 ;
  LAYER M3 ;
        RECT 13.232 23.82 13.264 26.328 ;
  LAYER M3 ;
        RECT 13.296 23.82 13.328 26.328 ;
  LAYER M3 ;
        RECT 13.36 23.82 13.392 26.328 ;
  LAYER M3 ;
        RECT 13.424 23.82 13.456 26.328 ;
  LAYER M3 ;
        RECT 13.488 23.82 13.52 26.328 ;
  LAYER M3 ;
        RECT 13.552 23.82 13.584 26.328 ;
  LAYER M3 ;
        RECT 13.616 23.82 13.648 26.328 ;
  LAYER M3 ;
        RECT 13.68 23.82 13.712 26.328 ;
  LAYER M3 ;
        RECT 13.744 23.82 13.776 26.328 ;
  LAYER M3 ;
        RECT 13.808 23.82 13.84 26.328 ;
  LAYER M3 ;
        RECT 13.872 23.82 13.904 26.328 ;
  LAYER M3 ;
        RECT 13.936 23.82 13.968 26.328 ;
  LAYER M3 ;
        RECT 14 23.82 14.032 26.328 ;
  LAYER M3 ;
        RECT 14.064 23.82 14.096 26.328 ;
  LAYER M3 ;
        RECT 14.128 23.82 14.16 26.328 ;
  LAYER M3 ;
        RECT 14.192 23.82 14.224 26.328 ;
  LAYER M3 ;
        RECT 14.256 23.82 14.288 26.328 ;
  LAYER M3 ;
        RECT 14.32 23.82 14.352 26.328 ;
  LAYER M3 ;
        RECT 14.384 23.82 14.416 26.328 ;
  LAYER M3 ;
        RECT 14.448 23.82 14.48 26.328 ;
  LAYER M3 ;
        RECT 14.544 23.82 14.576 26.328 ;
  LAYER M1 ;
        RECT 12.159 23.856 12.161 26.292 ;
  LAYER M1 ;
        RECT 12.239 23.856 12.241 26.292 ;
  LAYER M1 ;
        RECT 12.319 23.856 12.321 26.292 ;
  LAYER M1 ;
        RECT 12.399 23.856 12.401 26.292 ;
  LAYER M1 ;
        RECT 12.479 23.856 12.481 26.292 ;
  LAYER M1 ;
        RECT 12.559 23.856 12.561 26.292 ;
  LAYER M1 ;
        RECT 12.639 23.856 12.641 26.292 ;
  LAYER M1 ;
        RECT 12.719 23.856 12.721 26.292 ;
  LAYER M1 ;
        RECT 12.799 23.856 12.801 26.292 ;
  LAYER M1 ;
        RECT 12.879 23.856 12.881 26.292 ;
  LAYER M1 ;
        RECT 12.959 23.856 12.961 26.292 ;
  LAYER M1 ;
        RECT 13.039 23.856 13.041 26.292 ;
  LAYER M1 ;
        RECT 13.119 23.856 13.121 26.292 ;
  LAYER M1 ;
        RECT 13.199 23.856 13.201 26.292 ;
  LAYER M1 ;
        RECT 13.279 23.856 13.281 26.292 ;
  LAYER M1 ;
        RECT 13.359 23.856 13.361 26.292 ;
  LAYER M1 ;
        RECT 13.439 23.856 13.441 26.292 ;
  LAYER M1 ;
        RECT 13.519 23.856 13.521 26.292 ;
  LAYER M1 ;
        RECT 13.599 23.856 13.601 26.292 ;
  LAYER M1 ;
        RECT 13.679 23.856 13.681 26.292 ;
  LAYER M1 ;
        RECT 13.759 23.856 13.761 26.292 ;
  LAYER M1 ;
        RECT 13.839 23.856 13.841 26.292 ;
  LAYER M1 ;
        RECT 13.919 23.856 13.921 26.292 ;
  LAYER M1 ;
        RECT 13.999 23.856 14.001 26.292 ;
  LAYER M1 ;
        RECT 14.079 23.856 14.081 26.292 ;
  LAYER M1 ;
        RECT 14.159 23.856 14.161 26.292 ;
  LAYER M1 ;
        RECT 14.239 23.856 14.241 26.292 ;
  LAYER M1 ;
        RECT 14.319 23.856 14.321 26.292 ;
  LAYER M1 ;
        RECT 14.399 23.856 14.401 26.292 ;
  LAYER M1 ;
        RECT 14.479 23.856 14.481 26.292 ;
  LAYER M2 ;
        RECT 12.16 23.855 14.56 23.857 ;
  LAYER M2 ;
        RECT 12.16 23.939 14.56 23.941 ;
  LAYER M2 ;
        RECT 12.16 24.023 14.56 24.025 ;
  LAYER M2 ;
        RECT 12.16 24.107 14.56 24.109 ;
  LAYER M2 ;
        RECT 12.16 24.191 14.56 24.193 ;
  LAYER M2 ;
        RECT 12.16 24.275 14.56 24.277 ;
  LAYER M2 ;
        RECT 12.16 24.359 14.56 24.361 ;
  LAYER M2 ;
        RECT 12.16 24.443 14.56 24.445 ;
  LAYER M2 ;
        RECT 12.16 24.527 14.56 24.529 ;
  LAYER M2 ;
        RECT 12.16 24.611 14.56 24.613 ;
  LAYER M2 ;
        RECT 12.16 24.695 14.56 24.697 ;
  LAYER M2 ;
        RECT 12.16 24.779 14.56 24.781 ;
  LAYER M2 ;
        RECT 12.16 24.8625 14.56 24.8645 ;
  LAYER M2 ;
        RECT 12.16 24.947 14.56 24.949 ;
  LAYER M2 ;
        RECT 12.16 25.031 14.56 25.033 ;
  LAYER M2 ;
        RECT 12.16 25.115 14.56 25.117 ;
  LAYER M2 ;
        RECT 12.16 25.199 14.56 25.201 ;
  LAYER M2 ;
        RECT 12.16 25.283 14.56 25.285 ;
  LAYER M2 ;
        RECT 12.16 25.367 14.56 25.369 ;
  LAYER M2 ;
        RECT 12.16 25.451 14.56 25.453 ;
  LAYER M2 ;
        RECT 12.16 25.535 14.56 25.537 ;
  LAYER M2 ;
        RECT 12.16 25.619 14.56 25.621 ;
  LAYER M2 ;
        RECT 12.16 25.703 14.56 25.705 ;
  LAYER M2 ;
        RECT 12.16 25.787 14.56 25.789 ;
  LAYER M2 ;
        RECT 12.16 25.871 14.56 25.873 ;
  LAYER M2 ;
        RECT 12.16 25.955 14.56 25.957 ;
  LAYER M2 ;
        RECT 12.16 26.039 14.56 26.041 ;
  LAYER M2 ;
        RECT 12.16 26.123 14.56 26.125 ;
  LAYER M2 ;
        RECT 12.16 26.207 14.56 26.209 ;
  LAYER M1 ;
        RECT 12.144 26.76 12.176 29.268 ;
  LAYER M1 ;
        RECT 12.208 26.76 12.24 29.268 ;
  LAYER M1 ;
        RECT 12.272 26.76 12.304 29.268 ;
  LAYER M1 ;
        RECT 12.336 26.76 12.368 29.268 ;
  LAYER M1 ;
        RECT 12.4 26.76 12.432 29.268 ;
  LAYER M1 ;
        RECT 12.464 26.76 12.496 29.268 ;
  LAYER M1 ;
        RECT 12.528 26.76 12.56 29.268 ;
  LAYER M1 ;
        RECT 12.592 26.76 12.624 29.268 ;
  LAYER M1 ;
        RECT 12.656 26.76 12.688 29.268 ;
  LAYER M1 ;
        RECT 12.72 26.76 12.752 29.268 ;
  LAYER M1 ;
        RECT 12.784 26.76 12.816 29.268 ;
  LAYER M1 ;
        RECT 12.848 26.76 12.88 29.268 ;
  LAYER M1 ;
        RECT 12.912 26.76 12.944 29.268 ;
  LAYER M1 ;
        RECT 12.976 26.76 13.008 29.268 ;
  LAYER M1 ;
        RECT 13.04 26.76 13.072 29.268 ;
  LAYER M1 ;
        RECT 13.104 26.76 13.136 29.268 ;
  LAYER M1 ;
        RECT 13.168 26.76 13.2 29.268 ;
  LAYER M1 ;
        RECT 13.232 26.76 13.264 29.268 ;
  LAYER M1 ;
        RECT 13.296 26.76 13.328 29.268 ;
  LAYER M1 ;
        RECT 13.36 26.76 13.392 29.268 ;
  LAYER M1 ;
        RECT 13.424 26.76 13.456 29.268 ;
  LAYER M1 ;
        RECT 13.488 26.76 13.52 29.268 ;
  LAYER M1 ;
        RECT 13.552 26.76 13.584 29.268 ;
  LAYER M1 ;
        RECT 13.616 26.76 13.648 29.268 ;
  LAYER M1 ;
        RECT 13.68 26.76 13.712 29.268 ;
  LAYER M1 ;
        RECT 13.744 26.76 13.776 29.268 ;
  LAYER M1 ;
        RECT 13.808 26.76 13.84 29.268 ;
  LAYER M1 ;
        RECT 13.872 26.76 13.904 29.268 ;
  LAYER M1 ;
        RECT 13.936 26.76 13.968 29.268 ;
  LAYER M1 ;
        RECT 14 26.76 14.032 29.268 ;
  LAYER M1 ;
        RECT 14.064 26.76 14.096 29.268 ;
  LAYER M1 ;
        RECT 14.128 26.76 14.16 29.268 ;
  LAYER M1 ;
        RECT 14.192 26.76 14.224 29.268 ;
  LAYER M1 ;
        RECT 14.256 26.76 14.288 29.268 ;
  LAYER M1 ;
        RECT 14.32 26.76 14.352 29.268 ;
  LAYER M1 ;
        RECT 14.384 26.76 14.416 29.268 ;
  LAYER M1 ;
        RECT 14.448 26.76 14.48 29.268 ;
  LAYER M2 ;
        RECT 12.124 26.844 14.596 26.876 ;
  LAYER M2 ;
        RECT 12.124 26.908 14.596 26.94 ;
  LAYER M2 ;
        RECT 12.124 26.972 14.596 27.004 ;
  LAYER M2 ;
        RECT 12.124 27.036 14.596 27.068 ;
  LAYER M2 ;
        RECT 12.124 27.1 14.596 27.132 ;
  LAYER M2 ;
        RECT 12.124 27.164 14.596 27.196 ;
  LAYER M2 ;
        RECT 12.124 27.228 14.596 27.26 ;
  LAYER M2 ;
        RECT 12.124 27.292 14.596 27.324 ;
  LAYER M2 ;
        RECT 12.124 27.356 14.596 27.388 ;
  LAYER M2 ;
        RECT 12.124 27.42 14.596 27.452 ;
  LAYER M2 ;
        RECT 12.124 27.484 14.596 27.516 ;
  LAYER M2 ;
        RECT 12.124 27.548 14.596 27.58 ;
  LAYER M2 ;
        RECT 12.124 27.612 14.596 27.644 ;
  LAYER M2 ;
        RECT 12.124 27.676 14.596 27.708 ;
  LAYER M2 ;
        RECT 12.124 27.74 14.596 27.772 ;
  LAYER M2 ;
        RECT 12.124 27.804 14.596 27.836 ;
  LAYER M2 ;
        RECT 12.124 27.868 14.596 27.9 ;
  LAYER M2 ;
        RECT 12.124 27.932 14.596 27.964 ;
  LAYER M2 ;
        RECT 12.124 27.996 14.596 28.028 ;
  LAYER M2 ;
        RECT 12.124 28.06 14.596 28.092 ;
  LAYER M2 ;
        RECT 12.124 28.124 14.596 28.156 ;
  LAYER M2 ;
        RECT 12.124 28.188 14.596 28.22 ;
  LAYER M2 ;
        RECT 12.124 28.252 14.596 28.284 ;
  LAYER M2 ;
        RECT 12.124 28.316 14.596 28.348 ;
  LAYER M2 ;
        RECT 12.124 28.38 14.596 28.412 ;
  LAYER M2 ;
        RECT 12.124 28.444 14.596 28.476 ;
  LAYER M2 ;
        RECT 12.124 28.508 14.596 28.54 ;
  LAYER M2 ;
        RECT 12.124 28.572 14.596 28.604 ;
  LAYER M2 ;
        RECT 12.124 28.636 14.596 28.668 ;
  LAYER M2 ;
        RECT 12.124 28.7 14.596 28.732 ;
  LAYER M2 ;
        RECT 12.124 28.764 14.596 28.796 ;
  LAYER M2 ;
        RECT 12.124 28.828 14.596 28.86 ;
  LAYER M2 ;
        RECT 12.124 28.892 14.596 28.924 ;
  LAYER M2 ;
        RECT 12.124 28.956 14.596 28.988 ;
  LAYER M2 ;
        RECT 12.124 29.02 14.596 29.052 ;
  LAYER M2 ;
        RECT 12.124 29.084 14.596 29.116 ;
  LAYER M3 ;
        RECT 12.144 26.76 12.176 29.268 ;
  LAYER M3 ;
        RECT 12.208 26.76 12.24 29.268 ;
  LAYER M3 ;
        RECT 12.272 26.76 12.304 29.268 ;
  LAYER M3 ;
        RECT 12.336 26.76 12.368 29.268 ;
  LAYER M3 ;
        RECT 12.4 26.76 12.432 29.268 ;
  LAYER M3 ;
        RECT 12.464 26.76 12.496 29.268 ;
  LAYER M3 ;
        RECT 12.528 26.76 12.56 29.268 ;
  LAYER M3 ;
        RECT 12.592 26.76 12.624 29.268 ;
  LAYER M3 ;
        RECT 12.656 26.76 12.688 29.268 ;
  LAYER M3 ;
        RECT 12.72 26.76 12.752 29.268 ;
  LAYER M3 ;
        RECT 12.784 26.76 12.816 29.268 ;
  LAYER M3 ;
        RECT 12.848 26.76 12.88 29.268 ;
  LAYER M3 ;
        RECT 12.912 26.76 12.944 29.268 ;
  LAYER M3 ;
        RECT 12.976 26.76 13.008 29.268 ;
  LAYER M3 ;
        RECT 13.04 26.76 13.072 29.268 ;
  LAYER M3 ;
        RECT 13.104 26.76 13.136 29.268 ;
  LAYER M3 ;
        RECT 13.168 26.76 13.2 29.268 ;
  LAYER M3 ;
        RECT 13.232 26.76 13.264 29.268 ;
  LAYER M3 ;
        RECT 13.296 26.76 13.328 29.268 ;
  LAYER M3 ;
        RECT 13.36 26.76 13.392 29.268 ;
  LAYER M3 ;
        RECT 13.424 26.76 13.456 29.268 ;
  LAYER M3 ;
        RECT 13.488 26.76 13.52 29.268 ;
  LAYER M3 ;
        RECT 13.552 26.76 13.584 29.268 ;
  LAYER M3 ;
        RECT 13.616 26.76 13.648 29.268 ;
  LAYER M3 ;
        RECT 13.68 26.76 13.712 29.268 ;
  LAYER M3 ;
        RECT 13.744 26.76 13.776 29.268 ;
  LAYER M3 ;
        RECT 13.808 26.76 13.84 29.268 ;
  LAYER M3 ;
        RECT 13.872 26.76 13.904 29.268 ;
  LAYER M3 ;
        RECT 13.936 26.76 13.968 29.268 ;
  LAYER M3 ;
        RECT 14 26.76 14.032 29.268 ;
  LAYER M3 ;
        RECT 14.064 26.76 14.096 29.268 ;
  LAYER M3 ;
        RECT 14.128 26.76 14.16 29.268 ;
  LAYER M3 ;
        RECT 14.192 26.76 14.224 29.268 ;
  LAYER M3 ;
        RECT 14.256 26.76 14.288 29.268 ;
  LAYER M3 ;
        RECT 14.32 26.76 14.352 29.268 ;
  LAYER M3 ;
        RECT 14.384 26.76 14.416 29.268 ;
  LAYER M3 ;
        RECT 14.448 26.76 14.48 29.268 ;
  LAYER M3 ;
        RECT 14.544 26.76 14.576 29.268 ;
  LAYER M1 ;
        RECT 12.159 26.796 12.161 29.232 ;
  LAYER M1 ;
        RECT 12.239 26.796 12.241 29.232 ;
  LAYER M1 ;
        RECT 12.319 26.796 12.321 29.232 ;
  LAYER M1 ;
        RECT 12.399 26.796 12.401 29.232 ;
  LAYER M1 ;
        RECT 12.479 26.796 12.481 29.232 ;
  LAYER M1 ;
        RECT 12.559 26.796 12.561 29.232 ;
  LAYER M1 ;
        RECT 12.639 26.796 12.641 29.232 ;
  LAYER M1 ;
        RECT 12.719 26.796 12.721 29.232 ;
  LAYER M1 ;
        RECT 12.799 26.796 12.801 29.232 ;
  LAYER M1 ;
        RECT 12.879 26.796 12.881 29.232 ;
  LAYER M1 ;
        RECT 12.959 26.796 12.961 29.232 ;
  LAYER M1 ;
        RECT 13.039 26.796 13.041 29.232 ;
  LAYER M1 ;
        RECT 13.119 26.796 13.121 29.232 ;
  LAYER M1 ;
        RECT 13.199 26.796 13.201 29.232 ;
  LAYER M1 ;
        RECT 13.279 26.796 13.281 29.232 ;
  LAYER M1 ;
        RECT 13.359 26.796 13.361 29.232 ;
  LAYER M1 ;
        RECT 13.439 26.796 13.441 29.232 ;
  LAYER M1 ;
        RECT 13.519 26.796 13.521 29.232 ;
  LAYER M1 ;
        RECT 13.599 26.796 13.601 29.232 ;
  LAYER M1 ;
        RECT 13.679 26.796 13.681 29.232 ;
  LAYER M1 ;
        RECT 13.759 26.796 13.761 29.232 ;
  LAYER M1 ;
        RECT 13.839 26.796 13.841 29.232 ;
  LAYER M1 ;
        RECT 13.919 26.796 13.921 29.232 ;
  LAYER M1 ;
        RECT 13.999 26.796 14.001 29.232 ;
  LAYER M1 ;
        RECT 14.079 26.796 14.081 29.232 ;
  LAYER M1 ;
        RECT 14.159 26.796 14.161 29.232 ;
  LAYER M1 ;
        RECT 14.239 26.796 14.241 29.232 ;
  LAYER M1 ;
        RECT 14.319 26.796 14.321 29.232 ;
  LAYER M1 ;
        RECT 14.399 26.796 14.401 29.232 ;
  LAYER M1 ;
        RECT 14.479 26.796 14.481 29.232 ;
  LAYER M2 ;
        RECT 12.16 26.795 14.56 26.797 ;
  LAYER M2 ;
        RECT 12.16 26.879 14.56 26.881 ;
  LAYER M2 ;
        RECT 12.16 26.963 14.56 26.965 ;
  LAYER M2 ;
        RECT 12.16 27.047 14.56 27.049 ;
  LAYER M2 ;
        RECT 12.16 27.131 14.56 27.133 ;
  LAYER M2 ;
        RECT 12.16 27.215 14.56 27.217 ;
  LAYER M2 ;
        RECT 12.16 27.299 14.56 27.301 ;
  LAYER M2 ;
        RECT 12.16 27.383 14.56 27.385 ;
  LAYER M2 ;
        RECT 12.16 27.467 14.56 27.469 ;
  LAYER M2 ;
        RECT 12.16 27.551 14.56 27.553 ;
  LAYER M2 ;
        RECT 12.16 27.635 14.56 27.637 ;
  LAYER M2 ;
        RECT 12.16 27.719 14.56 27.721 ;
  LAYER M2 ;
        RECT 12.16 27.8025 14.56 27.8045 ;
  LAYER M2 ;
        RECT 12.16 27.887 14.56 27.889 ;
  LAYER M2 ;
        RECT 12.16 27.971 14.56 27.973 ;
  LAYER M2 ;
        RECT 12.16 28.055 14.56 28.057 ;
  LAYER M2 ;
        RECT 12.16 28.139 14.56 28.141 ;
  LAYER M2 ;
        RECT 12.16 28.223 14.56 28.225 ;
  LAYER M2 ;
        RECT 12.16 28.307 14.56 28.309 ;
  LAYER M2 ;
        RECT 12.16 28.391 14.56 28.393 ;
  LAYER M2 ;
        RECT 12.16 28.475 14.56 28.477 ;
  LAYER M2 ;
        RECT 12.16 28.559 14.56 28.561 ;
  LAYER M2 ;
        RECT 12.16 28.643 14.56 28.645 ;
  LAYER M2 ;
        RECT 12.16 28.727 14.56 28.729 ;
  LAYER M2 ;
        RECT 12.16 28.811 14.56 28.813 ;
  LAYER M2 ;
        RECT 12.16 28.895 14.56 28.897 ;
  LAYER M2 ;
        RECT 12.16 28.979 14.56 28.981 ;
  LAYER M2 ;
        RECT 12.16 29.063 14.56 29.065 ;
  LAYER M2 ;
        RECT 12.16 29.147 14.56 29.149 ;
  LAYER M1 ;
        RECT 5.104 0.3 5.136 0.96 ;
  LAYER M1 ;
        RECT 5.024 0.3 5.056 0.96 ;
  LAYER M1 ;
        RECT 5.184 0.3 5.216 0.96 ;
  LAYER M2 ;
        RECT 4.924 0.908 5.236 0.94 ;
  LAYER M2 ;
        RECT 4.924 0.656 5.236 0.688 ;
  LAYER M2 ;
        RECT 5.004 0.824 5.316 0.856 ;
  LAYER M2 ;
        RECT 5.004 0.572 5.316 0.604 ;
  LAYER M2 ;
        RECT 5.004 0.74 5.396 0.772 ;
  LAYER M2 ;
        RECT 5.004 0.488 5.396 0.52 ;
  LAYER M1 ;
        RECT 15.184 17.352 15.216 18.012 ;
  LAYER M1 ;
        RECT 15.104 17.352 15.136 18.012 ;
  LAYER M1 ;
        RECT 15.264 17.352 15.296 18.012 ;
  LAYER M2 ;
        RECT 15.004 17.96 15.316 17.992 ;
  LAYER M2 ;
        RECT 15.004 17.708 15.316 17.74 ;
  LAYER M2 ;
        RECT 15.084 17.876 15.396 17.908 ;
  LAYER M2 ;
        RECT 15.084 17.624 15.396 17.656 ;
  LAYER M2 ;
        RECT 15.084 17.792 15.476 17.824 ;
  LAYER M2 ;
        RECT 15.084 17.54 15.476 17.572 ;
  LAYER M1 ;
        RECT 6.464 0.3 6.496 0.96 ;
  LAYER M1 ;
        RECT 6.544 0.3 6.576 0.96 ;
  LAYER M1 ;
        RECT 6.384 0.3 6.416 0.96 ;
  LAYER M1 ;
        RECT 5.824 0.3 5.856 0.96 ;
  LAYER M1 ;
        RECT 5.904 0.3 5.936 0.96 ;
  LAYER M1 ;
        RECT 5.744 0.3 5.776 0.96 ;
  LAYER M1 ;
        RECT 7.184 0.3 7.216 0.96 ;
  LAYER M1 ;
        RECT 7.104 0.3 7.136 0.96 ;
  LAYER M1 ;
        RECT 7.264 0.3 7.296 0.96 ;
  LAYER M1 ;
        RECT 7.824 0.3 7.856 0.96 ;
  LAYER M1 ;
        RECT 7.744 0.3 7.776 0.96 ;
  LAYER M1 ;
        RECT 7.904 0.3 7.936 0.96 ;
  LAYER M1 ;
        RECT 8.704 10.296 8.736 10.368 ;
  LAYER M2 ;
        RECT 8.684 10.316 8.756 10.348 ;
  LAYER M2 ;
        RECT 8.72 10.316 9.04 10.348 ;
  LAYER M1 ;
        RECT 9.024 10.296 9.056 10.368 ;
  LAYER M2 ;
        RECT 9.004 10.316 9.076 10.348 ;
  LAYER M1 ;
        RECT 11.584 7.356 11.616 7.428 ;
  LAYER M2 ;
        RECT 11.564 7.376 11.636 7.408 ;
  LAYER M1 ;
        RECT 11.584 7.392 11.616 7.56 ;
  LAYER M1 ;
        RECT 11.584 7.524 11.616 7.596 ;
  LAYER M2 ;
        RECT 11.564 7.544 11.636 7.576 ;
  LAYER M2 ;
        RECT 9.04 7.544 11.6 7.576 ;
  LAYER M1 ;
        RECT 9.024 7.524 9.056 7.596 ;
  LAYER M2 ;
        RECT 9.004 7.544 9.076 7.576 ;
  LAYER M1 ;
        RECT 9.024 16.68 9.056 16.752 ;
  LAYER M2 ;
        RECT 9.004 16.7 9.076 16.732 ;
  LAYER M1 ;
        RECT 9.024 16.548 9.056 16.716 ;
  LAYER M1 ;
        RECT 9.024 7.56 9.056 16.548 ;
  LAYER M1 ;
        RECT 5.824 13.236 5.856 13.308 ;
  LAYER M2 ;
        RECT 5.804 13.256 5.876 13.288 ;
  LAYER M2 ;
        RECT 5.84 13.256 6.16 13.288 ;
  LAYER M1 ;
        RECT 6.144 13.236 6.176 13.308 ;
  LAYER M2 ;
        RECT 6.124 13.256 6.196 13.288 ;
  LAYER M1 ;
        RECT 6.144 16.68 6.176 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.7 6.196 16.732 ;
  LAYER M1 ;
        RECT 6.144 16.548 6.176 16.716 ;
  LAYER M1 ;
        RECT 6.144 13.272 6.176 16.548 ;
  LAYER M2 ;
        RECT 6.16 16.7 9.04 16.732 ;
  LAYER M1 ;
        RECT 11.584 10.296 11.616 10.368 ;
  LAYER M2 ;
        RECT 11.564 10.316 11.636 10.348 ;
  LAYER M2 ;
        RECT 11.6 10.316 11.92 10.348 ;
  LAYER M1 ;
        RECT 11.904 10.296 11.936 10.368 ;
  LAYER M2 ;
        RECT 11.884 10.316 11.956 10.348 ;
  LAYER M1 ;
        RECT 11.584 13.236 11.616 13.308 ;
  LAYER M2 ;
        RECT 11.564 13.256 11.636 13.288 ;
  LAYER M2 ;
        RECT 11.6 13.256 11.92 13.288 ;
  LAYER M1 ;
        RECT 11.904 13.236 11.936 13.308 ;
  LAYER M2 ;
        RECT 11.884 13.256 11.956 13.288 ;
  LAYER M1 ;
        RECT 11.904 16.848 11.936 16.92 ;
  LAYER M2 ;
        RECT 11.884 16.868 11.956 16.9 ;
  LAYER M1 ;
        RECT 11.904 16.548 11.936 16.884 ;
  LAYER M1 ;
        RECT 11.904 10.332 11.936 16.548 ;
  LAYER M1 ;
        RECT 5.824 10.296 5.856 10.368 ;
  LAYER M2 ;
        RECT 5.804 10.316 5.876 10.348 ;
  LAYER M1 ;
        RECT 5.824 10.332 5.856 10.5 ;
  LAYER M1 ;
        RECT 5.824 10.464 5.856 10.536 ;
  LAYER M2 ;
        RECT 5.804 10.484 5.876 10.516 ;
  LAYER M2 ;
        RECT 3.28 10.484 5.84 10.516 ;
  LAYER M1 ;
        RECT 3.264 10.464 3.296 10.536 ;
  LAYER M2 ;
        RECT 3.244 10.484 3.316 10.516 ;
  LAYER M1 ;
        RECT 5.824 7.356 5.856 7.428 ;
  LAYER M2 ;
        RECT 5.804 7.376 5.876 7.408 ;
  LAYER M1 ;
        RECT 5.824 7.392 5.856 7.56 ;
  LAYER M1 ;
        RECT 5.824 7.524 5.856 7.596 ;
  LAYER M2 ;
        RECT 5.804 7.544 5.876 7.576 ;
  LAYER M2 ;
        RECT 3.28 7.544 5.84 7.576 ;
  LAYER M1 ;
        RECT 3.264 7.524 3.296 7.596 ;
  LAYER M2 ;
        RECT 3.244 7.544 3.316 7.576 ;
  LAYER M1 ;
        RECT 3.264 16.848 3.296 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.868 3.316 16.9 ;
  LAYER M1 ;
        RECT 3.264 16.548 3.296 16.884 ;
  LAYER M1 ;
        RECT 3.264 7.56 3.296 16.548 ;
  LAYER M2 ;
        RECT 3.28 16.868 11.92 16.9 ;
  LAYER M1 ;
        RECT 8.704 13.236 8.736 13.308 ;
  LAYER M2 ;
        RECT 8.684 13.256 8.756 13.288 ;
  LAYER M2 ;
        RECT 8.72 13.256 11.6 13.288 ;
  LAYER M1 ;
        RECT 11.584 13.236 11.616 13.308 ;
  LAYER M2 ;
        RECT 11.564 13.256 11.636 13.288 ;
  LAYER M1 ;
        RECT 8.704 7.356 8.736 7.428 ;
  LAYER M2 ;
        RECT 8.684 7.376 8.756 7.408 ;
  LAYER M2 ;
        RECT 5.84 7.376 8.72 7.408 ;
  LAYER M1 ;
        RECT 5.824 7.356 5.856 7.428 ;
  LAYER M2 ;
        RECT 5.804 7.376 5.876 7.408 ;
  LAYER M1 ;
        RECT 14.464 16.176 14.496 16.248 ;
  LAYER M2 ;
        RECT 14.444 16.196 14.516 16.228 ;
  LAYER M2 ;
        RECT 14.48 16.196 14.8 16.228 ;
  LAYER M1 ;
        RECT 14.784 16.176 14.816 16.248 ;
  LAYER M2 ;
        RECT 14.764 16.196 14.836 16.228 ;
  LAYER M1 ;
        RECT 14.464 13.236 14.496 13.308 ;
  LAYER M2 ;
        RECT 14.444 13.256 14.516 13.288 ;
  LAYER M2 ;
        RECT 14.48 13.256 14.8 13.288 ;
  LAYER M1 ;
        RECT 14.784 13.236 14.816 13.308 ;
  LAYER M2 ;
        RECT 14.764 13.256 14.836 13.288 ;
  LAYER M1 ;
        RECT 14.464 10.296 14.496 10.368 ;
  LAYER M2 ;
        RECT 14.444 10.316 14.516 10.348 ;
  LAYER M2 ;
        RECT 14.48 10.316 14.8 10.348 ;
  LAYER M1 ;
        RECT 14.784 10.296 14.816 10.368 ;
  LAYER M2 ;
        RECT 14.764 10.316 14.836 10.348 ;
  LAYER M1 ;
        RECT 14.464 7.356 14.496 7.428 ;
  LAYER M2 ;
        RECT 14.444 7.376 14.516 7.408 ;
  LAYER M2 ;
        RECT 14.48 7.376 14.8 7.408 ;
  LAYER M1 ;
        RECT 14.784 7.356 14.816 7.428 ;
  LAYER M2 ;
        RECT 14.764 7.376 14.836 7.408 ;
  LAYER M1 ;
        RECT 14.464 4.416 14.496 4.488 ;
  LAYER M2 ;
        RECT 14.444 4.436 14.516 4.468 ;
  LAYER M2 ;
        RECT 14.48 4.436 14.8 4.468 ;
  LAYER M1 ;
        RECT 14.784 4.416 14.816 4.488 ;
  LAYER M2 ;
        RECT 14.764 4.436 14.836 4.468 ;
  LAYER M1 ;
        RECT 14.784 17.016 14.816 17.088 ;
  LAYER M2 ;
        RECT 14.764 17.036 14.836 17.068 ;
  LAYER M1 ;
        RECT 14.784 16.548 14.816 17.052 ;
  LAYER M1 ;
        RECT 14.784 4.452 14.816 16.548 ;
  LAYER M1 ;
        RECT 2.944 16.176 2.976 16.248 ;
  LAYER M2 ;
        RECT 2.924 16.196 2.996 16.228 ;
  LAYER M1 ;
        RECT 2.944 16.212 2.976 16.38 ;
  LAYER M1 ;
        RECT 2.944 16.344 2.976 16.416 ;
  LAYER M2 ;
        RECT 2.924 16.364 2.996 16.396 ;
  LAYER M2 ;
        RECT 0.4 16.364 2.96 16.396 ;
  LAYER M1 ;
        RECT 0.384 16.344 0.416 16.416 ;
  LAYER M2 ;
        RECT 0.364 16.364 0.436 16.396 ;
  LAYER M1 ;
        RECT 2.944 13.236 2.976 13.308 ;
  LAYER M2 ;
        RECT 2.924 13.256 2.996 13.288 ;
  LAYER M1 ;
        RECT 2.944 13.272 2.976 13.44 ;
  LAYER M1 ;
        RECT 2.944 13.404 2.976 13.476 ;
  LAYER M2 ;
        RECT 2.924 13.424 2.996 13.456 ;
  LAYER M2 ;
        RECT 0.4 13.424 2.96 13.456 ;
  LAYER M1 ;
        RECT 0.384 13.404 0.416 13.476 ;
  LAYER M2 ;
        RECT 0.364 13.424 0.436 13.456 ;
  LAYER M1 ;
        RECT 2.944 10.296 2.976 10.368 ;
  LAYER M2 ;
        RECT 2.924 10.316 2.996 10.348 ;
  LAYER M1 ;
        RECT 2.944 10.332 2.976 10.5 ;
  LAYER M1 ;
        RECT 2.944 10.464 2.976 10.536 ;
  LAYER M2 ;
        RECT 2.924 10.484 2.996 10.516 ;
  LAYER M2 ;
        RECT 0.4 10.484 2.96 10.516 ;
  LAYER M1 ;
        RECT 0.384 10.464 0.416 10.536 ;
  LAYER M2 ;
        RECT 0.364 10.484 0.436 10.516 ;
  LAYER M1 ;
        RECT 2.944 7.356 2.976 7.428 ;
  LAYER M2 ;
        RECT 2.924 7.376 2.996 7.408 ;
  LAYER M1 ;
        RECT 2.944 7.392 2.976 7.56 ;
  LAYER M1 ;
        RECT 2.944 7.524 2.976 7.596 ;
  LAYER M2 ;
        RECT 2.924 7.544 2.996 7.576 ;
  LAYER M2 ;
        RECT 0.4 7.544 2.96 7.576 ;
  LAYER M1 ;
        RECT 0.384 7.524 0.416 7.596 ;
  LAYER M2 ;
        RECT 0.364 7.544 0.436 7.576 ;
  LAYER M1 ;
        RECT 2.944 4.416 2.976 4.488 ;
  LAYER M2 ;
        RECT 2.924 4.436 2.996 4.468 ;
  LAYER M1 ;
        RECT 2.944 4.452 2.976 4.62 ;
  LAYER M1 ;
        RECT 2.944 4.584 2.976 4.656 ;
  LAYER M2 ;
        RECT 2.924 4.604 2.996 4.636 ;
  LAYER M2 ;
        RECT 0.4 4.604 2.96 4.636 ;
  LAYER M1 ;
        RECT 0.384 4.584 0.416 4.656 ;
  LAYER M2 ;
        RECT 0.364 4.604 0.436 4.636 ;
  LAYER M1 ;
        RECT 0.384 17.016 0.416 17.088 ;
  LAYER M2 ;
        RECT 0.364 17.036 0.436 17.068 ;
  LAYER M1 ;
        RECT 0.384 16.548 0.416 17.052 ;
  LAYER M1 ;
        RECT 0.384 4.62 0.416 16.548 ;
  LAYER M2 ;
        RECT 0.4 17.036 14.8 17.068 ;
  LAYER M1 ;
        RECT 11.584 16.176 11.616 16.248 ;
  LAYER M2 ;
        RECT 11.564 16.196 11.636 16.228 ;
  LAYER M2 ;
        RECT 11.6 16.196 14.48 16.228 ;
  LAYER M1 ;
        RECT 14.464 16.176 14.496 16.248 ;
  LAYER M2 ;
        RECT 14.444 16.196 14.516 16.228 ;
  LAYER M1 ;
        RECT 11.584 4.416 11.616 4.488 ;
  LAYER M2 ;
        RECT 11.564 4.436 11.636 4.468 ;
  LAYER M2 ;
        RECT 11.6 4.436 14.48 4.468 ;
  LAYER M1 ;
        RECT 14.464 4.416 14.496 4.488 ;
  LAYER M2 ;
        RECT 14.444 4.436 14.516 4.468 ;
  LAYER M1 ;
        RECT 8.704 4.416 8.736 4.488 ;
  LAYER M2 ;
        RECT 8.684 4.436 8.756 4.468 ;
  LAYER M2 ;
        RECT 8.72 4.436 11.6 4.468 ;
  LAYER M1 ;
        RECT 11.584 4.416 11.616 4.488 ;
  LAYER M2 ;
        RECT 11.564 4.436 11.636 4.468 ;
  LAYER M1 ;
        RECT 5.824 4.416 5.856 4.488 ;
  LAYER M2 ;
        RECT 5.804 4.436 5.876 4.468 ;
  LAYER M2 ;
        RECT 5.84 4.436 8.72 4.468 ;
  LAYER M1 ;
        RECT 8.704 4.416 8.736 4.488 ;
  LAYER M2 ;
        RECT 8.684 4.436 8.756 4.468 ;
  LAYER M1 ;
        RECT 5.824 16.176 5.856 16.248 ;
  LAYER M2 ;
        RECT 5.804 16.196 5.876 16.228 ;
  LAYER M2 ;
        RECT 2.96 16.196 5.84 16.228 ;
  LAYER M1 ;
        RECT 2.944 16.176 2.976 16.248 ;
  LAYER M2 ;
        RECT 2.924 16.196 2.996 16.228 ;
  LAYER M1 ;
        RECT 8.704 16.176 8.736 16.248 ;
  LAYER M2 ;
        RECT 8.684 16.196 8.756 16.228 ;
  LAYER M2 ;
        RECT 5.84 16.196 8.72 16.228 ;
  LAYER M1 ;
        RECT 5.824 16.176 5.856 16.248 ;
  LAYER M2 ;
        RECT 5.804 16.196 5.876 16.228 ;
  LAYER M1 ;
        RECT 6.304 7.86 6.336 7.932 ;
  LAYER M2 ;
        RECT 6.284 7.88 6.356 7.912 ;
  LAYER M2 ;
        RECT 6.32 7.88 8.88 7.912 ;
  LAYER M1 ;
        RECT 8.864 7.86 8.896 7.932 ;
  LAYER M2 ;
        RECT 8.844 7.88 8.916 7.912 ;
  LAYER M1 ;
        RECT 9.184 4.92 9.216 4.992 ;
  LAYER M2 ;
        RECT 9.164 4.94 9.236 4.972 ;
  LAYER M1 ;
        RECT 9.184 4.788 9.216 4.956 ;
  LAYER M1 ;
        RECT 9.184 4.752 9.216 4.824 ;
  LAYER M2 ;
        RECT 9.164 4.772 9.236 4.804 ;
  LAYER M2 ;
        RECT 8.88 4.772 9.2 4.804 ;
  LAYER M1 ;
        RECT 8.864 4.752 8.896 4.824 ;
  LAYER M2 ;
        RECT 8.844 4.772 8.916 4.804 ;
  LAYER M1 ;
        RECT 8.864 1.476 8.896 1.548 ;
  LAYER M2 ;
        RECT 8.844 1.496 8.916 1.528 ;
  LAYER M1 ;
        RECT 8.864 1.512 8.896 1.68 ;
  LAYER M1 ;
        RECT 8.864 1.68 8.896 7.896 ;
  LAYER M1 ;
        RECT 3.424 10.8 3.456 10.872 ;
  LAYER M2 ;
        RECT 3.404 10.82 3.476 10.852 ;
  LAYER M2 ;
        RECT 3.44 10.82 6 10.852 ;
  LAYER M1 ;
        RECT 5.984 10.8 6.016 10.872 ;
  LAYER M2 ;
        RECT 5.964 10.82 6.036 10.852 ;
  LAYER M1 ;
        RECT 5.984 1.476 6.016 1.548 ;
  LAYER M2 ;
        RECT 5.964 1.496 6.036 1.528 ;
  LAYER M1 ;
        RECT 5.984 1.512 6.016 1.68 ;
  LAYER M1 ;
        RECT 5.984 1.68 6.016 10.836 ;
  LAYER M2 ;
        RECT 6 1.496 8.88 1.528 ;
  LAYER M1 ;
        RECT 9.184 7.86 9.216 7.932 ;
  LAYER M2 ;
        RECT 9.164 7.88 9.236 7.912 ;
  LAYER M2 ;
        RECT 9.2 7.88 11.76 7.912 ;
  LAYER M1 ;
        RECT 11.744 7.86 11.776 7.932 ;
  LAYER M2 ;
        RECT 11.724 7.88 11.796 7.912 ;
  LAYER M1 ;
        RECT 9.184 10.8 9.216 10.872 ;
  LAYER M2 ;
        RECT 9.164 10.82 9.236 10.852 ;
  LAYER M2 ;
        RECT 9.2 10.82 11.76 10.852 ;
  LAYER M1 ;
        RECT 11.744 10.8 11.776 10.872 ;
  LAYER M2 ;
        RECT 11.724 10.82 11.796 10.852 ;
  LAYER M1 ;
        RECT 11.744 1.308 11.776 1.38 ;
  LAYER M2 ;
        RECT 11.724 1.328 11.796 1.36 ;
  LAYER M1 ;
        RECT 11.744 1.344 11.776 1.68 ;
  LAYER M1 ;
        RECT 11.744 1.68 11.776 10.836 ;
  LAYER M1 ;
        RECT 3.424 7.86 3.456 7.932 ;
  LAYER M2 ;
        RECT 3.404 7.88 3.476 7.912 ;
  LAYER M1 ;
        RECT 3.424 7.728 3.456 7.896 ;
  LAYER M1 ;
        RECT 3.424 7.692 3.456 7.764 ;
  LAYER M2 ;
        RECT 3.404 7.712 3.476 7.744 ;
  LAYER M2 ;
        RECT 3.12 7.712 3.44 7.744 ;
  LAYER M1 ;
        RECT 3.104 7.692 3.136 7.764 ;
  LAYER M2 ;
        RECT 3.084 7.712 3.156 7.744 ;
  LAYER M1 ;
        RECT 3.424 4.92 3.456 4.992 ;
  LAYER M2 ;
        RECT 3.404 4.94 3.476 4.972 ;
  LAYER M1 ;
        RECT 3.424 4.788 3.456 4.956 ;
  LAYER M1 ;
        RECT 3.424 4.752 3.456 4.824 ;
  LAYER M2 ;
        RECT 3.404 4.772 3.476 4.804 ;
  LAYER M2 ;
        RECT 3.12 4.772 3.44 4.804 ;
  LAYER M1 ;
        RECT 3.104 4.752 3.136 4.824 ;
  LAYER M2 ;
        RECT 3.084 4.772 3.156 4.804 ;
  LAYER M1 ;
        RECT 3.104 1.308 3.136 1.38 ;
  LAYER M2 ;
        RECT 3.084 1.328 3.156 1.36 ;
  LAYER M1 ;
        RECT 3.104 1.344 3.136 1.68 ;
  LAYER M1 ;
        RECT 3.104 1.68 3.136 7.728 ;
  LAYER M2 ;
        RECT 3.12 1.328 11.76 1.36 ;
  LAYER M1 ;
        RECT 6.304 10.8 6.336 10.872 ;
  LAYER M2 ;
        RECT 6.284 10.82 6.356 10.852 ;
  LAYER M2 ;
        RECT 6.32 10.82 9.2 10.852 ;
  LAYER M1 ;
        RECT 9.184 10.8 9.216 10.872 ;
  LAYER M2 ;
        RECT 9.164 10.82 9.236 10.852 ;
  LAYER M1 ;
        RECT 6.304 4.92 6.336 4.992 ;
  LAYER M2 ;
        RECT 6.284 4.94 6.356 4.972 ;
  LAYER M2 ;
        RECT 3.44 4.94 6.32 4.972 ;
  LAYER M1 ;
        RECT 3.424 4.92 3.456 4.992 ;
  LAYER M2 ;
        RECT 3.404 4.94 3.476 4.972 ;
  LAYER M1 ;
        RECT 12.064 13.74 12.096 13.812 ;
  LAYER M2 ;
        RECT 12.044 13.76 12.116 13.792 ;
  LAYER M2 ;
        RECT 12.08 13.76 14.64 13.792 ;
  LAYER M1 ;
        RECT 14.624 13.74 14.656 13.812 ;
  LAYER M2 ;
        RECT 14.604 13.76 14.676 13.792 ;
  LAYER M1 ;
        RECT 12.064 10.8 12.096 10.872 ;
  LAYER M2 ;
        RECT 12.044 10.82 12.116 10.852 ;
  LAYER M2 ;
        RECT 12.08 10.82 14.64 10.852 ;
  LAYER M1 ;
        RECT 14.624 10.8 14.656 10.872 ;
  LAYER M2 ;
        RECT 14.604 10.82 14.676 10.852 ;
  LAYER M1 ;
        RECT 12.064 7.86 12.096 7.932 ;
  LAYER M2 ;
        RECT 12.044 7.88 12.116 7.912 ;
  LAYER M2 ;
        RECT 12.08 7.88 14.64 7.912 ;
  LAYER M1 ;
        RECT 14.624 7.86 14.656 7.932 ;
  LAYER M2 ;
        RECT 14.604 7.88 14.676 7.912 ;
  LAYER M1 ;
        RECT 12.064 4.92 12.096 4.992 ;
  LAYER M2 ;
        RECT 12.044 4.94 12.116 4.972 ;
  LAYER M2 ;
        RECT 12.08 4.94 14.64 4.972 ;
  LAYER M1 ;
        RECT 14.624 4.92 14.656 4.992 ;
  LAYER M2 ;
        RECT 14.604 4.94 14.676 4.972 ;
  LAYER M1 ;
        RECT 12.064 1.98 12.096 2.052 ;
  LAYER M2 ;
        RECT 12.044 2 12.116 2.032 ;
  LAYER M2 ;
        RECT 12.08 2 14.64 2.032 ;
  LAYER M1 ;
        RECT 14.624 1.98 14.656 2.052 ;
  LAYER M2 ;
        RECT 14.604 2 14.676 2.032 ;
  LAYER M1 ;
        RECT 14.624 1.14 14.656 1.212 ;
  LAYER M2 ;
        RECT 14.604 1.16 14.676 1.192 ;
  LAYER M1 ;
        RECT 14.624 1.176 14.656 1.68 ;
  LAYER M1 ;
        RECT 14.624 1.68 14.656 13.776 ;
  LAYER M1 ;
        RECT 0.544 13.74 0.576 13.812 ;
  LAYER M2 ;
        RECT 0.524 13.76 0.596 13.792 ;
  LAYER M1 ;
        RECT 0.544 13.608 0.576 13.776 ;
  LAYER M1 ;
        RECT 0.544 13.572 0.576 13.644 ;
  LAYER M2 ;
        RECT 0.524 13.592 0.596 13.624 ;
  LAYER M2 ;
        RECT 0.24 13.592 0.56 13.624 ;
  LAYER M1 ;
        RECT 0.224 13.572 0.256 13.644 ;
  LAYER M2 ;
        RECT 0.204 13.592 0.276 13.624 ;
  LAYER M1 ;
        RECT 0.544 10.8 0.576 10.872 ;
  LAYER M2 ;
        RECT 0.524 10.82 0.596 10.852 ;
  LAYER M1 ;
        RECT 0.544 10.668 0.576 10.836 ;
  LAYER M1 ;
        RECT 0.544 10.632 0.576 10.704 ;
  LAYER M2 ;
        RECT 0.524 10.652 0.596 10.684 ;
  LAYER M2 ;
        RECT 0.24 10.652 0.56 10.684 ;
  LAYER M1 ;
        RECT 0.224 10.632 0.256 10.704 ;
  LAYER M2 ;
        RECT 0.204 10.652 0.276 10.684 ;
  LAYER M1 ;
        RECT 0.544 7.86 0.576 7.932 ;
  LAYER M2 ;
        RECT 0.524 7.88 0.596 7.912 ;
  LAYER M1 ;
        RECT 0.544 7.728 0.576 7.896 ;
  LAYER M1 ;
        RECT 0.544 7.692 0.576 7.764 ;
  LAYER M2 ;
        RECT 0.524 7.712 0.596 7.744 ;
  LAYER M2 ;
        RECT 0.24 7.712 0.56 7.744 ;
  LAYER M1 ;
        RECT 0.224 7.692 0.256 7.764 ;
  LAYER M2 ;
        RECT 0.204 7.712 0.276 7.744 ;
  LAYER M1 ;
        RECT 0.544 4.92 0.576 4.992 ;
  LAYER M2 ;
        RECT 0.524 4.94 0.596 4.972 ;
  LAYER M1 ;
        RECT 0.544 4.788 0.576 4.956 ;
  LAYER M1 ;
        RECT 0.544 4.752 0.576 4.824 ;
  LAYER M2 ;
        RECT 0.524 4.772 0.596 4.804 ;
  LAYER M2 ;
        RECT 0.24 4.772 0.56 4.804 ;
  LAYER M1 ;
        RECT 0.224 4.752 0.256 4.824 ;
  LAYER M2 ;
        RECT 0.204 4.772 0.276 4.804 ;
  LAYER M1 ;
        RECT 0.544 1.98 0.576 2.052 ;
  LAYER M2 ;
        RECT 0.524 2 0.596 2.032 ;
  LAYER M1 ;
        RECT 0.544 1.848 0.576 2.016 ;
  LAYER M1 ;
        RECT 0.544 1.812 0.576 1.884 ;
  LAYER M2 ;
        RECT 0.524 1.832 0.596 1.864 ;
  LAYER M2 ;
        RECT 0.24 1.832 0.56 1.864 ;
  LAYER M1 ;
        RECT 0.224 1.812 0.256 1.884 ;
  LAYER M2 ;
        RECT 0.204 1.832 0.276 1.864 ;
  LAYER M1 ;
        RECT 0.224 1.14 0.256 1.212 ;
  LAYER M2 ;
        RECT 0.204 1.16 0.276 1.192 ;
  LAYER M1 ;
        RECT 0.224 1.176 0.256 1.68 ;
  LAYER M1 ;
        RECT 0.224 1.68 0.256 13.608 ;
  LAYER M2 ;
        RECT 0.24 1.16 14.64 1.192 ;
  LAYER M1 ;
        RECT 9.184 13.74 9.216 13.812 ;
  LAYER M2 ;
        RECT 9.164 13.76 9.236 13.792 ;
  LAYER M2 ;
        RECT 9.2 13.76 12.08 13.792 ;
  LAYER M1 ;
        RECT 12.064 13.74 12.096 13.812 ;
  LAYER M2 ;
        RECT 12.044 13.76 12.116 13.792 ;
  LAYER M1 ;
        RECT 9.184 1.98 9.216 2.052 ;
  LAYER M2 ;
        RECT 9.164 2 9.236 2.032 ;
  LAYER M2 ;
        RECT 9.2 2 12.08 2.032 ;
  LAYER M1 ;
        RECT 12.064 1.98 12.096 2.052 ;
  LAYER M2 ;
        RECT 12.044 2 12.116 2.032 ;
  LAYER M1 ;
        RECT 6.304 1.98 6.336 2.052 ;
  LAYER M2 ;
        RECT 6.284 2 6.356 2.032 ;
  LAYER M2 ;
        RECT 6.32 2 9.2 2.032 ;
  LAYER M1 ;
        RECT 9.184 1.98 9.216 2.052 ;
  LAYER M2 ;
        RECT 9.164 2 9.236 2.032 ;
  LAYER M1 ;
        RECT 3.424 1.98 3.456 2.052 ;
  LAYER M2 ;
        RECT 3.404 2 3.476 2.032 ;
  LAYER M2 ;
        RECT 3.44 2 6.32 2.032 ;
  LAYER M1 ;
        RECT 6.304 1.98 6.336 2.052 ;
  LAYER M2 ;
        RECT 6.284 2 6.356 2.032 ;
  LAYER M1 ;
        RECT 3.424 13.74 3.456 13.812 ;
  LAYER M2 ;
        RECT 3.404 13.76 3.476 13.792 ;
  LAYER M2 ;
        RECT 0.56 13.76 3.44 13.792 ;
  LAYER M1 ;
        RECT 0.544 13.74 0.576 13.812 ;
  LAYER M2 ;
        RECT 0.524 13.76 0.596 13.792 ;
  LAYER M1 ;
        RECT 6.304 13.74 6.336 13.812 ;
  LAYER M2 ;
        RECT 6.284 13.76 6.356 13.792 ;
  LAYER M2 ;
        RECT 3.44 13.76 6.32 13.792 ;
  LAYER M1 ;
        RECT 3.424 13.74 3.456 13.812 ;
  LAYER M2 ;
        RECT 3.404 13.76 3.476 13.792 ;
  LAYER M1 ;
        RECT 14.464 13.74 14.496 16.248 ;
  LAYER M1 ;
        RECT 14.4 13.74 14.432 16.248 ;
  LAYER M1 ;
        RECT 14.336 13.74 14.368 16.248 ;
  LAYER M1 ;
        RECT 14.272 13.74 14.304 16.248 ;
  LAYER M1 ;
        RECT 14.208 13.74 14.24 16.248 ;
  LAYER M1 ;
        RECT 14.144 13.74 14.176 16.248 ;
  LAYER M1 ;
        RECT 14.08 13.74 14.112 16.248 ;
  LAYER M1 ;
        RECT 14.016 13.74 14.048 16.248 ;
  LAYER M1 ;
        RECT 13.952 13.74 13.984 16.248 ;
  LAYER M1 ;
        RECT 13.888 13.74 13.92 16.248 ;
  LAYER M1 ;
        RECT 13.824 13.74 13.856 16.248 ;
  LAYER M1 ;
        RECT 13.76 13.74 13.792 16.248 ;
  LAYER M1 ;
        RECT 13.696 13.74 13.728 16.248 ;
  LAYER M1 ;
        RECT 13.632 13.74 13.664 16.248 ;
  LAYER M1 ;
        RECT 13.568 13.74 13.6 16.248 ;
  LAYER M1 ;
        RECT 13.504 13.74 13.536 16.248 ;
  LAYER M1 ;
        RECT 13.44 13.74 13.472 16.248 ;
  LAYER M1 ;
        RECT 13.376 13.74 13.408 16.248 ;
  LAYER M1 ;
        RECT 13.312 13.74 13.344 16.248 ;
  LAYER M1 ;
        RECT 13.248 13.74 13.28 16.248 ;
  LAYER M1 ;
        RECT 13.184 13.74 13.216 16.248 ;
  LAYER M1 ;
        RECT 13.12 13.74 13.152 16.248 ;
  LAYER M1 ;
        RECT 13.056 13.74 13.088 16.248 ;
  LAYER M1 ;
        RECT 12.992 13.74 13.024 16.248 ;
  LAYER M1 ;
        RECT 12.928 13.74 12.96 16.248 ;
  LAYER M1 ;
        RECT 12.864 13.74 12.896 16.248 ;
  LAYER M1 ;
        RECT 12.8 13.74 12.832 16.248 ;
  LAYER M1 ;
        RECT 12.736 13.74 12.768 16.248 ;
  LAYER M1 ;
        RECT 12.672 13.74 12.704 16.248 ;
  LAYER M1 ;
        RECT 12.608 13.74 12.64 16.248 ;
  LAYER M1 ;
        RECT 12.544 13.74 12.576 16.248 ;
  LAYER M1 ;
        RECT 12.48 13.74 12.512 16.248 ;
  LAYER M1 ;
        RECT 12.416 13.74 12.448 16.248 ;
  LAYER M1 ;
        RECT 12.352 13.74 12.384 16.248 ;
  LAYER M1 ;
        RECT 12.288 13.74 12.32 16.248 ;
  LAYER M1 ;
        RECT 12.224 13.74 12.256 16.248 ;
  LAYER M1 ;
        RECT 12.16 13.74 12.192 16.248 ;
  LAYER M2 ;
        RECT 12.044 16.132 14.516 16.164 ;
  LAYER M2 ;
        RECT 12.044 16.068 14.516 16.1 ;
  LAYER M2 ;
        RECT 12.044 16.004 14.516 16.036 ;
  LAYER M2 ;
        RECT 12.044 15.94 14.516 15.972 ;
  LAYER M2 ;
        RECT 12.044 15.876 14.516 15.908 ;
  LAYER M2 ;
        RECT 12.044 15.812 14.516 15.844 ;
  LAYER M2 ;
        RECT 12.044 15.748 14.516 15.78 ;
  LAYER M2 ;
        RECT 12.044 15.684 14.516 15.716 ;
  LAYER M2 ;
        RECT 12.044 15.62 14.516 15.652 ;
  LAYER M2 ;
        RECT 12.044 15.556 14.516 15.588 ;
  LAYER M2 ;
        RECT 12.044 15.492 14.516 15.524 ;
  LAYER M2 ;
        RECT 12.044 15.428 14.516 15.46 ;
  LAYER M2 ;
        RECT 12.044 15.364 14.516 15.396 ;
  LAYER M2 ;
        RECT 12.044 15.3 14.516 15.332 ;
  LAYER M2 ;
        RECT 12.044 15.236 14.516 15.268 ;
  LAYER M2 ;
        RECT 12.044 15.172 14.516 15.204 ;
  LAYER M2 ;
        RECT 12.044 15.108 14.516 15.14 ;
  LAYER M2 ;
        RECT 12.044 15.044 14.516 15.076 ;
  LAYER M2 ;
        RECT 12.044 14.98 14.516 15.012 ;
  LAYER M2 ;
        RECT 12.044 14.916 14.516 14.948 ;
  LAYER M2 ;
        RECT 12.044 14.852 14.516 14.884 ;
  LAYER M2 ;
        RECT 12.044 14.788 14.516 14.82 ;
  LAYER M2 ;
        RECT 12.044 14.724 14.516 14.756 ;
  LAYER M2 ;
        RECT 12.044 14.66 14.516 14.692 ;
  LAYER M2 ;
        RECT 12.044 14.596 14.516 14.628 ;
  LAYER M2 ;
        RECT 12.044 14.532 14.516 14.564 ;
  LAYER M2 ;
        RECT 12.044 14.468 14.516 14.5 ;
  LAYER M2 ;
        RECT 12.044 14.404 14.516 14.436 ;
  LAYER M2 ;
        RECT 12.044 14.34 14.516 14.372 ;
  LAYER M2 ;
        RECT 12.044 14.276 14.516 14.308 ;
  LAYER M2 ;
        RECT 12.044 14.212 14.516 14.244 ;
  LAYER M2 ;
        RECT 12.044 14.148 14.516 14.18 ;
  LAYER M2 ;
        RECT 12.044 14.084 14.516 14.116 ;
  LAYER M2 ;
        RECT 12.044 14.02 14.516 14.052 ;
  LAYER M2 ;
        RECT 12.044 13.956 14.516 13.988 ;
  LAYER M2 ;
        RECT 12.044 13.892 14.516 13.924 ;
  LAYER M3 ;
        RECT 14.464 13.74 14.496 16.248 ;
  LAYER M3 ;
        RECT 14.4 13.74 14.432 16.248 ;
  LAYER M3 ;
        RECT 14.336 13.74 14.368 16.248 ;
  LAYER M3 ;
        RECT 14.272 13.74 14.304 16.248 ;
  LAYER M3 ;
        RECT 14.208 13.74 14.24 16.248 ;
  LAYER M3 ;
        RECT 14.144 13.74 14.176 16.248 ;
  LAYER M3 ;
        RECT 14.08 13.74 14.112 16.248 ;
  LAYER M3 ;
        RECT 14.016 13.74 14.048 16.248 ;
  LAYER M3 ;
        RECT 13.952 13.74 13.984 16.248 ;
  LAYER M3 ;
        RECT 13.888 13.74 13.92 16.248 ;
  LAYER M3 ;
        RECT 13.824 13.74 13.856 16.248 ;
  LAYER M3 ;
        RECT 13.76 13.74 13.792 16.248 ;
  LAYER M3 ;
        RECT 13.696 13.74 13.728 16.248 ;
  LAYER M3 ;
        RECT 13.632 13.74 13.664 16.248 ;
  LAYER M3 ;
        RECT 13.568 13.74 13.6 16.248 ;
  LAYER M3 ;
        RECT 13.504 13.74 13.536 16.248 ;
  LAYER M3 ;
        RECT 13.44 13.74 13.472 16.248 ;
  LAYER M3 ;
        RECT 13.376 13.74 13.408 16.248 ;
  LAYER M3 ;
        RECT 13.312 13.74 13.344 16.248 ;
  LAYER M3 ;
        RECT 13.248 13.74 13.28 16.248 ;
  LAYER M3 ;
        RECT 13.184 13.74 13.216 16.248 ;
  LAYER M3 ;
        RECT 13.12 13.74 13.152 16.248 ;
  LAYER M3 ;
        RECT 13.056 13.74 13.088 16.248 ;
  LAYER M3 ;
        RECT 12.992 13.74 13.024 16.248 ;
  LAYER M3 ;
        RECT 12.928 13.74 12.96 16.248 ;
  LAYER M3 ;
        RECT 12.864 13.74 12.896 16.248 ;
  LAYER M3 ;
        RECT 12.8 13.74 12.832 16.248 ;
  LAYER M3 ;
        RECT 12.736 13.74 12.768 16.248 ;
  LAYER M3 ;
        RECT 12.672 13.74 12.704 16.248 ;
  LAYER M3 ;
        RECT 12.608 13.74 12.64 16.248 ;
  LAYER M3 ;
        RECT 12.544 13.74 12.576 16.248 ;
  LAYER M3 ;
        RECT 12.48 13.74 12.512 16.248 ;
  LAYER M3 ;
        RECT 12.416 13.74 12.448 16.248 ;
  LAYER M3 ;
        RECT 12.352 13.74 12.384 16.248 ;
  LAYER M3 ;
        RECT 12.288 13.74 12.32 16.248 ;
  LAYER M3 ;
        RECT 12.224 13.74 12.256 16.248 ;
  LAYER M3 ;
        RECT 12.16 13.74 12.192 16.248 ;
  LAYER M3 ;
        RECT 12.064 13.74 12.096 16.248 ;
  LAYER M1 ;
        RECT 14.479 13.776 14.481 16.212 ;
  LAYER M1 ;
        RECT 14.399 13.776 14.401 16.212 ;
  LAYER M1 ;
        RECT 14.319 13.776 14.321 16.212 ;
  LAYER M1 ;
        RECT 14.239 13.776 14.241 16.212 ;
  LAYER M1 ;
        RECT 14.159 13.776 14.161 16.212 ;
  LAYER M1 ;
        RECT 14.079 13.776 14.081 16.212 ;
  LAYER M1 ;
        RECT 13.999 13.776 14.001 16.212 ;
  LAYER M1 ;
        RECT 13.919 13.776 13.921 16.212 ;
  LAYER M1 ;
        RECT 13.839 13.776 13.841 16.212 ;
  LAYER M1 ;
        RECT 13.759 13.776 13.761 16.212 ;
  LAYER M1 ;
        RECT 13.679 13.776 13.681 16.212 ;
  LAYER M1 ;
        RECT 13.599 13.776 13.601 16.212 ;
  LAYER M1 ;
        RECT 13.519 13.776 13.521 16.212 ;
  LAYER M1 ;
        RECT 13.439 13.776 13.441 16.212 ;
  LAYER M1 ;
        RECT 13.359 13.776 13.361 16.212 ;
  LAYER M1 ;
        RECT 13.279 13.776 13.281 16.212 ;
  LAYER M1 ;
        RECT 13.199 13.776 13.201 16.212 ;
  LAYER M1 ;
        RECT 13.119 13.776 13.121 16.212 ;
  LAYER M1 ;
        RECT 13.039 13.776 13.041 16.212 ;
  LAYER M1 ;
        RECT 12.959 13.776 12.961 16.212 ;
  LAYER M1 ;
        RECT 12.879 13.776 12.881 16.212 ;
  LAYER M1 ;
        RECT 12.799 13.776 12.801 16.212 ;
  LAYER M1 ;
        RECT 12.719 13.776 12.721 16.212 ;
  LAYER M1 ;
        RECT 12.639 13.776 12.641 16.212 ;
  LAYER M1 ;
        RECT 12.559 13.776 12.561 16.212 ;
  LAYER M1 ;
        RECT 12.479 13.776 12.481 16.212 ;
  LAYER M1 ;
        RECT 12.399 13.776 12.401 16.212 ;
  LAYER M1 ;
        RECT 12.319 13.776 12.321 16.212 ;
  LAYER M1 ;
        RECT 12.239 13.776 12.241 16.212 ;
  LAYER M1 ;
        RECT 12.159 13.776 12.161 16.212 ;
  LAYER M2 ;
        RECT 12.08 16.211 14.48 16.213 ;
  LAYER M2 ;
        RECT 12.08 16.127 14.48 16.129 ;
  LAYER M2 ;
        RECT 12.08 16.043 14.48 16.045 ;
  LAYER M2 ;
        RECT 12.08 15.959 14.48 15.961 ;
  LAYER M2 ;
        RECT 12.08 15.875 14.48 15.877 ;
  LAYER M2 ;
        RECT 12.08 15.791 14.48 15.793 ;
  LAYER M2 ;
        RECT 12.08 15.707 14.48 15.709 ;
  LAYER M2 ;
        RECT 12.08 15.623 14.48 15.625 ;
  LAYER M2 ;
        RECT 12.08 15.539 14.48 15.541 ;
  LAYER M2 ;
        RECT 12.08 15.455 14.48 15.457 ;
  LAYER M2 ;
        RECT 12.08 15.371 14.48 15.373 ;
  LAYER M2 ;
        RECT 12.08 15.287 14.48 15.289 ;
  LAYER M2 ;
        RECT 12.08 15.2035 14.48 15.2055 ;
  LAYER M2 ;
        RECT 12.08 15.119 14.48 15.121 ;
  LAYER M2 ;
        RECT 12.08 15.035 14.48 15.037 ;
  LAYER M2 ;
        RECT 12.08 14.951 14.48 14.953 ;
  LAYER M2 ;
        RECT 12.08 14.867 14.48 14.869 ;
  LAYER M2 ;
        RECT 12.08 14.783 14.48 14.785 ;
  LAYER M2 ;
        RECT 12.08 14.699 14.48 14.701 ;
  LAYER M2 ;
        RECT 12.08 14.615 14.48 14.617 ;
  LAYER M2 ;
        RECT 12.08 14.531 14.48 14.533 ;
  LAYER M2 ;
        RECT 12.08 14.447 14.48 14.449 ;
  LAYER M2 ;
        RECT 12.08 14.363 14.48 14.365 ;
  LAYER M2 ;
        RECT 12.08 14.279 14.48 14.281 ;
  LAYER M2 ;
        RECT 12.08 14.195 14.48 14.197 ;
  LAYER M2 ;
        RECT 12.08 14.111 14.48 14.113 ;
  LAYER M2 ;
        RECT 12.08 14.027 14.48 14.029 ;
  LAYER M2 ;
        RECT 12.08 13.943 14.48 13.945 ;
  LAYER M2 ;
        RECT 12.08 13.859 14.48 13.861 ;
  LAYER M1 ;
        RECT 14.464 10.8 14.496 13.308 ;
  LAYER M1 ;
        RECT 14.4 10.8 14.432 13.308 ;
  LAYER M1 ;
        RECT 14.336 10.8 14.368 13.308 ;
  LAYER M1 ;
        RECT 14.272 10.8 14.304 13.308 ;
  LAYER M1 ;
        RECT 14.208 10.8 14.24 13.308 ;
  LAYER M1 ;
        RECT 14.144 10.8 14.176 13.308 ;
  LAYER M1 ;
        RECT 14.08 10.8 14.112 13.308 ;
  LAYER M1 ;
        RECT 14.016 10.8 14.048 13.308 ;
  LAYER M1 ;
        RECT 13.952 10.8 13.984 13.308 ;
  LAYER M1 ;
        RECT 13.888 10.8 13.92 13.308 ;
  LAYER M1 ;
        RECT 13.824 10.8 13.856 13.308 ;
  LAYER M1 ;
        RECT 13.76 10.8 13.792 13.308 ;
  LAYER M1 ;
        RECT 13.696 10.8 13.728 13.308 ;
  LAYER M1 ;
        RECT 13.632 10.8 13.664 13.308 ;
  LAYER M1 ;
        RECT 13.568 10.8 13.6 13.308 ;
  LAYER M1 ;
        RECT 13.504 10.8 13.536 13.308 ;
  LAYER M1 ;
        RECT 13.44 10.8 13.472 13.308 ;
  LAYER M1 ;
        RECT 13.376 10.8 13.408 13.308 ;
  LAYER M1 ;
        RECT 13.312 10.8 13.344 13.308 ;
  LAYER M1 ;
        RECT 13.248 10.8 13.28 13.308 ;
  LAYER M1 ;
        RECT 13.184 10.8 13.216 13.308 ;
  LAYER M1 ;
        RECT 13.12 10.8 13.152 13.308 ;
  LAYER M1 ;
        RECT 13.056 10.8 13.088 13.308 ;
  LAYER M1 ;
        RECT 12.992 10.8 13.024 13.308 ;
  LAYER M1 ;
        RECT 12.928 10.8 12.96 13.308 ;
  LAYER M1 ;
        RECT 12.864 10.8 12.896 13.308 ;
  LAYER M1 ;
        RECT 12.8 10.8 12.832 13.308 ;
  LAYER M1 ;
        RECT 12.736 10.8 12.768 13.308 ;
  LAYER M1 ;
        RECT 12.672 10.8 12.704 13.308 ;
  LAYER M1 ;
        RECT 12.608 10.8 12.64 13.308 ;
  LAYER M1 ;
        RECT 12.544 10.8 12.576 13.308 ;
  LAYER M1 ;
        RECT 12.48 10.8 12.512 13.308 ;
  LAYER M1 ;
        RECT 12.416 10.8 12.448 13.308 ;
  LAYER M1 ;
        RECT 12.352 10.8 12.384 13.308 ;
  LAYER M1 ;
        RECT 12.288 10.8 12.32 13.308 ;
  LAYER M1 ;
        RECT 12.224 10.8 12.256 13.308 ;
  LAYER M1 ;
        RECT 12.16 10.8 12.192 13.308 ;
  LAYER M2 ;
        RECT 12.044 13.192 14.516 13.224 ;
  LAYER M2 ;
        RECT 12.044 13.128 14.516 13.16 ;
  LAYER M2 ;
        RECT 12.044 13.064 14.516 13.096 ;
  LAYER M2 ;
        RECT 12.044 13 14.516 13.032 ;
  LAYER M2 ;
        RECT 12.044 12.936 14.516 12.968 ;
  LAYER M2 ;
        RECT 12.044 12.872 14.516 12.904 ;
  LAYER M2 ;
        RECT 12.044 12.808 14.516 12.84 ;
  LAYER M2 ;
        RECT 12.044 12.744 14.516 12.776 ;
  LAYER M2 ;
        RECT 12.044 12.68 14.516 12.712 ;
  LAYER M2 ;
        RECT 12.044 12.616 14.516 12.648 ;
  LAYER M2 ;
        RECT 12.044 12.552 14.516 12.584 ;
  LAYER M2 ;
        RECT 12.044 12.488 14.516 12.52 ;
  LAYER M2 ;
        RECT 12.044 12.424 14.516 12.456 ;
  LAYER M2 ;
        RECT 12.044 12.36 14.516 12.392 ;
  LAYER M2 ;
        RECT 12.044 12.296 14.516 12.328 ;
  LAYER M2 ;
        RECT 12.044 12.232 14.516 12.264 ;
  LAYER M2 ;
        RECT 12.044 12.168 14.516 12.2 ;
  LAYER M2 ;
        RECT 12.044 12.104 14.516 12.136 ;
  LAYER M2 ;
        RECT 12.044 12.04 14.516 12.072 ;
  LAYER M2 ;
        RECT 12.044 11.976 14.516 12.008 ;
  LAYER M2 ;
        RECT 12.044 11.912 14.516 11.944 ;
  LAYER M2 ;
        RECT 12.044 11.848 14.516 11.88 ;
  LAYER M2 ;
        RECT 12.044 11.784 14.516 11.816 ;
  LAYER M2 ;
        RECT 12.044 11.72 14.516 11.752 ;
  LAYER M2 ;
        RECT 12.044 11.656 14.516 11.688 ;
  LAYER M2 ;
        RECT 12.044 11.592 14.516 11.624 ;
  LAYER M2 ;
        RECT 12.044 11.528 14.516 11.56 ;
  LAYER M2 ;
        RECT 12.044 11.464 14.516 11.496 ;
  LAYER M2 ;
        RECT 12.044 11.4 14.516 11.432 ;
  LAYER M2 ;
        RECT 12.044 11.336 14.516 11.368 ;
  LAYER M2 ;
        RECT 12.044 11.272 14.516 11.304 ;
  LAYER M2 ;
        RECT 12.044 11.208 14.516 11.24 ;
  LAYER M2 ;
        RECT 12.044 11.144 14.516 11.176 ;
  LAYER M2 ;
        RECT 12.044 11.08 14.516 11.112 ;
  LAYER M2 ;
        RECT 12.044 11.016 14.516 11.048 ;
  LAYER M2 ;
        RECT 12.044 10.952 14.516 10.984 ;
  LAYER M3 ;
        RECT 14.464 10.8 14.496 13.308 ;
  LAYER M3 ;
        RECT 14.4 10.8 14.432 13.308 ;
  LAYER M3 ;
        RECT 14.336 10.8 14.368 13.308 ;
  LAYER M3 ;
        RECT 14.272 10.8 14.304 13.308 ;
  LAYER M3 ;
        RECT 14.208 10.8 14.24 13.308 ;
  LAYER M3 ;
        RECT 14.144 10.8 14.176 13.308 ;
  LAYER M3 ;
        RECT 14.08 10.8 14.112 13.308 ;
  LAYER M3 ;
        RECT 14.016 10.8 14.048 13.308 ;
  LAYER M3 ;
        RECT 13.952 10.8 13.984 13.308 ;
  LAYER M3 ;
        RECT 13.888 10.8 13.92 13.308 ;
  LAYER M3 ;
        RECT 13.824 10.8 13.856 13.308 ;
  LAYER M3 ;
        RECT 13.76 10.8 13.792 13.308 ;
  LAYER M3 ;
        RECT 13.696 10.8 13.728 13.308 ;
  LAYER M3 ;
        RECT 13.632 10.8 13.664 13.308 ;
  LAYER M3 ;
        RECT 13.568 10.8 13.6 13.308 ;
  LAYER M3 ;
        RECT 13.504 10.8 13.536 13.308 ;
  LAYER M3 ;
        RECT 13.44 10.8 13.472 13.308 ;
  LAYER M3 ;
        RECT 13.376 10.8 13.408 13.308 ;
  LAYER M3 ;
        RECT 13.312 10.8 13.344 13.308 ;
  LAYER M3 ;
        RECT 13.248 10.8 13.28 13.308 ;
  LAYER M3 ;
        RECT 13.184 10.8 13.216 13.308 ;
  LAYER M3 ;
        RECT 13.12 10.8 13.152 13.308 ;
  LAYER M3 ;
        RECT 13.056 10.8 13.088 13.308 ;
  LAYER M3 ;
        RECT 12.992 10.8 13.024 13.308 ;
  LAYER M3 ;
        RECT 12.928 10.8 12.96 13.308 ;
  LAYER M3 ;
        RECT 12.864 10.8 12.896 13.308 ;
  LAYER M3 ;
        RECT 12.8 10.8 12.832 13.308 ;
  LAYER M3 ;
        RECT 12.736 10.8 12.768 13.308 ;
  LAYER M3 ;
        RECT 12.672 10.8 12.704 13.308 ;
  LAYER M3 ;
        RECT 12.608 10.8 12.64 13.308 ;
  LAYER M3 ;
        RECT 12.544 10.8 12.576 13.308 ;
  LAYER M3 ;
        RECT 12.48 10.8 12.512 13.308 ;
  LAYER M3 ;
        RECT 12.416 10.8 12.448 13.308 ;
  LAYER M3 ;
        RECT 12.352 10.8 12.384 13.308 ;
  LAYER M3 ;
        RECT 12.288 10.8 12.32 13.308 ;
  LAYER M3 ;
        RECT 12.224 10.8 12.256 13.308 ;
  LAYER M3 ;
        RECT 12.16 10.8 12.192 13.308 ;
  LAYER M3 ;
        RECT 12.064 10.8 12.096 13.308 ;
  LAYER M1 ;
        RECT 14.479 10.836 14.481 13.272 ;
  LAYER M1 ;
        RECT 14.399 10.836 14.401 13.272 ;
  LAYER M1 ;
        RECT 14.319 10.836 14.321 13.272 ;
  LAYER M1 ;
        RECT 14.239 10.836 14.241 13.272 ;
  LAYER M1 ;
        RECT 14.159 10.836 14.161 13.272 ;
  LAYER M1 ;
        RECT 14.079 10.836 14.081 13.272 ;
  LAYER M1 ;
        RECT 13.999 10.836 14.001 13.272 ;
  LAYER M1 ;
        RECT 13.919 10.836 13.921 13.272 ;
  LAYER M1 ;
        RECT 13.839 10.836 13.841 13.272 ;
  LAYER M1 ;
        RECT 13.759 10.836 13.761 13.272 ;
  LAYER M1 ;
        RECT 13.679 10.836 13.681 13.272 ;
  LAYER M1 ;
        RECT 13.599 10.836 13.601 13.272 ;
  LAYER M1 ;
        RECT 13.519 10.836 13.521 13.272 ;
  LAYER M1 ;
        RECT 13.439 10.836 13.441 13.272 ;
  LAYER M1 ;
        RECT 13.359 10.836 13.361 13.272 ;
  LAYER M1 ;
        RECT 13.279 10.836 13.281 13.272 ;
  LAYER M1 ;
        RECT 13.199 10.836 13.201 13.272 ;
  LAYER M1 ;
        RECT 13.119 10.836 13.121 13.272 ;
  LAYER M1 ;
        RECT 13.039 10.836 13.041 13.272 ;
  LAYER M1 ;
        RECT 12.959 10.836 12.961 13.272 ;
  LAYER M1 ;
        RECT 12.879 10.836 12.881 13.272 ;
  LAYER M1 ;
        RECT 12.799 10.836 12.801 13.272 ;
  LAYER M1 ;
        RECT 12.719 10.836 12.721 13.272 ;
  LAYER M1 ;
        RECT 12.639 10.836 12.641 13.272 ;
  LAYER M1 ;
        RECT 12.559 10.836 12.561 13.272 ;
  LAYER M1 ;
        RECT 12.479 10.836 12.481 13.272 ;
  LAYER M1 ;
        RECT 12.399 10.836 12.401 13.272 ;
  LAYER M1 ;
        RECT 12.319 10.836 12.321 13.272 ;
  LAYER M1 ;
        RECT 12.239 10.836 12.241 13.272 ;
  LAYER M1 ;
        RECT 12.159 10.836 12.161 13.272 ;
  LAYER M2 ;
        RECT 12.08 13.271 14.48 13.273 ;
  LAYER M2 ;
        RECT 12.08 13.187 14.48 13.189 ;
  LAYER M2 ;
        RECT 12.08 13.103 14.48 13.105 ;
  LAYER M2 ;
        RECT 12.08 13.019 14.48 13.021 ;
  LAYER M2 ;
        RECT 12.08 12.935 14.48 12.937 ;
  LAYER M2 ;
        RECT 12.08 12.851 14.48 12.853 ;
  LAYER M2 ;
        RECT 12.08 12.767 14.48 12.769 ;
  LAYER M2 ;
        RECT 12.08 12.683 14.48 12.685 ;
  LAYER M2 ;
        RECT 12.08 12.599 14.48 12.601 ;
  LAYER M2 ;
        RECT 12.08 12.515 14.48 12.517 ;
  LAYER M2 ;
        RECT 12.08 12.431 14.48 12.433 ;
  LAYER M2 ;
        RECT 12.08 12.347 14.48 12.349 ;
  LAYER M2 ;
        RECT 12.08 12.2635 14.48 12.2655 ;
  LAYER M2 ;
        RECT 12.08 12.179 14.48 12.181 ;
  LAYER M2 ;
        RECT 12.08 12.095 14.48 12.097 ;
  LAYER M2 ;
        RECT 12.08 12.011 14.48 12.013 ;
  LAYER M2 ;
        RECT 12.08 11.927 14.48 11.929 ;
  LAYER M2 ;
        RECT 12.08 11.843 14.48 11.845 ;
  LAYER M2 ;
        RECT 12.08 11.759 14.48 11.761 ;
  LAYER M2 ;
        RECT 12.08 11.675 14.48 11.677 ;
  LAYER M2 ;
        RECT 12.08 11.591 14.48 11.593 ;
  LAYER M2 ;
        RECT 12.08 11.507 14.48 11.509 ;
  LAYER M2 ;
        RECT 12.08 11.423 14.48 11.425 ;
  LAYER M2 ;
        RECT 12.08 11.339 14.48 11.341 ;
  LAYER M2 ;
        RECT 12.08 11.255 14.48 11.257 ;
  LAYER M2 ;
        RECT 12.08 11.171 14.48 11.173 ;
  LAYER M2 ;
        RECT 12.08 11.087 14.48 11.089 ;
  LAYER M2 ;
        RECT 12.08 11.003 14.48 11.005 ;
  LAYER M2 ;
        RECT 12.08 10.919 14.48 10.921 ;
  LAYER M1 ;
        RECT 14.464 7.86 14.496 10.368 ;
  LAYER M1 ;
        RECT 14.4 7.86 14.432 10.368 ;
  LAYER M1 ;
        RECT 14.336 7.86 14.368 10.368 ;
  LAYER M1 ;
        RECT 14.272 7.86 14.304 10.368 ;
  LAYER M1 ;
        RECT 14.208 7.86 14.24 10.368 ;
  LAYER M1 ;
        RECT 14.144 7.86 14.176 10.368 ;
  LAYER M1 ;
        RECT 14.08 7.86 14.112 10.368 ;
  LAYER M1 ;
        RECT 14.016 7.86 14.048 10.368 ;
  LAYER M1 ;
        RECT 13.952 7.86 13.984 10.368 ;
  LAYER M1 ;
        RECT 13.888 7.86 13.92 10.368 ;
  LAYER M1 ;
        RECT 13.824 7.86 13.856 10.368 ;
  LAYER M1 ;
        RECT 13.76 7.86 13.792 10.368 ;
  LAYER M1 ;
        RECT 13.696 7.86 13.728 10.368 ;
  LAYER M1 ;
        RECT 13.632 7.86 13.664 10.368 ;
  LAYER M1 ;
        RECT 13.568 7.86 13.6 10.368 ;
  LAYER M1 ;
        RECT 13.504 7.86 13.536 10.368 ;
  LAYER M1 ;
        RECT 13.44 7.86 13.472 10.368 ;
  LAYER M1 ;
        RECT 13.376 7.86 13.408 10.368 ;
  LAYER M1 ;
        RECT 13.312 7.86 13.344 10.368 ;
  LAYER M1 ;
        RECT 13.248 7.86 13.28 10.368 ;
  LAYER M1 ;
        RECT 13.184 7.86 13.216 10.368 ;
  LAYER M1 ;
        RECT 13.12 7.86 13.152 10.368 ;
  LAYER M1 ;
        RECT 13.056 7.86 13.088 10.368 ;
  LAYER M1 ;
        RECT 12.992 7.86 13.024 10.368 ;
  LAYER M1 ;
        RECT 12.928 7.86 12.96 10.368 ;
  LAYER M1 ;
        RECT 12.864 7.86 12.896 10.368 ;
  LAYER M1 ;
        RECT 12.8 7.86 12.832 10.368 ;
  LAYER M1 ;
        RECT 12.736 7.86 12.768 10.368 ;
  LAYER M1 ;
        RECT 12.672 7.86 12.704 10.368 ;
  LAYER M1 ;
        RECT 12.608 7.86 12.64 10.368 ;
  LAYER M1 ;
        RECT 12.544 7.86 12.576 10.368 ;
  LAYER M1 ;
        RECT 12.48 7.86 12.512 10.368 ;
  LAYER M1 ;
        RECT 12.416 7.86 12.448 10.368 ;
  LAYER M1 ;
        RECT 12.352 7.86 12.384 10.368 ;
  LAYER M1 ;
        RECT 12.288 7.86 12.32 10.368 ;
  LAYER M1 ;
        RECT 12.224 7.86 12.256 10.368 ;
  LAYER M1 ;
        RECT 12.16 7.86 12.192 10.368 ;
  LAYER M2 ;
        RECT 12.044 10.252 14.516 10.284 ;
  LAYER M2 ;
        RECT 12.044 10.188 14.516 10.22 ;
  LAYER M2 ;
        RECT 12.044 10.124 14.516 10.156 ;
  LAYER M2 ;
        RECT 12.044 10.06 14.516 10.092 ;
  LAYER M2 ;
        RECT 12.044 9.996 14.516 10.028 ;
  LAYER M2 ;
        RECT 12.044 9.932 14.516 9.964 ;
  LAYER M2 ;
        RECT 12.044 9.868 14.516 9.9 ;
  LAYER M2 ;
        RECT 12.044 9.804 14.516 9.836 ;
  LAYER M2 ;
        RECT 12.044 9.74 14.516 9.772 ;
  LAYER M2 ;
        RECT 12.044 9.676 14.516 9.708 ;
  LAYER M2 ;
        RECT 12.044 9.612 14.516 9.644 ;
  LAYER M2 ;
        RECT 12.044 9.548 14.516 9.58 ;
  LAYER M2 ;
        RECT 12.044 9.484 14.516 9.516 ;
  LAYER M2 ;
        RECT 12.044 9.42 14.516 9.452 ;
  LAYER M2 ;
        RECT 12.044 9.356 14.516 9.388 ;
  LAYER M2 ;
        RECT 12.044 9.292 14.516 9.324 ;
  LAYER M2 ;
        RECT 12.044 9.228 14.516 9.26 ;
  LAYER M2 ;
        RECT 12.044 9.164 14.516 9.196 ;
  LAYER M2 ;
        RECT 12.044 9.1 14.516 9.132 ;
  LAYER M2 ;
        RECT 12.044 9.036 14.516 9.068 ;
  LAYER M2 ;
        RECT 12.044 8.972 14.516 9.004 ;
  LAYER M2 ;
        RECT 12.044 8.908 14.516 8.94 ;
  LAYER M2 ;
        RECT 12.044 8.844 14.516 8.876 ;
  LAYER M2 ;
        RECT 12.044 8.78 14.516 8.812 ;
  LAYER M2 ;
        RECT 12.044 8.716 14.516 8.748 ;
  LAYER M2 ;
        RECT 12.044 8.652 14.516 8.684 ;
  LAYER M2 ;
        RECT 12.044 8.588 14.516 8.62 ;
  LAYER M2 ;
        RECT 12.044 8.524 14.516 8.556 ;
  LAYER M2 ;
        RECT 12.044 8.46 14.516 8.492 ;
  LAYER M2 ;
        RECT 12.044 8.396 14.516 8.428 ;
  LAYER M2 ;
        RECT 12.044 8.332 14.516 8.364 ;
  LAYER M2 ;
        RECT 12.044 8.268 14.516 8.3 ;
  LAYER M2 ;
        RECT 12.044 8.204 14.516 8.236 ;
  LAYER M2 ;
        RECT 12.044 8.14 14.516 8.172 ;
  LAYER M2 ;
        RECT 12.044 8.076 14.516 8.108 ;
  LAYER M2 ;
        RECT 12.044 8.012 14.516 8.044 ;
  LAYER M3 ;
        RECT 14.464 7.86 14.496 10.368 ;
  LAYER M3 ;
        RECT 14.4 7.86 14.432 10.368 ;
  LAYER M3 ;
        RECT 14.336 7.86 14.368 10.368 ;
  LAYER M3 ;
        RECT 14.272 7.86 14.304 10.368 ;
  LAYER M3 ;
        RECT 14.208 7.86 14.24 10.368 ;
  LAYER M3 ;
        RECT 14.144 7.86 14.176 10.368 ;
  LAYER M3 ;
        RECT 14.08 7.86 14.112 10.368 ;
  LAYER M3 ;
        RECT 14.016 7.86 14.048 10.368 ;
  LAYER M3 ;
        RECT 13.952 7.86 13.984 10.368 ;
  LAYER M3 ;
        RECT 13.888 7.86 13.92 10.368 ;
  LAYER M3 ;
        RECT 13.824 7.86 13.856 10.368 ;
  LAYER M3 ;
        RECT 13.76 7.86 13.792 10.368 ;
  LAYER M3 ;
        RECT 13.696 7.86 13.728 10.368 ;
  LAYER M3 ;
        RECT 13.632 7.86 13.664 10.368 ;
  LAYER M3 ;
        RECT 13.568 7.86 13.6 10.368 ;
  LAYER M3 ;
        RECT 13.504 7.86 13.536 10.368 ;
  LAYER M3 ;
        RECT 13.44 7.86 13.472 10.368 ;
  LAYER M3 ;
        RECT 13.376 7.86 13.408 10.368 ;
  LAYER M3 ;
        RECT 13.312 7.86 13.344 10.368 ;
  LAYER M3 ;
        RECT 13.248 7.86 13.28 10.368 ;
  LAYER M3 ;
        RECT 13.184 7.86 13.216 10.368 ;
  LAYER M3 ;
        RECT 13.12 7.86 13.152 10.368 ;
  LAYER M3 ;
        RECT 13.056 7.86 13.088 10.368 ;
  LAYER M3 ;
        RECT 12.992 7.86 13.024 10.368 ;
  LAYER M3 ;
        RECT 12.928 7.86 12.96 10.368 ;
  LAYER M3 ;
        RECT 12.864 7.86 12.896 10.368 ;
  LAYER M3 ;
        RECT 12.8 7.86 12.832 10.368 ;
  LAYER M3 ;
        RECT 12.736 7.86 12.768 10.368 ;
  LAYER M3 ;
        RECT 12.672 7.86 12.704 10.368 ;
  LAYER M3 ;
        RECT 12.608 7.86 12.64 10.368 ;
  LAYER M3 ;
        RECT 12.544 7.86 12.576 10.368 ;
  LAYER M3 ;
        RECT 12.48 7.86 12.512 10.368 ;
  LAYER M3 ;
        RECT 12.416 7.86 12.448 10.368 ;
  LAYER M3 ;
        RECT 12.352 7.86 12.384 10.368 ;
  LAYER M3 ;
        RECT 12.288 7.86 12.32 10.368 ;
  LAYER M3 ;
        RECT 12.224 7.86 12.256 10.368 ;
  LAYER M3 ;
        RECT 12.16 7.86 12.192 10.368 ;
  LAYER M3 ;
        RECT 12.064 7.86 12.096 10.368 ;
  LAYER M1 ;
        RECT 14.479 7.896 14.481 10.332 ;
  LAYER M1 ;
        RECT 14.399 7.896 14.401 10.332 ;
  LAYER M1 ;
        RECT 14.319 7.896 14.321 10.332 ;
  LAYER M1 ;
        RECT 14.239 7.896 14.241 10.332 ;
  LAYER M1 ;
        RECT 14.159 7.896 14.161 10.332 ;
  LAYER M1 ;
        RECT 14.079 7.896 14.081 10.332 ;
  LAYER M1 ;
        RECT 13.999 7.896 14.001 10.332 ;
  LAYER M1 ;
        RECT 13.919 7.896 13.921 10.332 ;
  LAYER M1 ;
        RECT 13.839 7.896 13.841 10.332 ;
  LAYER M1 ;
        RECT 13.759 7.896 13.761 10.332 ;
  LAYER M1 ;
        RECT 13.679 7.896 13.681 10.332 ;
  LAYER M1 ;
        RECT 13.599 7.896 13.601 10.332 ;
  LAYER M1 ;
        RECT 13.519 7.896 13.521 10.332 ;
  LAYER M1 ;
        RECT 13.439 7.896 13.441 10.332 ;
  LAYER M1 ;
        RECT 13.359 7.896 13.361 10.332 ;
  LAYER M1 ;
        RECT 13.279 7.896 13.281 10.332 ;
  LAYER M1 ;
        RECT 13.199 7.896 13.201 10.332 ;
  LAYER M1 ;
        RECT 13.119 7.896 13.121 10.332 ;
  LAYER M1 ;
        RECT 13.039 7.896 13.041 10.332 ;
  LAYER M1 ;
        RECT 12.959 7.896 12.961 10.332 ;
  LAYER M1 ;
        RECT 12.879 7.896 12.881 10.332 ;
  LAYER M1 ;
        RECT 12.799 7.896 12.801 10.332 ;
  LAYER M1 ;
        RECT 12.719 7.896 12.721 10.332 ;
  LAYER M1 ;
        RECT 12.639 7.896 12.641 10.332 ;
  LAYER M1 ;
        RECT 12.559 7.896 12.561 10.332 ;
  LAYER M1 ;
        RECT 12.479 7.896 12.481 10.332 ;
  LAYER M1 ;
        RECT 12.399 7.896 12.401 10.332 ;
  LAYER M1 ;
        RECT 12.319 7.896 12.321 10.332 ;
  LAYER M1 ;
        RECT 12.239 7.896 12.241 10.332 ;
  LAYER M1 ;
        RECT 12.159 7.896 12.161 10.332 ;
  LAYER M2 ;
        RECT 12.08 10.331 14.48 10.333 ;
  LAYER M2 ;
        RECT 12.08 10.247 14.48 10.249 ;
  LAYER M2 ;
        RECT 12.08 10.163 14.48 10.165 ;
  LAYER M2 ;
        RECT 12.08 10.079 14.48 10.081 ;
  LAYER M2 ;
        RECT 12.08 9.995 14.48 9.997 ;
  LAYER M2 ;
        RECT 12.08 9.911 14.48 9.913 ;
  LAYER M2 ;
        RECT 12.08 9.827 14.48 9.829 ;
  LAYER M2 ;
        RECT 12.08 9.743 14.48 9.745 ;
  LAYER M2 ;
        RECT 12.08 9.659 14.48 9.661 ;
  LAYER M2 ;
        RECT 12.08 9.575 14.48 9.577 ;
  LAYER M2 ;
        RECT 12.08 9.491 14.48 9.493 ;
  LAYER M2 ;
        RECT 12.08 9.407 14.48 9.409 ;
  LAYER M2 ;
        RECT 12.08 9.3235 14.48 9.3255 ;
  LAYER M2 ;
        RECT 12.08 9.239 14.48 9.241 ;
  LAYER M2 ;
        RECT 12.08 9.155 14.48 9.157 ;
  LAYER M2 ;
        RECT 12.08 9.071 14.48 9.073 ;
  LAYER M2 ;
        RECT 12.08 8.987 14.48 8.989 ;
  LAYER M2 ;
        RECT 12.08 8.903 14.48 8.905 ;
  LAYER M2 ;
        RECT 12.08 8.819 14.48 8.821 ;
  LAYER M2 ;
        RECT 12.08 8.735 14.48 8.737 ;
  LAYER M2 ;
        RECT 12.08 8.651 14.48 8.653 ;
  LAYER M2 ;
        RECT 12.08 8.567 14.48 8.569 ;
  LAYER M2 ;
        RECT 12.08 8.483 14.48 8.485 ;
  LAYER M2 ;
        RECT 12.08 8.399 14.48 8.401 ;
  LAYER M2 ;
        RECT 12.08 8.315 14.48 8.317 ;
  LAYER M2 ;
        RECT 12.08 8.231 14.48 8.233 ;
  LAYER M2 ;
        RECT 12.08 8.147 14.48 8.149 ;
  LAYER M2 ;
        RECT 12.08 8.063 14.48 8.065 ;
  LAYER M2 ;
        RECT 12.08 7.979 14.48 7.981 ;
  LAYER M1 ;
        RECT 14.464 4.92 14.496 7.428 ;
  LAYER M1 ;
        RECT 14.4 4.92 14.432 7.428 ;
  LAYER M1 ;
        RECT 14.336 4.92 14.368 7.428 ;
  LAYER M1 ;
        RECT 14.272 4.92 14.304 7.428 ;
  LAYER M1 ;
        RECT 14.208 4.92 14.24 7.428 ;
  LAYER M1 ;
        RECT 14.144 4.92 14.176 7.428 ;
  LAYER M1 ;
        RECT 14.08 4.92 14.112 7.428 ;
  LAYER M1 ;
        RECT 14.016 4.92 14.048 7.428 ;
  LAYER M1 ;
        RECT 13.952 4.92 13.984 7.428 ;
  LAYER M1 ;
        RECT 13.888 4.92 13.92 7.428 ;
  LAYER M1 ;
        RECT 13.824 4.92 13.856 7.428 ;
  LAYER M1 ;
        RECT 13.76 4.92 13.792 7.428 ;
  LAYER M1 ;
        RECT 13.696 4.92 13.728 7.428 ;
  LAYER M1 ;
        RECT 13.632 4.92 13.664 7.428 ;
  LAYER M1 ;
        RECT 13.568 4.92 13.6 7.428 ;
  LAYER M1 ;
        RECT 13.504 4.92 13.536 7.428 ;
  LAYER M1 ;
        RECT 13.44 4.92 13.472 7.428 ;
  LAYER M1 ;
        RECT 13.376 4.92 13.408 7.428 ;
  LAYER M1 ;
        RECT 13.312 4.92 13.344 7.428 ;
  LAYER M1 ;
        RECT 13.248 4.92 13.28 7.428 ;
  LAYER M1 ;
        RECT 13.184 4.92 13.216 7.428 ;
  LAYER M1 ;
        RECT 13.12 4.92 13.152 7.428 ;
  LAYER M1 ;
        RECT 13.056 4.92 13.088 7.428 ;
  LAYER M1 ;
        RECT 12.992 4.92 13.024 7.428 ;
  LAYER M1 ;
        RECT 12.928 4.92 12.96 7.428 ;
  LAYER M1 ;
        RECT 12.864 4.92 12.896 7.428 ;
  LAYER M1 ;
        RECT 12.8 4.92 12.832 7.428 ;
  LAYER M1 ;
        RECT 12.736 4.92 12.768 7.428 ;
  LAYER M1 ;
        RECT 12.672 4.92 12.704 7.428 ;
  LAYER M1 ;
        RECT 12.608 4.92 12.64 7.428 ;
  LAYER M1 ;
        RECT 12.544 4.92 12.576 7.428 ;
  LAYER M1 ;
        RECT 12.48 4.92 12.512 7.428 ;
  LAYER M1 ;
        RECT 12.416 4.92 12.448 7.428 ;
  LAYER M1 ;
        RECT 12.352 4.92 12.384 7.428 ;
  LAYER M1 ;
        RECT 12.288 4.92 12.32 7.428 ;
  LAYER M1 ;
        RECT 12.224 4.92 12.256 7.428 ;
  LAYER M1 ;
        RECT 12.16 4.92 12.192 7.428 ;
  LAYER M2 ;
        RECT 12.044 7.312 14.516 7.344 ;
  LAYER M2 ;
        RECT 12.044 7.248 14.516 7.28 ;
  LAYER M2 ;
        RECT 12.044 7.184 14.516 7.216 ;
  LAYER M2 ;
        RECT 12.044 7.12 14.516 7.152 ;
  LAYER M2 ;
        RECT 12.044 7.056 14.516 7.088 ;
  LAYER M2 ;
        RECT 12.044 6.992 14.516 7.024 ;
  LAYER M2 ;
        RECT 12.044 6.928 14.516 6.96 ;
  LAYER M2 ;
        RECT 12.044 6.864 14.516 6.896 ;
  LAYER M2 ;
        RECT 12.044 6.8 14.516 6.832 ;
  LAYER M2 ;
        RECT 12.044 6.736 14.516 6.768 ;
  LAYER M2 ;
        RECT 12.044 6.672 14.516 6.704 ;
  LAYER M2 ;
        RECT 12.044 6.608 14.516 6.64 ;
  LAYER M2 ;
        RECT 12.044 6.544 14.516 6.576 ;
  LAYER M2 ;
        RECT 12.044 6.48 14.516 6.512 ;
  LAYER M2 ;
        RECT 12.044 6.416 14.516 6.448 ;
  LAYER M2 ;
        RECT 12.044 6.352 14.516 6.384 ;
  LAYER M2 ;
        RECT 12.044 6.288 14.516 6.32 ;
  LAYER M2 ;
        RECT 12.044 6.224 14.516 6.256 ;
  LAYER M2 ;
        RECT 12.044 6.16 14.516 6.192 ;
  LAYER M2 ;
        RECT 12.044 6.096 14.516 6.128 ;
  LAYER M2 ;
        RECT 12.044 6.032 14.516 6.064 ;
  LAYER M2 ;
        RECT 12.044 5.968 14.516 6 ;
  LAYER M2 ;
        RECT 12.044 5.904 14.516 5.936 ;
  LAYER M2 ;
        RECT 12.044 5.84 14.516 5.872 ;
  LAYER M2 ;
        RECT 12.044 5.776 14.516 5.808 ;
  LAYER M2 ;
        RECT 12.044 5.712 14.516 5.744 ;
  LAYER M2 ;
        RECT 12.044 5.648 14.516 5.68 ;
  LAYER M2 ;
        RECT 12.044 5.584 14.516 5.616 ;
  LAYER M2 ;
        RECT 12.044 5.52 14.516 5.552 ;
  LAYER M2 ;
        RECT 12.044 5.456 14.516 5.488 ;
  LAYER M2 ;
        RECT 12.044 5.392 14.516 5.424 ;
  LAYER M2 ;
        RECT 12.044 5.328 14.516 5.36 ;
  LAYER M2 ;
        RECT 12.044 5.264 14.516 5.296 ;
  LAYER M2 ;
        RECT 12.044 5.2 14.516 5.232 ;
  LAYER M2 ;
        RECT 12.044 5.136 14.516 5.168 ;
  LAYER M2 ;
        RECT 12.044 5.072 14.516 5.104 ;
  LAYER M3 ;
        RECT 14.464 4.92 14.496 7.428 ;
  LAYER M3 ;
        RECT 14.4 4.92 14.432 7.428 ;
  LAYER M3 ;
        RECT 14.336 4.92 14.368 7.428 ;
  LAYER M3 ;
        RECT 14.272 4.92 14.304 7.428 ;
  LAYER M3 ;
        RECT 14.208 4.92 14.24 7.428 ;
  LAYER M3 ;
        RECT 14.144 4.92 14.176 7.428 ;
  LAYER M3 ;
        RECT 14.08 4.92 14.112 7.428 ;
  LAYER M3 ;
        RECT 14.016 4.92 14.048 7.428 ;
  LAYER M3 ;
        RECT 13.952 4.92 13.984 7.428 ;
  LAYER M3 ;
        RECT 13.888 4.92 13.92 7.428 ;
  LAYER M3 ;
        RECT 13.824 4.92 13.856 7.428 ;
  LAYER M3 ;
        RECT 13.76 4.92 13.792 7.428 ;
  LAYER M3 ;
        RECT 13.696 4.92 13.728 7.428 ;
  LAYER M3 ;
        RECT 13.632 4.92 13.664 7.428 ;
  LAYER M3 ;
        RECT 13.568 4.92 13.6 7.428 ;
  LAYER M3 ;
        RECT 13.504 4.92 13.536 7.428 ;
  LAYER M3 ;
        RECT 13.44 4.92 13.472 7.428 ;
  LAYER M3 ;
        RECT 13.376 4.92 13.408 7.428 ;
  LAYER M3 ;
        RECT 13.312 4.92 13.344 7.428 ;
  LAYER M3 ;
        RECT 13.248 4.92 13.28 7.428 ;
  LAYER M3 ;
        RECT 13.184 4.92 13.216 7.428 ;
  LAYER M3 ;
        RECT 13.12 4.92 13.152 7.428 ;
  LAYER M3 ;
        RECT 13.056 4.92 13.088 7.428 ;
  LAYER M3 ;
        RECT 12.992 4.92 13.024 7.428 ;
  LAYER M3 ;
        RECT 12.928 4.92 12.96 7.428 ;
  LAYER M3 ;
        RECT 12.864 4.92 12.896 7.428 ;
  LAYER M3 ;
        RECT 12.8 4.92 12.832 7.428 ;
  LAYER M3 ;
        RECT 12.736 4.92 12.768 7.428 ;
  LAYER M3 ;
        RECT 12.672 4.92 12.704 7.428 ;
  LAYER M3 ;
        RECT 12.608 4.92 12.64 7.428 ;
  LAYER M3 ;
        RECT 12.544 4.92 12.576 7.428 ;
  LAYER M3 ;
        RECT 12.48 4.92 12.512 7.428 ;
  LAYER M3 ;
        RECT 12.416 4.92 12.448 7.428 ;
  LAYER M3 ;
        RECT 12.352 4.92 12.384 7.428 ;
  LAYER M3 ;
        RECT 12.288 4.92 12.32 7.428 ;
  LAYER M3 ;
        RECT 12.224 4.92 12.256 7.428 ;
  LAYER M3 ;
        RECT 12.16 4.92 12.192 7.428 ;
  LAYER M3 ;
        RECT 12.064 4.92 12.096 7.428 ;
  LAYER M1 ;
        RECT 14.479 4.956 14.481 7.392 ;
  LAYER M1 ;
        RECT 14.399 4.956 14.401 7.392 ;
  LAYER M1 ;
        RECT 14.319 4.956 14.321 7.392 ;
  LAYER M1 ;
        RECT 14.239 4.956 14.241 7.392 ;
  LAYER M1 ;
        RECT 14.159 4.956 14.161 7.392 ;
  LAYER M1 ;
        RECT 14.079 4.956 14.081 7.392 ;
  LAYER M1 ;
        RECT 13.999 4.956 14.001 7.392 ;
  LAYER M1 ;
        RECT 13.919 4.956 13.921 7.392 ;
  LAYER M1 ;
        RECT 13.839 4.956 13.841 7.392 ;
  LAYER M1 ;
        RECT 13.759 4.956 13.761 7.392 ;
  LAYER M1 ;
        RECT 13.679 4.956 13.681 7.392 ;
  LAYER M1 ;
        RECT 13.599 4.956 13.601 7.392 ;
  LAYER M1 ;
        RECT 13.519 4.956 13.521 7.392 ;
  LAYER M1 ;
        RECT 13.439 4.956 13.441 7.392 ;
  LAYER M1 ;
        RECT 13.359 4.956 13.361 7.392 ;
  LAYER M1 ;
        RECT 13.279 4.956 13.281 7.392 ;
  LAYER M1 ;
        RECT 13.199 4.956 13.201 7.392 ;
  LAYER M1 ;
        RECT 13.119 4.956 13.121 7.392 ;
  LAYER M1 ;
        RECT 13.039 4.956 13.041 7.392 ;
  LAYER M1 ;
        RECT 12.959 4.956 12.961 7.392 ;
  LAYER M1 ;
        RECT 12.879 4.956 12.881 7.392 ;
  LAYER M1 ;
        RECT 12.799 4.956 12.801 7.392 ;
  LAYER M1 ;
        RECT 12.719 4.956 12.721 7.392 ;
  LAYER M1 ;
        RECT 12.639 4.956 12.641 7.392 ;
  LAYER M1 ;
        RECT 12.559 4.956 12.561 7.392 ;
  LAYER M1 ;
        RECT 12.479 4.956 12.481 7.392 ;
  LAYER M1 ;
        RECT 12.399 4.956 12.401 7.392 ;
  LAYER M1 ;
        RECT 12.319 4.956 12.321 7.392 ;
  LAYER M1 ;
        RECT 12.239 4.956 12.241 7.392 ;
  LAYER M1 ;
        RECT 12.159 4.956 12.161 7.392 ;
  LAYER M2 ;
        RECT 12.08 7.391 14.48 7.393 ;
  LAYER M2 ;
        RECT 12.08 7.307 14.48 7.309 ;
  LAYER M2 ;
        RECT 12.08 7.223 14.48 7.225 ;
  LAYER M2 ;
        RECT 12.08 7.139 14.48 7.141 ;
  LAYER M2 ;
        RECT 12.08 7.055 14.48 7.057 ;
  LAYER M2 ;
        RECT 12.08 6.971 14.48 6.973 ;
  LAYER M2 ;
        RECT 12.08 6.887 14.48 6.889 ;
  LAYER M2 ;
        RECT 12.08 6.803 14.48 6.805 ;
  LAYER M2 ;
        RECT 12.08 6.719 14.48 6.721 ;
  LAYER M2 ;
        RECT 12.08 6.635 14.48 6.637 ;
  LAYER M2 ;
        RECT 12.08 6.551 14.48 6.553 ;
  LAYER M2 ;
        RECT 12.08 6.467 14.48 6.469 ;
  LAYER M2 ;
        RECT 12.08 6.3835 14.48 6.3855 ;
  LAYER M2 ;
        RECT 12.08 6.299 14.48 6.301 ;
  LAYER M2 ;
        RECT 12.08 6.215 14.48 6.217 ;
  LAYER M2 ;
        RECT 12.08 6.131 14.48 6.133 ;
  LAYER M2 ;
        RECT 12.08 6.047 14.48 6.049 ;
  LAYER M2 ;
        RECT 12.08 5.963 14.48 5.965 ;
  LAYER M2 ;
        RECT 12.08 5.879 14.48 5.881 ;
  LAYER M2 ;
        RECT 12.08 5.795 14.48 5.797 ;
  LAYER M2 ;
        RECT 12.08 5.711 14.48 5.713 ;
  LAYER M2 ;
        RECT 12.08 5.627 14.48 5.629 ;
  LAYER M2 ;
        RECT 12.08 5.543 14.48 5.545 ;
  LAYER M2 ;
        RECT 12.08 5.459 14.48 5.461 ;
  LAYER M2 ;
        RECT 12.08 5.375 14.48 5.377 ;
  LAYER M2 ;
        RECT 12.08 5.291 14.48 5.293 ;
  LAYER M2 ;
        RECT 12.08 5.207 14.48 5.209 ;
  LAYER M2 ;
        RECT 12.08 5.123 14.48 5.125 ;
  LAYER M2 ;
        RECT 12.08 5.039 14.48 5.041 ;
  LAYER M1 ;
        RECT 14.464 1.98 14.496 4.488 ;
  LAYER M1 ;
        RECT 14.4 1.98 14.432 4.488 ;
  LAYER M1 ;
        RECT 14.336 1.98 14.368 4.488 ;
  LAYER M1 ;
        RECT 14.272 1.98 14.304 4.488 ;
  LAYER M1 ;
        RECT 14.208 1.98 14.24 4.488 ;
  LAYER M1 ;
        RECT 14.144 1.98 14.176 4.488 ;
  LAYER M1 ;
        RECT 14.08 1.98 14.112 4.488 ;
  LAYER M1 ;
        RECT 14.016 1.98 14.048 4.488 ;
  LAYER M1 ;
        RECT 13.952 1.98 13.984 4.488 ;
  LAYER M1 ;
        RECT 13.888 1.98 13.92 4.488 ;
  LAYER M1 ;
        RECT 13.824 1.98 13.856 4.488 ;
  LAYER M1 ;
        RECT 13.76 1.98 13.792 4.488 ;
  LAYER M1 ;
        RECT 13.696 1.98 13.728 4.488 ;
  LAYER M1 ;
        RECT 13.632 1.98 13.664 4.488 ;
  LAYER M1 ;
        RECT 13.568 1.98 13.6 4.488 ;
  LAYER M1 ;
        RECT 13.504 1.98 13.536 4.488 ;
  LAYER M1 ;
        RECT 13.44 1.98 13.472 4.488 ;
  LAYER M1 ;
        RECT 13.376 1.98 13.408 4.488 ;
  LAYER M1 ;
        RECT 13.312 1.98 13.344 4.488 ;
  LAYER M1 ;
        RECT 13.248 1.98 13.28 4.488 ;
  LAYER M1 ;
        RECT 13.184 1.98 13.216 4.488 ;
  LAYER M1 ;
        RECT 13.12 1.98 13.152 4.488 ;
  LAYER M1 ;
        RECT 13.056 1.98 13.088 4.488 ;
  LAYER M1 ;
        RECT 12.992 1.98 13.024 4.488 ;
  LAYER M1 ;
        RECT 12.928 1.98 12.96 4.488 ;
  LAYER M1 ;
        RECT 12.864 1.98 12.896 4.488 ;
  LAYER M1 ;
        RECT 12.8 1.98 12.832 4.488 ;
  LAYER M1 ;
        RECT 12.736 1.98 12.768 4.488 ;
  LAYER M1 ;
        RECT 12.672 1.98 12.704 4.488 ;
  LAYER M1 ;
        RECT 12.608 1.98 12.64 4.488 ;
  LAYER M1 ;
        RECT 12.544 1.98 12.576 4.488 ;
  LAYER M1 ;
        RECT 12.48 1.98 12.512 4.488 ;
  LAYER M1 ;
        RECT 12.416 1.98 12.448 4.488 ;
  LAYER M1 ;
        RECT 12.352 1.98 12.384 4.488 ;
  LAYER M1 ;
        RECT 12.288 1.98 12.32 4.488 ;
  LAYER M1 ;
        RECT 12.224 1.98 12.256 4.488 ;
  LAYER M1 ;
        RECT 12.16 1.98 12.192 4.488 ;
  LAYER M2 ;
        RECT 12.044 4.372 14.516 4.404 ;
  LAYER M2 ;
        RECT 12.044 4.308 14.516 4.34 ;
  LAYER M2 ;
        RECT 12.044 4.244 14.516 4.276 ;
  LAYER M2 ;
        RECT 12.044 4.18 14.516 4.212 ;
  LAYER M2 ;
        RECT 12.044 4.116 14.516 4.148 ;
  LAYER M2 ;
        RECT 12.044 4.052 14.516 4.084 ;
  LAYER M2 ;
        RECT 12.044 3.988 14.516 4.02 ;
  LAYER M2 ;
        RECT 12.044 3.924 14.516 3.956 ;
  LAYER M2 ;
        RECT 12.044 3.86 14.516 3.892 ;
  LAYER M2 ;
        RECT 12.044 3.796 14.516 3.828 ;
  LAYER M2 ;
        RECT 12.044 3.732 14.516 3.764 ;
  LAYER M2 ;
        RECT 12.044 3.668 14.516 3.7 ;
  LAYER M2 ;
        RECT 12.044 3.604 14.516 3.636 ;
  LAYER M2 ;
        RECT 12.044 3.54 14.516 3.572 ;
  LAYER M2 ;
        RECT 12.044 3.476 14.516 3.508 ;
  LAYER M2 ;
        RECT 12.044 3.412 14.516 3.444 ;
  LAYER M2 ;
        RECT 12.044 3.348 14.516 3.38 ;
  LAYER M2 ;
        RECT 12.044 3.284 14.516 3.316 ;
  LAYER M2 ;
        RECT 12.044 3.22 14.516 3.252 ;
  LAYER M2 ;
        RECT 12.044 3.156 14.516 3.188 ;
  LAYER M2 ;
        RECT 12.044 3.092 14.516 3.124 ;
  LAYER M2 ;
        RECT 12.044 3.028 14.516 3.06 ;
  LAYER M2 ;
        RECT 12.044 2.964 14.516 2.996 ;
  LAYER M2 ;
        RECT 12.044 2.9 14.516 2.932 ;
  LAYER M2 ;
        RECT 12.044 2.836 14.516 2.868 ;
  LAYER M2 ;
        RECT 12.044 2.772 14.516 2.804 ;
  LAYER M2 ;
        RECT 12.044 2.708 14.516 2.74 ;
  LAYER M2 ;
        RECT 12.044 2.644 14.516 2.676 ;
  LAYER M2 ;
        RECT 12.044 2.58 14.516 2.612 ;
  LAYER M2 ;
        RECT 12.044 2.516 14.516 2.548 ;
  LAYER M2 ;
        RECT 12.044 2.452 14.516 2.484 ;
  LAYER M2 ;
        RECT 12.044 2.388 14.516 2.42 ;
  LAYER M2 ;
        RECT 12.044 2.324 14.516 2.356 ;
  LAYER M2 ;
        RECT 12.044 2.26 14.516 2.292 ;
  LAYER M2 ;
        RECT 12.044 2.196 14.516 2.228 ;
  LAYER M2 ;
        RECT 12.044 2.132 14.516 2.164 ;
  LAYER M3 ;
        RECT 14.464 1.98 14.496 4.488 ;
  LAYER M3 ;
        RECT 14.4 1.98 14.432 4.488 ;
  LAYER M3 ;
        RECT 14.336 1.98 14.368 4.488 ;
  LAYER M3 ;
        RECT 14.272 1.98 14.304 4.488 ;
  LAYER M3 ;
        RECT 14.208 1.98 14.24 4.488 ;
  LAYER M3 ;
        RECT 14.144 1.98 14.176 4.488 ;
  LAYER M3 ;
        RECT 14.08 1.98 14.112 4.488 ;
  LAYER M3 ;
        RECT 14.016 1.98 14.048 4.488 ;
  LAYER M3 ;
        RECT 13.952 1.98 13.984 4.488 ;
  LAYER M3 ;
        RECT 13.888 1.98 13.92 4.488 ;
  LAYER M3 ;
        RECT 13.824 1.98 13.856 4.488 ;
  LAYER M3 ;
        RECT 13.76 1.98 13.792 4.488 ;
  LAYER M3 ;
        RECT 13.696 1.98 13.728 4.488 ;
  LAYER M3 ;
        RECT 13.632 1.98 13.664 4.488 ;
  LAYER M3 ;
        RECT 13.568 1.98 13.6 4.488 ;
  LAYER M3 ;
        RECT 13.504 1.98 13.536 4.488 ;
  LAYER M3 ;
        RECT 13.44 1.98 13.472 4.488 ;
  LAYER M3 ;
        RECT 13.376 1.98 13.408 4.488 ;
  LAYER M3 ;
        RECT 13.312 1.98 13.344 4.488 ;
  LAYER M3 ;
        RECT 13.248 1.98 13.28 4.488 ;
  LAYER M3 ;
        RECT 13.184 1.98 13.216 4.488 ;
  LAYER M3 ;
        RECT 13.12 1.98 13.152 4.488 ;
  LAYER M3 ;
        RECT 13.056 1.98 13.088 4.488 ;
  LAYER M3 ;
        RECT 12.992 1.98 13.024 4.488 ;
  LAYER M3 ;
        RECT 12.928 1.98 12.96 4.488 ;
  LAYER M3 ;
        RECT 12.864 1.98 12.896 4.488 ;
  LAYER M3 ;
        RECT 12.8 1.98 12.832 4.488 ;
  LAYER M3 ;
        RECT 12.736 1.98 12.768 4.488 ;
  LAYER M3 ;
        RECT 12.672 1.98 12.704 4.488 ;
  LAYER M3 ;
        RECT 12.608 1.98 12.64 4.488 ;
  LAYER M3 ;
        RECT 12.544 1.98 12.576 4.488 ;
  LAYER M3 ;
        RECT 12.48 1.98 12.512 4.488 ;
  LAYER M3 ;
        RECT 12.416 1.98 12.448 4.488 ;
  LAYER M3 ;
        RECT 12.352 1.98 12.384 4.488 ;
  LAYER M3 ;
        RECT 12.288 1.98 12.32 4.488 ;
  LAYER M3 ;
        RECT 12.224 1.98 12.256 4.488 ;
  LAYER M3 ;
        RECT 12.16 1.98 12.192 4.488 ;
  LAYER M3 ;
        RECT 12.064 1.98 12.096 4.488 ;
  LAYER M1 ;
        RECT 14.479 2.016 14.481 4.452 ;
  LAYER M1 ;
        RECT 14.399 2.016 14.401 4.452 ;
  LAYER M1 ;
        RECT 14.319 2.016 14.321 4.452 ;
  LAYER M1 ;
        RECT 14.239 2.016 14.241 4.452 ;
  LAYER M1 ;
        RECT 14.159 2.016 14.161 4.452 ;
  LAYER M1 ;
        RECT 14.079 2.016 14.081 4.452 ;
  LAYER M1 ;
        RECT 13.999 2.016 14.001 4.452 ;
  LAYER M1 ;
        RECT 13.919 2.016 13.921 4.452 ;
  LAYER M1 ;
        RECT 13.839 2.016 13.841 4.452 ;
  LAYER M1 ;
        RECT 13.759 2.016 13.761 4.452 ;
  LAYER M1 ;
        RECT 13.679 2.016 13.681 4.452 ;
  LAYER M1 ;
        RECT 13.599 2.016 13.601 4.452 ;
  LAYER M1 ;
        RECT 13.519 2.016 13.521 4.452 ;
  LAYER M1 ;
        RECT 13.439 2.016 13.441 4.452 ;
  LAYER M1 ;
        RECT 13.359 2.016 13.361 4.452 ;
  LAYER M1 ;
        RECT 13.279 2.016 13.281 4.452 ;
  LAYER M1 ;
        RECT 13.199 2.016 13.201 4.452 ;
  LAYER M1 ;
        RECT 13.119 2.016 13.121 4.452 ;
  LAYER M1 ;
        RECT 13.039 2.016 13.041 4.452 ;
  LAYER M1 ;
        RECT 12.959 2.016 12.961 4.452 ;
  LAYER M1 ;
        RECT 12.879 2.016 12.881 4.452 ;
  LAYER M1 ;
        RECT 12.799 2.016 12.801 4.452 ;
  LAYER M1 ;
        RECT 12.719 2.016 12.721 4.452 ;
  LAYER M1 ;
        RECT 12.639 2.016 12.641 4.452 ;
  LAYER M1 ;
        RECT 12.559 2.016 12.561 4.452 ;
  LAYER M1 ;
        RECT 12.479 2.016 12.481 4.452 ;
  LAYER M1 ;
        RECT 12.399 2.016 12.401 4.452 ;
  LAYER M1 ;
        RECT 12.319 2.016 12.321 4.452 ;
  LAYER M1 ;
        RECT 12.239 2.016 12.241 4.452 ;
  LAYER M1 ;
        RECT 12.159 2.016 12.161 4.452 ;
  LAYER M2 ;
        RECT 12.08 4.451 14.48 4.453 ;
  LAYER M2 ;
        RECT 12.08 4.367 14.48 4.369 ;
  LAYER M2 ;
        RECT 12.08 4.283 14.48 4.285 ;
  LAYER M2 ;
        RECT 12.08 4.199 14.48 4.201 ;
  LAYER M2 ;
        RECT 12.08 4.115 14.48 4.117 ;
  LAYER M2 ;
        RECT 12.08 4.031 14.48 4.033 ;
  LAYER M2 ;
        RECT 12.08 3.947 14.48 3.949 ;
  LAYER M2 ;
        RECT 12.08 3.863 14.48 3.865 ;
  LAYER M2 ;
        RECT 12.08 3.779 14.48 3.781 ;
  LAYER M2 ;
        RECT 12.08 3.695 14.48 3.697 ;
  LAYER M2 ;
        RECT 12.08 3.611 14.48 3.613 ;
  LAYER M2 ;
        RECT 12.08 3.527 14.48 3.529 ;
  LAYER M2 ;
        RECT 12.08 3.4435 14.48 3.4455 ;
  LAYER M2 ;
        RECT 12.08 3.359 14.48 3.361 ;
  LAYER M2 ;
        RECT 12.08 3.275 14.48 3.277 ;
  LAYER M2 ;
        RECT 12.08 3.191 14.48 3.193 ;
  LAYER M2 ;
        RECT 12.08 3.107 14.48 3.109 ;
  LAYER M2 ;
        RECT 12.08 3.023 14.48 3.025 ;
  LAYER M2 ;
        RECT 12.08 2.939 14.48 2.941 ;
  LAYER M2 ;
        RECT 12.08 2.855 14.48 2.857 ;
  LAYER M2 ;
        RECT 12.08 2.771 14.48 2.773 ;
  LAYER M2 ;
        RECT 12.08 2.687 14.48 2.689 ;
  LAYER M2 ;
        RECT 12.08 2.603 14.48 2.605 ;
  LAYER M2 ;
        RECT 12.08 2.519 14.48 2.521 ;
  LAYER M2 ;
        RECT 12.08 2.435 14.48 2.437 ;
  LAYER M2 ;
        RECT 12.08 2.351 14.48 2.353 ;
  LAYER M2 ;
        RECT 12.08 2.267 14.48 2.269 ;
  LAYER M2 ;
        RECT 12.08 2.183 14.48 2.185 ;
  LAYER M2 ;
        RECT 12.08 2.099 14.48 2.101 ;
  LAYER M1 ;
        RECT 11.584 13.74 11.616 16.248 ;
  LAYER M1 ;
        RECT 11.52 13.74 11.552 16.248 ;
  LAYER M1 ;
        RECT 11.456 13.74 11.488 16.248 ;
  LAYER M1 ;
        RECT 11.392 13.74 11.424 16.248 ;
  LAYER M1 ;
        RECT 11.328 13.74 11.36 16.248 ;
  LAYER M1 ;
        RECT 11.264 13.74 11.296 16.248 ;
  LAYER M1 ;
        RECT 11.2 13.74 11.232 16.248 ;
  LAYER M1 ;
        RECT 11.136 13.74 11.168 16.248 ;
  LAYER M1 ;
        RECT 11.072 13.74 11.104 16.248 ;
  LAYER M1 ;
        RECT 11.008 13.74 11.04 16.248 ;
  LAYER M1 ;
        RECT 10.944 13.74 10.976 16.248 ;
  LAYER M1 ;
        RECT 10.88 13.74 10.912 16.248 ;
  LAYER M1 ;
        RECT 10.816 13.74 10.848 16.248 ;
  LAYER M1 ;
        RECT 10.752 13.74 10.784 16.248 ;
  LAYER M1 ;
        RECT 10.688 13.74 10.72 16.248 ;
  LAYER M1 ;
        RECT 10.624 13.74 10.656 16.248 ;
  LAYER M1 ;
        RECT 10.56 13.74 10.592 16.248 ;
  LAYER M1 ;
        RECT 10.496 13.74 10.528 16.248 ;
  LAYER M1 ;
        RECT 10.432 13.74 10.464 16.248 ;
  LAYER M1 ;
        RECT 10.368 13.74 10.4 16.248 ;
  LAYER M1 ;
        RECT 10.304 13.74 10.336 16.248 ;
  LAYER M1 ;
        RECT 10.24 13.74 10.272 16.248 ;
  LAYER M1 ;
        RECT 10.176 13.74 10.208 16.248 ;
  LAYER M1 ;
        RECT 10.112 13.74 10.144 16.248 ;
  LAYER M1 ;
        RECT 10.048 13.74 10.08 16.248 ;
  LAYER M1 ;
        RECT 9.984 13.74 10.016 16.248 ;
  LAYER M1 ;
        RECT 9.92 13.74 9.952 16.248 ;
  LAYER M1 ;
        RECT 9.856 13.74 9.888 16.248 ;
  LAYER M1 ;
        RECT 9.792 13.74 9.824 16.248 ;
  LAYER M1 ;
        RECT 9.728 13.74 9.76 16.248 ;
  LAYER M1 ;
        RECT 9.664 13.74 9.696 16.248 ;
  LAYER M1 ;
        RECT 9.6 13.74 9.632 16.248 ;
  LAYER M1 ;
        RECT 9.536 13.74 9.568 16.248 ;
  LAYER M1 ;
        RECT 9.472 13.74 9.504 16.248 ;
  LAYER M1 ;
        RECT 9.408 13.74 9.44 16.248 ;
  LAYER M1 ;
        RECT 9.344 13.74 9.376 16.248 ;
  LAYER M1 ;
        RECT 9.28 13.74 9.312 16.248 ;
  LAYER M2 ;
        RECT 9.164 16.132 11.636 16.164 ;
  LAYER M2 ;
        RECT 9.164 16.068 11.636 16.1 ;
  LAYER M2 ;
        RECT 9.164 16.004 11.636 16.036 ;
  LAYER M2 ;
        RECT 9.164 15.94 11.636 15.972 ;
  LAYER M2 ;
        RECT 9.164 15.876 11.636 15.908 ;
  LAYER M2 ;
        RECT 9.164 15.812 11.636 15.844 ;
  LAYER M2 ;
        RECT 9.164 15.748 11.636 15.78 ;
  LAYER M2 ;
        RECT 9.164 15.684 11.636 15.716 ;
  LAYER M2 ;
        RECT 9.164 15.62 11.636 15.652 ;
  LAYER M2 ;
        RECT 9.164 15.556 11.636 15.588 ;
  LAYER M2 ;
        RECT 9.164 15.492 11.636 15.524 ;
  LAYER M2 ;
        RECT 9.164 15.428 11.636 15.46 ;
  LAYER M2 ;
        RECT 9.164 15.364 11.636 15.396 ;
  LAYER M2 ;
        RECT 9.164 15.3 11.636 15.332 ;
  LAYER M2 ;
        RECT 9.164 15.236 11.636 15.268 ;
  LAYER M2 ;
        RECT 9.164 15.172 11.636 15.204 ;
  LAYER M2 ;
        RECT 9.164 15.108 11.636 15.14 ;
  LAYER M2 ;
        RECT 9.164 15.044 11.636 15.076 ;
  LAYER M2 ;
        RECT 9.164 14.98 11.636 15.012 ;
  LAYER M2 ;
        RECT 9.164 14.916 11.636 14.948 ;
  LAYER M2 ;
        RECT 9.164 14.852 11.636 14.884 ;
  LAYER M2 ;
        RECT 9.164 14.788 11.636 14.82 ;
  LAYER M2 ;
        RECT 9.164 14.724 11.636 14.756 ;
  LAYER M2 ;
        RECT 9.164 14.66 11.636 14.692 ;
  LAYER M2 ;
        RECT 9.164 14.596 11.636 14.628 ;
  LAYER M2 ;
        RECT 9.164 14.532 11.636 14.564 ;
  LAYER M2 ;
        RECT 9.164 14.468 11.636 14.5 ;
  LAYER M2 ;
        RECT 9.164 14.404 11.636 14.436 ;
  LAYER M2 ;
        RECT 9.164 14.34 11.636 14.372 ;
  LAYER M2 ;
        RECT 9.164 14.276 11.636 14.308 ;
  LAYER M2 ;
        RECT 9.164 14.212 11.636 14.244 ;
  LAYER M2 ;
        RECT 9.164 14.148 11.636 14.18 ;
  LAYER M2 ;
        RECT 9.164 14.084 11.636 14.116 ;
  LAYER M2 ;
        RECT 9.164 14.02 11.636 14.052 ;
  LAYER M2 ;
        RECT 9.164 13.956 11.636 13.988 ;
  LAYER M2 ;
        RECT 9.164 13.892 11.636 13.924 ;
  LAYER M3 ;
        RECT 11.584 13.74 11.616 16.248 ;
  LAYER M3 ;
        RECT 11.52 13.74 11.552 16.248 ;
  LAYER M3 ;
        RECT 11.456 13.74 11.488 16.248 ;
  LAYER M3 ;
        RECT 11.392 13.74 11.424 16.248 ;
  LAYER M3 ;
        RECT 11.328 13.74 11.36 16.248 ;
  LAYER M3 ;
        RECT 11.264 13.74 11.296 16.248 ;
  LAYER M3 ;
        RECT 11.2 13.74 11.232 16.248 ;
  LAYER M3 ;
        RECT 11.136 13.74 11.168 16.248 ;
  LAYER M3 ;
        RECT 11.072 13.74 11.104 16.248 ;
  LAYER M3 ;
        RECT 11.008 13.74 11.04 16.248 ;
  LAYER M3 ;
        RECT 10.944 13.74 10.976 16.248 ;
  LAYER M3 ;
        RECT 10.88 13.74 10.912 16.248 ;
  LAYER M3 ;
        RECT 10.816 13.74 10.848 16.248 ;
  LAYER M3 ;
        RECT 10.752 13.74 10.784 16.248 ;
  LAYER M3 ;
        RECT 10.688 13.74 10.72 16.248 ;
  LAYER M3 ;
        RECT 10.624 13.74 10.656 16.248 ;
  LAYER M3 ;
        RECT 10.56 13.74 10.592 16.248 ;
  LAYER M3 ;
        RECT 10.496 13.74 10.528 16.248 ;
  LAYER M3 ;
        RECT 10.432 13.74 10.464 16.248 ;
  LAYER M3 ;
        RECT 10.368 13.74 10.4 16.248 ;
  LAYER M3 ;
        RECT 10.304 13.74 10.336 16.248 ;
  LAYER M3 ;
        RECT 10.24 13.74 10.272 16.248 ;
  LAYER M3 ;
        RECT 10.176 13.74 10.208 16.248 ;
  LAYER M3 ;
        RECT 10.112 13.74 10.144 16.248 ;
  LAYER M3 ;
        RECT 10.048 13.74 10.08 16.248 ;
  LAYER M3 ;
        RECT 9.984 13.74 10.016 16.248 ;
  LAYER M3 ;
        RECT 9.92 13.74 9.952 16.248 ;
  LAYER M3 ;
        RECT 9.856 13.74 9.888 16.248 ;
  LAYER M3 ;
        RECT 9.792 13.74 9.824 16.248 ;
  LAYER M3 ;
        RECT 9.728 13.74 9.76 16.248 ;
  LAYER M3 ;
        RECT 9.664 13.74 9.696 16.248 ;
  LAYER M3 ;
        RECT 9.6 13.74 9.632 16.248 ;
  LAYER M3 ;
        RECT 9.536 13.74 9.568 16.248 ;
  LAYER M3 ;
        RECT 9.472 13.74 9.504 16.248 ;
  LAYER M3 ;
        RECT 9.408 13.74 9.44 16.248 ;
  LAYER M3 ;
        RECT 9.344 13.74 9.376 16.248 ;
  LAYER M3 ;
        RECT 9.28 13.74 9.312 16.248 ;
  LAYER M3 ;
        RECT 9.184 13.74 9.216 16.248 ;
  LAYER M1 ;
        RECT 11.599 13.776 11.601 16.212 ;
  LAYER M1 ;
        RECT 11.519 13.776 11.521 16.212 ;
  LAYER M1 ;
        RECT 11.439 13.776 11.441 16.212 ;
  LAYER M1 ;
        RECT 11.359 13.776 11.361 16.212 ;
  LAYER M1 ;
        RECT 11.279 13.776 11.281 16.212 ;
  LAYER M1 ;
        RECT 11.199 13.776 11.201 16.212 ;
  LAYER M1 ;
        RECT 11.119 13.776 11.121 16.212 ;
  LAYER M1 ;
        RECT 11.039 13.776 11.041 16.212 ;
  LAYER M1 ;
        RECT 10.959 13.776 10.961 16.212 ;
  LAYER M1 ;
        RECT 10.879 13.776 10.881 16.212 ;
  LAYER M1 ;
        RECT 10.799 13.776 10.801 16.212 ;
  LAYER M1 ;
        RECT 10.719 13.776 10.721 16.212 ;
  LAYER M1 ;
        RECT 10.639 13.776 10.641 16.212 ;
  LAYER M1 ;
        RECT 10.559 13.776 10.561 16.212 ;
  LAYER M1 ;
        RECT 10.479 13.776 10.481 16.212 ;
  LAYER M1 ;
        RECT 10.399 13.776 10.401 16.212 ;
  LAYER M1 ;
        RECT 10.319 13.776 10.321 16.212 ;
  LAYER M1 ;
        RECT 10.239 13.776 10.241 16.212 ;
  LAYER M1 ;
        RECT 10.159 13.776 10.161 16.212 ;
  LAYER M1 ;
        RECT 10.079 13.776 10.081 16.212 ;
  LAYER M1 ;
        RECT 9.999 13.776 10.001 16.212 ;
  LAYER M1 ;
        RECT 9.919 13.776 9.921 16.212 ;
  LAYER M1 ;
        RECT 9.839 13.776 9.841 16.212 ;
  LAYER M1 ;
        RECT 9.759 13.776 9.761 16.212 ;
  LAYER M1 ;
        RECT 9.679 13.776 9.681 16.212 ;
  LAYER M1 ;
        RECT 9.599 13.776 9.601 16.212 ;
  LAYER M1 ;
        RECT 9.519 13.776 9.521 16.212 ;
  LAYER M1 ;
        RECT 9.439 13.776 9.441 16.212 ;
  LAYER M1 ;
        RECT 9.359 13.776 9.361 16.212 ;
  LAYER M1 ;
        RECT 9.279 13.776 9.281 16.212 ;
  LAYER M2 ;
        RECT 9.2 16.211 11.6 16.213 ;
  LAYER M2 ;
        RECT 9.2 16.127 11.6 16.129 ;
  LAYER M2 ;
        RECT 9.2 16.043 11.6 16.045 ;
  LAYER M2 ;
        RECT 9.2 15.959 11.6 15.961 ;
  LAYER M2 ;
        RECT 9.2 15.875 11.6 15.877 ;
  LAYER M2 ;
        RECT 9.2 15.791 11.6 15.793 ;
  LAYER M2 ;
        RECT 9.2 15.707 11.6 15.709 ;
  LAYER M2 ;
        RECT 9.2 15.623 11.6 15.625 ;
  LAYER M2 ;
        RECT 9.2 15.539 11.6 15.541 ;
  LAYER M2 ;
        RECT 9.2 15.455 11.6 15.457 ;
  LAYER M2 ;
        RECT 9.2 15.371 11.6 15.373 ;
  LAYER M2 ;
        RECT 9.2 15.287 11.6 15.289 ;
  LAYER M2 ;
        RECT 9.2 15.2035 11.6 15.2055 ;
  LAYER M2 ;
        RECT 9.2 15.119 11.6 15.121 ;
  LAYER M2 ;
        RECT 9.2 15.035 11.6 15.037 ;
  LAYER M2 ;
        RECT 9.2 14.951 11.6 14.953 ;
  LAYER M2 ;
        RECT 9.2 14.867 11.6 14.869 ;
  LAYER M2 ;
        RECT 9.2 14.783 11.6 14.785 ;
  LAYER M2 ;
        RECT 9.2 14.699 11.6 14.701 ;
  LAYER M2 ;
        RECT 9.2 14.615 11.6 14.617 ;
  LAYER M2 ;
        RECT 9.2 14.531 11.6 14.533 ;
  LAYER M2 ;
        RECT 9.2 14.447 11.6 14.449 ;
  LAYER M2 ;
        RECT 9.2 14.363 11.6 14.365 ;
  LAYER M2 ;
        RECT 9.2 14.279 11.6 14.281 ;
  LAYER M2 ;
        RECT 9.2 14.195 11.6 14.197 ;
  LAYER M2 ;
        RECT 9.2 14.111 11.6 14.113 ;
  LAYER M2 ;
        RECT 9.2 14.027 11.6 14.029 ;
  LAYER M2 ;
        RECT 9.2 13.943 11.6 13.945 ;
  LAYER M2 ;
        RECT 9.2 13.859 11.6 13.861 ;
  LAYER M1 ;
        RECT 11.584 10.8 11.616 13.308 ;
  LAYER M1 ;
        RECT 11.52 10.8 11.552 13.308 ;
  LAYER M1 ;
        RECT 11.456 10.8 11.488 13.308 ;
  LAYER M1 ;
        RECT 11.392 10.8 11.424 13.308 ;
  LAYER M1 ;
        RECT 11.328 10.8 11.36 13.308 ;
  LAYER M1 ;
        RECT 11.264 10.8 11.296 13.308 ;
  LAYER M1 ;
        RECT 11.2 10.8 11.232 13.308 ;
  LAYER M1 ;
        RECT 11.136 10.8 11.168 13.308 ;
  LAYER M1 ;
        RECT 11.072 10.8 11.104 13.308 ;
  LAYER M1 ;
        RECT 11.008 10.8 11.04 13.308 ;
  LAYER M1 ;
        RECT 10.944 10.8 10.976 13.308 ;
  LAYER M1 ;
        RECT 10.88 10.8 10.912 13.308 ;
  LAYER M1 ;
        RECT 10.816 10.8 10.848 13.308 ;
  LAYER M1 ;
        RECT 10.752 10.8 10.784 13.308 ;
  LAYER M1 ;
        RECT 10.688 10.8 10.72 13.308 ;
  LAYER M1 ;
        RECT 10.624 10.8 10.656 13.308 ;
  LAYER M1 ;
        RECT 10.56 10.8 10.592 13.308 ;
  LAYER M1 ;
        RECT 10.496 10.8 10.528 13.308 ;
  LAYER M1 ;
        RECT 10.432 10.8 10.464 13.308 ;
  LAYER M1 ;
        RECT 10.368 10.8 10.4 13.308 ;
  LAYER M1 ;
        RECT 10.304 10.8 10.336 13.308 ;
  LAYER M1 ;
        RECT 10.24 10.8 10.272 13.308 ;
  LAYER M1 ;
        RECT 10.176 10.8 10.208 13.308 ;
  LAYER M1 ;
        RECT 10.112 10.8 10.144 13.308 ;
  LAYER M1 ;
        RECT 10.048 10.8 10.08 13.308 ;
  LAYER M1 ;
        RECT 9.984 10.8 10.016 13.308 ;
  LAYER M1 ;
        RECT 9.92 10.8 9.952 13.308 ;
  LAYER M1 ;
        RECT 9.856 10.8 9.888 13.308 ;
  LAYER M1 ;
        RECT 9.792 10.8 9.824 13.308 ;
  LAYER M1 ;
        RECT 9.728 10.8 9.76 13.308 ;
  LAYER M1 ;
        RECT 9.664 10.8 9.696 13.308 ;
  LAYER M1 ;
        RECT 9.6 10.8 9.632 13.308 ;
  LAYER M1 ;
        RECT 9.536 10.8 9.568 13.308 ;
  LAYER M1 ;
        RECT 9.472 10.8 9.504 13.308 ;
  LAYER M1 ;
        RECT 9.408 10.8 9.44 13.308 ;
  LAYER M1 ;
        RECT 9.344 10.8 9.376 13.308 ;
  LAYER M1 ;
        RECT 9.28 10.8 9.312 13.308 ;
  LAYER M2 ;
        RECT 9.164 13.192 11.636 13.224 ;
  LAYER M2 ;
        RECT 9.164 13.128 11.636 13.16 ;
  LAYER M2 ;
        RECT 9.164 13.064 11.636 13.096 ;
  LAYER M2 ;
        RECT 9.164 13 11.636 13.032 ;
  LAYER M2 ;
        RECT 9.164 12.936 11.636 12.968 ;
  LAYER M2 ;
        RECT 9.164 12.872 11.636 12.904 ;
  LAYER M2 ;
        RECT 9.164 12.808 11.636 12.84 ;
  LAYER M2 ;
        RECT 9.164 12.744 11.636 12.776 ;
  LAYER M2 ;
        RECT 9.164 12.68 11.636 12.712 ;
  LAYER M2 ;
        RECT 9.164 12.616 11.636 12.648 ;
  LAYER M2 ;
        RECT 9.164 12.552 11.636 12.584 ;
  LAYER M2 ;
        RECT 9.164 12.488 11.636 12.52 ;
  LAYER M2 ;
        RECT 9.164 12.424 11.636 12.456 ;
  LAYER M2 ;
        RECT 9.164 12.36 11.636 12.392 ;
  LAYER M2 ;
        RECT 9.164 12.296 11.636 12.328 ;
  LAYER M2 ;
        RECT 9.164 12.232 11.636 12.264 ;
  LAYER M2 ;
        RECT 9.164 12.168 11.636 12.2 ;
  LAYER M2 ;
        RECT 9.164 12.104 11.636 12.136 ;
  LAYER M2 ;
        RECT 9.164 12.04 11.636 12.072 ;
  LAYER M2 ;
        RECT 9.164 11.976 11.636 12.008 ;
  LAYER M2 ;
        RECT 9.164 11.912 11.636 11.944 ;
  LAYER M2 ;
        RECT 9.164 11.848 11.636 11.88 ;
  LAYER M2 ;
        RECT 9.164 11.784 11.636 11.816 ;
  LAYER M2 ;
        RECT 9.164 11.72 11.636 11.752 ;
  LAYER M2 ;
        RECT 9.164 11.656 11.636 11.688 ;
  LAYER M2 ;
        RECT 9.164 11.592 11.636 11.624 ;
  LAYER M2 ;
        RECT 9.164 11.528 11.636 11.56 ;
  LAYER M2 ;
        RECT 9.164 11.464 11.636 11.496 ;
  LAYER M2 ;
        RECT 9.164 11.4 11.636 11.432 ;
  LAYER M2 ;
        RECT 9.164 11.336 11.636 11.368 ;
  LAYER M2 ;
        RECT 9.164 11.272 11.636 11.304 ;
  LAYER M2 ;
        RECT 9.164 11.208 11.636 11.24 ;
  LAYER M2 ;
        RECT 9.164 11.144 11.636 11.176 ;
  LAYER M2 ;
        RECT 9.164 11.08 11.636 11.112 ;
  LAYER M2 ;
        RECT 9.164 11.016 11.636 11.048 ;
  LAYER M2 ;
        RECT 9.164 10.952 11.636 10.984 ;
  LAYER M3 ;
        RECT 11.584 10.8 11.616 13.308 ;
  LAYER M3 ;
        RECT 11.52 10.8 11.552 13.308 ;
  LAYER M3 ;
        RECT 11.456 10.8 11.488 13.308 ;
  LAYER M3 ;
        RECT 11.392 10.8 11.424 13.308 ;
  LAYER M3 ;
        RECT 11.328 10.8 11.36 13.308 ;
  LAYER M3 ;
        RECT 11.264 10.8 11.296 13.308 ;
  LAYER M3 ;
        RECT 11.2 10.8 11.232 13.308 ;
  LAYER M3 ;
        RECT 11.136 10.8 11.168 13.308 ;
  LAYER M3 ;
        RECT 11.072 10.8 11.104 13.308 ;
  LAYER M3 ;
        RECT 11.008 10.8 11.04 13.308 ;
  LAYER M3 ;
        RECT 10.944 10.8 10.976 13.308 ;
  LAYER M3 ;
        RECT 10.88 10.8 10.912 13.308 ;
  LAYER M3 ;
        RECT 10.816 10.8 10.848 13.308 ;
  LAYER M3 ;
        RECT 10.752 10.8 10.784 13.308 ;
  LAYER M3 ;
        RECT 10.688 10.8 10.72 13.308 ;
  LAYER M3 ;
        RECT 10.624 10.8 10.656 13.308 ;
  LAYER M3 ;
        RECT 10.56 10.8 10.592 13.308 ;
  LAYER M3 ;
        RECT 10.496 10.8 10.528 13.308 ;
  LAYER M3 ;
        RECT 10.432 10.8 10.464 13.308 ;
  LAYER M3 ;
        RECT 10.368 10.8 10.4 13.308 ;
  LAYER M3 ;
        RECT 10.304 10.8 10.336 13.308 ;
  LAYER M3 ;
        RECT 10.24 10.8 10.272 13.308 ;
  LAYER M3 ;
        RECT 10.176 10.8 10.208 13.308 ;
  LAYER M3 ;
        RECT 10.112 10.8 10.144 13.308 ;
  LAYER M3 ;
        RECT 10.048 10.8 10.08 13.308 ;
  LAYER M3 ;
        RECT 9.984 10.8 10.016 13.308 ;
  LAYER M3 ;
        RECT 9.92 10.8 9.952 13.308 ;
  LAYER M3 ;
        RECT 9.856 10.8 9.888 13.308 ;
  LAYER M3 ;
        RECT 9.792 10.8 9.824 13.308 ;
  LAYER M3 ;
        RECT 9.728 10.8 9.76 13.308 ;
  LAYER M3 ;
        RECT 9.664 10.8 9.696 13.308 ;
  LAYER M3 ;
        RECT 9.6 10.8 9.632 13.308 ;
  LAYER M3 ;
        RECT 9.536 10.8 9.568 13.308 ;
  LAYER M3 ;
        RECT 9.472 10.8 9.504 13.308 ;
  LAYER M3 ;
        RECT 9.408 10.8 9.44 13.308 ;
  LAYER M3 ;
        RECT 9.344 10.8 9.376 13.308 ;
  LAYER M3 ;
        RECT 9.28 10.8 9.312 13.308 ;
  LAYER M3 ;
        RECT 9.184 10.8 9.216 13.308 ;
  LAYER M1 ;
        RECT 11.599 10.836 11.601 13.272 ;
  LAYER M1 ;
        RECT 11.519 10.836 11.521 13.272 ;
  LAYER M1 ;
        RECT 11.439 10.836 11.441 13.272 ;
  LAYER M1 ;
        RECT 11.359 10.836 11.361 13.272 ;
  LAYER M1 ;
        RECT 11.279 10.836 11.281 13.272 ;
  LAYER M1 ;
        RECT 11.199 10.836 11.201 13.272 ;
  LAYER M1 ;
        RECT 11.119 10.836 11.121 13.272 ;
  LAYER M1 ;
        RECT 11.039 10.836 11.041 13.272 ;
  LAYER M1 ;
        RECT 10.959 10.836 10.961 13.272 ;
  LAYER M1 ;
        RECT 10.879 10.836 10.881 13.272 ;
  LAYER M1 ;
        RECT 10.799 10.836 10.801 13.272 ;
  LAYER M1 ;
        RECT 10.719 10.836 10.721 13.272 ;
  LAYER M1 ;
        RECT 10.639 10.836 10.641 13.272 ;
  LAYER M1 ;
        RECT 10.559 10.836 10.561 13.272 ;
  LAYER M1 ;
        RECT 10.479 10.836 10.481 13.272 ;
  LAYER M1 ;
        RECT 10.399 10.836 10.401 13.272 ;
  LAYER M1 ;
        RECT 10.319 10.836 10.321 13.272 ;
  LAYER M1 ;
        RECT 10.239 10.836 10.241 13.272 ;
  LAYER M1 ;
        RECT 10.159 10.836 10.161 13.272 ;
  LAYER M1 ;
        RECT 10.079 10.836 10.081 13.272 ;
  LAYER M1 ;
        RECT 9.999 10.836 10.001 13.272 ;
  LAYER M1 ;
        RECT 9.919 10.836 9.921 13.272 ;
  LAYER M1 ;
        RECT 9.839 10.836 9.841 13.272 ;
  LAYER M1 ;
        RECT 9.759 10.836 9.761 13.272 ;
  LAYER M1 ;
        RECT 9.679 10.836 9.681 13.272 ;
  LAYER M1 ;
        RECT 9.599 10.836 9.601 13.272 ;
  LAYER M1 ;
        RECT 9.519 10.836 9.521 13.272 ;
  LAYER M1 ;
        RECT 9.439 10.836 9.441 13.272 ;
  LAYER M1 ;
        RECT 9.359 10.836 9.361 13.272 ;
  LAYER M1 ;
        RECT 9.279 10.836 9.281 13.272 ;
  LAYER M2 ;
        RECT 9.2 13.271 11.6 13.273 ;
  LAYER M2 ;
        RECT 9.2 13.187 11.6 13.189 ;
  LAYER M2 ;
        RECT 9.2 13.103 11.6 13.105 ;
  LAYER M2 ;
        RECT 9.2 13.019 11.6 13.021 ;
  LAYER M2 ;
        RECT 9.2 12.935 11.6 12.937 ;
  LAYER M2 ;
        RECT 9.2 12.851 11.6 12.853 ;
  LAYER M2 ;
        RECT 9.2 12.767 11.6 12.769 ;
  LAYER M2 ;
        RECT 9.2 12.683 11.6 12.685 ;
  LAYER M2 ;
        RECT 9.2 12.599 11.6 12.601 ;
  LAYER M2 ;
        RECT 9.2 12.515 11.6 12.517 ;
  LAYER M2 ;
        RECT 9.2 12.431 11.6 12.433 ;
  LAYER M2 ;
        RECT 9.2 12.347 11.6 12.349 ;
  LAYER M2 ;
        RECT 9.2 12.2635 11.6 12.2655 ;
  LAYER M2 ;
        RECT 9.2 12.179 11.6 12.181 ;
  LAYER M2 ;
        RECT 9.2 12.095 11.6 12.097 ;
  LAYER M2 ;
        RECT 9.2 12.011 11.6 12.013 ;
  LAYER M2 ;
        RECT 9.2 11.927 11.6 11.929 ;
  LAYER M2 ;
        RECT 9.2 11.843 11.6 11.845 ;
  LAYER M2 ;
        RECT 9.2 11.759 11.6 11.761 ;
  LAYER M2 ;
        RECT 9.2 11.675 11.6 11.677 ;
  LAYER M2 ;
        RECT 9.2 11.591 11.6 11.593 ;
  LAYER M2 ;
        RECT 9.2 11.507 11.6 11.509 ;
  LAYER M2 ;
        RECT 9.2 11.423 11.6 11.425 ;
  LAYER M2 ;
        RECT 9.2 11.339 11.6 11.341 ;
  LAYER M2 ;
        RECT 9.2 11.255 11.6 11.257 ;
  LAYER M2 ;
        RECT 9.2 11.171 11.6 11.173 ;
  LAYER M2 ;
        RECT 9.2 11.087 11.6 11.089 ;
  LAYER M2 ;
        RECT 9.2 11.003 11.6 11.005 ;
  LAYER M2 ;
        RECT 9.2 10.919 11.6 10.921 ;
  LAYER M1 ;
        RECT 11.584 7.86 11.616 10.368 ;
  LAYER M1 ;
        RECT 11.52 7.86 11.552 10.368 ;
  LAYER M1 ;
        RECT 11.456 7.86 11.488 10.368 ;
  LAYER M1 ;
        RECT 11.392 7.86 11.424 10.368 ;
  LAYER M1 ;
        RECT 11.328 7.86 11.36 10.368 ;
  LAYER M1 ;
        RECT 11.264 7.86 11.296 10.368 ;
  LAYER M1 ;
        RECT 11.2 7.86 11.232 10.368 ;
  LAYER M1 ;
        RECT 11.136 7.86 11.168 10.368 ;
  LAYER M1 ;
        RECT 11.072 7.86 11.104 10.368 ;
  LAYER M1 ;
        RECT 11.008 7.86 11.04 10.368 ;
  LAYER M1 ;
        RECT 10.944 7.86 10.976 10.368 ;
  LAYER M1 ;
        RECT 10.88 7.86 10.912 10.368 ;
  LAYER M1 ;
        RECT 10.816 7.86 10.848 10.368 ;
  LAYER M1 ;
        RECT 10.752 7.86 10.784 10.368 ;
  LAYER M1 ;
        RECT 10.688 7.86 10.72 10.368 ;
  LAYER M1 ;
        RECT 10.624 7.86 10.656 10.368 ;
  LAYER M1 ;
        RECT 10.56 7.86 10.592 10.368 ;
  LAYER M1 ;
        RECT 10.496 7.86 10.528 10.368 ;
  LAYER M1 ;
        RECT 10.432 7.86 10.464 10.368 ;
  LAYER M1 ;
        RECT 10.368 7.86 10.4 10.368 ;
  LAYER M1 ;
        RECT 10.304 7.86 10.336 10.368 ;
  LAYER M1 ;
        RECT 10.24 7.86 10.272 10.368 ;
  LAYER M1 ;
        RECT 10.176 7.86 10.208 10.368 ;
  LAYER M1 ;
        RECT 10.112 7.86 10.144 10.368 ;
  LAYER M1 ;
        RECT 10.048 7.86 10.08 10.368 ;
  LAYER M1 ;
        RECT 9.984 7.86 10.016 10.368 ;
  LAYER M1 ;
        RECT 9.92 7.86 9.952 10.368 ;
  LAYER M1 ;
        RECT 9.856 7.86 9.888 10.368 ;
  LAYER M1 ;
        RECT 9.792 7.86 9.824 10.368 ;
  LAYER M1 ;
        RECT 9.728 7.86 9.76 10.368 ;
  LAYER M1 ;
        RECT 9.664 7.86 9.696 10.368 ;
  LAYER M1 ;
        RECT 9.6 7.86 9.632 10.368 ;
  LAYER M1 ;
        RECT 9.536 7.86 9.568 10.368 ;
  LAYER M1 ;
        RECT 9.472 7.86 9.504 10.368 ;
  LAYER M1 ;
        RECT 9.408 7.86 9.44 10.368 ;
  LAYER M1 ;
        RECT 9.344 7.86 9.376 10.368 ;
  LAYER M1 ;
        RECT 9.28 7.86 9.312 10.368 ;
  LAYER M2 ;
        RECT 9.164 10.252 11.636 10.284 ;
  LAYER M2 ;
        RECT 9.164 10.188 11.636 10.22 ;
  LAYER M2 ;
        RECT 9.164 10.124 11.636 10.156 ;
  LAYER M2 ;
        RECT 9.164 10.06 11.636 10.092 ;
  LAYER M2 ;
        RECT 9.164 9.996 11.636 10.028 ;
  LAYER M2 ;
        RECT 9.164 9.932 11.636 9.964 ;
  LAYER M2 ;
        RECT 9.164 9.868 11.636 9.9 ;
  LAYER M2 ;
        RECT 9.164 9.804 11.636 9.836 ;
  LAYER M2 ;
        RECT 9.164 9.74 11.636 9.772 ;
  LAYER M2 ;
        RECT 9.164 9.676 11.636 9.708 ;
  LAYER M2 ;
        RECT 9.164 9.612 11.636 9.644 ;
  LAYER M2 ;
        RECT 9.164 9.548 11.636 9.58 ;
  LAYER M2 ;
        RECT 9.164 9.484 11.636 9.516 ;
  LAYER M2 ;
        RECT 9.164 9.42 11.636 9.452 ;
  LAYER M2 ;
        RECT 9.164 9.356 11.636 9.388 ;
  LAYER M2 ;
        RECT 9.164 9.292 11.636 9.324 ;
  LAYER M2 ;
        RECT 9.164 9.228 11.636 9.26 ;
  LAYER M2 ;
        RECT 9.164 9.164 11.636 9.196 ;
  LAYER M2 ;
        RECT 9.164 9.1 11.636 9.132 ;
  LAYER M2 ;
        RECT 9.164 9.036 11.636 9.068 ;
  LAYER M2 ;
        RECT 9.164 8.972 11.636 9.004 ;
  LAYER M2 ;
        RECT 9.164 8.908 11.636 8.94 ;
  LAYER M2 ;
        RECT 9.164 8.844 11.636 8.876 ;
  LAYER M2 ;
        RECT 9.164 8.78 11.636 8.812 ;
  LAYER M2 ;
        RECT 9.164 8.716 11.636 8.748 ;
  LAYER M2 ;
        RECT 9.164 8.652 11.636 8.684 ;
  LAYER M2 ;
        RECT 9.164 8.588 11.636 8.62 ;
  LAYER M2 ;
        RECT 9.164 8.524 11.636 8.556 ;
  LAYER M2 ;
        RECT 9.164 8.46 11.636 8.492 ;
  LAYER M2 ;
        RECT 9.164 8.396 11.636 8.428 ;
  LAYER M2 ;
        RECT 9.164 8.332 11.636 8.364 ;
  LAYER M2 ;
        RECT 9.164 8.268 11.636 8.3 ;
  LAYER M2 ;
        RECT 9.164 8.204 11.636 8.236 ;
  LAYER M2 ;
        RECT 9.164 8.14 11.636 8.172 ;
  LAYER M2 ;
        RECT 9.164 8.076 11.636 8.108 ;
  LAYER M2 ;
        RECT 9.164 8.012 11.636 8.044 ;
  LAYER M3 ;
        RECT 11.584 7.86 11.616 10.368 ;
  LAYER M3 ;
        RECT 11.52 7.86 11.552 10.368 ;
  LAYER M3 ;
        RECT 11.456 7.86 11.488 10.368 ;
  LAYER M3 ;
        RECT 11.392 7.86 11.424 10.368 ;
  LAYER M3 ;
        RECT 11.328 7.86 11.36 10.368 ;
  LAYER M3 ;
        RECT 11.264 7.86 11.296 10.368 ;
  LAYER M3 ;
        RECT 11.2 7.86 11.232 10.368 ;
  LAYER M3 ;
        RECT 11.136 7.86 11.168 10.368 ;
  LAYER M3 ;
        RECT 11.072 7.86 11.104 10.368 ;
  LAYER M3 ;
        RECT 11.008 7.86 11.04 10.368 ;
  LAYER M3 ;
        RECT 10.944 7.86 10.976 10.368 ;
  LAYER M3 ;
        RECT 10.88 7.86 10.912 10.368 ;
  LAYER M3 ;
        RECT 10.816 7.86 10.848 10.368 ;
  LAYER M3 ;
        RECT 10.752 7.86 10.784 10.368 ;
  LAYER M3 ;
        RECT 10.688 7.86 10.72 10.368 ;
  LAYER M3 ;
        RECT 10.624 7.86 10.656 10.368 ;
  LAYER M3 ;
        RECT 10.56 7.86 10.592 10.368 ;
  LAYER M3 ;
        RECT 10.496 7.86 10.528 10.368 ;
  LAYER M3 ;
        RECT 10.432 7.86 10.464 10.368 ;
  LAYER M3 ;
        RECT 10.368 7.86 10.4 10.368 ;
  LAYER M3 ;
        RECT 10.304 7.86 10.336 10.368 ;
  LAYER M3 ;
        RECT 10.24 7.86 10.272 10.368 ;
  LAYER M3 ;
        RECT 10.176 7.86 10.208 10.368 ;
  LAYER M3 ;
        RECT 10.112 7.86 10.144 10.368 ;
  LAYER M3 ;
        RECT 10.048 7.86 10.08 10.368 ;
  LAYER M3 ;
        RECT 9.984 7.86 10.016 10.368 ;
  LAYER M3 ;
        RECT 9.92 7.86 9.952 10.368 ;
  LAYER M3 ;
        RECT 9.856 7.86 9.888 10.368 ;
  LAYER M3 ;
        RECT 9.792 7.86 9.824 10.368 ;
  LAYER M3 ;
        RECT 9.728 7.86 9.76 10.368 ;
  LAYER M3 ;
        RECT 9.664 7.86 9.696 10.368 ;
  LAYER M3 ;
        RECT 9.6 7.86 9.632 10.368 ;
  LAYER M3 ;
        RECT 9.536 7.86 9.568 10.368 ;
  LAYER M3 ;
        RECT 9.472 7.86 9.504 10.368 ;
  LAYER M3 ;
        RECT 9.408 7.86 9.44 10.368 ;
  LAYER M3 ;
        RECT 9.344 7.86 9.376 10.368 ;
  LAYER M3 ;
        RECT 9.28 7.86 9.312 10.368 ;
  LAYER M3 ;
        RECT 9.184 7.86 9.216 10.368 ;
  LAYER M1 ;
        RECT 11.599 7.896 11.601 10.332 ;
  LAYER M1 ;
        RECT 11.519 7.896 11.521 10.332 ;
  LAYER M1 ;
        RECT 11.439 7.896 11.441 10.332 ;
  LAYER M1 ;
        RECT 11.359 7.896 11.361 10.332 ;
  LAYER M1 ;
        RECT 11.279 7.896 11.281 10.332 ;
  LAYER M1 ;
        RECT 11.199 7.896 11.201 10.332 ;
  LAYER M1 ;
        RECT 11.119 7.896 11.121 10.332 ;
  LAYER M1 ;
        RECT 11.039 7.896 11.041 10.332 ;
  LAYER M1 ;
        RECT 10.959 7.896 10.961 10.332 ;
  LAYER M1 ;
        RECT 10.879 7.896 10.881 10.332 ;
  LAYER M1 ;
        RECT 10.799 7.896 10.801 10.332 ;
  LAYER M1 ;
        RECT 10.719 7.896 10.721 10.332 ;
  LAYER M1 ;
        RECT 10.639 7.896 10.641 10.332 ;
  LAYER M1 ;
        RECT 10.559 7.896 10.561 10.332 ;
  LAYER M1 ;
        RECT 10.479 7.896 10.481 10.332 ;
  LAYER M1 ;
        RECT 10.399 7.896 10.401 10.332 ;
  LAYER M1 ;
        RECT 10.319 7.896 10.321 10.332 ;
  LAYER M1 ;
        RECT 10.239 7.896 10.241 10.332 ;
  LAYER M1 ;
        RECT 10.159 7.896 10.161 10.332 ;
  LAYER M1 ;
        RECT 10.079 7.896 10.081 10.332 ;
  LAYER M1 ;
        RECT 9.999 7.896 10.001 10.332 ;
  LAYER M1 ;
        RECT 9.919 7.896 9.921 10.332 ;
  LAYER M1 ;
        RECT 9.839 7.896 9.841 10.332 ;
  LAYER M1 ;
        RECT 9.759 7.896 9.761 10.332 ;
  LAYER M1 ;
        RECT 9.679 7.896 9.681 10.332 ;
  LAYER M1 ;
        RECT 9.599 7.896 9.601 10.332 ;
  LAYER M1 ;
        RECT 9.519 7.896 9.521 10.332 ;
  LAYER M1 ;
        RECT 9.439 7.896 9.441 10.332 ;
  LAYER M1 ;
        RECT 9.359 7.896 9.361 10.332 ;
  LAYER M1 ;
        RECT 9.279 7.896 9.281 10.332 ;
  LAYER M2 ;
        RECT 9.2 10.331 11.6 10.333 ;
  LAYER M2 ;
        RECT 9.2 10.247 11.6 10.249 ;
  LAYER M2 ;
        RECT 9.2 10.163 11.6 10.165 ;
  LAYER M2 ;
        RECT 9.2 10.079 11.6 10.081 ;
  LAYER M2 ;
        RECT 9.2 9.995 11.6 9.997 ;
  LAYER M2 ;
        RECT 9.2 9.911 11.6 9.913 ;
  LAYER M2 ;
        RECT 9.2 9.827 11.6 9.829 ;
  LAYER M2 ;
        RECT 9.2 9.743 11.6 9.745 ;
  LAYER M2 ;
        RECT 9.2 9.659 11.6 9.661 ;
  LAYER M2 ;
        RECT 9.2 9.575 11.6 9.577 ;
  LAYER M2 ;
        RECT 9.2 9.491 11.6 9.493 ;
  LAYER M2 ;
        RECT 9.2 9.407 11.6 9.409 ;
  LAYER M2 ;
        RECT 9.2 9.3235 11.6 9.3255 ;
  LAYER M2 ;
        RECT 9.2 9.239 11.6 9.241 ;
  LAYER M2 ;
        RECT 9.2 9.155 11.6 9.157 ;
  LAYER M2 ;
        RECT 9.2 9.071 11.6 9.073 ;
  LAYER M2 ;
        RECT 9.2 8.987 11.6 8.989 ;
  LAYER M2 ;
        RECT 9.2 8.903 11.6 8.905 ;
  LAYER M2 ;
        RECT 9.2 8.819 11.6 8.821 ;
  LAYER M2 ;
        RECT 9.2 8.735 11.6 8.737 ;
  LAYER M2 ;
        RECT 9.2 8.651 11.6 8.653 ;
  LAYER M2 ;
        RECT 9.2 8.567 11.6 8.569 ;
  LAYER M2 ;
        RECT 9.2 8.483 11.6 8.485 ;
  LAYER M2 ;
        RECT 9.2 8.399 11.6 8.401 ;
  LAYER M2 ;
        RECT 9.2 8.315 11.6 8.317 ;
  LAYER M2 ;
        RECT 9.2 8.231 11.6 8.233 ;
  LAYER M2 ;
        RECT 9.2 8.147 11.6 8.149 ;
  LAYER M2 ;
        RECT 9.2 8.063 11.6 8.065 ;
  LAYER M2 ;
        RECT 9.2 7.979 11.6 7.981 ;
  LAYER M1 ;
        RECT 11.584 4.92 11.616 7.428 ;
  LAYER M1 ;
        RECT 11.52 4.92 11.552 7.428 ;
  LAYER M1 ;
        RECT 11.456 4.92 11.488 7.428 ;
  LAYER M1 ;
        RECT 11.392 4.92 11.424 7.428 ;
  LAYER M1 ;
        RECT 11.328 4.92 11.36 7.428 ;
  LAYER M1 ;
        RECT 11.264 4.92 11.296 7.428 ;
  LAYER M1 ;
        RECT 11.2 4.92 11.232 7.428 ;
  LAYER M1 ;
        RECT 11.136 4.92 11.168 7.428 ;
  LAYER M1 ;
        RECT 11.072 4.92 11.104 7.428 ;
  LAYER M1 ;
        RECT 11.008 4.92 11.04 7.428 ;
  LAYER M1 ;
        RECT 10.944 4.92 10.976 7.428 ;
  LAYER M1 ;
        RECT 10.88 4.92 10.912 7.428 ;
  LAYER M1 ;
        RECT 10.816 4.92 10.848 7.428 ;
  LAYER M1 ;
        RECT 10.752 4.92 10.784 7.428 ;
  LAYER M1 ;
        RECT 10.688 4.92 10.72 7.428 ;
  LAYER M1 ;
        RECT 10.624 4.92 10.656 7.428 ;
  LAYER M1 ;
        RECT 10.56 4.92 10.592 7.428 ;
  LAYER M1 ;
        RECT 10.496 4.92 10.528 7.428 ;
  LAYER M1 ;
        RECT 10.432 4.92 10.464 7.428 ;
  LAYER M1 ;
        RECT 10.368 4.92 10.4 7.428 ;
  LAYER M1 ;
        RECT 10.304 4.92 10.336 7.428 ;
  LAYER M1 ;
        RECT 10.24 4.92 10.272 7.428 ;
  LAYER M1 ;
        RECT 10.176 4.92 10.208 7.428 ;
  LAYER M1 ;
        RECT 10.112 4.92 10.144 7.428 ;
  LAYER M1 ;
        RECT 10.048 4.92 10.08 7.428 ;
  LAYER M1 ;
        RECT 9.984 4.92 10.016 7.428 ;
  LAYER M1 ;
        RECT 9.92 4.92 9.952 7.428 ;
  LAYER M1 ;
        RECT 9.856 4.92 9.888 7.428 ;
  LAYER M1 ;
        RECT 9.792 4.92 9.824 7.428 ;
  LAYER M1 ;
        RECT 9.728 4.92 9.76 7.428 ;
  LAYER M1 ;
        RECT 9.664 4.92 9.696 7.428 ;
  LAYER M1 ;
        RECT 9.6 4.92 9.632 7.428 ;
  LAYER M1 ;
        RECT 9.536 4.92 9.568 7.428 ;
  LAYER M1 ;
        RECT 9.472 4.92 9.504 7.428 ;
  LAYER M1 ;
        RECT 9.408 4.92 9.44 7.428 ;
  LAYER M1 ;
        RECT 9.344 4.92 9.376 7.428 ;
  LAYER M1 ;
        RECT 9.28 4.92 9.312 7.428 ;
  LAYER M2 ;
        RECT 9.164 7.312 11.636 7.344 ;
  LAYER M2 ;
        RECT 9.164 7.248 11.636 7.28 ;
  LAYER M2 ;
        RECT 9.164 7.184 11.636 7.216 ;
  LAYER M2 ;
        RECT 9.164 7.12 11.636 7.152 ;
  LAYER M2 ;
        RECT 9.164 7.056 11.636 7.088 ;
  LAYER M2 ;
        RECT 9.164 6.992 11.636 7.024 ;
  LAYER M2 ;
        RECT 9.164 6.928 11.636 6.96 ;
  LAYER M2 ;
        RECT 9.164 6.864 11.636 6.896 ;
  LAYER M2 ;
        RECT 9.164 6.8 11.636 6.832 ;
  LAYER M2 ;
        RECT 9.164 6.736 11.636 6.768 ;
  LAYER M2 ;
        RECT 9.164 6.672 11.636 6.704 ;
  LAYER M2 ;
        RECT 9.164 6.608 11.636 6.64 ;
  LAYER M2 ;
        RECT 9.164 6.544 11.636 6.576 ;
  LAYER M2 ;
        RECT 9.164 6.48 11.636 6.512 ;
  LAYER M2 ;
        RECT 9.164 6.416 11.636 6.448 ;
  LAYER M2 ;
        RECT 9.164 6.352 11.636 6.384 ;
  LAYER M2 ;
        RECT 9.164 6.288 11.636 6.32 ;
  LAYER M2 ;
        RECT 9.164 6.224 11.636 6.256 ;
  LAYER M2 ;
        RECT 9.164 6.16 11.636 6.192 ;
  LAYER M2 ;
        RECT 9.164 6.096 11.636 6.128 ;
  LAYER M2 ;
        RECT 9.164 6.032 11.636 6.064 ;
  LAYER M2 ;
        RECT 9.164 5.968 11.636 6 ;
  LAYER M2 ;
        RECT 9.164 5.904 11.636 5.936 ;
  LAYER M2 ;
        RECT 9.164 5.84 11.636 5.872 ;
  LAYER M2 ;
        RECT 9.164 5.776 11.636 5.808 ;
  LAYER M2 ;
        RECT 9.164 5.712 11.636 5.744 ;
  LAYER M2 ;
        RECT 9.164 5.648 11.636 5.68 ;
  LAYER M2 ;
        RECT 9.164 5.584 11.636 5.616 ;
  LAYER M2 ;
        RECT 9.164 5.52 11.636 5.552 ;
  LAYER M2 ;
        RECT 9.164 5.456 11.636 5.488 ;
  LAYER M2 ;
        RECT 9.164 5.392 11.636 5.424 ;
  LAYER M2 ;
        RECT 9.164 5.328 11.636 5.36 ;
  LAYER M2 ;
        RECT 9.164 5.264 11.636 5.296 ;
  LAYER M2 ;
        RECT 9.164 5.2 11.636 5.232 ;
  LAYER M2 ;
        RECT 9.164 5.136 11.636 5.168 ;
  LAYER M2 ;
        RECT 9.164 5.072 11.636 5.104 ;
  LAYER M3 ;
        RECT 11.584 4.92 11.616 7.428 ;
  LAYER M3 ;
        RECT 11.52 4.92 11.552 7.428 ;
  LAYER M3 ;
        RECT 11.456 4.92 11.488 7.428 ;
  LAYER M3 ;
        RECT 11.392 4.92 11.424 7.428 ;
  LAYER M3 ;
        RECT 11.328 4.92 11.36 7.428 ;
  LAYER M3 ;
        RECT 11.264 4.92 11.296 7.428 ;
  LAYER M3 ;
        RECT 11.2 4.92 11.232 7.428 ;
  LAYER M3 ;
        RECT 11.136 4.92 11.168 7.428 ;
  LAYER M3 ;
        RECT 11.072 4.92 11.104 7.428 ;
  LAYER M3 ;
        RECT 11.008 4.92 11.04 7.428 ;
  LAYER M3 ;
        RECT 10.944 4.92 10.976 7.428 ;
  LAYER M3 ;
        RECT 10.88 4.92 10.912 7.428 ;
  LAYER M3 ;
        RECT 10.816 4.92 10.848 7.428 ;
  LAYER M3 ;
        RECT 10.752 4.92 10.784 7.428 ;
  LAYER M3 ;
        RECT 10.688 4.92 10.72 7.428 ;
  LAYER M3 ;
        RECT 10.624 4.92 10.656 7.428 ;
  LAYER M3 ;
        RECT 10.56 4.92 10.592 7.428 ;
  LAYER M3 ;
        RECT 10.496 4.92 10.528 7.428 ;
  LAYER M3 ;
        RECT 10.432 4.92 10.464 7.428 ;
  LAYER M3 ;
        RECT 10.368 4.92 10.4 7.428 ;
  LAYER M3 ;
        RECT 10.304 4.92 10.336 7.428 ;
  LAYER M3 ;
        RECT 10.24 4.92 10.272 7.428 ;
  LAYER M3 ;
        RECT 10.176 4.92 10.208 7.428 ;
  LAYER M3 ;
        RECT 10.112 4.92 10.144 7.428 ;
  LAYER M3 ;
        RECT 10.048 4.92 10.08 7.428 ;
  LAYER M3 ;
        RECT 9.984 4.92 10.016 7.428 ;
  LAYER M3 ;
        RECT 9.92 4.92 9.952 7.428 ;
  LAYER M3 ;
        RECT 9.856 4.92 9.888 7.428 ;
  LAYER M3 ;
        RECT 9.792 4.92 9.824 7.428 ;
  LAYER M3 ;
        RECT 9.728 4.92 9.76 7.428 ;
  LAYER M3 ;
        RECT 9.664 4.92 9.696 7.428 ;
  LAYER M3 ;
        RECT 9.6 4.92 9.632 7.428 ;
  LAYER M3 ;
        RECT 9.536 4.92 9.568 7.428 ;
  LAYER M3 ;
        RECT 9.472 4.92 9.504 7.428 ;
  LAYER M3 ;
        RECT 9.408 4.92 9.44 7.428 ;
  LAYER M3 ;
        RECT 9.344 4.92 9.376 7.428 ;
  LAYER M3 ;
        RECT 9.28 4.92 9.312 7.428 ;
  LAYER M3 ;
        RECT 9.184 4.92 9.216 7.428 ;
  LAYER M1 ;
        RECT 11.599 4.956 11.601 7.392 ;
  LAYER M1 ;
        RECT 11.519 4.956 11.521 7.392 ;
  LAYER M1 ;
        RECT 11.439 4.956 11.441 7.392 ;
  LAYER M1 ;
        RECT 11.359 4.956 11.361 7.392 ;
  LAYER M1 ;
        RECT 11.279 4.956 11.281 7.392 ;
  LAYER M1 ;
        RECT 11.199 4.956 11.201 7.392 ;
  LAYER M1 ;
        RECT 11.119 4.956 11.121 7.392 ;
  LAYER M1 ;
        RECT 11.039 4.956 11.041 7.392 ;
  LAYER M1 ;
        RECT 10.959 4.956 10.961 7.392 ;
  LAYER M1 ;
        RECT 10.879 4.956 10.881 7.392 ;
  LAYER M1 ;
        RECT 10.799 4.956 10.801 7.392 ;
  LAYER M1 ;
        RECT 10.719 4.956 10.721 7.392 ;
  LAYER M1 ;
        RECT 10.639 4.956 10.641 7.392 ;
  LAYER M1 ;
        RECT 10.559 4.956 10.561 7.392 ;
  LAYER M1 ;
        RECT 10.479 4.956 10.481 7.392 ;
  LAYER M1 ;
        RECT 10.399 4.956 10.401 7.392 ;
  LAYER M1 ;
        RECT 10.319 4.956 10.321 7.392 ;
  LAYER M1 ;
        RECT 10.239 4.956 10.241 7.392 ;
  LAYER M1 ;
        RECT 10.159 4.956 10.161 7.392 ;
  LAYER M1 ;
        RECT 10.079 4.956 10.081 7.392 ;
  LAYER M1 ;
        RECT 9.999 4.956 10.001 7.392 ;
  LAYER M1 ;
        RECT 9.919 4.956 9.921 7.392 ;
  LAYER M1 ;
        RECT 9.839 4.956 9.841 7.392 ;
  LAYER M1 ;
        RECT 9.759 4.956 9.761 7.392 ;
  LAYER M1 ;
        RECT 9.679 4.956 9.681 7.392 ;
  LAYER M1 ;
        RECT 9.599 4.956 9.601 7.392 ;
  LAYER M1 ;
        RECT 9.519 4.956 9.521 7.392 ;
  LAYER M1 ;
        RECT 9.439 4.956 9.441 7.392 ;
  LAYER M1 ;
        RECT 9.359 4.956 9.361 7.392 ;
  LAYER M1 ;
        RECT 9.279 4.956 9.281 7.392 ;
  LAYER M2 ;
        RECT 9.2 7.391 11.6 7.393 ;
  LAYER M2 ;
        RECT 9.2 7.307 11.6 7.309 ;
  LAYER M2 ;
        RECT 9.2 7.223 11.6 7.225 ;
  LAYER M2 ;
        RECT 9.2 7.139 11.6 7.141 ;
  LAYER M2 ;
        RECT 9.2 7.055 11.6 7.057 ;
  LAYER M2 ;
        RECT 9.2 6.971 11.6 6.973 ;
  LAYER M2 ;
        RECT 9.2 6.887 11.6 6.889 ;
  LAYER M2 ;
        RECT 9.2 6.803 11.6 6.805 ;
  LAYER M2 ;
        RECT 9.2 6.719 11.6 6.721 ;
  LAYER M2 ;
        RECT 9.2 6.635 11.6 6.637 ;
  LAYER M2 ;
        RECT 9.2 6.551 11.6 6.553 ;
  LAYER M2 ;
        RECT 9.2 6.467 11.6 6.469 ;
  LAYER M2 ;
        RECT 9.2 6.3835 11.6 6.3855 ;
  LAYER M2 ;
        RECT 9.2 6.299 11.6 6.301 ;
  LAYER M2 ;
        RECT 9.2 6.215 11.6 6.217 ;
  LAYER M2 ;
        RECT 9.2 6.131 11.6 6.133 ;
  LAYER M2 ;
        RECT 9.2 6.047 11.6 6.049 ;
  LAYER M2 ;
        RECT 9.2 5.963 11.6 5.965 ;
  LAYER M2 ;
        RECT 9.2 5.879 11.6 5.881 ;
  LAYER M2 ;
        RECT 9.2 5.795 11.6 5.797 ;
  LAYER M2 ;
        RECT 9.2 5.711 11.6 5.713 ;
  LAYER M2 ;
        RECT 9.2 5.627 11.6 5.629 ;
  LAYER M2 ;
        RECT 9.2 5.543 11.6 5.545 ;
  LAYER M2 ;
        RECT 9.2 5.459 11.6 5.461 ;
  LAYER M2 ;
        RECT 9.2 5.375 11.6 5.377 ;
  LAYER M2 ;
        RECT 9.2 5.291 11.6 5.293 ;
  LAYER M2 ;
        RECT 9.2 5.207 11.6 5.209 ;
  LAYER M2 ;
        RECT 9.2 5.123 11.6 5.125 ;
  LAYER M2 ;
        RECT 9.2 5.039 11.6 5.041 ;
  LAYER M1 ;
        RECT 11.584 1.98 11.616 4.488 ;
  LAYER M1 ;
        RECT 11.52 1.98 11.552 4.488 ;
  LAYER M1 ;
        RECT 11.456 1.98 11.488 4.488 ;
  LAYER M1 ;
        RECT 11.392 1.98 11.424 4.488 ;
  LAYER M1 ;
        RECT 11.328 1.98 11.36 4.488 ;
  LAYER M1 ;
        RECT 11.264 1.98 11.296 4.488 ;
  LAYER M1 ;
        RECT 11.2 1.98 11.232 4.488 ;
  LAYER M1 ;
        RECT 11.136 1.98 11.168 4.488 ;
  LAYER M1 ;
        RECT 11.072 1.98 11.104 4.488 ;
  LAYER M1 ;
        RECT 11.008 1.98 11.04 4.488 ;
  LAYER M1 ;
        RECT 10.944 1.98 10.976 4.488 ;
  LAYER M1 ;
        RECT 10.88 1.98 10.912 4.488 ;
  LAYER M1 ;
        RECT 10.816 1.98 10.848 4.488 ;
  LAYER M1 ;
        RECT 10.752 1.98 10.784 4.488 ;
  LAYER M1 ;
        RECT 10.688 1.98 10.72 4.488 ;
  LAYER M1 ;
        RECT 10.624 1.98 10.656 4.488 ;
  LAYER M1 ;
        RECT 10.56 1.98 10.592 4.488 ;
  LAYER M1 ;
        RECT 10.496 1.98 10.528 4.488 ;
  LAYER M1 ;
        RECT 10.432 1.98 10.464 4.488 ;
  LAYER M1 ;
        RECT 10.368 1.98 10.4 4.488 ;
  LAYER M1 ;
        RECT 10.304 1.98 10.336 4.488 ;
  LAYER M1 ;
        RECT 10.24 1.98 10.272 4.488 ;
  LAYER M1 ;
        RECT 10.176 1.98 10.208 4.488 ;
  LAYER M1 ;
        RECT 10.112 1.98 10.144 4.488 ;
  LAYER M1 ;
        RECT 10.048 1.98 10.08 4.488 ;
  LAYER M1 ;
        RECT 9.984 1.98 10.016 4.488 ;
  LAYER M1 ;
        RECT 9.92 1.98 9.952 4.488 ;
  LAYER M1 ;
        RECT 9.856 1.98 9.888 4.488 ;
  LAYER M1 ;
        RECT 9.792 1.98 9.824 4.488 ;
  LAYER M1 ;
        RECT 9.728 1.98 9.76 4.488 ;
  LAYER M1 ;
        RECT 9.664 1.98 9.696 4.488 ;
  LAYER M1 ;
        RECT 9.6 1.98 9.632 4.488 ;
  LAYER M1 ;
        RECT 9.536 1.98 9.568 4.488 ;
  LAYER M1 ;
        RECT 9.472 1.98 9.504 4.488 ;
  LAYER M1 ;
        RECT 9.408 1.98 9.44 4.488 ;
  LAYER M1 ;
        RECT 9.344 1.98 9.376 4.488 ;
  LAYER M1 ;
        RECT 9.28 1.98 9.312 4.488 ;
  LAYER M2 ;
        RECT 9.164 4.372 11.636 4.404 ;
  LAYER M2 ;
        RECT 9.164 4.308 11.636 4.34 ;
  LAYER M2 ;
        RECT 9.164 4.244 11.636 4.276 ;
  LAYER M2 ;
        RECT 9.164 4.18 11.636 4.212 ;
  LAYER M2 ;
        RECT 9.164 4.116 11.636 4.148 ;
  LAYER M2 ;
        RECT 9.164 4.052 11.636 4.084 ;
  LAYER M2 ;
        RECT 9.164 3.988 11.636 4.02 ;
  LAYER M2 ;
        RECT 9.164 3.924 11.636 3.956 ;
  LAYER M2 ;
        RECT 9.164 3.86 11.636 3.892 ;
  LAYER M2 ;
        RECT 9.164 3.796 11.636 3.828 ;
  LAYER M2 ;
        RECT 9.164 3.732 11.636 3.764 ;
  LAYER M2 ;
        RECT 9.164 3.668 11.636 3.7 ;
  LAYER M2 ;
        RECT 9.164 3.604 11.636 3.636 ;
  LAYER M2 ;
        RECT 9.164 3.54 11.636 3.572 ;
  LAYER M2 ;
        RECT 9.164 3.476 11.636 3.508 ;
  LAYER M2 ;
        RECT 9.164 3.412 11.636 3.444 ;
  LAYER M2 ;
        RECT 9.164 3.348 11.636 3.38 ;
  LAYER M2 ;
        RECT 9.164 3.284 11.636 3.316 ;
  LAYER M2 ;
        RECT 9.164 3.22 11.636 3.252 ;
  LAYER M2 ;
        RECT 9.164 3.156 11.636 3.188 ;
  LAYER M2 ;
        RECT 9.164 3.092 11.636 3.124 ;
  LAYER M2 ;
        RECT 9.164 3.028 11.636 3.06 ;
  LAYER M2 ;
        RECT 9.164 2.964 11.636 2.996 ;
  LAYER M2 ;
        RECT 9.164 2.9 11.636 2.932 ;
  LAYER M2 ;
        RECT 9.164 2.836 11.636 2.868 ;
  LAYER M2 ;
        RECT 9.164 2.772 11.636 2.804 ;
  LAYER M2 ;
        RECT 9.164 2.708 11.636 2.74 ;
  LAYER M2 ;
        RECT 9.164 2.644 11.636 2.676 ;
  LAYER M2 ;
        RECT 9.164 2.58 11.636 2.612 ;
  LAYER M2 ;
        RECT 9.164 2.516 11.636 2.548 ;
  LAYER M2 ;
        RECT 9.164 2.452 11.636 2.484 ;
  LAYER M2 ;
        RECT 9.164 2.388 11.636 2.42 ;
  LAYER M2 ;
        RECT 9.164 2.324 11.636 2.356 ;
  LAYER M2 ;
        RECT 9.164 2.26 11.636 2.292 ;
  LAYER M2 ;
        RECT 9.164 2.196 11.636 2.228 ;
  LAYER M2 ;
        RECT 9.164 2.132 11.636 2.164 ;
  LAYER M3 ;
        RECT 11.584 1.98 11.616 4.488 ;
  LAYER M3 ;
        RECT 11.52 1.98 11.552 4.488 ;
  LAYER M3 ;
        RECT 11.456 1.98 11.488 4.488 ;
  LAYER M3 ;
        RECT 11.392 1.98 11.424 4.488 ;
  LAYER M3 ;
        RECT 11.328 1.98 11.36 4.488 ;
  LAYER M3 ;
        RECT 11.264 1.98 11.296 4.488 ;
  LAYER M3 ;
        RECT 11.2 1.98 11.232 4.488 ;
  LAYER M3 ;
        RECT 11.136 1.98 11.168 4.488 ;
  LAYER M3 ;
        RECT 11.072 1.98 11.104 4.488 ;
  LAYER M3 ;
        RECT 11.008 1.98 11.04 4.488 ;
  LAYER M3 ;
        RECT 10.944 1.98 10.976 4.488 ;
  LAYER M3 ;
        RECT 10.88 1.98 10.912 4.488 ;
  LAYER M3 ;
        RECT 10.816 1.98 10.848 4.488 ;
  LAYER M3 ;
        RECT 10.752 1.98 10.784 4.488 ;
  LAYER M3 ;
        RECT 10.688 1.98 10.72 4.488 ;
  LAYER M3 ;
        RECT 10.624 1.98 10.656 4.488 ;
  LAYER M3 ;
        RECT 10.56 1.98 10.592 4.488 ;
  LAYER M3 ;
        RECT 10.496 1.98 10.528 4.488 ;
  LAYER M3 ;
        RECT 10.432 1.98 10.464 4.488 ;
  LAYER M3 ;
        RECT 10.368 1.98 10.4 4.488 ;
  LAYER M3 ;
        RECT 10.304 1.98 10.336 4.488 ;
  LAYER M3 ;
        RECT 10.24 1.98 10.272 4.488 ;
  LAYER M3 ;
        RECT 10.176 1.98 10.208 4.488 ;
  LAYER M3 ;
        RECT 10.112 1.98 10.144 4.488 ;
  LAYER M3 ;
        RECT 10.048 1.98 10.08 4.488 ;
  LAYER M3 ;
        RECT 9.984 1.98 10.016 4.488 ;
  LAYER M3 ;
        RECT 9.92 1.98 9.952 4.488 ;
  LAYER M3 ;
        RECT 9.856 1.98 9.888 4.488 ;
  LAYER M3 ;
        RECT 9.792 1.98 9.824 4.488 ;
  LAYER M3 ;
        RECT 9.728 1.98 9.76 4.488 ;
  LAYER M3 ;
        RECT 9.664 1.98 9.696 4.488 ;
  LAYER M3 ;
        RECT 9.6 1.98 9.632 4.488 ;
  LAYER M3 ;
        RECT 9.536 1.98 9.568 4.488 ;
  LAYER M3 ;
        RECT 9.472 1.98 9.504 4.488 ;
  LAYER M3 ;
        RECT 9.408 1.98 9.44 4.488 ;
  LAYER M3 ;
        RECT 9.344 1.98 9.376 4.488 ;
  LAYER M3 ;
        RECT 9.28 1.98 9.312 4.488 ;
  LAYER M3 ;
        RECT 9.184 1.98 9.216 4.488 ;
  LAYER M1 ;
        RECT 11.599 2.016 11.601 4.452 ;
  LAYER M1 ;
        RECT 11.519 2.016 11.521 4.452 ;
  LAYER M1 ;
        RECT 11.439 2.016 11.441 4.452 ;
  LAYER M1 ;
        RECT 11.359 2.016 11.361 4.452 ;
  LAYER M1 ;
        RECT 11.279 2.016 11.281 4.452 ;
  LAYER M1 ;
        RECT 11.199 2.016 11.201 4.452 ;
  LAYER M1 ;
        RECT 11.119 2.016 11.121 4.452 ;
  LAYER M1 ;
        RECT 11.039 2.016 11.041 4.452 ;
  LAYER M1 ;
        RECT 10.959 2.016 10.961 4.452 ;
  LAYER M1 ;
        RECT 10.879 2.016 10.881 4.452 ;
  LAYER M1 ;
        RECT 10.799 2.016 10.801 4.452 ;
  LAYER M1 ;
        RECT 10.719 2.016 10.721 4.452 ;
  LAYER M1 ;
        RECT 10.639 2.016 10.641 4.452 ;
  LAYER M1 ;
        RECT 10.559 2.016 10.561 4.452 ;
  LAYER M1 ;
        RECT 10.479 2.016 10.481 4.452 ;
  LAYER M1 ;
        RECT 10.399 2.016 10.401 4.452 ;
  LAYER M1 ;
        RECT 10.319 2.016 10.321 4.452 ;
  LAYER M1 ;
        RECT 10.239 2.016 10.241 4.452 ;
  LAYER M1 ;
        RECT 10.159 2.016 10.161 4.452 ;
  LAYER M1 ;
        RECT 10.079 2.016 10.081 4.452 ;
  LAYER M1 ;
        RECT 9.999 2.016 10.001 4.452 ;
  LAYER M1 ;
        RECT 9.919 2.016 9.921 4.452 ;
  LAYER M1 ;
        RECT 9.839 2.016 9.841 4.452 ;
  LAYER M1 ;
        RECT 9.759 2.016 9.761 4.452 ;
  LAYER M1 ;
        RECT 9.679 2.016 9.681 4.452 ;
  LAYER M1 ;
        RECT 9.599 2.016 9.601 4.452 ;
  LAYER M1 ;
        RECT 9.519 2.016 9.521 4.452 ;
  LAYER M1 ;
        RECT 9.439 2.016 9.441 4.452 ;
  LAYER M1 ;
        RECT 9.359 2.016 9.361 4.452 ;
  LAYER M1 ;
        RECT 9.279 2.016 9.281 4.452 ;
  LAYER M2 ;
        RECT 9.2 4.451 11.6 4.453 ;
  LAYER M2 ;
        RECT 9.2 4.367 11.6 4.369 ;
  LAYER M2 ;
        RECT 9.2 4.283 11.6 4.285 ;
  LAYER M2 ;
        RECT 9.2 4.199 11.6 4.201 ;
  LAYER M2 ;
        RECT 9.2 4.115 11.6 4.117 ;
  LAYER M2 ;
        RECT 9.2 4.031 11.6 4.033 ;
  LAYER M2 ;
        RECT 9.2 3.947 11.6 3.949 ;
  LAYER M2 ;
        RECT 9.2 3.863 11.6 3.865 ;
  LAYER M2 ;
        RECT 9.2 3.779 11.6 3.781 ;
  LAYER M2 ;
        RECT 9.2 3.695 11.6 3.697 ;
  LAYER M2 ;
        RECT 9.2 3.611 11.6 3.613 ;
  LAYER M2 ;
        RECT 9.2 3.527 11.6 3.529 ;
  LAYER M2 ;
        RECT 9.2 3.4435 11.6 3.4455 ;
  LAYER M2 ;
        RECT 9.2 3.359 11.6 3.361 ;
  LAYER M2 ;
        RECT 9.2 3.275 11.6 3.277 ;
  LAYER M2 ;
        RECT 9.2 3.191 11.6 3.193 ;
  LAYER M2 ;
        RECT 9.2 3.107 11.6 3.109 ;
  LAYER M2 ;
        RECT 9.2 3.023 11.6 3.025 ;
  LAYER M2 ;
        RECT 9.2 2.939 11.6 2.941 ;
  LAYER M2 ;
        RECT 9.2 2.855 11.6 2.857 ;
  LAYER M2 ;
        RECT 9.2 2.771 11.6 2.773 ;
  LAYER M2 ;
        RECT 9.2 2.687 11.6 2.689 ;
  LAYER M2 ;
        RECT 9.2 2.603 11.6 2.605 ;
  LAYER M2 ;
        RECT 9.2 2.519 11.6 2.521 ;
  LAYER M2 ;
        RECT 9.2 2.435 11.6 2.437 ;
  LAYER M2 ;
        RECT 9.2 2.351 11.6 2.353 ;
  LAYER M2 ;
        RECT 9.2 2.267 11.6 2.269 ;
  LAYER M2 ;
        RECT 9.2 2.183 11.6 2.185 ;
  LAYER M2 ;
        RECT 9.2 2.099 11.6 2.101 ;
  LAYER M1 ;
        RECT 8.704 13.74 8.736 16.248 ;
  LAYER M1 ;
        RECT 8.64 13.74 8.672 16.248 ;
  LAYER M1 ;
        RECT 8.576 13.74 8.608 16.248 ;
  LAYER M1 ;
        RECT 8.512 13.74 8.544 16.248 ;
  LAYER M1 ;
        RECT 8.448 13.74 8.48 16.248 ;
  LAYER M1 ;
        RECT 8.384 13.74 8.416 16.248 ;
  LAYER M1 ;
        RECT 8.32 13.74 8.352 16.248 ;
  LAYER M1 ;
        RECT 8.256 13.74 8.288 16.248 ;
  LAYER M1 ;
        RECT 8.192 13.74 8.224 16.248 ;
  LAYER M1 ;
        RECT 8.128 13.74 8.16 16.248 ;
  LAYER M1 ;
        RECT 8.064 13.74 8.096 16.248 ;
  LAYER M1 ;
        RECT 8 13.74 8.032 16.248 ;
  LAYER M1 ;
        RECT 7.936 13.74 7.968 16.248 ;
  LAYER M1 ;
        RECT 7.872 13.74 7.904 16.248 ;
  LAYER M1 ;
        RECT 7.808 13.74 7.84 16.248 ;
  LAYER M1 ;
        RECT 7.744 13.74 7.776 16.248 ;
  LAYER M1 ;
        RECT 7.68 13.74 7.712 16.248 ;
  LAYER M1 ;
        RECT 7.616 13.74 7.648 16.248 ;
  LAYER M1 ;
        RECT 7.552 13.74 7.584 16.248 ;
  LAYER M1 ;
        RECT 7.488 13.74 7.52 16.248 ;
  LAYER M1 ;
        RECT 7.424 13.74 7.456 16.248 ;
  LAYER M1 ;
        RECT 7.36 13.74 7.392 16.248 ;
  LAYER M1 ;
        RECT 7.296 13.74 7.328 16.248 ;
  LAYER M1 ;
        RECT 7.232 13.74 7.264 16.248 ;
  LAYER M1 ;
        RECT 7.168 13.74 7.2 16.248 ;
  LAYER M1 ;
        RECT 7.104 13.74 7.136 16.248 ;
  LAYER M1 ;
        RECT 7.04 13.74 7.072 16.248 ;
  LAYER M1 ;
        RECT 6.976 13.74 7.008 16.248 ;
  LAYER M1 ;
        RECT 6.912 13.74 6.944 16.248 ;
  LAYER M1 ;
        RECT 6.848 13.74 6.88 16.248 ;
  LAYER M1 ;
        RECT 6.784 13.74 6.816 16.248 ;
  LAYER M1 ;
        RECT 6.72 13.74 6.752 16.248 ;
  LAYER M1 ;
        RECT 6.656 13.74 6.688 16.248 ;
  LAYER M1 ;
        RECT 6.592 13.74 6.624 16.248 ;
  LAYER M1 ;
        RECT 6.528 13.74 6.56 16.248 ;
  LAYER M1 ;
        RECT 6.464 13.74 6.496 16.248 ;
  LAYER M1 ;
        RECT 6.4 13.74 6.432 16.248 ;
  LAYER M2 ;
        RECT 6.284 16.132 8.756 16.164 ;
  LAYER M2 ;
        RECT 6.284 16.068 8.756 16.1 ;
  LAYER M2 ;
        RECT 6.284 16.004 8.756 16.036 ;
  LAYER M2 ;
        RECT 6.284 15.94 8.756 15.972 ;
  LAYER M2 ;
        RECT 6.284 15.876 8.756 15.908 ;
  LAYER M2 ;
        RECT 6.284 15.812 8.756 15.844 ;
  LAYER M2 ;
        RECT 6.284 15.748 8.756 15.78 ;
  LAYER M2 ;
        RECT 6.284 15.684 8.756 15.716 ;
  LAYER M2 ;
        RECT 6.284 15.62 8.756 15.652 ;
  LAYER M2 ;
        RECT 6.284 15.556 8.756 15.588 ;
  LAYER M2 ;
        RECT 6.284 15.492 8.756 15.524 ;
  LAYER M2 ;
        RECT 6.284 15.428 8.756 15.46 ;
  LAYER M2 ;
        RECT 6.284 15.364 8.756 15.396 ;
  LAYER M2 ;
        RECT 6.284 15.3 8.756 15.332 ;
  LAYER M2 ;
        RECT 6.284 15.236 8.756 15.268 ;
  LAYER M2 ;
        RECT 6.284 15.172 8.756 15.204 ;
  LAYER M2 ;
        RECT 6.284 15.108 8.756 15.14 ;
  LAYER M2 ;
        RECT 6.284 15.044 8.756 15.076 ;
  LAYER M2 ;
        RECT 6.284 14.98 8.756 15.012 ;
  LAYER M2 ;
        RECT 6.284 14.916 8.756 14.948 ;
  LAYER M2 ;
        RECT 6.284 14.852 8.756 14.884 ;
  LAYER M2 ;
        RECT 6.284 14.788 8.756 14.82 ;
  LAYER M2 ;
        RECT 6.284 14.724 8.756 14.756 ;
  LAYER M2 ;
        RECT 6.284 14.66 8.756 14.692 ;
  LAYER M2 ;
        RECT 6.284 14.596 8.756 14.628 ;
  LAYER M2 ;
        RECT 6.284 14.532 8.756 14.564 ;
  LAYER M2 ;
        RECT 6.284 14.468 8.756 14.5 ;
  LAYER M2 ;
        RECT 6.284 14.404 8.756 14.436 ;
  LAYER M2 ;
        RECT 6.284 14.34 8.756 14.372 ;
  LAYER M2 ;
        RECT 6.284 14.276 8.756 14.308 ;
  LAYER M2 ;
        RECT 6.284 14.212 8.756 14.244 ;
  LAYER M2 ;
        RECT 6.284 14.148 8.756 14.18 ;
  LAYER M2 ;
        RECT 6.284 14.084 8.756 14.116 ;
  LAYER M2 ;
        RECT 6.284 14.02 8.756 14.052 ;
  LAYER M2 ;
        RECT 6.284 13.956 8.756 13.988 ;
  LAYER M2 ;
        RECT 6.284 13.892 8.756 13.924 ;
  LAYER M3 ;
        RECT 8.704 13.74 8.736 16.248 ;
  LAYER M3 ;
        RECT 8.64 13.74 8.672 16.248 ;
  LAYER M3 ;
        RECT 8.576 13.74 8.608 16.248 ;
  LAYER M3 ;
        RECT 8.512 13.74 8.544 16.248 ;
  LAYER M3 ;
        RECT 8.448 13.74 8.48 16.248 ;
  LAYER M3 ;
        RECT 8.384 13.74 8.416 16.248 ;
  LAYER M3 ;
        RECT 8.32 13.74 8.352 16.248 ;
  LAYER M3 ;
        RECT 8.256 13.74 8.288 16.248 ;
  LAYER M3 ;
        RECT 8.192 13.74 8.224 16.248 ;
  LAYER M3 ;
        RECT 8.128 13.74 8.16 16.248 ;
  LAYER M3 ;
        RECT 8.064 13.74 8.096 16.248 ;
  LAYER M3 ;
        RECT 8 13.74 8.032 16.248 ;
  LAYER M3 ;
        RECT 7.936 13.74 7.968 16.248 ;
  LAYER M3 ;
        RECT 7.872 13.74 7.904 16.248 ;
  LAYER M3 ;
        RECT 7.808 13.74 7.84 16.248 ;
  LAYER M3 ;
        RECT 7.744 13.74 7.776 16.248 ;
  LAYER M3 ;
        RECT 7.68 13.74 7.712 16.248 ;
  LAYER M3 ;
        RECT 7.616 13.74 7.648 16.248 ;
  LAYER M3 ;
        RECT 7.552 13.74 7.584 16.248 ;
  LAYER M3 ;
        RECT 7.488 13.74 7.52 16.248 ;
  LAYER M3 ;
        RECT 7.424 13.74 7.456 16.248 ;
  LAYER M3 ;
        RECT 7.36 13.74 7.392 16.248 ;
  LAYER M3 ;
        RECT 7.296 13.74 7.328 16.248 ;
  LAYER M3 ;
        RECT 7.232 13.74 7.264 16.248 ;
  LAYER M3 ;
        RECT 7.168 13.74 7.2 16.248 ;
  LAYER M3 ;
        RECT 7.104 13.74 7.136 16.248 ;
  LAYER M3 ;
        RECT 7.04 13.74 7.072 16.248 ;
  LAYER M3 ;
        RECT 6.976 13.74 7.008 16.248 ;
  LAYER M3 ;
        RECT 6.912 13.74 6.944 16.248 ;
  LAYER M3 ;
        RECT 6.848 13.74 6.88 16.248 ;
  LAYER M3 ;
        RECT 6.784 13.74 6.816 16.248 ;
  LAYER M3 ;
        RECT 6.72 13.74 6.752 16.248 ;
  LAYER M3 ;
        RECT 6.656 13.74 6.688 16.248 ;
  LAYER M3 ;
        RECT 6.592 13.74 6.624 16.248 ;
  LAYER M3 ;
        RECT 6.528 13.74 6.56 16.248 ;
  LAYER M3 ;
        RECT 6.464 13.74 6.496 16.248 ;
  LAYER M3 ;
        RECT 6.4 13.74 6.432 16.248 ;
  LAYER M3 ;
        RECT 6.304 13.74 6.336 16.248 ;
  LAYER M1 ;
        RECT 8.719 13.776 8.721 16.212 ;
  LAYER M1 ;
        RECT 8.639 13.776 8.641 16.212 ;
  LAYER M1 ;
        RECT 8.559 13.776 8.561 16.212 ;
  LAYER M1 ;
        RECT 8.479 13.776 8.481 16.212 ;
  LAYER M1 ;
        RECT 8.399 13.776 8.401 16.212 ;
  LAYER M1 ;
        RECT 8.319 13.776 8.321 16.212 ;
  LAYER M1 ;
        RECT 8.239 13.776 8.241 16.212 ;
  LAYER M1 ;
        RECT 8.159 13.776 8.161 16.212 ;
  LAYER M1 ;
        RECT 8.079 13.776 8.081 16.212 ;
  LAYER M1 ;
        RECT 7.999 13.776 8.001 16.212 ;
  LAYER M1 ;
        RECT 7.919 13.776 7.921 16.212 ;
  LAYER M1 ;
        RECT 7.839 13.776 7.841 16.212 ;
  LAYER M1 ;
        RECT 7.759 13.776 7.761 16.212 ;
  LAYER M1 ;
        RECT 7.679 13.776 7.681 16.212 ;
  LAYER M1 ;
        RECT 7.599 13.776 7.601 16.212 ;
  LAYER M1 ;
        RECT 7.519 13.776 7.521 16.212 ;
  LAYER M1 ;
        RECT 7.439 13.776 7.441 16.212 ;
  LAYER M1 ;
        RECT 7.359 13.776 7.361 16.212 ;
  LAYER M1 ;
        RECT 7.279 13.776 7.281 16.212 ;
  LAYER M1 ;
        RECT 7.199 13.776 7.201 16.212 ;
  LAYER M1 ;
        RECT 7.119 13.776 7.121 16.212 ;
  LAYER M1 ;
        RECT 7.039 13.776 7.041 16.212 ;
  LAYER M1 ;
        RECT 6.959 13.776 6.961 16.212 ;
  LAYER M1 ;
        RECT 6.879 13.776 6.881 16.212 ;
  LAYER M1 ;
        RECT 6.799 13.776 6.801 16.212 ;
  LAYER M1 ;
        RECT 6.719 13.776 6.721 16.212 ;
  LAYER M1 ;
        RECT 6.639 13.776 6.641 16.212 ;
  LAYER M1 ;
        RECT 6.559 13.776 6.561 16.212 ;
  LAYER M1 ;
        RECT 6.479 13.776 6.481 16.212 ;
  LAYER M1 ;
        RECT 6.399 13.776 6.401 16.212 ;
  LAYER M2 ;
        RECT 6.32 16.211 8.72 16.213 ;
  LAYER M2 ;
        RECT 6.32 16.127 8.72 16.129 ;
  LAYER M2 ;
        RECT 6.32 16.043 8.72 16.045 ;
  LAYER M2 ;
        RECT 6.32 15.959 8.72 15.961 ;
  LAYER M2 ;
        RECT 6.32 15.875 8.72 15.877 ;
  LAYER M2 ;
        RECT 6.32 15.791 8.72 15.793 ;
  LAYER M2 ;
        RECT 6.32 15.707 8.72 15.709 ;
  LAYER M2 ;
        RECT 6.32 15.623 8.72 15.625 ;
  LAYER M2 ;
        RECT 6.32 15.539 8.72 15.541 ;
  LAYER M2 ;
        RECT 6.32 15.455 8.72 15.457 ;
  LAYER M2 ;
        RECT 6.32 15.371 8.72 15.373 ;
  LAYER M2 ;
        RECT 6.32 15.287 8.72 15.289 ;
  LAYER M2 ;
        RECT 6.32 15.2035 8.72 15.2055 ;
  LAYER M2 ;
        RECT 6.32 15.119 8.72 15.121 ;
  LAYER M2 ;
        RECT 6.32 15.035 8.72 15.037 ;
  LAYER M2 ;
        RECT 6.32 14.951 8.72 14.953 ;
  LAYER M2 ;
        RECT 6.32 14.867 8.72 14.869 ;
  LAYER M2 ;
        RECT 6.32 14.783 8.72 14.785 ;
  LAYER M2 ;
        RECT 6.32 14.699 8.72 14.701 ;
  LAYER M2 ;
        RECT 6.32 14.615 8.72 14.617 ;
  LAYER M2 ;
        RECT 6.32 14.531 8.72 14.533 ;
  LAYER M2 ;
        RECT 6.32 14.447 8.72 14.449 ;
  LAYER M2 ;
        RECT 6.32 14.363 8.72 14.365 ;
  LAYER M2 ;
        RECT 6.32 14.279 8.72 14.281 ;
  LAYER M2 ;
        RECT 6.32 14.195 8.72 14.197 ;
  LAYER M2 ;
        RECT 6.32 14.111 8.72 14.113 ;
  LAYER M2 ;
        RECT 6.32 14.027 8.72 14.029 ;
  LAYER M2 ;
        RECT 6.32 13.943 8.72 13.945 ;
  LAYER M2 ;
        RECT 6.32 13.859 8.72 13.861 ;
  LAYER M1 ;
        RECT 8.704 10.8 8.736 13.308 ;
  LAYER M1 ;
        RECT 8.64 10.8 8.672 13.308 ;
  LAYER M1 ;
        RECT 8.576 10.8 8.608 13.308 ;
  LAYER M1 ;
        RECT 8.512 10.8 8.544 13.308 ;
  LAYER M1 ;
        RECT 8.448 10.8 8.48 13.308 ;
  LAYER M1 ;
        RECT 8.384 10.8 8.416 13.308 ;
  LAYER M1 ;
        RECT 8.32 10.8 8.352 13.308 ;
  LAYER M1 ;
        RECT 8.256 10.8 8.288 13.308 ;
  LAYER M1 ;
        RECT 8.192 10.8 8.224 13.308 ;
  LAYER M1 ;
        RECT 8.128 10.8 8.16 13.308 ;
  LAYER M1 ;
        RECT 8.064 10.8 8.096 13.308 ;
  LAYER M1 ;
        RECT 8 10.8 8.032 13.308 ;
  LAYER M1 ;
        RECT 7.936 10.8 7.968 13.308 ;
  LAYER M1 ;
        RECT 7.872 10.8 7.904 13.308 ;
  LAYER M1 ;
        RECT 7.808 10.8 7.84 13.308 ;
  LAYER M1 ;
        RECT 7.744 10.8 7.776 13.308 ;
  LAYER M1 ;
        RECT 7.68 10.8 7.712 13.308 ;
  LAYER M1 ;
        RECT 7.616 10.8 7.648 13.308 ;
  LAYER M1 ;
        RECT 7.552 10.8 7.584 13.308 ;
  LAYER M1 ;
        RECT 7.488 10.8 7.52 13.308 ;
  LAYER M1 ;
        RECT 7.424 10.8 7.456 13.308 ;
  LAYER M1 ;
        RECT 7.36 10.8 7.392 13.308 ;
  LAYER M1 ;
        RECT 7.296 10.8 7.328 13.308 ;
  LAYER M1 ;
        RECT 7.232 10.8 7.264 13.308 ;
  LAYER M1 ;
        RECT 7.168 10.8 7.2 13.308 ;
  LAYER M1 ;
        RECT 7.104 10.8 7.136 13.308 ;
  LAYER M1 ;
        RECT 7.04 10.8 7.072 13.308 ;
  LAYER M1 ;
        RECT 6.976 10.8 7.008 13.308 ;
  LAYER M1 ;
        RECT 6.912 10.8 6.944 13.308 ;
  LAYER M1 ;
        RECT 6.848 10.8 6.88 13.308 ;
  LAYER M1 ;
        RECT 6.784 10.8 6.816 13.308 ;
  LAYER M1 ;
        RECT 6.72 10.8 6.752 13.308 ;
  LAYER M1 ;
        RECT 6.656 10.8 6.688 13.308 ;
  LAYER M1 ;
        RECT 6.592 10.8 6.624 13.308 ;
  LAYER M1 ;
        RECT 6.528 10.8 6.56 13.308 ;
  LAYER M1 ;
        RECT 6.464 10.8 6.496 13.308 ;
  LAYER M1 ;
        RECT 6.4 10.8 6.432 13.308 ;
  LAYER M2 ;
        RECT 6.284 13.192 8.756 13.224 ;
  LAYER M2 ;
        RECT 6.284 13.128 8.756 13.16 ;
  LAYER M2 ;
        RECT 6.284 13.064 8.756 13.096 ;
  LAYER M2 ;
        RECT 6.284 13 8.756 13.032 ;
  LAYER M2 ;
        RECT 6.284 12.936 8.756 12.968 ;
  LAYER M2 ;
        RECT 6.284 12.872 8.756 12.904 ;
  LAYER M2 ;
        RECT 6.284 12.808 8.756 12.84 ;
  LAYER M2 ;
        RECT 6.284 12.744 8.756 12.776 ;
  LAYER M2 ;
        RECT 6.284 12.68 8.756 12.712 ;
  LAYER M2 ;
        RECT 6.284 12.616 8.756 12.648 ;
  LAYER M2 ;
        RECT 6.284 12.552 8.756 12.584 ;
  LAYER M2 ;
        RECT 6.284 12.488 8.756 12.52 ;
  LAYER M2 ;
        RECT 6.284 12.424 8.756 12.456 ;
  LAYER M2 ;
        RECT 6.284 12.36 8.756 12.392 ;
  LAYER M2 ;
        RECT 6.284 12.296 8.756 12.328 ;
  LAYER M2 ;
        RECT 6.284 12.232 8.756 12.264 ;
  LAYER M2 ;
        RECT 6.284 12.168 8.756 12.2 ;
  LAYER M2 ;
        RECT 6.284 12.104 8.756 12.136 ;
  LAYER M2 ;
        RECT 6.284 12.04 8.756 12.072 ;
  LAYER M2 ;
        RECT 6.284 11.976 8.756 12.008 ;
  LAYER M2 ;
        RECT 6.284 11.912 8.756 11.944 ;
  LAYER M2 ;
        RECT 6.284 11.848 8.756 11.88 ;
  LAYER M2 ;
        RECT 6.284 11.784 8.756 11.816 ;
  LAYER M2 ;
        RECT 6.284 11.72 8.756 11.752 ;
  LAYER M2 ;
        RECT 6.284 11.656 8.756 11.688 ;
  LAYER M2 ;
        RECT 6.284 11.592 8.756 11.624 ;
  LAYER M2 ;
        RECT 6.284 11.528 8.756 11.56 ;
  LAYER M2 ;
        RECT 6.284 11.464 8.756 11.496 ;
  LAYER M2 ;
        RECT 6.284 11.4 8.756 11.432 ;
  LAYER M2 ;
        RECT 6.284 11.336 8.756 11.368 ;
  LAYER M2 ;
        RECT 6.284 11.272 8.756 11.304 ;
  LAYER M2 ;
        RECT 6.284 11.208 8.756 11.24 ;
  LAYER M2 ;
        RECT 6.284 11.144 8.756 11.176 ;
  LAYER M2 ;
        RECT 6.284 11.08 8.756 11.112 ;
  LAYER M2 ;
        RECT 6.284 11.016 8.756 11.048 ;
  LAYER M2 ;
        RECT 6.284 10.952 8.756 10.984 ;
  LAYER M3 ;
        RECT 8.704 10.8 8.736 13.308 ;
  LAYER M3 ;
        RECT 8.64 10.8 8.672 13.308 ;
  LAYER M3 ;
        RECT 8.576 10.8 8.608 13.308 ;
  LAYER M3 ;
        RECT 8.512 10.8 8.544 13.308 ;
  LAYER M3 ;
        RECT 8.448 10.8 8.48 13.308 ;
  LAYER M3 ;
        RECT 8.384 10.8 8.416 13.308 ;
  LAYER M3 ;
        RECT 8.32 10.8 8.352 13.308 ;
  LAYER M3 ;
        RECT 8.256 10.8 8.288 13.308 ;
  LAYER M3 ;
        RECT 8.192 10.8 8.224 13.308 ;
  LAYER M3 ;
        RECT 8.128 10.8 8.16 13.308 ;
  LAYER M3 ;
        RECT 8.064 10.8 8.096 13.308 ;
  LAYER M3 ;
        RECT 8 10.8 8.032 13.308 ;
  LAYER M3 ;
        RECT 7.936 10.8 7.968 13.308 ;
  LAYER M3 ;
        RECT 7.872 10.8 7.904 13.308 ;
  LAYER M3 ;
        RECT 7.808 10.8 7.84 13.308 ;
  LAYER M3 ;
        RECT 7.744 10.8 7.776 13.308 ;
  LAYER M3 ;
        RECT 7.68 10.8 7.712 13.308 ;
  LAYER M3 ;
        RECT 7.616 10.8 7.648 13.308 ;
  LAYER M3 ;
        RECT 7.552 10.8 7.584 13.308 ;
  LAYER M3 ;
        RECT 7.488 10.8 7.52 13.308 ;
  LAYER M3 ;
        RECT 7.424 10.8 7.456 13.308 ;
  LAYER M3 ;
        RECT 7.36 10.8 7.392 13.308 ;
  LAYER M3 ;
        RECT 7.296 10.8 7.328 13.308 ;
  LAYER M3 ;
        RECT 7.232 10.8 7.264 13.308 ;
  LAYER M3 ;
        RECT 7.168 10.8 7.2 13.308 ;
  LAYER M3 ;
        RECT 7.104 10.8 7.136 13.308 ;
  LAYER M3 ;
        RECT 7.04 10.8 7.072 13.308 ;
  LAYER M3 ;
        RECT 6.976 10.8 7.008 13.308 ;
  LAYER M3 ;
        RECT 6.912 10.8 6.944 13.308 ;
  LAYER M3 ;
        RECT 6.848 10.8 6.88 13.308 ;
  LAYER M3 ;
        RECT 6.784 10.8 6.816 13.308 ;
  LAYER M3 ;
        RECT 6.72 10.8 6.752 13.308 ;
  LAYER M3 ;
        RECT 6.656 10.8 6.688 13.308 ;
  LAYER M3 ;
        RECT 6.592 10.8 6.624 13.308 ;
  LAYER M3 ;
        RECT 6.528 10.8 6.56 13.308 ;
  LAYER M3 ;
        RECT 6.464 10.8 6.496 13.308 ;
  LAYER M3 ;
        RECT 6.4 10.8 6.432 13.308 ;
  LAYER M3 ;
        RECT 6.304 10.8 6.336 13.308 ;
  LAYER M1 ;
        RECT 8.719 10.836 8.721 13.272 ;
  LAYER M1 ;
        RECT 8.639 10.836 8.641 13.272 ;
  LAYER M1 ;
        RECT 8.559 10.836 8.561 13.272 ;
  LAYER M1 ;
        RECT 8.479 10.836 8.481 13.272 ;
  LAYER M1 ;
        RECT 8.399 10.836 8.401 13.272 ;
  LAYER M1 ;
        RECT 8.319 10.836 8.321 13.272 ;
  LAYER M1 ;
        RECT 8.239 10.836 8.241 13.272 ;
  LAYER M1 ;
        RECT 8.159 10.836 8.161 13.272 ;
  LAYER M1 ;
        RECT 8.079 10.836 8.081 13.272 ;
  LAYER M1 ;
        RECT 7.999 10.836 8.001 13.272 ;
  LAYER M1 ;
        RECT 7.919 10.836 7.921 13.272 ;
  LAYER M1 ;
        RECT 7.839 10.836 7.841 13.272 ;
  LAYER M1 ;
        RECT 7.759 10.836 7.761 13.272 ;
  LAYER M1 ;
        RECT 7.679 10.836 7.681 13.272 ;
  LAYER M1 ;
        RECT 7.599 10.836 7.601 13.272 ;
  LAYER M1 ;
        RECT 7.519 10.836 7.521 13.272 ;
  LAYER M1 ;
        RECT 7.439 10.836 7.441 13.272 ;
  LAYER M1 ;
        RECT 7.359 10.836 7.361 13.272 ;
  LAYER M1 ;
        RECT 7.279 10.836 7.281 13.272 ;
  LAYER M1 ;
        RECT 7.199 10.836 7.201 13.272 ;
  LAYER M1 ;
        RECT 7.119 10.836 7.121 13.272 ;
  LAYER M1 ;
        RECT 7.039 10.836 7.041 13.272 ;
  LAYER M1 ;
        RECT 6.959 10.836 6.961 13.272 ;
  LAYER M1 ;
        RECT 6.879 10.836 6.881 13.272 ;
  LAYER M1 ;
        RECT 6.799 10.836 6.801 13.272 ;
  LAYER M1 ;
        RECT 6.719 10.836 6.721 13.272 ;
  LAYER M1 ;
        RECT 6.639 10.836 6.641 13.272 ;
  LAYER M1 ;
        RECT 6.559 10.836 6.561 13.272 ;
  LAYER M1 ;
        RECT 6.479 10.836 6.481 13.272 ;
  LAYER M1 ;
        RECT 6.399 10.836 6.401 13.272 ;
  LAYER M2 ;
        RECT 6.32 13.271 8.72 13.273 ;
  LAYER M2 ;
        RECT 6.32 13.187 8.72 13.189 ;
  LAYER M2 ;
        RECT 6.32 13.103 8.72 13.105 ;
  LAYER M2 ;
        RECT 6.32 13.019 8.72 13.021 ;
  LAYER M2 ;
        RECT 6.32 12.935 8.72 12.937 ;
  LAYER M2 ;
        RECT 6.32 12.851 8.72 12.853 ;
  LAYER M2 ;
        RECT 6.32 12.767 8.72 12.769 ;
  LAYER M2 ;
        RECT 6.32 12.683 8.72 12.685 ;
  LAYER M2 ;
        RECT 6.32 12.599 8.72 12.601 ;
  LAYER M2 ;
        RECT 6.32 12.515 8.72 12.517 ;
  LAYER M2 ;
        RECT 6.32 12.431 8.72 12.433 ;
  LAYER M2 ;
        RECT 6.32 12.347 8.72 12.349 ;
  LAYER M2 ;
        RECT 6.32 12.2635 8.72 12.2655 ;
  LAYER M2 ;
        RECT 6.32 12.179 8.72 12.181 ;
  LAYER M2 ;
        RECT 6.32 12.095 8.72 12.097 ;
  LAYER M2 ;
        RECT 6.32 12.011 8.72 12.013 ;
  LAYER M2 ;
        RECT 6.32 11.927 8.72 11.929 ;
  LAYER M2 ;
        RECT 6.32 11.843 8.72 11.845 ;
  LAYER M2 ;
        RECT 6.32 11.759 8.72 11.761 ;
  LAYER M2 ;
        RECT 6.32 11.675 8.72 11.677 ;
  LAYER M2 ;
        RECT 6.32 11.591 8.72 11.593 ;
  LAYER M2 ;
        RECT 6.32 11.507 8.72 11.509 ;
  LAYER M2 ;
        RECT 6.32 11.423 8.72 11.425 ;
  LAYER M2 ;
        RECT 6.32 11.339 8.72 11.341 ;
  LAYER M2 ;
        RECT 6.32 11.255 8.72 11.257 ;
  LAYER M2 ;
        RECT 6.32 11.171 8.72 11.173 ;
  LAYER M2 ;
        RECT 6.32 11.087 8.72 11.089 ;
  LAYER M2 ;
        RECT 6.32 11.003 8.72 11.005 ;
  LAYER M2 ;
        RECT 6.32 10.919 8.72 10.921 ;
  LAYER M1 ;
        RECT 8.704 7.86 8.736 10.368 ;
  LAYER M1 ;
        RECT 8.64 7.86 8.672 10.368 ;
  LAYER M1 ;
        RECT 8.576 7.86 8.608 10.368 ;
  LAYER M1 ;
        RECT 8.512 7.86 8.544 10.368 ;
  LAYER M1 ;
        RECT 8.448 7.86 8.48 10.368 ;
  LAYER M1 ;
        RECT 8.384 7.86 8.416 10.368 ;
  LAYER M1 ;
        RECT 8.32 7.86 8.352 10.368 ;
  LAYER M1 ;
        RECT 8.256 7.86 8.288 10.368 ;
  LAYER M1 ;
        RECT 8.192 7.86 8.224 10.368 ;
  LAYER M1 ;
        RECT 8.128 7.86 8.16 10.368 ;
  LAYER M1 ;
        RECT 8.064 7.86 8.096 10.368 ;
  LAYER M1 ;
        RECT 8 7.86 8.032 10.368 ;
  LAYER M1 ;
        RECT 7.936 7.86 7.968 10.368 ;
  LAYER M1 ;
        RECT 7.872 7.86 7.904 10.368 ;
  LAYER M1 ;
        RECT 7.808 7.86 7.84 10.368 ;
  LAYER M1 ;
        RECT 7.744 7.86 7.776 10.368 ;
  LAYER M1 ;
        RECT 7.68 7.86 7.712 10.368 ;
  LAYER M1 ;
        RECT 7.616 7.86 7.648 10.368 ;
  LAYER M1 ;
        RECT 7.552 7.86 7.584 10.368 ;
  LAYER M1 ;
        RECT 7.488 7.86 7.52 10.368 ;
  LAYER M1 ;
        RECT 7.424 7.86 7.456 10.368 ;
  LAYER M1 ;
        RECT 7.36 7.86 7.392 10.368 ;
  LAYER M1 ;
        RECT 7.296 7.86 7.328 10.368 ;
  LAYER M1 ;
        RECT 7.232 7.86 7.264 10.368 ;
  LAYER M1 ;
        RECT 7.168 7.86 7.2 10.368 ;
  LAYER M1 ;
        RECT 7.104 7.86 7.136 10.368 ;
  LAYER M1 ;
        RECT 7.04 7.86 7.072 10.368 ;
  LAYER M1 ;
        RECT 6.976 7.86 7.008 10.368 ;
  LAYER M1 ;
        RECT 6.912 7.86 6.944 10.368 ;
  LAYER M1 ;
        RECT 6.848 7.86 6.88 10.368 ;
  LAYER M1 ;
        RECT 6.784 7.86 6.816 10.368 ;
  LAYER M1 ;
        RECT 6.72 7.86 6.752 10.368 ;
  LAYER M1 ;
        RECT 6.656 7.86 6.688 10.368 ;
  LAYER M1 ;
        RECT 6.592 7.86 6.624 10.368 ;
  LAYER M1 ;
        RECT 6.528 7.86 6.56 10.368 ;
  LAYER M1 ;
        RECT 6.464 7.86 6.496 10.368 ;
  LAYER M1 ;
        RECT 6.4 7.86 6.432 10.368 ;
  LAYER M2 ;
        RECT 6.284 10.252 8.756 10.284 ;
  LAYER M2 ;
        RECT 6.284 10.188 8.756 10.22 ;
  LAYER M2 ;
        RECT 6.284 10.124 8.756 10.156 ;
  LAYER M2 ;
        RECT 6.284 10.06 8.756 10.092 ;
  LAYER M2 ;
        RECT 6.284 9.996 8.756 10.028 ;
  LAYER M2 ;
        RECT 6.284 9.932 8.756 9.964 ;
  LAYER M2 ;
        RECT 6.284 9.868 8.756 9.9 ;
  LAYER M2 ;
        RECT 6.284 9.804 8.756 9.836 ;
  LAYER M2 ;
        RECT 6.284 9.74 8.756 9.772 ;
  LAYER M2 ;
        RECT 6.284 9.676 8.756 9.708 ;
  LAYER M2 ;
        RECT 6.284 9.612 8.756 9.644 ;
  LAYER M2 ;
        RECT 6.284 9.548 8.756 9.58 ;
  LAYER M2 ;
        RECT 6.284 9.484 8.756 9.516 ;
  LAYER M2 ;
        RECT 6.284 9.42 8.756 9.452 ;
  LAYER M2 ;
        RECT 6.284 9.356 8.756 9.388 ;
  LAYER M2 ;
        RECT 6.284 9.292 8.756 9.324 ;
  LAYER M2 ;
        RECT 6.284 9.228 8.756 9.26 ;
  LAYER M2 ;
        RECT 6.284 9.164 8.756 9.196 ;
  LAYER M2 ;
        RECT 6.284 9.1 8.756 9.132 ;
  LAYER M2 ;
        RECT 6.284 9.036 8.756 9.068 ;
  LAYER M2 ;
        RECT 6.284 8.972 8.756 9.004 ;
  LAYER M2 ;
        RECT 6.284 8.908 8.756 8.94 ;
  LAYER M2 ;
        RECT 6.284 8.844 8.756 8.876 ;
  LAYER M2 ;
        RECT 6.284 8.78 8.756 8.812 ;
  LAYER M2 ;
        RECT 6.284 8.716 8.756 8.748 ;
  LAYER M2 ;
        RECT 6.284 8.652 8.756 8.684 ;
  LAYER M2 ;
        RECT 6.284 8.588 8.756 8.62 ;
  LAYER M2 ;
        RECT 6.284 8.524 8.756 8.556 ;
  LAYER M2 ;
        RECT 6.284 8.46 8.756 8.492 ;
  LAYER M2 ;
        RECT 6.284 8.396 8.756 8.428 ;
  LAYER M2 ;
        RECT 6.284 8.332 8.756 8.364 ;
  LAYER M2 ;
        RECT 6.284 8.268 8.756 8.3 ;
  LAYER M2 ;
        RECT 6.284 8.204 8.756 8.236 ;
  LAYER M2 ;
        RECT 6.284 8.14 8.756 8.172 ;
  LAYER M2 ;
        RECT 6.284 8.076 8.756 8.108 ;
  LAYER M2 ;
        RECT 6.284 8.012 8.756 8.044 ;
  LAYER M3 ;
        RECT 8.704 7.86 8.736 10.368 ;
  LAYER M3 ;
        RECT 8.64 7.86 8.672 10.368 ;
  LAYER M3 ;
        RECT 8.576 7.86 8.608 10.368 ;
  LAYER M3 ;
        RECT 8.512 7.86 8.544 10.368 ;
  LAYER M3 ;
        RECT 8.448 7.86 8.48 10.368 ;
  LAYER M3 ;
        RECT 8.384 7.86 8.416 10.368 ;
  LAYER M3 ;
        RECT 8.32 7.86 8.352 10.368 ;
  LAYER M3 ;
        RECT 8.256 7.86 8.288 10.368 ;
  LAYER M3 ;
        RECT 8.192 7.86 8.224 10.368 ;
  LAYER M3 ;
        RECT 8.128 7.86 8.16 10.368 ;
  LAYER M3 ;
        RECT 8.064 7.86 8.096 10.368 ;
  LAYER M3 ;
        RECT 8 7.86 8.032 10.368 ;
  LAYER M3 ;
        RECT 7.936 7.86 7.968 10.368 ;
  LAYER M3 ;
        RECT 7.872 7.86 7.904 10.368 ;
  LAYER M3 ;
        RECT 7.808 7.86 7.84 10.368 ;
  LAYER M3 ;
        RECT 7.744 7.86 7.776 10.368 ;
  LAYER M3 ;
        RECT 7.68 7.86 7.712 10.368 ;
  LAYER M3 ;
        RECT 7.616 7.86 7.648 10.368 ;
  LAYER M3 ;
        RECT 7.552 7.86 7.584 10.368 ;
  LAYER M3 ;
        RECT 7.488 7.86 7.52 10.368 ;
  LAYER M3 ;
        RECT 7.424 7.86 7.456 10.368 ;
  LAYER M3 ;
        RECT 7.36 7.86 7.392 10.368 ;
  LAYER M3 ;
        RECT 7.296 7.86 7.328 10.368 ;
  LAYER M3 ;
        RECT 7.232 7.86 7.264 10.368 ;
  LAYER M3 ;
        RECT 7.168 7.86 7.2 10.368 ;
  LAYER M3 ;
        RECT 7.104 7.86 7.136 10.368 ;
  LAYER M3 ;
        RECT 7.04 7.86 7.072 10.368 ;
  LAYER M3 ;
        RECT 6.976 7.86 7.008 10.368 ;
  LAYER M3 ;
        RECT 6.912 7.86 6.944 10.368 ;
  LAYER M3 ;
        RECT 6.848 7.86 6.88 10.368 ;
  LAYER M3 ;
        RECT 6.784 7.86 6.816 10.368 ;
  LAYER M3 ;
        RECT 6.72 7.86 6.752 10.368 ;
  LAYER M3 ;
        RECT 6.656 7.86 6.688 10.368 ;
  LAYER M3 ;
        RECT 6.592 7.86 6.624 10.368 ;
  LAYER M3 ;
        RECT 6.528 7.86 6.56 10.368 ;
  LAYER M3 ;
        RECT 6.464 7.86 6.496 10.368 ;
  LAYER M3 ;
        RECT 6.4 7.86 6.432 10.368 ;
  LAYER M3 ;
        RECT 6.304 7.86 6.336 10.368 ;
  LAYER M1 ;
        RECT 8.719 7.896 8.721 10.332 ;
  LAYER M1 ;
        RECT 8.639 7.896 8.641 10.332 ;
  LAYER M1 ;
        RECT 8.559 7.896 8.561 10.332 ;
  LAYER M1 ;
        RECT 8.479 7.896 8.481 10.332 ;
  LAYER M1 ;
        RECT 8.399 7.896 8.401 10.332 ;
  LAYER M1 ;
        RECT 8.319 7.896 8.321 10.332 ;
  LAYER M1 ;
        RECT 8.239 7.896 8.241 10.332 ;
  LAYER M1 ;
        RECT 8.159 7.896 8.161 10.332 ;
  LAYER M1 ;
        RECT 8.079 7.896 8.081 10.332 ;
  LAYER M1 ;
        RECT 7.999 7.896 8.001 10.332 ;
  LAYER M1 ;
        RECT 7.919 7.896 7.921 10.332 ;
  LAYER M1 ;
        RECT 7.839 7.896 7.841 10.332 ;
  LAYER M1 ;
        RECT 7.759 7.896 7.761 10.332 ;
  LAYER M1 ;
        RECT 7.679 7.896 7.681 10.332 ;
  LAYER M1 ;
        RECT 7.599 7.896 7.601 10.332 ;
  LAYER M1 ;
        RECT 7.519 7.896 7.521 10.332 ;
  LAYER M1 ;
        RECT 7.439 7.896 7.441 10.332 ;
  LAYER M1 ;
        RECT 7.359 7.896 7.361 10.332 ;
  LAYER M1 ;
        RECT 7.279 7.896 7.281 10.332 ;
  LAYER M1 ;
        RECT 7.199 7.896 7.201 10.332 ;
  LAYER M1 ;
        RECT 7.119 7.896 7.121 10.332 ;
  LAYER M1 ;
        RECT 7.039 7.896 7.041 10.332 ;
  LAYER M1 ;
        RECT 6.959 7.896 6.961 10.332 ;
  LAYER M1 ;
        RECT 6.879 7.896 6.881 10.332 ;
  LAYER M1 ;
        RECT 6.799 7.896 6.801 10.332 ;
  LAYER M1 ;
        RECT 6.719 7.896 6.721 10.332 ;
  LAYER M1 ;
        RECT 6.639 7.896 6.641 10.332 ;
  LAYER M1 ;
        RECT 6.559 7.896 6.561 10.332 ;
  LAYER M1 ;
        RECT 6.479 7.896 6.481 10.332 ;
  LAYER M1 ;
        RECT 6.399 7.896 6.401 10.332 ;
  LAYER M2 ;
        RECT 6.32 10.331 8.72 10.333 ;
  LAYER M2 ;
        RECT 6.32 10.247 8.72 10.249 ;
  LAYER M2 ;
        RECT 6.32 10.163 8.72 10.165 ;
  LAYER M2 ;
        RECT 6.32 10.079 8.72 10.081 ;
  LAYER M2 ;
        RECT 6.32 9.995 8.72 9.997 ;
  LAYER M2 ;
        RECT 6.32 9.911 8.72 9.913 ;
  LAYER M2 ;
        RECT 6.32 9.827 8.72 9.829 ;
  LAYER M2 ;
        RECT 6.32 9.743 8.72 9.745 ;
  LAYER M2 ;
        RECT 6.32 9.659 8.72 9.661 ;
  LAYER M2 ;
        RECT 6.32 9.575 8.72 9.577 ;
  LAYER M2 ;
        RECT 6.32 9.491 8.72 9.493 ;
  LAYER M2 ;
        RECT 6.32 9.407 8.72 9.409 ;
  LAYER M2 ;
        RECT 6.32 9.3235 8.72 9.3255 ;
  LAYER M2 ;
        RECT 6.32 9.239 8.72 9.241 ;
  LAYER M2 ;
        RECT 6.32 9.155 8.72 9.157 ;
  LAYER M2 ;
        RECT 6.32 9.071 8.72 9.073 ;
  LAYER M2 ;
        RECT 6.32 8.987 8.72 8.989 ;
  LAYER M2 ;
        RECT 6.32 8.903 8.72 8.905 ;
  LAYER M2 ;
        RECT 6.32 8.819 8.72 8.821 ;
  LAYER M2 ;
        RECT 6.32 8.735 8.72 8.737 ;
  LAYER M2 ;
        RECT 6.32 8.651 8.72 8.653 ;
  LAYER M2 ;
        RECT 6.32 8.567 8.72 8.569 ;
  LAYER M2 ;
        RECT 6.32 8.483 8.72 8.485 ;
  LAYER M2 ;
        RECT 6.32 8.399 8.72 8.401 ;
  LAYER M2 ;
        RECT 6.32 8.315 8.72 8.317 ;
  LAYER M2 ;
        RECT 6.32 8.231 8.72 8.233 ;
  LAYER M2 ;
        RECT 6.32 8.147 8.72 8.149 ;
  LAYER M2 ;
        RECT 6.32 8.063 8.72 8.065 ;
  LAYER M2 ;
        RECT 6.32 7.979 8.72 7.981 ;
  LAYER M1 ;
        RECT 8.704 4.92 8.736 7.428 ;
  LAYER M1 ;
        RECT 8.64 4.92 8.672 7.428 ;
  LAYER M1 ;
        RECT 8.576 4.92 8.608 7.428 ;
  LAYER M1 ;
        RECT 8.512 4.92 8.544 7.428 ;
  LAYER M1 ;
        RECT 8.448 4.92 8.48 7.428 ;
  LAYER M1 ;
        RECT 8.384 4.92 8.416 7.428 ;
  LAYER M1 ;
        RECT 8.32 4.92 8.352 7.428 ;
  LAYER M1 ;
        RECT 8.256 4.92 8.288 7.428 ;
  LAYER M1 ;
        RECT 8.192 4.92 8.224 7.428 ;
  LAYER M1 ;
        RECT 8.128 4.92 8.16 7.428 ;
  LAYER M1 ;
        RECT 8.064 4.92 8.096 7.428 ;
  LAYER M1 ;
        RECT 8 4.92 8.032 7.428 ;
  LAYER M1 ;
        RECT 7.936 4.92 7.968 7.428 ;
  LAYER M1 ;
        RECT 7.872 4.92 7.904 7.428 ;
  LAYER M1 ;
        RECT 7.808 4.92 7.84 7.428 ;
  LAYER M1 ;
        RECT 7.744 4.92 7.776 7.428 ;
  LAYER M1 ;
        RECT 7.68 4.92 7.712 7.428 ;
  LAYER M1 ;
        RECT 7.616 4.92 7.648 7.428 ;
  LAYER M1 ;
        RECT 7.552 4.92 7.584 7.428 ;
  LAYER M1 ;
        RECT 7.488 4.92 7.52 7.428 ;
  LAYER M1 ;
        RECT 7.424 4.92 7.456 7.428 ;
  LAYER M1 ;
        RECT 7.36 4.92 7.392 7.428 ;
  LAYER M1 ;
        RECT 7.296 4.92 7.328 7.428 ;
  LAYER M1 ;
        RECT 7.232 4.92 7.264 7.428 ;
  LAYER M1 ;
        RECT 7.168 4.92 7.2 7.428 ;
  LAYER M1 ;
        RECT 7.104 4.92 7.136 7.428 ;
  LAYER M1 ;
        RECT 7.04 4.92 7.072 7.428 ;
  LAYER M1 ;
        RECT 6.976 4.92 7.008 7.428 ;
  LAYER M1 ;
        RECT 6.912 4.92 6.944 7.428 ;
  LAYER M1 ;
        RECT 6.848 4.92 6.88 7.428 ;
  LAYER M1 ;
        RECT 6.784 4.92 6.816 7.428 ;
  LAYER M1 ;
        RECT 6.72 4.92 6.752 7.428 ;
  LAYER M1 ;
        RECT 6.656 4.92 6.688 7.428 ;
  LAYER M1 ;
        RECT 6.592 4.92 6.624 7.428 ;
  LAYER M1 ;
        RECT 6.528 4.92 6.56 7.428 ;
  LAYER M1 ;
        RECT 6.464 4.92 6.496 7.428 ;
  LAYER M1 ;
        RECT 6.4 4.92 6.432 7.428 ;
  LAYER M2 ;
        RECT 6.284 7.312 8.756 7.344 ;
  LAYER M2 ;
        RECT 6.284 7.248 8.756 7.28 ;
  LAYER M2 ;
        RECT 6.284 7.184 8.756 7.216 ;
  LAYER M2 ;
        RECT 6.284 7.12 8.756 7.152 ;
  LAYER M2 ;
        RECT 6.284 7.056 8.756 7.088 ;
  LAYER M2 ;
        RECT 6.284 6.992 8.756 7.024 ;
  LAYER M2 ;
        RECT 6.284 6.928 8.756 6.96 ;
  LAYER M2 ;
        RECT 6.284 6.864 8.756 6.896 ;
  LAYER M2 ;
        RECT 6.284 6.8 8.756 6.832 ;
  LAYER M2 ;
        RECT 6.284 6.736 8.756 6.768 ;
  LAYER M2 ;
        RECT 6.284 6.672 8.756 6.704 ;
  LAYER M2 ;
        RECT 6.284 6.608 8.756 6.64 ;
  LAYER M2 ;
        RECT 6.284 6.544 8.756 6.576 ;
  LAYER M2 ;
        RECT 6.284 6.48 8.756 6.512 ;
  LAYER M2 ;
        RECT 6.284 6.416 8.756 6.448 ;
  LAYER M2 ;
        RECT 6.284 6.352 8.756 6.384 ;
  LAYER M2 ;
        RECT 6.284 6.288 8.756 6.32 ;
  LAYER M2 ;
        RECT 6.284 6.224 8.756 6.256 ;
  LAYER M2 ;
        RECT 6.284 6.16 8.756 6.192 ;
  LAYER M2 ;
        RECT 6.284 6.096 8.756 6.128 ;
  LAYER M2 ;
        RECT 6.284 6.032 8.756 6.064 ;
  LAYER M2 ;
        RECT 6.284 5.968 8.756 6 ;
  LAYER M2 ;
        RECT 6.284 5.904 8.756 5.936 ;
  LAYER M2 ;
        RECT 6.284 5.84 8.756 5.872 ;
  LAYER M2 ;
        RECT 6.284 5.776 8.756 5.808 ;
  LAYER M2 ;
        RECT 6.284 5.712 8.756 5.744 ;
  LAYER M2 ;
        RECT 6.284 5.648 8.756 5.68 ;
  LAYER M2 ;
        RECT 6.284 5.584 8.756 5.616 ;
  LAYER M2 ;
        RECT 6.284 5.52 8.756 5.552 ;
  LAYER M2 ;
        RECT 6.284 5.456 8.756 5.488 ;
  LAYER M2 ;
        RECT 6.284 5.392 8.756 5.424 ;
  LAYER M2 ;
        RECT 6.284 5.328 8.756 5.36 ;
  LAYER M2 ;
        RECT 6.284 5.264 8.756 5.296 ;
  LAYER M2 ;
        RECT 6.284 5.2 8.756 5.232 ;
  LAYER M2 ;
        RECT 6.284 5.136 8.756 5.168 ;
  LAYER M2 ;
        RECT 6.284 5.072 8.756 5.104 ;
  LAYER M3 ;
        RECT 8.704 4.92 8.736 7.428 ;
  LAYER M3 ;
        RECT 8.64 4.92 8.672 7.428 ;
  LAYER M3 ;
        RECT 8.576 4.92 8.608 7.428 ;
  LAYER M3 ;
        RECT 8.512 4.92 8.544 7.428 ;
  LAYER M3 ;
        RECT 8.448 4.92 8.48 7.428 ;
  LAYER M3 ;
        RECT 8.384 4.92 8.416 7.428 ;
  LAYER M3 ;
        RECT 8.32 4.92 8.352 7.428 ;
  LAYER M3 ;
        RECT 8.256 4.92 8.288 7.428 ;
  LAYER M3 ;
        RECT 8.192 4.92 8.224 7.428 ;
  LAYER M3 ;
        RECT 8.128 4.92 8.16 7.428 ;
  LAYER M3 ;
        RECT 8.064 4.92 8.096 7.428 ;
  LAYER M3 ;
        RECT 8 4.92 8.032 7.428 ;
  LAYER M3 ;
        RECT 7.936 4.92 7.968 7.428 ;
  LAYER M3 ;
        RECT 7.872 4.92 7.904 7.428 ;
  LAYER M3 ;
        RECT 7.808 4.92 7.84 7.428 ;
  LAYER M3 ;
        RECT 7.744 4.92 7.776 7.428 ;
  LAYER M3 ;
        RECT 7.68 4.92 7.712 7.428 ;
  LAYER M3 ;
        RECT 7.616 4.92 7.648 7.428 ;
  LAYER M3 ;
        RECT 7.552 4.92 7.584 7.428 ;
  LAYER M3 ;
        RECT 7.488 4.92 7.52 7.428 ;
  LAYER M3 ;
        RECT 7.424 4.92 7.456 7.428 ;
  LAYER M3 ;
        RECT 7.36 4.92 7.392 7.428 ;
  LAYER M3 ;
        RECT 7.296 4.92 7.328 7.428 ;
  LAYER M3 ;
        RECT 7.232 4.92 7.264 7.428 ;
  LAYER M3 ;
        RECT 7.168 4.92 7.2 7.428 ;
  LAYER M3 ;
        RECT 7.104 4.92 7.136 7.428 ;
  LAYER M3 ;
        RECT 7.04 4.92 7.072 7.428 ;
  LAYER M3 ;
        RECT 6.976 4.92 7.008 7.428 ;
  LAYER M3 ;
        RECT 6.912 4.92 6.944 7.428 ;
  LAYER M3 ;
        RECT 6.848 4.92 6.88 7.428 ;
  LAYER M3 ;
        RECT 6.784 4.92 6.816 7.428 ;
  LAYER M3 ;
        RECT 6.72 4.92 6.752 7.428 ;
  LAYER M3 ;
        RECT 6.656 4.92 6.688 7.428 ;
  LAYER M3 ;
        RECT 6.592 4.92 6.624 7.428 ;
  LAYER M3 ;
        RECT 6.528 4.92 6.56 7.428 ;
  LAYER M3 ;
        RECT 6.464 4.92 6.496 7.428 ;
  LAYER M3 ;
        RECT 6.4 4.92 6.432 7.428 ;
  LAYER M3 ;
        RECT 6.304 4.92 6.336 7.428 ;
  LAYER M1 ;
        RECT 8.719 4.956 8.721 7.392 ;
  LAYER M1 ;
        RECT 8.639 4.956 8.641 7.392 ;
  LAYER M1 ;
        RECT 8.559 4.956 8.561 7.392 ;
  LAYER M1 ;
        RECT 8.479 4.956 8.481 7.392 ;
  LAYER M1 ;
        RECT 8.399 4.956 8.401 7.392 ;
  LAYER M1 ;
        RECT 8.319 4.956 8.321 7.392 ;
  LAYER M1 ;
        RECT 8.239 4.956 8.241 7.392 ;
  LAYER M1 ;
        RECT 8.159 4.956 8.161 7.392 ;
  LAYER M1 ;
        RECT 8.079 4.956 8.081 7.392 ;
  LAYER M1 ;
        RECT 7.999 4.956 8.001 7.392 ;
  LAYER M1 ;
        RECT 7.919 4.956 7.921 7.392 ;
  LAYER M1 ;
        RECT 7.839 4.956 7.841 7.392 ;
  LAYER M1 ;
        RECT 7.759 4.956 7.761 7.392 ;
  LAYER M1 ;
        RECT 7.679 4.956 7.681 7.392 ;
  LAYER M1 ;
        RECT 7.599 4.956 7.601 7.392 ;
  LAYER M1 ;
        RECT 7.519 4.956 7.521 7.392 ;
  LAYER M1 ;
        RECT 7.439 4.956 7.441 7.392 ;
  LAYER M1 ;
        RECT 7.359 4.956 7.361 7.392 ;
  LAYER M1 ;
        RECT 7.279 4.956 7.281 7.392 ;
  LAYER M1 ;
        RECT 7.199 4.956 7.201 7.392 ;
  LAYER M1 ;
        RECT 7.119 4.956 7.121 7.392 ;
  LAYER M1 ;
        RECT 7.039 4.956 7.041 7.392 ;
  LAYER M1 ;
        RECT 6.959 4.956 6.961 7.392 ;
  LAYER M1 ;
        RECT 6.879 4.956 6.881 7.392 ;
  LAYER M1 ;
        RECT 6.799 4.956 6.801 7.392 ;
  LAYER M1 ;
        RECT 6.719 4.956 6.721 7.392 ;
  LAYER M1 ;
        RECT 6.639 4.956 6.641 7.392 ;
  LAYER M1 ;
        RECT 6.559 4.956 6.561 7.392 ;
  LAYER M1 ;
        RECT 6.479 4.956 6.481 7.392 ;
  LAYER M1 ;
        RECT 6.399 4.956 6.401 7.392 ;
  LAYER M2 ;
        RECT 6.32 7.391 8.72 7.393 ;
  LAYER M2 ;
        RECT 6.32 7.307 8.72 7.309 ;
  LAYER M2 ;
        RECT 6.32 7.223 8.72 7.225 ;
  LAYER M2 ;
        RECT 6.32 7.139 8.72 7.141 ;
  LAYER M2 ;
        RECT 6.32 7.055 8.72 7.057 ;
  LAYER M2 ;
        RECT 6.32 6.971 8.72 6.973 ;
  LAYER M2 ;
        RECT 6.32 6.887 8.72 6.889 ;
  LAYER M2 ;
        RECT 6.32 6.803 8.72 6.805 ;
  LAYER M2 ;
        RECT 6.32 6.719 8.72 6.721 ;
  LAYER M2 ;
        RECT 6.32 6.635 8.72 6.637 ;
  LAYER M2 ;
        RECT 6.32 6.551 8.72 6.553 ;
  LAYER M2 ;
        RECT 6.32 6.467 8.72 6.469 ;
  LAYER M2 ;
        RECT 6.32 6.3835 8.72 6.3855 ;
  LAYER M2 ;
        RECT 6.32 6.299 8.72 6.301 ;
  LAYER M2 ;
        RECT 6.32 6.215 8.72 6.217 ;
  LAYER M2 ;
        RECT 6.32 6.131 8.72 6.133 ;
  LAYER M2 ;
        RECT 6.32 6.047 8.72 6.049 ;
  LAYER M2 ;
        RECT 6.32 5.963 8.72 5.965 ;
  LAYER M2 ;
        RECT 6.32 5.879 8.72 5.881 ;
  LAYER M2 ;
        RECT 6.32 5.795 8.72 5.797 ;
  LAYER M2 ;
        RECT 6.32 5.711 8.72 5.713 ;
  LAYER M2 ;
        RECT 6.32 5.627 8.72 5.629 ;
  LAYER M2 ;
        RECT 6.32 5.543 8.72 5.545 ;
  LAYER M2 ;
        RECT 6.32 5.459 8.72 5.461 ;
  LAYER M2 ;
        RECT 6.32 5.375 8.72 5.377 ;
  LAYER M2 ;
        RECT 6.32 5.291 8.72 5.293 ;
  LAYER M2 ;
        RECT 6.32 5.207 8.72 5.209 ;
  LAYER M2 ;
        RECT 6.32 5.123 8.72 5.125 ;
  LAYER M2 ;
        RECT 6.32 5.039 8.72 5.041 ;
  LAYER M1 ;
        RECT 8.704 1.98 8.736 4.488 ;
  LAYER M1 ;
        RECT 8.64 1.98 8.672 4.488 ;
  LAYER M1 ;
        RECT 8.576 1.98 8.608 4.488 ;
  LAYER M1 ;
        RECT 8.512 1.98 8.544 4.488 ;
  LAYER M1 ;
        RECT 8.448 1.98 8.48 4.488 ;
  LAYER M1 ;
        RECT 8.384 1.98 8.416 4.488 ;
  LAYER M1 ;
        RECT 8.32 1.98 8.352 4.488 ;
  LAYER M1 ;
        RECT 8.256 1.98 8.288 4.488 ;
  LAYER M1 ;
        RECT 8.192 1.98 8.224 4.488 ;
  LAYER M1 ;
        RECT 8.128 1.98 8.16 4.488 ;
  LAYER M1 ;
        RECT 8.064 1.98 8.096 4.488 ;
  LAYER M1 ;
        RECT 8 1.98 8.032 4.488 ;
  LAYER M1 ;
        RECT 7.936 1.98 7.968 4.488 ;
  LAYER M1 ;
        RECT 7.872 1.98 7.904 4.488 ;
  LAYER M1 ;
        RECT 7.808 1.98 7.84 4.488 ;
  LAYER M1 ;
        RECT 7.744 1.98 7.776 4.488 ;
  LAYER M1 ;
        RECT 7.68 1.98 7.712 4.488 ;
  LAYER M1 ;
        RECT 7.616 1.98 7.648 4.488 ;
  LAYER M1 ;
        RECT 7.552 1.98 7.584 4.488 ;
  LAYER M1 ;
        RECT 7.488 1.98 7.52 4.488 ;
  LAYER M1 ;
        RECT 7.424 1.98 7.456 4.488 ;
  LAYER M1 ;
        RECT 7.36 1.98 7.392 4.488 ;
  LAYER M1 ;
        RECT 7.296 1.98 7.328 4.488 ;
  LAYER M1 ;
        RECT 7.232 1.98 7.264 4.488 ;
  LAYER M1 ;
        RECT 7.168 1.98 7.2 4.488 ;
  LAYER M1 ;
        RECT 7.104 1.98 7.136 4.488 ;
  LAYER M1 ;
        RECT 7.04 1.98 7.072 4.488 ;
  LAYER M1 ;
        RECT 6.976 1.98 7.008 4.488 ;
  LAYER M1 ;
        RECT 6.912 1.98 6.944 4.488 ;
  LAYER M1 ;
        RECT 6.848 1.98 6.88 4.488 ;
  LAYER M1 ;
        RECT 6.784 1.98 6.816 4.488 ;
  LAYER M1 ;
        RECT 6.72 1.98 6.752 4.488 ;
  LAYER M1 ;
        RECT 6.656 1.98 6.688 4.488 ;
  LAYER M1 ;
        RECT 6.592 1.98 6.624 4.488 ;
  LAYER M1 ;
        RECT 6.528 1.98 6.56 4.488 ;
  LAYER M1 ;
        RECT 6.464 1.98 6.496 4.488 ;
  LAYER M1 ;
        RECT 6.4 1.98 6.432 4.488 ;
  LAYER M2 ;
        RECT 6.284 4.372 8.756 4.404 ;
  LAYER M2 ;
        RECT 6.284 4.308 8.756 4.34 ;
  LAYER M2 ;
        RECT 6.284 4.244 8.756 4.276 ;
  LAYER M2 ;
        RECT 6.284 4.18 8.756 4.212 ;
  LAYER M2 ;
        RECT 6.284 4.116 8.756 4.148 ;
  LAYER M2 ;
        RECT 6.284 4.052 8.756 4.084 ;
  LAYER M2 ;
        RECT 6.284 3.988 8.756 4.02 ;
  LAYER M2 ;
        RECT 6.284 3.924 8.756 3.956 ;
  LAYER M2 ;
        RECT 6.284 3.86 8.756 3.892 ;
  LAYER M2 ;
        RECT 6.284 3.796 8.756 3.828 ;
  LAYER M2 ;
        RECT 6.284 3.732 8.756 3.764 ;
  LAYER M2 ;
        RECT 6.284 3.668 8.756 3.7 ;
  LAYER M2 ;
        RECT 6.284 3.604 8.756 3.636 ;
  LAYER M2 ;
        RECT 6.284 3.54 8.756 3.572 ;
  LAYER M2 ;
        RECT 6.284 3.476 8.756 3.508 ;
  LAYER M2 ;
        RECT 6.284 3.412 8.756 3.444 ;
  LAYER M2 ;
        RECT 6.284 3.348 8.756 3.38 ;
  LAYER M2 ;
        RECT 6.284 3.284 8.756 3.316 ;
  LAYER M2 ;
        RECT 6.284 3.22 8.756 3.252 ;
  LAYER M2 ;
        RECT 6.284 3.156 8.756 3.188 ;
  LAYER M2 ;
        RECT 6.284 3.092 8.756 3.124 ;
  LAYER M2 ;
        RECT 6.284 3.028 8.756 3.06 ;
  LAYER M2 ;
        RECT 6.284 2.964 8.756 2.996 ;
  LAYER M2 ;
        RECT 6.284 2.9 8.756 2.932 ;
  LAYER M2 ;
        RECT 6.284 2.836 8.756 2.868 ;
  LAYER M2 ;
        RECT 6.284 2.772 8.756 2.804 ;
  LAYER M2 ;
        RECT 6.284 2.708 8.756 2.74 ;
  LAYER M2 ;
        RECT 6.284 2.644 8.756 2.676 ;
  LAYER M2 ;
        RECT 6.284 2.58 8.756 2.612 ;
  LAYER M2 ;
        RECT 6.284 2.516 8.756 2.548 ;
  LAYER M2 ;
        RECT 6.284 2.452 8.756 2.484 ;
  LAYER M2 ;
        RECT 6.284 2.388 8.756 2.42 ;
  LAYER M2 ;
        RECT 6.284 2.324 8.756 2.356 ;
  LAYER M2 ;
        RECT 6.284 2.26 8.756 2.292 ;
  LAYER M2 ;
        RECT 6.284 2.196 8.756 2.228 ;
  LAYER M2 ;
        RECT 6.284 2.132 8.756 2.164 ;
  LAYER M3 ;
        RECT 8.704 1.98 8.736 4.488 ;
  LAYER M3 ;
        RECT 8.64 1.98 8.672 4.488 ;
  LAYER M3 ;
        RECT 8.576 1.98 8.608 4.488 ;
  LAYER M3 ;
        RECT 8.512 1.98 8.544 4.488 ;
  LAYER M3 ;
        RECT 8.448 1.98 8.48 4.488 ;
  LAYER M3 ;
        RECT 8.384 1.98 8.416 4.488 ;
  LAYER M3 ;
        RECT 8.32 1.98 8.352 4.488 ;
  LAYER M3 ;
        RECT 8.256 1.98 8.288 4.488 ;
  LAYER M3 ;
        RECT 8.192 1.98 8.224 4.488 ;
  LAYER M3 ;
        RECT 8.128 1.98 8.16 4.488 ;
  LAYER M3 ;
        RECT 8.064 1.98 8.096 4.488 ;
  LAYER M3 ;
        RECT 8 1.98 8.032 4.488 ;
  LAYER M3 ;
        RECT 7.936 1.98 7.968 4.488 ;
  LAYER M3 ;
        RECT 7.872 1.98 7.904 4.488 ;
  LAYER M3 ;
        RECT 7.808 1.98 7.84 4.488 ;
  LAYER M3 ;
        RECT 7.744 1.98 7.776 4.488 ;
  LAYER M3 ;
        RECT 7.68 1.98 7.712 4.488 ;
  LAYER M3 ;
        RECT 7.616 1.98 7.648 4.488 ;
  LAYER M3 ;
        RECT 7.552 1.98 7.584 4.488 ;
  LAYER M3 ;
        RECT 7.488 1.98 7.52 4.488 ;
  LAYER M3 ;
        RECT 7.424 1.98 7.456 4.488 ;
  LAYER M3 ;
        RECT 7.36 1.98 7.392 4.488 ;
  LAYER M3 ;
        RECT 7.296 1.98 7.328 4.488 ;
  LAYER M3 ;
        RECT 7.232 1.98 7.264 4.488 ;
  LAYER M3 ;
        RECT 7.168 1.98 7.2 4.488 ;
  LAYER M3 ;
        RECT 7.104 1.98 7.136 4.488 ;
  LAYER M3 ;
        RECT 7.04 1.98 7.072 4.488 ;
  LAYER M3 ;
        RECT 6.976 1.98 7.008 4.488 ;
  LAYER M3 ;
        RECT 6.912 1.98 6.944 4.488 ;
  LAYER M3 ;
        RECT 6.848 1.98 6.88 4.488 ;
  LAYER M3 ;
        RECT 6.784 1.98 6.816 4.488 ;
  LAYER M3 ;
        RECT 6.72 1.98 6.752 4.488 ;
  LAYER M3 ;
        RECT 6.656 1.98 6.688 4.488 ;
  LAYER M3 ;
        RECT 6.592 1.98 6.624 4.488 ;
  LAYER M3 ;
        RECT 6.528 1.98 6.56 4.488 ;
  LAYER M3 ;
        RECT 6.464 1.98 6.496 4.488 ;
  LAYER M3 ;
        RECT 6.4 1.98 6.432 4.488 ;
  LAYER M3 ;
        RECT 6.304 1.98 6.336 4.488 ;
  LAYER M1 ;
        RECT 8.719 2.016 8.721 4.452 ;
  LAYER M1 ;
        RECT 8.639 2.016 8.641 4.452 ;
  LAYER M1 ;
        RECT 8.559 2.016 8.561 4.452 ;
  LAYER M1 ;
        RECT 8.479 2.016 8.481 4.452 ;
  LAYER M1 ;
        RECT 8.399 2.016 8.401 4.452 ;
  LAYER M1 ;
        RECT 8.319 2.016 8.321 4.452 ;
  LAYER M1 ;
        RECT 8.239 2.016 8.241 4.452 ;
  LAYER M1 ;
        RECT 8.159 2.016 8.161 4.452 ;
  LAYER M1 ;
        RECT 8.079 2.016 8.081 4.452 ;
  LAYER M1 ;
        RECT 7.999 2.016 8.001 4.452 ;
  LAYER M1 ;
        RECT 7.919 2.016 7.921 4.452 ;
  LAYER M1 ;
        RECT 7.839 2.016 7.841 4.452 ;
  LAYER M1 ;
        RECT 7.759 2.016 7.761 4.452 ;
  LAYER M1 ;
        RECT 7.679 2.016 7.681 4.452 ;
  LAYER M1 ;
        RECT 7.599 2.016 7.601 4.452 ;
  LAYER M1 ;
        RECT 7.519 2.016 7.521 4.452 ;
  LAYER M1 ;
        RECT 7.439 2.016 7.441 4.452 ;
  LAYER M1 ;
        RECT 7.359 2.016 7.361 4.452 ;
  LAYER M1 ;
        RECT 7.279 2.016 7.281 4.452 ;
  LAYER M1 ;
        RECT 7.199 2.016 7.201 4.452 ;
  LAYER M1 ;
        RECT 7.119 2.016 7.121 4.452 ;
  LAYER M1 ;
        RECT 7.039 2.016 7.041 4.452 ;
  LAYER M1 ;
        RECT 6.959 2.016 6.961 4.452 ;
  LAYER M1 ;
        RECT 6.879 2.016 6.881 4.452 ;
  LAYER M1 ;
        RECT 6.799 2.016 6.801 4.452 ;
  LAYER M1 ;
        RECT 6.719 2.016 6.721 4.452 ;
  LAYER M1 ;
        RECT 6.639 2.016 6.641 4.452 ;
  LAYER M1 ;
        RECT 6.559 2.016 6.561 4.452 ;
  LAYER M1 ;
        RECT 6.479 2.016 6.481 4.452 ;
  LAYER M1 ;
        RECT 6.399 2.016 6.401 4.452 ;
  LAYER M2 ;
        RECT 6.32 4.451 8.72 4.453 ;
  LAYER M2 ;
        RECT 6.32 4.367 8.72 4.369 ;
  LAYER M2 ;
        RECT 6.32 4.283 8.72 4.285 ;
  LAYER M2 ;
        RECT 6.32 4.199 8.72 4.201 ;
  LAYER M2 ;
        RECT 6.32 4.115 8.72 4.117 ;
  LAYER M2 ;
        RECT 6.32 4.031 8.72 4.033 ;
  LAYER M2 ;
        RECT 6.32 3.947 8.72 3.949 ;
  LAYER M2 ;
        RECT 6.32 3.863 8.72 3.865 ;
  LAYER M2 ;
        RECT 6.32 3.779 8.72 3.781 ;
  LAYER M2 ;
        RECT 6.32 3.695 8.72 3.697 ;
  LAYER M2 ;
        RECT 6.32 3.611 8.72 3.613 ;
  LAYER M2 ;
        RECT 6.32 3.527 8.72 3.529 ;
  LAYER M2 ;
        RECT 6.32 3.4435 8.72 3.4455 ;
  LAYER M2 ;
        RECT 6.32 3.359 8.72 3.361 ;
  LAYER M2 ;
        RECT 6.32 3.275 8.72 3.277 ;
  LAYER M2 ;
        RECT 6.32 3.191 8.72 3.193 ;
  LAYER M2 ;
        RECT 6.32 3.107 8.72 3.109 ;
  LAYER M2 ;
        RECT 6.32 3.023 8.72 3.025 ;
  LAYER M2 ;
        RECT 6.32 2.939 8.72 2.941 ;
  LAYER M2 ;
        RECT 6.32 2.855 8.72 2.857 ;
  LAYER M2 ;
        RECT 6.32 2.771 8.72 2.773 ;
  LAYER M2 ;
        RECT 6.32 2.687 8.72 2.689 ;
  LAYER M2 ;
        RECT 6.32 2.603 8.72 2.605 ;
  LAYER M2 ;
        RECT 6.32 2.519 8.72 2.521 ;
  LAYER M2 ;
        RECT 6.32 2.435 8.72 2.437 ;
  LAYER M2 ;
        RECT 6.32 2.351 8.72 2.353 ;
  LAYER M2 ;
        RECT 6.32 2.267 8.72 2.269 ;
  LAYER M2 ;
        RECT 6.32 2.183 8.72 2.185 ;
  LAYER M2 ;
        RECT 6.32 2.099 8.72 2.101 ;
  LAYER M1 ;
        RECT 5.824 13.74 5.856 16.248 ;
  LAYER M1 ;
        RECT 5.76 13.74 5.792 16.248 ;
  LAYER M1 ;
        RECT 5.696 13.74 5.728 16.248 ;
  LAYER M1 ;
        RECT 5.632 13.74 5.664 16.248 ;
  LAYER M1 ;
        RECT 5.568 13.74 5.6 16.248 ;
  LAYER M1 ;
        RECT 5.504 13.74 5.536 16.248 ;
  LAYER M1 ;
        RECT 5.44 13.74 5.472 16.248 ;
  LAYER M1 ;
        RECT 5.376 13.74 5.408 16.248 ;
  LAYER M1 ;
        RECT 5.312 13.74 5.344 16.248 ;
  LAYER M1 ;
        RECT 5.248 13.74 5.28 16.248 ;
  LAYER M1 ;
        RECT 5.184 13.74 5.216 16.248 ;
  LAYER M1 ;
        RECT 5.12 13.74 5.152 16.248 ;
  LAYER M1 ;
        RECT 5.056 13.74 5.088 16.248 ;
  LAYER M1 ;
        RECT 4.992 13.74 5.024 16.248 ;
  LAYER M1 ;
        RECT 4.928 13.74 4.96 16.248 ;
  LAYER M1 ;
        RECT 4.864 13.74 4.896 16.248 ;
  LAYER M1 ;
        RECT 4.8 13.74 4.832 16.248 ;
  LAYER M1 ;
        RECT 4.736 13.74 4.768 16.248 ;
  LAYER M1 ;
        RECT 4.672 13.74 4.704 16.248 ;
  LAYER M1 ;
        RECT 4.608 13.74 4.64 16.248 ;
  LAYER M1 ;
        RECT 4.544 13.74 4.576 16.248 ;
  LAYER M1 ;
        RECT 4.48 13.74 4.512 16.248 ;
  LAYER M1 ;
        RECT 4.416 13.74 4.448 16.248 ;
  LAYER M1 ;
        RECT 4.352 13.74 4.384 16.248 ;
  LAYER M1 ;
        RECT 4.288 13.74 4.32 16.248 ;
  LAYER M1 ;
        RECT 4.224 13.74 4.256 16.248 ;
  LAYER M1 ;
        RECT 4.16 13.74 4.192 16.248 ;
  LAYER M1 ;
        RECT 4.096 13.74 4.128 16.248 ;
  LAYER M1 ;
        RECT 4.032 13.74 4.064 16.248 ;
  LAYER M1 ;
        RECT 3.968 13.74 4 16.248 ;
  LAYER M1 ;
        RECT 3.904 13.74 3.936 16.248 ;
  LAYER M1 ;
        RECT 3.84 13.74 3.872 16.248 ;
  LAYER M1 ;
        RECT 3.776 13.74 3.808 16.248 ;
  LAYER M1 ;
        RECT 3.712 13.74 3.744 16.248 ;
  LAYER M1 ;
        RECT 3.648 13.74 3.68 16.248 ;
  LAYER M1 ;
        RECT 3.584 13.74 3.616 16.248 ;
  LAYER M1 ;
        RECT 3.52 13.74 3.552 16.248 ;
  LAYER M2 ;
        RECT 3.404 16.132 5.876 16.164 ;
  LAYER M2 ;
        RECT 3.404 16.068 5.876 16.1 ;
  LAYER M2 ;
        RECT 3.404 16.004 5.876 16.036 ;
  LAYER M2 ;
        RECT 3.404 15.94 5.876 15.972 ;
  LAYER M2 ;
        RECT 3.404 15.876 5.876 15.908 ;
  LAYER M2 ;
        RECT 3.404 15.812 5.876 15.844 ;
  LAYER M2 ;
        RECT 3.404 15.748 5.876 15.78 ;
  LAYER M2 ;
        RECT 3.404 15.684 5.876 15.716 ;
  LAYER M2 ;
        RECT 3.404 15.62 5.876 15.652 ;
  LAYER M2 ;
        RECT 3.404 15.556 5.876 15.588 ;
  LAYER M2 ;
        RECT 3.404 15.492 5.876 15.524 ;
  LAYER M2 ;
        RECT 3.404 15.428 5.876 15.46 ;
  LAYER M2 ;
        RECT 3.404 15.364 5.876 15.396 ;
  LAYER M2 ;
        RECT 3.404 15.3 5.876 15.332 ;
  LAYER M2 ;
        RECT 3.404 15.236 5.876 15.268 ;
  LAYER M2 ;
        RECT 3.404 15.172 5.876 15.204 ;
  LAYER M2 ;
        RECT 3.404 15.108 5.876 15.14 ;
  LAYER M2 ;
        RECT 3.404 15.044 5.876 15.076 ;
  LAYER M2 ;
        RECT 3.404 14.98 5.876 15.012 ;
  LAYER M2 ;
        RECT 3.404 14.916 5.876 14.948 ;
  LAYER M2 ;
        RECT 3.404 14.852 5.876 14.884 ;
  LAYER M2 ;
        RECT 3.404 14.788 5.876 14.82 ;
  LAYER M2 ;
        RECT 3.404 14.724 5.876 14.756 ;
  LAYER M2 ;
        RECT 3.404 14.66 5.876 14.692 ;
  LAYER M2 ;
        RECT 3.404 14.596 5.876 14.628 ;
  LAYER M2 ;
        RECT 3.404 14.532 5.876 14.564 ;
  LAYER M2 ;
        RECT 3.404 14.468 5.876 14.5 ;
  LAYER M2 ;
        RECT 3.404 14.404 5.876 14.436 ;
  LAYER M2 ;
        RECT 3.404 14.34 5.876 14.372 ;
  LAYER M2 ;
        RECT 3.404 14.276 5.876 14.308 ;
  LAYER M2 ;
        RECT 3.404 14.212 5.876 14.244 ;
  LAYER M2 ;
        RECT 3.404 14.148 5.876 14.18 ;
  LAYER M2 ;
        RECT 3.404 14.084 5.876 14.116 ;
  LAYER M2 ;
        RECT 3.404 14.02 5.876 14.052 ;
  LAYER M2 ;
        RECT 3.404 13.956 5.876 13.988 ;
  LAYER M2 ;
        RECT 3.404 13.892 5.876 13.924 ;
  LAYER M3 ;
        RECT 5.824 13.74 5.856 16.248 ;
  LAYER M3 ;
        RECT 5.76 13.74 5.792 16.248 ;
  LAYER M3 ;
        RECT 5.696 13.74 5.728 16.248 ;
  LAYER M3 ;
        RECT 5.632 13.74 5.664 16.248 ;
  LAYER M3 ;
        RECT 5.568 13.74 5.6 16.248 ;
  LAYER M3 ;
        RECT 5.504 13.74 5.536 16.248 ;
  LAYER M3 ;
        RECT 5.44 13.74 5.472 16.248 ;
  LAYER M3 ;
        RECT 5.376 13.74 5.408 16.248 ;
  LAYER M3 ;
        RECT 5.312 13.74 5.344 16.248 ;
  LAYER M3 ;
        RECT 5.248 13.74 5.28 16.248 ;
  LAYER M3 ;
        RECT 5.184 13.74 5.216 16.248 ;
  LAYER M3 ;
        RECT 5.12 13.74 5.152 16.248 ;
  LAYER M3 ;
        RECT 5.056 13.74 5.088 16.248 ;
  LAYER M3 ;
        RECT 4.992 13.74 5.024 16.248 ;
  LAYER M3 ;
        RECT 4.928 13.74 4.96 16.248 ;
  LAYER M3 ;
        RECT 4.864 13.74 4.896 16.248 ;
  LAYER M3 ;
        RECT 4.8 13.74 4.832 16.248 ;
  LAYER M3 ;
        RECT 4.736 13.74 4.768 16.248 ;
  LAYER M3 ;
        RECT 4.672 13.74 4.704 16.248 ;
  LAYER M3 ;
        RECT 4.608 13.74 4.64 16.248 ;
  LAYER M3 ;
        RECT 4.544 13.74 4.576 16.248 ;
  LAYER M3 ;
        RECT 4.48 13.74 4.512 16.248 ;
  LAYER M3 ;
        RECT 4.416 13.74 4.448 16.248 ;
  LAYER M3 ;
        RECT 4.352 13.74 4.384 16.248 ;
  LAYER M3 ;
        RECT 4.288 13.74 4.32 16.248 ;
  LAYER M3 ;
        RECT 4.224 13.74 4.256 16.248 ;
  LAYER M3 ;
        RECT 4.16 13.74 4.192 16.248 ;
  LAYER M3 ;
        RECT 4.096 13.74 4.128 16.248 ;
  LAYER M3 ;
        RECT 4.032 13.74 4.064 16.248 ;
  LAYER M3 ;
        RECT 3.968 13.74 4 16.248 ;
  LAYER M3 ;
        RECT 3.904 13.74 3.936 16.248 ;
  LAYER M3 ;
        RECT 3.84 13.74 3.872 16.248 ;
  LAYER M3 ;
        RECT 3.776 13.74 3.808 16.248 ;
  LAYER M3 ;
        RECT 3.712 13.74 3.744 16.248 ;
  LAYER M3 ;
        RECT 3.648 13.74 3.68 16.248 ;
  LAYER M3 ;
        RECT 3.584 13.74 3.616 16.248 ;
  LAYER M3 ;
        RECT 3.52 13.74 3.552 16.248 ;
  LAYER M3 ;
        RECT 3.424 13.74 3.456 16.248 ;
  LAYER M1 ;
        RECT 5.839 13.776 5.841 16.212 ;
  LAYER M1 ;
        RECT 5.759 13.776 5.761 16.212 ;
  LAYER M1 ;
        RECT 5.679 13.776 5.681 16.212 ;
  LAYER M1 ;
        RECT 5.599 13.776 5.601 16.212 ;
  LAYER M1 ;
        RECT 5.519 13.776 5.521 16.212 ;
  LAYER M1 ;
        RECT 5.439 13.776 5.441 16.212 ;
  LAYER M1 ;
        RECT 5.359 13.776 5.361 16.212 ;
  LAYER M1 ;
        RECT 5.279 13.776 5.281 16.212 ;
  LAYER M1 ;
        RECT 5.199 13.776 5.201 16.212 ;
  LAYER M1 ;
        RECT 5.119 13.776 5.121 16.212 ;
  LAYER M1 ;
        RECT 5.039 13.776 5.041 16.212 ;
  LAYER M1 ;
        RECT 4.959 13.776 4.961 16.212 ;
  LAYER M1 ;
        RECT 4.879 13.776 4.881 16.212 ;
  LAYER M1 ;
        RECT 4.799 13.776 4.801 16.212 ;
  LAYER M1 ;
        RECT 4.719 13.776 4.721 16.212 ;
  LAYER M1 ;
        RECT 4.639 13.776 4.641 16.212 ;
  LAYER M1 ;
        RECT 4.559 13.776 4.561 16.212 ;
  LAYER M1 ;
        RECT 4.479 13.776 4.481 16.212 ;
  LAYER M1 ;
        RECT 4.399 13.776 4.401 16.212 ;
  LAYER M1 ;
        RECT 4.319 13.776 4.321 16.212 ;
  LAYER M1 ;
        RECT 4.239 13.776 4.241 16.212 ;
  LAYER M1 ;
        RECT 4.159 13.776 4.161 16.212 ;
  LAYER M1 ;
        RECT 4.079 13.776 4.081 16.212 ;
  LAYER M1 ;
        RECT 3.999 13.776 4.001 16.212 ;
  LAYER M1 ;
        RECT 3.919 13.776 3.921 16.212 ;
  LAYER M1 ;
        RECT 3.839 13.776 3.841 16.212 ;
  LAYER M1 ;
        RECT 3.759 13.776 3.761 16.212 ;
  LAYER M1 ;
        RECT 3.679 13.776 3.681 16.212 ;
  LAYER M1 ;
        RECT 3.599 13.776 3.601 16.212 ;
  LAYER M1 ;
        RECT 3.519 13.776 3.521 16.212 ;
  LAYER M2 ;
        RECT 3.44 16.211 5.84 16.213 ;
  LAYER M2 ;
        RECT 3.44 16.127 5.84 16.129 ;
  LAYER M2 ;
        RECT 3.44 16.043 5.84 16.045 ;
  LAYER M2 ;
        RECT 3.44 15.959 5.84 15.961 ;
  LAYER M2 ;
        RECT 3.44 15.875 5.84 15.877 ;
  LAYER M2 ;
        RECT 3.44 15.791 5.84 15.793 ;
  LAYER M2 ;
        RECT 3.44 15.707 5.84 15.709 ;
  LAYER M2 ;
        RECT 3.44 15.623 5.84 15.625 ;
  LAYER M2 ;
        RECT 3.44 15.539 5.84 15.541 ;
  LAYER M2 ;
        RECT 3.44 15.455 5.84 15.457 ;
  LAYER M2 ;
        RECT 3.44 15.371 5.84 15.373 ;
  LAYER M2 ;
        RECT 3.44 15.287 5.84 15.289 ;
  LAYER M2 ;
        RECT 3.44 15.2035 5.84 15.2055 ;
  LAYER M2 ;
        RECT 3.44 15.119 5.84 15.121 ;
  LAYER M2 ;
        RECT 3.44 15.035 5.84 15.037 ;
  LAYER M2 ;
        RECT 3.44 14.951 5.84 14.953 ;
  LAYER M2 ;
        RECT 3.44 14.867 5.84 14.869 ;
  LAYER M2 ;
        RECT 3.44 14.783 5.84 14.785 ;
  LAYER M2 ;
        RECT 3.44 14.699 5.84 14.701 ;
  LAYER M2 ;
        RECT 3.44 14.615 5.84 14.617 ;
  LAYER M2 ;
        RECT 3.44 14.531 5.84 14.533 ;
  LAYER M2 ;
        RECT 3.44 14.447 5.84 14.449 ;
  LAYER M2 ;
        RECT 3.44 14.363 5.84 14.365 ;
  LAYER M2 ;
        RECT 3.44 14.279 5.84 14.281 ;
  LAYER M2 ;
        RECT 3.44 14.195 5.84 14.197 ;
  LAYER M2 ;
        RECT 3.44 14.111 5.84 14.113 ;
  LAYER M2 ;
        RECT 3.44 14.027 5.84 14.029 ;
  LAYER M2 ;
        RECT 3.44 13.943 5.84 13.945 ;
  LAYER M2 ;
        RECT 3.44 13.859 5.84 13.861 ;
  LAYER M1 ;
        RECT 5.824 10.8 5.856 13.308 ;
  LAYER M1 ;
        RECT 5.76 10.8 5.792 13.308 ;
  LAYER M1 ;
        RECT 5.696 10.8 5.728 13.308 ;
  LAYER M1 ;
        RECT 5.632 10.8 5.664 13.308 ;
  LAYER M1 ;
        RECT 5.568 10.8 5.6 13.308 ;
  LAYER M1 ;
        RECT 5.504 10.8 5.536 13.308 ;
  LAYER M1 ;
        RECT 5.44 10.8 5.472 13.308 ;
  LAYER M1 ;
        RECT 5.376 10.8 5.408 13.308 ;
  LAYER M1 ;
        RECT 5.312 10.8 5.344 13.308 ;
  LAYER M1 ;
        RECT 5.248 10.8 5.28 13.308 ;
  LAYER M1 ;
        RECT 5.184 10.8 5.216 13.308 ;
  LAYER M1 ;
        RECT 5.12 10.8 5.152 13.308 ;
  LAYER M1 ;
        RECT 5.056 10.8 5.088 13.308 ;
  LAYER M1 ;
        RECT 4.992 10.8 5.024 13.308 ;
  LAYER M1 ;
        RECT 4.928 10.8 4.96 13.308 ;
  LAYER M1 ;
        RECT 4.864 10.8 4.896 13.308 ;
  LAYER M1 ;
        RECT 4.8 10.8 4.832 13.308 ;
  LAYER M1 ;
        RECT 4.736 10.8 4.768 13.308 ;
  LAYER M1 ;
        RECT 4.672 10.8 4.704 13.308 ;
  LAYER M1 ;
        RECT 4.608 10.8 4.64 13.308 ;
  LAYER M1 ;
        RECT 4.544 10.8 4.576 13.308 ;
  LAYER M1 ;
        RECT 4.48 10.8 4.512 13.308 ;
  LAYER M1 ;
        RECT 4.416 10.8 4.448 13.308 ;
  LAYER M1 ;
        RECT 4.352 10.8 4.384 13.308 ;
  LAYER M1 ;
        RECT 4.288 10.8 4.32 13.308 ;
  LAYER M1 ;
        RECT 4.224 10.8 4.256 13.308 ;
  LAYER M1 ;
        RECT 4.16 10.8 4.192 13.308 ;
  LAYER M1 ;
        RECT 4.096 10.8 4.128 13.308 ;
  LAYER M1 ;
        RECT 4.032 10.8 4.064 13.308 ;
  LAYER M1 ;
        RECT 3.968 10.8 4 13.308 ;
  LAYER M1 ;
        RECT 3.904 10.8 3.936 13.308 ;
  LAYER M1 ;
        RECT 3.84 10.8 3.872 13.308 ;
  LAYER M1 ;
        RECT 3.776 10.8 3.808 13.308 ;
  LAYER M1 ;
        RECT 3.712 10.8 3.744 13.308 ;
  LAYER M1 ;
        RECT 3.648 10.8 3.68 13.308 ;
  LAYER M1 ;
        RECT 3.584 10.8 3.616 13.308 ;
  LAYER M1 ;
        RECT 3.52 10.8 3.552 13.308 ;
  LAYER M2 ;
        RECT 3.404 13.192 5.876 13.224 ;
  LAYER M2 ;
        RECT 3.404 13.128 5.876 13.16 ;
  LAYER M2 ;
        RECT 3.404 13.064 5.876 13.096 ;
  LAYER M2 ;
        RECT 3.404 13 5.876 13.032 ;
  LAYER M2 ;
        RECT 3.404 12.936 5.876 12.968 ;
  LAYER M2 ;
        RECT 3.404 12.872 5.876 12.904 ;
  LAYER M2 ;
        RECT 3.404 12.808 5.876 12.84 ;
  LAYER M2 ;
        RECT 3.404 12.744 5.876 12.776 ;
  LAYER M2 ;
        RECT 3.404 12.68 5.876 12.712 ;
  LAYER M2 ;
        RECT 3.404 12.616 5.876 12.648 ;
  LAYER M2 ;
        RECT 3.404 12.552 5.876 12.584 ;
  LAYER M2 ;
        RECT 3.404 12.488 5.876 12.52 ;
  LAYER M2 ;
        RECT 3.404 12.424 5.876 12.456 ;
  LAYER M2 ;
        RECT 3.404 12.36 5.876 12.392 ;
  LAYER M2 ;
        RECT 3.404 12.296 5.876 12.328 ;
  LAYER M2 ;
        RECT 3.404 12.232 5.876 12.264 ;
  LAYER M2 ;
        RECT 3.404 12.168 5.876 12.2 ;
  LAYER M2 ;
        RECT 3.404 12.104 5.876 12.136 ;
  LAYER M2 ;
        RECT 3.404 12.04 5.876 12.072 ;
  LAYER M2 ;
        RECT 3.404 11.976 5.876 12.008 ;
  LAYER M2 ;
        RECT 3.404 11.912 5.876 11.944 ;
  LAYER M2 ;
        RECT 3.404 11.848 5.876 11.88 ;
  LAYER M2 ;
        RECT 3.404 11.784 5.876 11.816 ;
  LAYER M2 ;
        RECT 3.404 11.72 5.876 11.752 ;
  LAYER M2 ;
        RECT 3.404 11.656 5.876 11.688 ;
  LAYER M2 ;
        RECT 3.404 11.592 5.876 11.624 ;
  LAYER M2 ;
        RECT 3.404 11.528 5.876 11.56 ;
  LAYER M2 ;
        RECT 3.404 11.464 5.876 11.496 ;
  LAYER M2 ;
        RECT 3.404 11.4 5.876 11.432 ;
  LAYER M2 ;
        RECT 3.404 11.336 5.876 11.368 ;
  LAYER M2 ;
        RECT 3.404 11.272 5.876 11.304 ;
  LAYER M2 ;
        RECT 3.404 11.208 5.876 11.24 ;
  LAYER M2 ;
        RECT 3.404 11.144 5.876 11.176 ;
  LAYER M2 ;
        RECT 3.404 11.08 5.876 11.112 ;
  LAYER M2 ;
        RECT 3.404 11.016 5.876 11.048 ;
  LAYER M2 ;
        RECT 3.404 10.952 5.876 10.984 ;
  LAYER M3 ;
        RECT 5.824 10.8 5.856 13.308 ;
  LAYER M3 ;
        RECT 5.76 10.8 5.792 13.308 ;
  LAYER M3 ;
        RECT 5.696 10.8 5.728 13.308 ;
  LAYER M3 ;
        RECT 5.632 10.8 5.664 13.308 ;
  LAYER M3 ;
        RECT 5.568 10.8 5.6 13.308 ;
  LAYER M3 ;
        RECT 5.504 10.8 5.536 13.308 ;
  LAYER M3 ;
        RECT 5.44 10.8 5.472 13.308 ;
  LAYER M3 ;
        RECT 5.376 10.8 5.408 13.308 ;
  LAYER M3 ;
        RECT 5.312 10.8 5.344 13.308 ;
  LAYER M3 ;
        RECT 5.248 10.8 5.28 13.308 ;
  LAYER M3 ;
        RECT 5.184 10.8 5.216 13.308 ;
  LAYER M3 ;
        RECT 5.12 10.8 5.152 13.308 ;
  LAYER M3 ;
        RECT 5.056 10.8 5.088 13.308 ;
  LAYER M3 ;
        RECT 4.992 10.8 5.024 13.308 ;
  LAYER M3 ;
        RECT 4.928 10.8 4.96 13.308 ;
  LAYER M3 ;
        RECT 4.864 10.8 4.896 13.308 ;
  LAYER M3 ;
        RECT 4.8 10.8 4.832 13.308 ;
  LAYER M3 ;
        RECT 4.736 10.8 4.768 13.308 ;
  LAYER M3 ;
        RECT 4.672 10.8 4.704 13.308 ;
  LAYER M3 ;
        RECT 4.608 10.8 4.64 13.308 ;
  LAYER M3 ;
        RECT 4.544 10.8 4.576 13.308 ;
  LAYER M3 ;
        RECT 4.48 10.8 4.512 13.308 ;
  LAYER M3 ;
        RECT 4.416 10.8 4.448 13.308 ;
  LAYER M3 ;
        RECT 4.352 10.8 4.384 13.308 ;
  LAYER M3 ;
        RECT 4.288 10.8 4.32 13.308 ;
  LAYER M3 ;
        RECT 4.224 10.8 4.256 13.308 ;
  LAYER M3 ;
        RECT 4.16 10.8 4.192 13.308 ;
  LAYER M3 ;
        RECT 4.096 10.8 4.128 13.308 ;
  LAYER M3 ;
        RECT 4.032 10.8 4.064 13.308 ;
  LAYER M3 ;
        RECT 3.968 10.8 4 13.308 ;
  LAYER M3 ;
        RECT 3.904 10.8 3.936 13.308 ;
  LAYER M3 ;
        RECT 3.84 10.8 3.872 13.308 ;
  LAYER M3 ;
        RECT 3.776 10.8 3.808 13.308 ;
  LAYER M3 ;
        RECT 3.712 10.8 3.744 13.308 ;
  LAYER M3 ;
        RECT 3.648 10.8 3.68 13.308 ;
  LAYER M3 ;
        RECT 3.584 10.8 3.616 13.308 ;
  LAYER M3 ;
        RECT 3.52 10.8 3.552 13.308 ;
  LAYER M3 ;
        RECT 3.424 10.8 3.456 13.308 ;
  LAYER M1 ;
        RECT 5.839 10.836 5.841 13.272 ;
  LAYER M1 ;
        RECT 5.759 10.836 5.761 13.272 ;
  LAYER M1 ;
        RECT 5.679 10.836 5.681 13.272 ;
  LAYER M1 ;
        RECT 5.599 10.836 5.601 13.272 ;
  LAYER M1 ;
        RECT 5.519 10.836 5.521 13.272 ;
  LAYER M1 ;
        RECT 5.439 10.836 5.441 13.272 ;
  LAYER M1 ;
        RECT 5.359 10.836 5.361 13.272 ;
  LAYER M1 ;
        RECT 5.279 10.836 5.281 13.272 ;
  LAYER M1 ;
        RECT 5.199 10.836 5.201 13.272 ;
  LAYER M1 ;
        RECT 5.119 10.836 5.121 13.272 ;
  LAYER M1 ;
        RECT 5.039 10.836 5.041 13.272 ;
  LAYER M1 ;
        RECT 4.959 10.836 4.961 13.272 ;
  LAYER M1 ;
        RECT 4.879 10.836 4.881 13.272 ;
  LAYER M1 ;
        RECT 4.799 10.836 4.801 13.272 ;
  LAYER M1 ;
        RECT 4.719 10.836 4.721 13.272 ;
  LAYER M1 ;
        RECT 4.639 10.836 4.641 13.272 ;
  LAYER M1 ;
        RECT 4.559 10.836 4.561 13.272 ;
  LAYER M1 ;
        RECT 4.479 10.836 4.481 13.272 ;
  LAYER M1 ;
        RECT 4.399 10.836 4.401 13.272 ;
  LAYER M1 ;
        RECT 4.319 10.836 4.321 13.272 ;
  LAYER M1 ;
        RECT 4.239 10.836 4.241 13.272 ;
  LAYER M1 ;
        RECT 4.159 10.836 4.161 13.272 ;
  LAYER M1 ;
        RECT 4.079 10.836 4.081 13.272 ;
  LAYER M1 ;
        RECT 3.999 10.836 4.001 13.272 ;
  LAYER M1 ;
        RECT 3.919 10.836 3.921 13.272 ;
  LAYER M1 ;
        RECT 3.839 10.836 3.841 13.272 ;
  LAYER M1 ;
        RECT 3.759 10.836 3.761 13.272 ;
  LAYER M1 ;
        RECT 3.679 10.836 3.681 13.272 ;
  LAYER M1 ;
        RECT 3.599 10.836 3.601 13.272 ;
  LAYER M1 ;
        RECT 3.519 10.836 3.521 13.272 ;
  LAYER M2 ;
        RECT 3.44 13.271 5.84 13.273 ;
  LAYER M2 ;
        RECT 3.44 13.187 5.84 13.189 ;
  LAYER M2 ;
        RECT 3.44 13.103 5.84 13.105 ;
  LAYER M2 ;
        RECT 3.44 13.019 5.84 13.021 ;
  LAYER M2 ;
        RECT 3.44 12.935 5.84 12.937 ;
  LAYER M2 ;
        RECT 3.44 12.851 5.84 12.853 ;
  LAYER M2 ;
        RECT 3.44 12.767 5.84 12.769 ;
  LAYER M2 ;
        RECT 3.44 12.683 5.84 12.685 ;
  LAYER M2 ;
        RECT 3.44 12.599 5.84 12.601 ;
  LAYER M2 ;
        RECT 3.44 12.515 5.84 12.517 ;
  LAYER M2 ;
        RECT 3.44 12.431 5.84 12.433 ;
  LAYER M2 ;
        RECT 3.44 12.347 5.84 12.349 ;
  LAYER M2 ;
        RECT 3.44 12.2635 5.84 12.2655 ;
  LAYER M2 ;
        RECT 3.44 12.179 5.84 12.181 ;
  LAYER M2 ;
        RECT 3.44 12.095 5.84 12.097 ;
  LAYER M2 ;
        RECT 3.44 12.011 5.84 12.013 ;
  LAYER M2 ;
        RECT 3.44 11.927 5.84 11.929 ;
  LAYER M2 ;
        RECT 3.44 11.843 5.84 11.845 ;
  LAYER M2 ;
        RECT 3.44 11.759 5.84 11.761 ;
  LAYER M2 ;
        RECT 3.44 11.675 5.84 11.677 ;
  LAYER M2 ;
        RECT 3.44 11.591 5.84 11.593 ;
  LAYER M2 ;
        RECT 3.44 11.507 5.84 11.509 ;
  LAYER M2 ;
        RECT 3.44 11.423 5.84 11.425 ;
  LAYER M2 ;
        RECT 3.44 11.339 5.84 11.341 ;
  LAYER M2 ;
        RECT 3.44 11.255 5.84 11.257 ;
  LAYER M2 ;
        RECT 3.44 11.171 5.84 11.173 ;
  LAYER M2 ;
        RECT 3.44 11.087 5.84 11.089 ;
  LAYER M2 ;
        RECT 3.44 11.003 5.84 11.005 ;
  LAYER M2 ;
        RECT 3.44 10.919 5.84 10.921 ;
  LAYER M1 ;
        RECT 5.824 7.86 5.856 10.368 ;
  LAYER M1 ;
        RECT 5.76 7.86 5.792 10.368 ;
  LAYER M1 ;
        RECT 5.696 7.86 5.728 10.368 ;
  LAYER M1 ;
        RECT 5.632 7.86 5.664 10.368 ;
  LAYER M1 ;
        RECT 5.568 7.86 5.6 10.368 ;
  LAYER M1 ;
        RECT 5.504 7.86 5.536 10.368 ;
  LAYER M1 ;
        RECT 5.44 7.86 5.472 10.368 ;
  LAYER M1 ;
        RECT 5.376 7.86 5.408 10.368 ;
  LAYER M1 ;
        RECT 5.312 7.86 5.344 10.368 ;
  LAYER M1 ;
        RECT 5.248 7.86 5.28 10.368 ;
  LAYER M1 ;
        RECT 5.184 7.86 5.216 10.368 ;
  LAYER M1 ;
        RECT 5.12 7.86 5.152 10.368 ;
  LAYER M1 ;
        RECT 5.056 7.86 5.088 10.368 ;
  LAYER M1 ;
        RECT 4.992 7.86 5.024 10.368 ;
  LAYER M1 ;
        RECT 4.928 7.86 4.96 10.368 ;
  LAYER M1 ;
        RECT 4.864 7.86 4.896 10.368 ;
  LAYER M1 ;
        RECT 4.8 7.86 4.832 10.368 ;
  LAYER M1 ;
        RECT 4.736 7.86 4.768 10.368 ;
  LAYER M1 ;
        RECT 4.672 7.86 4.704 10.368 ;
  LAYER M1 ;
        RECT 4.608 7.86 4.64 10.368 ;
  LAYER M1 ;
        RECT 4.544 7.86 4.576 10.368 ;
  LAYER M1 ;
        RECT 4.48 7.86 4.512 10.368 ;
  LAYER M1 ;
        RECT 4.416 7.86 4.448 10.368 ;
  LAYER M1 ;
        RECT 4.352 7.86 4.384 10.368 ;
  LAYER M1 ;
        RECT 4.288 7.86 4.32 10.368 ;
  LAYER M1 ;
        RECT 4.224 7.86 4.256 10.368 ;
  LAYER M1 ;
        RECT 4.16 7.86 4.192 10.368 ;
  LAYER M1 ;
        RECT 4.096 7.86 4.128 10.368 ;
  LAYER M1 ;
        RECT 4.032 7.86 4.064 10.368 ;
  LAYER M1 ;
        RECT 3.968 7.86 4 10.368 ;
  LAYER M1 ;
        RECT 3.904 7.86 3.936 10.368 ;
  LAYER M1 ;
        RECT 3.84 7.86 3.872 10.368 ;
  LAYER M1 ;
        RECT 3.776 7.86 3.808 10.368 ;
  LAYER M1 ;
        RECT 3.712 7.86 3.744 10.368 ;
  LAYER M1 ;
        RECT 3.648 7.86 3.68 10.368 ;
  LAYER M1 ;
        RECT 3.584 7.86 3.616 10.368 ;
  LAYER M1 ;
        RECT 3.52 7.86 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.404 10.252 5.876 10.284 ;
  LAYER M2 ;
        RECT 3.404 10.188 5.876 10.22 ;
  LAYER M2 ;
        RECT 3.404 10.124 5.876 10.156 ;
  LAYER M2 ;
        RECT 3.404 10.06 5.876 10.092 ;
  LAYER M2 ;
        RECT 3.404 9.996 5.876 10.028 ;
  LAYER M2 ;
        RECT 3.404 9.932 5.876 9.964 ;
  LAYER M2 ;
        RECT 3.404 9.868 5.876 9.9 ;
  LAYER M2 ;
        RECT 3.404 9.804 5.876 9.836 ;
  LAYER M2 ;
        RECT 3.404 9.74 5.876 9.772 ;
  LAYER M2 ;
        RECT 3.404 9.676 5.876 9.708 ;
  LAYER M2 ;
        RECT 3.404 9.612 5.876 9.644 ;
  LAYER M2 ;
        RECT 3.404 9.548 5.876 9.58 ;
  LAYER M2 ;
        RECT 3.404 9.484 5.876 9.516 ;
  LAYER M2 ;
        RECT 3.404 9.42 5.876 9.452 ;
  LAYER M2 ;
        RECT 3.404 9.356 5.876 9.388 ;
  LAYER M2 ;
        RECT 3.404 9.292 5.876 9.324 ;
  LAYER M2 ;
        RECT 3.404 9.228 5.876 9.26 ;
  LAYER M2 ;
        RECT 3.404 9.164 5.876 9.196 ;
  LAYER M2 ;
        RECT 3.404 9.1 5.876 9.132 ;
  LAYER M2 ;
        RECT 3.404 9.036 5.876 9.068 ;
  LAYER M2 ;
        RECT 3.404 8.972 5.876 9.004 ;
  LAYER M2 ;
        RECT 3.404 8.908 5.876 8.94 ;
  LAYER M2 ;
        RECT 3.404 8.844 5.876 8.876 ;
  LAYER M2 ;
        RECT 3.404 8.78 5.876 8.812 ;
  LAYER M2 ;
        RECT 3.404 8.716 5.876 8.748 ;
  LAYER M2 ;
        RECT 3.404 8.652 5.876 8.684 ;
  LAYER M2 ;
        RECT 3.404 8.588 5.876 8.62 ;
  LAYER M2 ;
        RECT 3.404 8.524 5.876 8.556 ;
  LAYER M2 ;
        RECT 3.404 8.46 5.876 8.492 ;
  LAYER M2 ;
        RECT 3.404 8.396 5.876 8.428 ;
  LAYER M2 ;
        RECT 3.404 8.332 5.876 8.364 ;
  LAYER M2 ;
        RECT 3.404 8.268 5.876 8.3 ;
  LAYER M2 ;
        RECT 3.404 8.204 5.876 8.236 ;
  LAYER M2 ;
        RECT 3.404 8.14 5.876 8.172 ;
  LAYER M2 ;
        RECT 3.404 8.076 5.876 8.108 ;
  LAYER M2 ;
        RECT 3.404 8.012 5.876 8.044 ;
  LAYER M3 ;
        RECT 5.824 7.86 5.856 10.368 ;
  LAYER M3 ;
        RECT 5.76 7.86 5.792 10.368 ;
  LAYER M3 ;
        RECT 5.696 7.86 5.728 10.368 ;
  LAYER M3 ;
        RECT 5.632 7.86 5.664 10.368 ;
  LAYER M3 ;
        RECT 5.568 7.86 5.6 10.368 ;
  LAYER M3 ;
        RECT 5.504 7.86 5.536 10.368 ;
  LAYER M3 ;
        RECT 5.44 7.86 5.472 10.368 ;
  LAYER M3 ;
        RECT 5.376 7.86 5.408 10.368 ;
  LAYER M3 ;
        RECT 5.312 7.86 5.344 10.368 ;
  LAYER M3 ;
        RECT 5.248 7.86 5.28 10.368 ;
  LAYER M3 ;
        RECT 5.184 7.86 5.216 10.368 ;
  LAYER M3 ;
        RECT 5.12 7.86 5.152 10.368 ;
  LAYER M3 ;
        RECT 5.056 7.86 5.088 10.368 ;
  LAYER M3 ;
        RECT 4.992 7.86 5.024 10.368 ;
  LAYER M3 ;
        RECT 4.928 7.86 4.96 10.368 ;
  LAYER M3 ;
        RECT 4.864 7.86 4.896 10.368 ;
  LAYER M3 ;
        RECT 4.8 7.86 4.832 10.368 ;
  LAYER M3 ;
        RECT 4.736 7.86 4.768 10.368 ;
  LAYER M3 ;
        RECT 4.672 7.86 4.704 10.368 ;
  LAYER M3 ;
        RECT 4.608 7.86 4.64 10.368 ;
  LAYER M3 ;
        RECT 4.544 7.86 4.576 10.368 ;
  LAYER M3 ;
        RECT 4.48 7.86 4.512 10.368 ;
  LAYER M3 ;
        RECT 4.416 7.86 4.448 10.368 ;
  LAYER M3 ;
        RECT 4.352 7.86 4.384 10.368 ;
  LAYER M3 ;
        RECT 4.288 7.86 4.32 10.368 ;
  LAYER M3 ;
        RECT 4.224 7.86 4.256 10.368 ;
  LAYER M3 ;
        RECT 4.16 7.86 4.192 10.368 ;
  LAYER M3 ;
        RECT 4.096 7.86 4.128 10.368 ;
  LAYER M3 ;
        RECT 4.032 7.86 4.064 10.368 ;
  LAYER M3 ;
        RECT 3.968 7.86 4 10.368 ;
  LAYER M3 ;
        RECT 3.904 7.86 3.936 10.368 ;
  LAYER M3 ;
        RECT 3.84 7.86 3.872 10.368 ;
  LAYER M3 ;
        RECT 3.776 7.86 3.808 10.368 ;
  LAYER M3 ;
        RECT 3.712 7.86 3.744 10.368 ;
  LAYER M3 ;
        RECT 3.648 7.86 3.68 10.368 ;
  LAYER M3 ;
        RECT 3.584 7.86 3.616 10.368 ;
  LAYER M3 ;
        RECT 3.52 7.86 3.552 10.368 ;
  LAYER M3 ;
        RECT 3.424 7.86 3.456 10.368 ;
  LAYER M1 ;
        RECT 5.839 7.896 5.841 10.332 ;
  LAYER M1 ;
        RECT 5.759 7.896 5.761 10.332 ;
  LAYER M1 ;
        RECT 5.679 7.896 5.681 10.332 ;
  LAYER M1 ;
        RECT 5.599 7.896 5.601 10.332 ;
  LAYER M1 ;
        RECT 5.519 7.896 5.521 10.332 ;
  LAYER M1 ;
        RECT 5.439 7.896 5.441 10.332 ;
  LAYER M1 ;
        RECT 5.359 7.896 5.361 10.332 ;
  LAYER M1 ;
        RECT 5.279 7.896 5.281 10.332 ;
  LAYER M1 ;
        RECT 5.199 7.896 5.201 10.332 ;
  LAYER M1 ;
        RECT 5.119 7.896 5.121 10.332 ;
  LAYER M1 ;
        RECT 5.039 7.896 5.041 10.332 ;
  LAYER M1 ;
        RECT 4.959 7.896 4.961 10.332 ;
  LAYER M1 ;
        RECT 4.879 7.896 4.881 10.332 ;
  LAYER M1 ;
        RECT 4.799 7.896 4.801 10.332 ;
  LAYER M1 ;
        RECT 4.719 7.896 4.721 10.332 ;
  LAYER M1 ;
        RECT 4.639 7.896 4.641 10.332 ;
  LAYER M1 ;
        RECT 4.559 7.896 4.561 10.332 ;
  LAYER M1 ;
        RECT 4.479 7.896 4.481 10.332 ;
  LAYER M1 ;
        RECT 4.399 7.896 4.401 10.332 ;
  LAYER M1 ;
        RECT 4.319 7.896 4.321 10.332 ;
  LAYER M1 ;
        RECT 4.239 7.896 4.241 10.332 ;
  LAYER M1 ;
        RECT 4.159 7.896 4.161 10.332 ;
  LAYER M1 ;
        RECT 4.079 7.896 4.081 10.332 ;
  LAYER M1 ;
        RECT 3.999 7.896 4.001 10.332 ;
  LAYER M1 ;
        RECT 3.919 7.896 3.921 10.332 ;
  LAYER M1 ;
        RECT 3.839 7.896 3.841 10.332 ;
  LAYER M1 ;
        RECT 3.759 7.896 3.761 10.332 ;
  LAYER M1 ;
        RECT 3.679 7.896 3.681 10.332 ;
  LAYER M1 ;
        RECT 3.599 7.896 3.601 10.332 ;
  LAYER M1 ;
        RECT 3.519 7.896 3.521 10.332 ;
  LAYER M2 ;
        RECT 3.44 10.331 5.84 10.333 ;
  LAYER M2 ;
        RECT 3.44 10.247 5.84 10.249 ;
  LAYER M2 ;
        RECT 3.44 10.163 5.84 10.165 ;
  LAYER M2 ;
        RECT 3.44 10.079 5.84 10.081 ;
  LAYER M2 ;
        RECT 3.44 9.995 5.84 9.997 ;
  LAYER M2 ;
        RECT 3.44 9.911 5.84 9.913 ;
  LAYER M2 ;
        RECT 3.44 9.827 5.84 9.829 ;
  LAYER M2 ;
        RECT 3.44 9.743 5.84 9.745 ;
  LAYER M2 ;
        RECT 3.44 9.659 5.84 9.661 ;
  LAYER M2 ;
        RECT 3.44 9.575 5.84 9.577 ;
  LAYER M2 ;
        RECT 3.44 9.491 5.84 9.493 ;
  LAYER M2 ;
        RECT 3.44 9.407 5.84 9.409 ;
  LAYER M2 ;
        RECT 3.44 9.3235 5.84 9.3255 ;
  LAYER M2 ;
        RECT 3.44 9.239 5.84 9.241 ;
  LAYER M2 ;
        RECT 3.44 9.155 5.84 9.157 ;
  LAYER M2 ;
        RECT 3.44 9.071 5.84 9.073 ;
  LAYER M2 ;
        RECT 3.44 8.987 5.84 8.989 ;
  LAYER M2 ;
        RECT 3.44 8.903 5.84 8.905 ;
  LAYER M2 ;
        RECT 3.44 8.819 5.84 8.821 ;
  LAYER M2 ;
        RECT 3.44 8.735 5.84 8.737 ;
  LAYER M2 ;
        RECT 3.44 8.651 5.84 8.653 ;
  LAYER M2 ;
        RECT 3.44 8.567 5.84 8.569 ;
  LAYER M2 ;
        RECT 3.44 8.483 5.84 8.485 ;
  LAYER M2 ;
        RECT 3.44 8.399 5.84 8.401 ;
  LAYER M2 ;
        RECT 3.44 8.315 5.84 8.317 ;
  LAYER M2 ;
        RECT 3.44 8.231 5.84 8.233 ;
  LAYER M2 ;
        RECT 3.44 8.147 5.84 8.149 ;
  LAYER M2 ;
        RECT 3.44 8.063 5.84 8.065 ;
  LAYER M2 ;
        RECT 3.44 7.979 5.84 7.981 ;
  LAYER M1 ;
        RECT 5.824 4.92 5.856 7.428 ;
  LAYER M1 ;
        RECT 5.76 4.92 5.792 7.428 ;
  LAYER M1 ;
        RECT 5.696 4.92 5.728 7.428 ;
  LAYER M1 ;
        RECT 5.632 4.92 5.664 7.428 ;
  LAYER M1 ;
        RECT 5.568 4.92 5.6 7.428 ;
  LAYER M1 ;
        RECT 5.504 4.92 5.536 7.428 ;
  LAYER M1 ;
        RECT 5.44 4.92 5.472 7.428 ;
  LAYER M1 ;
        RECT 5.376 4.92 5.408 7.428 ;
  LAYER M1 ;
        RECT 5.312 4.92 5.344 7.428 ;
  LAYER M1 ;
        RECT 5.248 4.92 5.28 7.428 ;
  LAYER M1 ;
        RECT 5.184 4.92 5.216 7.428 ;
  LAYER M1 ;
        RECT 5.12 4.92 5.152 7.428 ;
  LAYER M1 ;
        RECT 5.056 4.92 5.088 7.428 ;
  LAYER M1 ;
        RECT 4.992 4.92 5.024 7.428 ;
  LAYER M1 ;
        RECT 4.928 4.92 4.96 7.428 ;
  LAYER M1 ;
        RECT 4.864 4.92 4.896 7.428 ;
  LAYER M1 ;
        RECT 4.8 4.92 4.832 7.428 ;
  LAYER M1 ;
        RECT 4.736 4.92 4.768 7.428 ;
  LAYER M1 ;
        RECT 4.672 4.92 4.704 7.428 ;
  LAYER M1 ;
        RECT 4.608 4.92 4.64 7.428 ;
  LAYER M1 ;
        RECT 4.544 4.92 4.576 7.428 ;
  LAYER M1 ;
        RECT 4.48 4.92 4.512 7.428 ;
  LAYER M1 ;
        RECT 4.416 4.92 4.448 7.428 ;
  LAYER M1 ;
        RECT 4.352 4.92 4.384 7.428 ;
  LAYER M1 ;
        RECT 4.288 4.92 4.32 7.428 ;
  LAYER M1 ;
        RECT 4.224 4.92 4.256 7.428 ;
  LAYER M1 ;
        RECT 4.16 4.92 4.192 7.428 ;
  LAYER M1 ;
        RECT 4.096 4.92 4.128 7.428 ;
  LAYER M1 ;
        RECT 4.032 4.92 4.064 7.428 ;
  LAYER M1 ;
        RECT 3.968 4.92 4 7.428 ;
  LAYER M1 ;
        RECT 3.904 4.92 3.936 7.428 ;
  LAYER M1 ;
        RECT 3.84 4.92 3.872 7.428 ;
  LAYER M1 ;
        RECT 3.776 4.92 3.808 7.428 ;
  LAYER M1 ;
        RECT 3.712 4.92 3.744 7.428 ;
  LAYER M1 ;
        RECT 3.648 4.92 3.68 7.428 ;
  LAYER M1 ;
        RECT 3.584 4.92 3.616 7.428 ;
  LAYER M1 ;
        RECT 3.52 4.92 3.552 7.428 ;
  LAYER M2 ;
        RECT 3.404 7.312 5.876 7.344 ;
  LAYER M2 ;
        RECT 3.404 7.248 5.876 7.28 ;
  LAYER M2 ;
        RECT 3.404 7.184 5.876 7.216 ;
  LAYER M2 ;
        RECT 3.404 7.12 5.876 7.152 ;
  LAYER M2 ;
        RECT 3.404 7.056 5.876 7.088 ;
  LAYER M2 ;
        RECT 3.404 6.992 5.876 7.024 ;
  LAYER M2 ;
        RECT 3.404 6.928 5.876 6.96 ;
  LAYER M2 ;
        RECT 3.404 6.864 5.876 6.896 ;
  LAYER M2 ;
        RECT 3.404 6.8 5.876 6.832 ;
  LAYER M2 ;
        RECT 3.404 6.736 5.876 6.768 ;
  LAYER M2 ;
        RECT 3.404 6.672 5.876 6.704 ;
  LAYER M2 ;
        RECT 3.404 6.608 5.876 6.64 ;
  LAYER M2 ;
        RECT 3.404 6.544 5.876 6.576 ;
  LAYER M2 ;
        RECT 3.404 6.48 5.876 6.512 ;
  LAYER M2 ;
        RECT 3.404 6.416 5.876 6.448 ;
  LAYER M2 ;
        RECT 3.404 6.352 5.876 6.384 ;
  LAYER M2 ;
        RECT 3.404 6.288 5.876 6.32 ;
  LAYER M2 ;
        RECT 3.404 6.224 5.876 6.256 ;
  LAYER M2 ;
        RECT 3.404 6.16 5.876 6.192 ;
  LAYER M2 ;
        RECT 3.404 6.096 5.876 6.128 ;
  LAYER M2 ;
        RECT 3.404 6.032 5.876 6.064 ;
  LAYER M2 ;
        RECT 3.404 5.968 5.876 6 ;
  LAYER M2 ;
        RECT 3.404 5.904 5.876 5.936 ;
  LAYER M2 ;
        RECT 3.404 5.84 5.876 5.872 ;
  LAYER M2 ;
        RECT 3.404 5.776 5.876 5.808 ;
  LAYER M2 ;
        RECT 3.404 5.712 5.876 5.744 ;
  LAYER M2 ;
        RECT 3.404 5.648 5.876 5.68 ;
  LAYER M2 ;
        RECT 3.404 5.584 5.876 5.616 ;
  LAYER M2 ;
        RECT 3.404 5.52 5.876 5.552 ;
  LAYER M2 ;
        RECT 3.404 5.456 5.876 5.488 ;
  LAYER M2 ;
        RECT 3.404 5.392 5.876 5.424 ;
  LAYER M2 ;
        RECT 3.404 5.328 5.876 5.36 ;
  LAYER M2 ;
        RECT 3.404 5.264 5.876 5.296 ;
  LAYER M2 ;
        RECT 3.404 5.2 5.876 5.232 ;
  LAYER M2 ;
        RECT 3.404 5.136 5.876 5.168 ;
  LAYER M2 ;
        RECT 3.404 5.072 5.876 5.104 ;
  LAYER M3 ;
        RECT 5.824 4.92 5.856 7.428 ;
  LAYER M3 ;
        RECT 5.76 4.92 5.792 7.428 ;
  LAYER M3 ;
        RECT 5.696 4.92 5.728 7.428 ;
  LAYER M3 ;
        RECT 5.632 4.92 5.664 7.428 ;
  LAYER M3 ;
        RECT 5.568 4.92 5.6 7.428 ;
  LAYER M3 ;
        RECT 5.504 4.92 5.536 7.428 ;
  LAYER M3 ;
        RECT 5.44 4.92 5.472 7.428 ;
  LAYER M3 ;
        RECT 5.376 4.92 5.408 7.428 ;
  LAYER M3 ;
        RECT 5.312 4.92 5.344 7.428 ;
  LAYER M3 ;
        RECT 5.248 4.92 5.28 7.428 ;
  LAYER M3 ;
        RECT 5.184 4.92 5.216 7.428 ;
  LAYER M3 ;
        RECT 5.12 4.92 5.152 7.428 ;
  LAYER M3 ;
        RECT 5.056 4.92 5.088 7.428 ;
  LAYER M3 ;
        RECT 4.992 4.92 5.024 7.428 ;
  LAYER M3 ;
        RECT 4.928 4.92 4.96 7.428 ;
  LAYER M3 ;
        RECT 4.864 4.92 4.896 7.428 ;
  LAYER M3 ;
        RECT 4.8 4.92 4.832 7.428 ;
  LAYER M3 ;
        RECT 4.736 4.92 4.768 7.428 ;
  LAYER M3 ;
        RECT 4.672 4.92 4.704 7.428 ;
  LAYER M3 ;
        RECT 4.608 4.92 4.64 7.428 ;
  LAYER M3 ;
        RECT 4.544 4.92 4.576 7.428 ;
  LAYER M3 ;
        RECT 4.48 4.92 4.512 7.428 ;
  LAYER M3 ;
        RECT 4.416 4.92 4.448 7.428 ;
  LAYER M3 ;
        RECT 4.352 4.92 4.384 7.428 ;
  LAYER M3 ;
        RECT 4.288 4.92 4.32 7.428 ;
  LAYER M3 ;
        RECT 4.224 4.92 4.256 7.428 ;
  LAYER M3 ;
        RECT 4.16 4.92 4.192 7.428 ;
  LAYER M3 ;
        RECT 4.096 4.92 4.128 7.428 ;
  LAYER M3 ;
        RECT 4.032 4.92 4.064 7.428 ;
  LAYER M3 ;
        RECT 3.968 4.92 4 7.428 ;
  LAYER M3 ;
        RECT 3.904 4.92 3.936 7.428 ;
  LAYER M3 ;
        RECT 3.84 4.92 3.872 7.428 ;
  LAYER M3 ;
        RECT 3.776 4.92 3.808 7.428 ;
  LAYER M3 ;
        RECT 3.712 4.92 3.744 7.428 ;
  LAYER M3 ;
        RECT 3.648 4.92 3.68 7.428 ;
  LAYER M3 ;
        RECT 3.584 4.92 3.616 7.428 ;
  LAYER M3 ;
        RECT 3.52 4.92 3.552 7.428 ;
  LAYER M3 ;
        RECT 3.424 4.92 3.456 7.428 ;
  LAYER M1 ;
        RECT 5.839 4.956 5.841 7.392 ;
  LAYER M1 ;
        RECT 5.759 4.956 5.761 7.392 ;
  LAYER M1 ;
        RECT 5.679 4.956 5.681 7.392 ;
  LAYER M1 ;
        RECT 5.599 4.956 5.601 7.392 ;
  LAYER M1 ;
        RECT 5.519 4.956 5.521 7.392 ;
  LAYER M1 ;
        RECT 5.439 4.956 5.441 7.392 ;
  LAYER M1 ;
        RECT 5.359 4.956 5.361 7.392 ;
  LAYER M1 ;
        RECT 5.279 4.956 5.281 7.392 ;
  LAYER M1 ;
        RECT 5.199 4.956 5.201 7.392 ;
  LAYER M1 ;
        RECT 5.119 4.956 5.121 7.392 ;
  LAYER M1 ;
        RECT 5.039 4.956 5.041 7.392 ;
  LAYER M1 ;
        RECT 4.959 4.956 4.961 7.392 ;
  LAYER M1 ;
        RECT 4.879 4.956 4.881 7.392 ;
  LAYER M1 ;
        RECT 4.799 4.956 4.801 7.392 ;
  LAYER M1 ;
        RECT 4.719 4.956 4.721 7.392 ;
  LAYER M1 ;
        RECT 4.639 4.956 4.641 7.392 ;
  LAYER M1 ;
        RECT 4.559 4.956 4.561 7.392 ;
  LAYER M1 ;
        RECT 4.479 4.956 4.481 7.392 ;
  LAYER M1 ;
        RECT 4.399 4.956 4.401 7.392 ;
  LAYER M1 ;
        RECT 4.319 4.956 4.321 7.392 ;
  LAYER M1 ;
        RECT 4.239 4.956 4.241 7.392 ;
  LAYER M1 ;
        RECT 4.159 4.956 4.161 7.392 ;
  LAYER M1 ;
        RECT 4.079 4.956 4.081 7.392 ;
  LAYER M1 ;
        RECT 3.999 4.956 4.001 7.392 ;
  LAYER M1 ;
        RECT 3.919 4.956 3.921 7.392 ;
  LAYER M1 ;
        RECT 3.839 4.956 3.841 7.392 ;
  LAYER M1 ;
        RECT 3.759 4.956 3.761 7.392 ;
  LAYER M1 ;
        RECT 3.679 4.956 3.681 7.392 ;
  LAYER M1 ;
        RECT 3.599 4.956 3.601 7.392 ;
  LAYER M1 ;
        RECT 3.519 4.956 3.521 7.392 ;
  LAYER M2 ;
        RECT 3.44 7.391 5.84 7.393 ;
  LAYER M2 ;
        RECT 3.44 7.307 5.84 7.309 ;
  LAYER M2 ;
        RECT 3.44 7.223 5.84 7.225 ;
  LAYER M2 ;
        RECT 3.44 7.139 5.84 7.141 ;
  LAYER M2 ;
        RECT 3.44 7.055 5.84 7.057 ;
  LAYER M2 ;
        RECT 3.44 6.971 5.84 6.973 ;
  LAYER M2 ;
        RECT 3.44 6.887 5.84 6.889 ;
  LAYER M2 ;
        RECT 3.44 6.803 5.84 6.805 ;
  LAYER M2 ;
        RECT 3.44 6.719 5.84 6.721 ;
  LAYER M2 ;
        RECT 3.44 6.635 5.84 6.637 ;
  LAYER M2 ;
        RECT 3.44 6.551 5.84 6.553 ;
  LAYER M2 ;
        RECT 3.44 6.467 5.84 6.469 ;
  LAYER M2 ;
        RECT 3.44 6.3835 5.84 6.3855 ;
  LAYER M2 ;
        RECT 3.44 6.299 5.84 6.301 ;
  LAYER M2 ;
        RECT 3.44 6.215 5.84 6.217 ;
  LAYER M2 ;
        RECT 3.44 6.131 5.84 6.133 ;
  LAYER M2 ;
        RECT 3.44 6.047 5.84 6.049 ;
  LAYER M2 ;
        RECT 3.44 5.963 5.84 5.965 ;
  LAYER M2 ;
        RECT 3.44 5.879 5.84 5.881 ;
  LAYER M2 ;
        RECT 3.44 5.795 5.84 5.797 ;
  LAYER M2 ;
        RECT 3.44 5.711 5.84 5.713 ;
  LAYER M2 ;
        RECT 3.44 5.627 5.84 5.629 ;
  LAYER M2 ;
        RECT 3.44 5.543 5.84 5.545 ;
  LAYER M2 ;
        RECT 3.44 5.459 5.84 5.461 ;
  LAYER M2 ;
        RECT 3.44 5.375 5.84 5.377 ;
  LAYER M2 ;
        RECT 3.44 5.291 5.84 5.293 ;
  LAYER M2 ;
        RECT 3.44 5.207 5.84 5.209 ;
  LAYER M2 ;
        RECT 3.44 5.123 5.84 5.125 ;
  LAYER M2 ;
        RECT 3.44 5.039 5.84 5.041 ;
  LAYER M1 ;
        RECT 5.824 1.98 5.856 4.488 ;
  LAYER M1 ;
        RECT 5.76 1.98 5.792 4.488 ;
  LAYER M1 ;
        RECT 5.696 1.98 5.728 4.488 ;
  LAYER M1 ;
        RECT 5.632 1.98 5.664 4.488 ;
  LAYER M1 ;
        RECT 5.568 1.98 5.6 4.488 ;
  LAYER M1 ;
        RECT 5.504 1.98 5.536 4.488 ;
  LAYER M1 ;
        RECT 5.44 1.98 5.472 4.488 ;
  LAYER M1 ;
        RECT 5.376 1.98 5.408 4.488 ;
  LAYER M1 ;
        RECT 5.312 1.98 5.344 4.488 ;
  LAYER M1 ;
        RECT 5.248 1.98 5.28 4.488 ;
  LAYER M1 ;
        RECT 5.184 1.98 5.216 4.488 ;
  LAYER M1 ;
        RECT 5.12 1.98 5.152 4.488 ;
  LAYER M1 ;
        RECT 5.056 1.98 5.088 4.488 ;
  LAYER M1 ;
        RECT 4.992 1.98 5.024 4.488 ;
  LAYER M1 ;
        RECT 4.928 1.98 4.96 4.488 ;
  LAYER M1 ;
        RECT 4.864 1.98 4.896 4.488 ;
  LAYER M1 ;
        RECT 4.8 1.98 4.832 4.488 ;
  LAYER M1 ;
        RECT 4.736 1.98 4.768 4.488 ;
  LAYER M1 ;
        RECT 4.672 1.98 4.704 4.488 ;
  LAYER M1 ;
        RECT 4.608 1.98 4.64 4.488 ;
  LAYER M1 ;
        RECT 4.544 1.98 4.576 4.488 ;
  LAYER M1 ;
        RECT 4.48 1.98 4.512 4.488 ;
  LAYER M1 ;
        RECT 4.416 1.98 4.448 4.488 ;
  LAYER M1 ;
        RECT 4.352 1.98 4.384 4.488 ;
  LAYER M1 ;
        RECT 4.288 1.98 4.32 4.488 ;
  LAYER M1 ;
        RECT 4.224 1.98 4.256 4.488 ;
  LAYER M1 ;
        RECT 4.16 1.98 4.192 4.488 ;
  LAYER M1 ;
        RECT 4.096 1.98 4.128 4.488 ;
  LAYER M1 ;
        RECT 4.032 1.98 4.064 4.488 ;
  LAYER M1 ;
        RECT 3.968 1.98 4 4.488 ;
  LAYER M1 ;
        RECT 3.904 1.98 3.936 4.488 ;
  LAYER M1 ;
        RECT 3.84 1.98 3.872 4.488 ;
  LAYER M1 ;
        RECT 3.776 1.98 3.808 4.488 ;
  LAYER M1 ;
        RECT 3.712 1.98 3.744 4.488 ;
  LAYER M1 ;
        RECT 3.648 1.98 3.68 4.488 ;
  LAYER M1 ;
        RECT 3.584 1.98 3.616 4.488 ;
  LAYER M1 ;
        RECT 3.52 1.98 3.552 4.488 ;
  LAYER M2 ;
        RECT 3.404 4.372 5.876 4.404 ;
  LAYER M2 ;
        RECT 3.404 4.308 5.876 4.34 ;
  LAYER M2 ;
        RECT 3.404 4.244 5.876 4.276 ;
  LAYER M2 ;
        RECT 3.404 4.18 5.876 4.212 ;
  LAYER M2 ;
        RECT 3.404 4.116 5.876 4.148 ;
  LAYER M2 ;
        RECT 3.404 4.052 5.876 4.084 ;
  LAYER M2 ;
        RECT 3.404 3.988 5.876 4.02 ;
  LAYER M2 ;
        RECT 3.404 3.924 5.876 3.956 ;
  LAYER M2 ;
        RECT 3.404 3.86 5.876 3.892 ;
  LAYER M2 ;
        RECT 3.404 3.796 5.876 3.828 ;
  LAYER M2 ;
        RECT 3.404 3.732 5.876 3.764 ;
  LAYER M2 ;
        RECT 3.404 3.668 5.876 3.7 ;
  LAYER M2 ;
        RECT 3.404 3.604 5.876 3.636 ;
  LAYER M2 ;
        RECT 3.404 3.54 5.876 3.572 ;
  LAYER M2 ;
        RECT 3.404 3.476 5.876 3.508 ;
  LAYER M2 ;
        RECT 3.404 3.412 5.876 3.444 ;
  LAYER M2 ;
        RECT 3.404 3.348 5.876 3.38 ;
  LAYER M2 ;
        RECT 3.404 3.284 5.876 3.316 ;
  LAYER M2 ;
        RECT 3.404 3.22 5.876 3.252 ;
  LAYER M2 ;
        RECT 3.404 3.156 5.876 3.188 ;
  LAYER M2 ;
        RECT 3.404 3.092 5.876 3.124 ;
  LAYER M2 ;
        RECT 3.404 3.028 5.876 3.06 ;
  LAYER M2 ;
        RECT 3.404 2.964 5.876 2.996 ;
  LAYER M2 ;
        RECT 3.404 2.9 5.876 2.932 ;
  LAYER M2 ;
        RECT 3.404 2.836 5.876 2.868 ;
  LAYER M2 ;
        RECT 3.404 2.772 5.876 2.804 ;
  LAYER M2 ;
        RECT 3.404 2.708 5.876 2.74 ;
  LAYER M2 ;
        RECT 3.404 2.644 5.876 2.676 ;
  LAYER M2 ;
        RECT 3.404 2.58 5.876 2.612 ;
  LAYER M2 ;
        RECT 3.404 2.516 5.876 2.548 ;
  LAYER M2 ;
        RECT 3.404 2.452 5.876 2.484 ;
  LAYER M2 ;
        RECT 3.404 2.388 5.876 2.42 ;
  LAYER M2 ;
        RECT 3.404 2.324 5.876 2.356 ;
  LAYER M2 ;
        RECT 3.404 2.26 5.876 2.292 ;
  LAYER M2 ;
        RECT 3.404 2.196 5.876 2.228 ;
  LAYER M2 ;
        RECT 3.404 2.132 5.876 2.164 ;
  LAYER M3 ;
        RECT 5.824 1.98 5.856 4.488 ;
  LAYER M3 ;
        RECT 5.76 1.98 5.792 4.488 ;
  LAYER M3 ;
        RECT 5.696 1.98 5.728 4.488 ;
  LAYER M3 ;
        RECT 5.632 1.98 5.664 4.488 ;
  LAYER M3 ;
        RECT 5.568 1.98 5.6 4.488 ;
  LAYER M3 ;
        RECT 5.504 1.98 5.536 4.488 ;
  LAYER M3 ;
        RECT 5.44 1.98 5.472 4.488 ;
  LAYER M3 ;
        RECT 5.376 1.98 5.408 4.488 ;
  LAYER M3 ;
        RECT 5.312 1.98 5.344 4.488 ;
  LAYER M3 ;
        RECT 5.248 1.98 5.28 4.488 ;
  LAYER M3 ;
        RECT 5.184 1.98 5.216 4.488 ;
  LAYER M3 ;
        RECT 5.12 1.98 5.152 4.488 ;
  LAYER M3 ;
        RECT 5.056 1.98 5.088 4.488 ;
  LAYER M3 ;
        RECT 4.992 1.98 5.024 4.488 ;
  LAYER M3 ;
        RECT 4.928 1.98 4.96 4.488 ;
  LAYER M3 ;
        RECT 4.864 1.98 4.896 4.488 ;
  LAYER M3 ;
        RECT 4.8 1.98 4.832 4.488 ;
  LAYER M3 ;
        RECT 4.736 1.98 4.768 4.488 ;
  LAYER M3 ;
        RECT 4.672 1.98 4.704 4.488 ;
  LAYER M3 ;
        RECT 4.608 1.98 4.64 4.488 ;
  LAYER M3 ;
        RECT 4.544 1.98 4.576 4.488 ;
  LAYER M3 ;
        RECT 4.48 1.98 4.512 4.488 ;
  LAYER M3 ;
        RECT 4.416 1.98 4.448 4.488 ;
  LAYER M3 ;
        RECT 4.352 1.98 4.384 4.488 ;
  LAYER M3 ;
        RECT 4.288 1.98 4.32 4.488 ;
  LAYER M3 ;
        RECT 4.224 1.98 4.256 4.488 ;
  LAYER M3 ;
        RECT 4.16 1.98 4.192 4.488 ;
  LAYER M3 ;
        RECT 4.096 1.98 4.128 4.488 ;
  LAYER M3 ;
        RECT 4.032 1.98 4.064 4.488 ;
  LAYER M3 ;
        RECT 3.968 1.98 4 4.488 ;
  LAYER M3 ;
        RECT 3.904 1.98 3.936 4.488 ;
  LAYER M3 ;
        RECT 3.84 1.98 3.872 4.488 ;
  LAYER M3 ;
        RECT 3.776 1.98 3.808 4.488 ;
  LAYER M3 ;
        RECT 3.712 1.98 3.744 4.488 ;
  LAYER M3 ;
        RECT 3.648 1.98 3.68 4.488 ;
  LAYER M3 ;
        RECT 3.584 1.98 3.616 4.488 ;
  LAYER M3 ;
        RECT 3.52 1.98 3.552 4.488 ;
  LAYER M3 ;
        RECT 3.424 1.98 3.456 4.488 ;
  LAYER M1 ;
        RECT 5.839 2.016 5.841 4.452 ;
  LAYER M1 ;
        RECT 5.759 2.016 5.761 4.452 ;
  LAYER M1 ;
        RECT 5.679 2.016 5.681 4.452 ;
  LAYER M1 ;
        RECT 5.599 2.016 5.601 4.452 ;
  LAYER M1 ;
        RECT 5.519 2.016 5.521 4.452 ;
  LAYER M1 ;
        RECT 5.439 2.016 5.441 4.452 ;
  LAYER M1 ;
        RECT 5.359 2.016 5.361 4.452 ;
  LAYER M1 ;
        RECT 5.279 2.016 5.281 4.452 ;
  LAYER M1 ;
        RECT 5.199 2.016 5.201 4.452 ;
  LAYER M1 ;
        RECT 5.119 2.016 5.121 4.452 ;
  LAYER M1 ;
        RECT 5.039 2.016 5.041 4.452 ;
  LAYER M1 ;
        RECT 4.959 2.016 4.961 4.452 ;
  LAYER M1 ;
        RECT 4.879 2.016 4.881 4.452 ;
  LAYER M1 ;
        RECT 4.799 2.016 4.801 4.452 ;
  LAYER M1 ;
        RECT 4.719 2.016 4.721 4.452 ;
  LAYER M1 ;
        RECT 4.639 2.016 4.641 4.452 ;
  LAYER M1 ;
        RECT 4.559 2.016 4.561 4.452 ;
  LAYER M1 ;
        RECT 4.479 2.016 4.481 4.452 ;
  LAYER M1 ;
        RECT 4.399 2.016 4.401 4.452 ;
  LAYER M1 ;
        RECT 4.319 2.016 4.321 4.452 ;
  LAYER M1 ;
        RECT 4.239 2.016 4.241 4.452 ;
  LAYER M1 ;
        RECT 4.159 2.016 4.161 4.452 ;
  LAYER M1 ;
        RECT 4.079 2.016 4.081 4.452 ;
  LAYER M1 ;
        RECT 3.999 2.016 4.001 4.452 ;
  LAYER M1 ;
        RECT 3.919 2.016 3.921 4.452 ;
  LAYER M1 ;
        RECT 3.839 2.016 3.841 4.452 ;
  LAYER M1 ;
        RECT 3.759 2.016 3.761 4.452 ;
  LAYER M1 ;
        RECT 3.679 2.016 3.681 4.452 ;
  LAYER M1 ;
        RECT 3.599 2.016 3.601 4.452 ;
  LAYER M1 ;
        RECT 3.519 2.016 3.521 4.452 ;
  LAYER M2 ;
        RECT 3.44 4.451 5.84 4.453 ;
  LAYER M2 ;
        RECT 3.44 4.367 5.84 4.369 ;
  LAYER M2 ;
        RECT 3.44 4.283 5.84 4.285 ;
  LAYER M2 ;
        RECT 3.44 4.199 5.84 4.201 ;
  LAYER M2 ;
        RECT 3.44 4.115 5.84 4.117 ;
  LAYER M2 ;
        RECT 3.44 4.031 5.84 4.033 ;
  LAYER M2 ;
        RECT 3.44 3.947 5.84 3.949 ;
  LAYER M2 ;
        RECT 3.44 3.863 5.84 3.865 ;
  LAYER M2 ;
        RECT 3.44 3.779 5.84 3.781 ;
  LAYER M2 ;
        RECT 3.44 3.695 5.84 3.697 ;
  LAYER M2 ;
        RECT 3.44 3.611 5.84 3.613 ;
  LAYER M2 ;
        RECT 3.44 3.527 5.84 3.529 ;
  LAYER M2 ;
        RECT 3.44 3.4435 5.84 3.4455 ;
  LAYER M2 ;
        RECT 3.44 3.359 5.84 3.361 ;
  LAYER M2 ;
        RECT 3.44 3.275 5.84 3.277 ;
  LAYER M2 ;
        RECT 3.44 3.191 5.84 3.193 ;
  LAYER M2 ;
        RECT 3.44 3.107 5.84 3.109 ;
  LAYER M2 ;
        RECT 3.44 3.023 5.84 3.025 ;
  LAYER M2 ;
        RECT 3.44 2.939 5.84 2.941 ;
  LAYER M2 ;
        RECT 3.44 2.855 5.84 2.857 ;
  LAYER M2 ;
        RECT 3.44 2.771 5.84 2.773 ;
  LAYER M2 ;
        RECT 3.44 2.687 5.84 2.689 ;
  LAYER M2 ;
        RECT 3.44 2.603 5.84 2.605 ;
  LAYER M2 ;
        RECT 3.44 2.519 5.84 2.521 ;
  LAYER M2 ;
        RECT 3.44 2.435 5.84 2.437 ;
  LAYER M2 ;
        RECT 3.44 2.351 5.84 2.353 ;
  LAYER M2 ;
        RECT 3.44 2.267 5.84 2.269 ;
  LAYER M2 ;
        RECT 3.44 2.183 5.84 2.185 ;
  LAYER M2 ;
        RECT 3.44 2.099 5.84 2.101 ;
  LAYER M1 ;
        RECT 2.944 13.74 2.976 16.248 ;
  LAYER M1 ;
        RECT 2.88 13.74 2.912 16.248 ;
  LAYER M1 ;
        RECT 2.816 13.74 2.848 16.248 ;
  LAYER M1 ;
        RECT 2.752 13.74 2.784 16.248 ;
  LAYER M1 ;
        RECT 2.688 13.74 2.72 16.248 ;
  LAYER M1 ;
        RECT 2.624 13.74 2.656 16.248 ;
  LAYER M1 ;
        RECT 2.56 13.74 2.592 16.248 ;
  LAYER M1 ;
        RECT 2.496 13.74 2.528 16.248 ;
  LAYER M1 ;
        RECT 2.432 13.74 2.464 16.248 ;
  LAYER M1 ;
        RECT 2.368 13.74 2.4 16.248 ;
  LAYER M1 ;
        RECT 2.304 13.74 2.336 16.248 ;
  LAYER M1 ;
        RECT 2.24 13.74 2.272 16.248 ;
  LAYER M1 ;
        RECT 2.176 13.74 2.208 16.248 ;
  LAYER M1 ;
        RECT 2.112 13.74 2.144 16.248 ;
  LAYER M1 ;
        RECT 2.048 13.74 2.08 16.248 ;
  LAYER M1 ;
        RECT 1.984 13.74 2.016 16.248 ;
  LAYER M1 ;
        RECT 1.92 13.74 1.952 16.248 ;
  LAYER M1 ;
        RECT 1.856 13.74 1.888 16.248 ;
  LAYER M1 ;
        RECT 1.792 13.74 1.824 16.248 ;
  LAYER M1 ;
        RECT 1.728 13.74 1.76 16.248 ;
  LAYER M1 ;
        RECT 1.664 13.74 1.696 16.248 ;
  LAYER M1 ;
        RECT 1.6 13.74 1.632 16.248 ;
  LAYER M1 ;
        RECT 1.536 13.74 1.568 16.248 ;
  LAYER M1 ;
        RECT 1.472 13.74 1.504 16.248 ;
  LAYER M1 ;
        RECT 1.408 13.74 1.44 16.248 ;
  LAYER M1 ;
        RECT 1.344 13.74 1.376 16.248 ;
  LAYER M1 ;
        RECT 1.28 13.74 1.312 16.248 ;
  LAYER M1 ;
        RECT 1.216 13.74 1.248 16.248 ;
  LAYER M1 ;
        RECT 1.152 13.74 1.184 16.248 ;
  LAYER M1 ;
        RECT 1.088 13.74 1.12 16.248 ;
  LAYER M1 ;
        RECT 1.024 13.74 1.056 16.248 ;
  LAYER M1 ;
        RECT 0.96 13.74 0.992 16.248 ;
  LAYER M1 ;
        RECT 0.896 13.74 0.928 16.248 ;
  LAYER M1 ;
        RECT 0.832 13.74 0.864 16.248 ;
  LAYER M1 ;
        RECT 0.768 13.74 0.8 16.248 ;
  LAYER M1 ;
        RECT 0.704 13.74 0.736 16.248 ;
  LAYER M1 ;
        RECT 0.64 13.74 0.672 16.248 ;
  LAYER M2 ;
        RECT 0.524 16.132 2.996 16.164 ;
  LAYER M2 ;
        RECT 0.524 16.068 2.996 16.1 ;
  LAYER M2 ;
        RECT 0.524 16.004 2.996 16.036 ;
  LAYER M2 ;
        RECT 0.524 15.94 2.996 15.972 ;
  LAYER M2 ;
        RECT 0.524 15.876 2.996 15.908 ;
  LAYER M2 ;
        RECT 0.524 15.812 2.996 15.844 ;
  LAYER M2 ;
        RECT 0.524 15.748 2.996 15.78 ;
  LAYER M2 ;
        RECT 0.524 15.684 2.996 15.716 ;
  LAYER M2 ;
        RECT 0.524 15.62 2.996 15.652 ;
  LAYER M2 ;
        RECT 0.524 15.556 2.996 15.588 ;
  LAYER M2 ;
        RECT 0.524 15.492 2.996 15.524 ;
  LAYER M2 ;
        RECT 0.524 15.428 2.996 15.46 ;
  LAYER M2 ;
        RECT 0.524 15.364 2.996 15.396 ;
  LAYER M2 ;
        RECT 0.524 15.3 2.996 15.332 ;
  LAYER M2 ;
        RECT 0.524 15.236 2.996 15.268 ;
  LAYER M2 ;
        RECT 0.524 15.172 2.996 15.204 ;
  LAYER M2 ;
        RECT 0.524 15.108 2.996 15.14 ;
  LAYER M2 ;
        RECT 0.524 15.044 2.996 15.076 ;
  LAYER M2 ;
        RECT 0.524 14.98 2.996 15.012 ;
  LAYER M2 ;
        RECT 0.524 14.916 2.996 14.948 ;
  LAYER M2 ;
        RECT 0.524 14.852 2.996 14.884 ;
  LAYER M2 ;
        RECT 0.524 14.788 2.996 14.82 ;
  LAYER M2 ;
        RECT 0.524 14.724 2.996 14.756 ;
  LAYER M2 ;
        RECT 0.524 14.66 2.996 14.692 ;
  LAYER M2 ;
        RECT 0.524 14.596 2.996 14.628 ;
  LAYER M2 ;
        RECT 0.524 14.532 2.996 14.564 ;
  LAYER M2 ;
        RECT 0.524 14.468 2.996 14.5 ;
  LAYER M2 ;
        RECT 0.524 14.404 2.996 14.436 ;
  LAYER M2 ;
        RECT 0.524 14.34 2.996 14.372 ;
  LAYER M2 ;
        RECT 0.524 14.276 2.996 14.308 ;
  LAYER M2 ;
        RECT 0.524 14.212 2.996 14.244 ;
  LAYER M2 ;
        RECT 0.524 14.148 2.996 14.18 ;
  LAYER M2 ;
        RECT 0.524 14.084 2.996 14.116 ;
  LAYER M2 ;
        RECT 0.524 14.02 2.996 14.052 ;
  LAYER M2 ;
        RECT 0.524 13.956 2.996 13.988 ;
  LAYER M2 ;
        RECT 0.524 13.892 2.996 13.924 ;
  LAYER M3 ;
        RECT 2.944 13.74 2.976 16.248 ;
  LAYER M3 ;
        RECT 2.88 13.74 2.912 16.248 ;
  LAYER M3 ;
        RECT 2.816 13.74 2.848 16.248 ;
  LAYER M3 ;
        RECT 2.752 13.74 2.784 16.248 ;
  LAYER M3 ;
        RECT 2.688 13.74 2.72 16.248 ;
  LAYER M3 ;
        RECT 2.624 13.74 2.656 16.248 ;
  LAYER M3 ;
        RECT 2.56 13.74 2.592 16.248 ;
  LAYER M3 ;
        RECT 2.496 13.74 2.528 16.248 ;
  LAYER M3 ;
        RECT 2.432 13.74 2.464 16.248 ;
  LAYER M3 ;
        RECT 2.368 13.74 2.4 16.248 ;
  LAYER M3 ;
        RECT 2.304 13.74 2.336 16.248 ;
  LAYER M3 ;
        RECT 2.24 13.74 2.272 16.248 ;
  LAYER M3 ;
        RECT 2.176 13.74 2.208 16.248 ;
  LAYER M3 ;
        RECT 2.112 13.74 2.144 16.248 ;
  LAYER M3 ;
        RECT 2.048 13.74 2.08 16.248 ;
  LAYER M3 ;
        RECT 1.984 13.74 2.016 16.248 ;
  LAYER M3 ;
        RECT 1.92 13.74 1.952 16.248 ;
  LAYER M3 ;
        RECT 1.856 13.74 1.888 16.248 ;
  LAYER M3 ;
        RECT 1.792 13.74 1.824 16.248 ;
  LAYER M3 ;
        RECT 1.728 13.74 1.76 16.248 ;
  LAYER M3 ;
        RECT 1.664 13.74 1.696 16.248 ;
  LAYER M3 ;
        RECT 1.6 13.74 1.632 16.248 ;
  LAYER M3 ;
        RECT 1.536 13.74 1.568 16.248 ;
  LAYER M3 ;
        RECT 1.472 13.74 1.504 16.248 ;
  LAYER M3 ;
        RECT 1.408 13.74 1.44 16.248 ;
  LAYER M3 ;
        RECT 1.344 13.74 1.376 16.248 ;
  LAYER M3 ;
        RECT 1.28 13.74 1.312 16.248 ;
  LAYER M3 ;
        RECT 1.216 13.74 1.248 16.248 ;
  LAYER M3 ;
        RECT 1.152 13.74 1.184 16.248 ;
  LAYER M3 ;
        RECT 1.088 13.74 1.12 16.248 ;
  LAYER M3 ;
        RECT 1.024 13.74 1.056 16.248 ;
  LAYER M3 ;
        RECT 0.96 13.74 0.992 16.248 ;
  LAYER M3 ;
        RECT 0.896 13.74 0.928 16.248 ;
  LAYER M3 ;
        RECT 0.832 13.74 0.864 16.248 ;
  LAYER M3 ;
        RECT 0.768 13.74 0.8 16.248 ;
  LAYER M3 ;
        RECT 0.704 13.74 0.736 16.248 ;
  LAYER M3 ;
        RECT 0.64 13.74 0.672 16.248 ;
  LAYER M3 ;
        RECT 0.544 13.74 0.576 16.248 ;
  LAYER M1 ;
        RECT 2.959 13.776 2.961 16.212 ;
  LAYER M1 ;
        RECT 2.879 13.776 2.881 16.212 ;
  LAYER M1 ;
        RECT 2.799 13.776 2.801 16.212 ;
  LAYER M1 ;
        RECT 2.719 13.776 2.721 16.212 ;
  LAYER M1 ;
        RECT 2.639 13.776 2.641 16.212 ;
  LAYER M1 ;
        RECT 2.559 13.776 2.561 16.212 ;
  LAYER M1 ;
        RECT 2.479 13.776 2.481 16.212 ;
  LAYER M1 ;
        RECT 2.399 13.776 2.401 16.212 ;
  LAYER M1 ;
        RECT 2.319 13.776 2.321 16.212 ;
  LAYER M1 ;
        RECT 2.239 13.776 2.241 16.212 ;
  LAYER M1 ;
        RECT 2.159 13.776 2.161 16.212 ;
  LAYER M1 ;
        RECT 2.079 13.776 2.081 16.212 ;
  LAYER M1 ;
        RECT 1.999 13.776 2.001 16.212 ;
  LAYER M1 ;
        RECT 1.919 13.776 1.921 16.212 ;
  LAYER M1 ;
        RECT 1.839 13.776 1.841 16.212 ;
  LAYER M1 ;
        RECT 1.759 13.776 1.761 16.212 ;
  LAYER M1 ;
        RECT 1.679 13.776 1.681 16.212 ;
  LAYER M1 ;
        RECT 1.599 13.776 1.601 16.212 ;
  LAYER M1 ;
        RECT 1.519 13.776 1.521 16.212 ;
  LAYER M1 ;
        RECT 1.439 13.776 1.441 16.212 ;
  LAYER M1 ;
        RECT 1.359 13.776 1.361 16.212 ;
  LAYER M1 ;
        RECT 1.279 13.776 1.281 16.212 ;
  LAYER M1 ;
        RECT 1.199 13.776 1.201 16.212 ;
  LAYER M1 ;
        RECT 1.119 13.776 1.121 16.212 ;
  LAYER M1 ;
        RECT 1.039 13.776 1.041 16.212 ;
  LAYER M1 ;
        RECT 0.959 13.776 0.961 16.212 ;
  LAYER M1 ;
        RECT 0.879 13.776 0.881 16.212 ;
  LAYER M1 ;
        RECT 0.799 13.776 0.801 16.212 ;
  LAYER M1 ;
        RECT 0.719 13.776 0.721 16.212 ;
  LAYER M1 ;
        RECT 0.639 13.776 0.641 16.212 ;
  LAYER M2 ;
        RECT 0.56 16.211 2.96 16.213 ;
  LAYER M2 ;
        RECT 0.56 16.127 2.96 16.129 ;
  LAYER M2 ;
        RECT 0.56 16.043 2.96 16.045 ;
  LAYER M2 ;
        RECT 0.56 15.959 2.96 15.961 ;
  LAYER M2 ;
        RECT 0.56 15.875 2.96 15.877 ;
  LAYER M2 ;
        RECT 0.56 15.791 2.96 15.793 ;
  LAYER M2 ;
        RECT 0.56 15.707 2.96 15.709 ;
  LAYER M2 ;
        RECT 0.56 15.623 2.96 15.625 ;
  LAYER M2 ;
        RECT 0.56 15.539 2.96 15.541 ;
  LAYER M2 ;
        RECT 0.56 15.455 2.96 15.457 ;
  LAYER M2 ;
        RECT 0.56 15.371 2.96 15.373 ;
  LAYER M2 ;
        RECT 0.56 15.287 2.96 15.289 ;
  LAYER M2 ;
        RECT 0.56 15.2035 2.96 15.2055 ;
  LAYER M2 ;
        RECT 0.56 15.119 2.96 15.121 ;
  LAYER M2 ;
        RECT 0.56 15.035 2.96 15.037 ;
  LAYER M2 ;
        RECT 0.56 14.951 2.96 14.953 ;
  LAYER M2 ;
        RECT 0.56 14.867 2.96 14.869 ;
  LAYER M2 ;
        RECT 0.56 14.783 2.96 14.785 ;
  LAYER M2 ;
        RECT 0.56 14.699 2.96 14.701 ;
  LAYER M2 ;
        RECT 0.56 14.615 2.96 14.617 ;
  LAYER M2 ;
        RECT 0.56 14.531 2.96 14.533 ;
  LAYER M2 ;
        RECT 0.56 14.447 2.96 14.449 ;
  LAYER M2 ;
        RECT 0.56 14.363 2.96 14.365 ;
  LAYER M2 ;
        RECT 0.56 14.279 2.96 14.281 ;
  LAYER M2 ;
        RECT 0.56 14.195 2.96 14.197 ;
  LAYER M2 ;
        RECT 0.56 14.111 2.96 14.113 ;
  LAYER M2 ;
        RECT 0.56 14.027 2.96 14.029 ;
  LAYER M2 ;
        RECT 0.56 13.943 2.96 13.945 ;
  LAYER M2 ;
        RECT 0.56 13.859 2.96 13.861 ;
  LAYER M1 ;
        RECT 2.944 10.8 2.976 13.308 ;
  LAYER M1 ;
        RECT 2.88 10.8 2.912 13.308 ;
  LAYER M1 ;
        RECT 2.816 10.8 2.848 13.308 ;
  LAYER M1 ;
        RECT 2.752 10.8 2.784 13.308 ;
  LAYER M1 ;
        RECT 2.688 10.8 2.72 13.308 ;
  LAYER M1 ;
        RECT 2.624 10.8 2.656 13.308 ;
  LAYER M1 ;
        RECT 2.56 10.8 2.592 13.308 ;
  LAYER M1 ;
        RECT 2.496 10.8 2.528 13.308 ;
  LAYER M1 ;
        RECT 2.432 10.8 2.464 13.308 ;
  LAYER M1 ;
        RECT 2.368 10.8 2.4 13.308 ;
  LAYER M1 ;
        RECT 2.304 10.8 2.336 13.308 ;
  LAYER M1 ;
        RECT 2.24 10.8 2.272 13.308 ;
  LAYER M1 ;
        RECT 2.176 10.8 2.208 13.308 ;
  LAYER M1 ;
        RECT 2.112 10.8 2.144 13.308 ;
  LAYER M1 ;
        RECT 2.048 10.8 2.08 13.308 ;
  LAYER M1 ;
        RECT 1.984 10.8 2.016 13.308 ;
  LAYER M1 ;
        RECT 1.92 10.8 1.952 13.308 ;
  LAYER M1 ;
        RECT 1.856 10.8 1.888 13.308 ;
  LAYER M1 ;
        RECT 1.792 10.8 1.824 13.308 ;
  LAYER M1 ;
        RECT 1.728 10.8 1.76 13.308 ;
  LAYER M1 ;
        RECT 1.664 10.8 1.696 13.308 ;
  LAYER M1 ;
        RECT 1.6 10.8 1.632 13.308 ;
  LAYER M1 ;
        RECT 1.536 10.8 1.568 13.308 ;
  LAYER M1 ;
        RECT 1.472 10.8 1.504 13.308 ;
  LAYER M1 ;
        RECT 1.408 10.8 1.44 13.308 ;
  LAYER M1 ;
        RECT 1.344 10.8 1.376 13.308 ;
  LAYER M1 ;
        RECT 1.28 10.8 1.312 13.308 ;
  LAYER M1 ;
        RECT 1.216 10.8 1.248 13.308 ;
  LAYER M1 ;
        RECT 1.152 10.8 1.184 13.308 ;
  LAYER M1 ;
        RECT 1.088 10.8 1.12 13.308 ;
  LAYER M1 ;
        RECT 1.024 10.8 1.056 13.308 ;
  LAYER M1 ;
        RECT 0.96 10.8 0.992 13.308 ;
  LAYER M1 ;
        RECT 0.896 10.8 0.928 13.308 ;
  LAYER M1 ;
        RECT 0.832 10.8 0.864 13.308 ;
  LAYER M1 ;
        RECT 0.768 10.8 0.8 13.308 ;
  LAYER M1 ;
        RECT 0.704 10.8 0.736 13.308 ;
  LAYER M1 ;
        RECT 0.64 10.8 0.672 13.308 ;
  LAYER M2 ;
        RECT 0.524 13.192 2.996 13.224 ;
  LAYER M2 ;
        RECT 0.524 13.128 2.996 13.16 ;
  LAYER M2 ;
        RECT 0.524 13.064 2.996 13.096 ;
  LAYER M2 ;
        RECT 0.524 13 2.996 13.032 ;
  LAYER M2 ;
        RECT 0.524 12.936 2.996 12.968 ;
  LAYER M2 ;
        RECT 0.524 12.872 2.996 12.904 ;
  LAYER M2 ;
        RECT 0.524 12.808 2.996 12.84 ;
  LAYER M2 ;
        RECT 0.524 12.744 2.996 12.776 ;
  LAYER M2 ;
        RECT 0.524 12.68 2.996 12.712 ;
  LAYER M2 ;
        RECT 0.524 12.616 2.996 12.648 ;
  LAYER M2 ;
        RECT 0.524 12.552 2.996 12.584 ;
  LAYER M2 ;
        RECT 0.524 12.488 2.996 12.52 ;
  LAYER M2 ;
        RECT 0.524 12.424 2.996 12.456 ;
  LAYER M2 ;
        RECT 0.524 12.36 2.996 12.392 ;
  LAYER M2 ;
        RECT 0.524 12.296 2.996 12.328 ;
  LAYER M2 ;
        RECT 0.524 12.232 2.996 12.264 ;
  LAYER M2 ;
        RECT 0.524 12.168 2.996 12.2 ;
  LAYER M2 ;
        RECT 0.524 12.104 2.996 12.136 ;
  LAYER M2 ;
        RECT 0.524 12.04 2.996 12.072 ;
  LAYER M2 ;
        RECT 0.524 11.976 2.996 12.008 ;
  LAYER M2 ;
        RECT 0.524 11.912 2.996 11.944 ;
  LAYER M2 ;
        RECT 0.524 11.848 2.996 11.88 ;
  LAYER M2 ;
        RECT 0.524 11.784 2.996 11.816 ;
  LAYER M2 ;
        RECT 0.524 11.72 2.996 11.752 ;
  LAYER M2 ;
        RECT 0.524 11.656 2.996 11.688 ;
  LAYER M2 ;
        RECT 0.524 11.592 2.996 11.624 ;
  LAYER M2 ;
        RECT 0.524 11.528 2.996 11.56 ;
  LAYER M2 ;
        RECT 0.524 11.464 2.996 11.496 ;
  LAYER M2 ;
        RECT 0.524 11.4 2.996 11.432 ;
  LAYER M2 ;
        RECT 0.524 11.336 2.996 11.368 ;
  LAYER M2 ;
        RECT 0.524 11.272 2.996 11.304 ;
  LAYER M2 ;
        RECT 0.524 11.208 2.996 11.24 ;
  LAYER M2 ;
        RECT 0.524 11.144 2.996 11.176 ;
  LAYER M2 ;
        RECT 0.524 11.08 2.996 11.112 ;
  LAYER M2 ;
        RECT 0.524 11.016 2.996 11.048 ;
  LAYER M2 ;
        RECT 0.524 10.952 2.996 10.984 ;
  LAYER M3 ;
        RECT 2.944 10.8 2.976 13.308 ;
  LAYER M3 ;
        RECT 2.88 10.8 2.912 13.308 ;
  LAYER M3 ;
        RECT 2.816 10.8 2.848 13.308 ;
  LAYER M3 ;
        RECT 2.752 10.8 2.784 13.308 ;
  LAYER M3 ;
        RECT 2.688 10.8 2.72 13.308 ;
  LAYER M3 ;
        RECT 2.624 10.8 2.656 13.308 ;
  LAYER M3 ;
        RECT 2.56 10.8 2.592 13.308 ;
  LAYER M3 ;
        RECT 2.496 10.8 2.528 13.308 ;
  LAYER M3 ;
        RECT 2.432 10.8 2.464 13.308 ;
  LAYER M3 ;
        RECT 2.368 10.8 2.4 13.308 ;
  LAYER M3 ;
        RECT 2.304 10.8 2.336 13.308 ;
  LAYER M3 ;
        RECT 2.24 10.8 2.272 13.308 ;
  LAYER M3 ;
        RECT 2.176 10.8 2.208 13.308 ;
  LAYER M3 ;
        RECT 2.112 10.8 2.144 13.308 ;
  LAYER M3 ;
        RECT 2.048 10.8 2.08 13.308 ;
  LAYER M3 ;
        RECT 1.984 10.8 2.016 13.308 ;
  LAYER M3 ;
        RECT 1.92 10.8 1.952 13.308 ;
  LAYER M3 ;
        RECT 1.856 10.8 1.888 13.308 ;
  LAYER M3 ;
        RECT 1.792 10.8 1.824 13.308 ;
  LAYER M3 ;
        RECT 1.728 10.8 1.76 13.308 ;
  LAYER M3 ;
        RECT 1.664 10.8 1.696 13.308 ;
  LAYER M3 ;
        RECT 1.6 10.8 1.632 13.308 ;
  LAYER M3 ;
        RECT 1.536 10.8 1.568 13.308 ;
  LAYER M3 ;
        RECT 1.472 10.8 1.504 13.308 ;
  LAYER M3 ;
        RECT 1.408 10.8 1.44 13.308 ;
  LAYER M3 ;
        RECT 1.344 10.8 1.376 13.308 ;
  LAYER M3 ;
        RECT 1.28 10.8 1.312 13.308 ;
  LAYER M3 ;
        RECT 1.216 10.8 1.248 13.308 ;
  LAYER M3 ;
        RECT 1.152 10.8 1.184 13.308 ;
  LAYER M3 ;
        RECT 1.088 10.8 1.12 13.308 ;
  LAYER M3 ;
        RECT 1.024 10.8 1.056 13.308 ;
  LAYER M3 ;
        RECT 0.96 10.8 0.992 13.308 ;
  LAYER M3 ;
        RECT 0.896 10.8 0.928 13.308 ;
  LAYER M3 ;
        RECT 0.832 10.8 0.864 13.308 ;
  LAYER M3 ;
        RECT 0.768 10.8 0.8 13.308 ;
  LAYER M3 ;
        RECT 0.704 10.8 0.736 13.308 ;
  LAYER M3 ;
        RECT 0.64 10.8 0.672 13.308 ;
  LAYER M3 ;
        RECT 0.544 10.8 0.576 13.308 ;
  LAYER M1 ;
        RECT 2.959 10.836 2.961 13.272 ;
  LAYER M1 ;
        RECT 2.879 10.836 2.881 13.272 ;
  LAYER M1 ;
        RECT 2.799 10.836 2.801 13.272 ;
  LAYER M1 ;
        RECT 2.719 10.836 2.721 13.272 ;
  LAYER M1 ;
        RECT 2.639 10.836 2.641 13.272 ;
  LAYER M1 ;
        RECT 2.559 10.836 2.561 13.272 ;
  LAYER M1 ;
        RECT 2.479 10.836 2.481 13.272 ;
  LAYER M1 ;
        RECT 2.399 10.836 2.401 13.272 ;
  LAYER M1 ;
        RECT 2.319 10.836 2.321 13.272 ;
  LAYER M1 ;
        RECT 2.239 10.836 2.241 13.272 ;
  LAYER M1 ;
        RECT 2.159 10.836 2.161 13.272 ;
  LAYER M1 ;
        RECT 2.079 10.836 2.081 13.272 ;
  LAYER M1 ;
        RECT 1.999 10.836 2.001 13.272 ;
  LAYER M1 ;
        RECT 1.919 10.836 1.921 13.272 ;
  LAYER M1 ;
        RECT 1.839 10.836 1.841 13.272 ;
  LAYER M1 ;
        RECT 1.759 10.836 1.761 13.272 ;
  LAYER M1 ;
        RECT 1.679 10.836 1.681 13.272 ;
  LAYER M1 ;
        RECT 1.599 10.836 1.601 13.272 ;
  LAYER M1 ;
        RECT 1.519 10.836 1.521 13.272 ;
  LAYER M1 ;
        RECT 1.439 10.836 1.441 13.272 ;
  LAYER M1 ;
        RECT 1.359 10.836 1.361 13.272 ;
  LAYER M1 ;
        RECT 1.279 10.836 1.281 13.272 ;
  LAYER M1 ;
        RECT 1.199 10.836 1.201 13.272 ;
  LAYER M1 ;
        RECT 1.119 10.836 1.121 13.272 ;
  LAYER M1 ;
        RECT 1.039 10.836 1.041 13.272 ;
  LAYER M1 ;
        RECT 0.959 10.836 0.961 13.272 ;
  LAYER M1 ;
        RECT 0.879 10.836 0.881 13.272 ;
  LAYER M1 ;
        RECT 0.799 10.836 0.801 13.272 ;
  LAYER M1 ;
        RECT 0.719 10.836 0.721 13.272 ;
  LAYER M1 ;
        RECT 0.639 10.836 0.641 13.272 ;
  LAYER M2 ;
        RECT 0.56 13.271 2.96 13.273 ;
  LAYER M2 ;
        RECT 0.56 13.187 2.96 13.189 ;
  LAYER M2 ;
        RECT 0.56 13.103 2.96 13.105 ;
  LAYER M2 ;
        RECT 0.56 13.019 2.96 13.021 ;
  LAYER M2 ;
        RECT 0.56 12.935 2.96 12.937 ;
  LAYER M2 ;
        RECT 0.56 12.851 2.96 12.853 ;
  LAYER M2 ;
        RECT 0.56 12.767 2.96 12.769 ;
  LAYER M2 ;
        RECT 0.56 12.683 2.96 12.685 ;
  LAYER M2 ;
        RECT 0.56 12.599 2.96 12.601 ;
  LAYER M2 ;
        RECT 0.56 12.515 2.96 12.517 ;
  LAYER M2 ;
        RECT 0.56 12.431 2.96 12.433 ;
  LAYER M2 ;
        RECT 0.56 12.347 2.96 12.349 ;
  LAYER M2 ;
        RECT 0.56 12.2635 2.96 12.2655 ;
  LAYER M2 ;
        RECT 0.56 12.179 2.96 12.181 ;
  LAYER M2 ;
        RECT 0.56 12.095 2.96 12.097 ;
  LAYER M2 ;
        RECT 0.56 12.011 2.96 12.013 ;
  LAYER M2 ;
        RECT 0.56 11.927 2.96 11.929 ;
  LAYER M2 ;
        RECT 0.56 11.843 2.96 11.845 ;
  LAYER M2 ;
        RECT 0.56 11.759 2.96 11.761 ;
  LAYER M2 ;
        RECT 0.56 11.675 2.96 11.677 ;
  LAYER M2 ;
        RECT 0.56 11.591 2.96 11.593 ;
  LAYER M2 ;
        RECT 0.56 11.507 2.96 11.509 ;
  LAYER M2 ;
        RECT 0.56 11.423 2.96 11.425 ;
  LAYER M2 ;
        RECT 0.56 11.339 2.96 11.341 ;
  LAYER M2 ;
        RECT 0.56 11.255 2.96 11.257 ;
  LAYER M2 ;
        RECT 0.56 11.171 2.96 11.173 ;
  LAYER M2 ;
        RECT 0.56 11.087 2.96 11.089 ;
  LAYER M2 ;
        RECT 0.56 11.003 2.96 11.005 ;
  LAYER M2 ;
        RECT 0.56 10.919 2.96 10.921 ;
  LAYER M1 ;
        RECT 2.944 7.86 2.976 10.368 ;
  LAYER M1 ;
        RECT 2.88 7.86 2.912 10.368 ;
  LAYER M1 ;
        RECT 2.816 7.86 2.848 10.368 ;
  LAYER M1 ;
        RECT 2.752 7.86 2.784 10.368 ;
  LAYER M1 ;
        RECT 2.688 7.86 2.72 10.368 ;
  LAYER M1 ;
        RECT 2.624 7.86 2.656 10.368 ;
  LAYER M1 ;
        RECT 2.56 7.86 2.592 10.368 ;
  LAYER M1 ;
        RECT 2.496 7.86 2.528 10.368 ;
  LAYER M1 ;
        RECT 2.432 7.86 2.464 10.368 ;
  LAYER M1 ;
        RECT 2.368 7.86 2.4 10.368 ;
  LAYER M1 ;
        RECT 2.304 7.86 2.336 10.368 ;
  LAYER M1 ;
        RECT 2.24 7.86 2.272 10.368 ;
  LAYER M1 ;
        RECT 2.176 7.86 2.208 10.368 ;
  LAYER M1 ;
        RECT 2.112 7.86 2.144 10.368 ;
  LAYER M1 ;
        RECT 2.048 7.86 2.08 10.368 ;
  LAYER M1 ;
        RECT 1.984 7.86 2.016 10.368 ;
  LAYER M1 ;
        RECT 1.92 7.86 1.952 10.368 ;
  LAYER M1 ;
        RECT 1.856 7.86 1.888 10.368 ;
  LAYER M1 ;
        RECT 1.792 7.86 1.824 10.368 ;
  LAYER M1 ;
        RECT 1.728 7.86 1.76 10.368 ;
  LAYER M1 ;
        RECT 1.664 7.86 1.696 10.368 ;
  LAYER M1 ;
        RECT 1.6 7.86 1.632 10.368 ;
  LAYER M1 ;
        RECT 1.536 7.86 1.568 10.368 ;
  LAYER M1 ;
        RECT 1.472 7.86 1.504 10.368 ;
  LAYER M1 ;
        RECT 1.408 7.86 1.44 10.368 ;
  LAYER M1 ;
        RECT 1.344 7.86 1.376 10.368 ;
  LAYER M1 ;
        RECT 1.28 7.86 1.312 10.368 ;
  LAYER M1 ;
        RECT 1.216 7.86 1.248 10.368 ;
  LAYER M1 ;
        RECT 1.152 7.86 1.184 10.368 ;
  LAYER M1 ;
        RECT 1.088 7.86 1.12 10.368 ;
  LAYER M1 ;
        RECT 1.024 7.86 1.056 10.368 ;
  LAYER M1 ;
        RECT 0.96 7.86 0.992 10.368 ;
  LAYER M1 ;
        RECT 0.896 7.86 0.928 10.368 ;
  LAYER M1 ;
        RECT 0.832 7.86 0.864 10.368 ;
  LAYER M1 ;
        RECT 0.768 7.86 0.8 10.368 ;
  LAYER M1 ;
        RECT 0.704 7.86 0.736 10.368 ;
  LAYER M1 ;
        RECT 0.64 7.86 0.672 10.368 ;
  LAYER M2 ;
        RECT 0.524 10.252 2.996 10.284 ;
  LAYER M2 ;
        RECT 0.524 10.188 2.996 10.22 ;
  LAYER M2 ;
        RECT 0.524 10.124 2.996 10.156 ;
  LAYER M2 ;
        RECT 0.524 10.06 2.996 10.092 ;
  LAYER M2 ;
        RECT 0.524 9.996 2.996 10.028 ;
  LAYER M2 ;
        RECT 0.524 9.932 2.996 9.964 ;
  LAYER M2 ;
        RECT 0.524 9.868 2.996 9.9 ;
  LAYER M2 ;
        RECT 0.524 9.804 2.996 9.836 ;
  LAYER M2 ;
        RECT 0.524 9.74 2.996 9.772 ;
  LAYER M2 ;
        RECT 0.524 9.676 2.996 9.708 ;
  LAYER M2 ;
        RECT 0.524 9.612 2.996 9.644 ;
  LAYER M2 ;
        RECT 0.524 9.548 2.996 9.58 ;
  LAYER M2 ;
        RECT 0.524 9.484 2.996 9.516 ;
  LAYER M2 ;
        RECT 0.524 9.42 2.996 9.452 ;
  LAYER M2 ;
        RECT 0.524 9.356 2.996 9.388 ;
  LAYER M2 ;
        RECT 0.524 9.292 2.996 9.324 ;
  LAYER M2 ;
        RECT 0.524 9.228 2.996 9.26 ;
  LAYER M2 ;
        RECT 0.524 9.164 2.996 9.196 ;
  LAYER M2 ;
        RECT 0.524 9.1 2.996 9.132 ;
  LAYER M2 ;
        RECT 0.524 9.036 2.996 9.068 ;
  LAYER M2 ;
        RECT 0.524 8.972 2.996 9.004 ;
  LAYER M2 ;
        RECT 0.524 8.908 2.996 8.94 ;
  LAYER M2 ;
        RECT 0.524 8.844 2.996 8.876 ;
  LAYER M2 ;
        RECT 0.524 8.78 2.996 8.812 ;
  LAYER M2 ;
        RECT 0.524 8.716 2.996 8.748 ;
  LAYER M2 ;
        RECT 0.524 8.652 2.996 8.684 ;
  LAYER M2 ;
        RECT 0.524 8.588 2.996 8.62 ;
  LAYER M2 ;
        RECT 0.524 8.524 2.996 8.556 ;
  LAYER M2 ;
        RECT 0.524 8.46 2.996 8.492 ;
  LAYER M2 ;
        RECT 0.524 8.396 2.996 8.428 ;
  LAYER M2 ;
        RECT 0.524 8.332 2.996 8.364 ;
  LAYER M2 ;
        RECT 0.524 8.268 2.996 8.3 ;
  LAYER M2 ;
        RECT 0.524 8.204 2.996 8.236 ;
  LAYER M2 ;
        RECT 0.524 8.14 2.996 8.172 ;
  LAYER M2 ;
        RECT 0.524 8.076 2.996 8.108 ;
  LAYER M2 ;
        RECT 0.524 8.012 2.996 8.044 ;
  LAYER M3 ;
        RECT 2.944 7.86 2.976 10.368 ;
  LAYER M3 ;
        RECT 2.88 7.86 2.912 10.368 ;
  LAYER M3 ;
        RECT 2.816 7.86 2.848 10.368 ;
  LAYER M3 ;
        RECT 2.752 7.86 2.784 10.368 ;
  LAYER M3 ;
        RECT 2.688 7.86 2.72 10.368 ;
  LAYER M3 ;
        RECT 2.624 7.86 2.656 10.368 ;
  LAYER M3 ;
        RECT 2.56 7.86 2.592 10.368 ;
  LAYER M3 ;
        RECT 2.496 7.86 2.528 10.368 ;
  LAYER M3 ;
        RECT 2.432 7.86 2.464 10.368 ;
  LAYER M3 ;
        RECT 2.368 7.86 2.4 10.368 ;
  LAYER M3 ;
        RECT 2.304 7.86 2.336 10.368 ;
  LAYER M3 ;
        RECT 2.24 7.86 2.272 10.368 ;
  LAYER M3 ;
        RECT 2.176 7.86 2.208 10.368 ;
  LAYER M3 ;
        RECT 2.112 7.86 2.144 10.368 ;
  LAYER M3 ;
        RECT 2.048 7.86 2.08 10.368 ;
  LAYER M3 ;
        RECT 1.984 7.86 2.016 10.368 ;
  LAYER M3 ;
        RECT 1.92 7.86 1.952 10.368 ;
  LAYER M3 ;
        RECT 1.856 7.86 1.888 10.368 ;
  LAYER M3 ;
        RECT 1.792 7.86 1.824 10.368 ;
  LAYER M3 ;
        RECT 1.728 7.86 1.76 10.368 ;
  LAYER M3 ;
        RECT 1.664 7.86 1.696 10.368 ;
  LAYER M3 ;
        RECT 1.6 7.86 1.632 10.368 ;
  LAYER M3 ;
        RECT 1.536 7.86 1.568 10.368 ;
  LAYER M3 ;
        RECT 1.472 7.86 1.504 10.368 ;
  LAYER M3 ;
        RECT 1.408 7.86 1.44 10.368 ;
  LAYER M3 ;
        RECT 1.344 7.86 1.376 10.368 ;
  LAYER M3 ;
        RECT 1.28 7.86 1.312 10.368 ;
  LAYER M3 ;
        RECT 1.216 7.86 1.248 10.368 ;
  LAYER M3 ;
        RECT 1.152 7.86 1.184 10.368 ;
  LAYER M3 ;
        RECT 1.088 7.86 1.12 10.368 ;
  LAYER M3 ;
        RECT 1.024 7.86 1.056 10.368 ;
  LAYER M3 ;
        RECT 0.96 7.86 0.992 10.368 ;
  LAYER M3 ;
        RECT 0.896 7.86 0.928 10.368 ;
  LAYER M3 ;
        RECT 0.832 7.86 0.864 10.368 ;
  LAYER M3 ;
        RECT 0.768 7.86 0.8 10.368 ;
  LAYER M3 ;
        RECT 0.704 7.86 0.736 10.368 ;
  LAYER M3 ;
        RECT 0.64 7.86 0.672 10.368 ;
  LAYER M3 ;
        RECT 0.544 7.86 0.576 10.368 ;
  LAYER M1 ;
        RECT 2.959 7.896 2.961 10.332 ;
  LAYER M1 ;
        RECT 2.879 7.896 2.881 10.332 ;
  LAYER M1 ;
        RECT 2.799 7.896 2.801 10.332 ;
  LAYER M1 ;
        RECT 2.719 7.896 2.721 10.332 ;
  LAYER M1 ;
        RECT 2.639 7.896 2.641 10.332 ;
  LAYER M1 ;
        RECT 2.559 7.896 2.561 10.332 ;
  LAYER M1 ;
        RECT 2.479 7.896 2.481 10.332 ;
  LAYER M1 ;
        RECT 2.399 7.896 2.401 10.332 ;
  LAYER M1 ;
        RECT 2.319 7.896 2.321 10.332 ;
  LAYER M1 ;
        RECT 2.239 7.896 2.241 10.332 ;
  LAYER M1 ;
        RECT 2.159 7.896 2.161 10.332 ;
  LAYER M1 ;
        RECT 2.079 7.896 2.081 10.332 ;
  LAYER M1 ;
        RECT 1.999 7.896 2.001 10.332 ;
  LAYER M1 ;
        RECT 1.919 7.896 1.921 10.332 ;
  LAYER M1 ;
        RECT 1.839 7.896 1.841 10.332 ;
  LAYER M1 ;
        RECT 1.759 7.896 1.761 10.332 ;
  LAYER M1 ;
        RECT 1.679 7.896 1.681 10.332 ;
  LAYER M1 ;
        RECT 1.599 7.896 1.601 10.332 ;
  LAYER M1 ;
        RECT 1.519 7.896 1.521 10.332 ;
  LAYER M1 ;
        RECT 1.439 7.896 1.441 10.332 ;
  LAYER M1 ;
        RECT 1.359 7.896 1.361 10.332 ;
  LAYER M1 ;
        RECT 1.279 7.896 1.281 10.332 ;
  LAYER M1 ;
        RECT 1.199 7.896 1.201 10.332 ;
  LAYER M1 ;
        RECT 1.119 7.896 1.121 10.332 ;
  LAYER M1 ;
        RECT 1.039 7.896 1.041 10.332 ;
  LAYER M1 ;
        RECT 0.959 7.896 0.961 10.332 ;
  LAYER M1 ;
        RECT 0.879 7.896 0.881 10.332 ;
  LAYER M1 ;
        RECT 0.799 7.896 0.801 10.332 ;
  LAYER M1 ;
        RECT 0.719 7.896 0.721 10.332 ;
  LAYER M1 ;
        RECT 0.639 7.896 0.641 10.332 ;
  LAYER M2 ;
        RECT 0.56 10.331 2.96 10.333 ;
  LAYER M2 ;
        RECT 0.56 10.247 2.96 10.249 ;
  LAYER M2 ;
        RECT 0.56 10.163 2.96 10.165 ;
  LAYER M2 ;
        RECT 0.56 10.079 2.96 10.081 ;
  LAYER M2 ;
        RECT 0.56 9.995 2.96 9.997 ;
  LAYER M2 ;
        RECT 0.56 9.911 2.96 9.913 ;
  LAYER M2 ;
        RECT 0.56 9.827 2.96 9.829 ;
  LAYER M2 ;
        RECT 0.56 9.743 2.96 9.745 ;
  LAYER M2 ;
        RECT 0.56 9.659 2.96 9.661 ;
  LAYER M2 ;
        RECT 0.56 9.575 2.96 9.577 ;
  LAYER M2 ;
        RECT 0.56 9.491 2.96 9.493 ;
  LAYER M2 ;
        RECT 0.56 9.407 2.96 9.409 ;
  LAYER M2 ;
        RECT 0.56 9.3235 2.96 9.3255 ;
  LAYER M2 ;
        RECT 0.56 9.239 2.96 9.241 ;
  LAYER M2 ;
        RECT 0.56 9.155 2.96 9.157 ;
  LAYER M2 ;
        RECT 0.56 9.071 2.96 9.073 ;
  LAYER M2 ;
        RECT 0.56 8.987 2.96 8.989 ;
  LAYER M2 ;
        RECT 0.56 8.903 2.96 8.905 ;
  LAYER M2 ;
        RECT 0.56 8.819 2.96 8.821 ;
  LAYER M2 ;
        RECT 0.56 8.735 2.96 8.737 ;
  LAYER M2 ;
        RECT 0.56 8.651 2.96 8.653 ;
  LAYER M2 ;
        RECT 0.56 8.567 2.96 8.569 ;
  LAYER M2 ;
        RECT 0.56 8.483 2.96 8.485 ;
  LAYER M2 ;
        RECT 0.56 8.399 2.96 8.401 ;
  LAYER M2 ;
        RECT 0.56 8.315 2.96 8.317 ;
  LAYER M2 ;
        RECT 0.56 8.231 2.96 8.233 ;
  LAYER M2 ;
        RECT 0.56 8.147 2.96 8.149 ;
  LAYER M2 ;
        RECT 0.56 8.063 2.96 8.065 ;
  LAYER M2 ;
        RECT 0.56 7.979 2.96 7.981 ;
  LAYER M1 ;
        RECT 2.944 4.92 2.976 7.428 ;
  LAYER M1 ;
        RECT 2.88 4.92 2.912 7.428 ;
  LAYER M1 ;
        RECT 2.816 4.92 2.848 7.428 ;
  LAYER M1 ;
        RECT 2.752 4.92 2.784 7.428 ;
  LAYER M1 ;
        RECT 2.688 4.92 2.72 7.428 ;
  LAYER M1 ;
        RECT 2.624 4.92 2.656 7.428 ;
  LAYER M1 ;
        RECT 2.56 4.92 2.592 7.428 ;
  LAYER M1 ;
        RECT 2.496 4.92 2.528 7.428 ;
  LAYER M1 ;
        RECT 2.432 4.92 2.464 7.428 ;
  LAYER M1 ;
        RECT 2.368 4.92 2.4 7.428 ;
  LAYER M1 ;
        RECT 2.304 4.92 2.336 7.428 ;
  LAYER M1 ;
        RECT 2.24 4.92 2.272 7.428 ;
  LAYER M1 ;
        RECT 2.176 4.92 2.208 7.428 ;
  LAYER M1 ;
        RECT 2.112 4.92 2.144 7.428 ;
  LAYER M1 ;
        RECT 2.048 4.92 2.08 7.428 ;
  LAYER M1 ;
        RECT 1.984 4.92 2.016 7.428 ;
  LAYER M1 ;
        RECT 1.92 4.92 1.952 7.428 ;
  LAYER M1 ;
        RECT 1.856 4.92 1.888 7.428 ;
  LAYER M1 ;
        RECT 1.792 4.92 1.824 7.428 ;
  LAYER M1 ;
        RECT 1.728 4.92 1.76 7.428 ;
  LAYER M1 ;
        RECT 1.664 4.92 1.696 7.428 ;
  LAYER M1 ;
        RECT 1.6 4.92 1.632 7.428 ;
  LAYER M1 ;
        RECT 1.536 4.92 1.568 7.428 ;
  LAYER M1 ;
        RECT 1.472 4.92 1.504 7.428 ;
  LAYER M1 ;
        RECT 1.408 4.92 1.44 7.428 ;
  LAYER M1 ;
        RECT 1.344 4.92 1.376 7.428 ;
  LAYER M1 ;
        RECT 1.28 4.92 1.312 7.428 ;
  LAYER M1 ;
        RECT 1.216 4.92 1.248 7.428 ;
  LAYER M1 ;
        RECT 1.152 4.92 1.184 7.428 ;
  LAYER M1 ;
        RECT 1.088 4.92 1.12 7.428 ;
  LAYER M1 ;
        RECT 1.024 4.92 1.056 7.428 ;
  LAYER M1 ;
        RECT 0.96 4.92 0.992 7.428 ;
  LAYER M1 ;
        RECT 0.896 4.92 0.928 7.428 ;
  LAYER M1 ;
        RECT 0.832 4.92 0.864 7.428 ;
  LAYER M1 ;
        RECT 0.768 4.92 0.8 7.428 ;
  LAYER M1 ;
        RECT 0.704 4.92 0.736 7.428 ;
  LAYER M1 ;
        RECT 0.64 4.92 0.672 7.428 ;
  LAYER M2 ;
        RECT 0.524 7.312 2.996 7.344 ;
  LAYER M2 ;
        RECT 0.524 7.248 2.996 7.28 ;
  LAYER M2 ;
        RECT 0.524 7.184 2.996 7.216 ;
  LAYER M2 ;
        RECT 0.524 7.12 2.996 7.152 ;
  LAYER M2 ;
        RECT 0.524 7.056 2.996 7.088 ;
  LAYER M2 ;
        RECT 0.524 6.992 2.996 7.024 ;
  LAYER M2 ;
        RECT 0.524 6.928 2.996 6.96 ;
  LAYER M2 ;
        RECT 0.524 6.864 2.996 6.896 ;
  LAYER M2 ;
        RECT 0.524 6.8 2.996 6.832 ;
  LAYER M2 ;
        RECT 0.524 6.736 2.996 6.768 ;
  LAYER M2 ;
        RECT 0.524 6.672 2.996 6.704 ;
  LAYER M2 ;
        RECT 0.524 6.608 2.996 6.64 ;
  LAYER M2 ;
        RECT 0.524 6.544 2.996 6.576 ;
  LAYER M2 ;
        RECT 0.524 6.48 2.996 6.512 ;
  LAYER M2 ;
        RECT 0.524 6.416 2.996 6.448 ;
  LAYER M2 ;
        RECT 0.524 6.352 2.996 6.384 ;
  LAYER M2 ;
        RECT 0.524 6.288 2.996 6.32 ;
  LAYER M2 ;
        RECT 0.524 6.224 2.996 6.256 ;
  LAYER M2 ;
        RECT 0.524 6.16 2.996 6.192 ;
  LAYER M2 ;
        RECT 0.524 6.096 2.996 6.128 ;
  LAYER M2 ;
        RECT 0.524 6.032 2.996 6.064 ;
  LAYER M2 ;
        RECT 0.524 5.968 2.996 6 ;
  LAYER M2 ;
        RECT 0.524 5.904 2.996 5.936 ;
  LAYER M2 ;
        RECT 0.524 5.84 2.996 5.872 ;
  LAYER M2 ;
        RECT 0.524 5.776 2.996 5.808 ;
  LAYER M2 ;
        RECT 0.524 5.712 2.996 5.744 ;
  LAYER M2 ;
        RECT 0.524 5.648 2.996 5.68 ;
  LAYER M2 ;
        RECT 0.524 5.584 2.996 5.616 ;
  LAYER M2 ;
        RECT 0.524 5.52 2.996 5.552 ;
  LAYER M2 ;
        RECT 0.524 5.456 2.996 5.488 ;
  LAYER M2 ;
        RECT 0.524 5.392 2.996 5.424 ;
  LAYER M2 ;
        RECT 0.524 5.328 2.996 5.36 ;
  LAYER M2 ;
        RECT 0.524 5.264 2.996 5.296 ;
  LAYER M2 ;
        RECT 0.524 5.2 2.996 5.232 ;
  LAYER M2 ;
        RECT 0.524 5.136 2.996 5.168 ;
  LAYER M2 ;
        RECT 0.524 5.072 2.996 5.104 ;
  LAYER M3 ;
        RECT 2.944 4.92 2.976 7.428 ;
  LAYER M3 ;
        RECT 2.88 4.92 2.912 7.428 ;
  LAYER M3 ;
        RECT 2.816 4.92 2.848 7.428 ;
  LAYER M3 ;
        RECT 2.752 4.92 2.784 7.428 ;
  LAYER M3 ;
        RECT 2.688 4.92 2.72 7.428 ;
  LAYER M3 ;
        RECT 2.624 4.92 2.656 7.428 ;
  LAYER M3 ;
        RECT 2.56 4.92 2.592 7.428 ;
  LAYER M3 ;
        RECT 2.496 4.92 2.528 7.428 ;
  LAYER M3 ;
        RECT 2.432 4.92 2.464 7.428 ;
  LAYER M3 ;
        RECT 2.368 4.92 2.4 7.428 ;
  LAYER M3 ;
        RECT 2.304 4.92 2.336 7.428 ;
  LAYER M3 ;
        RECT 2.24 4.92 2.272 7.428 ;
  LAYER M3 ;
        RECT 2.176 4.92 2.208 7.428 ;
  LAYER M3 ;
        RECT 2.112 4.92 2.144 7.428 ;
  LAYER M3 ;
        RECT 2.048 4.92 2.08 7.428 ;
  LAYER M3 ;
        RECT 1.984 4.92 2.016 7.428 ;
  LAYER M3 ;
        RECT 1.92 4.92 1.952 7.428 ;
  LAYER M3 ;
        RECT 1.856 4.92 1.888 7.428 ;
  LAYER M3 ;
        RECT 1.792 4.92 1.824 7.428 ;
  LAYER M3 ;
        RECT 1.728 4.92 1.76 7.428 ;
  LAYER M3 ;
        RECT 1.664 4.92 1.696 7.428 ;
  LAYER M3 ;
        RECT 1.6 4.92 1.632 7.428 ;
  LAYER M3 ;
        RECT 1.536 4.92 1.568 7.428 ;
  LAYER M3 ;
        RECT 1.472 4.92 1.504 7.428 ;
  LAYER M3 ;
        RECT 1.408 4.92 1.44 7.428 ;
  LAYER M3 ;
        RECT 1.344 4.92 1.376 7.428 ;
  LAYER M3 ;
        RECT 1.28 4.92 1.312 7.428 ;
  LAYER M3 ;
        RECT 1.216 4.92 1.248 7.428 ;
  LAYER M3 ;
        RECT 1.152 4.92 1.184 7.428 ;
  LAYER M3 ;
        RECT 1.088 4.92 1.12 7.428 ;
  LAYER M3 ;
        RECT 1.024 4.92 1.056 7.428 ;
  LAYER M3 ;
        RECT 0.96 4.92 0.992 7.428 ;
  LAYER M3 ;
        RECT 0.896 4.92 0.928 7.428 ;
  LAYER M3 ;
        RECT 0.832 4.92 0.864 7.428 ;
  LAYER M3 ;
        RECT 0.768 4.92 0.8 7.428 ;
  LAYER M3 ;
        RECT 0.704 4.92 0.736 7.428 ;
  LAYER M3 ;
        RECT 0.64 4.92 0.672 7.428 ;
  LAYER M3 ;
        RECT 0.544 4.92 0.576 7.428 ;
  LAYER M1 ;
        RECT 2.959 4.956 2.961 7.392 ;
  LAYER M1 ;
        RECT 2.879 4.956 2.881 7.392 ;
  LAYER M1 ;
        RECT 2.799 4.956 2.801 7.392 ;
  LAYER M1 ;
        RECT 2.719 4.956 2.721 7.392 ;
  LAYER M1 ;
        RECT 2.639 4.956 2.641 7.392 ;
  LAYER M1 ;
        RECT 2.559 4.956 2.561 7.392 ;
  LAYER M1 ;
        RECT 2.479 4.956 2.481 7.392 ;
  LAYER M1 ;
        RECT 2.399 4.956 2.401 7.392 ;
  LAYER M1 ;
        RECT 2.319 4.956 2.321 7.392 ;
  LAYER M1 ;
        RECT 2.239 4.956 2.241 7.392 ;
  LAYER M1 ;
        RECT 2.159 4.956 2.161 7.392 ;
  LAYER M1 ;
        RECT 2.079 4.956 2.081 7.392 ;
  LAYER M1 ;
        RECT 1.999 4.956 2.001 7.392 ;
  LAYER M1 ;
        RECT 1.919 4.956 1.921 7.392 ;
  LAYER M1 ;
        RECT 1.839 4.956 1.841 7.392 ;
  LAYER M1 ;
        RECT 1.759 4.956 1.761 7.392 ;
  LAYER M1 ;
        RECT 1.679 4.956 1.681 7.392 ;
  LAYER M1 ;
        RECT 1.599 4.956 1.601 7.392 ;
  LAYER M1 ;
        RECT 1.519 4.956 1.521 7.392 ;
  LAYER M1 ;
        RECT 1.439 4.956 1.441 7.392 ;
  LAYER M1 ;
        RECT 1.359 4.956 1.361 7.392 ;
  LAYER M1 ;
        RECT 1.279 4.956 1.281 7.392 ;
  LAYER M1 ;
        RECT 1.199 4.956 1.201 7.392 ;
  LAYER M1 ;
        RECT 1.119 4.956 1.121 7.392 ;
  LAYER M1 ;
        RECT 1.039 4.956 1.041 7.392 ;
  LAYER M1 ;
        RECT 0.959 4.956 0.961 7.392 ;
  LAYER M1 ;
        RECT 0.879 4.956 0.881 7.392 ;
  LAYER M1 ;
        RECT 0.799 4.956 0.801 7.392 ;
  LAYER M1 ;
        RECT 0.719 4.956 0.721 7.392 ;
  LAYER M1 ;
        RECT 0.639 4.956 0.641 7.392 ;
  LAYER M2 ;
        RECT 0.56 7.391 2.96 7.393 ;
  LAYER M2 ;
        RECT 0.56 7.307 2.96 7.309 ;
  LAYER M2 ;
        RECT 0.56 7.223 2.96 7.225 ;
  LAYER M2 ;
        RECT 0.56 7.139 2.96 7.141 ;
  LAYER M2 ;
        RECT 0.56 7.055 2.96 7.057 ;
  LAYER M2 ;
        RECT 0.56 6.971 2.96 6.973 ;
  LAYER M2 ;
        RECT 0.56 6.887 2.96 6.889 ;
  LAYER M2 ;
        RECT 0.56 6.803 2.96 6.805 ;
  LAYER M2 ;
        RECT 0.56 6.719 2.96 6.721 ;
  LAYER M2 ;
        RECT 0.56 6.635 2.96 6.637 ;
  LAYER M2 ;
        RECT 0.56 6.551 2.96 6.553 ;
  LAYER M2 ;
        RECT 0.56 6.467 2.96 6.469 ;
  LAYER M2 ;
        RECT 0.56 6.3835 2.96 6.3855 ;
  LAYER M2 ;
        RECT 0.56 6.299 2.96 6.301 ;
  LAYER M2 ;
        RECT 0.56 6.215 2.96 6.217 ;
  LAYER M2 ;
        RECT 0.56 6.131 2.96 6.133 ;
  LAYER M2 ;
        RECT 0.56 6.047 2.96 6.049 ;
  LAYER M2 ;
        RECT 0.56 5.963 2.96 5.965 ;
  LAYER M2 ;
        RECT 0.56 5.879 2.96 5.881 ;
  LAYER M2 ;
        RECT 0.56 5.795 2.96 5.797 ;
  LAYER M2 ;
        RECT 0.56 5.711 2.96 5.713 ;
  LAYER M2 ;
        RECT 0.56 5.627 2.96 5.629 ;
  LAYER M2 ;
        RECT 0.56 5.543 2.96 5.545 ;
  LAYER M2 ;
        RECT 0.56 5.459 2.96 5.461 ;
  LAYER M2 ;
        RECT 0.56 5.375 2.96 5.377 ;
  LAYER M2 ;
        RECT 0.56 5.291 2.96 5.293 ;
  LAYER M2 ;
        RECT 0.56 5.207 2.96 5.209 ;
  LAYER M2 ;
        RECT 0.56 5.123 2.96 5.125 ;
  LAYER M2 ;
        RECT 0.56 5.039 2.96 5.041 ;
  LAYER M1 ;
        RECT 2.944 1.98 2.976 4.488 ;
  LAYER M1 ;
        RECT 2.88 1.98 2.912 4.488 ;
  LAYER M1 ;
        RECT 2.816 1.98 2.848 4.488 ;
  LAYER M1 ;
        RECT 2.752 1.98 2.784 4.488 ;
  LAYER M1 ;
        RECT 2.688 1.98 2.72 4.488 ;
  LAYER M1 ;
        RECT 2.624 1.98 2.656 4.488 ;
  LAYER M1 ;
        RECT 2.56 1.98 2.592 4.488 ;
  LAYER M1 ;
        RECT 2.496 1.98 2.528 4.488 ;
  LAYER M1 ;
        RECT 2.432 1.98 2.464 4.488 ;
  LAYER M1 ;
        RECT 2.368 1.98 2.4 4.488 ;
  LAYER M1 ;
        RECT 2.304 1.98 2.336 4.488 ;
  LAYER M1 ;
        RECT 2.24 1.98 2.272 4.488 ;
  LAYER M1 ;
        RECT 2.176 1.98 2.208 4.488 ;
  LAYER M1 ;
        RECT 2.112 1.98 2.144 4.488 ;
  LAYER M1 ;
        RECT 2.048 1.98 2.08 4.488 ;
  LAYER M1 ;
        RECT 1.984 1.98 2.016 4.488 ;
  LAYER M1 ;
        RECT 1.92 1.98 1.952 4.488 ;
  LAYER M1 ;
        RECT 1.856 1.98 1.888 4.488 ;
  LAYER M1 ;
        RECT 1.792 1.98 1.824 4.488 ;
  LAYER M1 ;
        RECT 1.728 1.98 1.76 4.488 ;
  LAYER M1 ;
        RECT 1.664 1.98 1.696 4.488 ;
  LAYER M1 ;
        RECT 1.6 1.98 1.632 4.488 ;
  LAYER M1 ;
        RECT 1.536 1.98 1.568 4.488 ;
  LAYER M1 ;
        RECT 1.472 1.98 1.504 4.488 ;
  LAYER M1 ;
        RECT 1.408 1.98 1.44 4.488 ;
  LAYER M1 ;
        RECT 1.344 1.98 1.376 4.488 ;
  LAYER M1 ;
        RECT 1.28 1.98 1.312 4.488 ;
  LAYER M1 ;
        RECT 1.216 1.98 1.248 4.488 ;
  LAYER M1 ;
        RECT 1.152 1.98 1.184 4.488 ;
  LAYER M1 ;
        RECT 1.088 1.98 1.12 4.488 ;
  LAYER M1 ;
        RECT 1.024 1.98 1.056 4.488 ;
  LAYER M1 ;
        RECT 0.96 1.98 0.992 4.488 ;
  LAYER M1 ;
        RECT 0.896 1.98 0.928 4.488 ;
  LAYER M1 ;
        RECT 0.832 1.98 0.864 4.488 ;
  LAYER M1 ;
        RECT 0.768 1.98 0.8 4.488 ;
  LAYER M1 ;
        RECT 0.704 1.98 0.736 4.488 ;
  LAYER M1 ;
        RECT 0.64 1.98 0.672 4.488 ;
  LAYER M2 ;
        RECT 0.524 4.372 2.996 4.404 ;
  LAYER M2 ;
        RECT 0.524 4.308 2.996 4.34 ;
  LAYER M2 ;
        RECT 0.524 4.244 2.996 4.276 ;
  LAYER M2 ;
        RECT 0.524 4.18 2.996 4.212 ;
  LAYER M2 ;
        RECT 0.524 4.116 2.996 4.148 ;
  LAYER M2 ;
        RECT 0.524 4.052 2.996 4.084 ;
  LAYER M2 ;
        RECT 0.524 3.988 2.996 4.02 ;
  LAYER M2 ;
        RECT 0.524 3.924 2.996 3.956 ;
  LAYER M2 ;
        RECT 0.524 3.86 2.996 3.892 ;
  LAYER M2 ;
        RECT 0.524 3.796 2.996 3.828 ;
  LAYER M2 ;
        RECT 0.524 3.732 2.996 3.764 ;
  LAYER M2 ;
        RECT 0.524 3.668 2.996 3.7 ;
  LAYER M2 ;
        RECT 0.524 3.604 2.996 3.636 ;
  LAYER M2 ;
        RECT 0.524 3.54 2.996 3.572 ;
  LAYER M2 ;
        RECT 0.524 3.476 2.996 3.508 ;
  LAYER M2 ;
        RECT 0.524 3.412 2.996 3.444 ;
  LAYER M2 ;
        RECT 0.524 3.348 2.996 3.38 ;
  LAYER M2 ;
        RECT 0.524 3.284 2.996 3.316 ;
  LAYER M2 ;
        RECT 0.524 3.22 2.996 3.252 ;
  LAYER M2 ;
        RECT 0.524 3.156 2.996 3.188 ;
  LAYER M2 ;
        RECT 0.524 3.092 2.996 3.124 ;
  LAYER M2 ;
        RECT 0.524 3.028 2.996 3.06 ;
  LAYER M2 ;
        RECT 0.524 2.964 2.996 2.996 ;
  LAYER M2 ;
        RECT 0.524 2.9 2.996 2.932 ;
  LAYER M2 ;
        RECT 0.524 2.836 2.996 2.868 ;
  LAYER M2 ;
        RECT 0.524 2.772 2.996 2.804 ;
  LAYER M2 ;
        RECT 0.524 2.708 2.996 2.74 ;
  LAYER M2 ;
        RECT 0.524 2.644 2.996 2.676 ;
  LAYER M2 ;
        RECT 0.524 2.58 2.996 2.612 ;
  LAYER M2 ;
        RECT 0.524 2.516 2.996 2.548 ;
  LAYER M2 ;
        RECT 0.524 2.452 2.996 2.484 ;
  LAYER M2 ;
        RECT 0.524 2.388 2.996 2.42 ;
  LAYER M2 ;
        RECT 0.524 2.324 2.996 2.356 ;
  LAYER M2 ;
        RECT 0.524 2.26 2.996 2.292 ;
  LAYER M2 ;
        RECT 0.524 2.196 2.996 2.228 ;
  LAYER M2 ;
        RECT 0.524 2.132 2.996 2.164 ;
  LAYER M3 ;
        RECT 2.944 1.98 2.976 4.488 ;
  LAYER M3 ;
        RECT 2.88 1.98 2.912 4.488 ;
  LAYER M3 ;
        RECT 2.816 1.98 2.848 4.488 ;
  LAYER M3 ;
        RECT 2.752 1.98 2.784 4.488 ;
  LAYER M3 ;
        RECT 2.688 1.98 2.72 4.488 ;
  LAYER M3 ;
        RECT 2.624 1.98 2.656 4.488 ;
  LAYER M3 ;
        RECT 2.56 1.98 2.592 4.488 ;
  LAYER M3 ;
        RECT 2.496 1.98 2.528 4.488 ;
  LAYER M3 ;
        RECT 2.432 1.98 2.464 4.488 ;
  LAYER M3 ;
        RECT 2.368 1.98 2.4 4.488 ;
  LAYER M3 ;
        RECT 2.304 1.98 2.336 4.488 ;
  LAYER M3 ;
        RECT 2.24 1.98 2.272 4.488 ;
  LAYER M3 ;
        RECT 2.176 1.98 2.208 4.488 ;
  LAYER M3 ;
        RECT 2.112 1.98 2.144 4.488 ;
  LAYER M3 ;
        RECT 2.048 1.98 2.08 4.488 ;
  LAYER M3 ;
        RECT 1.984 1.98 2.016 4.488 ;
  LAYER M3 ;
        RECT 1.92 1.98 1.952 4.488 ;
  LAYER M3 ;
        RECT 1.856 1.98 1.888 4.488 ;
  LAYER M3 ;
        RECT 1.792 1.98 1.824 4.488 ;
  LAYER M3 ;
        RECT 1.728 1.98 1.76 4.488 ;
  LAYER M3 ;
        RECT 1.664 1.98 1.696 4.488 ;
  LAYER M3 ;
        RECT 1.6 1.98 1.632 4.488 ;
  LAYER M3 ;
        RECT 1.536 1.98 1.568 4.488 ;
  LAYER M3 ;
        RECT 1.472 1.98 1.504 4.488 ;
  LAYER M3 ;
        RECT 1.408 1.98 1.44 4.488 ;
  LAYER M3 ;
        RECT 1.344 1.98 1.376 4.488 ;
  LAYER M3 ;
        RECT 1.28 1.98 1.312 4.488 ;
  LAYER M3 ;
        RECT 1.216 1.98 1.248 4.488 ;
  LAYER M3 ;
        RECT 1.152 1.98 1.184 4.488 ;
  LAYER M3 ;
        RECT 1.088 1.98 1.12 4.488 ;
  LAYER M3 ;
        RECT 1.024 1.98 1.056 4.488 ;
  LAYER M3 ;
        RECT 0.96 1.98 0.992 4.488 ;
  LAYER M3 ;
        RECT 0.896 1.98 0.928 4.488 ;
  LAYER M3 ;
        RECT 0.832 1.98 0.864 4.488 ;
  LAYER M3 ;
        RECT 0.768 1.98 0.8 4.488 ;
  LAYER M3 ;
        RECT 0.704 1.98 0.736 4.488 ;
  LAYER M3 ;
        RECT 0.64 1.98 0.672 4.488 ;
  LAYER M3 ;
        RECT 0.544 1.98 0.576 4.488 ;
  LAYER M1 ;
        RECT 2.959 2.016 2.961 4.452 ;
  LAYER M1 ;
        RECT 2.879 2.016 2.881 4.452 ;
  LAYER M1 ;
        RECT 2.799 2.016 2.801 4.452 ;
  LAYER M1 ;
        RECT 2.719 2.016 2.721 4.452 ;
  LAYER M1 ;
        RECT 2.639 2.016 2.641 4.452 ;
  LAYER M1 ;
        RECT 2.559 2.016 2.561 4.452 ;
  LAYER M1 ;
        RECT 2.479 2.016 2.481 4.452 ;
  LAYER M1 ;
        RECT 2.399 2.016 2.401 4.452 ;
  LAYER M1 ;
        RECT 2.319 2.016 2.321 4.452 ;
  LAYER M1 ;
        RECT 2.239 2.016 2.241 4.452 ;
  LAYER M1 ;
        RECT 2.159 2.016 2.161 4.452 ;
  LAYER M1 ;
        RECT 2.079 2.016 2.081 4.452 ;
  LAYER M1 ;
        RECT 1.999 2.016 2.001 4.452 ;
  LAYER M1 ;
        RECT 1.919 2.016 1.921 4.452 ;
  LAYER M1 ;
        RECT 1.839 2.016 1.841 4.452 ;
  LAYER M1 ;
        RECT 1.759 2.016 1.761 4.452 ;
  LAYER M1 ;
        RECT 1.679 2.016 1.681 4.452 ;
  LAYER M1 ;
        RECT 1.599 2.016 1.601 4.452 ;
  LAYER M1 ;
        RECT 1.519 2.016 1.521 4.452 ;
  LAYER M1 ;
        RECT 1.439 2.016 1.441 4.452 ;
  LAYER M1 ;
        RECT 1.359 2.016 1.361 4.452 ;
  LAYER M1 ;
        RECT 1.279 2.016 1.281 4.452 ;
  LAYER M1 ;
        RECT 1.199 2.016 1.201 4.452 ;
  LAYER M1 ;
        RECT 1.119 2.016 1.121 4.452 ;
  LAYER M1 ;
        RECT 1.039 2.016 1.041 4.452 ;
  LAYER M1 ;
        RECT 0.959 2.016 0.961 4.452 ;
  LAYER M1 ;
        RECT 0.879 2.016 0.881 4.452 ;
  LAYER M1 ;
        RECT 0.799 2.016 0.801 4.452 ;
  LAYER M1 ;
        RECT 0.719 2.016 0.721 4.452 ;
  LAYER M1 ;
        RECT 0.639 2.016 0.641 4.452 ;
  LAYER M2 ;
        RECT 0.56 4.451 2.96 4.453 ;
  LAYER M2 ;
        RECT 0.56 4.367 2.96 4.369 ;
  LAYER M2 ;
        RECT 0.56 4.283 2.96 4.285 ;
  LAYER M2 ;
        RECT 0.56 4.199 2.96 4.201 ;
  LAYER M2 ;
        RECT 0.56 4.115 2.96 4.117 ;
  LAYER M2 ;
        RECT 0.56 4.031 2.96 4.033 ;
  LAYER M2 ;
        RECT 0.56 3.947 2.96 3.949 ;
  LAYER M2 ;
        RECT 0.56 3.863 2.96 3.865 ;
  LAYER M2 ;
        RECT 0.56 3.779 2.96 3.781 ;
  LAYER M2 ;
        RECT 0.56 3.695 2.96 3.697 ;
  LAYER M2 ;
        RECT 0.56 3.611 2.96 3.613 ;
  LAYER M2 ;
        RECT 0.56 3.527 2.96 3.529 ;
  LAYER M2 ;
        RECT 0.56 3.4435 2.96 3.4455 ;
  LAYER M2 ;
        RECT 0.56 3.359 2.96 3.361 ;
  LAYER M2 ;
        RECT 0.56 3.275 2.96 3.277 ;
  LAYER M2 ;
        RECT 0.56 3.191 2.96 3.193 ;
  LAYER M2 ;
        RECT 0.56 3.107 2.96 3.109 ;
  LAYER M2 ;
        RECT 0.56 3.023 2.96 3.025 ;
  LAYER M2 ;
        RECT 0.56 2.939 2.96 2.941 ;
  LAYER M2 ;
        RECT 0.56 2.855 2.96 2.857 ;
  LAYER M2 ;
        RECT 0.56 2.771 2.96 2.773 ;
  LAYER M2 ;
        RECT 0.56 2.687 2.96 2.689 ;
  LAYER M2 ;
        RECT 0.56 2.603 2.96 2.605 ;
  LAYER M2 ;
        RECT 0.56 2.519 2.96 2.521 ;
  LAYER M2 ;
        RECT 0.56 2.435 2.96 2.437 ;
  LAYER M2 ;
        RECT 0.56 2.351 2.96 2.353 ;
  LAYER M2 ;
        RECT 0.56 2.267 2.96 2.269 ;
  LAYER M2 ;
        RECT 0.56 2.183 2.96 2.185 ;
  LAYER M2 ;
        RECT 0.56 2.099 2.96 2.101 ;
  LAYER M1 ;
        RECT 39.824 29.7 39.856 29.772 ;
  LAYER M2 ;
        RECT 39.804 29.72 39.876 29.752 ;
  LAYER M1 ;
        RECT 36.944 29.7 36.976 29.772 ;
  LAYER M2 ;
        RECT 36.924 29.72 36.996 29.752 ;
  LAYER M2 ;
        RECT 36.96 29.72 39.84 29.752 ;
  LAYER M2 ;
        RECT 39.484 0.908 40.196 0.94 ;
  LAYER M1 ;
        RECT 37.024 16.68 37.056 16.752 ;
  LAYER M2 ;
        RECT 37.004 16.7 37.076 16.732 ;
  LAYER M1 ;
        RECT 39.904 16.68 39.936 16.752 ;
  LAYER M2 ;
        RECT 39.884 16.7 39.956 16.732 ;
  LAYER M2 ;
        RECT 37.04 16.7 39.92 16.732 ;
  LAYER M2 ;
        RECT 37.664 29.72 37.696 29.752 ;
  LAYER M3 ;
        RECT 37.66 29.484 37.7 29.736 ;
  LAYER M4 ;
        RECT 37.66 29.464 37.7 29.504 ;
  LAYER M5 ;
        RECT 37.648 16.968 37.712 29.484 ;
  LAYER M4 ;
        RECT 37.66 16.948 37.7 16.988 ;
  LAYER M3 ;
        RECT 37.66 16.716 37.7 16.968 ;
  LAYER M2 ;
        RECT 37.664 16.7 37.696 16.732 ;
  LAYER M2 ;
        RECT 39.824 16.7 39.856 16.732 ;
  LAYER M3 ;
        RECT 39.82 1.596 39.86 16.716 ;
  LAYER M4 ;
        RECT 39.82 1.576 39.86 1.616 ;
  LAYER M5 ;
        RECT 39.808 1.428 39.872 1.596 ;
  LAYER M4 ;
        RECT 39.82 1.408 39.86 1.448 ;
  LAYER M3 ;
        RECT 39.82 0.924 39.86 1.428 ;
  LAYER M2 ;
        RECT 39.824 0.908 39.856 0.94 ;
  LAYER M1 ;
        RECT 39.984 17.436 40.016 17.508 ;
  LAYER M2 ;
        RECT 39.964 17.456 40.036 17.488 ;
  LAYER M1 ;
        RECT 37.104 17.436 37.136 17.508 ;
  LAYER M2 ;
        RECT 37.084 17.456 37.156 17.488 ;
  LAYER M2 ;
        RECT 37.12 17.456 40 17.488 ;
  LAYER M3 ;
        RECT 41.02 0.552 41.06 0.876 ;
  LAYER M3 ;
        RECT 40.78 0.552 40.82 0.876 ;
  LAYER M3 ;
        RECT 30.94 17.604 30.98 17.928 ;
  LAYER M3 ;
        RECT 30.7 17.604 30.74 17.928 ;
  LAYER M2 ;
        RECT 30.96 17.456 37.2 17.488 ;
  LAYER M3 ;
        RECT 30.94 17.472 30.98 17.724 ;
  LAYER M2 ;
        RECT 39.984 17.456 40.016 17.488 ;
  LAYER M3 ;
        RECT 39.98 0.84 40.02 17.472 ;
  LAYER M4 ;
        RECT 40 0.82 40.8 0.86 ;
  LAYER M3 ;
        RECT 40.78 0.82 40.82 0.86 ;
  LAYER M2 ;
        RECT 38.284 0.908 38.996 0.94 ;
  LAYER M1 ;
        RECT 37.184 1.476 37.216 1.548 ;
  LAYER M2 ;
        RECT 37.164 1.496 37.236 1.528 ;
  LAYER M1 ;
        RECT 40.064 1.476 40.096 1.548 ;
  LAYER M2 ;
        RECT 40.044 1.496 40.116 1.528 ;
  LAYER M2 ;
        RECT 37.2 1.496 40.08 1.528 ;
  LAYER M2 ;
        RECT 38.384 0.908 38.416 0.94 ;
  LAYER M3 ;
        RECT 38.38 0.924 38.42 1.428 ;
  LAYER M4 ;
        RECT 38.38 1.408 38.42 1.448 ;
  LAYER M5 ;
        RECT 38.368 1.428 38.432 1.512 ;
  LAYER M4 ;
        RECT 38.38 1.492 38.42 1.532 ;
  LAYER M3 ;
        RECT 38.38 1.492 38.42 1.532 ;
  LAYER M2 ;
        RECT 38.384 1.496 38.416 1.528 ;
  LAYER M1 ;
        RECT 39.664 20.88 39.696 20.952 ;
  LAYER M2 ;
        RECT 39.644 20.9 39.716 20.932 ;
  LAYER M2 ;
        RECT 39.68 20.9 40 20.932 ;
  LAYER M1 ;
        RECT 39.984 20.88 40.016 20.952 ;
  LAYER M2 ;
        RECT 39.964 20.9 40.036 20.932 ;
  LAYER M1 ;
        RECT 39.664 23.82 39.696 23.892 ;
  LAYER M2 ;
        RECT 39.644 23.84 39.716 23.872 ;
  LAYER M2 ;
        RECT 39.68 23.84 40 23.872 ;
  LAYER M1 ;
        RECT 39.984 23.82 40.016 23.892 ;
  LAYER M2 ;
        RECT 39.964 23.84 40.036 23.872 ;
  LAYER M1 ;
        RECT 42.544 20.88 42.576 20.952 ;
  LAYER M2 ;
        RECT 42.524 20.9 42.596 20.932 ;
  LAYER M1 ;
        RECT 42.544 20.748 42.576 20.916 ;
  LAYER M1 ;
        RECT 42.544 20.712 42.576 20.784 ;
  LAYER M2 ;
        RECT 42.524 20.732 42.596 20.764 ;
  LAYER M2 ;
        RECT 40 20.732 42.56 20.764 ;
  LAYER M1 ;
        RECT 39.984 20.712 40.016 20.784 ;
  LAYER M2 ;
        RECT 39.964 20.732 40.036 20.764 ;
  LAYER M1 ;
        RECT 42.544 23.82 42.576 23.892 ;
  LAYER M2 ;
        RECT 42.524 23.84 42.596 23.872 ;
  LAYER M1 ;
        RECT 42.544 23.688 42.576 23.856 ;
  LAYER M1 ;
        RECT 42.544 23.652 42.576 23.724 ;
  LAYER M2 ;
        RECT 42.524 23.672 42.596 23.704 ;
  LAYER M2 ;
        RECT 40 23.672 42.56 23.704 ;
  LAYER M1 ;
        RECT 39.984 23.652 40.016 23.724 ;
  LAYER M2 ;
        RECT 39.964 23.672 40.036 23.704 ;
  LAYER M1 ;
        RECT 39.984 17.436 40.016 17.508 ;
  LAYER M2 ;
        RECT 39.964 17.456 40.036 17.488 ;
  LAYER M1 ;
        RECT 39.984 17.472 40.016 17.64 ;
  LAYER M1 ;
        RECT 39.984 17.64 40.016 23.856 ;
  LAYER M1 ;
        RECT 36.784 23.82 36.816 23.892 ;
  LAYER M2 ;
        RECT 36.764 23.84 36.836 23.872 ;
  LAYER M2 ;
        RECT 36.8 23.84 37.12 23.872 ;
  LAYER M1 ;
        RECT 37.104 23.82 37.136 23.892 ;
  LAYER M2 ;
        RECT 37.084 23.84 37.156 23.872 ;
  LAYER M1 ;
        RECT 36.784 20.88 36.816 20.952 ;
  LAYER M2 ;
        RECT 36.764 20.9 36.836 20.932 ;
  LAYER M2 ;
        RECT 36.8 20.9 37.12 20.932 ;
  LAYER M1 ;
        RECT 37.104 20.88 37.136 20.952 ;
  LAYER M2 ;
        RECT 37.084 20.9 37.156 20.932 ;
  LAYER M1 ;
        RECT 37.104 17.436 37.136 17.508 ;
  LAYER M2 ;
        RECT 37.084 17.456 37.156 17.488 ;
  LAYER M1 ;
        RECT 37.104 17.472 37.136 17.64 ;
  LAYER M1 ;
        RECT 37.104 17.64 37.136 23.856 ;
  LAYER M2 ;
        RECT 37.12 17.456 40 17.488 ;
  LAYER M1 ;
        RECT 45.424 17.94 45.456 18.012 ;
  LAYER M2 ;
        RECT 45.404 17.96 45.476 17.992 ;
  LAYER M1 ;
        RECT 45.424 17.808 45.456 17.976 ;
  LAYER M1 ;
        RECT 45.424 17.772 45.456 17.844 ;
  LAYER M2 ;
        RECT 45.404 17.792 45.476 17.824 ;
  LAYER M2 ;
        RECT 42.88 17.792 45.44 17.824 ;
  LAYER M1 ;
        RECT 42.864 17.772 42.896 17.844 ;
  LAYER M2 ;
        RECT 42.844 17.792 42.916 17.824 ;
  LAYER M1 ;
        RECT 45.424 20.88 45.456 20.952 ;
  LAYER M2 ;
        RECT 45.404 20.9 45.476 20.932 ;
  LAYER M1 ;
        RECT 45.424 20.748 45.456 20.916 ;
  LAYER M1 ;
        RECT 45.424 20.712 45.456 20.784 ;
  LAYER M2 ;
        RECT 45.404 20.732 45.476 20.764 ;
  LAYER M2 ;
        RECT 42.88 20.732 45.44 20.764 ;
  LAYER M1 ;
        RECT 42.864 20.712 42.896 20.784 ;
  LAYER M2 ;
        RECT 42.844 20.732 42.916 20.764 ;
  LAYER M1 ;
        RECT 45.424 23.82 45.456 23.892 ;
  LAYER M2 ;
        RECT 45.404 23.84 45.476 23.872 ;
  LAYER M1 ;
        RECT 45.424 23.688 45.456 23.856 ;
  LAYER M1 ;
        RECT 45.424 23.652 45.456 23.724 ;
  LAYER M2 ;
        RECT 45.404 23.672 45.476 23.704 ;
  LAYER M2 ;
        RECT 42.88 23.672 45.44 23.704 ;
  LAYER M1 ;
        RECT 42.864 23.652 42.896 23.724 ;
  LAYER M2 ;
        RECT 42.844 23.672 42.916 23.704 ;
  LAYER M1 ;
        RECT 45.424 26.76 45.456 26.832 ;
  LAYER M2 ;
        RECT 45.404 26.78 45.476 26.812 ;
  LAYER M1 ;
        RECT 45.424 26.628 45.456 26.796 ;
  LAYER M1 ;
        RECT 45.424 26.592 45.456 26.664 ;
  LAYER M2 ;
        RECT 45.404 26.612 45.476 26.644 ;
  LAYER M2 ;
        RECT 42.88 26.612 45.44 26.644 ;
  LAYER M1 ;
        RECT 42.864 26.592 42.896 26.664 ;
  LAYER M2 ;
        RECT 42.844 26.612 42.916 26.644 ;
  LAYER M1 ;
        RECT 42.544 17.94 42.576 18.012 ;
  LAYER M2 ;
        RECT 42.524 17.96 42.596 17.992 ;
  LAYER M2 ;
        RECT 42.56 17.96 42.88 17.992 ;
  LAYER M1 ;
        RECT 42.864 17.94 42.896 18.012 ;
  LAYER M2 ;
        RECT 42.844 17.96 42.916 17.992 ;
  LAYER M1 ;
        RECT 42.544 26.76 42.576 26.832 ;
  LAYER M2 ;
        RECT 42.524 26.78 42.596 26.812 ;
  LAYER M2 ;
        RECT 42.56 26.78 42.88 26.812 ;
  LAYER M1 ;
        RECT 42.864 26.76 42.896 26.832 ;
  LAYER M2 ;
        RECT 42.844 26.78 42.916 26.812 ;
  LAYER M1 ;
        RECT 42.864 17.268 42.896 17.34 ;
  LAYER M2 ;
        RECT 42.844 17.288 42.916 17.32 ;
  LAYER M1 ;
        RECT 42.864 17.304 42.896 17.64 ;
  LAYER M1 ;
        RECT 42.864 17.64 42.896 26.796 ;
  LAYER M1 ;
        RECT 36.784 17.94 36.816 18.012 ;
  LAYER M2 ;
        RECT 36.764 17.96 36.836 17.992 ;
  LAYER M1 ;
        RECT 36.784 17.808 36.816 17.976 ;
  LAYER M1 ;
        RECT 36.784 17.772 36.816 17.844 ;
  LAYER M2 ;
        RECT 36.764 17.792 36.836 17.824 ;
  LAYER M2 ;
        RECT 34.24 17.792 36.8 17.824 ;
  LAYER M1 ;
        RECT 34.224 17.772 34.256 17.844 ;
  LAYER M2 ;
        RECT 34.204 17.792 34.276 17.824 ;
  LAYER M1 ;
        RECT 36.784 26.76 36.816 26.832 ;
  LAYER M2 ;
        RECT 36.764 26.78 36.836 26.812 ;
  LAYER M1 ;
        RECT 36.784 26.628 36.816 26.796 ;
  LAYER M1 ;
        RECT 36.784 26.592 36.816 26.664 ;
  LAYER M2 ;
        RECT 36.764 26.612 36.836 26.644 ;
  LAYER M2 ;
        RECT 34.24 26.612 36.8 26.644 ;
  LAYER M1 ;
        RECT 34.224 26.592 34.256 26.664 ;
  LAYER M2 ;
        RECT 34.204 26.612 34.276 26.644 ;
  LAYER M1 ;
        RECT 33.904 17.94 33.936 18.012 ;
  LAYER M2 ;
        RECT 33.884 17.96 33.956 17.992 ;
  LAYER M2 ;
        RECT 33.92 17.96 34.24 17.992 ;
  LAYER M1 ;
        RECT 34.224 17.94 34.256 18.012 ;
  LAYER M2 ;
        RECT 34.204 17.96 34.276 17.992 ;
  LAYER M1 ;
        RECT 33.904 20.88 33.936 20.952 ;
  LAYER M2 ;
        RECT 33.884 20.9 33.956 20.932 ;
  LAYER M2 ;
        RECT 33.92 20.9 34.24 20.932 ;
  LAYER M1 ;
        RECT 34.224 20.88 34.256 20.952 ;
  LAYER M2 ;
        RECT 34.204 20.9 34.276 20.932 ;
  LAYER M1 ;
        RECT 33.904 23.82 33.936 23.892 ;
  LAYER M2 ;
        RECT 33.884 23.84 33.956 23.872 ;
  LAYER M2 ;
        RECT 33.92 23.84 34.24 23.872 ;
  LAYER M1 ;
        RECT 34.224 23.82 34.256 23.892 ;
  LAYER M2 ;
        RECT 34.204 23.84 34.276 23.872 ;
  LAYER M1 ;
        RECT 33.904 26.76 33.936 26.832 ;
  LAYER M2 ;
        RECT 33.884 26.78 33.956 26.812 ;
  LAYER M2 ;
        RECT 33.92 26.78 34.24 26.812 ;
  LAYER M1 ;
        RECT 34.224 26.76 34.256 26.832 ;
  LAYER M2 ;
        RECT 34.204 26.78 34.276 26.812 ;
  LAYER M1 ;
        RECT 34.224 17.268 34.256 17.34 ;
  LAYER M2 ;
        RECT 34.204 17.288 34.276 17.32 ;
  LAYER M1 ;
        RECT 34.224 17.304 34.256 17.64 ;
  LAYER M1 ;
        RECT 34.224 17.64 34.256 26.796 ;
  LAYER M2 ;
        RECT 34.24 17.288 42.88 17.32 ;
  LAYER M1 ;
        RECT 39.664 26.76 39.696 26.832 ;
  LAYER M2 ;
        RECT 39.644 26.78 39.716 26.812 ;
  LAYER M2 ;
        RECT 39.68 26.78 42.56 26.812 ;
  LAYER M1 ;
        RECT 42.544 26.76 42.576 26.832 ;
  LAYER M2 ;
        RECT 42.524 26.78 42.596 26.812 ;
  LAYER M1 ;
        RECT 39.664 17.94 39.696 18.012 ;
  LAYER M2 ;
        RECT 39.644 17.96 39.716 17.992 ;
  LAYER M2 ;
        RECT 36.8 17.96 39.68 17.992 ;
  LAYER M1 ;
        RECT 36.784 17.94 36.816 18.012 ;
  LAYER M2 ;
        RECT 36.764 17.96 36.836 17.992 ;
  LAYER M1 ;
        RECT 37.264 23.316 37.296 23.388 ;
  LAYER M2 ;
        RECT 37.244 23.336 37.316 23.368 ;
  LAYER M2 ;
        RECT 37.28 23.336 39.84 23.368 ;
  LAYER M1 ;
        RECT 39.824 23.316 39.856 23.388 ;
  LAYER M2 ;
        RECT 39.804 23.336 39.876 23.368 ;
  LAYER M1 ;
        RECT 37.264 26.256 37.296 26.328 ;
  LAYER M2 ;
        RECT 37.244 26.276 37.316 26.308 ;
  LAYER M2 ;
        RECT 37.28 26.276 39.84 26.308 ;
  LAYER M1 ;
        RECT 39.824 26.256 39.856 26.328 ;
  LAYER M2 ;
        RECT 39.804 26.276 39.876 26.308 ;
  LAYER M1 ;
        RECT 40.144 23.316 40.176 23.388 ;
  LAYER M2 ;
        RECT 40.124 23.336 40.196 23.368 ;
  LAYER M1 ;
        RECT 40.144 23.352 40.176 23.52 ;
  LAYER M1 ;
        RECT 40.144 23.484 40.176 23.556 ;
  LAYER M2 ;
        RECT 40.124 23.504 40.196 23.536 ;
  LAYER M2 ;
        RECT 39.84 23.504 40.16 23.536 ;
  LAYER M1 ;
        RECT 39.824 23.484 39.856 23.556 ;
  LAYER M2 ;
        RECT 39.804 23.504 39.876 23.536 ;
  LAYER M1 ;
        RECT 40.144 26.256 40.176 26.328 ;
  LAYER M2 ;
        RECT 40.124 26.276 40.196 26.308 ;
  LAYER M1 ;
        RECT 40.144 26.292 40.176 26.46 ;
  LAYER M1 ;
        RECT 40.144 26.424 40.176 26.496 ;
  LAYER M2 ;
        RECT 40.124 26.444 40.196 26.476 ;
  LAYER M2 ;
        RECT 39.84 26.444 40.16 26.476 ;
  LAYER M1 ;
        RECT 39.824 26.424 39.856 26.496 ;
  LAYER M2 ;
        RECT 39.804 26.444 39.876 26.476 ;
  LAYER M1 ;
        RECT 39.824 29.7 39.856 29.772 ;
  LAYER M2 ;
        RECT 39.804 29.72 39.876 29.752 ;
  LAYER M1 ;
        RECT 39.824 29.568 39.856 29.736 ;
  LAYER M1 ;
        RECT 39.824 23.352 39.856 29.568 ;
  LAYER M1 ;
        RECT 34.384 26.256 34.416 26.328 ;
  LAYER M2 ;
        RECT 34.364 26.276 34.436 26.308 ;
  LAYER M2 ;
        RECT 34.4 26.276 36.96 26.308 ;
  LAYER M1 ;
        RECT 36.944 26.256 36.976 26.328 ;
  LAYER M2 ;
        RECT 36.924 26.276 36.996 26.308 ;
  LAYER M1 ;
        RECT 34.384 23.316 34.416 23.388 ;
  LAYER M2 ;
        RECT 34.364 23.336 34.436 23.368 ;
  LAYER M2 ;
        RECT 34.4 23.336 36.96 23.368 ;
  LAYER M1 ;
        RECT 36.944 23.316 36.976 23.388 ;
  LAYER M2 ;
        RECT 36.924 23.336 36.996 23.368 ;
  LAYER M1 ;
        RECT 36.944 29.7 36.976 29.772 ;
  LAYER M2 ;
        RECT 36.924 29.72 36.996 29.752 ;
  LAYER M1 ;
        RECT 36.944 29.568 36.976 29.736 ;
  LAYER M1 ;
        RECT 36.944 23.352 36.976 29.568 ;
  LAYER M2 ;
        RECT 36.96 29.72 39.84 29.752 ;
  LAYER M1 ;
        RECT 43.024 20.376 43.056 20.448 ;
  LAYER M2 ;
        RECT 43.004 20.396 43.076 20.428 ;
  LAYER M2 ;
        RECT 43.04 20.396 45.76 20.428 ;
  LAYER M1 ;
        RECT 45.744 20.376 45.776 20.448 ;
  LAYER M2 ;
        RECT 45.724 20.396 45.796 20.428 ;
  LAYER M1 ;
        RECT 43.024 23.316 43.056 23.388 ;
  LAYER M2 ;
        RECT 43.004 23.336 43.076 23.368 ;
  LAYER M2 ;
        RECT 43.04 23.336 45.76 23.368 ;
  LAYER M1 ;
        RECT 45.744 23.316 45.776 23.388 ;
  LAYER M2 ;
        RECT 45.724 23.336 45.796 23.368 ;
  LAYER M1 ;
        RECT 43.024 26.256 43.056 26.328 ;
  LAYER M2 ;
        RECT 43.004 26.276 43.076 26.308 ;
  LAYER M2 ;
        RECT 43.04 26.276 45.76 26.308 ;
  LAYER M1 ;
        RECT 45.744 26.256 45.776 26.328 ;
  LAYER M2 ;
        RECT 45.724 26.276 45.796 26.308 ;
  LAYER M1 ;
        RECT 43.024 29.196 43.056 29.268 ;
  LAYER M2 ;
        RECT 43.004 29.216 43.076 29.248 ;
  LAYER M2 ;
        RECT 43.04 29.216 45.76 29.248 ;
  LAYER M1 ;
        RECT 45.744 29.196 45.776 29.268 ;
  LAYER M2 ;
        RECT 45.724 29.216 45.796 29.248 ;
  LAYER M1 ;
        RECT 45.744 29.868 45.776 29.94 ;
  LAYER M2 ;
        RECT 45.724 29.888 45.796 29.92 ;
  LAYER M1 ;
        RECT 45.744 29.568 45.776 29.904 ;
  LAYER M1 ;
        RECT 45.744 20.412 45.776 29.568 ;
  LAYER M1 ;
        RECT 31.504 20.376 31.536 20.448 ;
  LAYER M2 ;
        RECT 31.484 20.396 31.556 20.428 ;
  LAYER M1 ;
        RECT 31.504 20.412 31.536 20.58 ;
  LAYER M1 ;
        RECT 31.504 20.544 31.536 20.616 ;
  LAYER M2 ;
        RECT 31.484 20.564 31.556 20.596 ;
  LAYER M2 ;
        RECT 31.36 20.564 31.52 20.596 ;
  LAYER M1 ;
        RECT 31.344 20.544 31.376 20.616 ;
  LAYER M2 ;
        RECT 31.324 20.564 31.396 20.596 ;
  LAYER M1 ;
        RECT 31.504 23.316 31.536 23.388 ;
  LAYER M2 ;
        RECT 31.484 23.336 31.556 23.368 ;
  LAYER M1 ;
        RECT 31.504 23.352 31.536 23.52 ;
  LAYER M1 ;
        RECT 31.504 23.484 31.536 23.556 ;
  LAYER M2 ;
        RECT 31.484 23.504 31.556 23.536 ;
  LAYER M2 ;
        RECT 31.36 23.504 31.52 23.536 ;
  LAYER M1 ;
        RECT 31.344 23.484 31.376 23.556 ;
  LAYER M2 ;
        RECT 31.324 23.504 31.396 23.536 ;
  LAYER M1 ;
        RECT 31.504 26.256 31.536 26.328 ;
  LAYER M2 ;
        RECT 31.484 26.276 31.556 26.308 ;
  LAYER M1 ;
        RECT 31.504 26.292 31.536 26.46 ;
  LAYER M1 ;
        RECT 31.504 26.424 31.536 26.496 ;
  LAYER M2 ;
        RECT 31.484 26.444 31.556 26.476 ;
  LAYER M2 ;
        RECT 31.36 26.444 31.52 26.476 ;
  LAYER M1 ;
        RECT 31.344 26.424 31.376 26.496 ;
  LAYER M2 ;
        RECT 31.324 26.444 31.396 26.476 ;
  LAYER M1 ;
        RECT 31.504 29.196 31.536 29.268 ;
  LAYER M2 ;
        RECT 31.484 29.216 31.556 29.248 ;
  LAYER M1 ;
        RECT 31.504 29.232 31.536 29.4 ;
  LAYER M1 ;
        RECT 31.504 29.364 31.536 29.436 ;
  LAYER M2 ;
        RECT 31.484 29.384 31.556 29.416 ;
  LAYER M2 ;
        RECT 31.36 29.384 31.52 29.416 ;
  LAYER M1 ;
        RECT 31.344 29.364 31.376 29.436 ;
  LAYER M2 ;
        RECT 31.324 29.384 31.396 29.416 ;
  LAYER M1 ;
        RECT 31.344 29.868 31.376 29.94 ;
  LAYER M2 ;
        RECT 31.324 29.888 31.396 29.92 ;
  LAYER M1 ;
        RECT 31.344 29.568 31.376 29.904 ;
  LAYER M1 ;
        RECT 31.344 20.58 31.376 29.568 ;
  LAYER M2 ;
        RECT 31.36 29.888 45.76 29.92 ;
  LAYER M1 ;
        RECT 40.144 20.376 40.176 20.448 ;
  LAYER M2 ;
        RECT 40.124 20.396 40.196 20.428 ;
  LAYER M2 ;
        RECT 40.16 20.396 43.04 20.428 ;
  LAYER M1 ;
        RECT 43.024 20.376 43.056 20.448 ;
  LAYER M2 ;
        RECT 43.004 20.396 43.076 20.428 ;
  LAYER M1 ;
        RECT 40.144 29.196 40.176 29.268 ;
  LAYER M2 ;
        RECT 40.124 29.216 40.196 29.248 ;
  LAYER M2 ;
        RECT 40.16 29.216 43.04 29.248 ;
  LAYER M1 ;
        RECT 43.024 29.196 43.056 29.268 ;
  LAYER M2 ;
        RECT 43.004 29.216 43.076 29.248 ;
  LAYER M1 ;
        RECT 37.264 29.196 37.296 29.268 ;
  LAYER M2 ;
        RECT 37.244 29.216 37.316 29.248 ;
  LAYER M2 ;
        RECT 37.28 29.216 40.16 29.248 ;
  LAYER M1 ;
        RECT 40.144 29.196 40.176 29.268 ;
  LAYER M2 ;
        RECT 40.124 29.216 40.196 29.248 ;
  LAYER M1 ;
        RECT 34.384 29.196 34.416 29.268 ;
  LAYER M2 ;
        RECT 34.364 29.216 34.436 29.248 ;
  LAYER M2 ;
        RECT 34.4 29.216 37.28 29.248 ;
  LAYER M1 ;
        RECT 37.264 29.196 37.296 29.268 ;
  LAYER M2 ;
        RECT 37.244 29.216 37.316 29.248 ;
  LAYER M1 ;
        RECT 34.384 20.376 34.416 20.448 ;
  LAYER M2 ;
        RECT 34.364 20.396 34.436 20.428 ;
  LAYER M2 ;
        RECT 31.52 20.396 34.4 20.428 ;
  LAYER M1 ;
        RECT 31.504 20.376 31.536 20.448 ;
  LAYER M2 ;
        RECT 31.484 20.396 31.556 20.428 ;
  LAYER M1 ;
        RECT 37.264 20.376 37.296 20.448 ;
  LAYER M2 ;
        RECT 37.244 20.396 37.316 20.428 ;
  LAYER M2 ;
        RECT 34.4 20.396 37.28 20.428 ;
  LAYER M1 ;
        RECT 34.384 20.376 34.416 20.448 ;
  LAYER M2 ;
        RECT 34.364 20.396 34.436 20.428 ;
  LAYER M1 ;
        RECT 45.424 17.94 45.456 20.448 ;
  LAYER M1 ;
        RECT 45.36 17.94 45.392 20.448 ;
  LAYER M1 ;
        RECT 45.296 17.94 45.328 20.448 ;
  LAYER M1 ;
        RECT 45.232 17.94 45.264 20.448 ;
  LAYER M1 ;
        RECT 45.168 17.94 45.2 20.448 ;
  LAYER M1 ;
        RECT 45.104 17.94 45.136 20.448 ;
  LAYER M1 ;
        RECT 45.04 17.94 45.072 20.448 ;
  LAYER M1 ;
        RECT 44.976 17.94 45.008 20.448 ;
  LAYER M1 ;
        RECT 44.912 17.94 44.944 20.448 ;
  LAYER M1 ;
        RECT 44.848 17.94 44.88 20.448 ;
  LAYER M1 ;
        RECT 44.784 17.94 44.816 20.448 ;
  LAYER M1 ;
        RECT 44.72 17.94 44.752 20.448 ;
  LAYER M1 ;
        RECT 44.656 17.94 44.688 20.448 ;
  LAYER M1 ;
        RECT 44.592 17.94 44.624 20.448 ;
  LAYER M1 ;
        RECT 44.528 17.94 44.56 20.448 ;
  LAYER M1 ;
        RECT 44.464 17.94 44.496 20.448 ;
  LAYER M1 ;
        RECT 44.4 17.94 44.432 20.448 ;
  LAYER M1 ;
        RECT 44.336 17.94 44.368 20.448 ;
  LAYER M1 ;
        RECT 44.272 17.94 44.304 20.448 ;
  LAYER M1 ;
        RECT 44.208 17.94 44.24 20.448 ;
  LAYER M1 ;
        RECT 44.144 17.94 44.176 20.448 ;
  LAYER M1 ;
        RECT 44.08 17.94 44.112 20.448 ;
  LAYER M1 ;
        RECT 44.016 17.94 44.048 20.448 ;
  LAYER M1 ;
        RECT 43.952 17.94 43.984 20.448 ;
  LAYER M1 ;
        RECT 43.888 17.94 43.92 20.448 ;
  LAYER M1 ;
        RECT 43.824 17.94 43.856 20.448 ;
  LAYER M1 ;
        RECT 43.76 17.94 43.792 20.448 ;
  LAYER M1 ;
        RECT 43.696 17.94 43.728 20.448 ;
  LAYER M1 ;
        RECT 43.632 17.94 43.664 20.448 ;
  LAYER M1 ;
        RECT 43.568 17.94 43.6 20.448 ;
  LAYER M1 ;
        RECT 43.504 17.94 43.536 20.448 ;
  LAYER M1 ;
        RECT 43.44 17.94 43.472 20.448 ;
  LAYER M1 ;
        RECT 43.376 17.94 43.408 20.448 ;
  LAYER M1 ;
        RECT 43.312 17.94 43.344 20.448 ;
  LAYER M1 ;
        RECT 43.248 17.94 43.28 20.448 ;
  LAYER M1 ;
        RECT 43.184 17.94 43.216 20.448 ;
  LAYER M1 ;
        RECT 43.12 17.94 43.152 20.448 ;
  LAYER M2 ;
        RECT 43.004 18.024 45.476 18.056 ;
  LAYER M2 ;
        RECT 43.004 18.088 45.476 18.12 ;
  LAYER M2 ;
        RECT 43.004 18.152 45.476 18.184 ;
  LAYER M2 ;
        RECT 43.004 18.216 45.476 18.248 ;
  LAYER M2 ;
        RECT 43.004 18.28 45.476 18.312 ;
  LAYER M2 ;
        RECT 43.004 18.344 45.476 18.376 ;
  LAYER M2 ;
        RECT 43.004 18.408 45.476 18.44 ;
  LAYER M2 ;
        RECT 43.004 18.472 45.476 18.504 ;
  LAYER M2 ;
        RECT 43.004 18.536 45.476 18.568 ;
  LAYER M2 ;
        RECT 43.004 18.6 45.476 18.632 ;
  LAYER M2 ;
        RECT 43.004 18.664 45.476 18.696 ;
  LAYER M2 ;
        RECT 43.004 18.728 45.476 18.76 ;
  LAYER M2 ;
        RECT 43.004 18.792 45.476 18.824 ;
  LAYER M2 ;
        RECT 43.004 18.856 45.476 18.888 ;
  LAYER M2 ;
        RECT 43.004 18.92 45.476 18.952 ;
  LAYER M2 ;
        RECT 43.004 18.984 45.476 19.016 ;
  LAYER M2 ;
        RECT 43.004 19.048 45.476 19.08 ;
  LAYER M2 ;
        RECT 43.004 19.112 45.476 19.144 ;
  LAYER M2 ;
        RECT 43.004 19.176 45.476 19.208 ;
  LAYER M2 ;
        RECT 43.004 19.24 45.476 19.272 ;
  LAYER M2 ;
        RECT 43.004 19.304 45.476 19.336 ;
  LAYER M2 ;
        RECT 43.004 19.368 45.476 19.4 ;
  LAYER M2 ;
        RECT 43.004 19.432 45.476 19.464 ;
  LAYER M2 ;
        RECT 43.004 19.496 45.476 19.528 ;
  LAYER M2 ;
        RECT 43.004 19.56 45.476 19.592 ;
  LAYER M2 ;
        RECT 43.004 19.624 45.476 19.656 ;
  LAYER M2 ;
        RECT 43.004 19.688 45.476 19.72 ;
  LAYER M2 ;
        RECT 43.004 19.752 45.476 19.784 ;
  LAYER M2 ;
        RECT 43.004 19.816 45.476 19.848 ;
  LAYER M2 ;
        RECT 43.004 19.88 45.476 19.912 ;
  LAYER M2 ;
        RECT 43.004 19.944 45.476 19.976 ;
  LAYER M2 ;
        RECT 43.004 20.008 45.476 20.04 ;
  LAYER M2 ;
        RECT 43.004 20.072 45.476 20.104 ;
  LAYER M2 ;
        RECT 43.004 20.136 45.476 20.168 ;
  LAYER M2 ;
        RECT 43.004 20.2 45.476 20.232 ;
  LAYER M2 ;
        RECT 43.004 20.264 45.476 20.296 ;
  LAYER M3 ;
        RECT 45.424 17.94 45.456 20.448 ;
  LAYER M3 ;
        RECT 45.36 17.94 45.392 20.448 ;
  LAYER M3 ;
        RECT 45.296 17.94 45.328 20.448 ;
  LAYER M3 ;
        RECT 45.232 17.94 45.264 20.448 ;
  LAYER M3 ;
        RECT 45.168 17.94 45.2 20.448 ;
  LAYER M3 ;
        RECT 45.104 17.94 45.136 20.448 ;
  LAYER M3 ;
        RECT 45.04 17.94 45.072 20.448 ;
  LAYER M3 ;
        RECT 44.976 17.94 45.008 20.448 ;
  LAYER M3 ;
        RECT 44.912 17.94 44.944 20.448 ;
  LAYER M3 ;
        RECT 44.848 17.94 44.88 20.448 ;
  LAYER M3 ;
        RECT 44.784 17.94 44.816 20.448 ;
  LAYER M3 ;
        RECT 44.72 17.94 44.752 20.448 ;
  LAYER M3 ;
        RECT 44.656 17.94 44.688 20.448 ;
  LAYER M3 ;
        RECT 44.592 17.94 44.624 20.448 ;
  LAYER M3 ;
        RECT 44.528 17.94 44.56 20.448 ;
  LAYER M3 ;
        RECT 44.464 17.94 44.496 20.448 ;
  LAYER M3 ;
        RECT 44.4 17.94 44.432 20.448 ;
  LAYER M3 ;
        RECT 44.336 17.94 44.368 20.448 ;
  LAYER M3 ;
        RECT 44.272 17.94 44.304 20.448 ;
  LAYER M3 ;
        RECT 44.208 17.94 44.24 20.448 ;
  LAYER M3 ;
        RECT 44.144 17.94 44.176 20.448 ;
  LAYER M3 ;
        RECT 44.08 17.94 44.112 20.448 ;
  LAYER M3 ;
        RECT 44.016 17.94 44.048 20.448 ;
  LAYER M3 ;
        RECT 43.952 17.94 43.984 20.448 ;
  LAYER M3 ;
        RECT 43.888 17.94 43.92 20.448 ;
  LAYER M3 ;
        RECT 43.824 17.94 43.856 20.448 ;
  LAYER M3 ;
        RECT 43.76 17.94 43.792 20.448 ;
  LAYER M3 ;
        RECT 43.696 17.94 43.728 20.448 ;
  LAYER M3 ;
        RECT 43.632 17.94 43.664 20.448 ;
  LAYER M3 ;
        RECT 43.568 17.94 43.6 20.448 ;
  LAYER M3 ;
        RECT 43.504 17.94 43.536 20.448 ;
  LAYER M3 ;
        RECT 43.44 17.94 43.472 20.448 ;
  LAYER M3 ;
        RECT 43.376 17.94 43.408 20.448 ;
  LAYER M3 ;
        RECT 43.312 17.94 43.344 20.448 ;
  LAYER M3 ;
        RECT 43.248 17.94 43.28 20.448 ;
  LAYER M3 ;
        RECT 43.184 17.94 43.216 20.448 ;
  LAYER M3 ;
        RECT 43.12 17.94 43.152 20.448 ;
  LAYER M3 ;
        RECT 43.024 17.94 43.056 20.448 ;
  LAYER M1 ;
        RECT 45.439 17.976 45.441 20.412 ;
  LAYER M1 ;
        RECT 45.359 17.976 45.361 20.412 ;
  LAYER M1 ;
        RECT 45.279 17.976 45.281 20.412 ;
  LAYER M1 ;
        RECT 45.199 17.976 45.201 20.412 ;
  LAYER M1 ;
        RECT 45.119 17.976 45.121 20.412 ;
  LAYER M1 ;
        RECT 45.039 17.976 45.041 20.412 ;
  LAYER M1 ;
        RECT 44.959 17.976 44.961 20.412 ;
  LAYER M1 ;
        RECT 44.879 17.976 44.881 20.412 ;
  LAYER M1 ;
        RECT 44.799 17.976 44.801 20.412 ;
  LAYER M1 ;
        RECT 44.719 17.976 44.721 20.412 ;
  LAYER M1 ;
        RECT 44.639 17.976 44.641 20.412 ;
  LAYER M1 ;
        RECT 44.559 17.976 44.561 20.412 ;
  LAYER M1 ;
        RECT 44.479 17.976 44.481 20.412 ;
  LAYER M1 ;
        RECT 44.399 17.976 44.401 20.412 ;
  LAYER M1 ;
        RECT 44.319 17.976 44.321 20.412 ;
  LAYER M1 ;
        RECT 44.239 17.976 44.241 20.412 ;
  LAYER M1 ;
        RECT 44.159 17.976 44.161 20.412 ;
  LAYER M1 ;
        RECT 44.079 17.976 44.081 20.412 ;
  LAYER M1 ;
        RECT 43.999 17.976 44.001 20.412 ;
  LAYER M1 ;
        RECT 43.919 17.976 43.921 20.412 ;
  LAYER M1 ;
        RECT 43.839 17.976 43.841 20.412 ;
  LAYER M1 ;
        RECT 43.759 17.976 43.761 20.412 ;
  LAYER M1 ;
        RECT 43.679 17.976 43.681 20.412 ;
  LAYER M1 ;
        RECT 43.599 17.976 43.601 20.412 ;
  LAYER M1 ;
        RECT 43.519 17.976 43.521 20.412 ;
  LAYER M1 ;
        RECT 43.439 17.976 43.441 20.412 ;
  LAYER M1 ;
        RECT 43.359 17.976 43.361 20.412 ;
  LAYER M1 ;
        RECT 43.279 17.976 43.281 20.412 ;
  LAYER M1 ;
        RECT 43.199 17.976 43.201 20.412 ;
  LAYER M1 ;
        RECT 43.119 17.976 43.121 20.412 ;
  LAYER M2 ;
        RECT 43.04 17.975 45.44 17.977 ;
  LAYER M2 ;
        RECT 43.04 18.059 45.44 18.061 ;
  LAYER M2 ;
        RECT 43.04 18.143 45.44 18.145 ;
  LAYER M2 ;
        RECT 43.04 18.227 45.44 18.229 ;
  LAYER M2 ;
        RECT 43.04 18.311 45.44 18.313 ;
  LAYER M2 ;
        RECT 43.04 18.395 45.44 18.397 ;
  LAYER M2 ;
        RECT 43.04 18.479 45.44 18.481 ;
  LAYER M2 ;
        RECT 43.04 18.563 45.44 18.565 ;
  LAYER M2 ;
        RECT 43.04 18.647 45.44 18.649 ;
  LAYER M2 ;
        RECT 43.04 18.731 45.44 18.733 ;
  LAYER M2 ;
        RECT 43.04 18.815 45.44 18.817 ;
  LAYER M2 ;
        RECT 43.04 18.899 45.44 18.901 ;
  LAYER M2 ;
        RECT 43.04 18.9825 45.44 18.9845 ;
  LAYER M2 ;
        RECT 43.04 19.067 45.44 19.069 ;
  LAYER M2 ;
        RECT 43.04 19.151 45.44 19.153 ;
  LAYER M2 ;
        RECT 43.04 19.235 45.44 19.237 ;
  LAYER M2 ;
        RECT 43.04 19.319 45.44 19.321 ;
  LAYER M2 ;
        RECT 43.04 19.403 45.44 19.405 ;
  LAYER M2 ;
        RECT 43.04 19.487 45.44 19.489 ;
  LAYER M2 ;
        RECT 43.04 19.571 45.44 19.573 ;
  LAYER M2 ;
        RECT 43.04 19.655 45.44 19.657 ;
  LAYER M2 ;
        RECT 43.04 19.739 45.44 19.741 ;
  LAYER M2 ;
        RECT 43.04 19.823 45.44 19.825 ;
  LAYER M2 ;
        RECT 43.04 19.907 45.44 19.909 ;
  LAYER M2 ;
        RECT 43.04 19.991 45.44 19.993 ;
  LAYER M2 ;
        RECT 43.04 20.075 45.44 20.077 ;
  LAYER M2 ;
        RECT 43.04 20.159 45.44 20.161 ;
  LAYER M2 ;
        RECT 43.04 20.243 45.44 20.245 ;
  LAYER M2 ;
        RECT 43.04 20.327 45.44 20.329 ;
  LAYER M1 ;
        RECT 45.424 20.88 45.456 23.388 ;
  LAYER M1 ;
        RECT 45.36 20.88 45.392 23.388 ;
  LAYER M1 ;
        RECT 45.296 20.88 45.328 23.388 ;
  LAYER M1 ;
        RECT 45.232 20.88 45.264 23.388 ;
  LAYER M1 ;
        RECT 45.168 20.88 45.2 23.388 ;
  LAYER M1 ;
        RECT 45.104 20.88 45.136 23.388 ;
  LAYER M1 ;
        RECT 45.04 20.88 45.072 23.388 ;
  LAYER M1 ;
        RECT 44.976 20.88 45.008 23.388 ;
  LAYER M1 ;
        RECT 44.912 20.88 44.944 23.388 ;
  LAYER M1 ;
        RECT 44.848 20.88 44.88 23.388 ;
  LAYER M1 ;
        RECT 44.784 20.88 44.816 23.388 ;
  LAYER M1 ;
        RECT 44.72 20.88 44.752 23.388 ;
  LAYER M1 ;
        RECT 44.656 20.88 44.688 23.388 ;
  LAYER M1 ;
        RECT 44.592 20.88 44.624 23.388 ;
  LAYER M1 ;
        RECT 44.528 20.88 44.56 23.388 ;
  LAYER M1 ;
        RECT 44.464 20.88 44.496 23.388 ;
  LAYER M1 ;
        RECT 44.4 20.88 44.432 23.388 ;
  LAYER M1 ;
        RECT 44.336 20.88 44.368 23.388 ;
  LAYER M1 ;
        RECT 44.272 20.88 44.304 23.388 ;
  LAYER M1 ;
        RECT 44.208 20.88 44.24 23.388 ;
  LAYER M1 ;
        RECT 44.144 20.88 44.176 23.388 ;
  LAYER M1 ;
        RECT 44.08 20.88 44.112 23.388 ;
  LAYER M1 ;
        RECT 44.016 20.88 44.048 23.388 ;
  LAYER M1 ;
        RECT 43.952 20.88 43.984 23.388 ;
  LAYER M1 ;
        RECT 43.888 20.88 43.92 23.388 ;
  LAYER M1 ;
        RECT 43.824 20.88 43.856 23.388 ;
  LAYER M1 ;
        RECT 43.76 20.88 43.792 23.388 ;
  LAYER M1 ;
        RECT 43.696 20.88 43.728 23.388 ;
  LAYER M1 ;
        RECT 43.632 20.88 43.664 23.388 ;
  LAYER M1 ;
        RECT 43.568 20.88 43.6 23.388 ;
  LAYER M1 ;
        RECT 43.504 20.88 43.536 23.388 ;
  LAYER M1 ;
        RECT 43.44 20.88 43.472 23.388 ;
  LAYER M1 ;
        RECT 43.376 20.88 43.408 23.388 ;
  LAYER M1 ;
        RECT 43.312 20.88 43.344 23.388 ;
  LAYER M1 ;
        RECT 43.248 20.88 43.28 23.388 ;
  LAYER M1 ;
        RECT 43.184 20.88 43.216 23.388 ;
  LAYER M1 ;
        RECT 43.12 20.88 43.152 23.388 ;
  LAYER M2 ;
        RECT 43.004 20.964 45.476 20.996 ;
  LAYER M2 ;
        RECT 43.004 21.028 45.476 21.06 ;
  LAYER M2 ;
        RECT 43.004 21.092 45.476 21.124 ;
  LAYER M2 ;
        RECT 43.004 21.156 45.476 21.188 ;
  LAYER M2 ;
        RECT 43.004 21.22 45.476 21.252 ;
  LAYER M2 ;
        RECT 43.004 21.284 45.476 21.316 ;
  LAYER M2 ;
        RECT 43.004 21.348 45.476 21.38 ;
  LAYER M2 ;
        RECT 43.004 21.412 45.476 21.444 ;
  LAYER M2 ;
        RECT 43.004 21.476 45.476 21.508 ;
  LAYER M2 ;
        RECT 43.004 21.54 45.476 21.572 ;
  LAYER M2 ;
        RECT 43.004 21.604 45.476 21.636 ;
  LAYER M2 ;
        RECT 43.004 21.668 45.476 21.7 ;
  LAYER M2 ;
        RECT 43.004 21.732 45.476 21.764 ;
  LAYER M2 ;
        RECT 43.004 21.796 45.476 21.828 ;
  LAYER M2 ;
        RECT 43.004 21.86 45.476 21.892 ;
  LAYER M2 ;
        RECT 43.004 21.924 45.476 21.956 ;
  LAYER M2 ;
        RECT 43.004 21.988 45.476 22.02 ;
  LAYER M2 ;
        RECT 43.004 22.052 45.476 22.084 ;
  LAYER M2 ;
        RECT 43.004 22.116 45.476 22.148 ;
  LAYER M2 ;
        RECT 43.004 22.18 45.476 22.212 ;
  LAYER M2 ;
        RECT 43.004 22.244 45.476 22.276 ;
  LAYER M2 ;
        RECT 43.004 22.308 45.476 22.34 ;
  LAYER M2 ;
        RECT 43.004 22.372 45.476 22.404 ;
  LAYER M2 ;
        RECT 43.004 22.436 45.476 22.468 ;
  LAYER M2 ;
        RECT 43.004 22.5 45.476 22.532 ;
  LAYER M2 ;
        RECT 43.004 22.564 45.476 22.596 ;
  LAYER M2 ;
        RECT 43.004 22.628 45.476 22.66 ;
  LAYER M2 ;
        RECT 43.004 22.692 45.476 22.724 ;
  LAYER M2 ;
        RECT 43.004 22.756 45.476 22.788 ;
  LAYER M2 ;
        RECT 43.004 22.82 45.476 22.852 ;
  LAYER M2 ;
        RECT 43.004 22.884 45.476 22.916 ;
  LAYER M2 ;
        RECT 43.004 22.948 45.476 22.98 ;
  LAYER M2 ;
        RECT 43.004 23.012 45.476 23.044 ;
  LAYER M2 ;
        RECT 43.004 23.076 45.476 23.108 ;
  LAYER M2 ;
        RECT 43.004 23.14 45.476 23.172 ;
  LAYER M2 ;
        RECT 43.004 23.204 45.476 23.236 ;
  LAYER M3 ;
        RECT 45.424 20.88 45.456 23.388 ;
  LAYER M3 ;
        RECT 45.36 20.88 45.392 23.388 ;
  LAYER M3 ;
        RECT 45.296 20.88 45.328 23.388 ;
  LAYER M3 ;
        RECT 45.232 20.88 45.264 23.388 ;
  LAYER M3 ;
        RECT 45.168 20.88 45.2 23.388 ;
  LAYER M3 ;
        RECT 45.104 20.88 45.136 23.388 ;
  LAYER M3 ;
        RECT 45.04 20.88 45.072 23.388 ;
  LAYER M3 ;
        RECT 44.976 20.88 45.008 23.388 ;
  LAYER M3 ;
        RECT 44.912 20.88 44.944 23.388 ;
  LAYER M3 ;
        RECT 44.848 20.88 44.88 23.388 ;
  LAYER M3 ;
        RECT 44.784 20.88 44.816 23.388 ;
  LAYER M3 ;
        RECT 44.72 20.88 44.752 23.388 ;
  LAYER M3 ;
        RECT 44.656 20.88 44.688 23.388 ;
  LAYER M3 ;
        RECT 44.592 20.88 44.624 23.388 ;
  LAYER M3 ;
        RECT 44.528 20.88 44.56 23.388 ;
  LAYER M3 ;
        RECT 44.464 20.88 44.496 23.388 ;
  LAYER M3 ;
        RECT 44.4 20.88 44.432 23.388 ;
  LAYER M3 ;
        RECT 44.336 20.88 44.368 23.388 ;
  LAYER M3 ;
        RECT 44.272 20.88 44.304 23.388 ;
  LAYER M3 ;
        RECT 44.208 20.88 44.24 23.388 ;
  LAYER M3 ;
        RECT 44.144 20.88 44.176 23.388 ;
  LAYER M3 ;
        RECT 44.08 20.88 44.112 23.388 ;
  LAYER M3 ;
        RECT 44.016 20.88 44.048 23.388 ;
  LAYER M3 ;
        RECT 43.952 20.88 43.984 23.388 ;
  LAYER M3 ;
        RECT 43.888 20.88 43.92 23.388 ;
  LAYER M3 ;
        RECT 43.824 20.88 43.856 23.388 ;
  LAYER M3 ;
        RECT 43.76 20.88 43.792 23.388 ;
  LAYER M3 ;
        RECT 43.696 20.88 43.728 23.388 ;
  LAYER M3 ;
        RECT 43.632 20.88 43.664 23.388 ;
  LAYER M3 ;
        RECT 43.568 20.88 43.6 23.388 ;
  LAYER M3 ;
        RECT 43.504 20.88 43.536 23.388 ;
  LAYER M3 ;
        RECT 43.44 20.88 43.472 23.388 ;
  LAYER M3 ;
        RECT 43.376 20.88 43.408 23.388 ;
  LAYER M3 ;
        RECT 43.312 20.88 43.344 23.388 ;
  LAYER M3 ;
        RECT 43.248 20.88 43.28 23.388 ;
  LAYER M3 ;
        RECT 43.184 20.88 43.216 23.388 ;
  LAYER M3 ;
        RECT 43.12 20.88 43.152 23.388 ;
  LAYER M3 ;
        RECT 43.024 20.88 43.056 23.388 ;
  LAYER M1 ;
        RECT 45.439 20.916 45.441 23.352 ;
  LAYER M1 ;
        RECT 45.359 20.916 45.361 23.352 ;
  LAYER M1 ;
        RECT 45.279 20.916 45.281 23.352 ;
  LAYER M1 ;
        RECT 45.199 20.916 45.201 23.352 ;
  LAYER M1 ;
        RECT 45.119 20.916 45.121 23.352 ;
  LAYER M1 ;
        RECT 45.039 20.916 45.041 23.352 ;
  LAYER M1 ;
        RECT 44.959 20.916 44.961 23.352 ;
  LAYER M1 ;
        RECT 44.879 20.916 44.881 23.352 ;
  LAYER M1 ;
        RECT 44.799 20.916 44.801 23.352 ;
  LAYER M1 ;
        RECT 44.719 20.916 44.721 23.352 ;
  LAYER M1 ;
        RECT 44.639 20.916 44.641 23.352 ;
  LAYER M1 ;
        RECT 44.559 20.916 44.561 23.352 ;
  LAYER M1 ;
        RECT 44.479 20.916 44.481 23.352 ;
  LAYER M1 ;
        RECT 44.399 20.916 44.401 23.352 ;
  LAYER M1 ;
        RECT 44.319 20.916 44.321 23.352 ;
  LAYER M1 ;
        RECT 44.239 20.916 44.241 23.352 ;
  LAYER M1 ;
        RECT 44.159 20.916 44.161 23.352 ;
  LAYER M1 ;
        RECT 44.079 20.916 44.081 23.352 ;
  LAYER M1 ;
        RECT 43.999 20.916 44.001 23.352 ;
  LAYER M1 ;
        RECT 43.919 20.916 43.921 23.352 ;
  LAYER M1 ;
        RECT 43.839 20.916 43.841 23.352 ;
  LAYER M1 ;
        RECT 43.759 20.916 43.761 23.352 ;
  LAYER M1 ;
        RECT 43.679 20.916 43.681 23.352 ;
  LAYER M1 ;
        RECT 43.599 20.916 43.601 23.352 ;
  LAYER M1 ;
        RECT 43.519 20.916 43.521 23.352 ;
  LAYER M1 ;
        RECT 43.439 20.916 43.441 23.352 ;
  LAYER M1 ;
        RECT 43.359 20.916 43.361 23.352 ;
  LAYER M1 ;
        RECT 43.279 20.916 43.281 23.352 ;
  LAYER M1 ;
        RECT 43.199 20.916 43.201 23.352 ;
  LAYER M1 ;
        RECT 43.119 20.916 43.121 23.352 ;
  LAYER M2 ;
        RECT 43.04 20.915 45.44 20.917 ;
  LAYER M2 ;
        RECT 43.04 20.999 45.44 21.001 ;
  LAYER M2 ;
        RECT 43.04 21.083 45.44 21.085 ;
  LAYER M2 ;
        RECT 43.04 21.167 45.44 21.169 ;
  LAYER M2 ;
        RECT 43.04 21.251 45.44 21.253 ;
  LAYER M2 ;
        RECT 43.04 21.335 45.44 21.337 ;
  LAYER M2 ;
        RECT 43.04 21.419 45.44 21.421 ;
  LAYER M2 ;
        RECT 43.04 21.503 45.44 21.505 ;
  LAYER M2 ;
        RECT 43.04 21.587 45.44 21.589 ;
  LAYER M2 ;
        RECT 43.04 21.671 45.44 21.673 ;
  LAYER M2 ;
        RECT 43.04 21.755 45.44 21.757 ;
  LAYER M2 ;
        RECT 43.04 21.839 45.44 21.841 ;
  LAYER M2 ;
        RECT 43.04 21.9225 45.44 21.9245 ;
  LAYER M2 ;
        RECT 43.04 22.007 45.44 22.009 ;
  LAYER M2 ;
        RECT 43.04 22.091 45.44 22.093 ;
  LAYER M2 ;
        RECT 43.04 22.175 45.44 22.177 ;
  LAYER M2 ;
        RECT 43.04 22.259 45.44 22.261 ;
  LAYER M2 ;
        RECT 43.04 22.343 45.44 22.345 ;
  LAYER M2 ;
        RECT 43.04 22.427 45.44 22.429 ;
  LAYER M2 ;
        RECT 43.04 22.511 45.44 22.513 ;
  LAYER M2 ;
        RECT 43.04 22.595 45.44 22.597 ;
  LAYER M2 ;
        RECT 43.04 22.679 45.44 22.681 ;
  LAYER M2 ;
        RECT 43.04 22.763 45.44 22.765 ;
  LAYER M2 ;
        RECT 43.04 22.847 45.44 22.849 ;
  LAYER M2 ;
        RECT 43.04 22.931 45.44 22.933 ;
  LAYER M2 ;
        RECT 43.04 23.015 45.44 23.017 ;
  LAYER M2 ;
        RECT 43.04 23.099 45.44 23.101 ;
  LAYER M2 ;
        RECT 43.04 23.183 45.44 23.185 ;
  LAYER M2 ;
        RECT 43.04 23.267 45.44 23.269 ;
  LAYER M1 ;
        RECT 45.424 23.82 45.456 26.328 ;
  LAYER M1 ;
        RECT 45.36 23.82 45.392 26.328 ;
  LAYER M1 ;
        RECT 45.296 23.82 45.328 26.328 ;
  LAYER M1 ;
        RECT 45.232 23.82 45.264 26.328 ;
  LAYER M1 ;
        RECT 45.168 23.82 45.2 26.328 ;
  LAYER M1 ;
        RECT 45.104 23.82 45.136 26.328 ;
  LAYER M1 ;
        RECT 45.04 23.82 45.072 26.328 ;
  LAYER M1 ;
        RECT 44.976 23.82 45.008 26.328 ;
  LAYER M1 ;
        RECT 44.912 23.82 44.944 26.328 ;
  LAYER M1 ;
        RECT 44.848 23.82 44.88 26.328 ;
  LAYER M1 ;
        RECT 44.784 23.82 44.816 26.328 ;
  LAYER M1 ;
        RECT 44.72 23.82 44.752 26.328 ;
  LAYER M1 ;
        RECT 44.656 23.82 44.688 26.328 ;
  LAYER M1 ;
        RECT 44.592 23.82 44.624 26.328 ;
  LAYER M1 ;
        RECT 44.528 23.82 44.56 26.328 ;
  LAYER M1 ;
        RECT 44.464 23.82 44.496 26.328 ;
  LAYER M1 ;
        RECT 44.4 23.82 44.432 26.328 ;
  LAYER M1 ;
        RECT 44.336 23.82 44.368 26.328 ;
  LAYER M1 ;
        RECT 44.272 23.82 44.304 26.328 ;
  LAYER M1 ;
        RECT 44.208 23.82 44.24 26.328 ;
  LAYER M1 ;
        RECT 44.144 23.82 44.176 26.328 ;
  LAYER M1 ;
        RECT 44.08 23.82 44.112 26.328 ;
  LAYER M1 ;
        RECT 44.016 23.82 44.048 26.328 ;
  LAYER M1 ;
        RECT 43.952 23.82 43.984 26.328 ;
  LAYER M1 ;
        RECT 43.888 23.82 43.92 26.328 ;
  LAYER M1 ;
        RECT 43.824 23.82 43.856 26.328 ;
  LAYER M1 ;
        RECT 43.76 23.82 43.792 26.328 ;
  LAYER M1 ;
        RECT 43.696 23.82 43.728 26.328 ;
  LAYER M1 ;
        RECT 43.632 23.82 43.664 26.328 ;
  LAYER M1 ;
        RECT 43.568 23.82 43.6 26.328 ;
  LAYER M1 ;
        RECT 43.504 23.82 43.536 26.328 ;
  LAYER M1 ;
        RECT 43.44 23.82 43.472 26.328 ;
  LAYER M1 ;
        RECT 43.376 23.82 43.408 26.328 ;
  LAYER M1 ;
        RECT 43.312 23.82 43.344 26.328 ;
  LAYER M1 ;
        RECT 43.248 23.82 43.28 26.328 ;
  LAYER M1 ;
        RECT 43.184 23.82 43.216 26.328 ;
  LAYER M1 ;
        RECT 43.12 23.82 43.152 26.328 ;
  LAYER M2 ;
        RECT 43.004 23.904 45.476 23.936 ;
  LAYER M2 ;
        RECT 43.004 23.968 45.476 24 ;
  LAYER M2 ;
        RECT 43.004 24.032 45.476 24.064 ;
  LAYER M2 ;
        RECT 43.004 24.096 45.476 24.128 ;
  LAYER M2 ;
        RECT 43.004 24.16 45.476 24.192 ;
  LAYER M2 ;
        RECT 43.004 24.224 45.476 24.256 ;
  LAYER M2 ;
        RECT 43.004 24.288 45.476 24.32 ;
  LAYER M2 ;
        RECT 43.004 24.352 45.476 24.384 ;
  LAYER M2 ;
        RECT 43.004 24.416 45.476 24.448 ;
  LAYER M2 ;
        RECT 43.004 24.48 45.476 24.512 ;
  LAYER M2 ;
        RECT 43.004 24.544 45.476 24.576 ;
  LAYER M2 ;
        RECT 43.004 24.608 45.476 24.64 ;
  LAYER M2 ;
        RECT 43.004 24.672 45.476 24.704 ;
  LAYER M2 ;
        RECT 43.004 24.736 45.476 24.768 ;
  LAYER M2 ;
        RECT 43.004 24.8 45.476 24.832 ;
  LAYER M2 ;
        RECT 43.004 24.864 45.476 24.896 ;
  LAYER M2 ;
        RECT 43.004 24.928 45.476 24.96 ;
  LAYER M2 ;
        RECT 43.004 24.992 45.476 25.024 ;
  LAYER M2 ;
        RECT 43.004 25.056 45.476 25.088 ;
  LAYER M2 ;
        RECT 43.004 25.12 45.476 25.152 ;
  LAYER M2 ;
        RECT 43.004 25.184 45.476 25.216 ;
  LAYER M2 ;
        RECT 43.004 25.248 45.476 25.28 ;
  LAYER M2 ;
        RECT 43.004 25.312 45.476 25.344 ;
  LAYER M2 ;
        RECT 43.004 25.376 45.476 25.408 ;
  LAYER M2 ;
        RECT 43.004 25.44 45.476 25.472 ;
  LAYER M2 ;
        RECT 43.004 25.504 45.476 25.536 ;
  LAYER M2 ;
        RECT 43.004 25.568 45.476 25.6 ;
  LAYER M2 ;
        RECT 43.004 25.632 45.476 25.664 ;
  LAYER M2 ;
        RECT 43.004 25.696 45.476 25.728 ;
  LAYER M2 ;
        RECT 43.004 25.76 45.476 25.792 ;
  LAYER M2 ;
        RECT 43.004 25.824 45.476 25.856 ;
  LAYER M2 ;
        RECT 43.004 25.888 45.476 25.92 ;
  LAYER M2 ;
        RECT 43.004 25.952 45.476 25.984 ;
  LAYER M2 ;
        RECT 43.004 26.016 45.476 26.048 ;
  LAYER M2 ;
        RECT 43.004 26.08 45.476 26.112 ;
  LAYER M2 ;
        RECT 43.004 26.144 45.476 26.176 ;
  LAYER M3 ;
        RECT 45.424 23.82 45.456 26.328 ;
  LAYER M3 ;
        RECT 45.36 23.82 45.392 26.328 ;
  LAYER M3 ;
        RECT 45.296 23.82 45.328 26.328 ;
  LAYER M3 ;
        RECT 45.232 23.82 45.264 26.328 ;
  LAYER M3 ;
        RECT 45.168 23.82 45.2 26.328 ;
  LAYER M3 ;
        RECT 45.104 23.82 45.136 26.328 ;
  LAYER M3 ;
        RECT 45.04 23.82 45.072 26.328 ;
  LAYER M3 ;
        RECT 44.976 23.82 45.008 26.328 ;
  LAYER M3 ;
        RECT 44.912 23.82 44.944 26.328 ;
  LAYER M3 ;
        RECT 44.848 23.82 44.88 26.328 ;
  LAYER M3 ;
        RECT 44.784 23.82 44.816 26.328 ;
  LAYER M3 ;
        RECT 44.72 23.82 44.752 26.328 ;
  LAYER M3 ;
        RECT 44.656 23.82 44.688 26.328 ;
  LAYER M3 ;
        RECT 44.592 23.82 44.624 26.328 ;
  LAYER M3 ;
        RECT 44.528 23.82 44.56 26.328 ;
  LAYER M3 ;
        RECT 44.464 23.82 44.496 26.328 ;
  LAYER M3 ;
        RECT 44.4 23.82 44.432 26.328 ;
  LAYER M3 ;
        RECT 44.336 23.82 44.368 26.328 ;
  LAYER M3 ;
        RECT 44.272 23.82 44.304 26.328 ;
  LAYER M3 ;
        RECT 44.208 23.82 44.24 26.328 ;
  LAYER M3 ;
        RECT 44.144 23.82 44.176 26.328 ;
  LAYER M3 ;
        RECT 44.08 23.82 44.112 26.328 ;
  LAYER M3 ;
        RECT 44.016 23.82 44.048 26.328 ;
  LAYER M3 ;
        RECT 43.952 23.82 43.984 26.328 ;
  LAYER M3 ;
        RECT 43.888 23.82 43.92 26.328 ;
  LAYER M3 ;
        RECT 43.824 23.82 43.856 26.328 ;
  LAYER M3 ;
        RECT 43.76 23.82 43.792 26.328 ;
  LAYER M3 ;
        RECT 43.696 23.82 43.728 26.328 ;
  LAYER M3 ;
        RECT 43.632 23.82 43.664 26.328 ;
  LAYER M3 ;
        RECT 43.568 23.82 43.6 26.328 ;
  LAYER M3 ;
        RECT 43.504 23.82 43.536 26.328 ;
  LAYER M3 ;
        RECT 43.44 23.82 43.472 26.328 ;
  LAYER M3 ;
        RECT 43.376 23.82 43.408 26.328 ;
  LAYER M3 ;
        RECT 43.312 23.82 43.344 26.328 ;
  LAYER M3 ;
        RECT 43.248 23.82 43.28 26.328 ;
  LAYER M3 ;
        RECT 43.184 23.82 43.216 26.328 ;
  LAYER M3 ;
        RECT 43.12 23.82 43.152 26.328 ;
  LAYER M3 ;
        RECT 43.024 23.82 43.056 26.328 ;
  LAYER M1 ;
        RECT 45.439 23.856 45.441 26.292 ;
  LAYER M1 ;
        RECT 45.359 23.856 45.361 26.292 ;
  LAYER M1 ;
        RECT 45.279 23.856 45.281 26.292 ;
  LAYER M1 ;
        RECT 45.199 23.856 45.201 26.292 ;
  LAYER M1 ;
        RECT 45.119 23.856 45.121 26.292 ;
  LAYER M1 ;
        RECT 45.039 23.856 45.041 26.292 ;
  LAYER M1 ;
        RECT 44.959 23.856 44.961 26.292 ;
  LAYER M1 ;
        RECT 44.879 23.856 44.881 26.292 ;
  LAYER M1 ;
        RECT 44.799 23.856 44.801 26.292 ;
  LAYER M1 ;
        RECT 44.719 23.856 44.721 26.292 ;
  LAYER M1 ;
        RECT 44.639 23.856 44.641 26.292 ;
  LAYER M1 ;
        RECT 44.559 23.856 44.561 26.292 ;
  LAYER M1 ;
        RECT 44.479 23.856 44.481 26.292 ;
  LAYER M1 ;
        RECT 44.399 23.856 44.401 26.292 ;
  LAYER M1 ;
        RECT 44.319 23.856 44.321 26.292 ;
  LAYER M1 ;
        RECT 44.239 23.856 44.241 26.292 ;
  LAYER M1 ;
        RECT 44.159 23.856 44.161 26.292 ;
  LAYER M1 ;
        RECT 44.079 23.856 44.081 26.292 ;
  LAYER M1 ;
        RECT 43.999 23.856 44.001 26.292 ;
  LAYER M1 ;
        RECT 43.919 23.856 43.921 26.292 ;
  LAYER M1 ;
        RECT 43.839 23.856 43.841 26.292 ;
  LAYER M1 ;
        RECT 43.759 23.856 43.761 26.292 ;
  LAYER M1 ;
        RECT 43.679 23.856 43.681 26.292 ;
  LAYER M1 ;
        RECT 43.599 23.856 43.601 26.292 ;
  LAYER M1 ;
        RECT 43.519 23.856 43.521 26.292 ;
  LAYER M1 ;
        RECT 43.439 23.856 43.441 26.292 ;
  LAYER M1 ;
        RECT 43.359 23.856 43.361 26.292 ;
  LAYER M1 ;
        RECT 43.279 23.856 43.281 26.292 ;
  LAYER M1 ;
        RECT 43.199 23.856 43.201 26.292 ;
  LAYER M1 ;
        RECT 43.119 23.856 43.121 26.292 ;
  LAYER M2 ;
        RECT 43.04 23.855 45.44 23.857 ;
  LAYER M2 ;
        RECT 43.04 23.939 45.44 23.941 ;
  LAYER M2 ;
        RECT 43.04 24.023 45.44 24.025 ;
  LAYER M2 ;
        RECT 43.04 24.107 45.44 24.109 ;
  LAYER M2 ;
        RECT 43.04 24.191 45.44 24.193 ;
  LAYER M2 ;
        RECT 43.04 24.275 45.44 24.277 ;
  LAYER M2 ;
        RECT 43.04 24.359 45.44 24.361 ;
  LAYER M2 ;
        RECT 43.04 24.443 45.44 24.445 ;
  LAYER M2 ;
        RECT 43.04 24.527 45.44 24.529 ;
  LAYER M2 ;
        RECT 43.04 24.611 45.44 24.613 ;
  LAYER M2 ;
        RECT 43.04 24.695 45.44 24.697 ;
  LAYER M2 ;
        RECT 43.04 24.779 45.44 24.781 ;
  LAYER M2 ;
        RECT 43.04 24.8625 45.44 24.8645 ;
  LAYER M2 ;
        RECT 43.04 24.947 45.44 24.949 ;
  LAYER M2 ;
        RECT 43.04 25.031 45.44 25.033 ;
  LAYER M2 ;
        RECT 43.04 25.115 45.44 25.117 ;
  LAYER M2 ;
        RECT 43.04 25.199 45.44 25.201 ;
  LAYER M2 ;
        RECT 43.04 25.283 45.44 25.285 ;
  LAYER M2 ;
        RECT 43.04 25.367 45.44 25.369 ;
  LAYER M2 ;
        RECT 43.04 25.451 45.44 25.453 ;
  LAYER M2 ;
        RECT 43.04 25.535 45.44 25.537 ;
  LAYER M2 ;
        RECT 43.04 25.619 45.44 25.621 ;
  LAYER M2 ;
        RECT 43.04 25.703 45.44 25.705 ;
  LAYER M2 ;
        RECT 43.04 25.787 45.44 25.789 ;
  LAYER M2 ;
        RECT 43.04 25.871 45.44 25.873 ;
  LAYER M2 ;
        RECT 43.04 25.955 45.44 25.957 ;
  LAYER M2 ;
        RECT 43.04 26.039 45.44 26.041 ;
  LAYER M2 ;
        RECT 43.04 26.123 45.44 26.125 ;
  LAYER M2 ;
        RECT 43.04 26.207 45.44 26.209 ;
  LAYER M1 ;
        RECT 45.424 26.76 45.456 29.268 ;
  LAYER M1 ;
        RECT 45.36 26.76 45.392 29.268 ;
  LAYER M1 ;
        RECT 45.296 26.76 45.328 29.268 ;
  LAYER M1 ;
        RECT 45.232 26.76 45.264 29.268 ;
  LAYER M1 ;
        RECT 45.168 26.76 45.2 29.268 ;
  LAYER M1 ;
        RECT 45.104 26.76 45.136 29.268 ;
  LAYER M1 ;
        RECT 45.04 26.76 45.072 29.268 ;
  LAYER M1 ;
        RECT 44.976 26.76 45.008 29.268 ;
  LAYER M1 ;
        RECT 44.912 26.76 44.944 29.268 ;
  LAYER M1 ;
        RECT 44.848 26.76 44.88 29.268 ;
  LAYER M1 ;
        RECT 44.784 26.76 44.816 29.268 ;
  LAYER M1 ;
        RECT 44.72 26.76 44.752 29.268 ;
  LAYER M1 ;
        RECT 44.656 26.76 44.688 29.268 ;
  LAYER M1 ;
        RECT 44.592 26.76 44.624 29.268 ;
  LAYER M1 ;
        RECT 44.528 26.76 44.56 29.268 ;
  LAYER M1 ;
        RECT 44.464 26.76 44.496 29.268 ;
  LAYER M1 ;
        RECT 44.4 26.76 44.432 29.268 ;
  LAYER M1 ;
        RECT 44.336 26.76 44.368 29.268 ;
  LAYER M1 ;
        RECT 44.272 26.76 44.304 29.268 ;
  LAYER M1 ;
        RECT 44.208 26.76 44.24 29.268 ;
  LAYER M1 ;
        RECT 44.144 26.76 44.176 29.268 ;
  LAYER M1 ;
        RECT 44.08 26.76 44.112 29.268 ;
  LAYER M1 ;
        RECT 44.016 26.76 44.048 29.268 ;
  LAYER M1 ;
        RECT 43.952 26.76 43.984 29.268 ;
  LAYER M1 ;
        RECT 43.888 26.76 43.92 29.268 ;
  LAYER M1 ;
        RECT 43.824 26.76 43.856 29.268 ;
  LAYER M1 ;
        RECT 43.76 26.76 43.792 29.268 ;
  LAYER M1 ;
        RECT 43.696 26.76 43.728 29.268 ;
  LAYER M1 ;
        RECT 43.632 26.76 43.664 29.268 ;
  LAYER M1 ;
        RECT 43.568 26.76 43.6 29.268 ;
  LAYER M1 ;
        RECT 43.504 26.76 43.536 29.268 ;
  LAYER M1 ;
        RECT 43.44 26.76 43.472 29.268 ;
  LAYER M1 ;
        RECT 43.376 26.76 43.408 29.268 ;
  LAYER M1 ;
        RECT 43.312 26.76 43.344 29.268 ;
  LAYER M1 ;
        RECT 43.248 26.76 43.28 29.268 ;
  LAYER M1 ;
        RECT 43.184 26.76 43.216 29.268 ;
  LAYER M1 ;
        RECT 43.12 26.76 43.152 29.268 ;
  LAYER M2 ;
        RECT 43.004 26.844 45.476 26.876 ;
  LAYER M2 ;
        RECT 43.004 26.908 45.476 26.94 ;
  LAYER M2 ;
        RECT 43.004 26.972 45.476 27.004 ;
  LAYER M2 ;
        RECT 43.004 27.036 45.476 27.068 ;
  LAYER M2 ;
        RECT 43.004 27.1 45.476 27.132 ;
  LAYER M2 ;
        RECT 43.004 27.164 45.476 27.196 ;
  LAYER M2 ;
        RECT 43.004 27.228 45.476 27.26 ;
  LAYER M2 ;
        RECT 43.004 27.292 45.476 27.324 ;
  LAYER M2 ;
        RECT 43.004 27.356 45.476 27.388 ;
  LAYER M2 ;
        RECT 43.004 27.42 45.476 27.452 ;
  LAYER M2 ;
        RECT 43.004 27.484 45.476 27.516 ;
  LAYER M2 ;
        RECT 43.004 27.548 45.476 27.58 ;
  LAYER M2 ;
        RECT 43.004 27.612 45.476 27.644 ;
  LAYER M2 ;
        RECT 43.004 27.676 45.476 27.708 ;
  LAYER M2 ;
        RECT 43.004 27.74 45.476 27.772 ;
  LAYER M2 ;
        RECT 43.004 27.804 45.476 27.836 ;
  LAYER M2 ;
        RECT 43.004 27.868 45.476 27.9 ;
  LAYER M2 ;
        RECT 43.004 27.932 45.476 27.964 ;
  LAYER M2 ;
        RECT 43.004 27.996 45.476 28.028 ;
  LAYER M2 ;
        RECT 43.004 28.06 45.476 28.092 ;
  LAYER M2 ;
        RECT 43.004 28.124 45.476 28.156 ;
  LAYER M2 ;
        RECT 43.004 28.188 45.476 28.22 ;
  LAYER M2 ;
        RECT 43.004 28.252 45.476 28.284 ;
  LAYER M2 ;
        RECT 43.004 28.316 45.476 28.348 ;
  LAYER M2 ;
        RECT 43.004 28.38 45.476 28.412 ;
  LAYER M2 ;
        RECT 43.004 28.444 45.476 28.476 ;
  LAYER M2 ;
        RECT 43.004 28.508 45.476 28.54 ;
  LAYER M2 ;
        RECT 43.004 28.572 45.476 28.604 ;
  LAYER M2 ;
        RECT 43.004 28.636 45.476 28.668 ;
  LAYER M2 ;
        RECT 43.004 28.7 45.476 28.732 ;
  LAYER M2 ;
        RECT 43.004 28.764 45.476 28.796 ;
  LAYER M2 ;
        RECT 43.004 28.828 45.476 28.86 ;
  LAYER M2 ;
        RECT 43.004 28.892 45.476 28.924 ;
  LAYER M2 ;
        RECT 43.004 28.956 45.476 28.988 ;
  LAYER M2 ;
        RECT 43.004 29.02 45.476 29.052 ;
  LAYER M2 ;
        RECT 43.004 29.084 45.476 29.116 ;
  LAYER M3 ;
        RECT 45.424 26.76 45.456 29.268 ;
  LAYER M3 ;
        RECT 45.36 26.76 45.392 29.268 ;
  LAYER M3 ;
        RECT 45.296 26.76 45.328 29.268 ;
  LAYER M3 ;
        RECT 45.232 26.76 45.264 29.268 ;
  LAYER M3 ;
        RECT 45.168 26.76 45.2 29.268 ;
  LAYER M3 ;
        RECT 45.104 26.76 45.136 29.268 ;
  LAYER M3 ;
        RECT 45.04 26.76 45.072 29.268 ;
  LAYER M3 ;
        RECT 44.976 26.76 45.008 29.268 ;
  LAYER M3 ;
        RECT 44.912 26.76 44.944 29.268 ;
  LAYER M3 ;
        RECT 44.848 26.76 44.88 29.268 ;
  LAYER M3 ;
        RECT 44.784 26.76 44.816 29.268 ;
  LAYER M3 ;
        RECT 44.72 26.76 44.752 29.268 ;
  LAYER M3 ;
        RECT 44.656 26.76 44.688 29.268 ;
  LAYER M3 ;
        RECT 44.592 26.76 44.624 29.268 ;
  LAYER M3 ;
        RECT 44.528 26.76 44.56 29.268 ;
  LAYER M3 ;
        RECT 44.464 26.76 44.496 29.268 ;
  LAYER M3 ;
        RECT 44.4 26.76 44.432 29.268 ;
  LAYER M3 ;
        RECT 44.336 26.76 44.368 29.268 ;
  LAYER M3 ;
        RECT 44.272 26.76 44.304 29.268 ;
  LAYER M3 ;
        RECT 44.208 26.76 44.24 29.268 ;
  LAYER M3 ;
        RECT 44.144 26.76 44.176 29.268 ;
  LAYER M3 ;
        RECT 44.08 26.76 44.112 29.268 ;
  LAYER M3 ;
        RECT 44.016 26.76 44.048 29.268 ;
  LAYER M3 ;
        RECT 43.952 26.76 43.984 29.268 ;
  LAYER M3 ;
        RECT 43.888 26.76 43.92 29.268 ;
  LAYER M3 ;
        RECT 43.824 26.76 43.856 29.268 ;
  LAYER M3 ;
        RECT 43.76 26.76 43.792 29.268 ;
  LAYER M3 ;
        RECT 43.696 26.76 43.728 29.268 ;
  LAYER M3 ;
        RECT 43.632 26.76 43.664 29.268 ;
  LAYER M3 ;
        RECT 43.568 26.76 43.6 29.268 ;
  LAYER M3 ;
        RECT 43.504 26.76 43.536 29.268 ;
  LAYER M3 ;
        RECT 43.44 26.76 43.472 29.268 ;
  LAYER M3 ;
        RECT 43.376 26.76 43.408 29.268 ;
  LAYER M3 ;
        RECT 43.312 26.76 43.344 29.268 ;
  LAYER M3 ;
        RECT 43.248 26.76 43.28 29.268 ;
  LAYER M3 ;
        RECT 43.184 26.76 43.216 29.268 ;
  LAYER M3 ;
        RECT 43.12 26.76 43.152 29.268 ;
  LAYER M3 ;
        RECT 43.024 26.76 43.056 29.268 ;
  LAYER M1 ;
        RECT 45.439 26.796 45.441 29.232 ;
  LAYER M1 ;
        RECT 45.359 26.796 45.361 29.232 ;
  LAYER M1 ;
        RECT 45.279 26.796 45.281 29.232 ;
  LAYER M1 ;
        RECT 45.199 26.796 45.201 29.232 ;
  LAYER M1 ;
        RECT 45.119 26.796 45.121 29.232 ;
  LAYER M1 ;
        RECT 45.039 26.796 45.041 29.232 ;
  LAYER M1 ;
        RECT 44.959 26.796 44.961 29.232 ;
  LAYER M1 ;
        RECT 44.879 26.796 44.881 29.232 ;
  LAYER M1 ;
        RECT 44.799 26.796 44.801 29.232 ;
  LAYER M1 ;
        RECT 44.719 26.796 44.721 29.232 ;
  LAYER M1 ;
        RECT 44.639 26.796 44.641 29.232 ;
  LAYER M1 ;
        RECT 44.559 26.796 44.561 29.232 ;
  LAYER M1 ;
        RECT 44.479 26.796 44.481 29.232 ;
  LAYER M1 ;
        RECT 44.399 26.796 44.401 29.232 ;
  LAYER M1 ;
        RECT 44.319 26.796 44.321 29.232 ;
  LAYER M1 ;
        RECT 44.239 26.796 44.241 29.232 ;
  LAYER M1 ;
        RECT 44.159 26.796 44.161 29.232 ;
  LAYER M1 ;
        RECT 44.079 26.796 44.081 29.232 ;
  LAYER M1 ;
        RECT 43.999 26.796 44.001 29.232 ;
  LAYER M1 ;
        RECT 43.919 26.796 43.921 29.232 ;
  LAYER M1 ;
        RECT 43.839 26.796 43.841 29.232 ;
  LAYER M1 ;
        RECT 43.759 26.796 43.761 29.232 ;
  LAYER M1 ;
        RECT 43.679 26.796 43.681 29.232 ;
  LAYER M1 ;
        RECT 43.599 26.796 43.601 29.232 ;
  LAYER M1 ;
        RECT 43.519 26.796 43.521 29.232 ;
  LAYER M1 ;
        RECT 43.439 26.796 43.441 29.232 ;
  LAYER M1 ;
        RECT 43.359 26.796 43.361 29.232 ;
  LAYER M1 ;
        RECT 43.279 26.796 43.281 29.232 ;
  LAYER M1 ;
        RECT 43.199 26.796 43.201 29.232 ;
  LAYER M1 ;
        RECT 43.119 26.796 43.121 29.232 ;
  LAYER M2 ;
        RECT 43.04 26.795 45.44 26.797 ;
  LAYER M2 ;
        RECT 43.04 26.879 45.44 26.881 ;
  LAYER M2 ;
        RECT 43.04 26.963 45.44 26.965 ;
  LAYER M2 ;
        RECT 43.04 27.047 45.44 27.049 ;
  LAYER M2 ;
        RECT 43.04 27.131 45.44 27.133 ;
  LAYER M2 ;
        RECT 43.04 27.215 45.44 27.217 ;
  LAYER M2 ;
        RECT 43.04 27.299 45.44 27.301 ;
  LAYER M2 ;
        RECT 43.04 27.383 45.44 27.385 ;
  LAYER M2 ;
        RECT 43.04 27.467 45.44 27.469 ;
  LAYER M2 ;
        RECT 43.04 27.551 45.44 27.553 ;
  LAYER M2 ;
        RECT 43.04 27.635 45.44 27.637 ;
  LAYER M2 ;
        RECT 43.04 27.719 45.44 27.721 ;
  LAYER M2 ;
        RECT 43.04 27.8025 45.44 27.8045 ;
  LAYER M2 ;
        RECT 43.04 27.887 45.44 27.889 ;
  LAYER M2 ;
        RECT 43.04 27.971 45.44 27.973 ;
  LAYER M2 ;
        RECT 43.04 28.055 45.44 28.057 ;
  LAYER M2 ;
        RECT 43.04 28.139 45.44 28.141 ;
  LAYER M2 ;
        RECT 43.04 28.223 45.44 28.225 ;
  LAYER M2 ;
        RECT 43.04 28.307 45.44 28.309 ;
  LAYER M2 ;
        RECT 43.04 28.391 45.44 28.393 ;
  LAYER M2 ;
        RECT 43.04 28.475 45.44 28.477 ;
  LAYER M2 ;
        RECT 43.04 28.559 45.44 28.561 ;
  LAYER M2 ;
        RECT 43.04 28.643 45.44 28.645 ;
  LAYER M2 ;
        RECT 43.04 28.727 45.44 28.729 ;
  LAYER M2 ;
        RECT 43.04 28.811 45.44 28.813 ;
  LAYER M2 ;
        RECT 43.04 28.895 45.44 28.897 ;
  LAYER M2 ;
        RECT 43.04 28.979 45.44 28.981 ;
  LAYER M2 ;
        RECT 43.04 29.063 45.44 29.065 ;
  LAYER M2 ;
        RECT 43.04 29.147 45.44 29.149 ;
  LAYER M1 ;
        RECT 42.544 17.94 42.576 20.448 ;
  LAYER M1 ;
        RECT 42.48 17.94 42.512 20.448 ;
  LAYER M1 ;
        RECT 42.416 17.94 42.448 20.448 ;
  LAYER M1 ;
        RECT 42.352 17.94 42.384 20.448 ;
  LAYER M1 ;
        RECT 42.288 17.94 42.32 20.448 ;
  LAYER M1 ;
        RECT 42.224 17.94 42.256 20.448 ;
  LAYER M1 ;
        RECT 42.16 17.94 42.192 20.448 ;
  LAYER M1 ;
        RECT 42.096 17.94 42.128 20.448 ;
  LAYER M1 ;
        RECT 42.032 17.94 42.064 20.448 ;
  LAYER M1 ;
        RECT 41.968 17.94 42 20.448 ;
  LAYER M1 ;
        RECT 41.904 17.94 41.936 20.448 ;
  LAYER M1 ;
        RECT 41.84 17.94 41.872 20.448 ;
  LAYER M1 ;
        RECT 41.776 17.94 41.808 20.448 ;
  LAYER M1 ;
        RECT 41.712 17.94 41.744 20.448 ;
  LAYER M1 ;
        RECT 41.648 17.94 41.68 20.448 ;
  LAYER M1 ;
        RECT 41.584 17.94 41.616 20.448 ;
  LAYER M1 ;
        RECT 41.52 17.94 41.552 20.448 ;
  LAYER M1 ;
        RECT 41.456 17.94 41.488 20.448 ;
  LAYER M1 ;
        RECT 41.392 17.94 41.424 20.448 ;
  LAYER M1 ;
        RECT 41.328 17.94 41.36 20.448 ;
  LAYER M1 ;
        RECT 41.264 17.94 41.296 20.448 ;
  LAYER M1 ;
        RECT 41.2 17.94 41.232 20.448 ;
  LAYER M1 ;
        RECT 41.136 17.94 41.168 20.448 ;
  LAYER M1 ;
        RECT 41.072 17.94 41.104 20.448 ;
  LAYER M1 ;
        RECT 41.008 17.94 41.04 20.448 ;
  LAYER M1 ;
        RECT 40.944 17.94 40.976 20.448 ;
  LAYER M1 ;
        RECT 40.88 17.94 40.912 20.448 ;
  LAYER M1 ;
        RECT 40.816 17.94 40.848 20.448 ;
  LAYER M1 ;
        RECT 40.752 17.94 40.784 20.448 ;
  LAYER M1 ;
        RECT 40.688 17.94 40.72 20.448 ;
  LAYER M1 ;
        RECT 40.624 17.94 40.656 20.448 ;
  LAYER M1 ;
        RECT 40.56 17.94 40.592 20.448 ;
  LAYER M1 ;
        RECT 40.496 17.94 40.528 20.448 ;
  LAYER M1 ;
        RECT 40.432 17.94 40.464 20.448 ;
  LAYER M1 ;
        RECT 40.368 17.94 40.4 20.448 ;
  LAYER M1 ;
        RECT 40.304 17.94 40.336 20.448 ;
  LAYER M1 ;
        RECT 40.24 17.94 40.272 20.448 ;
  LAYER M2 ;
        RECT 40.124 18.024 42.596 18.056 ;
  LAYER M2 ;
        RECT 40.124 18.088 42.596 18.12 ;
  LAYER M2 ;
        RECT 40.124 18.152 42.596 18.184 ;
  LAYER M2 ;
        RECT 40.124 18.216 42.596 18.248 ;
  LAYER M2 ;
        RECT 40.124 18.28 42.596 18.312 ;
  LAYER M2 ;
        RECT 40.124 18.344 42.596 18.376 ;
  LAYER M2 ;
        RECT 40.124 18.408 42.596 18.44 ;
  LAYER M2 ;
        RECT 40.124 18.472 42.596 18.504 ;
  LAYER M2 ;
        RECT 40.124 18.536 42.596 18.568 ;
  LAYER M2 ;
        RECT 40.124 18.6 42.596 18.632 ;
  LAYER M2 ;
        RECT 40.124 18.664 42.596 18.696 ;
  LAYER M2 ;
        RECT 40.124 18.728 42.596 18.76 ;
  LAYER M2 ;
        RECT 40.124 18.792 42.596 18.824 ;
  LAYER M2 ;
        RECT 40.124 18.856 42.596 18.888 ;
  LAYER M2 ;
        RECT 40.124 18.92 42.596 18.952 ;
  LAYER M2 ;
        RECT 40.124 18.984 42.596 19.016 ;
  LAYER M2 ;
        RECT 40.124 19.048 42.596 19.08 ;
  LAYER M2 ;
        RECT 40.124 19.112 42.596 19.144 ;
  LAYER M2 ;
        RECT 40.124 19.176 42.596 19.208 ;
  LAYER M2 ;
        RECT 40.124 19.24 42.596 19.272 ;
  LAYER M2 ;
        RECT 40.124 19.304 42.596 19.336 ;
  LAYER M2 ;
        RECT 40.124 19.368 42.596 19.4 ;
  LAYER M2 ;
        RECT 40.124 19.432 42.596 19.464 ;
  LAYER M2 ;
        RECT 40.124 19.496 42.596 19.528 ;
  LAYER M2 ;
        RECT 40.124 19.56 42.596 19.592 ;
  LAYER M2 ;
        RECT 40.124 19.624 42.596 19.656 ;
  LAYER M2 ;
        RECT 40.124 19.688 42.596 19.72 ;
  LAYER M2 ;
        RECT 40.124 19.752 42.596 19.784 ;
  LAYER M2 ;
        RECT 40.124 19.816 42.596 19.848 ;
  LAYER M2 ;
        RECT 40.124 19.88 42.596 19.912 ;
  LAYER M2 ;
        RECT 40.124 19.944 42.596 19.976 ;
  LAYER M2 ;
        RECT 40.124 20.008 42.596 20.04 ;
  LAYER M2 ;
        RECT 40.124 20.072 42.596 20.104 ;
  LAYER M2 ;
        RECT 40.124 20.136 42.596 20.168 ;
  LAYER M2 ;
        RECT 40.124 20.2 42.596 20.232 ;
  LAYER M2 ;
        RECT 40.124 20.264 42.596 20.296 ;
  LAYER M3 ;
        RECT 42.544 17.94 42.576 20.448 ;
  LAYER M3 ;
        RECT 42.48 17.94 42.512 20.448 ;
  LAYER M3 ;
        RECT 42.416 17.94 42.448 20.448 ;
  LAYER M3 ;
        RECT 42.352 17.94 42.384 20.448 ;
  LAYER M3 ;
        RECT 42.288 17.94 42.32 20.448 ;
  LAYER M3 ;
        RECT 42.224 17.94 42.256 20.448 ;
  LAYER M3 ;
        RECT 42.16 17.94 42.192 20.448 ;
  LAYER M3 ;
        RECT 42.096 17.94 42.128 20.448 ;
  LAYER M3 ;
        RECT 42.032 17.94 42.064 20.448 ;
  LAYER M3 ;
        RECT 41.968 17.94 42 20.448 ;
  LAYER M3 ;
        RECT 41.904 17.94 41.936 20.448 ;
  LAYER M3 ;
        RECT 41.84 17.94 41.872 20.448 ;
  LAYER M3 ;
        RECT 41.776 17.94 41.808 20.448 ;
  LAYER M3 ;
        RECT 41.712 17.94 41.744 20.448 ;
  LAYER M3 ;
        RECT 41.648 17.94 41.68 20.448 ;
  LAYER M3 ;
        RECT 41.584 17.94 41.616 20.448 ;
  LAYER M3 ;
        RECT 41.52 17.94 41.552 20.448 ;
  LAYER M3 ;
        RECT 41.456 17.94 41.488 20.448 ;
  LAYER M3 ;
        RECT 41.392 17.94 41.424 20.448 ;
  LAYER M3 ;
        RECT 41.328 17.94 41.36 20.448 ;
  LAYER M3 ;
        RECT 41.264 17.94 41.296 20.448 ;
  LAYER M3 ;
        RECT 41.2 17.94 41.232 20.448 ;
  LAYER M3 ;
        RECT 41.136 17.94 41.168 20.448 ;
  LAYER M3 ;
        RECT 41.072 17.94 41.104 20.448 ;
  LAYER M3 ;
        RECT 41.008 17.94 41.04 20.448 ;
  LAYER M3 ;
        RECT 40.944 17.94 40.976 20.448 ;
  LAYER M3 ;
        RECT 40.88 17.94 40.912 20.448 ;
  LAYER M3 ;
        RECT 40.816 17.94 40.848 20.448 ;
  LAYER M3 ;
        RECT 40.752 17.94 40.784 20.448 ;
  LAYER M3 ;
        RECT 40.688 17.94 40.72 20.448 ;
  LAYER M3 ;
        RECT 40.624 17.94 40.656 20.448 ;
  LAYER M3 ;
        RECT 40.56 17.94 40.592 20.448 ;
  LAYER M3 ;
        RECT 40.496 17.94 40.528 20.448 ;
  LAYER M3 ;
        RECT 40.432 17.94 40.464 20.448 ;
  LAYER M3 ;
        RECT 40.368 17.94 40.4 20.448 ;
  LAYER M3 ;
        RECT 40.304 17.94 40.336 20.448 ;
  LAYER M3 ;
        RECT 40.24 17.94 40.272 20.448 ;
  LAYER M3 ;
        RECT 40.144 17.94 40.176 20.448 ;
  LAYER M1 ;
        RECT 42.559 17.976 42.561 20.412 ;
  LAYER M1 ;
        RECT 42.479 17.976 42.481 20.412 ;
  LAYER M1 ;
        RECT 42.399 17.976 42.401 20.412 ;
  LAYER M1 ;
        RECT 42.319 17.976 42.321 20.412 ;
  LAYER M1 ;
        RECT 42.239 17.976 42.241 20.412 ;
  LAYER M1 ;
        RECT 42.159 17.976 42.161 20.412 ;
  LAYER M1 ;
        RECT 42.079 17.976 42.081 20.412 ;
  LAYER M1 ;
        RECT 41.999 17.976 42.001 20.412 ;
  LAYER M1 ;
        RECT 41.919 17.976 41.921 20.412 ;
  LAYER M1 ;
        RECT 41.839 17.976 41.841 20.412 ;
  LAYER M1 ;
        RECT 41.759 17.976 41.761 20.412 ;
  LAYER M1 ;
        RECT 41.679 17.976 41.681 20.412 ;
  LAYER M1 ;
        RECT 41.599 17.976 41.601 20.412 ;
  LAYER M1 ;
        RECT 41.519 17.976 41.521 20.412 ;
  LAYER M1 ;
        RECT 41.439 17.976 41.441 20.412 ;
  LAYER M1 ;
        RECT 41.359 17.976 41.361 20.412 ;
  LAYER M1 ;
        RECT 41.279 17.976 41.281 20.412 ;
  LAYER M1 ;
        RECT 41.199 17.976 41.201 20.412 ;
  LAYER M1 ;
        RECT 41.119 17.976 41.121 20.412 ;
  LAYER M1 ;
        RECT 41.039 17.976 41.041 20.412 ;
  LAYER M1 ;
        RECT 40.959 17.976 40.961 20.412 ;
  LAYER M1 ;
        RECT 40.879 17.976 40.881 20.412 ;
  LAYER M1 ;
        RECT 40.799 17.976 40.801 20.412 ;
  LAYER M1 ;
        RECT 40.719 17.976 40.721 20.412 ;
  LAYER M1 ;
        RECT 40.639 17.976 40.641 20.412 ;
  LAYER M1 ;
        RECT 40.559 17.976 40.561 20.412 ;
  LAYER M1 ;
        RECT 40.479 17.976 40.481 20.412 ;
  LAYER M1 ;
        RECT 40.399 17.976 40.401 20.412 ;
  LAYER M1 ;
        RECT 40.319 17.976 40.321 20.412 ;
  LAYER M1 ;
        RECT 40.239 17.976 40.241 20.412 ;
  LAYER M2 ;
        RECT 40.16 17.975 42.56 17.977 ;
  LAYER M2 ;
        RECT 40.16 18.059 42.56 18.061 ;
  LAYER M2 ;
        RECT 40.16 18.143 42.56 18.145 ;
  LAYER M2 ;
        RECT 40.16 18.227 42.56 18.229 ;
  LAYER M2 ;
        RECT 40.16 18.311 42.56 18.313 ;
  LAYER M2 ;
        RECT 40.16 18.395 42.56 18.397 ;
  LAYER M2 ;
        RECT 40.16 18.479 42.56 18.481 ;
  LAYER M2 ;
        RECT 40.16 18.563 42.56 18.565 ;
  LAYER M2 ;
        RECT 40.16 18.647 42.56 18.649 ;
  LAYER M2 ;
        RECT 40.16 18.731 42.56 18.733 ;
  LAYER M2 ;
        RECT 40.16 18.815 42.56 18.817 ;
  LAYER M2 ;
        RECT 40.16 18.899 42.56 18.901 ;
  LAYER M2 ;
        RECT 40.16 18.9825 42.56 18.9845 ;
  LAYER M2 ;
        RECT 40.16 19.067 42.56 19.069 ;
  LAYER M2 ;
        RECT 40.16 19.151 42.56 19.153 ;
  LAYER M2 ;
        RECT 40.16 19.235 42.56 19.237 ;
  LAYER M2 ;
        RECT 40.16 19.319 42.56 19.321 ;
  LAYER M2 ;
        RECT 40.16 19.403 42.56 19.405 ;
  LAYER M2 ;
        RECT 40.16 19.487 42.56 19.489 ;
  LAYER M2 ;
        RECT 40.16 19.571 42.56 19.573 ;
  LAYER M2 ;
        RECT 40.16 19.655 42.56 19.657 ;
  LAYER M2 ;
        RECT 40.16 19.739 42.56 19.741 ;
  LAYER M2 ;
        RECT 40.16 19.823 42.56 19.825 ;
  LAYER M2 ;
        RECT 40.16 19.907 42.56 19.909 ;
  LAYER M2 ;
        RECT 40.16 19.991 42.56 19.993 ;
  LAYER M2 ;
        RECT 40.16 20.075 42.56 20.077 ;
  LAYER M2 ;
        RECT 40.16 20.159 42.56 20.161 ;
  LAYER M2 ;
        RECT 40.16 20.243 42.56 20.245 ;
  LAYER M2 ;
        RECT 40.16 20.327 42.56 20.329 ;
  LAYER M1 ;
        RECT 42.544 20.88 42.576 23.388 ;
  LAYER M1 ;
        RECT 42.48 20.88 42.512 23.388 ;
  LAYER M1 ;
        RECT 42.416 20.88 42.448 23.388 ;
  LAYER M1 ;
        RECT 42.352 20.88 42.384 23.388 ;
  LAYER M1 ;
        RECT 42.288 20.88 42.32 23.388 ;
  LAYER M1 ;
        RECT 42.224 20.88 42.256 23.388 ;
  LAYER M1 ;
        RECT 42.16 20.88 42.192 23.388 ;
  LAYER M1 ;
        RECT 42.096 20.88 42.128 23.388 ;
  LAYER M1 ;
        RECT 42.032 20.88 42.064 23.388 ;
  LAYER M1 ;
        RECT 41.968 20.88 42 23.388 ;
  LAYER M1 ;
        RECT 41.904 20.88 41.936 23.388 ;
  LAYER M1 ;
        RECT 41.84 20.88 41.872 23.388 ;
  LAYER M1 ;
        RECT 41.776 20.88 41.808 23.388 ;
  LAYER M1 ;
        RECT 41.712 20.88 41.744 23.388 ;
  LAYER M1 ;
        RECT 41.648 20.88 41.68 23.388 ;
  LAYER M1 ;
        RECT 41.584 20.88 41.616 23.388 ;
  LAYER M1 ;
        RECT 41.52 20.88 41.552 23.388 ;
  LAYER M1 ;
        RECT 41.456 20.88 41.488 23.388 ;
  LAYER M1 ;
        RECT 41.392 20.88 41.424 23.388 ;
  LAYER M1 ;
        RECT 41.328 20.88 41.36 23.388 ;
  LAYER M1 ;
        RECT 41.264 20.88 41.296 23.388 ;
  LAYER M1 ;
        RECT 41.2 20.88 41.232 23.388 ;
  LAYER M1 ;
        RECT 41.136 20.88 41.168 23.388 ;
  LAYER M1 ;
        RECT 41.072 20.88 41.104 23.388 ;
  LAYER M1 ;
        RECT 41.008 20.88 41.04 23.388 ;
  LAYER M1 ;
        RECT 40.944 20.88 40.976 23.388 ;
  LAYER M1 ;
        RECT 40.88 20.88 40.912 23.388 ;
  LAYER M1 ;
        RECT 40.816 20.88 40.848 23.388 ;
  LAYER M1 ;
        RECT 40.752 20.88 40.784 23.388 ;
  LAYER M1 ;
        RECT 40.688 20.88 40.72 23.388 ;
  LAYER M1 ;
        RECT 40.624 20.88 40.656 23.388 ;
  LAYER M1 ;
        RECT 40.56 20.88 40.592 23.388 ;
  LAYER M1 ;
        RECT 40.496 20.88 40.528 23.388 ;
  LAYER M1 ;
        RECT 40.432 20.88 40.464 23.388 ;
  LAYER M1 ;
        RECT 40.368 20.88 40.4 23.388 ;
  LAYER M1 ;
        RECT 40.304 20.88 40.336 23.388 ;
  LAYER M1 ;
        RECT 40.24 20.88 40.272 23.388 ;
  LAYER M2 ;
        RECT 40.124 20.964 42.596 20.996 ;
  LAYER M2 ;
        RECT 40.124 21.028 42.596 21.06 ;
  LAYER M2 ;
        RECT 40.124 21.092 42.596 21.124 ;
  LAYER M2 ;
        RECT 40.124 21.156 42.596 21.188 ;
  LAYER M2 ;
        RECT 40.124 21.22 42.596 21.252 ;
  LAYER M2 ;
        RECT 40.124 21.284 42.596 21.316 ;
  LAYER M2 ;
        RECT 40.124 21.348 42.596 21.38 ;
  LAYER M2 ;
        RECT 40.124 21.412 42.596 21.444 ;
  LAYER M2 ;
        RECT 40.124 21.476 42.596 21.508 ;
  LAYER M2 ;
        RECT 40.124 21.54 42.596 21.572 ;
  LAYER M2 ;
        RECT 40.124 21.604 42.596 21.636 ;
  LAYER M2 ;
        RECT 40.124 21.668 42.596 21.7 ;
  LAYER M2 ;
        RECT 40.124 21.732 42.596 21.764 ;
  LAYER M2 ;
        RECT 40.124 21.796 42.596 21.828 ;
  LAYER M2 ;
        RECT 40.124 21.86 42.596 21.892 ;
  LAYER M2 ;
        RECT 40.124 21.924 42.596 21.956 ;
  LAYER M2 ;
        RECT 40.124 21.988 42.596 22.02 ;
  LAYER M2 ;
        RECT 40.124 22.052 42.596 22.084 ;
  LAYER M2 ;
        RECT 40.124 22.116 42.596 22.148 ;
  LAYER M2 ;
        RECT 40.124 22.18 42.596 22.212 ;
  LAYER M2 ;
        RECT 40.124 22.244 42.596 22.276 ;
  LAYER M2 ;
        RECT 40.124 22.308 42.596 22.34 ;
  LAYER M2 ;
        RECT 40.124 22.372 42.596 22.404 ;
  LAYER M2 ;
        RECT 40.124 22.436 42.596 22.468 ;
  LAYER M2 ;
        RECT 40.124 22.5 42.596 22.532 ;
  LAYER M2 ;
        RECT 40.124 22.564 42.596 22.596 ;
  LAYER M2 ;
        RECT 40.124 22.628 42.596 22.66 ;
  LAYER M2 ;
        RECT 40.124 22.692 42.596 22.724 ;
  LAYER M2 ;
        RECT 40.124 22.756 42.596 22.788 ;
  LAYER M2 ;
        RECT 40.124 22.82 42.596 22.852 ;
  LAYER M2 ;
        RECT 40.124 22.884 42.596 22.916 ;
  LAYER M2 ;
        RECT 40.124 22.948 42.596 22.98 ;
  LAYER M2 ;
        RECT 40.124 23.012 42.596 23.044 ;
  LAYER M2 ;
        RECT 40.124 23.076 42.596 23.108 ;
  LAYER M2 ;
        RECT 40.124 23.14 42.596 23.172 ;
  LAYER M2 ;
        RECT 40.124 23.204 42.596 23.236 ;
  LAYER M3 ;
        RECT 42.544 20.88 42.576 23.388 ;
  LAYER M3 ;
        RECT 42.48 20.88 42.512 23.388 ;
  LAYER M3 ;
        RECT 42.416 20.88 42.448 23.388 ;
  LAYER M3 ;
        RECT 42.352 20.88 42.384 23.388 ;
  LAYER M3 ;
        RECT 42.288 20.88 42.32 23.388 ;
  LAYER M3 ;
        RECT 42.224 20.88 42.256 23.388 ;
  LAYER M3 ;
        RECT 42.16 20.88 42.192 23.388 ;
  LAYER M3 ;
        RECT 42.096 20.88 42.128 23.388 ;
  LAYER M3 ;
        RECT 42.032 20.88 42.064 23.388 ;
  LAYER M3 ;
        RECT 41.968 20.88 42 23.388 ;
  LAYER M3 ;
        RECT 41.904 20.88 41.936 23.388 ;
  LAYER M3 ;
        RECT 41.84 20.88 41.872 23.388 ;
  LAYER M3 ;
        RECT 41.776 20.88 41.808 23.388 ;
  LAYER M3 ;
        RECT 41.712 20.88 41.744 23.388 ;
  LAYER M3 ;
        RECT 41.648 20.88 41.68 23.388 ;
  LAYER M3 ;
        RECT 41.584 20.88 41.616 23.388 ;
  LAYER M3 ;
        RECT 41.52 20.88 41.552 23.388 ;
  LAYER M3 ;
        RECT 41.456 20.88 41.488 23.388 ;
  LAYER M3 ;
        RECT 41.392 20.88 41.424 23.388 ;
  LAYER M3 ;
        RECT 41.328 20.88 41.36 23.388 ;
  LAYER M3 ;
        RECT 41.264 20.88 41.296 23.388 ;
  LAYER M3 ;
        RECT 41.2 20.88 41.232 23.388 ;
  LAYER M3 ;
        RECT 41.136 20.88 41.168 23.388 ;
  LAYER M3 ;
        RECT 41.072 20.88 41.104 23.388 ;
  LAYER M3 ;
        RECT 41.008 20.88 41.04 23.388 ;
  LAYER M3 ;
        RECT 40.944 20.88 40.976 23.388 ;
  LAYER M3 ;
        RECT 40.88 20.88 40.912 23.388 ;
  LAYER M3 ;
        RECT 40.816 20.88 40.848 23.388 ;
  LAYER M3 ;
        RECT 40.752 20.88 40.784 23.388 ;
  LAYER M3 ;
        RECT 40.688 20.88 40.72 23.388 ;
  LAYER M3 ;
        RECT 40.624 20.88 40.656 23.388 ;
  LAYER M3 ;
        RECT 40.56 20.88 40.592 23.388 ;
  LAYER M3 ;
        RECT 40.496 20.88 40.528 23.388 ;
  LAYER M3 ;
        RECT 40.432 20.88 40.464 23.388 ;
  LAYER M3 ;
        RECT 40.368 20.88 40.4 23.388 ;
  LAYER M3 ;
        RECT 40.304 20.88 40.336 23.388 ;
  LAYER M3 ;
        RECT 40.24 20.88 40.272 23.388 ;
  LAYER M3 ;
        RECT 40.144 20.88 40.176 23.388 ;
  LAYER M1 ;
        RECT 42.559 20.916 42.561 23.352 ;
  LAYER M1 ;
        RECT 42.479 20.916 42.481 23.352 ;
  LAYER M1 ;
        RECT 42.399 20.916 42.401 23.352 ;
  LAYER M1 ;
        RECT 42.319 20.916 42.321 23.352 ;
  LAYER M1 ;
        RECT 42.239 20.916 42.241 23.352 ;
  LAYER M1 ;
        RECT 42.159 20.916 42.161 23.352 ;
  LAYER M1 ;
        RECT 42.079 20.916 42.081 23.352 ;
  LAYER M1 ;
        RECT 41.999 20.916 42.001 23.352 ;
  LAYER M1 ;
        RECT 41.919 20.916 41.921 23.352 ;
  LAYER M1 ;
        RECT 41.839 20.916 41.841 23.352 ;
  LAYER M1 ;
        RECT 41.759 20.916 41.761 23.352 ;
  LAYER M1 ;
        RECT 41.679 20.916 41.681 23.352 ;
  LAYER M1 ;
        RECT 41.599 20.916 41.601 23.352 ;
  LAYER M1 ;
        RECT 41.519 20.916 41.521 23.352 ;
  LAYER M1 ;
        RECT 41.439 20.916 41.441 23.352 ;
  LAYER M1 ;
        RECT 41.359 20.916 41.361 23.352 ;
  LAYER M1 ;
        RECT 41.279 20.916 41.281 23.352 ;
  LAYER M1 ;
        RECT 41.199 20.916 41.201 23.352 ;
  LAYER M1 ;
        RECT 41.119 20.916 41.121 23.352 ;
  LAYER M1 ;
        RECT 41.039 20.916 41.041 23.352 ;
  LAYER M1 ;
        RECT 40.959 20.916 40.961 23.352 ;
  LAYER M1 ;
        RECT 40.879 20.916 40.881 23.352 ;
  LAYER M1 ;
        RECT 40.799 20.916 40.801 23.352 ;
  LAYER M1 ;
        RECT 40.719 20.916 40.721 23.352 ;
  LAYER M1 ;
        RECT 40.639 20.916 40.641 23.352 ;
  LAYER M1 ;
        RECT 40.559 20.916 40.561 23.352 ;
  LAYER M1 ;
        RECT 40.479 20.916 40.481 23.352 ;
  LAYER M1 ;
        RECT 40.399 20.916 40.401 23.352 ;
  LAYER M1 ;
        RECT 40.319 20.916 40.321 23.352 ;
  LAYER M1 ;
        RECT 40.239 20.916 40.241 23.352 ;
  LAYER M2 ;
        RECT 40.16 20.915 42.56 20.917 ;
  LAYER M2 ;
        RECT 40.16 20.999 42.56 21.001 ;
  LAYER M2 ;
        RECT 40.16 21.083 42.56 21.085 ;
  LAYER M2 ;
        RECT 40.16 21.167 42.56 21.169 ;
  LAYER M2 ;
        RECT 40.16 21.251 42.56 21.253 ;
  LAYER M2 ;
        RECT 40.16 21.335 42.56 21.337 ;
  LAYER M2 ;
        RECT 40.16 21.419 42.56 21.421 ;
  LAYER M2 ;
        RECT 40.16 21.503 42.56 21.505 ;
  LAYER M2 ;
        RECT 40.16 21.587 42.56 21.589 ;
  LAYER M2 ;
        RECT 40.16 21.671 42.56 21.673 ;
  LAYER M2 ;
        RECT 40.16 21.755 42.56 21.757 ;
  LAYER M2 ;
        RECT 40.16 21.839 42.56 21.841 ;
  LAYER M2 ;
        RECT 40.16 21.9225 42.56 21.9245 ;
  LAYER M2 ;
        RECT 40.16 22.007 42.56 22.009 ;
  LAYER M2 ;
        RECT 40.16 22.091 42.56 22.093 ;
  LAYER M2 ;
        RECT 40.16 22.175 42.56 22.177 ;
  LAYER M2 ;
        RECT 40.16 22.259 42.56 22.261 ;
  LAYER M2 ;
        RECT 40.16 22.343 42.56 22.345 ;
  LAYER M2 ;
        RECT 40.16 22.427 42.56 22.429 ;
  LAYER M2 ;
        RECT 40.16 22.511 42.56 22.513 ;
  LAYER M2 ;
        RECT 40.16 22.595 42.56 22.597 ;
  LAYER M2 ;
        RECT 40.16 22.679 42.56 22.681 ;
  LAYER M2 ;
        RECT 40.16 22.763 42.56 22.765 ;
  LAYER M2 ;
        RECT 40.16 22.847 42.56 22.849 ;
  LAYER M2 ;
        RECT 40.16 22.931 42.56 22.933 ;
  LAYER M2 ;
        RECT 40.16 23.015 42.56 23.017 ;
  LAYER M2 ;
        RECT 40.16 23.099 42.56 23.101 ;
  LAYER M2 ;
        RECT 40.16 23.183 42.56 23.185 ;
  LAYER M2 ;
        RECT 40.16 23.267 42.56 23.269 ;
  LAYER M1 ;
        RECT 42.544 23.82 42.576 26.328 ;
  LAYER M1 ;
        RECT 42.48 23.82 42.512 26.328 ;
  LAYER M1 ;
        RECT 42.416 23.82 42.448 26.328 ;
  LAYER M1 ;
        RECT 42.352 23.82 42.384 26.328 ;
  LAYER M1 ;
        RECT 42.288 23.82 42.32 26.328 ;
  LAYER M1 ;
        RECT 42.224 23.82 42.256 26.328 ;
  LAYER M1 ;
        RECT 42.16 23.82 42.192 26.328 ;
  LAYER M1 ;
        RECT 42.096 23.82 42.128 26.328 ;
  LAYER M1 ;
        RECT 42.032 23.82 42.064 26.328 ;
  LAYER M1 ;
        RECT 41.968 23.82 42 26.328 ;
  LAYER M1 ;
        RECT 41.904 23.82 41.936 26.328 ;
  LAYER M1 ;
        RECT 41.84 23.82 41.872 26.328 ;
  LAYER M1 ;
        RECT 41.776 23.82 41.808 26.328 ;
  LAYER M1 ;
        RECT 41.712 23.82 41.744 26.328 ;
  LAYER M1 ;
        RECT 41.648 23.82 41.68 26.328 ;
  LAYER M1 ;
        RECT 41.584 23.82 41.616 26.328 ;
  LAYER M1 ;
        RECT 41.52 23.82 41.552 26.328 ;
  LAYER M1 ;
        RECT 41.456 23.82 41.488 26.328 ;
  LAYER M1 ;
        RECT 41.392 23.82 41.424 26.328 ;
  LAYER M1 ;
        RECT 41.328 23.82 41.36 26.328 ;
  LAYER M1 ;
        RECT 41.264 23.82 41.296 26.328 ;
  LAYER M1 ;
        RECT 41.2 23.82 41.232 26.328 ;
  LAYER M1 ;
        RECT 41.136 23.82 41.168 26.328 ;
  LAYER M1 ;
        RECT 41.072 23.82 41.104 26.328 ;
  LAYER M1 ;
        RECT 41.008 23.82 41.04 26.328 ;
  LAYER M1 ;
        RECT 40.944 23.82 40.976 26.328 ;
  LAYER M1 ;
        RECT 40.88 23.82 40.912 26.328 ;
  LAYER M1 ;
        RECT 40.816 23.82 40.848 26.328 ;
  LAYER M1 ;
        RECT 40.752 23.82 40.784 26.328 ;
  LAYER M1 ;
        RECT 40.688 23.82 40.72 26.328 ;
  LAYER M1 ;
        RECT 40.624 23.82 40.656 26.328 ;
  LAYER M1 ;
        RECT 40.56 23.82 40.592 26.328 ;
  LAYER M1 ;
        RECT 40.496 23.82 40.528 26.328 ;
  LAYER M1 ;
        RECT 40.432 23.82 40.464 26.328 ;
  LAYER M1 ;
        RECT 40.368 23.82 40.4 26.328 ;
  LAYER M1 ;
        RECT 40.304 23.82 40.336 26.328 ;
  LAYER M1 ;
        RECT 40.24 23.82 40.272 26.328 ;
  LAYER M2 ;
        RECT 40.124 23.904 42.596 23.936 ;
  LAYER M2 ;
        RECT 40.124 23.968 42.596 24 ;
  LAYER M2 ;
        RECT 40.124 24.032 42.596 24.064 ;
  LAYER M2 ;
        RECT 40.124 24.096 42.596 24.128 ;
  LAYER M2 ;
        RECT 40.124 24.16 42.596 24.192 ;
  LAYER M2 ;
        RECT 40.124 24.224 42.596 24.256 ;
  LAYER M2 ;
        RECT 40.124 24.288 42.596 24.32 ;
  LAYER M2 ;
        RECT 40.124 24.352 42.596 24.384 ;
  LAYER M2 ;
        RECT 40.124 24.416 42.596 24.448 ;
  LAYER M2 ;
        RECT 40.124 24.48 42.596 24.512 ;
  LAYER M2 ;
        RECT 40.124 24.544 42.596 24.576 ;
  LAYER M2 ;
        RECT 40.124 24.608 42.596 24.64 ;
  LAYER M2 ;
        RECT 40.124 24.672 42.596 24.704 ;
  LAYER M2 ;
        RECT 40.124 24.736 42.596 24.768 ;
  LAYER M2 ;
        RECT 40.124 24.8 42.596 24.832 ;
  LAYER M2 ;
        RECT 40.124 24.864 42.596 24.896 ;
  LAYER M2 ;
        RECT 40.124 24.928 42.596 24.96 ;
  LAYER M2 ;
        RECT 40.124 24.992 42.596 25.024 ;
  LAYER M2 ;
        RECT 40.124 25.056 42.596 25.088 ;
  LAYER M2 ;
        RECT 40.124 25.12 42.596 25.152 ;
  LAYER M2 ;
        RECT 40.124 25.184 42.596 25.216 ;
  LAYER M2 ;
        RECT 40.124 25.248 42.596 25.28 ;
  LAYER M2 ;
        RECT 40.124 25.312 42.596 25.344 ;
  LAYER M2 ;
        RECT 40.124 25.376 42.596 25.408 ;
  LAYER M2 ;
        RECT 40.124 25.44 42.596 25.472 ;
  LAYER M2 ;
        RECT 40.124 25.504 42.596 25.536 ;
  LAYER M2 ;
        RECT 40.124 25.568 42.596 25.6 ;
  LAYER M2 ;
        RECT 40.124 25.632 42.596 25.664 ;
  LAYER M2 ;
        RECT 40.124 25.696 42.596 25.728 ;
  LAYER M2 ;
        RECT 40.124 25.76 42.596 25.792 ;
  LAYER M2 ;
        RECT 40.124 25.824 42.596 25.856 ;
  LAYER M2 ;
        RECT 40.124 25.888 42.596 25.92 ;
  LAYER M2 ;
        RECT 40.124 25.952 42.596 25.984 ;
  LAYER M2 ;
        RECT 40.124 26.016 42.596 26.048 ;
  LAYER M2 ;
        RECT 40.124 26.08 42.596 26.112 ;
  LAYER M2 ;
        RECT 40.124 26.144 42.596 26.176 ;
  LAYER M3 ;
        RECT 42.544 23.82 42.576 26.328 ;
  LAYER M3 ;
        RECT 42.48 23.82 42.512 26.328 ;
  LAYER M3 ;
        RECT 42.416 23.82 42.448 26.328 ;
  LAYER M3 ;
        RECT 42.352 23.82 42.384 26.328 ;
  LAYER M3 ;
        RECT 42.288 23.82 42.32 26.328 ;
  LAYER M3 ;
        RECT 42.224 23.82 42.256 26.328 ;
  LAYER M3 ;
        RECT 42.16 23.82 42.192 26.328 ;
  LAYER M3 ;
        RECT 42.096 23.82 42.128 26.328 ;
  LAYER M3 ;
        RECT 42.032 23.82 42.064 26.328 ;
  LAYER M3 ;
        RECT 41.968 23.82 42 26.328 ;
  LAYER M3 ;
        RECT 41.904 23.82 41.936 26.328 ;
  LAYER M3 ;
        RECT 41.84 23.82 41.872 26.328 ;
  LAYER M3 ;
        RECT 41.776 23.82 41.808 26.328 ;
  LAYER M3 ;
        RECT 41.712 23.82 41.744 26.328 ;
  LAYER M3 ;
        RECT 41.648 23.82 41.68 26.328 ;
  LAYER M3 ;
        RECT 41.584 23.82 41.616 26.328 ;
  LAYER M3 ;
        RECT 41.52 23.82 41.552 26.328 ;
  LAYER M3 ;
        RECT 41.456 23.82 41.488 26.328 ;
  LAYER M3 ;
        RECT 41.392 23.82 41.424 26.328 ;
  LAYER M3 ;
        RECT 41.328 23.82 41.36 26.328 ;
  LAYER M3 ;
        RECT 41.264 23.82 41.296 26.328 ;
  LAYER M3 ;
        RECT 41.2 23.82 41.232 26.328 ;
  LAYER M3 ;
        RECT 41.136 23.82 41.168 26.328 ;
  LAYER M3 ;
        RECT 41.072 23.82 41.104 26.328 ;
  LAYER M3 ;
        RECT 41.008 23.82 41.04 26.328 ;
  LAYER M3 ;
        RECT 40.944 23.82 40.976 26.328 ;
  LAYER M3 ;
        RECT 40.88 23.82 40.912 26.328 ;
  LAYER M3 ;
        RECT 40.816 23.82 40.848 26.328 ;
  LAYER M3 ;
        RECT 40.752 23.82 40.784 26.328 ;
  LAYER M3 ;
        RECT 40.688 23.82 40.72 26.328 ;
  LAYER M3 ;
        RECT 40.624 23.82 40.656 26.328 ;
  LAYER M3 ;
        RECT 40.56 23.82 40.592 26.328 ;
  LAYER M3 ;
        RECT 40.496 23.82 40.528 26.328 ;
  LAYER M3 ;
        RECT 40.432 23.82 40.464 26.328 ;
  LAYER M3 ;
        RECT 40.368 23.82 40.4 26.328 ;
  LAYER M3 ;
        RECT 40.304 23.82 40.336 26.328 ;
  LAYER M3 ;
        RECT 40.24 23.82 40.272 26.328 ;
  LAYER M3 ;
        RECT 40.144 23.82 40.176 26.328 ;
  LAYER M1 ;
        RECT 42.559 23.856 42.561 26.292 ;
  LAYER M1 ;
        RECT 42.479 23.856 42.481 26.292 ;
  LAYER M1 ;
        RECT 42.399 23.856 42.401 26.292 ;
  LAYER M1 ;
        RECT 42.319 23.856 42.321 26.292 ;
  LAYER M1 ;
        RECT 42.239 23.856 42.241 26.292 ;
  LAYER M1 ;
        RECT 42.159 23.856 42.161 26.292 ;
  LAYER M1 ;
        RECT 42.079 23.856 42.081 26.292 ;
  LAYER M1 ;
        RECT 41.999 23.856 42.001 26.292 ;
  LAYER M1 ;
        RECT 41.919 23.856 41.921 26.292 ;
  LAYER M1 ;
        RECT 41.839 23.856 41.841 26.292 ;
  LAYER M1 ;
        RECT 41.759 23.856 41.761 26.292 ;
  LAYER M1 ;
        RECT 41.679 23.856 41.681 26.292 ;
  LAYER M1 ;
        RECT 41.599 23.856 41.601 26.292 ;
  LAYER M1 ;
        RECT 41.519 23.856 41.521 26.292 ;
  LAYER M1 ;
        RECT 41.439 23.856 41.441 26.292 ;
  LAYER M1 ;
        RECT 41.359 23.856 41.361 26.292 ;
  LAYER M1 ;
        RECT 41.279 23.856 41.281 26.292 ;
  LAYER M1 ;
        RECT 41.199 23.856 41.201 26.292 ;
  LAYER M1 ;
        RECT 41.119 23.856 41.121 26.292 ;
  LAYER M1 ;
        RECT 41.039 23.856 41.041 26.292 ;
  LAYER M1 ;
        RECT 40.959 23.856 40.961 26.292 ;
  LAYER M1 ;
        RECT 40.879 23.856 40.881 26.292 ;
  LAYER M1 ;
        RECT 40.799 23.856 40.801 26.292 ;
  LAYER M1 ;
        RECT 40.719 23.856 40.721 26.292 ;
  LAYER M1 ;
        RECT 40.639 23.856 40.641 26.292 ;
  LAYER M1 ;
        RECT 40.559 23.856 40.561 26.292 ;
  LAYER M1 ;
        RECT 40.479 23.856 40.481 26.292 ;
  LAYER M1 ;
        RECT 40.399 23.856 40.401 26.292 ;
  LAYER M1 ;
        RECT 40.319 23.856 40.321 26.292 ;
  LAYER M1 ;
        RECT 40.239 23.856 40.241 26.292 ;
  LAYER M2 ;
        RECT 40.16 23.855 42.56 23.857 ;
  LAYER M2 ;
        RECT 40.16 23.939 42.56 23.941 ;
  LAYER M2 ;
        RECT 40.16 24.023 42.56 24.025 ;
  LAYER M2 ;
        RECT 40.16 24.107 42.56 24.109 ;
  LAYER M2 ;
        RECT 40.16 24.191 42.56 24.193 ;
  LAYER M2 ;
        RECT 40.16 24.275 42.56 24.277 ;
  LAYER M2 ;
        RECT 40.16 24.359 42.56 24.361 ;
  LAYER M2 ;
        RECT 40.16 24.443 42.56 24.445 ;
  LAYER M2 ;
        RECT 40.16 24.527 42.56 24.529 ;
  LAYER M2 ;
        RECT 40.16 24.611 42.56 24.613 ;
  LAYER M2 ;
        RECT 40.16 24.695 42.56 24.697 ;
  LAYER M2 ;
        RECT 40.16 24.779 42.56 24.781 ;
  LAYER M2 ;
        RECT 40.16 24.8625 42.56 24.8645 ;
  LAYER M2 ;
        RECT 40.16 24.947 42.56 24.949 ;
  LAYER M2 ;
        RECT 40.16 25.031 42.56 25.033 ;
  LAYER M2 ;
        RECT 40.16 25.115 42.56 25.117 ;
  LAYER M2 ;
        RECT 40.16 25.199 42.56 25.201 ;
  LAYER M2 ;
        RECT 40.16 25.283 42.56 25.285 ;
  LAYER M2 ;
        RECT 40.16 25.367 42.56 25.369 ;
  LAYER M2 ;
        RECT 40.16 25.451 42.56 25.453 ;
  LAYER M2 ;
        RECT 40.16 25.535 42.56 25.537 ;
  LAYER M2 ;
        RECT 40.16 25.619 42.56 25.621 ;
  LAYER M2 ;
        RECT 40.16 25.703 42.56 25.705 ;
  LAYER M2 ;
        RECT 40.16 25.787 42.56 25.789 ;
  LAYER M2 ;
        RECT 40.16 25.871 42.56 25.873 ;
  LAYER M2 ;
        RECT 40.16 25.955 42.56 25.957 ;
  LAYER M2 ;
        RECT 40.16 26.039 42.56 26.041 ;
  LAYER M2 ;
        RECT 40.16 26.123 42.56 26.125 ;
  LAYER M2 ;
        RECT 40.16 26.207 42.56 26.209 ;
  LAYER M1 ;
        RECT 42.544 26.76 42.576 29.268 ;
  LAYER M1 ;
        RECT 42.48 26.76 42.512 29.268 ;
  LAYER M1 ;
        RECT 42.416 26.76 42.448 29.268 ;
  LAYER M1 ;
        RECT 42.352 26.76 42.384 29.268 ;
  LAYER M1 ;
        RECT 42.288 26.76 42.32 29.268 ;
  LAYER M1 ;
        RECT 42.224 26.76 42.256 29.268 ;
  LAYER M1 ;
        RECT 42.16 26.76 42.192 29.268 ;
  LAYER M1 ;
        RECT 42.096 26.76 42.128 29.268 ;
  LAYER M1 ;
        RECT 42.032 26.76 42.064 29.268 ;
  LAYER M1 ;
        RECT 41.968 26.76 42 29.268 ;
  LAYER M1 ;
        RECT 41.904 26.76 41.936 29.268 ;
  LAYER M1 ;
        RECT 41.84 26.76 41.872 29.268 ;
  LAYER M1 ;
        RECT 41.776 26.76 41.808 29.268 ;
  LAYER M1 ;
        RECT 41.712 26.76 41.744 29.268 ;
  LAYER M1 ;
        RECT 41.648 26.76 41.68 29.268 ;
  LAYER M1 ;
        RECT 41.584 26.76 41.616 29.268 ;
  LAYER M1 ;
        RECT 41.52 26.76 41.552 29.268 ;
  LAYER M1 ;
        RECT 41.456 26.76 41.488 29.268 ;
  LAYER M1 ;
        RECT 41.392 26.76 41.424 29.268 ;
  LAYER M1 ;
        RECT 41.328 26.76 41.36 29.268 ;
  LAYER M1 ;
        RECT 41.264 26.76 41.296 29.268 ;
  LAYER M1 ;
        RECT 41.2 26.76 41.232 29.268 ;
  LAYER M1 ;
        RECT 41.136 26.76 41.168 29.268 ;
  LAYER M1 ;
        RECT 41.072 26.76 41.104 29.268 ;
  LAYER M1 ;
        RECT 41.008 26.76 41.04 29.268 ;
  LAYER M1 ;
        RECT 40.944 26.76 40.976 29.268 ;
  LAYER M1 ;
        RECT 40.88 26.76 40.912 29.268 ;
  LAYER M1 ;
        RECT 40.816 26.76 40.848 29.268 ;
  LAYER M1 ;
        RECT 40.752 26.76 40.784 29.268 ;
  LAYER M1 ;
        RECT 40.688 26.76 40.72 29.268 ;
  LAYER M1 ;
        RECT 40.624 26.76 40.656 29.268 ;
  LAYER M1 ;
        RECT 40.56 26.76 40.592 29.268 ;
  LAYER M1 ;
        RECT 40.496 26.76 40.528 29.268 ;
  LAYER M1 ;
        RECT 40.432 26.76 40.464 29.268 ;
  LAYER M1 ;
        RECT 40.368 26.76 40.4 29.268 ;
  LAYER M1 ;
        RECT 40.304 26.76 40.336 29.268 ;
  LAYER M1 ;
        RECT 40.24 26.76 40.272 29.268 ;
  LAYER M2 ;
        RECT 40.124 26.844 42.596 26.876 ;
  LAYER M2 ;
        RECT 40.124 26.908 42.596 26.94 ;
  LAYER M2 ;
        RECT 40.124 26.972 42.596 27.004 ;
  LAYER M2 ;
        RECT 40.124 27.036 42.596 27.068 ;
  LAYER M2 ;
        RECT 40.124 27.1 42.596 27.132 ;
  LAYER M2 ;
        RECT 40.124 27.164 42.596 27.196 ;
  LAYER M2 ;
        RECT 40.124 27.228 42.596 27.26 ;
  LAYER M2 ;
        RECT 40.124 27.292 42.596 27.324 ;
  LAYER M2 ;
        RECT 40.124 27.356 42.596 27.388 ;
  LAYER M2 ;
        RECT 40.124 27.42 42.596 27.452 ;
  LAYER M2 ;
        RECT 40.124 27.484 42.596 27.516 ;
  LAYER M2 ;
        RECT 40.124 27.548 42.596 27.58 ;
  LAYER M2 ;
        RECT 40.124 27.612 42.596 27.644 ;
  LAYER M2 ;
        RECT 40.124 27.676 42.596 27.708 ;
  LAYER M2 ;
        RECT 40.124 27.74 42.596 27.772 ;
  LAYER M2 ;
        RECT 40.124 27.804 42.596 27.836 ;
  LAYER M2 ;
        RECT 40.124 27.868 42.596 27.9 ;
  LAYER M2 ;
        RECT 40.124 27.932 42.596 27.964 ;
  LAYER M2 ;
        RECT 40.124 27.996 42.596 28.028 ;
  LAYER M2 ;
        RECT 40.124 28.06 42.596 28.092 ;
  LAYER M2 ;
        RECT 40.124 28.124 42.596 28.156 ;
  LAYER M2 ;
        RECT 40.124 28.188 42.596 28.22 ;
  LAYER M2 ;
        RECT 40.124 28.252 42.596 28.284 ;
  LAYER M2 ;
        RECT 40.124 28.316 42.596 28.348 ;
  LAYER M2 ;
        RECT 40.124 28.38 42.596 28.412 ;
  LAYER M2 ;
        RECT 40.124 28.444 42.596 28.476 ;
  LAYER M2 ;
        RECT 40.124 28.508 42.596 28.54 ;
  LAYER M2 ;
        RECT 40.124 28.572 42.596 28.604 ;
  LAYER M2 ;
        RECT 40.124 28.636 42.596 28.668 ;
  LAYER M2 ;
        RECT 40.124 28.7 42.596 28.732 ;
  LAYER M2 ;
        RECT 40.124 28.764 42.596 28.796 ;
  LAYER M2 ;
        RECT 40.124 28.828 42.596 28.86 ;
  LAYER M2 ;
        RECT 40.124 28.892 42.596 28.924 ;
  LAYER M2 ;
        RECT 40.124 28.956 42.596 28.988 ;
  LAYER M2 ;
        RECT 40.124 29.02 42.596 29.052 ;
  LAYER M2 ;
        RECT 40.124 29.084 42.596 29.116 ;
  LAYER M3 ;
        RECT 42.544 26.76 42.576 29.268 ;
  LAYER M3 ;
        RECT 42.48 26.76 42.512 29.268 ;
  LAYER M3 ;
        RECT 42.416 26.76 42.448 29.268 ;
  LAYER M3 ;
        RECT 42.352 26.76 42.384 29.268 ;
  LAYER M3 ;
        RECT 42.288 26.76 42.32 29.268 ;
  LAYER M3 ;
        RECT 42.224 26.76 42.256 29.268 ;
  LAYER M3 ;
        RECT 42.16 26.76 42.192 29.268 ;
  LAYER M3 ;
        RECT 42.096 26.76 42.128 29.268 ;
  LAYER M3 ;
        RECT 42.032 26.76 42.064 29.268 ;
  LAYER M3 ;
        RECT 41.968 26.76 42 29.268 ;
  LAYER M3 ;
        RECT 41.904 26.76 41.936 29.268 ;
  LAYER M3 ;
        RECT 41.84 26.76 41.872 29.268 ;
  LAYER M3 ;
        RECT 41.776 26.76 41.808 29.268 ;
  LAYER M3 ;
        RECT 41.712 26.76 41.744 29.268 ;
  LAYER M3 ;
        RECT 41.648 26.76 41.68 29.268 ;
  LAYER M3 ;
        RECT 41.584 26.76 41.616 29.268 ;
  LAYER M3 ;
        RECT 41.52 26.76 41.552 29.268 ;
  LAYER M3 ;
        RECT 41.456 26.76 41.488 29.268 ;
  LAYER M3 ;
        RECT 41.392 26.76 41.424 29.268 ;
  LAYER M3 ;
        RECT 41.328 26.76 41.36 29.268 ;
  LAYER M3 ;
        RECT 41.264 26.76 41.296 29.268 ;
  LAYER M3 ;
        RECT 41.2 26.76 41.232 29.268 ;
  LAYER M3 ;
        RECT 41.136 26.76 41.168 29.268 ;
  LAYER M3 ;
        RECT 41.072 26.76 41.104 29.268 ;
  LAYER M3 ;
        RECT 41.008 26.76 41.04 29.268 ;
  LAYER M3 ;
        RECT 40.944 26.76 40.976 29.268 ;
  LAYER M3 ;
        RECT 40.88 26.76 40.912 29.268 ;
  LAYER M3 ;
        RECT 40.816 26.76 40.848 29.268 ;
  LAYER M3 ;
        RECT 40.752 26.76 40.784 29.268 ;
  LAYER M3 ;
        RECT 40.688 26.76 40.72 29.268 ;
  LAYER M3 ;
        RECT 40.624 26.76 40.656 29.268 ;
  LAYER M3 ;
        RECT 40.56 26.76 40.592 29.268 ;
  LAYER M3 ;
        RECT 40.496 26.76 40.528 29.268 ;
  LAYER M3 ;
        RECT 40.432 26.76 40.464 29.268 ;
  LAYER M3 ;
        RECT 40.368 26.76 40.4 29.268 ;
  LAYER M3 ;
        RECT 40.304 26.76 40.336 29.268 ;
  LAYER M3 ;
        RECT 40.24 26.76 40.272 29.268 ;
  LAYER M3 ;
        RECT 40.144 26.76 40.176 29.268 ;
  LAYER M1 ;
        RECT 42.559 26.796 42.561 29.232 ;
  LAYER M1 ;
        RECT 42.479 26.796 42.481 29.232 ;
  LAYER M1 ;
        RECT 42.399 26.796 42.401 29.232 ;
  LAYER M1 ;
        RECT 42.319 26.796 42.321 29.232 ;
  LAYER M1 ;
        RECT 42.239 26.796 42.241 29.232 ;
  LAYER M1 ;
        RECT 42.159 26.796 42.161 29.232 ;
  LAYER M1 ;
        RECT 42.079 26.796 42.081 29.232 ;
  LAYER M1 ;
        RECT 41.999 26.796 42.001 29.232 ;
  LAYER M1 ;
        RECT 41.919 26.796 41.921 29.232 ;
  LAYER M1 ;
        RECT 41.839 26.796 41.841 29.232 ;
  LAYER M1 ;
        RECT 41.759 26.796 41.761 29.232 ;
  LAYER M1 ;
        RECT 41.679 26.796 41.681 29.232 ;
  LAYER M1 ;
        RECT 41.599 26.796 41.601 29.232 ;
  LAYER M1 ;
        RECT 41.519 26.796 41.521 29.232 ;
  LAYER M1 ;
        RECT 41.439 26.796 41.441 29.232 ;
  LAYER M1 ;
        RECT 41.359 26.796 41.361 29.232 ;
  LAYER M1 ;
        RECT 41.279 26.796 41.281 29.232 ;
  LAYER M1 ;
        RECT 41.199 26.796 41.201 29.232 ;
  LAYER M1 ;
        RECT 41.119 26.796 41.121 29.232 ;
  LAYER M1 ;
        RECT 41.039 26.796 41.041 29.232 ;
  LAYER M1 ;
        RECT 40.959 26.796 40.961 29.232 ;
  LAYER M1 ;
        RECT 40.879 26.796 40.881 29.232 ;
  LAYER M1 ;
        RECT 40.799 26.796 40.801 29.232 ;
  LAYER M1 ;
        RECT 40.719 26.796 40.721 29.232 ;
  LAYER M1 ;
        RECT 40.639 26.796 40.641 29.232 ;
  LAYER M1 ;
        RECT 40.559 26.796 40.561 29.232 ;
  LAYER M1 ;
        RECT 40.479 26.796 40.481 29.232 ;
  LAYER M1 ;
        RECT 40.399 26.796 40.401 29.232 ;
  LAYER M1 ;
        RECT 40.319 26.796 40.321 29.232 ;
  LAYER M1 ;
        RECT 40.239 26.796 40.241 29.232 ;
  LAYER M2 ;
        RECT 40.16 26.795 42.56 26.797 ;
  LAYER M2 ;
        RECT 40.16 26.879 42.56 26.881 ;
  LAYER M2 ;
        RECT 40.16 26.963 42.56 26.965 ;
  LAYER M2 ;
        RECT 40.16 27.047 42.56 27.049 ;
  LAYER M2 ;
        RECT 40.16 27.131 42.56 27.133 ;
  LAYER M2 ;
        RECT 40.16 27.215 42.56 27.217 ;
  LAYER M2 ;
        RECT 40.16 27.299 42.56 27.301 ;
  LAYER M2 ;
        RECT 40.16 27.383 42.56 27.385 ;
  LAYER M2 ;
        RECT 40.16 27.467 42.56 27.469 ;
  LAYER M2 ;
        RECT 40.16 27.551 42.56 27.553 ;
  LAYER M2 ;
        RECT 40.16 27.635 42.56 27.637 ;
  LAYER M2 ;
        RECT 40.16 27.719 42.56 27.721 ;
  LAYER M2 ;
        RECT 40.16 27.8025 42.56 27.8045 ;
  LAYER M2 ;
        RECT 40.16 27.887 42.56 27.889 ;
  LAYER M2 ;
        RECT 40.16 27.971 42.56 27.973 ;
  LAYER M2 ;
        RECT 40.16 28.055 42.56 28.057 ;
  LAYER M2 ;
        RECT 40.16 28.139 42.56 28.141 ;
  LAYER M2 ;
        RECT 40.16 28.223 42.56 28.225 ;
  LAYER M2 ;
        RECT 40.16 28.307 42.56 28.309 ;
  LAYER M2 ;
        RECT 40.16 28.391 42.56 28.393 ;
  LAYER M2 ;
        RECT 40.16 28.475 42.56 28.477 ;
  LAYER M2 ;
        RECT 40.16 28.559 42.56 28.561 ;
  LAYER M2 ;
        RECT 40.16 28.643 42.56 28.645 ;
  LAYER M2 ;
        RECT 40.16 28.727 42.56 28.729 ;
  LAYER M2 ;
        RECT 40.16 28.811 42.56 28.813 ;
  LAYER M2 ;
        RECT 40.16 28.895 42.56 28.897 ;
  LAYER M2 ;
        RECT 40.16 28.979 42.56 28.981 ;
  LAYER M2 ;
        RECT 40.16 29.063 42.56 29.065 ;
  LAYER M2 ;
        RECT 40.16 29.147 42.56 29.149 ;
  LAYER M1 ;
        RECT 39.664 17.94 39.696 20.448 ;
  LAYER M1 ;
        RECT 39.6 17.94 39.632 20.448 ;
  LAYER M1 ;
        RECT 39.536 17.94 39.568 20.448 ;
  LAYER M1 ;
        RECT 39.472 17.94 39.504 20.448 ;
  LAYER M1 ;
        RECT 39.408 17.94 39.44 20.448 ;
  LAYER M1 ;
        RECT 39.344 17.94 39.376 20.448 ;
  LAYER M1 ;
        RECT 39.28 17.94 39.312 20.448 ;
  LAYER M1 ;
        RECT 39.216 17.94 39.248 20.448 ;
  LAYER M1 ;
        RECT 39.152 17.94 39.184 20.448 ;
  LAYER M1 ;
        RECT 39.088 17.94 39.12 20.448 ;
  LAYER M1 ;
        RECT 39.024 17.94 39.056 20.448 ;
  LAYER M1 ;
        RECT 38.96 17.94 38.992 20.448 ;
  LAYER M1 ;
        RECT 38.896 17.94 38.928 20.448 ;
  LAYER M1 ;
        RECT 38.832 17.94 38.864 20.448 ;
  LAYER M1 ;
        RECT 38.768 17.94 38.8 20.448 ;
  LAYER M1 ;
        RECT 38.704 17.94 38.736 20.448 ;
  LAYER M1 ;
        RECT 38.64 17.94 38.672 20.448 ;
  LAYER M1 ;
        RECT 38.576 17.94 38.608 20.448 ;
  LAYER M1 ;
        RECT 38.512 17.94 38.544 20.448 ;
  LAYER M1 ;
        RECT 38.448 17.94 38.48 20.448 ;
  LAYER M1 ;
        RECT 38.384 17.94 38.416 20.448 ;
  LAYER M1 ;
        RECT 38.32 17.94 38.352 20.448 ;
  LAYER M1 ;
        RECT 38.256 17.94 38.288 20.448 ;
  LAYER M1 ;
        RECT 38.192 17.94 38.224 20.448 ;
  LAYER M1 ;
        RECT 38.128 17.94 38.16 20.448 ;
  LAYER M1 ;
        RECT 38.064 17.94 38.096 20.448 ;
  LAYER M1 ;
        RECT 38 17.94 38.032 20.448 ;
  LAYER M1 ;
        RECT 37.936 17.94 37.968 20.448 ;
  LAYER M1 ;
        RECT 37.872 17.94 37.904 20.448 ;
  LAYER M1 ;
        RECT 37.808 17.94 37.84 20.448 ;
  LAYER M1 ;
        RECT 37.744 17.94 37.776 20.448 ;
  LAYER M1 ;
        RECT 37.68 17.94 37.712 20.448 ;
  LAYER M1 ;
        RECT 37.616 17.94 37.648 20.448 ;
  LAYER M1 ;
        RECT 37.552 17.94 37.584 20.448 ;
  LAYER M1 ;
        RECT 37.488 17.94 37.52 20.448 ;
  LAYER M1 ;
        RECT 37.424 17.94 37.456 20.448 ;
  LAYER M1 ;
        RECT 37.36 17.94 37.392 20.448 ;
  LAYER M2 ;
        RECT 37.244 18.024 39.716 18.056 ;
  LAYER M2 ;
        RECT 37.244 18.088 39.716 18.12 ;
  LAYER M2 ;
        RECT 37.244 18.152 39.716 18.184 ;
  LAYER M2 ;
        RECT 37.244 18.216 39.716 18.248 ;
  LAYER M2 ;
        RECT 37.244 18.28 39.716 18.312 ;
  LAYER M2 ;
        RECT 37.244 18.344 39.716 18.376 ;
  LAYER M2 ;
        RECT 37.244 18.408 39.716 18.44 ;
  LAYER M2 ;
        RECT 37.244 18.472 39.716 18.504 ;
  LAYER M2 ;
        RECT 37.244 18.536 39.716 18.568 ;
  LAYER M2 ;
        RECT 37.244 18.6 39.716 18.632 ;
  LAYER M2 ;
        RECT 37.244 18.664 39.716 18.696 ;
  LAYER M2 ;
        RECT 37.244 18.728 39.716 18.76 ;
  LAYER M2 ;
        RECT 37.244 18.792 39.716 18.824 ;
  LAYER M2 ;
        RECT 37.244 18.856 39.716 18.888 ;
  LAYER M2 ;
        RECT 37.244 18.92 39.716 18.952 ;
  LAYER M2 ;
        RECT 37.244 18.984 39.716 19.016 ;
  LAYER M2 ;
        RECT 37.244 19.048 39.716 19.08 ;
  LAYER M2 ;
        RECT 37.244 19.112 39.716 19.144 ;
  LAYER M2 ;
        RECT 37.244 19.176 39.716 19.208 ;
  LAYER M2 ;
        RECT 37.244 19.24 39.716 19.272 ;
  LAYER M2 ;
        RECT 37.244 19.304 39.716 19.336 ;
  LAYER M2 ;
        RECT 37.244 19.368 39.716 19.4 ;
  LAYER M2 ;
        RECT 37.244 19.432 39.716 19.464 ;
  LAYER M2 ;
        RECT 37.244 19.496 39.716 19.528 ;
  LAYER M2 ;
        RECT 37.244 19.56 39.716 19.592 ;
  LAYER M2 ;
        RECT 37.244 19.624 39.716 19.656 ;
  LAYER M2 ;
        RECT 37.244 19.688 39.716 19.72 ;
  LAYER M2 ;
        RECT 37.244 19.752 39.716 19.784 ;
  LAYER M2 ;
        RECT 37.244 19.816 39.716 19.848 ;
  LAYER M2 ;
        RECT 37.244 19.88 39.716 19.912 ;
  LAYER M2 ;
        RECT 37.244 19.944 39.716 19.976 ;
  LAYER M2 ;
        RECT 37.244 20.008 39.716 20.04 ;
  LAYER M2 ;
        RECT 37.244 20.072 39.716 20.104 ;
  LAYER M2 ;
        RECT 37.244 20.136 39.716 20.168 ;
  LAYER M2 ;
        RECT 37.244 20.2 39.716 20.232 ;
  LAYER M2 ;
        RECT 37.244 20.264 39.716 20.296 ;
  LAYER M3 ;
        RECT 39.664 17.94 39.696 20.448 ;
  LAYER M3 ;
        RECT 39.6 17.94 39.632 20.448 ;
  LAYER M3 ;
        RECT 39.536 17.94 39.568 20.448 ;
  LAYER M3 ;
        RECT 39.472 17.94 39.504 20.448 ;
  LAYER M3 ;
        RECT 39.408 17.94 39.44 20.448 ;
  LAYER M3 ;
        RECT 39.344 17.94 39.376 20.448 ;
  LAYER M3 ;
        RECT 39.28 17.94 39.312 20.448 ;
  LAYER M3 ;
        RECT 39.216 17.94 39.248 20.448 ;
  LAYER M3 ;
        RECT 39.152 17.94 39.184 20.448 ;
  LAYER M3 ;
        RECT 39.088 17.94 39.12 20.448 ;
  LAYER M3 ;
        RECT 39.024 17.94 39.056 20.448 ;
  LAYER M3 ;
        RECT 38.96 17.94 38.992 20.448 ;
  LAYER M3 ;
        RECT 38.896 17.94 38.928 20.448 ;
  LAYER M3 ;
        RECT 38.832 17.94 38.864 20.448 ;
  LAYER M3 ;
        RECT 38.768 17.94 38.8 20.448 ;
  LAYER M3 ;
        RECT 38.704 17.94 38.736 20.448 ;
  LAYER M3 ;
        RECT 38.64 17.94 38.672 20.448 ;
  LAYER M3 ;
        RECT 38.576 17.94 38.608 20.448 ;
  LAYER M3 ;
        RECT 38.512 17.94 38.544 20.448 ;
  LAYER M3 ;
        RECT 38.448 17.94 38.48 20.448 ;
  LAYER M3 ;
        RECT 38.384 17.94 38.416 20.448 ;
  LAYER M3 ;
        RECT 38.32 17.94 38.352 20.448 ;
  LAYER M3 ;
        RECT 38.256 17.94 38.288 20.448 ;
  LAYER M3 ;
        RECT 38.192 17.94 38.224 20.448 ;
  LAYER M3 ;
        RECT 38.128 17.94 38.16 20.448 ;
  LAYER M3 ;
        RECT 38.064 17.94 38.096 20.448 ;
  LAYER M3 ;
        RECT 38 17.94 38.032 20.448 ;
  LAYER M3 ;
        RECT 37.936 17.94 37.968 20.448 ;
  LAYER M3 ;
        RECT 37.872 17.94 37.904 20.448 ;
  LAYER M3 ;
        RECT 37.808 17.94 37.84 20.448 ;
  LAYER M3 ;
        RECT 37.744 17.94 37.776 20.448 ;
  LAYER M3 ;
        RECT 37.68 17.94 37.712 20.448 ;
  LAYER M3 ;
        RECT 37.616 17.94 37.648 20.448 ;
  LAYER M3 ;
        RECT 37.552 17.94 37.584 20.448 ;
  LAYER M3 ;
        RECT 37.488 17.94 37.52 20.448 ;
  LAYER M3 ;
        RECT 37.424 17.94 37.456 20.448 ;
  LAYER M3 ;
        RECT 37.36 17.94 37.392 20.448 ;
  LAYER M3 ;
        RECT 37.264 17.94 37.296 20.448 ;
  LAYER M1 ;
        RECT 39.679 17.976 39.681 20.412 ;
  LAYER M1 ;
        RECT 39.599 17.976 39.601 20.412 ;
  LAYER M1 ;
        RECT 39.519 17.976 39.521 20.412 ;
  LAYER M1 ;
        RECT 39.439 17.976 39.441 20.412 ;
  LAYER M1 ;
        RECT 39.359 17.976 39.361 20.412 ;
  LAYER M1 ;
        RECT 39.279 17.976 39.281 20.412 ;
  LAYER M1 ;
        RECT 39.199 17.976 39.201 20.412 ;
  LAYER M1 ;
        RECT 39.119 17.976 39.121 20.412 ;
  LAYER M1 ;
        RECT 39.039 17.976 39.041 20.412 ;
  LAYER M1 ;
        RECT 38.959 17.976 38.961 20.412 ;
  LAYER M1 ;
        RECT 38.879 17.976 38.881 20.412 ;
  LAYER M1 ;
        RECT 38.799 17.976 38.801 20.412 ;
  LAYER M1 ;
        RECT 38.719 17.976 38.721 20.412 ;
  LAYER M1 ;
        RECT 38.639 17.976 38.641 20.412 ;
  LAYER M1 ;
        RECT 38.559 17.976 38.561 20.412 ;
  LAYER M1 ;
        RECT 38.479 17.976 38.481 20.412 ;
  LAYER M1 ;
        RECT 38.399 17.976 38.401 20.412 ;
  LAYER M1 ;
        RECT 38.319 17.976 38.321 20.412 ;
  LAYER M1 ;
        RECT 38.239 17.976 38.241 20.412 ;
  LAYER M1 ;
        RECT 38.159 17.976 38.161 20.412 ;
  LAYER M1 ;
        RECT 38.079 17.976 38.081 20.412 ;
  LAYER M1 ;
        RECT 37.999 17.976 38.001 20.412 ;
  LAYER M1 ;
        RECT 37.919 17.976 37.921 20.412 ;
  LAYER M1 ;
        RECT 37.839 17.976 37.841 20.412 ;
  LAYER M1 ;
        RECT 37.759 17.976 37.761 20.412 ;
  LAYER M1 ;
        RECT 37.679 17.976 37.681 20.412 ;
  LAYER M1 ;
        RECT 37.599 17.976 37.601 20.412 ;
  LAYER M1 ;
        RECT 37.519 17.976 37.521 20.412 ;
  LAYER M1 ;
        RECT 37.439 17.976 37.441 20.412 ;
  LAYER M1 ;
        RECT 37.359 17.976 37.361 20.412 ;
  LAYER M2 ;
        RECT 37.28 17.975 39.68 17.977 ;
  LAYER M2 ;
        RECT 37.28 18.059 39.68 18.061 ;
  LAYER M2 ;
        RECT 37.28 18.143 39.68 18.145 ;
  LAYER M2 ;
        RECT 37.28 18.227 39.68 18.229 ;
  LAYER M2 ;
        RECT 37.28 18.311 39.68 18.313 ;
  LAYER M2 ;
        RECT 37.28 18.395 39.68 18.397 ;
  LAYER M2 ;
        RECT 37.28 18.479 39.68 18.481 ;
  LAYER M2 ;
        RECT 37.28 18.563 39.68 18.565 ;
  LAYER M2 ;
        RECT 37.28 18.647 39.68 18.649 ;
  LAYER M2 ;
        RECT 37.28 18.731 39.68 18.733 ;
  LAYER M2 ;
        RECT 37.28 18.815 39.68 18.817 ;
  LAYER M2 ;
        RECT 37.28 18.899 39.68 18.901 ;
  LAYER M2 ;
        RECT 37.28 18.9825 39.68 18.9845 ;
  LAYER M2 ;
        RECT 37.28 19.067 39.68 19.069 ;
  LAYER M2 ;
        RECT 37.28 19.151 39.68 19.153 ;
  LAYER M2 ;
        RECT 37.28 19.235 39.68 19.237 ;
  LAYER M2 ;
        RECT 37.28 19.319 39.68 19.321 ;
  LAYER M2 ;
        RECT 37.28 19.403 39.68 19.405 ;
  LAYER M2 ;
        RECT 37.28 19.487 39.68 19.489 ;
  LAYER M2 ;
        RECT 37.28 19.571 39.68 19.573 ;
  LAYER M2 ;
        RECT 37.28 19.655 39.68 19.657 ;
  LAYER M2 ;
        RECT 37.28 19.739 39.68 19.741 ;
  LAYER M2 ;
        RECT 37.28 19.823 39.68 19.825 ;
  LAYER M2 ;
        RECT 37.28 19.907 39.68 19.909 ;
  LAYER M2 ;
        RECT 37.28 19.991 39.68 19.993 ;
  LAYER M2 ;
        RECT 37.28 20.075 39.68 20.077 ;
  LAYER M2 ;
        RECT 37.28 20.159 39.68 20.161 ;
  LAYER M2 ;
        RECT 37.28 20.243 39.68 20.245 ;
  LAYER M2 ;
        RECT 37.28 20.327 39.68 20.329 ;
  LAYER M1 ;
        RECT 39.664 20.88 39.696 23.388 ;
  LAYER M1 ;
        RECT 39.6 20.88 39.632 23.388 ;
  LAYER M1 ;
        RECT 39.536 20.88 39.568 23.388 ;
  LAYER M1 ;
        RECT 39.472 20.88 39.504 23.388 ;
  LAYER M1 ;
        RECT 39.408 20.88 39.44 23.388 ;
  LAYER M1 ;
        RECT 39.344 20.88 39.376 23.388 ;
  LAYER M1 ;
        RECT 39.28 20.88 39.312 23.388 ;
  LAYER M1 ;
        RECT 39.216 20.88 39.248 23.388 ;
  LAYER M1 ;
        RECT 39.152 20.88 39.184 23.388 ;
  LAYER M1 ;
        RECT 39.088 20.88 39.12 23.388 ;
  LAYER M1 ;
        RECT 39.024 20.88 39.056 23.388 ;
  LAYER M1 ;
        RECT 38.96 20.88 38.992 23.388 ;
  LAYER M1 ;
        RECT 38.896 20.88 38.928 23.388 ;
  LAYER M1 ;
        RECT 38.832 20.88 38.864 23.388 ;
  LAYER M1 ;
        RECT 38.768 20.88 38.8 23.388 ;
  LAYER M1 ;
        RECT 38.704 20.88 38.736 23.388 ;
  LAYER M1 ;
        RECT 38.64 20.88 38.672 23.388 ;
  LAYER M1 ;
        RECT 38.576 20.88 38.608 23.388 ;
  LAYER M1 ;
        RECT 38.512 20.88 38.544 23.388 ;
  LAYER M1 ;
        RECT 38.448 20.88 38.48 23.388 ;
  LAYER M1 ;
        RECT 38.384 20.88 38.416 23.388 ;
  LAYER M1 ;
        RECT 38.32 20.88 38.352 23.388 ;
  LAYER M1 ;
        RECT 38.256 20.88 38.288 23.388 ;
  LAYER M1 ;
        RECT 38.192 20.88 38.224 23.388 ;
  LAYER M1 ;
        RECT 38.128 20.88 38.16 23.388 ;
  LAYER M1 ;
        RECT 38.064 20.88 38.096 23.388 ;
  LAYER M1 ;
        RECT 38 20.88 38.032 23.388 ;
  LAYER M1 ;
        RECT 37.936 20.88 37.968 23.388 ;
  LAYER M1 ;
        RECT 37.872 20.88 37.904 23.388 ;
  LAYER M1 ;
        RECT 37.808 20.88 37.84 23.388 ;
  LAYER M1 ;
        RECT 37.744 20.88 37.776 23.388 ;
  LAYER M1 ;
        RECT 37.68 20.88 37.712 23.388 ;
  LAYER M1 ;
        RECT 37.616 20.88 37.648 23.388 ;
  LAYER M1 ;
        RECT 37.552 20.88 37.584 23.388 ;
  LAYER M1 ;
        RECT 37.488 20.88 37.52 23.388 ;
  LAYER M1 ;
        RECT 37.424 20.88 37.456 23.388 ;
  LAYER M1 ;
        RECT 37.36 20.88 37.392 23.388 ;
  LAYER M2 ;
        RECT 37.244 20.964 39.716 20.996 ;
  LAYER M2 ;
        RECT 37.244 21.028 39.716 21.06 ;
  LAYER M2 ;
        RECT 37.244 21.092 39.716 21.124 ;
  LAYER M2 ;
        RECT 37.244 21.156 39.716 21.188 ;
  LAYER M2 ;
        RECT 37.244 21.22 39.716 21.252 ;
  LAYER M2 ;
        RECT 37.244 21.284 39.716 21.316 ;
  LAYER M2 ;
        RECT 37.244 21.348 39.716 21.38 ;
  LAYER M2 ;
        RECT 37.244 21.412 39.716 21.444 ;
  LAYER M2 ;
        RECT 37.244 21.476 39.716 21.508 ;
  LAYER M2 ;
        RECT 37.244 21.54 39.716 21.572 ;
  LAYER M2 ;
        RECT 37.244 21.604 39.716 21.636 ;
  LAYER M2 ;
        RECT 37.244 21.668 39.716 21.7 ;
  LAYER M2 ;
        RECT 37.244 21.732 39.716 21.764 ;
  LAYER M2 ;
        RECT 37.244 21.796 39.716 21.828 ;
  LAYER M2 ;
        RECT 37.244 21.86 39.716 21.892 ;
  LAYER M2 ;
        RECT 37.244 21.924 39.716 21.956 ;
  LAYER M2 ;
        RECT 37.244 21.988 39.716 22.02 ;
  LAYER M2 ;
        RECT 37.244 22.052 39.716 22.084 ;
  LAYER M2 ;
        RECT 37.244 22.116 39.716 22.148 ;
  LAYER M2 ;
        RECT 37.244 22.18 39.716 22.212 ;
  LAYER M2 ;
        RECT 37.244 22.244 39.716 22.276 ;
  LAYER M2 ;
        RECT 37.244 22.308 39.716 22.34 ;
  LAYER M2 ;
        RECT 37.244 22.372 39.716 22.404 ;
  LAYER M2 ;
        RECT 37.244 22.436 39.716 22.468 ;
  LAYER M2 ;
        RECT 37.244 22.5 39.716 22.532 ;
  LAYER M2 ;
        RECT 37.244 22.564 39.716 22.596 ;
  LAYER M2 ;
        RECT 37.244 22.628 39.716 22.66 ;
  LAYER M2 ;
        RECT 37.244 22.692 39.716 22.724 ;
  LAYER M2 ;
        RECT 37.244 22.756 39.716 22.788 ;
  LAYER M2 ;
        RECT 37.244 22.82 39.716 22.852 ;
  LAYER M2 ;
        RECT 37.244 22.884 39.716 22.916 ;
  LAYER M2 ;
        RECT 37.244 22.948 39.716 22.98 ;
  LAYER M2 ;
        RECT 37.244 23.012 39.716 23.044 ;
  LAYER M2 ;
        RECT 37.244 23.076 39.716 23.108 ;
  LAYER M2 ;
        RECT 37.244 23.14 39.716 23.172 ;
  LAYER M2 ;
        RECT 37.244 23.204 39.716 23.236 ;
  LAYER M3 ;
        RECT 39.664 20.88 39.696 23.388 ;
  LAYER M3 ;
        RECT 39.6 20.88 39.632 23.388 ;
  LAYER M3 ;
        RECT 39.536 20.88 39.568 23.388 ;
  LAYER M3 ;
        RECT 39.472 20.88 39.504 23.388 ;
  LAYER M3 ;
        RECT 39.408 20.88 39.44 23.388 ;
  LAYER M3 ;
        RECT 39.344 20.88 39.376 23.388 ;
  LAYER M3 ;
        RECT 39.28 20.88 39.312 23.388 ;
  LAYER M3 ;
        RECT 39.216 20.88 39.248 23.388 ;
  LAYER M3 ;
        RECT 39.152 20.88 39.184 23.388 ;
  LAYER M3 ;
        RECT 39.088 20.88 39.12 23.388 ;
  LAYER M3 ;
        RECT 39.024 20.88 39.056 23.388 ;
  LAYER M3 ;
        RECT 38.96 20.88 38.992 23.388 ;
  LAYER M3 ;
        RECT 38.896 20.88 38.928 23.388 ;
  LAYER M3 ;
        RECT 38.832 20.88 38.864 23.388 ;
  LAYER M3 ;
        RECT 38.768 20.88 38.8 23.388 ;
  LAYER M3 ;
        RECT 38.704 20.88 38.736 23.388 ;
  LAYER M3 ;
        RECT 38.64 20.88 38.672 23.388 ;
  LAYER M3 ;
        RECT 38.576 20.88 38.608 23.388 ;
  LAYER M3 ;
        RECT 38.512 20.88 38.544 23.388 ;
  LAYER M3 ;
        RECT 38.448 20.88 38.48 23.388 ;
  LAYER M3 ;
        RECT 38.384 20.88 38.416 23.388 ;
  LAYER M3 ;
        RECT 38.32 20.88 38.352 23.388 ;
  LAYER M3 ;
        RECT 38.256 20.88 38.288 23.388 ;
  LAYER M3 ;
        RECT 38.192 20.88 38.224 23.388 ;
  LAYER M3 ;
        RECT 38.128 20.88 38.16 23.388 ;
  LAYER M3 ;
        RECT 38.064 20.88 38.096 23.388 ;
  LAYER M3 ;
        RECT 38 20.88 38.032 23.388 ;
  LAYER M3 ;
        RECT 37.936 20.88 37.968 23.388 ;
  LAYER M3 ;
        RECT 37.872 20.88 37.904 23.388 ;
  LAYER M3 ;
        RECT 37.808 20.88 37.84 23.388 ;
  LAYER M3 ;
        RECT 37.744 20.88 37.776 23.388 ;
  LAYER M3 ;
        RECT 37.68 20.88 37.712 23.388 ;
  LAYER M3 ;
        RECT 37.616 20.88 37.648 23.388 ;
  LAYER M3 ;
        RECT 37.552 20.88 37.584 23.388 ;
  LAYER M3 ;
        RECT 37.488 20.88 37.52 23.388 ;
  LAYER M3 ;
        RECT 37.424 20.88 37.456 23.388 ;
  LAYER M3 ;
        RECT 37.36 20.88 37.392 23.388 ;
  LAYER M3 ;
        RECT 37.264 20.88 37.296 23.388 ;
  LAYER M1 ;
        RECT 39.679 20.916 39.681 23.352 ;
  LAYER M1 ;
        RECT 39.599 20.916 39.601 23.352 ;
  LAYER M1 ;
        RECT 39.519 20.916 39.521 23.352 ;
  LAYER M1 ;
        RECT 39.439 20.916 39.441 23.352 ;
  LAYER M1 ;
        RECT 39.359 20.916 39.361 23.352 ;
  LAYER M1 ;
        RECT 39.279 20.916 39.281 23.352 ;
  LAYER M1 ;
        RECT 39.199 20.916 39.201 23.352 ;
  LAYER M1 ;
        RECT 39.119 20.916 39.121 23.352 ;
  LAYER M1 ;
        RECT 39.039 20.916 39.041 23.352 ;
  LAYER M1 ;
        RECT 38.959 20.916 38.961 23.352 ;
  LAYER M1 ;
        RECT 38.879 20.916 38.881 23.352 ;
  LAYER M1 ;
        RECT 38.799 20.916 38.801 23.352 ;
  LAYER M1 ;
        RECT 38.719 20.916 38.721 23.352 ;
  LAYER M1 ;
        RECT 38.639 20.916 38.641 23.352 ;
  LAYER M1 ;
        RECT 38.559 20.916 38.561 23.352 ;
  LAYER M1 ;
        RECT 38.479 20.916 38.481 23.352 ;
  LAYER M1 ;
        RECT 38.399 20.916 38.401 23.352 ;
  LAYER M1 ;
        RECT 38.319 20.916 38.321 23.352 ;
  LAYER M1 ;
        RECT 38.239 20.916 38.241 23.352 ;
  LAYER M1 ;
        RECT 38.159 20.916 38.161 23.352 ;
  LAYER M1 ;
        RECT 38.079 20.916 38.081 23.352 ;
  LAYER M1 ;
        RECT 37.999 20.916 38.001 23.352 ;
  LAYER M1 ;
        RECT 37.919 20.916 37.921 23.352 ;
  LAYER M1 ;
        RECT 37.839 20.916 37.841 23.352 ;
  LAYER M1 ;
        RECT 37.759 20.916 37.761 23.352 ;
  LAYER M1 ;
        RECT 37.679 20.916 37.681 23.352 ;
  LAYER M1 ;
        RECT 37.599 20.916 37.601 23.352 ;
  LAYER M1 ;
        RECT 37.519 20.916 37.521 23.352 ;
  LAYER M1 ;
        RECT 37.439 20.916 37.441 23.352 ;
  LAYER M1 ;
        RECT 37.359 20.916 37.361 23.352 ;
  LAYER M2 ;
        RECT 37.28 20.915 39.68 20.917 ;
  LAYER M2 ;
        RECT 37.28 20.999 39.68 21.001 ;
  LAYER M2 ;
        RECT 37.28 21.083 39.68 21.085 ;
  LAYER M2 ;
        RECT 37.28 21.167 39.68 21.169 ;
  LAYER M2 ;
        RECT 37.28 21.251 39.68 21.253 ;
  LAYER M2 ;
        RECT 37.28 21.335 39.68 21.337 ;
  LAYER M2 ;
        RECT 37.28 21.419 39.68 21.421 ;
  LAYER M2 ;
        RECT 37.28 21.503 39.68 21.505 ;
  LAYER M2 ;
        RECT 37.28 21.587 39.68 21.589 ;
  LAYER M2 ;
        RECT 37.28 21.671 39.68 21.673 ;
  LAYER M2 ;
        RECT 37.28 21.755 39.68 21.757 ;
  LAYER M2 ;
        RECT 37.28 21.839 39.68 21.841 ;
  LAYER M2 ;
        RECT 37.28 21.9225 39.68 21.9245 ;
  LAYER M2 ;
        RECT 37.28 22.007 39.68 22.009 ;
  LAYER M2 ;
        RECT 37.28 22.091 39.68 22.093 ;
  LAYER M2 ;
        RECT 37.28 22.175 39.68 22.177 ;
  LAYER M2 ;
        RECT 37.28 22.259 39.68 22.261 ;
  LAYER M2 ;
        RECT 37.28 22.343 39.68 22.345 ;
  LAYER M2 ;
        RECT 37.28 22.427 39.68 22.429 ;
  LAYER M2 ;
        RECT 37.28 22.511 39.68 22.513 ;
  LAYER M2 ;
        RECT 37.28 22.595 39.68 22.597 ;
  LAYER M2 ;
        RECT 37.28 22.679 39.68 22.681 ;
  LAYER M2 ;
        RECT 37.28 22.763 39.68 22.765 ;
  LAYER M2 ;
        RECT 37.28 22.847 39.68 22.849 ;
  LAYER M2 ;
        RECT 37.28 22.931 39.68 22.933 ;
  LAYER M2 ;
        RECT 37.28 23.015 39.68 23.017 ;
  LAYER M2 ;
        RECT 37.28 23.099 39.68 23.101 ;
  LAYER M2 ;
        RECT 37.28 23.183 39.68 23.185 ;
  LAYER M2 ;
        RECT 37.28 23.267 39.68 23.269 ;
  LAYER M1 ;
        RECT 39.664 23.82 39.696 26.328 ;
  LAYER M1 ;
        RECT 39.6 23.82 39.632 26.328 ;
  LAYER M1 ;
        RECT 39.536 23.82 39.568 26.328 ;
  LAYER M1 ;
        RECT 39.472 23.82 39.504 26.328 ;
  LAYER M1 ;
        RECT 39.408 23.82 39.44 26.328 ;
  LAYER M1 ;
        RECT 39.344 23.82 39.376 26.328 ;
  LAYER M1 ;
        RECT 39.28 23.82 39.312 26.328 ;
  LAYER M1 ;
        RECT 39.216 23.82 39.248 26.328 ;
  LAYER M1 ;
        RECT 39.152 23.82 39.184 26.328 ;
  LAYER M1 ;
        RECT 39.088 23.82 39.12 26.328 ;
  LAYER M1 ;
        RECT 39.024 23.82 39.056 26.328 ;
  LAYER M1 ;
        RECT 38.96 23.82 38.992 26.328 ;
  LAYER M1 ;
        RECT 38.896 23.82 38.928 26.328 ;
  LAYER M1 ;
        RECT 38.832 23.82 38.864 26.328 ;
  LAYER M1 ;
        RECT 38.768 23.82 38.8 26.328 ;
  LAYER M1 ;
        RECT 38.704 23.82 38.736 26.328 ;
  LAYER M1 ;
        RECT 38.64 23.82 38.672 26.328 ;
  LAYER M1 ;
        RECT 38.576 23.82 38.608 26.328 ;
  LAYER M1 ;
        RECT 38.512 23.82 38.544 26.328 ;
  LAYER M1 ;
        RECT 38.448 23.82 38.48 26.328 ;
  LAYER M1 ;
        RECT 38.384 23.82 38.416 26.328 ;
  LAYER M1 ;
        RECT 38.32 23.82 38.352 26.328 ;
  LAYER M1 ;
        RECT 38.256 23.82 38.288 26.328 ;
  LAYER M1 ;
        RECT 38.192 23.82 38.224 26.328 ;
  LAYER M1 ;
        RECT 38.128 23.82 38.16 26.328 ;
  LAYER M1 ;
        RECT 38.064 23.82 38.096 26.328 ;
  LAYER M1 ;
        RECT 38 23.82 38.032 26.328 ;
  LAYER M1 ;
        RECT 37.936 23.82 37.968 26.328 ;
  LAYER M1 ;
        RECT 37.872 23.82 37.904 26.328 ;
  LAYER M1 ;
        RECT 37.808 23.82 37.84 26.328 ;
  LAYER M1 ;
        RECT 37.744 23.82 37.776 26.328 ;
  LAYER M1 ;
        RECT 37.68 23.82 37.712 26.328 ;
  LAYER M1 ;
        RECT 37.616 23.82 37.648 26.328 ;
  LAYER M1 ;
        RECT 37.552 23.82 37.584 26.328 ;
  LAYER M1 ;
        RECT 37.488 23.82 37.52 26.328 ;
  LAYER M1 ;
        RECT 37.424 23.82 37.456 26.328 ;
  LAYER M1 ;
        RECT 37.36 23.82 37.392 26.328 ;
  LAYER M2 ;
        RECT 37.244 23.904 39.716 23.936 ;
  LAYER M2 ;
        RECT 37.244 23.968 39.716 24 ;
  LAYER M2 ;
        RECT 37.244 24.032 39.716 24.064 ;
  LAYER M2 ;
        RECT 37.244 24.096 39.716 24.128 ;
  LAYER M2 ;
        RECT 37.244 24.16 39.716 24.192 ;
  LAYER M2 ;
        RECT 37.244 24.224 39.716 24.256 ;
  LAYER M2 ;
        RECT 37.244 24.288 39.716 24.32 ;
  LAYER M2 ;
        RECT 37.244 24.352 39.716 24.384 ;
  LAYER M2 ;
        RECT 37.244 24.416 39.716 24.448 ;
  LAYER M2 ;
        RECT 37.244 24.48 39.716 24.512 ;
  LAYER M2 ;
        RECT 37.244 24.544 39.716 24.576 ;
  LAYER M2 ;
        RECT 37.244 24.608 39.716 24.64 ;
  LAYER M2 ;
        RECT 37.244 24.672 39.716 24.704 ;
  LAYER M2 ;
        RECT 37.244 24.736 39.716 24.768 ;
  LAYER M2 ;
        RECT 37.244 24.8 39.716 24.832 ;
  LAYER M2 ;
        RECT 37.244 24.864 39.716 24.896 ;
  LAYER M2 ;
        RECT 37.244 24.928 39.716 24.96 ;
  LAYER M2 ;
        RECT 37.244 24.992 39.716 25.024 ;
  LAYER M2 ;
        RECT 37.244 25.056 39.716 25.088 ;
  LAYER M2 ;
        RECT 37.244 25.12 39.716 25.152 ;
  LAYER M2 ;
        RECT 37.244 25.184 39.716 25.216 ;
  LAYER M2 ;
        RECT 37.244 25.248 39.716 25.28 ;
  LAYER M2 ;
        RECT 37.244 25.312 39.716 25.344 ;
  LAYER M2 ;
        RECT 37.244 25.376 39.716 25.408 ;
  LAYER M2 ;
        RECT 37.244 25.44 39.716 25.472 ;
  LAYER M2 ;
        RECT 37.244 25.504 39.716 25.536 ;
  LAYER M2 ;
        RECT 37.244 25.568 39.716 25.6 ;
  LAYER M2 ;
        RECT 37.244 25.632 39.716 25.664 ;
  LAYER M2 ;
        RECT 37.244 25.696 39.716 25.728 ;
  LAYER M2 ;
        RECT 37.244 25.76 39.716 25.792 ;
  LAYER M2 ;
        RECT 37.244 25.824 39.716 25.856 ;
  LAYER M2 ;
        RECT 37.244 25.888 39.716 25.92 ;
  LAYER M2 ;
        RECT 37.244 25.952 39.716 25.984 ;
  LAYER M2 ;
        RECT 37.244 26.016 39.716 26.048 ;
  LAYER M2 ;
        RECT 37.244 26.08 39.716 26.112 ;
  LAYER M2 ;
        RECT 37.244 26.144 39.716 26.176 ;
  LAYER M3 ;
        RECT 39.664 23.82 39.696 26.328 ;
  LAYER M3 ;
        RECT 39.6 23.82 39.632 26.328 ;
  LAYER M3 ;
        RECT 39.536 23.82 39.568 26.328 ;
  LAYER M3 ;
        RECT 39.472 23.82 39.504 26.328 ;
  LAYER M3 ;
        RECT 39.408 23.82 39.44 26.328 ;
  LAYER M3 ;
        RECT 39.344 23.82 39.376 26.328 ;
  LAYER M3 ;
        RECT 39.28 23.82 39.312 26.328 ;
  LAYER M3 ;
        RECT 39.216 23.82 39.248 26.328 ;
  LAYER M3 ;
        RECT 39.152 23.82 39.184 26.328 ;
  LAYER M3 ;
        RECT 39.088 23.82 39.12 26.328 ;
  LAYER M3 ;
        RECT 39.024 23.82 39.056 26.328 ;
  LAYER M3 ;
        RECT 38.96 23.82 38.992 26.328 ;
  LAYER M3 ;
        RECT 38.896 23.82 38.928 26.328 ;
  LAYER M3 ;
        RECT 38.832 23.82 38.864 26.328 ;
  LAYER M3 ;
        RECT 38.768 23.82 38.8 26.328 ;
  LAYER M3 ;
        RECT 38.704 23.82 38.736 26.328 ;
  LAYER M3 ;
        RECT 38.64 23.82 38.672 26.328 ;
  LAYER M3 ;
        RECT 38.576 23.82 38.608 26.328 ;
  LAYER M3 ;
        RECT 38.512 23.82 38.544 26.328 ;
  LAYER M3 ;
        RECT 38.448 23.82 38.48 26.328 ;
  LAYER M3 ;
        RECT 38.384 23.82 38.416 26.328 ;
  LAYER M3 ;
        RECT 38.32 23.82 38.352 26.328 ;
  LAYER M3 ;
        RECT 38.256 23.82 38.288 26.328 ;
  LAYER M3 ;
        RECT 38.192 23.82 38.224 26.328 ;
  LAYER M3 ;
        RECT 38.128 23.82 38.16 26.328 ;
  LAYER M3 ;
        RECT 38.064 23.82 38.096 26.328 ;
  LAYER M3 ;
        RECT 38 23.82 38.032 26.328 ;
  LAYER M3 ;
        RECT 37.936 23.82 37.968 26.328 ;
  LAYER M3 ;
        RECT 37.872 23.82 37.904 26.328 ;
  LAYER M3 ;
        RECT 37.808 23.82 37.84 26.328 ;
  LAYER M3 ;
        RECT 37.744 23.82 37.776 26.328 ;
  LAYER M3 ;
        RECT 37.68 23.82 37.712 26.328 ;
  LAYER M3 ;
        RECT 37.616 23.82 37.648 26.328 ;
  LAYER M3 ;
        RECT 37.552 23.82 37.584 26.328 ;
  LAYER M3 ;
        RECT 37.488 23.82 37.52 26.328 ;
  LAYER M3 ;
        RECT 37.424 23.82 37.456 26.328 ;
  LAYER M3 ;
        RECT 37.36 23.82 37.392 26.328 ;
  LAYER M3 ;
        RECT 37.264 23.82 37.296 26.328 ;
  LAYER M1 ;
        RECT 39.679 23.856 39.681 26.292 ;
  LAYER M1 ;
        RECT 39.599 23.856 39.601 26.292 ;
  LAYER M1 ;
        RECT 39.519 23.856 39.521 26.292 ;
  LAYER M1 ;
        RECT 39.439 23.856 39.441 26.292 ;
  LAYER M1 ;
        RECT 39.359 23.856 39.361 26.292 ;
  LAYER M1 ;
        RECT 39.279 23.856 39.281 26.292 ;
  LAYER M1 ;
        RECT 39.199 23.856 39.201 26.292 ;
  LAYER M1 ;
        RECT 39.119 23.856 39.121 26.292 ;
  LAYER M1 ;
        RECT 39.039 23.856 39.041 26.292 ;
  LAYER M1 ;
        RECT 38.959 23.856 38.961 26.292 ;
  LAYER M1 ;
        RECT 38.879 23.856 38.881 26.292 ;
  LAYER M1 ;
        RECT 38.799 23.856 38.801 26.292 ;
  LAYER M1 ;
        RECT 38.719 23.856 38.721 26.292 ;
  LAYER M1 ;
        RECT 38.639 23.856 38.641 26.292 ;
  LAYER M1 ;
        RECT 38.559 23.856 38.561 26.292 ;
  LAYER M1 ;
        RECT 38.479 23.856 38.481 26.292 ;
  LAYER M1 ;
        RECT 38.399 23.856 38.401 26.292 ;
  LAYER M1 ;
        RECT 38.319 23.856 38.321 26.292 ;
  LAYER M1 ;
        RECT 38.239 23.856 38.241 26.292 ;
  LAYER M1 ;
        RECT 38.159 23.856 38.161 26.292 ;
  LAYER M1 ;
        RECT 38.079 23.856 38.081 26.292 ;
  LAYER M1 ;
        RECT 37.999 23.856 38.001 26.292 ;
  LAYER M1 ;
        RECT 37.919 23.856 37.921 26.292 ;
  LAYER M1 ;
        RECT 37.839 23.856 37.841 26.292 ;
  LAYER M1 ;
        RECT 37.759 23.856 37.761 26.292 ;
  LAYER M1 ;
        RECT 37.679 23.856 37.681 26.292 ;
  LAYER M1 ;
        RECT 37.599 23.856 37.601 26.292 ;
  LAYER M1 ;
        RECT 37.519 23.856 37.521 26.292 ;
  LAYER M1 ;
        RECT 37.439 23.856 37.441 26.292 ;
  LAYER M1 ;
        RECT 37.359 23.856 37.361 26.292 ;
  LAYER M2 ;
        RECT 37.28 23.855 39.68 23.857 ;
  LAYER M2 ;
        RECT 37.28 23.939 39.68 23.941 ;
  LAYER M2 ;
        RECT 37.28 24.023 39.68 24.025 ;
  LAYER M2 ;
        RECT 37.28 24.107 39.68 24.109 ;
  LAYER M2 ;
        RECT 37.28 24.191 39.68 24.193 ;
  LAYER M2 ;
        RECT 37.28 24.275 39.68 24.277 ;
  LAYER M2 ;
        RECT 37.28 24.359 39.68 24.361 ;
  LAYER M2 ;
        RECT 37.28 24.443 39.68 24.445 ;
  LAYER M2 ;
        RECT 37.28 24.527 39.68 24.529 ;
  LAYER M2 ;
        RECT 37.28 24.611 39.68 24.613 ;
  LAYER M2 ;
        RECT 37.28 24.695 39.68 24.697 ;
  LAYER M2 ;
        RECT 37.28 24.779 39.68 24.781 ;
  LAYER M2 ;
        RECT 37.28 24.8625 39.68 24.8645 ;
  LAYER M2 ;
        RECT 37.28 24.947 39.68 24.949 ;
  LAYER M2 ;
        RECT 37.28 25.031 39.68 25.033 ;
  LAYER M2 ;
        RECT 37.28 25.115 39.68 25.117 ;
  LAYER M2 ;
        RECT 37.28 25.199 39.68 25.201 ;
  LAYER M2 ;
        RECT 37.28 25.283 39.68 25.285 ;
  LAYER M2 ;
        RECT 37.28 25.367 39.68 25.369 ;
  LAYER M2 ;
        RECT 37.28 25.451 39.68 25.453 ;
  LAYER M2 ;
        RECT 37.28 25.535 39.68 25.537 ;
  LAYER M2 ;
        RECT 37.28 25.619 39.68 25.621 ;
  LAYER M2 ;
        RECT 37.28 25.703 39.68 25.705 ;
  LAYER M2 ;
        RECT 37.28 25.787 39.68 25.789 ;
  LAYER M2 ;
        RECT 37.28 25.871 39.68 25.873 ;
  LAYER M2 ;
        RECT 37.28 25.955 39.68 25.957 ;
  LAYER M2 ;
        RECT 37.28 26.039 39.68 26.041 ;
  LAYER M2 ;
        RECT 37.28 26.123 39.68 26.125 ;
  LAYER M2 ;
        RECT 37.28 26.207 39.68 26.209 ;
  LAYER M1 ;
        RECT 39.664 26.76 39.696 29.268 ;
  LAYER M1 ;
        RECT 39.6 26.76 39.632 29.268 ;
  LAYER M1 ;
        RECT 39.536 26.76 39.568 29.268 ;
  LAYER M1 ;
        RECT 39.472 26.76 39.504 29.268 ;
  LAYER M1 ;
        RECT 39.408 26.76 39.44 29.268 ;
  LAYER M1 ;
        RECT 39.344 26.76 39.376 29.268 ;
  LAYER M1 ;
        RECT 39.28 26.76 39.312 29.268 ;
  LAYER M1 ;
        RECT 39.216 26.76 39.248 29.268 ;
  LAYER M1 ;
        RECT 39.152 26.76 39.184 29.268 ;
  LAYER M1 ;
        RECT 39.088 26.76 39.12 29.268 ;
  LAYER M1 ;
        RECT 39.024 26.76 39.056 29.268 ;
  LAYER M1 ;
        RECT 38.96 26.76 38.992 29.268 ;
  LAYER M1 ;
        RECT 38.896 26.76 38.928 29.268 ;
  LAYER M1 ;
        RECT 38.832 26.76 38.864 29.268 ;
  LAYER M1 ;
        RECT 38.768 26.76 38.8 29.268 ;
  LAYER M1 ;
        RECT 38.704 26.76 38.736 29.268 ;
  LAYER M1 ;
        RECT 38.64 26.76 38.672 29.268 ;
  LAYER M1 ;
        RECT 38.576 26.76 38.608 29.268 ;
  LAYER M1 ;
        RECT 38.512 26.76 38.544 29.268 ;
  LAYER M1 ;
        RECT 38.448 26.76 38.48 29.268 ;
  LAYER M1 ;
        RECT 38.384 26.76 38.416 29.268 ;
  LAYER M1 ;
        RECT 38.32 26.76 38.352 29.268 ;
  LAYER M1 ;
        RECT 38.256 26.76 38.288 29.268 ;
  LAYER M1 ;
        RECT 38.192 26.76 38.224 29.268 ;
  LAYER M1 ;
        RECT 38.128 26.76 38.16 29.268 ;
  LAYER M1 ;
        RECT 38.064 26.76 38.096 29.268 ;
  LAYER M1 ;
        RECT 38 26.76 38.032 29.268 ;
  LAYER M1 ;
        RECT 37.936 26.76 37.968 29.268 ;
  LAYER M1 ;
        RECT 37.872 26.76 37.904 29.268 ;
  LAYER M1 ;
        RECT 37.808 26.76 37.84 29.268 ;
  LAYER M1 ;
        RECT 37.744 26.76 37.776 29.268 ;
  LAYER M1 ;
        RECT 37.68 26.76 37.712 29.268 ;
  LAYER M1 ;
        RECT 37.616 26.76 37.648 29.268 ;
  LAYER M1 ;
        RECT 37.552 26.76 37.584 29.268 ;
  LAYER M1 ;
        RECT 37.488 26.76 37.52 29.268 ;
  LAYER M1 ;
        RECT 37.424 26.76 37.456 29.268 ;
  LAYER M1 ;
        RECT 37.36 26.76 37.392 29.268 ;
  LAYER M2 ;
        RECT 37.244 26.844 39.716 26.876 ;
  LAYER M2 ;
        RECT 37.244 26.908 39.716 26.94 ;
  LAYER M2 ;
        RECT 37.244 26.972 39.716 27.004 ;
  LAYER M2 ;
        RECT 37.244 27.036 39.716 27.068 ;
  LAYER M2 ;
        RECT 37.244 27.1 39.716 27.132 ;
  LAYER M2 ;
        RECT 37.244 27.164 39.716 27.196 ;
  LAYER M2 ;
        RECT 37.244 27.228 39.716 27.26 ;
  LAYER M2 ;
        RECT 37.244 27.292 39.716 27.324 ;
  LAYER M2 ;
        RECT 37.244 27.356 39.716 27.388 ;
  LAYER M2 ;
        RECT 37.244 27.42 39.716 27.452 ;
  LAYER M2 ;
        RECT 37.244 27.484 39.716 27.516 ;
  LAYER M2 ;
        RECT 37.244 27.548 39.716 27.58 ;
  LAYER M2 ;
        RECT 37.244 27.612 39.716 27.644 ;
  LAYER M2 ;
        RECT 37.244 27.676 39.716 27.708 ;
  LAYER M2 ;
        RECT 37.244 27.74 39.716 27.772 ;
  LAYER M2 ;
        RECT 37.244 27.804 39.716 27.836 ;
  LAYER M2 ;
        RECT 37.244 27.868 39.716 27.9 ;
  LAYER M2 ;
        RECT 37.244 27.932 39.716 27.964 ;
  LAYER M2 ;
        RECT 37.244 27.996 39.716 28.028 ;
  LAYER M2 ;
        RECT 37.244 28.06 39.716 28.092 ;
  LAYER M2 ;
        RECT 37.244 28.124 39.716 28.156 ;
  LAYER M2 ;
        RECT 37.244 28.188 39.716 28.22 ;
  LAYER M2 ;
        RECT 37.244 28.252 39.716 28.284 ;
  LAYER M2 ;
        RECT 37.244 28.316 39.716 28.348 ;
  LAYER M2 ;
        RECT 37.244 28.38 39.716 28.412 ;
  LAYER M2 ;
        RECT 37.244 28.444 39.716 28.476 ;
  LAYER M2 ;
        RECT 37.244 28.508 39.716 28.54 ;
  LAYER M2 ;
        RECT 37.244 28.572 39.716 28.604 ;
  LAYER M2 ;
        RECT 37.244 28.636 39.716 28.668 ;
  LAYER M2 ;
        RECT 37.244 28.7 39.716 28.732 ;
  LAYER M2 ;
        RECT 37.244 28.764 39.716 28.796 ;
  LAYER M2 ;
        RECT 37.244 28.828 39.716 28.86 ;
  LAYER M2 ;
        RECT 37.244 28.892 39.716 28.924 ;
  LAYER M2 ;
        RECT 37.244 28.956 39.716 28.988 ;
  LAYER M2 ;
        RECT 37.244 29.02 39.716 29.052 ;
  LAYER M2 ;
        RECT 37.244 29.084 39.716 29.116 ;
  LAYER M3 ;
        RECT 39.664 26.76 39.696 29.268 ;
  LAYER M3 ;
        RECT 39.6 26.76 39.632 29.268 ;
  LAYER M3 ;
        RECT 39.536 26.76 39.568 29.268 ;
  LAYER M3 ;
        RECT 39.472 26.76 39.504 29.268 ;
  LAYER M3 ;
        RECT 39.408 26.76 39.44 29.268 ;
  LAYER M3 ;
        RECT 39.344 26.76 39.376 29.268 ;
  LAYER M3 ;
        RECT 39.28 26.76 39.312 29.268 ;
  LAYER M3 ;
        RECT 39.216 26.76 39.248 29.268 ;
  LAYER M3 ;
        RECT 39.152 26.76 39.184 29.268 ;
  LAYER M3 ;
        RECT 39.088 26.76 39.12 29.268 ;
  LAYER M3 ;
        RECT 39.024 26.76 39.056 29.268 ;
  LAYER M3 ;
        RECT 38.96 26.76 38.992 29.268 ;
  LAYER M3 ;
        RECT 38.896 26.76 38.928 29.268 ;
  LAYER M3 ;
        RECT 38.832 26.76 38.864 29.268 ;
  LAYER M3 ;
        RECT 38.768 26.76 38.8 29.268 ;
  LAYER M3 ;
        RECT 38.704 26.76 38.736 29.268 ;
  LAYER M3 ;
        RECT 38.64 26.76 38.672 29.268 ;
  LAYER M3 ;
        RECT 38.576 26.76 38.608 29.268 ;
  LAYER M3 ;
        RECT 38.512 26.76 38.544 29.268 ;
  LAYER M3 ;
        RECT 38.448 26.76 38.48 29.268 ;
  LAYER M3 ;
        RECT 38.384 26.76 38.416 29.268 ;
  LAYER M3 ;
        RECT 38.32 26.76 38.352 29.268 ;
  LAYER M3 ;
        RECT 38.256 26.76 38.288 29.268 ;
  LAYER M3 ;
        RECT 38.192 26.76 38.224 29.268 ;
  LAYER M3 ;
        RECT 38.128 26.76 38.16 29.268 ;
  LAYER M3 ;
        RECT 38.064 26.76 38.096 29.268 ;
  LAYER M3 ;
        RECT 38 26.76 38.032 29.268 ;
  LAYER M3 ;
        RECT 37.936 26.76 37.968 29.268 ;
  LAYER M3 ;
        RECT 37.872 26.76 37.904 29.268 ;
  LAYER M3 ;
        RECT 37.808 26.76 37.84 29.268 ;
  LAYER M3 ;
        RECT 37.744 26.76 37.776 29.268 ;
  LAYER M3 ;
        RECT 37.68 26.76 37.712 29.268 ;
  LAYER M3 ;
        RECT 37.616 26.76 37.648 29.268 ;
  LAYER M3 ;
        RECT 37.552 26.76 37.584 29.268 ;
  LAYER M3 ;
        RECT 37.488 26.76 37.52 29.268 ;
  LAYER M3 ;
        RECT 37.424 26.76 37.456 29.268 ;
  LAYER M3 ;
        RECT 37.36 26.76 37.392 29.268 ;
  LAYER M3 ;
        RECT 37.264 26.76 37.296 29.268 ;
  LAYER M1 ;
        RECT 39.679 26.796 39.681 29.232 ;
  LAYER M1 ;
        RECT 39.599 26.796 39.601 29.232 ;
  LAYER M1 ;
        RECT 39.519 26.796 39.521 29.232 ;
  LAYER M1 ;
        RECT 39.439 26.796 39.441 29.232 ;
  LAYER M1 ;
        RECT 39.359 26.796 39.361 29.232 ;
  LAYER M1 ;
        RECT 39.279 26.796 39.281 29.232 ;
  LAYER M1 ;
        RECT 39.199 26.796 39.201 29.232 ;
  LAYER M1 ;
        RECT 39.119 26.796 39.121 29.232 ;
  LAYER M1 ;
        RECT 39.039 26.796 39.041 29.232 ;
  LAYER M1 ;
        RECT 38.959 26.796 38.961 29.232 ;
  LAYER M1 ;
        RECT 38.879 26.796 38.881 29.232 ;
  LAYER M1 ;
        RECT 38.799 26.796 38.801 29.232 ;
  LAYER M1 ;
        RECT 38.719 26.796 38.721 29.232 ;
  LAYER M1 ;
        RECT 38.639 26.796 38.641 29.232 ;
  LAYER M1 ;
        RECT 38.559 26.796 38.561 29.232 ;
  LAYER M1 ;
        RECT 38.479 26.796 38.481 29.232 ;
  LAYER M1 ;
        RECT 38.399 26.796 38.401 29.232 ;
  LAYER M1 ;
        RECT 38.319 26.796 38.321 29.232 ;
  LAYER M1 ;
        RECT 38.239 26.796 38.241 29.232 ;
  LAYER M1 ;
        RECT 38.159 26.796 38.161 29.232 ;
  LAYER M1 ;
        RECT 38.079 26.796 38.081 29.232 ;
  LAYER M1 ;
        RECT 37.999 26.796 38.001 29.232 ;
  LAYER M1 ;
        RECT 37.919 26.796 37.921 29.232 ;
  LAYER M1 ;
        RECT 37.839 26.796 37.841 29.232 ;
  LAYER M1 ;
        RECT 37.759 26.796 37.761 29.232 ;
  LAYER M1 ;
        RECT 37.679 26.796 37.681 29.232 ;
  LAYER M1 ;
        RECT 37.599 26.796 37.601 29.232 ;
  LAYER M1 ;
        RECT 37.519 26.796 37.521 29.232 ;
  LAYER M1 ;
        RECT 37.439 26.796 37.441 29.232 ;
  LAYER M1 ;
        RECT 37.359 26.796 37.361 29.232 ;
  LAYER M2 ;
        RECT 37.28 26.795 39.68 26.797 ;
  LAYER M2 ;
        RECT 37.28 26.879 39.68 26.881 ;
  LAYER M2 ;
        RECT 37.28 26.963 39.68 26.965 ;
  LAYER M2 ;
        RECT 37.28 27.047 39.68 27.049 ;
  LAYER M2 ;
        RECT 37.28 27.131 39.68 27.133 ;
  LAYER M2 ;
        RECT 37.28 27.215 39.68 27.217 ;
  LAYER M2 ;
        RECT 37.28 27.299 39.68 27.301 ;
  LAYER M2 ;
        RECT 37.28 27.383 39.68 27.385 ;
  LAYER M2 ;
        RECT 37.28 27.467 39.68 27.469 ;
  LAYER M2 ;
        RECT 37.28 27.551 39.68 27.553 ;
  LAYER M2 ;
        RECT 37.28 27.635 39.68 27.637 ;
  LAYER M2 ;
        RECT 37.28 27.719 39.68 27.721 ;
  LAYER M2 ;
        RECT 37.28 27.8025 39.68 27.8045 ;
  LAYER M2 ;
        RECT 37.28 27.887 39.68 27.889 ;
  LAYER M2 ;
        RECT 37.28 27.971 39.68 27.973 ;
  LAYER M2 ;
        RECT 37.28 28.055 39.68 28.057 ;
  LAYER M2 ;
        RECT 37.28 28.139 39.68 28.141 ;
  LAYER M2 ;
        RECT 37.28 28.223 39.68 28.225 ;
  LAYER M2 ;
        RECT 37.28 28.307 39.68 28.309 ;
  LAYER M2 ;
        RECT 37.28 28.391 39.68 28.393 ;
  LAYER M2 ;
        RECT 37.28 28.475 39.68 28.477 ;
  LAYER M2 ;
        RECT 37.28 28.559 39.68 28.561 ;
  LAYER M2 ;
        RECT 37.28 28.643 39.68 28.645 ;
  LAYER M2 ;
        RECT 37.28 28.727 39.68 28.729 ;
  LAYER M2 ;
        RECT 37.28 28.811 39.68 28.813 ;
  LAYER M2 ;
        RECT 37.28 28.895 39.68 28.897 ;
  LAYER M2 ;
        RECT 37.28 28.979 39.68 28.981 ;
  LAYER M2 ;
        RECT 37.28 29.063 39.68 29.065 ;
  LAYER M2 ;
        RECT 37.28 29.147 39.68 29.149 ;
  LAYER M1 ;
        RECT 36.784 17.94 36.816 20.448 ;
  LAYER M1 ;
        RECT 36.72 17.94 36.752 20.448 ;
  LAYER M1 ;
        RECT 36.656 17.94 36.688 20.448 ;
  LAYER M1 ;
        RECT 36.592 17.94 36.624 20.448 ;
  LAYER M1 ;
        RECT 36.528 17.94 36.56 20.448 ;
  LAYER M1 ;
        RECT 36.464 17.94 36.496 20.448 ;
  LAYER M1 ;
        RECT 36.4 17.94 36.432 20.448 ;
  LAYER M1 ;
        RECT 36.336 17.94 36.368 20.448 ;
  LAYER M1 ;
        RECT 36.272 17.94 36.304 20.448 ;
  LAYER M1 ;
        RECT 36.208 17.94 36.24 20.448 ;
  LAYER M1 ;
        RECT 36.144 17.94 36.176 20.448 ;
  LAYER M1 ;
        RECT 36.08 17.94 36.112 20.448 ;
  LAYER M1 ;
        RECT 36.016 17.94 36.048 20.448 ;
  LAYER M1 ;
        RECT 35.952 17.94 35.984 20.448 ;
  LAYER M1 ;
        RECT 35.888 17.94 35.92 20.448 ;
  LAYER M1 ;
        RECT 35.824 17.94 35.856 20.448 ;
  LAYER M1 ;
        RECT 35.76 17.94 35.792 20.448 ;
  LAYER M1 ;
        RECT 35.696 17.94 35.728 20.448 ;
  LAYER M1 ;
        RECT 35.632 17.94 35.664 20.448 ;
  LAYER M1 ;
        RECT 35.568 17.94 35.6 20.448 ;
  LAYER M1 ;
        RECT 35.504 17.94 35.536 20.448 ;
  LAYER M1 ;
        RECT 35.44 17.94 35.472 20.448 ;
  LAYER M1 ;
        RECT 35.376 17.94 35.408 20.448 ;
  LAYER M1 ;
        RECT 35.312 17.94 35.344 20.448 ;
  LAYER M1 ;
        RECT 35.248 17.94 35.28 20.448 ;
  LAYER M1 ;
        RECT 35.184 17.94 35.216 20.448 ;
  LAYER M1 ;
        RECT 35.12 17.94 35.152 20.448 ;
  LAYER M1 ;
        RECT 35.056 17.94 35.088 20.448 ;
  LAYER M1 ;
        RECT 34.992 17.94 35.024 20.448 ;
  LAYER M1 ;
        RECT 34.928 17.94 34.96 20.448 ;
  LAYER M1 ;
        RECT 34.864 17.94 34.896 20.448 ;
  LAYER M1 ;
        RECT 34.8 17.94 34.832 20.448 ;
  LAYER M1 ;
        RECT 34.736 17.94 34.768 20.448 ;
  LAYER M1 ;
        RECT 34.672 17.94 34.704 20.448 ;
  LAYER M1 ;
        RECT 34.608 17.94 34.64 20.448 ;
  LAYER M1 ;
        RECT 34.544 17.94 34.576 20.448 ;
  LAYER M1 ;
        RECT 34.48 17.94 34.512 20.448 ;
  LAYER M2 ;
        RECT 34.364 18.024 36.836 18.056 ;
  LAYER M2 ;
        RECT 34.364 18.088 36.836 18.12 ;
  LAYER M2 ;
        RECT 34.364 18.152 36.836 18.184 ;
  LAYER M2 ;
        RECT 34.364 18.216 36.836 18.248 ;
  LAYER M2 ;
        RECT 34.364 18.28 36.836 18.312 ;
  LAYER M2 ;
        RECT 34.364 18.344 36.836 18.376 ;
  LAYER M2 ;
        RECT 34.364 18.408 36.836 18.44 ;
  LAYER M2 ;
        RECT 34.364 18.472 36.836 18.504 ;
  LAYER M2 ;
        RECT 34.364 18.536 36.836 18.568 ;
  LAYER M2 ;
        RECT 34.364 18.6 36.836 18.632 ;
  LAYER M2 ;
        RECT 34.364 18.664 36.836 18.696 ;
  LAYER M2 ;
        RECT 34.364 18.728 36.836 18.76 ;
  LAYER M2 ;
        RECT 34.364 18.792 36.836 18.824 ;
  LAYER M2 ;
        RECT 34.364 18.856 36.836 18.888 ;
  LAYER M2 ;
        RECT 34.364 18.92 36.836 18.952 ;
  LAYER M2 ;
        RECT 34.364 18.984 36.836 19.016 ;
  LAYER M2 ;
        RECT 34.364 19.048 36.836 19.08 ;
  LAYER M2 ;
        RECT 34.364 19.112 36.836 19.144 ;
  LAYER M2 ;
        RECT 34.364 19.176 36.836 19.208 ;
  LAYER M2 ;
        RECT 34.364 19.24 36.836 19.272 ;
  LAYER M2 ;
        RECT 34.364 19.304 36.836 19.336 ;
  LAYER M2 ;
        RECT 34.364 19.368 36.836 19.4 ;
  LAYER M2 ;
        RECT 34.364 19.432 36.836 19.464 ;
  LAYER M2 ;
        RECT 34.364 19.496 36.836 19.528 ;
  LAYER M2 ;
        RECT 34.364 19.56 36.836 19.592 ;
  LAYER M2 ;
        RECT 34.364 19.624 36.836 19.656 ;
  LAYER M2 ;
        RECT 34.364 19.688 36.836 19.72 ;
  LAYER M2 ;
        RECT 34.364 19.752 36.836 19.784 ;
  LAYER M2 ;
        RECT 34.364 19.816 36.836 19.848 ;
  LAYER M2 ;
        RECT 34.364 19.88 36.836 19.912 ;
  LAYER M2 ;
        RECT 34.364 19.944 36.836 19.976 ;
  LAYER M2 ;
        RECT 34.364 20.008 36.836 20.04 ;
  LAYER M2 ;
        RECT 34.364 20.072 36.836 20.104 ;
  LAYER M2 ;
        RECT 34.364 20.136 36.836 20.168 ;
  LAYER M2 ;
        RECT 34.364 20.2 36.836 20.232 ;
  LAYER M2 ;
        RECT 34.364 20.264 36.836 20.296 ;
  LAYER M3 ;
        RECT 36.784 17.94 36.816 20.448 ;
  LAYER M3 ;
        RECT 36.72 17.94 36.752 20.448 ;
  LAYER M3 ;
        RECT 36.656 17.94 36.688 20.448 ;
  LAYER M3 ;
        RECT 36.592 17.94 36.624 20.448 ;
  LAYER M3 ;
        RECT 36.528 17.94 36.56 20.448 ;
  LAYER M3 ;
        RECT 36.464 17.94 36.496 20.448 ;
  LAYER M3 ;
        RECT 36.4 17.94 36.432 20.448 ;
  LAYER M3 ;
        RECT 36.336 17.94 36.368 20.448 ;
  LAYER M3 ;
        RECT 36.272 17.94 36.304 20.448 ;
  LAYER M3 ;
        RECT 36.208 17.94 36.24 20.448 ;
  LAYER M3 ;
        RECT 36.144 17.94 36.176 20.448 ;
  LAYER M3 ;
        RECT 36.08 17.94 36.112 20.448 ;
  LAYER M3 ;
        RECT 36.016 17.94 36.048 20.448 ;
  LAYER M3 ;
        RECT 35.952 17.94 35.984 20.448 ;
  LAYER M3 ;
        RECT 35.888 17.94 35.92 20.448 ;
  LAYER M3 ;
        RECT 35.824 17.94 35.856 20.448 ;
  LAYER M3 ;
        RECT 35.76 17.94 35.792 20.448 ;
  LAYER M3 ;
        RECT 35.696 17.94 35.728 20.448 ;
  LAYER M3 ;
        RECT 35.632 17.94 35.664 20.448 ;
  LAYER M3 ;
        RECT 35.568 17.94 35.6 20.448 ;
  LAYER M3 ;
        RECT 35.504 17.94 35.536 20.448 ;
  LAYER M3 ;
        RECT 35.44 17.94 35.472 20.448 ;
  LAYER M3 ;
        RECT 35.376 17.94 35.408 20.448 ;
  LAYER M3 ;
        RECT 35.312 17.94 35.344 20.448 ;
  LAYER M3 ;
        RECT 35.248 17.94 35.28 20.448 ;
  LAYER M3 ;
        RECT 35.184 17.94 35.216 20.448 ;
  LAYER M3 ;
        RECT 35.12 17.94 35.152 20.448 ;
  LAYER M3 ;
        RECT 35.056 17.94 35.088 20.448 ;
  LAYER M3 ;
        RECT 34.992 17.94 35.024 20.448 ;
  LAYER M3 ;
        RECT 34.928 17.94 34.96 20.448 ;
  LAYER M3 ;
        RECT 34.864 17.94 34.896 20.448 ;
  LAYER M3 ;
        RECT 34.8 17.94 34.832 20.448 ;
  LAYER M3 ;
        RECT 34.736 17.94 34.768 20.448 ;
  LAYER M3 ;
        RECT 34.672 17.94 34.704 20.448 ;
  LAYER M3 ;
        RECT 34.608 17.94 34.64 20.448 ;
  LAYER M3 ;
        RECT 34.544 17.94 34.576 20.448 ;
  LAYER M3 ;
        RECT 34.48 17.94 34.512 20.448 ;
  LAYER M3 ;
        RECT 34.384 17.94 34.416 20.448 ;
  LAYER M1 ;
        RECT 36.799 17.976 36.801 20.412 ;
  LAYER M1 ;
        RECT 36.719 17.976 36.721 20.412 ;
  LAYER M1 ;
        RECT 36.639 17.976 36.641 20.412 ;
  LAYER M1 ;
        RECT 36.559 17.976 36.561 20.412 ;
  LAYER M1 ;
        RECT 36.479 17.976 36.481 20.412 ;
  LAYER M1 ;
        RECT 36.399 17.976 36.401 20.412 ;
  LAYER M1 ;
        RECT 36.319 17.976 36.321 20.412 ;
  LAYER M1 ;
        RECT 36.239 17.976 36.241 20.412 ;
  LAYER M1 ;
        RECT 36.159 17.976 36.161 20.412 ;
  LAYER M1 ;
        RECT 36.079 17.976 36.081 20.412 ;
  LAYER M1 ;
        RECT 35.999 17.976 36.001 20.412 ;
  LAYER M1 ;
        RECT 35.919 17.976 35.921 20.412 ;
  LAYER M1 ;
        RECT 35.839 17.976 35.841 20.412 ;
  LAYER M1 ;
        RECT 35.759 17.976 35.761 20.412 ;
  LAYER M1 ;
        RECT 35.679 17.976 35.681 20.412 ;
  LAYER M1 ;
        RECT 35.599 17.976 35.601 20.412 ;
  LAYER M1 ;
        RECT 35.519 17.976 35.521 20.412 ;
  LAYER M1 ;
        RECT 35.439 17.976 35.441 20.412 ;
  LAYER M1 ;
        RECT 35.359 17.976 35.361 20.412 ;
  LAYER M1 ;
        RECT 35.279 17.976 35.281 20.412 ;
  LAYER M1 ;
        RECT 35.199 17.976 35.201 20.412 ;
  LAYER M1 ;
        RECT 35.119 17.976 35.121 20.412 ;
  LAYER M1 ;
        RECT 35.039 17.976 35.041 20.412 ;
  LAYER M1 ;
        RECT 34.959 17.976 34.961 20.412 ;
  LAYER M1 ;
        RECT 34.879 17.976 34.881 20.412 ;
  LAYER M1 ;
        RECT 34.799 17.976 34.801 20.412 ;
  LAYER M1 ;
        RECT 34.719 17.976 34.721 20.412 ;
  LAYER M1 ;
        RECT 34.639 17.976 34.641 20.412 ;
  LAYER M1 ;
        RECT 34.559 17.976 34.561 20.412 ;
  LAYER M1 ;
        RECT 34.479 17.976 34.481 20.412 ;
  LAYER M2 ;
        RECT 34.4 17.975 36.8 17.977 ;
  LAYER M2 ;
        RECT 34.4 18.059 36.8 18.061 ;
  LAYER M2 ;
        RECT 34.4 18.143 36.8 18.145 ;
  LAYER M2 ;
        RECT 34.4 18.227 36.8 18.229 ;
  LAYER M2 ;
        RECT 34.4 18.311 36.8 18.313 ;
  LAYER M2 ;
        RECT 34.4 18.395 36.8 18.397 ;
  LAYER M2 ;
        RECT 34.4 18.479 36.8 18.481 ;
  LAYER M2 ;
        RECT 34.4 18.563 36.8 18.565 ;
  LAYER M2 ;
        RECT 34.4 18.647 36.8 18.649 ;
  LAYER M2 ;
        RECT 34.4 18.731 36.8 18.733 ;
  LAYER M2 ;
        RECT 34.4 18.815 36.8 18.817 ;
  LAYER M2 ;
        RECT 34.4 18.899 36.8 18.901 ;
  LAYER M2 ;
        RECT 34.4 18.9825 36.8 18.9845 ;
  LAYER M2 ;
        RECT 34.4 19.067 36.8 19.069 ;
  LAYER M2 ;
        RECT 34.4 19.151 36.8 19.153 ;
  LAYER M2 ;
        RECT 34.4 19.235 36.8 19.237 ;
  LAYER M2 ;
        RECT 34.4 19.319 36.8 19.321 ;
  LAYER M2 ;
        RECT 34.4 19.403 36.8 19.405 ;
  LAYER M2 ;
        RECT 34.4 19.487 36.8 19.489 ;
  LAYER M2 ;
        RECT 34.4 19.571 36.8 19.573 ;
  LAYER M2 ;
        RECT 34.4 19.655 36.8 19.657 ;
  LAYER M2 ;
        RECT 34.4 19.739 36.8 19.741 ;
  LAYER M2 ;
        RECT 34.4 19.823 36.8 19.825 ;
  LAYER M2 ;
        RECT 34.4 19.907 36.8 19.909 ;
  LAYER M2 ;
        RECT 34.4 19.991 36.8 19.993 ;
  LAYER M2 ;
        RECT 34.4 20.075 36.8 20.077 ;
  LAYER M2 ;
        RECT 34.4 20.159 36.8 20.161 ;
  LAYER M2 ;
        RECT 34.4 20.243 36.8 20.245 ;
  LAYER M2 ;
        RECT 34.4 20.327 36.8 20.329 ;
  LAYER M1 ;
        RECT 36.784 20.88 36.816 23.388 ;
  LAYER M1 ;
        RECT 36.72 20.88 36.752 23.388 ;
  LAYER M1 ;
        RECT 36.656 20.88 36.688 23.388 ;
  LAYER M1 ;
        RECT 36.592 20.88 36.624 23.388 ;
  LAYER M1 ;
        RECT 36.528 20.88 36.56 23.388 ;
  LAYER M1 ;
        RECT 36.464 20.88 36.496 23.388 ;
  LAYER M1 ;
        RECT 36.4 20.88 36.432 23.388 ;
  LAYER M1 ;
        RECT 36.336 20.88 36.368 23.388 ;
  LAYER M1 ;
        RECT 36.272 20.88 36.304 23.388 ;
  LAYER M1 ;
        RECT 36.208 20.88 36.24 23.388 ;
  LAYER M1 ;
        RECT 36.144 20.88 36.176 23.388 ;
  LAYER M1 ;
        RECT 36.08 20.88 36.112 23.388 ;
  LAYER M1 ;
        RECT 36.016 20.88 36.048 23.388 ;
  LAYER M1 ;
        RECT 35.952 20.88 35.984 23.388 ;
  LAYER M1 ;
        RECT 35.888 20.88 35.92 23.388 ;
  LAYER M1 ;
        RECT 35.824 20.88 35.856 23.388 ;
  LAYER M1 ;
        RECT 35.76 20.88 35.792 23.388 ;
  LAYER M1 ;
        RECT 35.696 20.88 35.728 23.388 ;
  LAYER M1 ;
        RECT 35.632 20.88 35.664 23.388 ;
  LAYER M1 ;
        RECT 35.568 20.88 35.6 23.388 ;
  LAYER M1 ;
        RECT 35.504 20.88 35.536 23.388 ;
  LAYER M1 ;
        RECT 35.44 20.88 35.472 23.388 ;
  LAYER M1 ;
        RECT 35.376 20.88 35.408 23.388 ;
  LAYER M1 ;
        RECT 35.312 20.88 35.344 23.388 ;
  LAYER M1 ;
        RECT 35.248 20.88 35.28 23.388 ;
  LAYER M1 ;
        RECT 35.184 20.88 35.216 23.388 ;
  LAYER M1 ;
        RECT 35.12 20.88 35.152 23.388 ;
  LAYER M1 ;
        RECT 35.056 20.88 35.088 23.388 ;
  LAYER M1 ;
        RECT 34.992 20.88 35.024 23.388 ;
  LAYER M1 ;
        RECT 34.928 20.88 34.96 23.388 ;
  LAYER M1 ;
        RECT 34.864 20.88 34.896 23.388 ;
  LAYER M1 ;
        RECT 34.8 20.88 34.832 23.388 ;
  LAYER M1 ;
        RECT 34.736 20.88 34.768 23.388 ;
  LAYER M1 ;
        RECT 34.672 20.88 34.704 23.388 ;
  LAYER M1 ;
        RECT 34.608 20.88 34.64 23.388 ;
  LAYER M1 ;
        RECT 34.544 20.88 34.576 23.388 ;
  LAYER M1 ;
        RECT 34.48 20.88 34.512 23.388 ;
  LAYER M2 ;
        RECT 34.364 20.964 36.836 20.996 ;
  LAYER M2 ;
        RECT 34.364 21.028 36.836 21.06 ;
  LAYER M2 ;
        RECT 34.364 21.092 36.836 21.124 ;
  LAYER M2 ;
        RECT 34.364 21.156 36.836 21.188 ;
  LAYER M2 ;
        RECT 34.364 21.22 36.836 21.252 ;
  LAYER M2 ;
        RECT 34.364 21.284 36.836 21.316 ;
  LAYER M2 ;
        RECT 34.364 21.348 36.836 21.38 ;
  LAYER M2 ;
        RECT 34.364 21.412 36.836 21.444 ;
  LAYER M2 ;
        RECT 34.364 21.476 36.836 21.508 ;
  LAYER M2 ;
        RECT 34.364 21.54 36.836 21.572 ;
  LAYER M2 ;
        RECT 34.364 21.604 36.836 21.636 ;
  LAYER M2 ;
        RECT 34.364 21.668 36.836 21.7 ;
  LAYER M2 ;
        RECT 34.364 21.732 36.836 21.764 ;
  LAYER M2 ;
        RECT 34.364 21.796 36.836 21.828 ;
  LAYER M2 ;
        RECT 34.364 21.86 36.836 21.892 ;
  LAYER M2 ;
        RECT 34.364 21.924 36.836 21.956 ;
  LAYER M2 ;
        RECT 34.364 21.988 36.836 22.02 ;
  LAYER M2 ;
        RECT 34.364 22.052 36.836 22.084 ;
  LAYER M2 ;
        RECT 34.364 22.116 36.836 22.148 ;
  LAYER M2 ;
        RECT 34.364 22.18 36.836 22.212 ;
  LAYER M2 ;
        RECT 34.364 22.244 36.836 22.276 ;
  LAYER M2 ;
        RECT 34.364 22.308 36.836 22.34 ;
  LAYER M2 ;
        RECT 34.364 22.372 36.836 22.404 ;
  LAYER M2 ;
        RECT 34.364 22.436 36.836 22.468 ;
  LAYER M2 ;
        RECT 34.364 22.5 36.836 22.532 ;
  LAYER M2 ;
        RECT 34.364 22.564 36.836 22.596 ;
  LAYER M2 ;
        RECT 34.364 22.628 36.836 22.66 ;
  LAYER M2 ;
        RECT 34.364 22.692 36.836 22.724 ;
  LAYER M2 ;
        RECT 34.364 22.756 36.836 22.788 ;
  LAYER M2 ;
        RECT 34.364 22.82 36.836 22.852 ;
  LAYER M2 ;
        RECT 34.364 22.884 36.836 22.916 ;
  LAYER M2 ;
        RECT 34.364 22.948 36.836 22.98 ;
  LAYER M2 ;
        RECT 34.364 23.012 36.836 23.044 ;
  LAYER M2 ;
        RECT 34.364 23.076 36.836 23.108 ;
  LAYER M2 ;
        RECT 34.364 23.14 36.836 23.172 ;
  LAYER M2 ;
        RECT 34.364 23.204 36.836 23.236 ;
  LAYER M3 ;
        RECT 36.784 20.88 36.816 23.388 ;
  LAYER M3 ;
        RECT 36.72 20.88 36.752 23.388 ;
  LAYER M3 ;
        RECT 36.656 20.88 36.688 23.388 ;
  LAYER M3 ;
        RECT 36.592 20.88 36.624 23.388 ;
  LAYER M3 ;
        RECT 36.528 20.88 36.56 23.388 ;
  LAYER M3 ;
        RECT 36.464 20.88 36.496 23.388 ;
  LAYER M3 ;
        RECT 36.4 20.88 36.432 23.388 ;
  LAYER M3 ;
        RECT 36.336 20.88 36.368 23.388 ;
  LAYER M3 ;
        RECT 36.272 20.88 36.304 23.388 ;
  LAYER M3 ;
        RECT 36.208 20.88 36.24 23.388 ;
  LAYER M3 ;
        RECT 36.144 20.88 36.176 23.388 ;
  LAYER M3 ;
        RECT 36.08 20.88 36.112 23.388 ;
  LAYER M3 ;
        RECT 36.016 20.88 36.048 23.388 ;
  LAYER M3 ;
        RECT 35.952 20.88 35.984 23.388 ;
  LAYER M3 ;
        RECT 35.888 20.88 35.92 23.388 ;
  LAYER M3 ;
        RECT 35.824 20.88 35.856 23.388 ;
  LAYER M3 ;
        RECT 35.76 20.88 35.792 23.388 ;
  LAYER M3 ;
        RECT 35.696 20.88 35.728 23.388 ;
  LAYER M3 ;
        RECT 35.632 20.88 35.664 23.388 ;
  LAYER M3 ;
        RECT 35.568 20.88 35.6 23.388 ;
  LAYER M3 ;
        RECT 35.504 20.88 35.536 23.388 ;
  LAYER M3 ;
        RECT 35.44 20.88 35.472 23.388 ;
  LAYER M3 ;
        RECT 35.376 20.88 35.408 23.388 ;
  LAYER M3 ;
        RECT 35.312 20.88 35.344 23.388 ;
  LAYER M3 ;
        RECT 35.248 20.88 35.28 23.388 ;
  LAYER M3 ;
        RECT 35.184 20.88 35.216 23.388 ;
  LAYER M3 ;
        RECT 35.12 20.88 35.152 23.388 ;
  LAYER M3 ;
        RECT 35.056 20.88 35.088 23.388 ;
  LAYER M3 ;
        RECT 34.992 20.88 35.024 23.388 ;
  LAYER M3 ;
        RECT 34.928 20.88 34.96 23.388 ;
  LAYER M3 ;
        RECT 34.864 20.88 34.896 23.388 ;
  LAYER M3 ;
        RECT 34.8 20.88 34.832 23.388 ;
  LAYER M3 ;
        RECT 34.736 20.88 34.768 23.388 ;
  LAYER M3 ;
        RECT 34.672 20.88 34.704 23.388 ;
  LAYER M3 ;
        RECT 34.608 20.88 34.64 23.388 ;
  LAYER M3 ;
        RECT 34.544 20.88 34.576 23.388 ;
  LAYER M3 ;
        RECT 34.48 20.88 34.512 23.388 ;
  LAYER M3 ;
        RECT 34.384 20.88 34.416 23.388 ;
  LAYER M1 ;
        RECT 36.799 20.916 36.801 23.352 ;
  LAYER M1 ;
        RECT 36.719 20.916 36.721 23.352 ;
  LAYER M1 ;
        RECT 36.639 20.916 36.641 23.352 ;
  LAYER M1 ;
        RECT 36.559 20.916 36.561 23.352 ;
  LAYER M1 ;
        RECT 36.479 20.916 36.481 23.352 ;
  LAYER M1 ;
        RECT 36.399 20.916 36.401 23.352 ;
  LAYER M1 ;
        RECT 36.319 20.916 36.321 23.352 ;
  LAYER M1 ;
        RECT 36.239 20.916 36.241 23.352 ;
  LAYER M1 ;
        RECT 36.159 20.916 36.161 23.352 ;
  LAYER M1 ;
        RECT 36.079 20.916 36.081 23.352 ;
  LAYER M1 ;
        RECT 35.999 20.916 36.001 23.352 ;
  LAYER M1 ;
        RECT 35.919 20.916 35.921 23.352 ;
  LAYER M1 ;
        RECT 35.839 20.916 35.841 23.352 ;
  LAYER M1 ;
        RECT 35.759 20.916 35.761 23.352 ;
  LAYER M1 ;
        RECT 35.679 20.916 35.681 23.352 ;
  LAYER M1 ;
        RECT 35.599 20.916 35.601 23.352 ;
  LAYER M1 ;
        RECT 35.519 20.916 35.521 23.352 ;
  LAYER M1 ;
        RECT 35.439 20.916 35.441 23.352 ;
  LAYER M1 ;
        RECT 35.359 20.916 35.361 23.352 ;
  LAYER M1 ;
        RECT 35.279 20.916 35.281 23.352 ;
  LAYER M1 ;
        RECT 35.199 20.916 35.201 23.352 ;
  LAYER M1 ;
        RECT 35.119 20.916 35.121 23.352 ;
  LAYER M1 ;
        RECT 35.039 20.916 35.041 23.352 ;
  LAYER M1 ;
        RECT 34.959 20.916 34.961 23.352 ;
  LAYER M1 ;
        RECT 34.879 20.916 34.881 23.352 ;
  LAYER M1 ;
        RECT 34.799 20.916 34.801 23.352 ;
  LAYER M1 ;
        RECT 34.719 20.916 34.721 23.352 ;
  LAYER M1 ;
        RECT 34.639 20.916 34.641 23.352 ;
  LAYER M1 ;
        RECT 34.559 20.916 34.561 23.352 ;
  LAYER M1 ;
        RECT 34.479 20.916 34.481 23.352 ;
  LAYER M2 ;
        RECT 34.4 20.915 36.8 20.917 ;
  LAYER M2 ;
        RECT 34.4 20.999 36.8 21.001 ;
  LAYER M2 ;
        RECT 34.4 21.083 36.8 21.085 ;
  LAYER M2 ;
        RECT 34.4 21.167 36.8 21.169 ;
  LAYER M2 ;
        RECT 34.4 21.251 36.8 21.253 ;
  LAYER M2 ;
        RECT 34.4 21.335 36.8 21.337 ;
  LAYER M2 ;
        RECT 34.4 21.419 36.8 21.421 ;
  LAYER M2 ;
        RECT 34.4 21.503 36.8 21.505 ;
  LAYER M2 ;
        RECT 34.4 21.587 36.8 21.589 ;
  LAYER M2 ;
        RECT 34.4 21.671 36.8 21.673 ;
  LAYER M2 ;
        RECT 34.4 21.755 36.8 21.757 ;
  LAYER M2 ;
        RECT 34.4 21.839 36.8 21.841 ;
  LAYER M2 ;
        RECT 34.4 21.9225 36.8 21.9245 ;
  LAYER M2 ;
        RECT 34.4 22.007 36.8 22.009 ;
  LAYER M2 ;
        RECT 34.4 22.091 36.8 22.093 ;
  LAYER M2 ;
        RECT 34.4 22.175 36.8 22.177 ;
  LAYER M2 ;
        RECT 34.4 22.259 36.8 22.261 ;
  LAYER M2 ;
        RECT 34.4 22.343 36.8 22.345 ;
  LAYER M2 ;
        RECT 34.4 22.427 36.8 22.429 ;
  LAYER M2 ;
        RECT 34.4 22.511 36.8 22.513 ;
  LAYER M2 ;
        RECT 34.4 22.595 36.8 22.597 ;
  LAYER M2 ;
        RECT 34.4 22.679 36.8 22.681 ;
  LAYER M2 ;
        RECT 34.4 22.763 36.8 22.765 ;
  LAYER M2 ;
        RECT 34.4 22.847 36.8 22.849 ;
  LAYER M2 ;
        RECT 34.4 22.931 36.8 22.933 ;
  LAYER M2 ;
        RECT 34.4 23.015 36.8 23.017 ;
  LAYER M2 ;
        RECT 34.4 23.099 36.8 23.101 ;
  LAYER M2 ;
        RECT 34.4 23.183 36.8 23.185 ;
  LAYER M2 ;
        RECT 34.4 23.267 36.8 23.269 ;
  LAYER M1 ;
        RECT 36.784 23.82 36.816 26.328 ;
  LAYER M1 ;
        RECT 36.72 23.82 36.752 26.328 ;
  LAYER M1 ;
        RECT 36.656 23.82 36.688 26.328 ;
  LAYER M1 ;
        RECT 36.592 23.82 36.624 26.328 ;
  LAYER M1 ;
        RECT 36.528 23.82 36.56 26.328 ;
  LAYER M1 ;
        RECT 36.464 23.82 36.496 26.328 ;
  LAYER M1 ;
        RECT 36.4 23.82 36.432 26.328 ;
  LAYER M1 ;
        RECT 36.336 23.82 36.368 26.328 ;
  LAYER M1 ;
        RECT 36.272 23.82 36.304 26.328 ;
  LAYER M1 ;
        RECT 36.208 23.82 36.24 26.328 ;
  LAYER M1 ;
        RECT 36.144 23.82 36.176 26.328 ;
  LAYER M1 ;
        RECT 36.08 23.82 36.112 26.328 ;
  LAYER M1 ;
        RECT 36.016 23.82 36.048 26.328 ;
  LAYER M1 ;
        RECT 35.952 23.82 35.984 26.328 ;
  LAYER M1 ;
        RECT 35.888 23.82 35.92 26.328 ;
  LAYER M1 ;
        RECT 35.824 23.82 35.856 26.328 ;
  LAYER M1 ;
        RECT 35.76 23.82 35.792 26.328 ;
  LAYER M1 ;
        RECT 35.696 23.82 35.728 26.328 ;
  LAYER M1 ;
        RECT 35.632 23.82 35.664 26.328 ;
  LAYER M1 ;
        RECT 35.568 23.82 35.6 26.328 ;
  LAYER M1 ;
        RECT 35.504 23.82 35.536 26.328 ;
  LAYER M1 ;
        RECT 35.44 23.82 35.472 26.328 ;
  LAYER M1 ;
        RECT 35.376 23.82 35.408 26.328 ;
  LAYER M1 ;
        RECT 35.312 23.82 35.344 26.328 ;
  LAYER M1 ;
        RECT 35.248 23.82 35.28 26.328 ;
  LAYER M1 ;
        RECT 35.184 23.82 35.216 26.328 ;
  LAYER M1 ;
        RECT 35.12 23.82 35.152 26.328 ;
  LAYER M1 ;
        RECT 35.056 23.82 35.088 26.328 ;
  LAYER M1 ;
        RECT 34.992 23.82 35.024 26.328 ;
  LAYER M1 ;
        RECT 34.928 23.82 34.96 26.328 ;
  LAYER M1 ;
        RECT 34.864 23.82 34.896 26.328 ;
  LAYER M1 ;
        RECT 34.8 23.82 34.832 26.328 ;
  LAYER M1 ;
        RECT 34.736 23.82 34.768 26.328 ;
  LAYER M1 ;
        RECT 34.672 23.82 34.704 26.328 ;
  LAYER M1 ;
        RECT 34.608 23.82 34.64 26.328 ;
  LAYER M1 ;
        RECT 34.544 23.82 34.576 26.328 ;
  LAYER M1 ;
        RECT 34.48 23.82 34.512 26.328 ;
  LAYER M2 ;
        RECT 34.364 23.904 36.836 23.936 ;
  LAYER M2 ;
        RECT 34.364 23.968 36.836 24 ;
  LAYER M2 ;
        RECT 34.364 24.032 36.836 24.064 ;
  LAYER M2 ;
        RECT 34.364 24.096 36.836 24.128 ;
  LAYER M2 ;
        RECT 34.364 24.16 36.836 24.192 ;
  LAYER M2 ;
        RECT 34.364 24.224 36.836 24.256 ;
  LAYER M2 ;
        RECT 34.364 24.288 36.836 24.32 ;
  LAYER M2 ;
        RECT 34.364 24.352 36.836 24.384 ;
  LAYER M2 ;
        RECT 34.364 24.416 36.836 24.448 ;
  LAYER M2 ;
        RECT 34.364 24.48 36.836 24.512 ;
  LAYER M2 ;
        RECT 34.364 24.544 36.836 24.576 ;
  LAYER M2 ;
        RECT 34.364 24.608 36.836 24.64 ;
  LAYER M2 ;
        RECT 34.364 24.672 36.836 24.704 ;
  LAYER M2 ;
        RECT 34.364 24.736 36.836 24.768 ;
  LAYER M2 ;
        RECT 34.364 24.8 36.836 24.832 ;
  LAYER M2 ;
        RECT 34.364 24.864 36.836 24.896 ;
  LAYER M2 ;
        RECT 34.364 24.928 36.836 24.96 ;
  LAYER M2 ;
        RECT 34.364 24.992 36.836 25.024 ;
  LAYER M2 ;
        RECT 34.364 25.056 36.836 25.088 ;
  LAYER M2 ;
        RECT 34.364 25.12 36.836 25.152 ;
  LAYER M2 ;
        RECT 34.364 25.184 36.836 25.216 ;
  LAYER M2 ;
        RECT 34.364 25.248 36.836 25.28 ;
  LAYER M2 ;
        RECT 34.364 25.312 36.836 25.344 ;
  LAYER M2 ;
        RECT 34.364 25.376 36.836 25.408 ;
  LAYER M2 ;
        RECT 34.364 25.44 36.836 25.472 ;
  LAYER M2 ;
        RECT 34.364 25.504 36.836 25.536 ;
  LAYER M2 ;
        RECT 34.364 25.568 36.836 25.6 ;
  LAYER M2 ;
        RECT 34.364 25.632 36.836 25.664 ;
  LAYER M2 ;
        RECT 34.364 25.696 36.836 25.728 ;
  LAYER M2 ;
        RECT 34.364 25.76 36.836 25.792 ;
  LAYER M2 ;
        RECT 34.364 25.824 36.836 25.856 ;
  LAYER M2 ;
        RECT 34.364 25.888 36.836 25.92 ;
  LAYER M2 ;
        RECT 34.364 25.952 36.836 25.984 ;
  LAYER M2 ;
        RECT 34.364 26.016 36.836 26.048 ;
  LAYER M2 ;
        RECT 34.364 26.08 36.836 26.112 ;
  LAYER M2 ;
        RECT 34.364 26.144 36.836 26.176 ;
  LAYER M3 ;
        RECT 36.784 23.82 36.816 26.328 ;
  LAYER M3 ;
        RECT 36.72 23.82 36.752 26.328 ;
  LAYER M3 ;
        RECT 36.656 23.82 36.688 26.328 ;
  LAYER M3 ;
        RECT 36.592 23.82 36.624 26.328 ;
  LAYER M3 ;
        RECT 36.528 23.82 36.56 26.328 ;
  LAYER M3 ;
        RECT 36.464 23.82 36.496 26.328 ;
  LAYER M3 ;
        RECT 36.4 23.82 36.432 26.328 ;
  LAYER M3 ;
        RECT 36.336 23.82 36.368 26.328 ;
  LAYER M3 ;
        RECT 36.272 23.82 36.304 26.328 ;
  LAYER M3 ;
        RECT 36.208 23.82 36.24 26.328 ;
  LAYER M3 ;
        RECT 36.144 23.82 36.176 26.328 ;
  LAYER M3 ;
        RECT 36.08 23.82 36.112 26.328 ;
  LAYER M3 ;
        RECT 36.016 23.82 36.048 26.328 ;
  LAYER M3 ;
        RECT 35.952 23.82 35.984 26.328 ;
  LAYER M3 ;
        RECT 35.888 23.82 35.92 26.328 ;
  LAYER M3 ;
        RECT 35.824 23.82 35.856 26.328 ;
  LAYER M3 ;
        RECT 35.76 23.82 35.792 26.328 ;
  LAYER M3 ;
        RECT 35.696 23.82 35.728 26.328 ;
  LAYER M3 ;
        RECT 35.632 23.82 35.664 26.328 ;
  LAYER M3 ;
        RECT 35.568 23.82 35.6 26.328 ;
  LAYER M3 ;
        RECT 35.504 23.82 35.536 26.328 ;
  LAYER M3 ;
        RECT 35.44 23.82 35.472 26.328 ;
  LAYER M3 ;
        RECT 35.376 23.82 35.408 26.328 ;
  LAYER M3 ;
        RECT 35.312 23.82 35.344 26.328 ;
  LAYER M3 ;
        RECT 35.248 23.82 35.28 26.328 ;
  LAYER M3 ;
        RECT 35.184 23.82 35.216 26.328 ;
  LAYER M3 ;
        RECT 35.12 23.82 35.152 26.328 ;
  LAYER M3 ;
        RECT 35.056 23.82 35.088 26.328 ;
  LAYER M3 ;
        RECT 34.992 23.82 35.024 26.328 ;
  LAYER M3 ;
        RECT 34.928 23.82 34.96 26.328 ;
  LAYER M3 ;
        RECT 34.864 23.82 34.896 26.328 ;
  LAYER M3 ;
        RECT 34.8 23.82 34.832 26.328 ;
  LAYER M3 ;
        RECT 34.736 23.82 34.768 26.328 ;
  LAYER M3 ;
        RECT 34.672 23.82 34.704 26.328 ;
  LAYER M3 ;
        RECT 34.608 23.82 34.64 26.328 ;
  LAYER M3 ;
        RECT 34.544 23.82 34.576 26.328 ;
  LAYER M3 ;
        RECT 34.48 23.82 34.512 26.328 ;
  LAYER M3 ;
        RECT 34.384 23.82 34.416 26.328 ;
  LAYER M1 ;
        RECT 36.799 23.856 36.801 26.292 ;
  LAYER M1 ;
        RECT 36.719 23.856 36.721 26.292 ;
  LAYER M1 ;
        RECT 36.639 23.856 36.641 26.292 ;
  LAYER M1 ;
        RECT 36.559 23.856 36.561 26.292 ;
  LAYER M1 ;
        RECT 36.479 23.856 36.481 26.292 ;
  LAYER M1 ;
        RECT 36.399 23.856 36.401 26.292 ;
  LAYER M1 ;
        RECT 36.319 23.856 36.321 26.292 ;
  LAYER M1 ;
        RECT 36.239 23.856 36.241 26.292 ;
  LAYER M1 ;
        RECT 36.159 23.856 36.161 26.292 ;
  LAYER M1 ;
        RECT 36.079 23.856 36.081 26.292 ;
  LAYER M1 ;
        RECT 35.999 23.856 36.001 26.292 ;
  LAYER M1 ;
        RECT 35.919 23.856 35.921 26.292 ;
  LAYER M1 ;
        RECT 35.839 23.856 35.841 26.292 ;
  LAYER M1 ;
        RECT 35.759 23.856 35.761 26.292 ;
  LAYER M1 ;
        RECT 35.679 23.856 35.681 26.292 ;
  LAYER M1 ;
        RECT 35.599 23.856 35.601 26.292 ;
  LAYER M1 ;
        RECT 35.519 23.856 35.521 26.292 ;
  LAYER M1 ;
        RECT 35.439 23.856 35.441 26.292 ;
  LAYER M1 ;
        RECT 35.359 23.856 35.361 26.292 ;
  LAYER M1 ;
        RECT 35.279 23.856 35.281 26.292 ;
  LAYER M1 ;
        RECT 35.199 23.856 35.201 26.292 ;
  LAYER M1 ;
        RECT 35.119 23.856 35.121 26.292 ;
  LAYER M1 ;
        RECT 35.039 23.856 35.041 26.292 ;
  LAYER M1 ;
        RECT 34.959 23.856 34.961 26.292 ;
  LAYER M1 ;
        RECT 34.879 23.856 34.881 26.292 ;
  LAYER M1 ;
        RECT 34.799 23.856 34.801 26.292 ;
  LAYER M1 ;
        RECT 34.719 23.856 34.721 26.292 ;
  LAYER M1 ;
        RECT 34.639 23.856 34.641 26.292 ;
  LAYER M1 ;
        RECT 34.559 23.856 34.561 26.292 ;
  LAYER M1 ;
        RECT 34.479 23.856 34.481 26.292 ;
  LAYER M2 ;
        RECT 34.4 23.855 36.8 23.857 ;
  LAYER M2 ;
        RECT 34.4 23.939 36.8 23.941 ;
  LAYER M2 ;
        RECT 34.4 24.023 36.8 24.025 ;
  LAYER M2 ;
        RECT 34.4 24.107 36.8 24.109 ;
  LAYER M2 ;
        RECT 34.4 24.191 36.8 24.193 ;
  LAYER M2 ;
        RECT 34.4 24.275 36.8 24.277 ;
  LAYER M2 ;
        RECT 34.4 24.359 36.8 24.361 ;
  LAYER M2 ;
        RECT 34.4 24.443 36.8 24.445 ;
  LAYER M2 ;
        RECT 34.4 24.527 36.8 24.529 ;
  LAYER M2 ;
        RECT 34.4 24.611 36.8 24.613 ;
  LAYER M2 ;
        RECT 34.4 24.695 36.8 24.697 ;
  LAYER M2 ;
        RECT 34.4 24.779 36.8 24.781 ;
  LAYER M2 ;
        RECT 34.4 24.8625 36.8 24.8645 ;
  LAYER M2 ;
        RECT 34.4 24.947 36.8 24.949 ;
  LAYER M2 ;
        RECT 34.4 25.031 36.8 25.033 ;
  LAYER M2 ;
        RECT 34.4 25.115 36.8 25.117 ;
  LAYER M2 ;
        RECT 34.4 25.199 36.8 25.201 ;
  LAYER M2 ;
        RECT 34.4 25.283 36.8 25.285 ;
  LAYER M2 ;
        RECT 34.4 25.367 36.8 25.369 ;
  LAYER M2 ;
        RECT 34.4 25.451 36.8 25.453 ;
  LAYER M2 ;
        RECT 34.4 25.535 36.8 25.537 ;
  LAYER M2 ;
        RECT 34.4 25.619 36.8 25.621 ;
  LAYER M2 ;
        RECT 34.4 25.703 36.8 25.705 ;
  LAYER M2 ;
        RECT 34.4 25.787 36.8 25.789 ;
  LAYER M2 ;
        RECT 34.4 25.871 36.8 25.873 ;
  LAYER M2 ;
        RECT 34.4 25.955 36.8 25.957 ;
  LAYER M2 ;
        RECT 34.4 26.039 36.8 26.041 ;
  LAYER M2 ;
        RECT 34.4 26.123 36.8 26.125 ;
  LAYER M2 ;
        RECT 34.4 26.207 36.8 26.209 ;
  LAYER M1 ;
        RECT 36.784 26.76 36.816 29.268 ;
  LAYER M1 ;
        RECT 36.72 26.76 36.752 29.268 ;
  LAYER M1 ;
        RECT 36.656 26.76 36.688 29.268 ;
  LAYER M1 ;
        RECT 36.592 26.76 36.624 29.268 ;
  LAYER M1 ;
        RECT 36.528 26.76 36.56 29.268 ;
  LAYER M1 ;
        RECT 36.464 26.76 36.496 29.268 ;
  LAYER M1 ;
        RECT 36.4 26.76 36.432 29.268 ;
  LAYER M1 ;
        RECT 36.336 26.76 36.368 29.268 ;
  LAYER M1 ;
        RECT 36.272 26.76 36.304 29.268 ;
  LAYER M1 ;
        RECT 36.208 26.76 36.24 29.268 ;
  LAYER M1 ;
        RECT 36.144 26.76 36.176 29.268 ;
  LAYER M1 ;
        RECT 36.08 26.76 36.112 29.268 ;
  LAYER M1 ;
        RECT 36.016 26.76 36.048 29.268 ;
  LAYER M1 ;
        RECT 35.952 26.76 35.984 29.268 ;
  LAYER M1 ;
        RECT 35.888 26.76 35.92 29.268 ;
  LAYER M1 ;
        RECT 35.824 26.76 35.856 29.268 ;
  LAYER M1 ;
        RECT 35.76 26.76 35.792 29.268 ;
  LAYER M1 ;
        RECT 35.696 26.76 35.728 29.268 ;
  LAYER M1 ;
        RECT 35.632 26.76 35.664 29.268 ;
  LAYER M1 ;
        RECT 35.568 26.76 35.6 29.268 ;
  LAYER M1 ;
        RECT 35.504 26.76 35.536 29.268 ;
  LAYER M1 ;
        RECT 35.44 26.76 35.472 29.268 ;
  LAYER M1 ;
        RECT 35.376 26.76 35.408 29.268 ;
  LAYER M1 ;
        RECT 35.312 26.76 35.344 29.268 ;
  LAYER M1 ;
        RECT 35.248 26.76 35.28 29.268 ;
  LAYER M1 ;
        RECT 35.184 26.76 35.216 29.268 ;
  LAYER M1 ;
        RECT 35.12 26.76 35.152 29.268 ;
  LAYER M1 ;
        RECT 35.056 26.76 35.088 29.268 ;
  LAYER M1 ;
        RECT 34.992 26.76 35.024 29.268 ;
  LAYER M1 ;
        RECT 34.928 26.76 34.96 29.268 ;
  LAYER M1 ;
        RECT 34.864 26.76 34.896 29.268 ;
  LAYER M1 ;
        RECT 34.8 26.76 34.832 29.268 ;
  LAYER M1 ;
        RECT 34.736 26.76 34.768 29.268 ;
  LAYER M1 ;
        RECT 34.672 26.76 34.704 29.268 ;
  LAYER M1 ;
        RECT 34.608 26.76 34.64 29.268 ;
  LAYER M1 ;
        RECT 34.544 26.76 34.576 29.268 ;
  LAYER M1 ;
        RECT 34.48 26.76 34.512 29.268 ;
  LAYER M2 ;
        RECT 34.364 26.844 36.836 26.876 ;
  LAYER M2 ;
        RECT 34.364 26.908 36.836 26.94 ;
  LAYER M2 ;
        RECT 34.364 26.972 36.836 27.004 ;
  LAYER M2 ;
        RECT 34.364 27.036 36.836 27.068 ;
  LAYER M2 ;
        RECT 34.364 27.1 36.836 27.132 ;
  LAYER M2 ;
        RECT 34.364 27.164 36.836 27.196 ;
  LAYER M2 ;
        RECT 34.364 27.228 36.836 27.26 ;
  LAYER M2 ;
        RECT 34.364 27.292 36.836 27.324 ;
  LAYER M2 ;
        RECT 34.364 27.356 36.836 27.388 ;
  LAYER M2 ;
        RECT 34.364 27.42 36.836 27.452 ;
  LAYER M2 ;
        RECT 34.364 27.484 36.836 27.516 ;
  LAYER M2 ;
        RECT 34.364 27.548 36.836 27.58 ;
  LAYER M2 ;
        RECT 34.364 27.612 36.836 27.644 ;
  LAYER M2 ;
        RECT 34.364 27.676 36.836 27.708 ;
  LAYER M2 ;
        RECT 34.364 27.74 36.836 27.772 ;
  LAYER M2 ;
        RECT 34.364 27.804 36.836 27.836 ;
  LAYER M2 ;
        RECT 34.364 27.868 36.836 27.9 ;
  LAYER M2 ;
        RECT 34.364 27.932 36.836 27.964 ;
  LAYER M2 ;
        RECT 34.364 27.996 36.836 28.028 ;
  LAYER M2 ;
        RECT 34.364 28.06 36.836 28.092 ;
  LAYER M2 ;
        RECT 34.364 28.124 36.836 28.156 ;
  LAYER M2 ;
        RECT 34.364 28.188 36.836 28.22 ;
  LAYER M2 ;
        RECT 34.364 28.252 36.836 28.284 ;
  LAYER M2 ;
        RECT 34.364 28.316 36.836 28.348 ;
  LAYER M2 ;
        RECT 34.364 28.38 36.836 28.412 ;
  LAYER M2 ;
        RECT 34.364 28.444 36.836 28.476 ;
  LAYER M2 ;
        RECT 34.364 28.508 36.836 28.54 ;
  LAYER M2 ;
        RECT 34.364 28.572 36.836 28.604 ;
  LAYER M2 ;
        RECT 34.364 28.636 36.836 28.668 ;
  LAYER M2 ;
        RECT 34.364 28.7 36.836 28.732 ;
  LAYER M2 ;
        RECT 34.364 28.764 36.836 28.796 ;
  LAYER M2 ;
        RECT 34.364 28.828 36.836 28.86 ;
  LAYER M2 ;
        RECT 34.364 28.892 36.836 28.924 ;
  LAYER M2 ;
        RECT 34.364 28.956 36.836 28.988 ;
  LAYER M2 ;
        RECT 34.364 29.02 36.836 29.052 ;
  LAYER M2 ;
        RECT 34.364 29.084 36.836 29.116 ;
  LAYER M3 ;
        RECT 36.784 26.76 36.816 29.268 ;
  LAYER M3 ;
        RECT 36.72 26.76 36.752 29.268 ;
  LAYER M3 ;
        RECT 36.656 26.76 36.688 29.268 ;
  LAYER M3 ;
        RECT 36.592 26.76 36.624 29.268 ;
  LAYER M3 ;
        RECT 36.528 26.76 36.56 29.268 ;
  LAYER M3 ;
        RECT 36.464 26.76 36.496 29.268 ;
  LAYER M3 ;
        RECT 36.4 26.76 36.432 29.268 ;
  LAYER M3 ;
        RECT 36.336 26.76 36.368 29.268 ;
  LAYER M3 ;
        RECT 36.272 26.76 36.304 29.268 ;
  LAYER M3 ;
        RECT 36.208 26.76 36.24 29.268 ;
  LAYER M3 ;
        RECT 36.144 26.76 36.176 29.268 ;
  LAYER M3 ;
        RECT 36.08 26.76 36.112 29.268 ;
  LAYER M3 ;
        RECT 36.016 26.76 36.048 29.268 ;
  LAYER M3 ;
        RECT 35.952 26.76 35.984 29.268 ;
  LAYER M3 ;
        RECT 35.888 26.76 35.92 29.268 ;
  LAYER M3 ;
        RECT 35.824 26.76 35.856 29.268 ;
  LAYER M3 ;
        RECT 35.76 26.76 35.792 29.268 ;
  LAYER M3 ;
        RECT 35.696 26.76 35.728 29.268 ;
  LAYER M3 ;
        RECT 35.632 26.76 35.664 29.268 ;
  LAYER M3 ;
        RECT 35.568 26.76 35.6 29.268 ;
  LAYER M3 ;
        RECT 35.504 26.76 35.536 29.268 ;
  LAYER M3 ;
        RECT 35.44 26.76 35.472 29.268 ;
  LAYER M3 ;
        RECT 35.376 26.76 35.408 29.268 ;
  LAYER M3 ;
        RECT 35.312 26.76 35.344 29.268 ;
  LAYER M3 ;
        RECT 35.248 26.76 35.28 29.268 ;
  LAYER M3 ;
        RECT 35.184 26.76 35.216 29.268 ;
  LAYER M3 ;
        RECT 35.12 26.76 35.152 29.268 ;
  LAYER M3 ;
        RECT 35.056 26.76 35.088 29.268 ;
  LAYER M3 ;
        RECT 34.992 26.76 35.024 29.268 ;
  LAYER M3 ;
        RECT 34.928 26.76 34.96 29.268 ;
  LAYER M3 ;
        RECT 34.864 26.76 34.896 29.268 ;
  LAYER M3 ;
        RECT 34.8 26.76 34.832 29.268 ;
  LAYER M3 ;
        RECT 34.736 26.76 34.768 29.268 ;
  LAYER M3 ;
        RECT 34.672 26.76 34.704 29.268 ;
  LAYER M3 ;
        RECT 34.608 26.76 34.64 29.268 ;
  LAYER M3 ;
        RECT 34.544 26.76 34.576 29.268 ;
  LAYER M3 ;
        RECT 34.48 26.76 34.512 29.268 ;
  LAYER M3 ;
        RECT 34.384 26.76 34.416 29.268 ;
  LAYER M1 ;
        RECT 36.799 26.796 36.801 29.232 ;
  LAYER M1 ;
        RECT 36.719 26.796 36.721 29.232 ;
  LAYER M1 ;
        RECT 36.639 26.796 36.641 29.232 ;
  LAYER M1 ;
        RECT 36.559 26.796 36.561 29.232 ;
  LAYER M1 ;
        RECT 36.479 26.796 36.481 29.232 ;
  LAYER M1 ;
        RECT 36.399 26.796 36.401 29.232 ;
  LAYER M1 ;
        RECT 36.319 26.796 36.321 29.232 ;
  LAYER M1 ;
        RECT 36.239 26.796 36.241 29.232 ;
  LAYER M1 ;
        RECT 36.159 26.796 36.161 29.232 ;
  LAYER M1 ;
        RECT 36.079 26.796 36.081 29.232 ;
  LAYER M1 ;
        RECT 35.999 26.796 36.001 29.232 ;
  LAYER M1 ;
        RECT 35.919 26.796 35.921 29.232 ;
  LAYER M1 ;
        RECT 35.839 26.796 35.841 29.232 ;
  LAYER M1 ;
        RECT 35.759 26.796 35.761 29.232 ;
  LAYER M1 ;
        RECT 35.679 26.796 35.681 29.232 ;
  LAYER M1 ;
        RECT 35.599 26.796 35.601 29.232 ;
  LAYER M1 ;
        RECT 35.519 26.796 35.521 29.232 ;
  LAYER M1 ;
        RECT 35.439 26.796 35.441 29.232 ;
  LAYER M1 ;
        RECT 35.359 26.796 35.361 29.232 ;
  LAYER M1 ;
        RECT 35.279 26.796 35.281 29.232 ;
  LAYER M1 ;
        RECT 35.199 26.796 35.201 29.232 ;
  LAYER M1 ;
        RECT 35.119 26.796 35.121 29.232 ;
  LAYER M1 ;
        RECT 35.039 26.796 35.041 29.232 ;
  LAYER M1 ;
        RECT 34.959 26.796 34.961 29.232 ;
  LAYER M1 ;
        RECT 34.879 26.796 34.881 29.232 ;
  LAYER M1 ;
        RECT 34.799 26.796 34.801 29.232 ;
  LAYER M1 ;
        RECT 34.719 26.796 34.721 29.232 ;
  LAYER M1 ;
        RECT 34.639 26.796 34.641 29.232 ;
  LAYER M1 ;
        RECT 34.559 26.796 34.561 29.232 ;
  LAYER M1 ;
        RECT 34.479 26.796 34.481 29.232 ;
  LAYER M2 ;
        RECT 34.4 26.795 36.8 26.797 ;
  LAYER M2 ;
        RECT 34.4 26.879 36.8 26.881 ;
  LAYER M2 ;
        RECT 34.4 26.963 36.8 26.965 ;
  LAYER M2 ;
        RECT 34.4 27.047 36.8 27.049 ;
  LAYER M2 ;
        RECT 34.4 27.131 36.8 27.133 ;
  LAYER M2 ;
        RECT 34.4 27.215 36.8 27.217 ;
  LAYER M2 ;
        RECT 34.4 27.299 36.8 27.301 ;
  LAYER M2 ;
        RECT 34.4 27.383 36.8 27.385 ;
  LAYER M2 ;
        RECT 34.4 27.467 36.8 27.469 ;
  LAYER M2 ;
        RECT 34.4 27.551 36.8 27.553 ;
  LAYER M2 ;
        RECT 34.4 27.635 36.8 27.637 ;
  LAYER M2 ;
        RECT 34.4 27.719 36.8 27.721 ;
  LAYER M2 ;
        RECT 34.4 27.8025 36.8 27.8045 ;
  LAYER M2 ;
        RECT 34.4 27.887 36.8 27.889 ;
  LAYER M2 ;
        RECT 34.4 27.971 36.8 27.973 ;
  LAYER M2 ;
        RECT 34.4 28.055 36.8 28.057 ;
  LAYER M2 ;
        RECT 34.4 28.139 36.8 28.141 ;
  LAYER M2 ;
        RECT 34.4 28.223 36.8 28.225 ;
  LAYER M2 ;
        RECT 34.4 28.307 36.8 28.309 ;
  LAYER M2 ;
        RECT 34.4 28.391 36.8 28.393 ;
  LAYER M2 ;
        RECT 34.4 28.475 36.8 28.477 ;
  LAYER M2 ;
        RECT 34.4 28.559 36.8 28.561 ;
  LAYER M2 ;
        RECT 34.4 28.643 36.8 28.645 ;
  LAYER M2 ;
        RECT 34.4 28.727 36.8 28.729 ;
  LAYER M2 ;
        RECT 34.4 28.811 36.8 28.813 ;
  LAYER M2 ;
        RECT 34.4 28.895 36.8 28.897 ;
  LAYER M2 ;
        RECT 34.4 28.979 36.8 28.981 ;
  LAYER M2 ;
        RECT 34.4 29.063 36.8 29.065 ;
  LAYER M2 ;
        RECT 34.4 29.147 36.8 29.149 ;
  LAYER M1 ;
        RECT 33.904 17.94 33.936 20.448 ;
  LAYER M1 ;
        RECT 33.84 17.94 33.872 20.448 ;
  LAYER M1 ;
        RECT 33.776 17.94 33.808 20.448 ;
  LAYER M1 ;
        RECT 33.712 17.94 33.744 20.448 ;
  LAYER M1 ;
        RECT 33.648 17.94 33.68 20.448 ;
  LAYER M1 ;
        RECT 33.584 17.94 33.616 20.448 ;
  LAYER M1 ;
        RECT 33.52 17.94 33.552 20.448 ;
  LAYER M1 ;
        RECT 33.456 17.94 33.488 20.448 ;
  LAYER M1 ;
        RECT 33.392 17.94 33.424 20.448 ;
  LAYER M1 ;
        RECT 33.328 17.94 33.36 20.448 ;
  LAYER M1 ;
        RECT 33.264 17.94 33.296 20.448 ;
  LAYER M1 ;
        RECT 33.2 17.94 33.232 20.448 ;
  LAYER M1 ;
        RECT 33.136 17.94 33.168 20.448 ;
  LAYER M1 ;
        RECT 33.072 17.94 33.104 20.448 ;
  LAYER M1 ;
        RECT 33.008 17.94 33.04 20.448 ;
  LAYER M1 ;
        RECT 32.944 17.94 32.976 20.448 ;
  LAYER M1 ;
        RECT 32.88 17.94 32.912 20.448 ;
  LAYER M1 ;
        RECT 32.816 17.94 32.848 20.448 ;
  LAYER M1 ;
        RECT 32.752 17.94 32.784 20.448 ;
  LAYER M1 ;
        RECT 32.688 17.94 32.72 20.448 ;
  LAYER M1 ;
        RECT 32.624 17.94 32.656 20.448 ;
  LAYER M1 ;
        RECT 32.56 17.94 32.592 20.448 ;
  LAYER M1 ;
        RECT 32.496 17.94 32.528 20.448 ;
  LAYER M1 ;
        RECT 32.432 17.94 32.464 20.448 ;
  LAYER M1 ;
        RECT 32.368 17.94 32.4 20.448 ;
  LAYER M1 ;
        RECT 32.304 17.94 32.336 20.448 ;
  LAYER M1 ;
        RECT 32.24 17.94 32.272 20.448 ;
  LAYER M1 ;
        RECT 32.176 17.94 32.208 20.448 ;
  LAYER M1 ;
        RECT 32.112 17.94 32.144 20.448 ;
  LAYER M1 ;
        RECT 32.048 17.94 32.08 20.448 ;
  LAYER M1 ;
        RECT 31.984 17.94 32.016 20.448 ;
  LAYER M1 ;
        RECT 31.92 17.94 31.952 20.448 ;
  LAYER M1 ;
        RECT 31.856 17.94 31.888 20.448 ;
  LAYER M1 ;
        RECT 31.792 17.94 31.824 20.448 ;
  LAYER M1 ;
        RECT 31.728 17.94 31.76 20.448 ;
  LAYER M1 ;
        RECT 31.664 17.94 31.696 20.448 ;
  LAYER M1 ;
        RECT 31.6 17.94 31.632 20.448 ;
  LAYER M2 ;
        RECT 31.484 18.024 33.956 18.056 ;
  LAYER M2 ;
        RECT 31.484 18.088 33.956 18.12 ;
  LAYER M2 ;
        RECT 31.484 18.152 33.956 18.184 ;
  LAYER M2 ;
        RECT 31.484 18.216 33.956 18.248 ;
  LAYER M2 ;
        RECT 31.484 18.28 33.956 18.312 ;
  LAYER M2 ;
        RECT 31.484 18.344 33.956 18.376 ;
  LAYER M2 ;
        RECT 31.484 18.408 33.956 18.44 ;
  LAYER M2 ;
        RECT 31.484 18.472 33.956 18.504 ;
  LAYER M2 ;
        RECT 31.484 18.536 33.956 18.568 ;
  LAYER M2 ;
        RECT 31.484 18.6 33.956 18.632 ;
  LAYER M2 ;
        RECT 31.484 18.664 33.956 18.696 ;
  LAYER M2 ;
        RECT 31.484 18.728 33.956 18.76 ;
  LAYER M2 ;
        RECT 31.484 18.792 33.956 18.824 ;
  LAYER M2 ;
        RECT 31.484 18.856 33.956 18.888 ;
  LAYER M2 ;
        RECT 31.484 18.92 33.956 18.952 ;
  LAYER M2 ;
        RECT 31.484 18.984 33.956 19.016 ;
  LAYER M2 ;
        RECT 31.484 19.048 33.956 19.08 ;
  LAYER M2 ;
        RECT 31.484 19.112 33.956 19.144 ;
  LAYER M2 ;
        RECT 31.484 19.176 33.956 19.208 ;
  LAYER M2 ;
        RECT 31.484 19.24 33.956 19.272 ;
  LAYER M2 ;
        RECT 31.484 19.304 33.956 19.336 ;
  LAYER M2 ;
        RECT 31.484 19.368 33.956 19.4 ;
  LAYER M2 ;
        RECT 31.484 19.432 33.956 19.464 ;
  LAYER M2 ;
        RECT 31.484 19.496 33.956 19.528 ;
  LAYER M2 ;
        RECT 31.484 19.56 33.956 19.592 ;
  LAYER M2 ;
        RECT 31.484 19.624 33.956 19.656 ;
  LAYER M2 ;
        RECT 31.484 19.688 33.956 19.72 ;
  LAYER M2 ;
        RECT 31.484 19.752 33.956 19.784 ;
  LAYER M2 ;
        RECT 31.484 19.816 33.956 19.848 ;
  LAYER M2 ;
        RECT 31.484 19.88 33.956 19.912 ;
  LAYER M2 ;
        RECT 31.484 19.944 33.956 19.976 ;
  LAYER M2 ;
        RECT 31.484 20.008 33.956 20.04 ;
  LAYER M2 ;
        RECT 31.484 20.072 33.956 20.104 ;
  LAYER M2 ;
        RECT 31.484 20.136 33.956 20.168 ;
  LAYER M2 ;
        RECT 31.484 20.2 33.956 20.232 ;
  LAYER M2 ;
        RECT 31.484 20.264 33.956 20.296 ;
  LAYER M3 ;
        RECT 33.904 17.94 33.936 20.448 ;
  LAYER M3 ;
        RECT 33.84 17.94 33.872 20.448 ;
  LAYER M3 ;
        RECT 33.776 17.94 33.808 20.448 ;
  LAYER M3 ;
        RECT 33.712 17.94 33.744 20.448 ;
  LAYER M3 ;
        RECT 33.648 17.94 33.68 20.448 ;
  LAYER M3 ;
        RECT 33.584 17.94 33.616 20.448 ;
  LAYER M3 ;
        RECT 33.52 17.94 33.552 20.448 ;
  LAYER M3 ;
        RECT 33.456 17.94 33.488 20.448 ;
  LAYER M3 ;
        RECT 33.392 17.94 33.424 20.448 ;
  LAYER M3 ;
        RECT 33.328 17.94 33.36 20.448 ;
  LAYER M3 ;
        RECT 33.264 17.94 33.296 20.448 ;
  LAYER M3 ;
        RECT 33.2 17.94 33.232 20.448 ;
  LAYER M3 ;
        RECT 33.136 17.94 33.168 20.448 ;
  LAYER M3 ;
        RECT 33.072 17.94 33.104 20.448 ;
  LAYER M3 ;
        RECT 33.008 17.94 33.04 20.448 ;
  LAYER M3 ;
        RECT 32.944 17.94 32.976 20.448 ;
  LAYER M3 ;
        RECT 32.88 17.94 32.912 20.448 ;
  LAYER M3 ;
        RECT 32.816 17.94 32.848 20.448 ;
  LAYER M3 ;
        RECT 32.752 17.94 32.784 20.448 ;
  LAYER M3 ;
        RECT 32.688 17.94 32.72 20.448 ;
  LAYER M3 ;
        RECT 32.624 17.94 32.656 20.448 ;
  LAYER M3 ;
        RECT 32.56 17.94 32.592 20.448 ;
  LAYER M3 ;
        RECT 32.496 17.94 32.528 20.448 ;
  LAYER M3 ;
        RECT 32.432 17.94 32.464 20.448 ;
  LAYER M3 ;
        RECT 32.368 17.94 32.4 20.448 ;
  LAYER M3 ;
        RECT 32.304 17.94 32.336 20.448 ;
  LAYER M3 ;
        RECT 32.24 17.94 32.272 20.448 ;
  LAYER M3 ;
        RECT 32.176 17.94 32.208 20.448 ;
  LAYER M3 ;
        RECT 32.112 17.94 32.144 20.448 ;
  LAYER M3 ;
        RECT 32.048 17.94 32.08 20.448 ;
  LAYER M3 ;
        RECT 31.984 17.94 32.016 20.448 ;
  LAYER M3 ;
        RECT 31.92 17.94 31.952 20.448 ;
  LAYER M3 ;
        RECT 31.856 17.94 31.888 20.448 ;
  LAYER M3 ;
        RECT 31.792 17.94 31.824 20.448 ;
  LAYER M3 ;
        RECT 31.728 17.94 31.76 20.448 ;
  LAYER M3 ;
        RECT 31.664 17.94 31.696 20.448 ;
  LAYER M3 ;
        RECT 31.6 17.94 31.632 20.448 ;
  LAYER M3 ;
        RECT 31.504 17.94 31.536 20.448 ;
  LAYER M1 ;
        RECT 33.919 17.976 33.921 20.412 ;
  LAYER M1 ;
        RECT 33.839 17.976 33.841 20.412 ;
  LAYER M1 ;
        RECT 33.759 17.976 33.761 20.412 ;
  LAYER M1 ;
        RECT 33.679 17.976 33.681 20.412 ;
  LAYER M1 ;
        RECT 33.599 17.976 33.601 20.412 ;
  LAYER M1 ;
        RECT 33.519 17.976 33.521 20.412 ;
  LAYER M1 ;
        RECT 33.439 17.976 33.441 20.412 ;
  LAYER M1 ;
        RECT 33.359 17.976 33.361 20.412 ;
  LAYER M1 ;
        RECT 33.279 17.976 33.281 20.412 ;
  LAYER M1 ;
        RECT 33.199 17.976 33.201 20.412 ;
  LAYER M1 ;
        RECT 33.119 17.976 33.121 20.412 ;
  LAYER M1 ;
        RECT 33.039 17.976 33.041 20.412 ;
  LAYER M1 ;
        RECT 32.959 17.976 32.961 20.412 ;
  LAYER M1 ;
        RECT 32.879 17.976 32.881 20.412 ;
  LAYER M1 ;
        RECT 32.799 17.976 32.801 20.412 ;
  LAYER M1 ;
        RECT 32.719 17.976 32.721 20.412 ;
  LAYER M1 ;
        RECT 32.639 17.976 32.641 20.412 ;
  LAYER M1 ;
        RECT 32.559 17.976 32.561 20.412 ;
  LAYER M1 ;
        RECT 32.479 17.976 32.481 20.412 ;
  LAYER M1 ;
        RECT 32.399 17.976 32.401 20.412 ;
  LAYER M1 ;
        RECT 32.319 17.976 32.321 20.412 ;
  LAYER M1 ;
        RECT 32.239 17.976 32.241 20.412 ;
  LAYER M1 ;
        RECT 32.159 17.976 32.161 20.412 ;
  LAYER M1 ;
        RECT 32.079 17.976 32.081 20.412 ;
  LAYER M1 ;
        RECT 31.999 17.976 32.001 20.412 ;
  LAYER M1 ;
        RECT 31.919 17.976 31.921 20.412 ;
  LAYER M1 ;
        RECT 31.839 17.976 31.841 20.412 ;
  LAYER M1 ;
        RECT 31.759 17.976 31.761 20.412 ;
  LAYER M1 ;
        RECT 31.679 17.976 31.681 20.412 ;
  LAYER M1 ;
        RECT 31.599 17.976 31.601 20.412 ;
  LAYER M2 ;
        RECT 31.52 17.975 33.92 17.977 ;
  LAYER M2 ;
        RECT 31.52 18.059 33.92 18.061 ;
  LAYER M2 ;
        RECT 31.52 18.143 33.92 18.145 ;
  LAYER M2 ;
        RECT 31.52 18.227 33.92 18.229 ;
  LAYER M2 ;
        RECT 31.52 18.311 33.92 18.313 ;
  LAYER M2 ;
        RECT 31.52 18.395 33.92 18.397 ;
  LAYER M2 ;
        RECT 31.52 18.479 33.92 18.481 ;
  LAYER M2 ;
        RECT 31.52 18.563 33.92 18.565 ;
  LAYER M2 ;
        RECT 31.52 18.647 33.92 18.649 ;
  LAYER M2 ;
        RECT 31.52 18.731 33.92 18.733 ;
  LAYER M2 ;
        RECT 31.52 18.815 33.92 18.817 ;
  LAYER M2 ;
        RECT 31.52 18.899 33.92 18.901 ;
  LAYER M2 ;
        RECT 31.52 18.9825 33.92 18.9845 ;
  LAYER M2 ;
        RECT 31.52 19.067 33.92 19.069 ;
  LAYER M2 ;
        RECT 31.52 19.151 33.92 19.153 ;
  LAYER M2 ;
        RECT 31.52 19.235 33.92 19.237 ;
  LAYER M2 ;
        RECT 31.52 19.319 33.92 19.321 ;
  LAYER M2 ;
        RECT 31.52 19.403 33.92 19.405 ;
  LAYER M2 ;
        RECT 31.52 19.487 33.92 19.489 ;
  LAYER M2 ;
        RECT 31.52 19.571 33.92 19.573 ;
  LAYER M2 ;
        RECT 31.52 19.655 33.92 19.657 ;
  LAYER M2 ;
        RECT 31.52 19.739 33.92 19.741 ;
  LAYER M2 ;
        RECT 31.52 19.823 33.92 19.825 ;
  LAYER M2 ;
        RECT 31.52 19.907 33.92 19.909 ;
  LAYER M2 ;
        RECT 31.52 19.991 33.92 19.993 ;
  LAYER M2 ;
        RECT 31.52 20.075 33.92 20.077 ;
  LAYER M2 ;
        RECT 31.52 20.159 33.92 20.161 ;
  LAYER M2 ;
        RECT 31.52 20.243 33.92 20.245 ;
  LAYER M2 ;
        RECT 31.52 20.327 33.92 20.329 ;
  LAYER M1 ;
        RECT 33.904 20.88 33.936 23.388 ;
  LAYER M1 ;
        RECT 33.84 20.88 33.872 23.388 ;
  LAYER M1 ;
        RECT 33.776 20.88 33.808 23.388 ;
  LAYER M1 ;
        RECT 33.712 20.88 33.744 23.388 ;
  LAYER M1 ;
        RECT 33.648 20.88 33.68 23.388 ;
  LAYER M1 ;
        RECT 33.584 20.88 33.616 23.388 ;
  LAYER M1 ;
        RECT 33.52 20.88 33.552 23.388 ;
  LAYER M1 ;
        RECT 33.456 20.88 33.488 23.388 ;
  LAYER M1 ;
        RECT 33.392 20.88 33.424 23.388 ;
  LAYER M1 ;
        RECT 33.328 20.88 33.36 23.388 ;
  LAYER M1 ;
        RECT 33.264 20.88 33.296 23.388 ;
  LAYER M1 ;
        RECT 33.2 20.88 33.232 23.388 ;
  LAYER M1 ;
        RECT 33.136 20.88 33.168 23.388 ;
  LAYER M1 ;
        RECT 33.072 20.88 33.104 23.388 ;
  LAYER M1 ;
        RECT 33.008 20.88 33.04 23.388 ;
  LAYER M1 ;
        RECT 32.944 20.88 32.976 23.388 ;
  LAYER M1 ;
        RECT 32.88 20.88 32.912 23.388 ;
  LAYER M1 ;
        RECT 32.816 20.88 32.848 23.388 ;
  LAYER M1 ;
        RECT 32.752 20.88 32.784 23.388 ;
  LAYER M1 ;
        RECT 32.688 20.88 32.72 23.388 ;
  LAYER M1 ;
        RECT 32.624 20.88 32.656 23.388 ;
  LAYER M1 ;
        RECT 32.56 20.88 32.592 23.388 ;
  LAYER M1 ;
        RECT 32.496 20.88 32.528 23.388 ;
  LAYER M1 ;
        RECT 32.432 20.88 32.464 23.388 ;
  LAYER M1 ;
        RECT 32.368 20.88 32.4 23.388 ;
  LAYER M1 ;
        RECT 32.304 20.88 32.336 23.388 ;
  LAYER M1 ;
        RECT 32.24 20.88 32.272 23.388 ;
  LAYER M1 ;
        RECT 32.176 20.88 32.208 23.388 ;
  LAYER M1 ;
        RECT 32.112 20.88 32.144 23.388 ;
  LAYER M1 ;
        RECT 32.048 20.88 32.08 23.388 ;
  LAYER M1 ;
        RECT 31.984 20.88 32.016 23.388 ;
  LAYER M1 ;
        RECT 31.92 20.88 31.952 23.388 ;
  LAYER M1 ;
        RECT 31.856 20.88 31.888 23.388 ;
  LAYER M1 ;
        RECT 31.792 20.88 31.824 23.388 ;
  LAYER M1 ;
        RECT 31.728 20.88 31.76 23.388 ;
  LAYER M1 ;
        RECT 31.664 20.88 31.696 23.388 ;
  LAYER M1 ;
        RECT 31.6 20.88 31.632 23.388 ;
  LAYER M2 ;
        RECT 31.484 20.964 33.956 20.996 ;
  LAYER M2 ;
        RECT 31.484 21.028 33.956 21.06 ;
  LAYER M2 ;
        RECT 31.484 21.092 33.956 21.124 ;
  LAYER M2 ;
        RECT 31.484 21.156 33.956 21.188 ;
  LAYER M2 ;
        RECT 31.484 21.22 33.956 21.252 ;
  LAYER M2 ;
        RECT 31.484 21.284 33.956 21.316 ;
  LAYER M2 ;
        RECT 31.484 21.348 33.956 21.38 ;
  LAYER M2 ;
        RECT 31.484 21.412 33.956 21.444 ;
  LAYER M2 ;
        RECT 31.484 21.476 33.956 21.508 ;
  LAYER M2 ;
        RECT 31.484 21.54 33.956 21.572 ;
  LAYER M2 ;
        RECT 31.484 21.604 33.956 21.636 ;
  LAYER M2 ;
        RECT 31.484 21.668 33.956 21.7 ;
  LAYER M2 ;
        RECT 31.484 21.732 33.956 21.764 ;
  LAYER M2 ;
        RECT 31.484 21.796 33.956 21.828 ;
  LAYER M2 ;
        RECT 31.484 21.86 33.956 21.892 ;
  LAYER M2 ;
        RECT 31.484 21.924 33.956 21.956 ;
  LAYER M2 ;
        RECT 31.484 21.988 33.956 22.02 ;
  LAYER M2 ;
        RECT 31.484 22.052 33.956 22.084 ;
  LAYER M2 ;
        RECT 31.484 22.116 33.956 22.148 ;
  LAYER M2 ;
        RECT 31.484 22.18 33.956 22.212 ;
  LAYER M2 ;
        RECT 31.484 22.244 33.956 22.276 ;
  LAYER M2 ;
        RECT 31.484 22.308 33.956 22.34 ;
  LAYER M2 ;
        RECT 31.484 22.372 33.956 22.404 ;
  LAYER M2 ;
        RECT 31.484 22.436 33.956 22.468 ;
  LAYER M2 ;
        RECT 31.484 22.5 33.956 22.532 ;
  LAYER M2 ;
        RECT 31.484 22.564 33.956 22.596 ;
  LAYER M2 ;
        RECT 31.484 22.628 33.956 22.66 ;
  LAYER M2 ;
        RECT 31.484 22.692 33.956 22.724 ;
  LAYER M2 ;
        RECT 31.484 22.756 33.956 22.788 ;
  LAYER M2 ;
        RECT 31.484 22.82 33.956 22.852 ;
  LAYER M2 ;
        RECT 31.484 22.884 33.956 22.916 ;
  LAYER M2 ;
        RECT 31.484 22.948 33.956 22.98 ;
  LAYER M2 ;
        RECT 31.484 23.012 33.956 23.044 ;
  LAYER M2 ;
        RECT 31.484 23.076 33.956 23.108 ;
  LAYER M2 ;
        RECT 31.484 23.14 33.956 23.172 ;
  LAYER M2 ;
        RECT 31.484 23.204 33.956 23.236 ;
  LAYER M3 ;
        RECT 33.904 20.88 33.936 23.388 ;
  LAYER M3 ;
        RECT 33.84 20.88 33.872 23.388 ;
  LAYER M3 ;
        RECT 33.776 20.88 33.808 23.388 ;
  LAYER M3 ;
        RECT 33.712 20.88 33.744 23.388 ;
  LAYER M3 ;
        RECT 33.648 20.88 33.68 23.388 ;
  LAYER M3 ;
        RECT 33.584 20.88 33.616 23.388 ;
  LAYER M3 ;
        RECT 33.52 20.88 33.552 23.388 ;
  LAYER M3 ;
        RECT 33.456 20.88 33.488 23.388 ;
  LAYER M3 ;
        RECT 33.392 20.88 33.424 23.388 ;
  LAYER M3 ;
        RECT 33.328 20.88 33.36 23.388 ;
  LAYER M3 ;
        RECT 33.264 20.88 33.296 23.388 ;
  LAYER M3 ;
        RECT 33.2 20.88 33.232 23.388 ;
  LAYER M3 ;
        RECT 33.136 20.88 33.168 23.388 ;
  LAYER M3 ;
        RECT 33.072 20.88 33.104 23.388 ;
  LAYER M3 ;
        RECT 33.008 20.88 33.04 23.388 ;
  LAYER M3 ;
        RECT 32.944 20.88 32.976 23.388 ;
  LAYER M3 ;
        RECT 32.88 20.88 32.912 23.388 ;
  LAYER M3 ;
        RECT 32.816 20.88 32.848 23.388 ;
  LAYER M3 ;
        RECT 32.752 20.88 32.784 23.388 ;
  LAYER M3 ;
        RECT 32.688 20.88 32.72 23.388 ;
  LAYER M3 ;
        RECT 32.624 20.88 32.656 23.388 ;
  LAYER M3 ;
        RECT 32.56 20.88 32.592 23.388 ;
  LAYER M3 ;
        RECT 32.496 20.88 32.528 23.388 ;
  LAYER M3 ;
        RECT 32.432 20.88 32.464 23.388 ;
  LAYER M3 ;
        RECT 32.368 20.88 32.4 23.388 ;
  LAYER M3 ;
        RECT 32.304 20.88 32.336 23.388 ;
  LAYER M3 ;
        RECT 32.24 20.88 32.272 23.388 ;
  LAYER M3 ;
        RECT 32.176 20.88 32.208 23.388 ;
  LAYER M3 ;
        RECT 32.112 20.88 32.144 23.388 ;
  LAYER M3 ;
        RECT 32.048 20.88 32.08 23.388 ;
  LAYER M3 ;
        RECT 31.984 20.88 32.016 23.388 ;
  LAYER M3 ;
        RECT 31.92 20.88 31.952 23.388 ;
  LAYER M3 ;
        RECT 31.856 20.88 31.888 23.388 ;
  LAYER M3 ;
        RECT 31.792 20.88 31.824 23.388 ;
  LAYER M3 ;
        RECT 31.728 20.88 31.76 23.388 ;
  LAYER M3 ;
        RECT 31.664 20.88 31.696 23.388 ;
  LAYER M3 ;
        RECT 31.6 20.88 31.632 23.388 ;
  LAYER M3 ;
        RECT 31.504 20.88 31.536 23.388 ;
  LAYER M1 ;
        RECT 33.919 20.916 33.921 23.352 ;
  LAYER M1 ;
        RECT 33.839 20.916 33.841 23.352 ;
  LAYER M1 ;
        RECT 33.759 20.916 33.761 23.352 ;
  LAYER M1 ;
        RECT 33.679 20.916 33.681 23.352 ;
  LAYER M1 ;
        RECT 33.599 20.916 33.601 23.352 ;
  LAYER M1 ;
        RECT 33.519 20.916 33.521 23.352 ;
  LAYER M1 ;
        RECT 33.439 20.916 33.441 23.352 ;
  LAYER M1 ;
        RECT 33.359 20.916 33.361 23.352 ;
  LAYER M1 ;
        RECT 33.279 20.916 33.281 23.352 ;
  LAYER M1 ;
        RECT 33.199 20.916 33.201 23.352 ;
  LAYER M1 ;
        RECT 33.119 20.916 33.121 23.352 ;
  LAYER M1 ;
        RECT 33.039 20.916 33.041 23.352 ;
  LAYER M1 ;
        RECT 32.959 20.916 32.961 23.352 ;
  LAYER M1 ;
        RECT 32.879 20.916 32.881 23.352 ;
  LAYER M1 ;
        RECT 32.799 20.916 32.801 23.352 ;
  LAYER M1 ;
        RECT 32.719 20.916 32.721 23.352 ;
  LAYER M1 ;
        RECT 32.639 20.916 32.641 23.352 ;
  LAYER M1 ;
        RECT 32.559 20.916 32.561 23.352 ;
  LAYER M1 ;
        RECT 32.479 20.916 32.481 23.352 ;
  LAYER M1 ;
        RECT 32.399 20.916 32.401 23.352 ;
  LAYER M1 ;
        RECT 32.319 20.916 32.321 23.352 ;
  LAYER M1 ;
        RECT 32.239 20.916 32.241 23.352 ;
  LAYER M1 ;
        RECT 32.159 20.916 32.161 23.352 ;
  LAYER M1 ;
        RECT 32.079 20.916 32.081 23.352 ;
  LAYER M1 ;
        RECT 31.999 20.916 32.001 23.352 ;
  LAYER M1 ;
        RECT 31.919 20.916 31.921 23.352 ;
  LAYER M1 ;
        RECT 31.839 20.916 31.841 23.352 ;
  LAYER M1 ;
        RECT 31.759 20.916 31.761 23.352 ;
  LAYER M1 ;
        RECT 31.679 20.916 31.681 23.352 ;
  LAYER M1 ;
        RECT 31.599 20.916 31.601 23.352 ;
  LAYER M2 ;
        RECT 31.52 20.915 33.92 20.917 ;
  LAYER M2 ;
        RECT 31.52 20.999 33.92 21.001 ;
  LAYER M2 ;
        RECT 31.52 21.083 33.92 21.085 ;
  LAYER M2 ;
        RECT 31.52 21.167 33.92 21.169 ;
  LAYER M2 ;
        RECT 31.52 21.251 33.92 21.253 ;
  LAYER M2 ;
        RECT 31.52 21.335 33.92 21.337 ;
  LAYER M2 ;
        RECT 31.52 21.419 33.92 21.421 ;
  LAYER M2 ;
        RECT 31.52 21.503 33.92 21.505 ;
  LAYER M2 ;
        RECT 31.52 21.587 33.92 21.589 ;
  LAYER M2 ;
        RECT 31.52 21.671 33.92 21.673 ;
  LAYER M2 ;
        RECT 31.52 21.755 33.92 21.757 ;
  LAYER M2 ;
        RECT 31.52 21.839 33.92 21.841 ;
  LAYER M2 ;
        RECT 31.52 21.9225 33.92 21.9245 ;
  LAYER M2 ;
        RECT 31.52 22.007 33.92 22.009 ;
  LAYER M2 ;
        RECT 31.52 22.091 33.92 22.093 ;
  LAYER M2 ;
        RECT 31.52 22.175 33.92 22.177 ;
  LAYER M2 ;
        RECT 31.52 22.259 33.92 22.261 ;
  LAYER M2 ;
        RECT 31.52 22.343 33.92 22.345 ;
  LAYER M2 ;
        RECT 31.52 22.427 33.92 22.429 ;
  LAYER M2 ;
        RECT 31.52 22.511 33.92 22.513 ;
  LAYER M2 ;
        RECT 31.52 22.595 33.92 22.597 ;
  LAYER M2 ;
        RECT 31.52 22.679 33.92 22.681 ;
  LAYER M2 ;
        RECT 31.52 22.763 33.92 22.765 ;
  LAYER M2 ;
        RECT 31.52 22.847 33.92 22.849 ;
  LAYER M2 ;
        RECT 31.52 22.931 33.92 22.933 ;
  LAYER M2 ;
        RECT 31.52 23.015 33.92 23.017 ;
  LAYER M2 ;
        RECT 31.52 23.099 33.92 23.101 ;
  LAYER M2 ;
        RECT 31.52 23.183 33.92 23.185 ;
  LAYER M2 ;
        RECT 31.52 23.267 33.92 23.269 ;
  LAYER M1 ;
        RECT 33.904 23.82 33.936 26.328 ;
  LAYER M1 ;
        RECT 33.84 23.82 33.872 26.328 ;
  LAYER M1 ;
        RECT 33.776 23.82 33.808 26.328 ;
  LAYER M1 ;
        RECT 33.712 23.82 33.744 26.328 ;
  LAYER M1 ;
        RECT 33.648 23.82 33.68 26.328 ;
  LAYER M1 ;
        RECT 33.584 23.82 33.616 26.328 ;
  LAYER M1 ;
        RECT 33.52 23.82 33.552 26.328 ;
  LAYER M1 ;
        RECT 33.456 23.82 33.488 26.328 ;
  LAYER M1 ;
        RECT 33.392 23.82 33.424 26.328 ;
  LAYER M1 ;
        RECT 33.328 23.82 33.36 26.328 ;
  LAYER M1 ;
        RECT 33.264 23.82 33.296 26.328 ;
  LAYER M1 ;
        RECT 33.2 23.82 33.232 26.328 ;
  LAYER M1 ;
        RECT 33.136 23.82 33.168 26.328 ;
  LAYER M1 ;
        RECT 33.072 23.82 33.104 26.328 ;
  LAYER M1 ;
        RECT 33.008 23.82 33.04 26.328 ;
  LAYER M1 ;
        RECT 32.944 23.82 32.976 26.328 ;
  LAYER M1 ;
        RECT 32.88 23.82 32.912 26.328 ;
  LAYER M1 ;
        RECT 32.816 23.82 32.848 26.328 ;
  LAYER M1 ;
        RECT 32.752 23.82 32.784 26.328 ;
  LAYER M1 ;
        RECT 32.688 23.82 32.72 26.328 ;
  LAYER M1 ;
        RECT 32.624 23.82 32.656 26.328 ;
  LAYER M1 ;
        RECT 32.56 23.82 32.592 26.328 ;
  LAYER M1 ;
        RECT 32.496 23.82 32.528 26.328 ;
  LAYER M1 ;
        RECT 32.432 23.82 32.464 26.328 ;
  LAYER M1 ;
        RECT 32.368 23.82 32.4 26.328 ;
  LAYER M1 ;
        RECT 32.304 23.82 32.336 26.328 ;
  LAYER M1 ;
        RECT 32.24 23.82 32.272 26.328 ;
  LAYER M1 ;
        RECT 32.176 23.82 32.208 26.328 ;
  LAYER M1 ;
        RECT 32.112 23.82 32.144 26.328 ;
  LAYER M1 ;
        RECT 32.048 23.82 32.08 26.328 ;
  LAYER M1 ;
        RECT 31.984 23.82 32.016 26.328 ;
  LAYER M1 ;
        RECT 31.92 23.82 31.952 26.328 ;
  LAYER M1 ;
        RECT 31.856 23.82 31.888 26.328 ;
  LAYER M1 ;
        RECT 31.792 23.82 31.824 26.328 ;
  LAYER M1 ;
        RECT 31.728 23.82 31.76 26.328 ;
  LAYER M1 ;
        RECT 31.664 23.82 31.696 26.328 ;
  LAYER M1 ;
        RECT 31.6 23.82 31.632 26.328 ;
  LAYER M2 ;
        RECT 31.484 23.904 33.956 23.936 ;
  LAYER M2 ;
        RECT 31.484 23.968 33.956 24 ;
  LAYER M2 ;
        RECT 31.484 24.032 33.956 24.064 ;
  LAYER M2 ;
        RECT 31.484 24.096 33.956 24.128 ;
  LAYER M2 ;
        RECT 31.484 24.16 33.956 24.192 ;
  LAYER M2 ;
        RECT 31.484 24.224 33.956 24.256 ;
  LAYER M2 ;
        RECT 31.484 24.288 33.956 24.32 ;
  LAYER M2 ;
        RECT 31.484 24.352 33.956 24.384 ;
  LAYER M2 ;
        RECT 31.484 24.416 33.956 24.448 ;
  LAYER M2 ;
        RECT 31.484 24.48 33.956 24.512 ;
  LAYER M2 ;
        RECT 31.484 24.544 33.956 24.576 ;
  LAYER M2 ;
        RECT 31.484 24.608 33.956 24.64 ;
  LAYER M2 ;
        RECT 31.484 24.672 33.956 24.704 ;
  LAYER M2 ;
        RECT 31.484 24.736 33.956 24.768 ;
  LAYER M2 ;
        RECT 31.484 24.8 33.956 24.832 ;
  LAYER M2 ;
        RECT 31.484 24.864 33.956 24.896 ;
  LAYER M2 ;
        RECT 31.484 24.928 33.956 24.96 ;
  LAYER M2 ;
        RECT 31.484 24.992 33.956 25.024 ;
  LAYER M2 ;
        RECT 31.484 25.056 33.956 25.088 ;
  LAYER M2 ;
        RECT 31.484 25.12 33.956 25.152 ;
  LAYER M2 ;
        RECT 31.484 25.184 33.956 25.216 ;
  LAYER M2 ;
        RECT 31.484 25.248 33.956 25.28 ;
  LAYER M2 ;
        RECT 31.484 25.312 33.956 25.344 ;
  LAYER M2 ;
        RECT 31.484 25.376 33.956 25.408 ;
  LAYER M2 ;
        RECT 31.484 25.44 33.956 25.472 ;
  LAYER M2 ;
        RECT 31.484 25.504 33.956 25.536 ;
  LAYER M2 ;
        RECT 31.484 25.568 33.956 25.6 ;
  LAYER M2 ;
        RECT 31.484 25.632 33.956 25.664 ;
  LAYER M2 ;
        RECT 31.484 25.696 33.956 25.728 ;
  LAYER M2 ;
        RECT 31.484 25.76 33.956 25.792 ;
  LAYER M2 ;
        RECT 31.484 25.824 33.956 25.856 ;
  LAYER M2 ;
        RECT 31.484 25.888 33.956 25.92 ;
  LAYER M2 ;
        RECT 31.484 25.952 33.956 25.984 ;
  LAYER M2 ;
        RECT 31.484 26.016 33.956 26.048 ;
  LAYER M2 ;
        RECT 31.484 26.08 33.956 26.112 ;
  LAYER M2 ;
        RECT 31.484 26.144 33.956 26.176 ;
  LAYER M3 ;
        RECT 33.904 23.82 33.936 26.328 ;
  LAYER M3 ;
        RECT 33.84 23.82 33.872 26.328 ;
  LAYER M3 ;
        RECT 33.776 23.82 33.808 26.328 ;
  LAYER M3 ;
        RECT 33.712 23.82 33.744 26.328 ;
  LAYER M3 ;
        RECT 33.648 23.82 33.68 26.328 ;
  LAYER M3 ;
        RECT 33.584 23.82 33.616 26.328 ;
  LAYER M3 ;
        RECT 33.52 23.82 33.552 26.328 ;
  LAYER M3 ;
        RECT 33.456 23.82 33.488 26.328 ;
  LAYER M3 ;
        RECT 33.392 23.82 33.424 26.328 ;
  LAYER M3 ;
        RECT 33.328 23.82 33.36 26.328 ;
  LAYER M3 ;
        RECT 33.264 23.82 33.296 26.328 ;
  LAYER M3 ;
        RECT 33.2 23.82 33.232 26.328 ;
  LAYER M3 ;
        RECT 33.136 23.82 33.168 26.328 ;
  LAYER M3 ;
        RECT 33.072 23.82 33.104 26.328 ;
  LAYER M3 ;
        RECT 33.008 23.82 33.04 26.328 ;
  LAYER M3 ;
        RECT 32.944 23.82 32.976 26.328 ;
  LAYER M3 ;
        RECT 32.88 23.82 32.912 26.328 ;
  LAYER M3 ;
        RECT 32.816 23.82 32.848 26.328 ;
  LAYER M3 ;
        RECT 32.752 23.82 32.784 26.328 ;
  LAYER M3 ;
        RECT 32.688 23.82 32.72 26.328 ;
  LAYER M3 ;
        RECT 32.624 23.82 32.656 26.328 ;
  LAYER M3 ;
        RECT 32.56 23.82 32.592 26.328 ;
  LAYER M3 ;
        RECT 32.496 23.82 32.528 26.328 ;
  LAYER M3 ;
        RECT 32.432 23.82 32.464 26.328 ;
  LAYER M3 ;
        RECT 32.368 23.82 32.4 26.328 ;
  LAYER M3 ;
        RECT 32.304 23.82 32.336 26.328 ;
  LAYER M3 ;
        RECT 32.24 23.82 32.272 26.328 ;
  LAYER M3 ;
        RECT 32.176 23.82 32.208 26.328 ;
  LAYER M3 ;
        RECT 32.112 23.82 32.144 26.328 ;
  LAYER M3 ;
        RECT 32.048 23.82 32.08 26.328 ;
  LAYER M3 ;
        RECT 31.984 23.82 32.016 26.328 ;
  LAYER M3 ;
        RECT 31.92 23.82 31.952 26.328 ;
  LAYER M3 ;
        RECT 31.856 23.82 31.888 26.328 ;
  LAYER M3 ;
        RECT 31.792 23.82 31.824 26.328 ;
  LAYER M3 ;
        RECT 31.728 23.82 31.76 26.328 ;
  LAYER M3 ;
        RECT 31.664 23.82 31.696 26.328 ;
  LAYER M3 ;
        RECT 31.6 23.82 31.632 26.328 ;
  LAYER M3 ;
        RECT 31.504 23.82 31.536 26.328 ;
  LAYER M1 ;
        RECT 33.919 23.856 33.921 26.292 ;
  LAYER M1 ;
        RECT 33.839 23.856 33.841 26.292 ;
  LAYER M1 ;
        RECT 33.759 23.856 33.761 26.292 ;
  LAYER M1 ;
        RECT 33.679 23.856 33.681 26.292 ;
  LAYER M1 ;
        RECT 33.599 23.856 33.601 26.292 ;
  LAYER M1 ;
        RECT 33.519 23.856 33.521 26.292 ;
  LAYER M1 ;
        RECT 33.439 23.856 33.441 26.292 ;
  LAYER M1 ;
        RECT 33.359 23.856 33.361 26.292 ;
  LAYER M1 ;
        RECT 33.279 23.856 33.281 26.292 ;
  LAYER M1 ;
        RECT 33.199 23.856 33.201 26.292 ;
  LAYER M1 ;
        RECT 33.119 23.856 33.121 26.292 ;
  LAYER M1 ;
        RECT 33.039 23.856 33.041 26.292 ;
  LAYER M1 ;
        RECT 32.959 23.856 32.961 26.292 ;
  LAYER M1 ;
        RECT 32.879 23.856 32.881 26.292 ;
  LAYER M1 ;
        RECT 32.799 23.856 32.801 26.292 ;
  LAYER M1 ;
        RECT 32.719 23.856 32.721 26.292 ;
  LAYER M1 ;
        RECT 32.639 23.856 32.641 26.292 ;
  LAYER M1 ;
        RECT 32.559 23.856 32.561 26.292 ;
  LAYER M1 ;
        RECT 32.479 23.856 32.481 26.292 ;
  LAYER M1 ;
        RECT 32.399 23.856 32.401 26.292 ;
  LAYER M1 ;
        RECT 32.319 23.856 32.321 26.292 ;
  LAYER M1 ;
        RECT 32.239 23.856 32.241 26.292 ;
  LAYER M1 ;
        RECT 32.159 23.856 32.161 26.292 ;
  LAYER M1 ;
        RECT 32.079 23.856 32.081 26.292 ;
  LAYER M1 ;
        RECT 31.999 23.856 32.001 26.292 ;
  LAYER M1 ;
        RECT 31.919 23.856 31.921 26.292 ;
  LAYER M1 ;
        RECT 31.839 23.856 31.841 26.292 ;
  LAYER M1 ;
        RECT 31.759 23.856 31.761 26.292 ;
  LAYER M1 ;
        RECT 31.679 23.856 31.681 26.292 ;
  LAYER M1 ;
        RECT 31.599 23.856 31.601 26.292 ;
  LAYER M2 ;
        RECT 31.52 23.855 33.92 23.857 ;
  LAYER M2 ;
        RECT 31.52 23.939 33.92 23.941 ;
  LAYER M2 ;
        RECT 31.52 24.023 33.92 24.025 ;
  LAYER M2 ;
        RECT 31.52 24.107 33.92 24.109 ;
  LAYER M2 ;
        RECT 31.52 24.191 33.92 24.193 ;
  LAYER M2 ;
        RECT 31.52 24.275 33.92 24.277 ;
  LAYER M2 ;
        RECT 31.52 24.359 33.92 24.361 ;
  LAYER M2 ;
        RECT 31.52 24.443 33.92 24.445 ;
  LAYER M2 ;
        RECT 31.52 24.527 33.92 24.529 ;
  LAYER M2 ;
        RECT 31.52 24.611 33.92 24.613 ;
  LAYER M2 ;
        RECT 31.52 24.695 33.92 24.697 ;
  LAYER M2 ;
        RECT 31.52 24.779 33.92 24.781 ;
  LAYER M2 ;
        RECT 31.52 24.8625 33.92 24.8645 ;
  LAYER M2 ;
        RECT 31.52 24.947 33.92 24.949 ;
  LAYER M2 ;
        RECT 31.52 25.031 33.92 25.033 ;
  LAYER M2 ;
        RECT 31.52 25.115 33.92 25.117 ;
  LAYER M2 ;
        RECT 31.52 25.199 33.92 25.201 ;
  LAYER M2 ;
        RECT 31.52 25.283 33.92 25.285 ;
  LAYER M2 ;
        RECT 31.52 25.367 33.92 25.369 ;
  LAYER M2 ;
        RECT 31.52 25.451 33.92 25.453 ;
  LAYER M2 ;
        RECT 31.52 25.535 33.92 25.537 ;
  LAYER M2 ;
        RECT 31.52 25.619 33.92 25.621 ;
  LAYER M2 ;
        RECT 31.52 25.703 33.92 25.705 ;
  LAYER M2 ;
        RECT 31.52 25.787 33.92 25.789 ;
  LAYER M2 ;
        RECT 31.52 25.871 33.92 25.873 ;
  LAYER M2 ;
        RECT 31.52 25.955 33.92 25.957 ;
  LAYER M2 ;
        RECT 31.52 26.039 33.92 26.041 ;
  LAYER M2 ;
        RECT 31.52 26.123 33.92 26.125 ;
  LAYER M2 ;
        RECT 31.52 26.207 33.92 26.209 ;
  LAYER M1 ;
        RECT 33.904 26.76 33.936 29.268 ;
  LAYER M1 ;
        RECT 33.84 26.76 33.872 29.268 ;
  LAYER M1 ;
        RECT 33.776 26.76 33.808 29.268 ;
  LAYER M1 ;
        RECT 33.712 26.76 33.744 29.268 ;
  LAYER M1 ;
        RECT 33.648 26.76 33.68 29.268 ;
  LAYER M1 ;
        RECT 33.584 26.76 33.616 29.268 ;
  LAYER M1 ;
        RECT 33.52 26.76 33.552 29.268 ;
  LAYER M1 ;
        RECT 33.456 26.76 33.488 29.268 ;
  LAYER M1 ;
        RECT 33.392 26.76 33.424 29.268 ;
  LAYER M1 ;
        RECT 33.328 26.76 33.36 29.268 ;
  LAYER M1 ;
        RECT 33.264 26.76 33.296 29.268 ;
  LAYER M1 ;
        RECT 33.2 26.76 33.232 29.268 ;
  LAYER M1 ;
        RECT 33.136 26.76 33.168 29.268 ;
  LAYER M1 ;
        RECT 33.072 26.76 33.104 29.268 ;
  LAYER M1 ;
        RECT 33.008 26.76 33.04 29.268 ;
  LAYER M1 ;
        RECT 32.944 26.76 32.976 29.268 ;
  LAYER M1 ;
        RECT 32.88 26.76 32.912 29.268 ;
  LAYER M1 ;
        RECT 32.816 26.76 32.848 29.268 ;
  LAYER M1 ;
        RECT 32.752 26.76 32.784 29.268 ;
  LAYER M1 ;
        RECT 32.688 26.76 32.72 29.268 ;
  LAYER M1 ;
        RECT 32.624 26.76 32.656 29.268 ;
  LAYER M1 ;
        RECT 32.56 26.76 32.592 29.268 ;
  LAYER M1 ;
        RECT 32.496 26.76 32.528 29.268 ;
  LAYER M1 ;
        RECT 32.432 26.76 32.464 29.268 ;
  LAYER M1 ;
        RECT 32.368 26.76 32.4 29.268 ;
  LAYER M1 ;
        RECT 32.304 26.76 32.336 29.268 ;
  LAYER M1 ;
        RECT 32.24 26.76 32.272 29.268 ;
  LAYER M1 ;
        RECT 32.176 26.76 32.208 29.268 ;
  LAYER M1 ;
        RECT 32.112 26.76 32.144 29.268 ;
  LAYER M1 ;
        RECT 32.048 26.76 32.08 29.268 ;
  LAYER M1 ;
        RECT 31.984 26.76 32.016 29.268 ;
  LAYER M1 ;
        RECT 31.92 26.76 31.952 29.268 ;
  LAYER M1 ;
        RECT 31.856 26.76 31.888 29.268 ;
  LAYER M1 ;
        RECT 31.792 26.76 31.824 29.268 ;
  LAYER M1 ;
        RECT 31.728 26.76 31.76 29.268 ;
  LAYER M1 ;
        RECT 31.664 26.76 31.696 29.268 ;
  LAYER M1 ;
        RECT 31.6 26.76 31.632 29.268 ;
  LAYER M2 ;
        RECT 31.484 26.844 33.956 26.876 ;
  LAYER M2 ;
        RECT 31.484 26.908 33.956 26.94 ;
  LAYER M2 ;
        RECT 31.484 26.972 33.956 27.004 ;
  LAYER M2 ;
        RECT 31.484 27.036 33.956 27.068 ;
  LAYER M2 ;
        RECT 31.484 27.1 33.956 27.132 ;
  LAYER M2 ;
        RECT 31.484 27.164 33.956 27.196 ;
  LAYER M2 ;
        RECT 31.484 27.228 33.956 27.26 ;
  LAYER M2 ;
        RECT 31.484 27.292 33.956 27.324 ;
  LAYER M2 ;
        RECT 31.484 27.356 33.956 27.388 ;
  LAYER M2 ;
        RECT 31.484 27.42 33.956 27.452 ;
  LAYER M2 ;
        RECT 31.484 27.484 33.956 27.516 ;
  LAYER M2 ;
        RECT 31.484 27.548 33.956 27.58 ;
  LAYER M2 ;
        RECT 31.484 27.612 33.956 27.644 ;
  LAYER M2 ;
        RECT 31.484 27.676 33.956 27.708 ;
  LAYER M2 ;
        RECT 31.484 27.74 33.956 27.772 ;
  LAYER M2 ;
        RECT 31.484 27.804 33.956 27.836 ;
  LAYER M2 ;
        RECT 31.484 27.868 33.956 27.9 ;
  LAYER M2 ;
        RECT 31.484 27.932 33.956 27.964 ;
  LAYER M2 ;
        RECT 31.484 27.996 33.956 28.028 ;
  LAYER M2 ;
        RECT 31.484 28.06 33.956 28.092 ;
  LAYER M2 ;
        RECT 31.484 28.124 33.956 28.156 ;
  LAYER M2 ;
        RECT 31.484 28.188 33.956 28.22 ;
  LAYER M2 ;
        RECT 31.484 28.252 33.956 28.284 ;
  LAYER M2 ;
        RECT 31.484 28.316 33.956 28.348 ;
  LAYER M2 ;
        RECT 31.484 28.38 33.956 28.412 ;
  LAYER M2 ;
        RECT 31.484 28.444 33.956 28.476 ;
  LAYER M2 ;
        RECT 31.484 28.508 33.956 28.54 ;
  LAYER M2 ;
        RECT 31.484 28.572 33.956 28.604 ;
  LAYER M2 ;
        RECT 31.484 28.636 33.956 28.668 ;
  LAYER M2 ;
        RECT 31.484 28.7 33.956 28.732 ;
  LAYER M2 ;
        RECT 31.484 28.764 33.956 28.796 ;
  LAYER M2 ;
        RECT 31.484 28.828 33.956 28.86 ;
  LAYER M2 ;
        RECT 31.484 28.892 33.956 28.924 ;
  LAYER M2 ;
        RECT 31.484 28.956 33.956 28.988 ;
  LAYER M2 ;
        RECT 31.484 29.02 33.956 29.052 ;
  LAYER M2 ;
        RECT 31.484 29.084 33.956 29.116 ;
  LAYER M3 ;
        RECT 33.904 26.76 33.936 29.268 ;
  LAYER M3 ;
        RECT 33.84 26.76 33.872 29.268 ;
  LAYER M3 ;
        RECT 33.776 26.76 33.808 29.268 ;
  LAYER M3 ;
        RECT 33.712 26.76 33.744 29.268 ;
  LAYER M3 ;
        RECT 33.648 26.76 33.68 29.268 ;
  LAYER M3 ;
        RECT 33.584 26.76 33.616 29.268 ;
  LAYER M3 ;
        RECT 33.52 26.76 33.552 29.268 ;
  LAYER M3 ;
        RECT 33.456 26.76 33.488 29.268 ;
  LAYER M3 ;
        RECT 33.392 26.76 33.424 29.268 ;
  LAYER M3 ;
        RECT 33.328 26.76 33.36 29.268 ;
  LAYER M3 ;
        RECT 33.264 26.76 33.296 29.268 ;
  LAYER M3 ;
        RECT 33.2 26.76 33.232 29.268 ;
  LAYER M3 ;
        RECT 33.136 26.76 33.168 29.268 ;
  LAYER M3 ;
        RECT 33.072 26.76 33.104 29.268 ;
  LAYER M3 ;
        RECT 33.008 26.76 33.04 29.268 ;
  LAYER M3 ;
        RECT 32.944 26.76 32.976 29.268 ;
  LAYER M3 ;
        RECT 32.88 26.76 32.912 29.268 ;
  LAYER M3 ;
        RECT 32.816 26.76 32.848 29.268 ;
  LAYER M3 ;
        RECT 32.752 26.76 32.784 29.268 ;
  LAYER M3 ;
        RECT 32.688 26.76 32.72 29.268 ;
  LAYER M3 ;
        RECT 32.624 26.76 32.656 29.268 ;
  LAYER M3 ;
        RECT 32.56 26.76 32.592 29.268 ;
  LAYER M3 ;
        RECT 32.496 26.76 32.528 29.268 ;
  LAYER M3 ;
        RECT 32.432 26.76 32.464 29.268 ;
  LAYER M3 ;
        RECT 32.368 26.76 32.4 29.268 ;
  LAYER M3 ;
        RECT 32.304 26.76 32.336 29.268 ;
  LAYER M3 ;
        RECT 32.24 26.76 32.272 29.268 ;
  LAYER M3 ;
        RECT 32.176 26.76 32.208 29.268 ;
  LAYER M3 ;
        RECT 32.112 26.76 32.144 29.268 ;
  LAYER M3 ;
        RECT 32.048 26.76 32.08 29.268 ;
  LAYER M3 ;
        RECT 31.984 26.76 32.016 29.268 ;
  LAYER M3 ;
        RECT 31.92 26.76 31.952 29.268 ;
  LAYER M3 ;
        RECT 31.856 26.76 31.888 29.268 ;
  LAYER M3 ;
        RECT 31.792 26.76 31.824 29.268 ;
  LAYER M3 ;
        RECT 31.728 26.76 31.76 29.268 ;
  LAYER M3 ;
        RECT 31.664 26.76 31.696 29.268 ;
  LAYER M3 ;
        RECT 31.6 26.76 31.632 29.268 ;
  LAYER M3 ;
        RECT 31.504 26.76 31.536 29.268 ;
  LAYER M1 ;
        RECT 33.919 26.796 33.921 29.232 ;
  LAYER M1 ;
        RECT 33.839 26.796 33.841 29.232 ;
  LAYER M1 ;
        RECT 33.759 26.796 33.761 29.232 ;
  LAYER M1 ;
        RECT 33.679 26.796 33.681 29.232 ;
  LAYER M1 ;
        RECT 33.599 26.796 33.601 29.232 ;
  LAYER M1 ;
        RECT 33.519 26.796 33.521 29.232 ;
  LAYER M1 ;
        RECT 33.439 26.796 33.441 29.232 ;
  LAYER M1 ;
        RECT 33.359 26.796 33.361 29.232 ;
  LAYER M1 ;
        RECT 33.279 26.796 33.281 29.232 ;
  LAYER M1 ;
        RECT 33.199 26.796 33.201 29.232 ;
  LAYER M1 ;
        RECT 33.119 26.796 33.121 29.232 ;
  LAYER M1 ;
        RECT 33.039 26.796 33.041 29.232 ;
  LAYER M1 ;
        RECT 32.959 26.796 32.961 29.232 ;
  LAYER M1 ;
        RECT 32.879 26.796 32.881 29.232 ;
  LAYER M1 ;
        RECT 32.799 26.796 32.801 29.232 ;
  LAYER M1 ;
        RECT 32.719 26.796 32.721 29.232 ;
  LAYER M1 ;
        RECT 32.639 26.796 32.641 29.232 ;
  LAYER M1 ;
        RECT 32.559 26.796 32.561 29.232 ;
  LAYER M1 ;
        RECT 32.479 26.796 32.481 29.232 ;
  LAYER M1 ;
        RECT 32.399 26.796 32.401 29.232 ;
  LAYER M1 ;
        RECT 32.319 26.796 32.321 29.232 ;
  LAYER M1 ;
        RECT 32.239 26.796 32.241 29.232 ;
  LAYER M1 ;
        RECT 32.159 26.796 32.161 29.232 ;
  LAYER M1 ;
        RECT 32.079 26.796 32.081 29.232 ;
  LAYER M1 ;
        RECT 31.999 26.796 32.001 29.232 ;
  LAYER M1 ;
        RECT 31.919 26.796 31.921 29.232 ;
  LAYER M1 ;
        RECT 31.839 26.796 31.841 29.232 ;
  LAYER M1 ;
        RECT 31.759 26.796 31.761 29.232 ;
  LAYER M1 ;
        RECT 31.679 26.796 31.681 29.232 ;
  LAYER M1 ;
        RECT 31.599 26.796 31.601 29.232 ;
  LAYER M2 ;
        RECT 31.52 26.795 33.92 26.797 ;
  LAYER M2 ;
        RECT 31.52 26.879 33.92 26.881 ;
  LAYER M2 ;
        RECT 31.52 26.963 33.92 26.965 ;
  LAYER M2 ;
        RECT 31.52 27.047 33.92 27.049 ;
  LAYER M2 ;
        RECT 31.52 27.131 33.92 27.133 ;
  LAYER M2 ;
        RECT 31.52 27.215 33.92 27.217 ;
  LAYER M2 ;
        RECT 31.52 27.299 33.92 27.301 ;
  LAYER M2 ;
        RECT 31.52 27.383 33.92 27.385 ;
  LAYER M2 ;
        RECT 31.52 27.467 33.92 27.469 ;
  LAYER M2 ;
        RECT 31.52 27.551 33.92 27.553 ;
  LAYER M2 ;
        RECT 31.52 27.635 33.92 27.637 ;
  LAYER M2 ;
        RECT 31.52 27.719 33.92 27.721 ;
  LAYER M2 ;
        RECT 31.52 27.8025 33.92 27.8045 ;
  LAYER M2 ;
        RECT 31.52 27.887 33.92 27.889 ;
  LAYER M2 ;
        RECT 31.52 27.971 33.92 27.973 ;
  LAYER M2 ;
        RECT 31.52 28.055 33.92 28.057 ;
  LAYER M2 ;
        RECT 31.52 28.139 33.92 28.141 ;
  LAYER M2 ;
        RECT 31.52 28.223 33.92 28.225 ;
  LAYER M2 ;
        RECT 31.52 28.307 33.92 28.309 ;
  LAYER M2 ;
        RECT 31.52 28.391 33.92 28.393 ;
  LAYER M2 ;
        RECT 31.52 28.475 33.92 28.477 ;
  LAYER M2 ;
        RECT 31.52 28.559 33.92 28.561 ;
  LAYER M2 ;
        RECT 31.52 28.643 33.92 28.645 ;
  LAYER M2 ;
        RECT 31.52 28.727 33.92 28.729 ;
  LAYER M2 ;
        RECT 31.52 28.811 33.92 28.813 ;
  LAYER M2 ;
        RECT 31.52 28.895 33.92 28.897 ;
  LAYER M2 ;
        RECT 31.52 28.979 33.92 28.981 ;
  LAYER M2 ;
        RECT 31.52 29.063 33.92 29.065 ;
  LAYER M2 ;
        RECT 31.52 29.147 33.92 29.149 ;
  LAYER M1 ;
        RECT 40.944 0.3 40.976 0.96 ;
  LAYER M1 ;
        RECT 41.024 0.3 41.056 0.96 ;
  LAYER M1 ;
        RECT 40.864 0.3 40.896 0.96 ;
  LAYER M2 ;
        RECT 40.844 0.908 41.156 0.94 ;
  LAYER M2 ;
        RECT 40.844 0.656 41.156 0.688 ;
  LAYER M2 ;
        RECT 40.764 0.824 41.076 0.856 ;
  LAYER M2 ;
        RECT 40.764 0.572 41.076 0.604 ;
  LAYER M2 ;
        RECT 40.684 0.74 41.076 0.772 ;
  LAYER M2 ;
        RECT 40.684 0.488 41.076 0.52 ;
  LAYER M1 ;
        RECT 30.864 17.352 30.896 18.012 ;
  LAYER M1 ;
        RECT 30.944 17.352 30.976 18.012 ;
  LAYER M1 ;
        RECT 30.784 17.352 30.816 18.012 ;
  LAYER M2 ;
        RECT 30.764 17.96 31.076 17.992 ;
  LAYER M2 ;
        RECT 30.764 17.708 31.076 17.74 ;
  LAYER M2 ;
        RECT 30.684 17.876 30.996 17.908 ;
  LAYER M2 ;
        RECT 30.684 17.624 30.996 17.656 ;
  LAYER M2 ;
        RECT 30.604 17.792 30.996 17.824 ;
  LAYER M2 ;
        RECT 30.604 17.54 30.996 17.572 ;
  LAYER M1 ;
        RECT 39.584 0.3 39.616 0.96 ;
  LAYER M1 ;
        RECT 39.504 0.3 39.536 0.96 ;
  LAYER M1 ;
        RECT 39.664 0.3 39.696 0.96 ;
  LAYER M1 ;
        RECT 40.224 0.3 40.256 0.96 ;
  LAYER M1 ;
        RECT 40.144 0.3 40.176 0.96 ;
  LAYER M1 ;
        RECT 40.304 0.3 40.336 0.96 ;
  LAYER M1 ;
        RECT 38.864 0.3 38.896 0.96 ;
  LAYER M1 ;
        RECT 38.944 0.3 38.976 0.96 ;
  LAYER M1 ;
        RECT 38.784 0.3 38.816 0.96 ;
  LAYER M1 ;
        RECT 38.224 0.3 38.256 0.96 ;
  LAYER M1 ;
        RECT 38.304 0.3 38.336 0.96 ;
  LAYER M1 ;
        RECT 38.144 0.3 38.176 0.96 ;
  LAYER M1 ;
        RECT 37.344 10.296 37.376 10.368 ;
  LAYER M2 ;
        RECT 37.324 10.316 37.396 10.348 ;
  LAYER M2 ;
        RECT 37.04 10.316 37.36 10.348 ;
  LAYER M1 ;
        RECT 37.024 10.296 37.056 10.368 ;
  LAYER M2 ;
        RECT 37.004 10.316 37.076 10.348 ;
  LAYER M1 ;
        RECT 34.464 7.356 34.496 7.428 ;
  LAYER M2 ;
        RECT 34.444 7.376 34.516 7.408 ;
  LAYER M1 ;
        RECT 34.464 7.392 34.496 7.56 ;
  LAYER M1 ;
        RECT 34.464 7.524 34.496 7.596 ;
  LAYER M2 ;
        RECT 34.444 7.544 34.516 7.576 ;
  LAYER M2 ;
        RECT 34.48 7.544 37.04 7.576 ;
  LAYER M1 ;
        RECT 37.024 7.524 37.056 7.596 ;
  LAYER M2 ;
        RECT 37.004 7.544 37.076 7.576 ;
  LAYER M1 ;
        RECT 37.024 16.68 37.056 16.752 ;
  LAYER M2 ;
        RECT 37.004 16.7 37.076 16.732 ;
  LAYER M1 ;
        RECT 37.024 16.548 37.056 16.716 ;
  LAYER M1 ;
        RECT 37.024 7.56 37.056 16.548 ;
  LAYER M1 ;
        RECT 40.224 13.236 40.256 13.308 ;
  LAYER M2 ;
        RECT 40.204 13.256 40.276 13.288 ;
  LAYER M2 ;
        RECT 39.92 13.256 40.24 13.288 ;
  LAYER M1 ;
        RECT 39.904 13.236 39.936 13.308 ;
  LAYER M2 ;
        RECT 39.884 13.256 39.956 13.288 ;
  LAYER M1 ;
        RECT 39.904 16.68 39.936 16.752 ;
  LAYER M2 ;
        RECT 39.884 16.7 39.956 16.732 ;
  LAYER M1 ;
        RECT 39.904 16.548 39.936 16.716 ;
  LAYER M1 ;
        RECT 39.904 13.272 39.936 16.548 ;
  LAYER M2 ;
        RECT 37.04 16.7 39.92 16.732 ;
  LAYER M1 ;
        RECT 34.464 10.296 34.496 10.368 ;
  LAYER M2 ;
        RECT 34.444 10.316 34.516 10.348 ;
  LAYER M2 ;
        RECT 34.16 10.316 34.48 10.348 ;
  LAYER M1 ;
        RECT 34.144 10.296 34.176 10.368 ;
  LAYER M2 ;
        RECT 34.124 10.316 34.196 10.348 ;
  LAYER M1 ;
        RECT 34.464 13.236 34.496 13.308 ;
  LAYER M2 ;
        RECT 34.444 13.256 34.516 13.288 ;
  LAYER M2 ;
        RECT 34.16 13.256 34.48 13.288 ;
  LAYER M1 ;
        RECT 34.144 13.236 34.176 13.308 ;
  LAYER M2 ;
        RECT 34.124 13.256 34.196 13.288 ;
  LAYER M1 ;
        RECT 34.144 16.848 34.176 16.92 ;
  LAYER M2 ;
        RECT 34.124 16.868 34.196 16.9 ;
  LAYER M1 ;
        RECT 34.144 16.548 34.176 16.884 ;
  LAYER M1 ;
        RECT 34.144 10.332 34.176 16.548 ;
  LAYER M1 ;
        RECT 40.224 10.296 40.256 10.368 ;
  LAYER M2 ;
        RECT 40.204 10.316 40.276 10.348 ;
  LAYER M1 ;
        RECT 40.224 10.332 40.256 10.5 ;
  LAYER M1 ;
        RECT 40.224 10.464 40.256 10.536 ;
  LAYER M2 ;
        RECT 40.204 10.484 40.276 10.516 ;
  LAYER M2 ;
        RECT 40.24 10.484 42.8 10.516 ;
  LAYER M1 ;
        RECT 42.784 10.464 42.816 10.536 ;
  LAYER M2 ;
        RECT 42.764 10.484 42.836 10.516 ;
  LAYER M1 ;
        RECT 40.224 7.356 40.256 7.428 ;
  LAYER M2 ;
        RECT 40.204 7.376 40.276 7.408 ;
  LAYER M1 ;
        RECT 40.224 7.392 40.256 7.56 ;
  LAYER M1 ;
        RECT 40.224 7.524 40.256 7.596 ;
  LAYER M2 ;
        RECT 40.204 7.544 40.276 7.576 ;
  LAYER M2 ;
        RECT 40.24 7.544 42.8 7.576 ;
  LAYER M1 ;
        RECT 42.784 7.524 42.816 7.596 ;
  LAYER M2 ;
        RECT 42.764 7.544 42.836 7.576 ;
  LAYER M1 ;
        RECT 42.784 16.848 42.816 16.92 ;
  LAYER M2 ;
        RECT 42.764 16.868 42.836 16.9 ;
  LAYER M1 ;
        RECT 42.784 16.548 42.816 16.884 ;
  LAYER M1 ;
        RECT 42.784 7.56 42.816 16.548 ;
  LAYER M2 ;
        RECT 34.16 16.868 42.8 16.9 ;
  LAYER M1 ;
        RECT 37.344 13.236 37.376 13.308 ;
  LAYER M2 ;
        RECT 37.324 13.256 37.396 13.288 ;
  LAYER M2 ;
        RECT 34.48 13.256 37.36 13.288 ;
  LAYER M1 ;
        RECT 34.464 13.236 34.496 13.308 ;
  LAYER M2 ;
        RECT 34.444 13.256 34.516 13.288 ;
  LAYER M1 ;
        RECT 37.344 7.356 37.376 7.428 ;
  LAYER M2 ;
        RECT 37.324 7.376 37.396 7.408 ;
  LAYER M2 ;
        RECT 37.36 7.376 40.24 7.408 ;
  LAYER M1 ;
        RECT 40.224 7.356 40.256 7.428 ;
  LAYER M2 ;
        RECT 40.204 7.376 40.276 7.408 ;
  LAYER M1 ;
        RECT 31.584 16.176 31.616 16.248 ;
  LAYER M2 ;
        RECT 31.564 16.196 31.636 16.228 ;
  LAYER M2 ;
        RECT 31.28 16.196 31.6 16.228 ;
  LAYER M1 ;
        RECT 31.264 16.176 31.296 16.248 ;
  LAYER M2 ;
        RECT 31.244 16.196 31.316 16.228 ;
  LAYER M1 ;
        RECT 31.584 13.236 31.616 13.308 ;
  LAYER M2 ;
        RECT 31.564 13.256 31.636 13.288 ;
  LAYER M2 ;
        RECT 31.28 13.256 31.6 13.288 ;
  LAYER M1 ;
        RECT 31.264 13.236 31.296 13.308 ;
  LAYER M2 ;
        RECT 31.244 13.256 31.316 13.288 ;
  LAYER M1 ;
        RECT 31.584 10.296 31.616 10.368 ;
  LAYER M2 ;
        RECT 31.564 10.316 31.636 10.348 ;
  LAYER M2 ;
        RECT 31.28 10.316 31.6 10.348 ;
  LAYER M1 ;
        RECT 31.264 10.296 31.296 10.368 ;
  LAYER M2 ;
        RECT 31.244 10.316 31.316 10.348 ;
  LAYER M1 ;
        RECT 31.584 7.356 31.616 7.428 ;
  LAYER M2 ;
        RECT 31.564 7.376 31.636 7.408 ;
  LAYER M2 ;
        RECT 31.28 7.376 31.6 7.408 ;
  LAYER M1 ;
        RECT 31.264 7.356 31.296 7.428 ;
  LAYER M2 ;
        RECT 31.244 7.376 31.316 7.408 ;
  LAYER M1 ;
        RECT 31.584 4.416 31.616 4.488 ;
  LAYER M2 ;
        RECT 31.564 4.436 31.636 4.468 ;
  LAYER M2 ;
        RECT 31.28 4.436 31.6 4.468 ;
  LAYER M1 ;
        RECT 31.264 4.416 31.296 4.488 ;
  LAYER M2 ;
        RECT 31.244 4.436 31.316 4.468 ;
  LAYER M1 ;
        RECT 31.264 17.016 31.296 17.088 ;
  LAYER M2 ;
        RECT 31.244 17.036 31.316 17.068 ;
  LAYER M1 ;
        RECT 31.264 16.548 31.296 17.052 ;
  LAYER M1 ;
        RECT 31.264 4.452 31.296 16.548 ;
  LAYER M1 ;
        RECT 43.104 16.176 43.136 16.248 ;
  LAYER M2 ;
        RECT 43.084 16.196 43.156 16.228 ;
  LAYER M1 ;
        RECT 43.104 16.212 43.136 16.38 ;
  LAYER M1 ;
        RECT 43.104 16.344 43.136 16.416 ;
  LAYER M2 ;
        RECT 43.084 16.364 43.156 16.396 ;
  LAYER M2 ;
        RECT 43.12 16.364 45.68 16.396 ;
  LAYER M1 ;
        RECT 45.664 16.344 45.696 16.416 ;
  LAYER M2 ;
        RECT 45.644 16.364 45.716 16.396 ;
  LAYER M1 ;
        RECT 43.104 13.236 43.136 13.308 ;
  LAYER M2 ;
        RECT 43.084 13.256 43.156 13.288 ;
  LAYER M1 ;
        RECT 43.104 13.272 43.136 13.44 ;
  LAYER M1 ;
        RECT 43.104 13.404 43.136 13.476 ;
  LAYER M2 ;
        RECT 43.084 13.424 43.156 13.456 ;
  LAYER M2 ;
        RECT 43.12 13.424 45.68 13.456 ;
  LAYER M1 ;
        RECT 45.664 13.404 45.696 13.476 ;
  LAYER M2 ;
        RECT 45.644 13.424 45.716 13.456 ;
  LAYER M1 ;
        RECT 43.104 10.296 43.136 10.368 ;
  LAYER M2 ;
        RECT 43.084 10.316 43.156 10.348 ;
  LAYER M1 ;
        RECT 43.104 10.332 43.136 10.5 ;
  LAYER M1 ;
        RECT 43.104 10.464 43.136 10.536 ;
  LAYER M2 ;
        RECT 43.084 10.484 43.156 10.516 ;
  LAYER M2 ;
        RECT 43.12 10.484 45.68 10.516 ;
  LAYER M1 ;
        RECT 45.664 10.464 45.696 10.536 ;
  LAYER M2 ;
        RECT 45.644 10.484 45.716 10.516 ;
  LAYER M1 ;
        RECT 43.104 7.356 43.136 7.428 ;
  LAYER M2 ;
        RECT 43.084 7.376 43.156 7.408 ;
  LAYER M1 ;
        RECT 43.104 7.392 43.136 7.56 ;
  LAYER M1 ;
        RECT 43.104 7.524 43.136 7.596 ;
  LAYER M2 ;
        RECT 43.084 7.544 43.156 7.576 ;
  LAYER M2 ;
        RECT 43.12 7.544 45.68 7.576 ;
  LAYER M1 ;
        RECT 45.664 7.524 45.696 7.596 ;
  LAYER M2 ;
        RECT 45.644 7.544 45.716 7.576 ;
  LAYER M1 ;
        RECT 43.104 4.416 43.136 4.488 ;
  LAYER M2 ;
        RECT 43.084 4.436 43.156 4.468 ;
  LAYER M1 ;
        RECT 43.104 4.452 43.136 4.62 ;
  LAYER M1 ;
        RECT 43.104 4.584 43.136 4.656 ;
  LAYER M2 ;
        RECT 43.084 4.604 43.156 4.636 ;
  LAYER M2 ;
        RECT 43.12 4.604 45.68 4.636 ;
  LAYER M1 ;
        RECT 45.664 4.584 45.696 4.656 ;
  LAYER M2 ;
        RECT 45.644 4.604 45.716 4.636 ;
  LAYER M1 ;
        RECT 45.664 17.016 45.696 17.088 ;
  LAYER M2 ;
        RECT 45.644 17.036 45.716 17.068 ;
  LAYER M1 ;
        RECT 45.664 16.548 45.696 17.052 ;
  LAYER M1 ;
        RECT 45.664 4.62 45.696 16.548 ;
  LAYER M2 ;
        RECT 31.28 17.036 45.68 17.068 ;
  LAYER M1 ;
        RECT 34.464 16.176 34.496 16.248 ;
  LAYER M2 ;
        RECT 34.444 16.196 34.516 16.228 ;
  LAYER M2 ;
        RECT 31.6 16.196 34.48 16.228 ;
  LAYER M1 ;
        RECT 31.584 16.176 31.616 16.248 ;
  LAYER M2 ;
        RECT 31.564 16.196 31.636 16.228 ;
  LAYER M1 ;
        RECT 34.464 4.416 34.496 4.488 ;
  LAYER M2 ;
        RECT 34.444 4.436 34.516 4.468 ;
  LAYER M2 ;
        RECT 31.6 4.436 34.48 4.468 ;
  LAYER M1 ;
        RECT 31.584 4.416 31.616 4.488 ;
  LAYER M2 ;
        RECT 31.564 4.436 31.636 4.468 ;
  LAYER M1 ;
        RECT 37.344 4.416 37.376 4.488 ;
  LAYER M2 ;
        RECT 37.324 4.436 37.396 4.468 ;
  LAYER M2 ;
        RECT 34.48 4.436 37.36 4.468 ;
  LAYER M1 ;
        RECT 34.464 4.416 34.496 4.488 ;
  LAYER M2 ;
        RECT 34.444 4.436 34.516 4.468 ;
  LAYER M1 ;
        RECT 40.224 4.416 40.256 4.488 ;
  LAYER M2 ;
        RECT 40.204 4.436 40.276 4.468 ;
  LAYER M2 ;
        RECT 37.36 4.436 40.24 4.468 ;
  LAYER M1 ;
        RECT 37.344 4.416 37.376 4.488 ;
  LAYER M2 ;
        RECT 37.324 4.436 37.396 4.468 ;
  LAYER M1 ;
        RECT 40.224 16.176 40.256 16.248 ;
  LAYER M2 ;
        RECT 40.204 16.196 40.276 16.228 ;
  LAYER M2 ;
        RECT 40.24 16.196 43.12 16.228 ;
  LAYER M1 ;
        RECT 43.104 16.176 43.136 16.248 ;
  LAYER M2 ;
        RECT 43.084 16.196 43.156 16.228 ;
  LAYER M1 ;
        RECT 37.344 16.176 37.376 16.248 ;
  LAYER M2 ;
        RECT 37.324 16.196 37.396 16.228 ;
  LAYER M2 ;
        RECT 37.36 16.196 40.24 16.228 ;
  LAYER M1 ;
        RECT 40.224 16.176 40.256 16.248 ;
  LAYER M2 ;
        RECT 40.204 16.196 40.276 16.228 ;
  LAYER M1 ;
        RECT 39.744 7.86 39.776 7.932 ;
  LAYER M2 ;
        RECT 39.724 7.88 39.796 7.912 ;
  LAYER M2 ;
        RECT 37.2 7.88 39.76 7.912 ;
  LAYER M1 ;
        RECT 37.184 7.86 37.216 7.932 ;
  LAYER M2 ;
        RECT 37.164 7.88 37.236 7.912 ;
  LAYER M1 ;
        RECT 36.864 4.92 36.896 4.992 ;
  LAYER M2 ;
        RECT 36.844 4.94 36.916 4.972 ;
  LAYER M1 ;
        RECT 36.864 4.788 36.896 4.956 ;
  LAYER M1 ;
        RECT 36.864 4.752 36.896 4.824 ;
  LAYER M2 ;
        RECT 36.844 4.772 36.916 4.804 ;
  LAYER M2 ;
        RECT 36.88 4.772 37.2 4.804 ;
  LAYER M1 ;
        RECT 37.184 4.752 37.216 4.824 ;
  LAYER M2 ;
        RECT 37.164 4.772 37.236 4.804 ;
  LAYER M1 ;
        RECT 37.184 1.476 37.216 1.548 ;
  LAYER M2 ;
        RECT 37.164 1.496 37.236 1.528 ;
  LAYER M1 ;
        RECT 37.184 1.512 37.216 1.68 ;
  LAYER M1 ;
        RECT 37.184 1.68 37.216 7.896 ;
  LAYER M1 ;
        RECT 42.624 10.8 42.656 10.872 ;
  LAYER M2 ;
        RECT 42.604 10.82 42.676 10.852 ;
  LAYER M2 ;
        RECT 40.08 10.82 42.64 10.852 ;
  LAYER M1 ;
        RECT 40.064 10.8 40.096 10.872 ;
  LAYER M2 ;
        RECT 40.044 10.82 40.116 10.852 ;
  LAYER M1 ;
        RECT 40.064 1.476 40.096 1.548 ;
  LAYER M2 ;
        RECT 40.044 1.496 40.116 1.528 ;
  LAYER M1 ;
        RECT 40.064 1.512 40.096 1.68 ;
  LAYER M1 ;
        RECT 40.064 1.68 40.096 10.836 ;
  LAYER M2 ;
        RECT 37.2 1.496 40.08 1.528 ;
  LAYER M1 ;
        RECT 36.864 7.86 36.896 7.932 ;
  LAYER M2 ;
        RECT 36.844 7.88 36.916 7.912 ;
  LAYER M2 ;
        RECT 34.32 7.88 36.88 7.912 ;
  LAYER M1 ;
        RECT 34.304 7.86 34.336 7.932 ;
  LAYER M2 ;
        RECT 34.284 7.88 34.356 7.912 ;
  LAYER M1 ;
        RECT 36.864 10.8 36.896 10.872 ;
  LAYER M2 ;
        RECT 36.844 10.82 36.916 10.852 ;
  LAYER M2 ;
        RECT 34.32 10.82 36.88 10.852 ;
  LAYER M1 ;
        RECT 34.304 10.8 34.336 10.872 ;
  LAYER M2 ;
        RECT 34.284 10.82 34.356 10.852 ;
  LAYER M1 ;
        RECT 34.304 1.308 34.336 1.38 ;
  LAYER M2 ;
        RECT 34.284 1.328 34.356 1.36 ;
  LAYER M1 ;
        RECT 34.304 1.344 34.336 1.68 ;
  LAYER M1 ;
        RECT 34.304 1.68 34.336 10.836 ;
  LAYER M1 ;
        RECT 42.624 7.86 42.656 7.932 ;
  LAYER M2 ;
        RECT 42.604 7.88 42.676 7.912 ;
  LAYER M1 ;
        RECT 42.624 7.728 42.656 7.896 ;
  LAYER M1 ;
        RECT 42.624 7.692 42.656 7.764 ;
  LAYER M2 ;
        RECT 42.604 7.712 42.676 7.744 ;
  LAYER M2 ;
        RECT 42.64 7.712 42.96 7.744 ;
  LAYER M1 ;
        RECT 42.944 7.692 42.976 7.764 ;
  LAYER M2 ;
        RECT 42.924 7.712 42.996 7.744 ;
  LAYER M1 ;
        RECT 42.624 4.92 42.656 4.992 ;
  LAYER M2 ;
        RECT 42.604 4.94 42.676 4.972 ;
  LAYER M1 ;
        RECT 42.624 4.788 42.656 4.956 ;
  LAYER M1 ;
        RECT 42.624 4.752 42.656 4.824 ;
  LAYER M2 ;
        RECT 42.604 4.772 42.676 4.804 ;
  LAYER M2 ;
        RECT 42.64 4.772 42.96 4.804 ;
  LAYER M1 ;
        RECT 42.944 4.752 42.976 4.824 ;
  LAYER M2 ;
        RECT 42.924 4.772 42.996 4.804 ;
  LAYER M1 ;
        RECT 42.944 1.308 42.976 1.38 ;
  LAYER M2 ;
        RECT 42.924 1.328 42.996 1.36 ;
  LAYER M1 ;
        RECT 42.944 1.344 42.976 1.68 ;
  LAYER M1 ;
        RECT 42.944 1.68 42.976 7.728 ;
  LAYER M2 ;
        RECT 34.32 1.328 42.96 1.36 ;
  LAYER M1 ;
        RECT 39.744 10.8 39.776 10.872 ;
  LAYER M2 ;
        RECT 39.724 10.82 39.796 10.852 ;
  LAYER M2 ;
        RECT 36.88 10.82 39.76 10.852 ;
  LAYER M1 ;
        RECT 36.864 10.8 36.896 10.872 ;
  LAYER M2 ;
        RECT 36.844 10.82 36.916 10.852 ;
  LAYER M1 ;
        RECT 39.744 4.92 39.776 4.992 ;
  LAYER M2 ;
        RECT 39.724 4.94 39.796 4.972 ;
  LAYER M2 ;
        RECT 39.76 4.94 42.64 4.972 ;
  LAYER M1 ;
        RECT 42.624 4.92 42.656 4.992 ;
  LAYER M2 ;
        RECT 42.604 4.94 42.676 4.972 ;
  LAYER M1 ;
        RECT 33.984 13.74 34.016 13.812 ;
  LAYER M2 ;
        RECT 33.964 13.76 34.036 13.792 ;
  LAYER M2 ;
        RECT 31.44 13.76 34 13.792 ;
  LAYER M1 ;
        RECT 31.424 13.74 31.456 13.812 ;
  LAYER M2 ;
        RECT 31.404 13.76 31.476 13.792 ;
  LAYER M1 ;
        RECT 33.984 10.8 34.016 10.872 ;
  LAYER M2 ;
        RECT 33.964 10.82 34.036 10.852 ;
  LAYER M2 ;
        RECT 31.44 10.82 34 10.852 ;
  LAYER M1 ;
        RECT 31.424 10.8 31.456 10.872 ;
  LAYER M2 ;
        RECT 31.404 10.82 31.476 10.852 ;
  LAYER M1 ;
        RECT 33.984 7.86 34.016 7.932 ;
  LAYER M2 ;
        RECT 33.964 7.88 34.036 7.912 ;
  LAYER M2 ;
        RECT 31.44 7.88 34 7.912 ;
  LAYER M1 ;
        RECT 31.424 7.86 31.456 7.932 ;
  LAYER M2 ;
        RECT 31.404 7.88 31.476 7.912 ;
  LAYER M1 ;
        RECT 33.984 4.92 34.016 4.992 ;
  LAYER M2 ;
        RECT 33.964 4.94 34.036 4.972 ;
  LAYER M2 ;
        RECT 31.44 4.94 34 4.972 ;
  LAYER M1 ;
        RECT 31.424 4.92 31.456 4.992 ;
  LAYER M2 ;
        RECT 31.404 4.94 31.476 4.972 ;
  LAYER M1 ;
        RECT 33.984 1.98 34.016 2.052 ;
  LAYER M2 ;
        RECT 33.964 2 34.036 2.032 ;
  LAYER M2 ;
        RECT 31.44 2 34 2.032 ;
  LAYER M1 ;
        RECT 31.424 1.98 31.456 2.052 ;
  LAYER M2 ;
        RECT 31.404 2 31.476 2.032 ;
  LAYER M1 ;
        RECT 31.424 1.14 31.456 1.212 ;
  LAYER M2 ;
        RECT 31.404 1.16 31.476 1.192 ;
  LAYER M1 ;
        RECT 31.424 1.176 31.456 1.68 ;
  LAYER M1 ;
        RECT 31.424 1.68 31.456 13.776 ;
  LAYER M1 ;
        RECT 45.504 13.74 45.536 13.812 ;
  LAYER M2 ;
        RECT 45.484 13.76 45.556 13.792 ;
  LAYER M1 ;
        RECT 45.504 13.608 45.536 13.776 ;
  LAYER M1 ;
        RECT 45.504 13.572 45.536 13.644 ;
  LAYER M2 ;
        RECT 45.484 13.592 45.556 13.624 ;
  LAYER M2 ;
        RECT 45.52 13.592 45.84 13.624 ;
  LAYER M1 ;
        RECT 45.824 13.572 45.856 13.644 ;
  LAYER M2 ;
        RECT 45.804 13.592 45.876 13.624 ;
  LAYER M1 ;
        RECT 45.504 10.8 45.536 10.872 ;
  LAYER M2 ;
        RECT 45.484 10.82 45.556 10.852 ;
  LAYER M1 ;
        RECT 45.504 10.668 45.536 10.836 ;
  LAYER M1 ;
        RECT 45.504 10.632 45.536 10.704 ;
  LAYER M2 ;
        RECT 45.484 10.652 45.556 10.684 ;
  LAYER M2 ;
        RECT 45.52 10.652 45.84 10.684 ;
  LAYER M1 ;
        RECT 45.824 10.632 45.856 10.704 ;
  LAYER M2 ;
        RECT 45.804 10.652 45.876 10.684 ;
  LAYER M1 ;
        RECT 45.504 7.86 45.536 7.932 ;
  LAYER M2 ;
        RECT 45.484 7.88 45.556 7.912 ;
  LAYER M1 ;
        RECT 45.504 7.728 45.536 7.896 ;
  LAYER M1 ;
        RECT 45.504 7.692 45.536 7.764 ;
  LAYER M2 ;
        RECT 45.484 7.712 45.556 7.744 ;
  LAYER M2 ;
        RECT 45.52 7.712 45.84 7.744 ;
  LAYER M1 ;
        RECT 45.824 7.692 45.856 7.764 ;
  LAYER M2 ;
        RECT 45.804 7.712 45.876 7.744 ;
  LAYER M1 ;
        RECT 45.504 4.92 45.536 4.992 ;
  LAYER M2 ;
        RECT 45.484 4.94 45.556 4.972 ;
  LAYER M1 ;
        RECT 45.504 4.788 45.536 4.956 ;
  LAYER M1 ;
        RECT 45.504 4.752 45.536 4.824 ;
  LAYER M2 ;
        RECT 45.484 4.772 45.556 4.804 ;
  LAYER M2 ;
        RECT 45.52 4.772 45.84 4.804 ;
  LAYER M1 ;
        RECT 45.824 4.752 45.856 4.824 ;
  LAYER M2 ;
        RECT 45.804 4.772 45.876 4.804 ;
  LAYER M1 ;
        RECT 45.504 1.98 45.536 2.052 ;
  LAYER M2 ;
        RECT 45.484 2 45.556 2.032 ;
  LAYER M1 ;
        RECT 45.504 1.848 45.536 2.016 ;
  LAYER M1 ;
        RECT 45.504 1.812 45.536 1.884 ;
  LAYER M2 ;
        RECT 45.484 1.832 45.556 1.864 ;
  LAYER M2 ;
        RECT 45.52 1.832 45.84 1.864 ;
  LAYER M1 ;
        RECT 45.824 1.812 45.856 1.884 ;
  LAYER M2 ;
        RECT 45.804 1.832 45.876 1.864 ;
  LAYER M1 ;
        RECT 45.824 1.14 45.856 1.212 ;
  LAYER M2 ;
        RECT 45.804 1.16 45.876 1.192 ;
  LAYER M1 ;
        RECT 45.824 1.176 45.856 1.68 ;
  LAYER M1 ;
        RECT 45.824 1.68 45.856 13.608 ;
  LAYER M2 ;
        RECT 31.44 1.16 45.84 1.192 ;
  LAYER M1 ;
        RECT 36.864 13.74 36.896 13.812 ;
  LAYER M2 ;
        RECT 36.844 13.76 36.916 13.792 ;
  LAYER M2 ;
        RECT 34 13.76 36.88 13.792 ;
  LAYER M1 ;
        RECT 33.984 13.74 34.016 13.812 ;
  LAYER M2 ;
        RECT 33.964 13.76 34.036 13.792 ;
  LAYER M1 ;
        RECT 36.864 1.98 36.896 2.052 ;
  LAYER M2 ;
        RECT 36.844 2 36.916 2.032 ;
  LAYER M2 ;
        RECT 34 2 36.88 2.032 ;
  LAYER M1 ;
        RECT 33.984 1.98 34.016 2.052 ;
  LAYER M2 ;
        RECT 33.964 2 34.036 2.032 ;
  LAYER M1 ;
        RECT 39.744 1.98 39.776 2.052 ;
  LAYER M2 ;
        RECT 39.724 2 39.796 2.032 ;
  LAYER M2 ;
        RECT 36.88 2 39.76 2.032 ;
  LAYER M1 ;
        RECT 36.864 1.98 36.896 2.052 ;
  LAYER M2 ;
        RECT 36.844 2 36.916 2.032 ;
  LAYER M1 ;
        RECT 42.624 1.98 42.656 2.052 ;
  LAYER M2 ;
        RECT 42.604 2 42.676 2.032 ;
  LAYER M2 ;
        RECT 39.76 2 42.64 2.032 ;
  LAYER M1 ;
        RECT 39.744 1.98 39.776 2.052 ;
  LAYER M2 ;
        RECT 39.724 2 39.796 2.032 ;
  LAYER M1 ;
        RECT 42.624 13.74 42.656 13.812 ;
  LAYER M2 ;
        RECT 42.604 13.76 42.676 13.792 ;
  LAYER M2 ;
        RECT 42.64 13.76 45.52 13.792 ;
  LAYER M1 ;
        RECT 45.504 13.74 45.536 13.812 ;
  LAYER M2 ;
        RECT 45.484 13.76 45.556 13.792 ;
  LAYER M1 ;
        RECT 39.744 13.74 39.776 13.812 ;
  LAYER M2 ;
        RECT 39.724 13.76 39.796 13.792 ;
  LAYER M2 ;
        RECT 39.76 13.76 42.64 13.792 ;
  LAYER M1 ;
        RECT 42.624 13.74 42.656 13.812 ;
  LAYER M2 ;
        RECT 42.604 13.76 42.676 13.792 ;
  LAYER M1 ;
        RECT 31.584 13.74 31.616 16.248 ;
  LAYER M1 ;
        RECT 31.648 13.74 31.68 16.248 ;
  LAYER M1 ;
        RECT 31.712 13.74 31.744 16.248 ;
  LAYER M1 ;
        RECT 31.776 13.74 31.808 16.248 ;
  LAYER M1 ;
        RECT 31.84 13.74 31.872 16.248 ;
  LAYER M1 ;
        RECT 31.904 13.74 31.936 16.248 ;
  LAYER M1 ;
        RECT 31.968 13.74 32 16.248 ;
  LAYER M1 ;
        RECT 32.032 13.74 32.064 16.248 ;
  LAYER M1 ;
        RECT 32.096 13.74 32.128 16.248 ;
  LAYER M1 ;
        RECT 32.16 13.74 32.192 16.248 ;
  LAYER M1 ;
        RECT 32.224 13.74 32.256 16.248 ;
  LAYER M1 ;
        RECT 32.288 13.74 32.32 16.248 ;
  LAYER M1 ;
        RECT 32.352 13.74 32.384 16.248 ;
  LAYER M1 ;
        RECT 32.416 13.74 32.448 16.248 ;
  LAYER M1 ;
        RECT 32.48 13.74 32.512 16.248 ;
  LAYER M1 ;
        RECT 32.544 13.74 32.576 16.248 ;
  LAYER M1 ;
        RECT 32.608 13.74 32.64 16.248 ;
  LAYER M1 ;
        RECT 32.672 13.74 32.704 16.248 ;
  LAYER M1 ;
        RECT 32.736 13.74 32.768 16.248 ;
  LAYER M1 ;
        RECT 32.8 13.74 32.832 16.248 ;
  LAYER M1 ;
        RECT 32.864 13.74 32.896 16.248 ;
  LAYER M1 ;
        RECT 32.928 13.74 32.96 16.248 ;
  LAYER M1 ;
        RECT 32.992 13.74 33.024 16.248 ;
  LAYER M1 ;
        RECT 33.056 13.74 33.088 16.248 ;
  LAYER M1 ;
        RECT 33.12 13.74 33.152 16.248 ;
  LAYER M1 ;
        RECT 33.184 13.74 33.216 16.248 ;
  LAYER M1 ;
        RECT 33.248 13.74 33.28 16.248 ;
  LAYER M1 ;
        RECT 33.312 13.74 33.344 16.248 ;
  LAYER M1 ;
        RECT 33.376 13.74 33.408 16.248 ;
  LAYER M1 ;
        RECT 33.44 13.74 33.472 16.248 ;
  LAYER M1 ;
        RECT 33.504 13.74 33.536 16.248 ;
  LAYER M1 ;
        RECT 33.568 13.74 33.6 16.248 ;
  LAYER M1 ;
        RECT 33.632 13.74 33.664 16.248 ;
  LAYER M1 ;
        RECT 33.696 13.74 33.728 16.248 ;
  LAYER M1 ;
        RECT 33.76 13.74 33.792 16.248 ;
  LAYER M1 ;
        RECT 33.824 13.74 33.856 16.248 ;
  LAYER M1 ;
        RECT 33.888 13.74 33.92 16.248 ;
  LAYER M2 ;
        RECT 31.564 16.132 34.036 16.164 ;
  LAYER M2 ;
        RECT 31.564 16.068 34.036 16.1 ;
  LAYER M2 ;
        RECT 31.564 16.004 34.036 16.036 ;
  LAYER M2 ;
        RECT 31.564 15.94 34.036 15.972 ;
  LAYER M2 ;
        RECT 31.564 15.876 34.036 15.908 ;
  LAYER M2 ;
        RECT 31.564 15.812 34.036 15.844 ;
  LAYER M2 ;
        RECT 31.564 15.748 34.036 15.78 ;
  LAYER M2 ;
        RECT 31.564 15.684 34.036 15.716 ;
  LAYER M2 ;
        RECT 31.564 15.62 34.036 15.652 ;
  LAYER M2 ;
        RECT 31.564 15.556 34.036 15.588 ;
  LAYER M2 ;
        RECT 31.564 15.492 34.036 15.524 ;
  LAYER M2 ;
        RECT 31.564 15.428 34.036 15.46 ;
  LAYER M2 ;
        RECT 31.564 15.364 34.036 15.396 ;
  LAYER M2 ;
        RECT 31.564 15.3 34.036 15.332 ;
  LAYER M2 ;
        RECT 31.564 15.236 34.036 15.268 ;
  LAYER M2 ;
        RECT 31.564 15.172 34.036 15.204 ;
  LAYER M2 ;
        RECT 31.564 15.108 34.036 15.14 ;
  LAYER M2 ;
        RECT 31.564 15.044 34.036 15.076 ;
  LAYER M2 ;
        RECT 31.564 14.98 34.036 15.012 ;
  LAYER M2 ;
        RECT 31.564 14.916 34.036 14.948 ;
  LAYER M2 ;
        RECT 31.564 14.852 34.036 14.884 ;
  LAYER M2 ;
        RECT 31.564 14.788 34.036 14.82 ;
  LAYER M2 ;
        RECT 31.564 14.724 34.036 14.756 ;
  LAYER M2 ;
        RECT 31.564 14.66 34.036 14.692 ;
  LAYER M2 ;
        RECT 31.564 14.596 34.036 14.628 ;
  LAYER M2 ;
        RECT 31.564 14.532 34.036 14.564 ;
  LAYER M2 ;
        RECT 31.564 14.468 34.036 14.5 ;
  LAYER M2 ;
        RECT 31.564 14.404 34.036 14.436 ;
  LAYER M2 ;
        RECT 31.564 14.34 34.036 14.372 ;
  LAYER M2 ;
        RECT 31.564 14.276 34.036 14.308 ;
  LAYER M2 ;
        RECT 31.564 14.212 34.036 14.244 ;
  LAYER M2 ;
        RECT 31.564 14.148 34.036 14.18 ;
  LAYER M2 ;
        RECT 31.564 14.084 34.036 14.116 ;
  LAYER M2 ;
        RECT 31.564 14.02 34.036 14.052 ;
  LAYER M2 ;
        RECT 31.564 13.956 34.036 13.988 ;
  LAYER M2 ;
        RECT 31.564 13.892 34.036 13.924 ;
  LAYER M3 ;
        RECT 31.584 13.74 31.616 16.248 ;
  LAYER M3 ;
        RECT 31.648 13.74 31.68 16.248 ;
  LAYER M3 ;
        RECT 31.712 13.74 31.744 16.248 ;
  LAYER M3 ;
        RECT 31.776 13.74 31.808 16.248 ;
  LAYER M3 ;
        RECT 31.84 13.74 31.872 16.248 ;
  LAYER M3 ;
        RECT 31.904 13.74 31.936 16.248 ;
  LAYER M3 ;
        RECT 31.968 13.74 32 16.248 ;
  LAYER M3 ;
        RECT 32.032 13.74 32.064 16.248 ;
  LAYER M3 ;
        RECT 32.096 13.74 32.128 16.248 ;
  LAYER M3 ;
        RECT 32.16 13.74 32.192 16.248 ;
  LAYER M3 ;
        RECT 32.224 13.74 32.256 16.248 ;
  LAYER M3 ;
        RECT 32.288 13.74 32.32 16.248 ;
  LAYER M3 ;
        RECT 32.352 13.74 32.384 16.248 ;
  LAYER M3 ;
        RECT 32.416 13.74 32.448 16.248 ;
  LAYER M3 ;
        RECT 32.48 13.74 32.512 16.248 ;
  LAYER M3 ;
        RECT 32.544 13.74 32.576 16.248 ;
  LAYER M3 ;
        RECT 32.608 13.74 32.64 16.248 ;
  LAYER M3 ;
        RECT 32.672 13.74 32.704 16.248 ;
  LAYER M3 ;
        RECT 32.736 13.74 32.768 16.248 ;
  LAYER M3 ;
        RECT 32.8 13.74 32.832 16.248 ;
  LAYER M3 ;
        RECT 32.864 13.74 32.896 16.248 ;
  LAYER M3 ;
        RECT 32.928 13.74 32.96 16.248 ;
  LAYER M3 ;
        RECT 32.992 13.74 33.024 16.248 ;
  LAYER M3 ;
        RECT 33.056 13.74 33.088 16.248 ;
  LAYER M3 ;
        RECT 33.12 13.74 33.152 16.248 ;
  LAYER M3 ;
        RECT 33.184 13.74 33.216 16.248 ;
  LAYER M3 ;
        RECT 33.248 13.74 33.28 16.248 ;
  LAYER M3 ;
        RECT 33.312 13.74 33.344 16.248 ;
  LAYER M3 ;
        RECT 33.376 13.74 33.408 16.248 ;
  LAYER M3 ;
        RECT 33.44 13.74 33.472 16.248 ;
  LAYER M3 ;
        RECT 33.504 13.74 33.536 16.248 ;
  LAYER M3 ;
        RECT 33.568 13.74 33.6 16.248 ;
  LAYER M3 ;
        RECT 33.632 13.74 33.664 16.248 ;
  LAYER M3 ;
        RECT 33.696 13.74 33.728 16.248 ;
  LAYER M3 ;
        RECT 33.76 13.74 33.792 16.248 ;
  LAYER M3 ;
        RECT 33.824 13.74 33.856 16.248 ;
  LAYER M3 ;
        RECT 33.888 13.74 33.92 16.248 ;
  LAYER M3 ;
        RECT 33.984 13.74 34.016 16.248 ;
  LAYER M1 ;
        RECT 31.599 13.776 31.601 16.212 ;
  LAYER M1 ;
        RECT 31.679 13.776 31.681 16.212 ;
  LAYER M1 ;
        RECT 31.759 13.776 31.761 16.212 ;
  LAYER M1 ;
        RECT 31.839 13.776 31.841 16.212 ;
  LAYER M1 ;
        RECT 31.919 13.776 31.921 16.212 ;
  LAYER M1 ;
        RECT 31.999 13.776 32.001 16.212 ;
  LAYER M1 ;
        RECT 32.079 13.776 32.081 16.212 ;
  LAYER M1 ;
        RECT 32.159 13.776 32.161 16.212 ;
  LAYER M1 ;
        RECT 32.239 13.776 32.241 16.212 ;
  LAYER M1 ;
        RECT 32.319 13.776 32.321 16.212 ;
  LAYER M1 ;
        RECT 32.399 13.776 32.401 16.212 ;
  LAYER M1 ;
        RECT 32.479 13.776 32.481 16.212 ;
  LAYER M1 ;
        RECT 32.559 13.776 32.561 16.212 ;
  LAYER M1 ;
        RECT 32.639 13.776 32.641 16.212 ;
  LAYER M1 ;
        RECT 32.719 13.776 32.721 16.212 ;
  LAYER M1 ;
        RECT 32.799 13.776 32.801 16.212 ;
  LAYER M1 ;
        RECT 32.879 13.776 32.881 16.212 ;
  LAYER M1 ;
        RECT 32.959 13.776 32.961 16.212 ;
  LAYER M1 ;
        RECT 33.039 13.776 33.041 16.212 ;
  LAYER M1 ;
        RECT 33.119 13.776 33.121 16.212 ;
  LAYER M1 ;
        RECT 33.199 13.776 33.201 16.212 ;
  LAYER M1 ;
        RECT 33.279 13.776 33.281 16.212 ;
  LAYER M1 ;
        RECT 33.359 13.776 33.361 16.212 ;
  LAYER M1 ;
        RECT 33.439 13.776 33.441 16.212 ;
  LAYER M1 ;
        RECT 33.519 13.776 33.521 16.212 ;
  LAYER M1 ;
        RECT 33.599 13.776 33.601 16.212 ;
  LAYER M1 ;
        RECT 33.679 13.776 33.681 16.212 ;
  LAYER M1 ;
        RECT 33.759 13.776 33.761 16.212 ;
  LAYER M1 ;
        RECT 33.839 13.776 33.841 16.212 ;
  LAYER M1 ;
        RECT 33.919 13.776 33.921 16.212 ;
  LAYER M2 ;
        RECT 31.6 16.211 34 16.213 ;
  LAYER M2 ;
        RECT 31.6 16.127 34 16.129 ;
  LAYER M2 ;
        RECT 31.6 16.043 34 16.045 ;
  LAYER M2 ;
        RECT 31.6 15.959 34 15.961 ;
  LAYER M2 ;
        RECT 31.6 15.875 34 15.877 ;
  LAYER M2 ;
        RECT 31.6 15.791 34 15.793 ;
  LAYER M2 ;
        RECT 31.6 15.707 34 15.709 ;
  LAYER M2 ;
        RECT 31.6 15.623 34 15.625 ;
  LAYER M2 ;
        RECT 31.6 15.539 34 15.541 ;
  LAYER M2 ;
        RECT 31.6 15.455 34 15.457 ;
  LAYER M2 ;
        RECT 31.6 15.371 34 15.373 ;
  LAYER M2 ;
        RECT 31.6 15.287 34 15.289 ;
  LAYER M2 ;
        RECT 31.6 15.2035 34 15.2055 ;
  LAYER M2 ;
        RECT 31.6 15.119 34 15.121 ;
  LAYER M2 ;
        RECT 31.6 15.035 34 15.037 ;
  LAYER M2 ;
        RECT 31.6 14.951 34 14.953 ;
  LAYER M2 ;
        RECT 31.6 14.867 34 14.869 ;
  LAYER M2 ;
        RECT 31.6 14.783 34 14.785 ;
  LAYER M2 ;
        RECT 31.6 14.699 34 14.701 ;
  LAYER M2 ;
        RECT 31.6 14.615 34 14.617 ;
  LAYER M2 ;
        RECT 31.6 14.531 34 14.533 ;
  LAYER M2 ;
        RECT 31.6 14.447 34 14.449 ;
  LAYER M2 ;
        RECT 31.6 14.363 34 14.365 ;
  LAYER M2 ;
        RECT 31.6 14.279 34 14.281 ;
  LAYER M2 ;
        RECT 31.6 14.195 34 14.197 ;
  LAYER M2 ;
        RECT 31.6 14.111 34 14.113 ;
  LAYER M2 ;
        RECT 31.6 14.027 34 14.029 ;
  LAYER M2 ;
        RECT 31.6 13.943 34 13.945 ;
  LAYER M2 ;
        RECT 31.6 13.859 34 13.861 ;
  LAYER M1 ;
        RECT 31.584 10.8 31.616 13.308 ;
  LAYER M1 ;
        RECT 31.648 10.8 31.68 13.308 ;
  LAYER M1 ;
        RECT 31.712 10.8 31.744 13.308 ;
  LAYER M1 ;
        RECT 31.776 10.8 31.808 13.308 ;
  LAYER M1 ;
        RECT 31.84 10.8 31.872 13.308 ;
  LAYER M1 ;
        RECT 31.904 10.8 31.936 13.308 ;
  LAYER M1 ;
        RECT 31.968 10.8 32 13.308 ;
  LAYER M1 ;
        RECT 32.032 10.8 32.064 13.308 ;
  LAYER M1 ;
        RECT 32.096 10.8 32.128 13.308 ;
  LAYER M1 ;
        RECT 32.16 10.8 32.192 13.308 ;
  LAYER M1 ;
        RECT 32.224 10.8 32.256 13.308 ;
  LAYER M1 ;
        RECT 32.288 10.8 32.32 13.308 ;
  LAYER M1 ;
        RECT 32.352 10.8 32.384 13.308 ;
  LAYER M1 ;
        RECT 32.416 10.8 32.448 13.308 ;
  LAYER M1 ;
        RECT 32.48 10.8 32.512 13.308 ;
  LAYER M1 ;
        RECT 32.544 10.8 32.576 13.308 ;
  LAYER M1 ;
        RECT 32.608 10.8 32.64 13.308 ;
  LAYER M1 ;
        RECT 32.672 10.8 32.704 13.308 ;
  LAYER M1 ;
        RECT 32.736 10.8 32.768 13.308 ;
  LAYER M1 ;
        RECT 32.8 10.8 32.832 13.308 ;
  LAYER M1 ;
        RECT 32.864 10.8 32.896 13.308 ;
  LAYER M1 ;
        RECT 32.928 10.8 32.96 13.308 ;
  LAYER M1 ;
        RECT 32.992 10.8 33.024 13.308 ;
  LAYER M1 ;
        RECT 33.056 10.8 33.088 13.308 ;
  LAYER M1 ;
        RECT 33.12 10.8 33.152 13.308 ;
  LAYER M1 ;
        RECT 33.184 10.8 33.216 13.308 ;
  LAYER M1 ;
        RECT 33.248 10.8 33.28 13.308 ;
  LAYER M1 ;
        RECT 33.312 10.8 33.344 13.308 ;
  LAYER M1 ;
        RECT 33.376 10.8 33.408 13.308 ;
  LAYER M1 ;
        RECT 33.44 10.8 33.472 13.308 ;
  LAYER M1 ;
        RECT 33.504 10.8 33.536 13.308 ;
  LAYER M1 ;
        RECT 33.568 10.8 33.6 13.308 ;
  LAYER M1 ;
        RECT 33.632 10.8 33.664 13.308 ;
  LAYER M1 ;
        RECT 33.696 10.8 33.728 13.308 ;
  LAYER M1 ;
        RECT 33.76 10.8 33.792 13.308 ;
  LAYER M1 ;
        RECT 33.824 10.8 33.856 13.308 ;
  LAYER M1 ;
        RECT 33.888 10.8 33.92 13.308 ;
  LAYER M2 ;
        RECT 31.564 13.192 34.036 13.224 ;
  LAYER M2 ;
        RECT 31.564 13.128 34.036 13.16 ;
  LAYER M2 ;
        RECT 31.564 13.064 34.036 13.096 ;
  LAYER M2 ;
        RECT 31.564 13 34.036 13.032 ;
  LAYER M2 ;
        RECT 31.564 12.936 34.036 12.968 ;
  LAYER M2 ;
        RECT 31.564 12.872 34.036 12.904 ;
  LAYER M2 ;
        RECT 31.564 12.808 34.036 12.84 ;
  LAYER M2 ;
        RECT 31.564 12.744 34.036 12.776 ;
  LAYER M2 ;
        RECT 31.564 12.68 34.036 12.712 ;
  LAYER M2 ;
        RECT 31.564 12.616 34.036 12.648 ;
  LAYER M2 ;
        RECT 31.564 12.552 34.036 12.584 ;
  LAYER M2 ;
        RECT 31.564 12.488 34.036 12.52 ;
  LAYER M2 ;
        RECT 31.564 12.424 34.036 12.456 ;
  LAYER M2 ;
        RECT 31.564 12.36 34.036 12.392 ;
  LAYER M2 ;
        RECT 31.564 12.296 34.036 12.328 ;
  LAYER M2 ;
        RECT 31.564 12.232 34.036 12.264 ;
  LAYER M2 ;
        RECT 31.564 12.168 34.036 12.2 ;
  LAYER M2 ;
        RECT 31.564 12.104 34.036 12.136 ;
  LAYER M2 ;
        RECT 31.564 12.04 34.036 12.072 ;
  LAYER M2 ;
        RECT 31.564 11.976 34.036 12.008 ;
  LAYER M2 ;
        RECT 31.564 11.912 34.036 11.944 ;
  LAYER M2 ;
        RECT 31.564 11.848 34.036 11.88 ;
  LAYER M2 ;
        RECT 31.564 11.784 34.036 11.816 ;
  LAYER M2 ;
        RECT 31.564 11.72 34.036 11.752 ;
  LAYER M2 ;
        RECT 31.564 11.656 34.036 11.688 ;
  LAYER M2 ;
        RECT 31.564 11.592 34.036 11.624 ;
  LAYER M2 ;
        RECT 31.564 11.528 34.036 11.56 ;
  LAYER M2 ;
        RECT 31.564 11.464 34.036 11.496 ;
  LAYER M2 ;
        RECT 31.564 11.4 34.036 11.432 ;
  LAYER M2 ;
        RECT 31.564 11.336 34.036 11.368 ;
  LAYER M2 ;
        RECT 31.564 11.272 34.036 11.304 ;
  LAYER M2 ;
        RECT 31.564 11.208 34.036 11.24 ;
  LAYER M2 ;
        RECT 31.564 11.144 34.036 11.176 ;
  LAYER M2 ;
        RECT 31.564 11.08 34.036 11.112 ;
  LAYER M2 ;
        RECT 31.564 11.016 34.036 11.048 ;
  LAYER M2 ;
        RECT 31.564 10.952 34.036 10.984 ;
  LAYER M3 ;
        RECT 31.584 10.8 31.616 13.308 ;
  LAYER M3 ;
        RECT 31.648 10.8 31.68 13.308 ;
  LAYER M3 ;
        RECT 31.712 10.8 31.744 13.308 ;
  LAYER M3 ;
        RECT 31.776 10.8 31.808 13.308 ;
  LAYER M3 ;
        RECT 31.84 10.8 31.872 13.308 ;
  LAYER M3 ;
        RECT 31.904 10.8 31.936 13.308 ;
  LAYER M3 ;
        RECT 31.968 10.8 32 13.308 ;
  LAYER M3 ;
        RECT 32.032 10.8 32.064 13.308 ;
  LAYER M3 ;
        RECT 32.096 10.8 32.128 13.308 ;
  LAYER M3 ;
        RECT 32.16 10.8 32.192 13.308 ;
  LAYER M3 ;
        RECT 32.224 10.8 32.256 13.308 ;
  LAYER M3 ;
        RECT 32.288 10.8 32.32 13.308 ;
  LAYER M3 ;
        RECT 32.352 10.8 32.384 13.308 ;
  LAYER M3 ;
        RECT 32.416 10.8 32.448 13.308 ;
  LAYER M3 ;
        RECT 32.48 10.8 32.512 13.308 ;
  LAYER M3 ;
        RECT 32.544 10.8 32.576 13.308 ;
  LAYER M3 ;
        RECT 32.608 10.8 32.64 13.308 ;
  LAYER M3 ;
        RECT 32.672 10.8 32.704 13.308 ;
  LAYER M3 ;
        RECT 32.736 10.8 32.768 13.308 ;
  LAYER M3 ;
        RECT 32.8 10.8 32.832 13.308 ;
  LAYER M3 ;
        RECT 32.864 10.8 32.896 13.308 ;
  LAYER M3 ;
        RECT 32.928 10.8 32.96 13.308 ;
  LAYER M3 ;
        RECT 32.992 10.8 33.024 13.308 ;
  LAYER M3 ;
        RECT 33.056 10.8 33.088 13.308 ;
  LAYER M3 ;
        RECT 33.12 10.8 33.152 13.308 ;
  LAYER M3 ;
        RECT 33.184 10.8 33.216 13.308 ;
  LAYER M3 ;
        RECT 33.248 10.8 33.28 13.308 ;
  LAYER M3 ;
        RECT 33.312 10.8 33.344 13.308 ;
  LAYER M3 ;
        RECT 33.376 10.8 33.408 13.308 ;
  LAYER M3 ;
        RECT 33.44 10.8 33.472 13.308 ;
  LAYER M3 ;
        RECT 33.504 10.8 33.536 13.308 ;
  LAYER M3 ;
        RECT 33.568 10.8 33.6 13.308 ;
  LAYER M3 ;
        RECT 33.632 10.8 33.664 13.308 ;
  LAYER M3 ;
        RECT 33.696 10.8 33.728 13.308 ;
  LAYER M3 ;
        RECT 33.76 10.8 33.792 13.308 ;
  LAYER M3 ;
        RECT 33.824 10.8 33.856 13.308 ;
  LAYER M3 ;
        RECT 33.888 10.8 33.92 13.308 ;
  LAYER M3 ;
        RECT 33.984 10.8 34.016 13.308 ;
  LAYER M1 ;
        RECT 31.599 10.836 31.601 13.272 ;
  LAYER M1 ;
        RECT 31.679 10.836 31.681 13.272 ;
  LAYER M1 ;
        RECT 31.759 10.836 31.761 13.272 ;
  LAYER M1 ;
        RECT 31.839 10.836 31.841 13.272 ;
  LAYER M1 ;
        RECT 31.919 10.836 31.921 13.272 ;
  LAYER M1 ;
        RECT 31.999 10.836 32.001 13.272 ;
  LAYER M1 ;
        RECT 32.079 10.836 32.081 13.272 ;
  LAYER M1 ;
        RECT 32.159 10.836 32.161 13.272 ;
  LAYER M1 ;
        RECT 32.239 10.836 32.241 13.272 ;
  LAYER M1 ;
        RECT 32.319 10.836 32.321 13.272 ;
  LAYER M1 ;
        RECT 32.399 10.836 32.401 13.272 ;
  LAYER M1 ;
        RECT 32.479 10.836 32.481 13.272 ;
  LAYER M1 ;
        RECT 32.559 10.836 32.561 13.272 ;
  LAYER M1 ;
        RECT 32.639 10.836 32.641 13.272 ;
  LAYER M1 ;
        RECT 32.719 10.836 32.721 13.272 ;
  LAYER M1 ;
        RECT 32.799 10.836 32.801 13.272 ;
  LAYER M1 ;
        RECT 32.879 10.836 32.881 13.272 ;
  LAYER M1 ;
        RECT 32.959 10.836 32.961 13.272 ;
  LAYER M1 ;
        RECT 33.039 10.836 33.041 13.272 ;
  LAYER M1 ;
        RECT 33.119 10.836 33.121 13.272 ;
  LAYER M1 ;
        RECT 33.199 10.836 33.201 13.272 ;
  LAYER M1 ;
        RECT 33.279 10.836 33.281 13.272 ;
  LAYER M1 ;
        RECT 33.359 10.836 33.361 13.272 ;
  LAYER M1 ;
        RECT 33.439 10.836 33.441 13.272 ;
  LAYER M1 ;
        RECT 33.519 10.836 33.521 13.272 ;
  LAYER M1 ;
        RECT 33.599 10.836 33.601 13.272 ;
  LAYER M1 ;
        RECT 33.679 10.836 33.681 13.272 ;
  LAYER M1 ;
        RECT 33.759 10.836 33.761 13.272 ;
  LAYER M1 ;
        RECT 33.839 10.836 33.841 13.272 ;
  LAYER M1 ;
        RECT 33.919 10.836 33.921 13.272 ;
  LAYER M2 ;
        RECT 31.6 13.271 34 13.273 ;
  LAYER M2 ;
        RECT 31.6 13.187 34 13.189 ;
  LAYER M2 ;
        RECT 31.6 13.103 34 13.105 ;
  LAYER M2 ;
        RECT 31.6 13.019 34 13.021 ;
  LAYER M2 ;
        RECT 31.6 12.935 34 12.937 ;
  LAYER M2 ;
        RECT 31.6 12.851 34 12.853 ;
  LAYER M2 ;
        RECT 31.6 12.767 34 12.769 ;
  LAYER M2 ;
        RECT 31.6 12.683 34 12.685 ;
  LAYER M2 ;
        RECT 31.6 12.599 34 12.601 ;
  LAYER M2 ;
        RECT 31.6 12.515 34 12.517 ;
  LAYER M2 ;
        RECT 31.6 12.431 34 12.433 ;
  LAYER M2 ;
        RECT 31.6 12.347 34 12.349 ;
  LAYER M2 ;
        RECT 31.6 12.2635 34 12.2655 ;
  LAYER M2 ;
        RECT 31.6 12.179 34 12.181 ;
  LAYER M2 ;
        RECT 31.6 12.095 34 12.097 ;
  LAYER M2 ;
        RECT 31.6 12.011 34 12.013 ;
  LAYER M2 ;
        RECT 31.6 11.927 34 11.929 ;
  LAYER M2 ;
        RECT 31.6 11.843 34 11.845 ;
  LAYER M2 ;
        RECT 31.6 11.759 34 11.761 ;
  LAYER M2 ;
        RECT 31.6 11.675 34 11.677 ;
  LAYER M2 ;
        RECT 31.6 11.591 34 11.593 ;
  LAYER M2 ;
        RECT 31.6 11.507 34 11.509 ;
  LAYER M2 ;
        RECT 31.6 11.423 34 11.425 ;
  LAYER M2 ;
        RECT 31.6 11.339 34 11.341 ;
  LAYER M2 ;
        RECT 31.6 11.255 34 11.257 ;
  LAYER M2 ;
        RECT 31.6 11.171 34 11.173 ;
  LAYER M2 ;
        RECT 31.6 11.087 34 11.089 ;
  LAYER M2 ;
        RECT 31.6 11.003 34 11.005 ;
  LAYER M2 ;
        RECT 31.6 10.919 34 10.921 ;
  LAYER M1 ;
        RECT 31.584 7.86 31.616 10.368 ;
  LAYER M1 ;
        RECT 31.648 7.86 31.68 10.368 ;
  LAYER M1 ;
        RECT 31.712 7.86 31.744 10.368 ;
  LAYER M1 ;
        RECT 31.776 7.86 31.808 10.368 ;
  LAYER M1 ;
        RECT 31.84 7.86 31.872 10.368 ;
  LAYER M1 ;
        RECT 31.904 7.86 31.936 10.368 ;
  LAYER M1 ;
        RECT 31.968 7.86 32 10.368 ;
  LAYER M1 ;
        RECT 32.032 7.86 32.064 10.368 ;
  LAYER M1 ;
        RECT 32.096 7.86 32.128 10.368 ;
  LAYER M1 ;
        RECT 32.16 7.86 32.192 10.368 ;
  LAYER M1 ;
        RECT 32.224 7.86 32.256 10.368 ;
  LAYER M1 ;
        RECT 32.288 7.86 32.32 10.368 ;
  LAYER M1 ;
        RECT 32.352 7.86 32.384 10.368 ;
  LAYER M1 ;
        RECT 32.416 7.86 32.448 10.368 ;
  LAYER M1 ;
        RECT 32.48 7.86 32.512 10.368 ;
  LAYER M1 ;
        RECT 32.544 7.86 32.576 10.368 ;
  LAYER M1 ;
        RECT 32.608 7.86 32.64 10.368 ;
  LAYER M1 ;
        RECT 32.672 7.86 32.704 10.368 ;
  LAYER M1 ;
        RECT 32.736 7.86 32.768 10.368 ;
  LAYER M1 ;
        RECT 32.8 7.86 32.832 10.368 ;
  LAYER M1 ;
        RECT 32.864 7.86 32.896 10.368 ;
  LAYER M1 ;
        RECT 32.928 7.86 32.96 10.368 ;
  LAYER M1 ;
        RECT 32.992 7.86 33.024 10.368 ;
  LAYER M1 ;
        RECT 33.056 7.86 33.088 10.368 ;
  LAYER M1 ;
        RECT 33.12 7.86 33.152 10.368 ;
  LAYER M1 ;
        RECT 33.184 7.86 33.216 10.368 ;
  LAYER M1 ;
        RECT 33.248 7.86 33.28 10.368 ;
  LAYER M1 ;
        RECT 33.312 7.86 33.344 10.368 ;
  LAYER M1 ;
        RECT 33.376 7.86 33.408 10.368 ;
  LAYER M1 ;
        RECT 33.44 7.86 33.472 10.368 ;
  LAYER M1 ;
        RECT 33.504 7.86 33.536 10.368 ;
  LAYER M1 ;
        RECT 33.568 7.86 33.6 10.368 ;
  LAYER M1 ;
        RECT 33.632 7.86 33.664 10.368 ;
  LAYER M1 ;
        RECT 33.696 7.86 33.728 10.368 ;
  LAYER M1 ;
        RECT 33.76 7.86 33.792 10.368 ;
  LAYER M1 ;
        RECT 33.824 7.86 33.856 10.368 ;
  LAYER M1 ;
        RECT 33.888 7.86 33.92 10.368 ;
  LAYER M2 ;
        RECT 31.564 10.252 34.036 10.284 ;
  LAYER M2 ;
        RECT 31.564 10.188 34.036 10.22 ;
  LAYER M2 ;
        RECT 31.564 10.124 34.036 10.156 ;
  LAYER M2 ;
        RECT 31.564 10.06 34.036 10.092 ;
  LAYER M2 ;
        RECT 31.564 9.996 34.036 10.028 ;
  LAYER M2 ;
        RECT 31.564 9.932 34.036 9.964 ;
  LAYER M2 ;
        RECT 31.564 9.868 34.036 9.9 ;
  LAYER M2 ;
        RECT 31.564 9.804 34.036 9.836 ;
  LAYER M2 ;
        RECT 31.564 9.74 34.036 9.772 ;
  LAYER M2 ;
        RECT 31.564 9.676 34.036 9.708 ;
  LAYER M2 ;
        RECT 31.564 9.612 34.036 9.644 ;
  LAYER M2 ;
        RECT 31.564 9.548 34.036 9.58 ;
  LAYER M2 ;
        RECT 31.564 9.484 34.036 9.516 ;
  LAYER M2 ;
        RECT 31.564 9.42 34.036 9.452 ;
  LAYER M2 ;
        RECT 31.564 9.356 34.036 9.388 ;
  LAYER M2 ;
        RECT 31.564 9.292 34.036 9.324 ;
  LAYER M2 ;
        RECT 31.564 9.228 34.036 9.26 ;
  LAYER M2 ;
        RECT 31.564 9.164 34.036 9.196 ;
  LAYER M2 ;
        RECT 31.564 9.1 34.036 9.132 ;
  LAYER M2 ;
        RECT 31.564 9.036 34.036 9.068 ;
  LAYER M2 ;
        RECT 31.564 8.972 34.036 9.004 ;
  LAYER M2 ;
        RECT 31.564 8.908 34.036 8.94 ;
  LAYER M2 ;
        RECT 31.564 8.844 34.036 8.876 ;
  LAYER M2 ;
        RECT 31.564 8.78 34.036 8.812 ;
  LAYER M2 ;
        RECT 31.564 8.716 34.036 8.748 ;
  LAYER M2 ;
        RECT 31.564 8.652 34.036 8.684 ;
  LAYER M2 ;
        RECT 31.564 8.588 34.036 8.62 ;
  LAYER M2 ;
        RECT 31.564 8.524 34.036 8.556 ;
  LAYER M2 ;
        RECT 31.564 8.46 34.036 8.492 ;
  LAYER M2 ;
        RECT 31.564 8.396 34.036 8.428 ;
  LAYER M2 ;
        RECT 31.564 8.332 34.036 8.364 ;
  LAYER M2 ;
        RECT 31.564 8.268 34.036 8.3 ;
  LAYER M2 ;
        RECT 31.564 8.204 34.036 8.236 ;
  LAYER M2 ;
        RECT 31.564 8.14 34.036 8.172 ;
  LAYER M2 ;
        RECT 31.564 8.076 34.036 8.108 ;
  LAYER M2 ;
        RECT 31.564 8.012 34.036 8.044 ;
  LAYER M3 ;
        RECT 31.584 7.86 31.616 10.368 ;
  LAYER M3 ;
        RECT 31.648 7.86 31.68 10.368 ;
  LAYER M3 ;
        RECT 31.712 7.86 31.744 10.368 ;
  LAYER M3 ;
        RECT 31.776 7.86 31.808 10.368 ;
  LAYER M3 ;
        RECT 31.84 7.86 31.872 10.368 ;
  LAYER M3 ;
        RECT 31.904 7.86 31.936 10.368 ;
  LAYER M3 ;
        RECT 31.968 7.86 32 10.368 ;
  LAYER M3 ;
        RECT 32.032 7.86 32.064 10.368 ;
  LAYER M3 ;
        RECT 32.096 7.86 32.128 10.368 ;
  LAYER M3 ;
        RECT 32.16 7.86 32.192 10.368 ;
  LAYER M3 ;
        RECT 32.224 7.86 32.256 10.368 ;
  LAYER M3 ;
        RECT 32.288 7.86 32.32 10.368 ;
  LAYER M3 ;
        RECT 32.352 7.86 32.384 10.368 ;
  LAYER M3 ;
        RECT 32.416 7.86 32.448 10.368 ;
  LAYER M3 ;
        RECT 32.48 7.86 32.512 10.368 ;
  LAYER M3 ;
        RECT 32.544 7.86 32.576 10.368 ;
  LAYER M3 ;
        RECT 32.608 7.86 32.64 10.368 ;
  LAYER M3 ;
        RECT 32.672 7.86 32.704 10.368 ;
  LAYER M3 ;
        RECT 32.736 7.86 32.768 10.368 ;
  LAYER M3 ;
        RECT 32.8 7.86 32.832 10.368 ;
  LAYER M3 ;
        RECT 32.864 7.86 32.896 10.368 ;
  LAYER M3 ;
        RECT 32.928 7.86 32.96 10.368 ;
  LAYER M3 ;
        RECT 32.992 7.86 33.024 10.368 ;
  LAYER M3 ;
        RECT 33.056 7.86 33.088 10.368 ;
  LAYER M3 ;
        RECT 33.12 7.86 33.152 10.368 ;
  LAYER M3 ;
        RECT 33.184 7.86 33.216 10.368 ;
  LAYER M3 ;
        RECT 33.248 7.86 33.28 10.368 ;
  LAYER M3 ;
        RECT 33.312 7.86 33.344 10.368 ;
  LAYER M3 ;
        RECT 33.376 7.86 33.408 10.368 ;
  LAYER M3 ;
        RECT 33.44 7.86 33.472 10.368 ;
  LAYER M3 ;
        RECT 33.504 7.86 33.536 10.368 ;
  LAYER M3 ;
        RECT 33.568 7.86 33.6 10.368 ;
  LAYER M3 ;
        RECT 33.632 7.86 33.664 10.368 ;
  LAYER M3 ;
        RECT 33.696 7.86 33.728 10.368 ;
  LAYER M3 ;
        RECT 33.76 7.86 33.792 10.368 ;
  LAYER M3 ;
        RECT 33.824 7.86 33.856 10.368 ;
  LAYER M3 ;
        RECT 33.888 7.86 33.92 10.368 ;
  LAYER M3 ;
        RECT 33.984 7.86 34.016 10.368 ;
  LAYER M1 ;
        RECT 31.599 7.896 31.601 10.332 ;
  LAYER M1 ;
        RECT 31.679 7.896 31.681 10.332 ;
  LAYER M1 ;
        RECT 31.759 7.896 31.761 10.332 ;
  LAYER M1 ;
        RECT 31.839 7.896 31.841 10.332 ;
  LAYER M1 ;
        RECT 31.919 7.896 31.921 10.332 ;
  LAYER M1 ;
        RECT 31.999 7.896 32.001 10.332 ;
  LAYER M1 ;
        RECT 32.079 7.896 32.081 10.332 ;
  LAYER M1 ;
        RECT 32.159 7.896 32.161 10.332 ;
  LAYER M1 ;
        RECT 32.239 7.896 32.241 10.332 ;
  LAYER M1 ;
        RECT 32.319 7.896 32.321 10.332 ;
  LAYER M1 ;
        RECT 32.399 7.896 32.401 10.332 ;
  LAYER M1 ;
        RECT 32.479 7.896 32.481 10.332 ;
  LAYER M1 ;
        RECT 32.559 7.896 32.561 10.332 ;
  LAYER M1 ;
        RECT 32.639 7.896 32.641 10.332 ;
  LAYER M1 ;
        RECT 32.719 7.896 32.721 10.332 ;
  LAYER M1 ;
        RECT 32.799 7.896 32.801 10.332 ;
  LAYER M1 ;
        RECT 32.879 7.896 32.881 10.332 ;
  LAYER M1 ;
        RECT 32.959 7.896 32.961 10.332 ;
  LAYER M1 ;
        RECT 33.039 7.896 33.041 10.332 ;
  LAYER M1 ;
        RECT 33.119 7.896 33.121 10.332 ;
  LAYER M1 ;
        RECT 33.199 7.896 33.201 10.332 ;
  LAYER M1 ;
        RECT 33.279 7.896 33.281 10.332 ;
  LAYER M1 ;
        RECT 33.359 7.896 33.361 10.332 ;
  LAYER M1 ;
        RECT 33.439 7.896 33.441 10.332 ;
  LAYER M1 ;
        RECT 33.519 7.896 33.521 10.332 ;
  LAYER M1 ;
        RECT 33.599 7.896 33.601 10.332 ;
  LAYER M1 ;
        RECT 33.679 7.896 33.681 10.332 ;
  LAYER M1 ;
        RECT 33.759 7.896 33.761 10.332 ;
  LAYER M1 ;
        RECT 33.839 7.896 33.841 10.332 ;
  LAYER M1 ;
        RECT 33.919 7.896 33.921 10.332 ;
  LAYER M2 ;
        RECT 31.6 10.331 34 10.333 ;
  LAYER M2 ;
        RECT 31.6 10.247 34 10.249 ;
  LAYER M2 ;
        RECT 31.6 10.163 34 10.165 ;
  LAYER M2 ;
        RECT 31.6 10.079 34 10.081 ;
  LAYER M2 ;
        RECT 31.6 9.995 34 9.997 ;
  LAYER M2 ;
        RECT 31.6 9.911 34 9.913 ;
  LAYER M2 ;
        RECT 31.6 9.827 34 9.829 ;
  LAYER M2 ;
        RECT 31.6 9.743 34 9.745 ;
  LAYER M2 ;
        RECT 31.6 9.659 34 9.661 ;
  LAYER M2 ;
        RECT 31.6 9.575 34 9.577 ;
  LAYER M2 ;
        RECT 31.6 9.491 34 9.493 ;
  LAYER M2 ;
        RECT 31.6 9.407 34 9.409 ;
  LAYER M2 ;
        RECT 31.6 9.3235 34 9.3255 ;
  LAYER M2 ;
        RECT 31.6 9.239 34 9.241 ;
  LAYER M2 ;
        RECT 31.6 9.155 34 9.157 ;
  LAYER M2 ;
        RECT 31.6 9.071 34 9.073 ;
  LAYER M2 ;
        RECT 31.6 8.987 34 8.989 ;
  LAYER M2 ;
        RECT 31.6 8.903 34 8.905 ;
  LAYER M2 ;
        RECT 31.6 8.819 34 8.821 ;
  LAYER M2 ;
        RECT 31.6 8.735 34 8.737 ;
  LAYER M2 ;
        RECT 31.6 8.651 34 8.653 ;
  LAYER M2 ;
        RECT 31.6 8.567 34 8.569 ;
  LAYER M2 ;
        RECT 31.6 8.483 34 8.485 ;
  LAYER M2 ;
        RECT 31.6 8.399 34 8.401 ;
  LAYER M2 ;
        RECT 31.6 8.315 34 8.317 ;
  LAYER M2 ;
        RECT 31.6 8.231 34 8.233 ;
  LAYER M2 ;
        RECT 31.6 8.147 34 8.149 ;
  LAYER M2 ;
        RECT 31.6 8.063 34 8.065 ;
  LAYER M2 ;
        RECT 31.6 7.979 34 7.981 ;
  LAYER M1 ;
        RECT 31.584 4.92 31.616 7.428 ;
  LAYER M1 ;
        RECT 31.648 4.92 31.68 7.428 ;
  LAYER M1 ;
        RECT 31.712 4.92 31.744 7.428 ;
  LAYER M1 ;
        RECT 31.776 4.92 31.808 7.428 ;
  LAYER M1 ;
        RECT 31.84 4.92 31.872 7.428 ;
  LAYER M1 ;
        RECT 31.904 4.92 31.936 7.428 ;
  LAYER M1 ;
        RECT 31.968 4.92 32 7.428 ;
  LAYER M1 ;
        RECT 32.032 4.92 32.064 7.428 ;
  LAYER M1 ;
        RECT 32.096 4.92 32.128 7.428 ;
  LAYER M1 ;
        RECT 32.16 4.92 32.192 7.428 ;
  LAYER M1 ;
        RECT 32.224 4.92 32.256 7.428 ;
  LAYER M1 ;
        RECT 32.288 4.92 32.32 7.428 ;
  LAYER M1 ;
        RECT 32.352 4.92 32.384 7.428 ;
  LAYER M1 ;
        RECT 32.416 4.92 32.448 7.428 ;
  LAYER M1 ;
        RECT 32.48 4.92 32.512 7.428 ;
  LAYER M1 ;
        RECT 32.544 4.92 32.576 7.428 ;
  LAYER M1 ;
        RECT 32.608 4.92 32.64 7.428 ;
  LAYER M1 ;
        RECT 32.672 4.92 32.704 7.428 ;
  LAYER M1 ;
        RECT 32.736 4.92 32.768 7.428 ;
  LAYER M1 ;
        RECT 32.8 4.92 32.832 7.428 ;
  LAYER M1 ;
        RECT 32.864 4.92 32.896 7.428 ;
  LAYER M1 ;
        RECT 32.928 4.92 32.96 7.428 ;
  LAYER M1 ;
        RECT 32.992 4.92 33.024 7.428 ;
  LAYER M1 ;
        RECT 33.056 4.92 33.088 7.428 ;
  LAYER M1 ;
        RECT 33.12 4.92 33.152 7.428 ;
  LAYER M1 ;
        RECT 33.184 4.92 33.216 7.428 ;
  LAYER M1 ;
        RECT 33.248 4.92 33.28 7.428 ;
  LAYER M1 ;
        RECT 33.312 4.92 33.344 7.428 ;
  LAYER M1 ;
        RECT 33.376 4.92 33.408 7.428 ;
  LAYER M1 ;
        RECT 33.44 4.92 33.472 7.428 ;
  LAYER M1 ;
        RECT 33.504 4.92 33.536 7.428 ;
  LAYER M1 ;
        RECT 33.568 4.92 33.6 7.428 ;
  LAYER M1 ;
        RECT 33.632 4.92 33.664 7.428 ;
  LAYER M1 ;
        RECT 33.696 4.92 33.728 7.428 ;
  LAYER M1 ;
        RECT 33.76 4.92 33.792 7.428 ;
  LAYER M1 ;
        RECT 33.824 4.92 33.856 7.428 ;
  LAYER M1 ;
        RECT 33.888 4.92 33.92 7.428 ;
  LAYER M2 ;
        RECT 31.564 7.312 34.036 7.344 ;
  LAYER M2 ;
        RECT 31.564 7.248 34.036 7.28 ;
  LAYER M2 ;
        RECT 31.564 7.184 34.036 7.216 ;
  LAYER M2 ;
        RECT 31.564 7.12 34.036 7.152 ;
  LAYER M2 ;
        RECT 31.564 7.056 34.036 7.088 ;
  LAYER M2 ;
        RECT 31.564 6.992 34.036 7.024 ;
  LAYER M2 ;
        RECT 31.564 6.928 34.036 6.96 ;
  LAYER M2 ;
        RECT 31.564 6.864 34.036 6.896 ;
  LAYER M2 ;
        RECT 31.564 6.8 34.036 6.832 ;
  LAYER M2 ;
        RECT 31.564 6.736 34.036 6.768 ;
  LAYER M2 ;
        RECT 31.564 6.672 34.036 6.704 ;
  LAYER M2 ;
        RECT 31.564 6.608 34.036 6.64 ;
  LAYER M2 ;
        RECT 31.564 6.544 34.036 6.576 ;
  LAYER M2 ;
        RECT 31.564 6.48 34.036 6.512 ;
  LAYER M2 ;
        RECT 31.564 6.416 34.036 6.448 ;
  LAYER M2 ;
        RECT 31.564 6.352 34.036 6.384 ;
  LAYER M2 ;
        RECT 31.564 6.288 34.036 6.32 ;
  LAYER M2 ;
        RECT 31.564 6.224 34.036 6.256 ;
  LAYER M2 ;
        RECT 31.564 6.16 34.036 6.192 ;
  LAYER M2 ;
        RECT 31.564 6.096 34.036 6.128 ;
  LAYER M2 ;
        RECT 31.564 6.032 34.036 6.064 ;
  LAYER M2 ;
        RECT 31.564 5.968 34.036 6 ;
  LAYER M2 ;
        RECT 31.564 5.904 34.036 5.936 ;
  LAYER M2 ;
        RECT 31.564 5.84 34.036 5.872 ;
  LAYER M2 ;
        RECT 31.564 5.776 34.036 5.808 ;
  LAYER M2 ;
        RECT 31.564 5.712 34.036 5.744 ;
  LAYER M2 ;
        RECT 31.564 5.648 34.036 5.68 ;
  LAYER M2 ;
        RECT 31.564 5.584 34.036 5.616 ;
  LAYER M2 ;
        RECT 31.564 5.52 34.036 5.552 ;
  LAYER M2 ;
        RECT 31.564 5.456 34.036 5.488 ;
  LAYER M2 ;
        RECT 31.564 5.392 34.036 5.424 ;
  LAYER M2 ;
        RECT 31.564 5.328 34.036 5.36 ;
  LAYER M2 ;
        RECT 31.564 5.264 34.036 5.296 ;
  LAYER M2 ;
        RECT 31.564 5.2 34.036 5.232 ;
  LAYER M2 ;
        RECT 31.564 5.136 34.036 5.168 ;
  LAYER M2 ;
        RECT 31.564 5.072 34.036 5.104 ;
  LAYER M3 ;
        RECT 31.584 4.92 31.616 7.428 ;
  LAYER M3 ;
        RECT 31.648 4.92 31.68 7.428 ;
  LAYER M3 ;
        RECT 31.712 4.92 31.744 7.428 ;
  LAYER M3 ;
        RECT 31.776 4.92 31.808 7.428 ;
  LAYER M3 ;
        RECT 31.84 4.92 31.872 7.428 ;
  LAYER M3 ;
        RECT 31.904 4.92 31.936 7.428 ;
  LAYER M3 ;
        RECT 31.968 4.92 32 7.428 ;
  LAYER M3 ;
        RECT 32.032 4.92 32.064 7.428 ;
  LAYER M3 ;
        RECT 32.096 4.92 32.128 7.428 ;
  LAYER M3 ;
        RECT 32.16 4.92 32.192 7.428 ;
  LAYER M3 ;
        RECT 32.224 4.92 32.256 7.428 ;
  LAYER M3 ;
        RECT 32.288 4.92 32.32 7.428 ;
  LAYER M3 ;
        RECT 32.352 4.92 32.384 7.428 ;
  LAYER M3 ;
        RECT 32.416 4.92 32.448 7.428 ;
  LAYER M3 ;
        RECT 32.48 4.92 32.512 7.428 ;
  LAYER M3 ;
        RECT 32.544 4.92 32.576 7.428 ;
  LAYER M3 ;
        RECT 32.608 4.92 32.64 7.428 ;
  LAYER M3 ;
        RECT 32.672 4.92 32.704 7.428 ;
  LAYER M3 ;
        RECT 32.736 4.92 32.768 7.428 ;
  LAYER M3 ;
        RECT 32.8 4.92 32.832 7.428 ;
  LAYER M3 ;
        RECT 32.864 4.92 32.896 7.428 ;
  LAYER M3 ;
        RECT 32.928 4.92 32.96 7.428 ;
  LAYER M3 ;
        RECT 32.992 4.92 33.024 7.428 ;
  LAYER M3 ;
        RECT 33.056 4.92 33.088 7.428 ;
  LAYER M3 ;
        RECT 33.12 4.92 33.152 7.428 ;
  LAYER M3 ;
        RECT 33.184 4.92 33.216 7.428 ;
  LAYER M3 ;
        RECT 33.248 4.92 33.28 7.428 ;
  LAYER M3 ;
        RECT 33.312 4.92 33.344 7.428 ;
  LAYER M3 ;
        RECT 33.376 4.92 33.408 7.428 ;
  LAYER M3 ;
        RECT 33.44 4.92 33.472 7.428 ;
  LAYER M3 ;
        RECT 33.504 4.92 33.536 7.428 ;
  LAYER M3 ;
        RECT 33.568 4.92 33.6 7.428 ;
  LAYER M3 ;
        RECT 33.632 4.92 33.664 7.428 ;
  LAYER M3 ;
        RECT 33.696 4.92 33.728 7.428 ;
  LAYER M3 ;
        RECT 33.76 4.92 33.792 7.428 ;
  LAYER M3 ;
        RECT 33.824 4.92 33.856 7.428 ;
  LAYER M3 ;
        RECT 33.888 4.92 33.92 7.428 ;
  LAYER M3 ;
        RECT 33.984 4.92 34.016 7.428 ;
  LAYER M1 ;
        RECT 31.599 4.956 31.601 7.392 ;
  LAYER M1 ;
        RECT 31.679 4.956 31.681 7.392 ;
  LAYER M1 ;
        RECT 31.759 4.956 31.761 7.392 ;
  LAYER M1 ;
        RECT 31.839 4.956 31.841 7.392 ;
  LAYER M1 ;
        RECT 31.919 4.956 31.921 7.392 ;
  LAYER M1 ;
        RECT 31.999 4.956 32.001 7.392 ;
  LAYER M1 ;
        RECT 32.079 4.956 32.081 7.392 ;
  LAYER M1 ;
        RECT 32.159 4.956 32.161 7.392 ;
  LAYER M1 ;
        RECT 32.239 4.956 32.241 7.392 ;
  LAYER M1 ;
        RECT 32.319 4.956 32.321 7.392 ;
  LAYER M1 ;
        RECT 32.399 4.956 32.401 7.392 ;
  LAYER M1 ;
        RECT 32.479 4.956 32.481 7.392 ;
  LAYER M1 ;
        RECT 32.559 4.956 32.561 7.392 ;
  LAYER M1 ;
        RECT 32.639 4.956 32.641 7.392 ;
  LAYER M1 ;
        RECT 32.719 4.956 32.721 7.392 ;
  LAYER M1 ;
        RECT 32.799 4.956 32.801 7.392 ;
  LAYER M1 ;
        RECT 32.879 4.956 32.881 7.392 ;
  LAYER M1 ;
        RECT 32.959 4.956 32.961 7.392 ;
  LAYER M1 ;
        RECT 33.039 4.956 33.041 7.392 ;
  LAYER M1 ;
        RECT 33.119 4.956 33.121 7.392 ;
  LAYER M1 ;
        RECT 33.199 4.956 33.201 7.392 ;
  LAYER M1 ;
        RECT 33.279 4.956 33.281 7.392 ;
  LAYER M1 ;
        RECT 33.359 4.956 33.361 7.392 ;
  LAYER M1 ;
        RECT 33.439 4.956 33.441 7.392 ;
  LAYER M1 ;
        RECT 33.519 4.956 33.521 7.392 ;
  LAYER M1 ;
        RECT 33.599 4.956 33.601 7.392 ;
  LAYER M1 ;
        RECT 33.679 4.956 33.681 7.392 ;
  LAYER M1 ;
        RECT 33.759 4.956 33.761 7.392 ;
  LAYER M1 ;
        RECT 33.839 4.956 33.841 7.392 ;
  LAYER M1 ;
        RECT 33.919 4.956 33.921 7.392 ;
  LAYER M2 ;
        RECT 31.6 7.391 34 7.393 ;
  LAYER M2 ;
        RECT 31.6 7.307 34 7.309 ;
  LAYER M2 ;
        RECT 31.6 7.223 34 7.225 ;
  LAYER M2 ;
        RECT 31.6 7.139 34 7.141 ;
  LAYER M2 ;
        RECT 31.6 7.055 34 7.057 ;
  LAYER M2 ;
        RECT 31.6 6.971 34 6.973 ;
  LAYER M2 ;
        RECT 31.6 6.887 34 6.889 ;
  LAYER M2 ;
        RECT 31.6 6.803 34 6.805 ;
  LAYER M2 ;
        RECT 31.6 6.719 34 6.721 ;
  LAYER M2 ;
        RECT 31.6 6.635 34 6.637 ;
  LAYER M2 ;
        RECT 31.6 6.551 34 6.553 ;
  LAYER M2 ;
        RECT 31.6 6.467 34 6.469 ;
  LAYER M2 ;
        RECT 31.6 6.3835 34 6.3855 ;
  LAYER M2 ;
        RECT 31.6 6.299 34 6.301 ;
  LAYER M2 ;
        RECT 31.6 6.215 34 6.217 ;
  LAYER M2 ;
        RECT 31.6 6.131 34 6.133 ;
  LAYER M2 ;
        RECT 31.6 6.047 34 6.049 ;
  LAYER M2 ;
        RECT 31.6 5.963 34 5.965 ;
  LAYER M2 ;
        RECT 31.6 5.879 34 5.881 ;
  LAYER M2 ;
        RECT 31.6 5.795 34 5.797 ;
  LAYER M2 ;
        RECT 31.6 5.711 34 5.713 ;
  LAYER M2 ;
        RECT 31.6 5.627 34 5.629 ;
  LAYER M2 ;
        RECT 31.6 5.543 34 5.545 ;
  LAYER M2 ;
        RECT 31.6 5.459 34 5.461 ;
  LAYER M2 ;
        RECT 31.6 5.375 34 5.377 ;
  LAYER M2 ;
        RECT 31.6 5.291 34 5.293 ;
  LAYER M2 ;
        RECT 31.6 5.207 34 5.209 ;
  LAYER M2 ;
        RECT 31.6 5.123 34 5.125 ;
  LAYER M2 ;
        RECT 31.6 5.039 34 5.041 ;
  LAYER M1 ;
        RECT 31.584 1.98 31.616 4.488 ;
  LAYER M1 ;
        RECT 31.648 1.98 31.68 4.488 ;
  LAYER M1 ;
        RECT 31.712 1.98 31.744 4.488 ;
  LAYER M1 ;
        RECT 31.776 1.98 31.808 4.488 ;
  LAYER M1 ;
        RECT 31.84 1.98 31.872 4.488 ;
  LAYER M1 ;
        RECT 31.904 1.98 31.936 4.488 ;
  LAYER M1 ;
        RECT 31.968 1.98 32 4.488 ;
  LAYER M1 ;
        RECT 32.032 1.98 32.064 4.488 ;
  LAYER M1 ;
        RECT 32.096 1.98 32.128 4.488 ;
  LAYER M1 ;
        RECT 32.16 1.98 32.192 4.488 ;
  LAYER M1 ;
        RECT 32.224 1.98 32.256 4.488 ;
  LAYER M1 ;
        RECT 32.288 1.98 32.32 4.488 ;
  LAYER M1 ;
        RECT 32.352 1.98 32.384 4.488 ;
  LAYER M1 ;
        RECT 32.416 1.98 32.448 4.488 ;
  LAYER M1 ;
        RECT 32.48 1.98 32.512 4.488 ;
  LAYER M1 ;
        RECT 32.544 1.98 32.576 4.488 ;
  LAYER M1 ;
        RECT 32.608 1.98 32.64 4.488 ;
  LAYER M1 ;
        RECT 32.672 1.98 32.704 4.488 ;
  LAYER M1 ;
        RECT 32.736 1.98 32.768 4.488 ;
  LAYER M1 ;
        RECT 32.8 1.98 32.832 4.488 ;
  LAYER M1 ;
        RECT 32.864 1.98 32.896 4.488 ;
  LAYER M1 ;
        RECT 32.928 1.98 32.96 4.488 ;
  LAYER M1 ;
        RECT 32.992 1.98 33.024 4.488 ;
  LAYER M1 ;
        RECT 33.056 1.98 33.088 4.488 ;
  LAYER M1 ;
        RECT 33.12 1.98 33.152 4.488 ;
  LAYER M1 ;
        RECT 33.184 1.98 33.216 4.488 ;
  LAYER M1 ;
        RECT 33.248 1.98 33.28 4.488 ;
  LAYER M1 ;
        RECT 33.312 1.98 33.344 4.488 ;
  LAYER M1 ;
        RECT 33.376 1.98 33.408 4.488 ;
  LAYER M1 ;
        RECT 33.44 1.98 33.472 4.488 ;
  LAYER M1 ;
        RECT 33.504 1.98 33.536 4.488 ;
  LAYER M1 ;
        RECT 33.568 1.98 33.6 4.488 ;
  LAYER M1 ;
        RECT 33.632 1.98 33.664 4.488 ;
  LAYER M1 ;
        RECT 33.696 1.98 33.728 4.488 ;
  LAYER M1 ;
        RECT 33.76 1.98 33.792 4.488 ;
  LAYER M1 ;
        RECT 33.824 1.98 33.856 4.488 ;
  LAYER M1 ;
        RECT 33.888 1.98 33.92 4.488 ;
  LAYER M2 ;
        RECT 31.564 4.372 34.036 4.404 ;
  LAYER M2 ;
        RECT 31.564 4.308 34.036 4.34 ;
  LAYER M2 ;
        RECT 31.564 4.244 34.036 4.276 ;
  LAYER M2 ;
        RECT 31.564 4.18 34.036 4.212 ;
  LAYER M2 ;
        RECT 31.564 4.116 34.036 4.148 ;
  LAYER M2 ;
        RECT 31.564 4.052 34.036 4.084 ;
  LAYER M2 ;
        RECT 31.564 3.988 34.036 4.02 ;
  LAYER M2 ;
        RECT 31.564 3.924 34.036 3.956 ;
  LAYER M2 ;
        RECT 31.564 3.86 34.036 3.892 ;
  LAYER M2 ;
        RECT 31.564 3.796 34.036 3.828 ;
  LAYER M2 ;
        RECT 31.564 3.732 34.036 3.764 ;
  LAYER M2 ;
        RECT 31.564 3.668 34.036 3.7 ;
  LAYER M2 ;
        RECT 31.564 3.604 34.036 3.636 ;
  LAYER M2 ;
        RECT 31.564 3.54 34.036 3.572 ;
  LAYER M2 ;
        RECT 31.564 3.476 34.036 3.508 ;
  LAYER M2 ;
        RECT 31.564 3.412 34.036 3.444 ;
  LAYER M2 ;
        RECT 31.564 3.348 34.036 3.38 ;
  LAYER M2 ;
        RECT 31.564 3.284 34.036 3.316 ;
  LAYER M2 ;
        RECT 31.564 3.22 34.036 3.252 ;
  LAYER M2 ;
        RECT 31.564 3.156 34.036 3.188 ;
  LAYER M2 ;
        RECT 31.564 3.092 34.036 3.124 ;
  LAYER M2 ;
        RECT 31.564 3.028 34.036 3.06 ;
  LAYER M2 ;
        RECT 31.564 2.964 34.036 2.996 ;
  LAYER M2 ;
        RECT 31.564 2.9 34.036 2.932 ;
  LAYER M2 ;
        RECT 31.564 2.836 34.036 2.868 ;
  LAYER M2 ;
        RECT 31.564 2.772 34.036 2.804 ;
  LAYER M2 ;
        RECT 31.564 2.708 34.036 2.74 ;
  LAYER M2 ;
        RECT 31.564 2.644 34.036 2.676 ;
  LAYER M2 ;
        RECT 31.564 2.58 34.036 2.612 ;
  LAYER M2 ;
        RECT 31.564 2.516 34.036 2.548 ;
  LAYER M2 ;
        RECT 31.564 2.452 34.036 2.484 ;
  LAYER M2 ;
        RECT 31.564 2.388 34.036 2.42 ;
  LAYER M2 ;
        RECT 31.564 2.324 34.036 2.356 ;
  LAYER M2 ;
        RECT 31.564 2.26 34.036 2.292 ;
  LAYER M2 ;
        RECT 31.564 2.196 34.036 2.228 ;
  LAYER M2 ;
        RECT 31.564 2.132 34.036 2.164 ;
  LAYER M3 ;
        RECT 31.584 1.98 31.616 4.488 ;
  LAYER M3 ;
        RECT 31.648 1.98 31.68 4.488 ;
  LAYER M3 ;
        RECT 31.712 1.98 31.744 4.488 ;
  LAYER M3 ;
        RECT 31.776 1.98 31.808 4.488 ;
  LAYER M3 ;
        RECT 31.84 1.98 31.872 4.488 ;
  LAYER M3 ;
        RECT 31.904 1.98 31.936 4.488 ;
  LAYER M3 ;
        RECT 31.968 1.98 32 4.488 ;
  LAYER M3 ;
        RECT 32.032 1.98 32.064 4.488 ;
  LAYER M3 ;
        RECT 32.096 1.98 32.128 4.488 ;
  LAYER M3 ;
        RECT 32.16 1.98 32.192 4.488 ;
  LAYER M3 ;
        RECT 32.224 1.98 32.256 4.488 ;
  LAYER M3 ;
        RECT 32.288 1.98 32.32 4.488 ;
  LAYER M3 ;
        RECT 32.352 1.98 32.384 4.488 ;
  LAYER M3 ;
        RECT 32.416 1.98 32.448 4.488 ;
  LAYER M3 ;
        RECT 32.48 1.98 32.512 4.488 ;
  LAYER M3 ;
        RECT 32.544 1.98 32.576 4.488 ;
  LAYER M3 ;
        RECT 32.608 1.98 32.64 4.488 ;
  LAYER M3 ;
        RECT 32.672 1.98 32.704 4.488 ;
  LAYER M3 ;
        RECT 32.736 1.98 32.768 4.488 ;
  LAYER M3 ;
        RECT 32.8 1.98 32.832 4.488 ;
  LAYER M3 ;
        RECT 32.864 1.98 32.896 4.488 ;
  LAYER M3 ;
        RECT 32.928 1.98 32.96 4.488 ;
  LAYER M3 ;
        RECT 32.992 1.98 33.024 4.488 ;
  LAYER M3 ;
        RECT 33.056 1.98 33.088 4.488 ;
  LAYER M3 ;
        RECT 33.12 1.98 33.152 4.488 ;
  LAYER M3 ;
        RECT 33.184 1.98 33.216 4.488 ;
  LAYER M3 ;
        RECT 33.248 1.98 33.28 4.488 ;
  LAYER M3 ;
        RECT 33.312 1.98 33.344 4.488 ;
  LAYER M3 ;
        RECT 33.376 1.98 33.408 4.488 ;
  LAYER M3 ;
        RECT 33.44 1.98 33.472 4.488 ;
  LAYER M3 ;
        RECT 33.504 1.98 33.536 4.488 ;
  LAYER M3 ;
        RECT 33.568 1.98 33.6 4.488 ;
  LAYER M3 ;
        RECT 33.632 1.98 33.664 4.488 ;
  LAYER M3 ;
        RECT 33.696 1.98 33.728 4.488 ;
  LAYER M3 ;
        RECT 33.76 1.98 33.792 4.488 ;
  LAYER M3 ;
        RECT 33.824 1.98 33.856 4.488 ;
  LAYER M3 ;
        RECT 33.888 1.98 33.92 4.488 ;
  LAYER M3 ;
        RECT 33.984 1.98 34.016 4.488 ;
  LAYER M1 ;
        RECT 31.599 2.016 31.601 4.452 ;
  LAYER M1 ;
        RECT 31.679 2.016 31.681 4.452 ;
  LAYER M1 ;
        RECT 31.759 2.016 31.761 4.452 ;
  LAYER M1 ;
        RECT 31.839 2.016 31.841 4.452 ;
  LAYER M1 ;
        RECT 31.919 2.016 31.921 4.452 ;
  LAYER M1 ;
        RECT 31.999 2.016 32.001 4.452 ;
  LAYER M1 ;
        RECT 32.079 2.016 32.081 4.452 ;
  LAYER M1 ;
        RECT 32.159 2.016 32.161 4.452 ;
  LAYER M1 ;
        RECT 32.239 2.016 32.241 4.452 ;
  LAYER M1 ;
        RECT 32.319 2.016 32.321 4.452 ;
  LAYER M1 ;
        RECT 32.399 2.016 32.401 4.452 ;
  LAYER M1 ;
        RECT 32.479 2.016 32.481 4.452 ;
  LAYER M1 ;
        RECT 32.559 2.016 32.561 4.452 ;
  LAYER M1 ;
        RECT 32.639 2.016 32.641 4.452 ;
  LAYER M1 ;
        RECT 32.719 2.016 32.721 4.452 ;
  LAYER M1 ;
        RECT 32.799 2.016 32.801 4.452 ;
  LAYER M1 ;
        RECT 32.879 2.016 32.881 4.452 ;
  LAYER M1 ;
        RECT 32.959 2.016 32.961 4.452 ;
  LAYER M1 ;
        RECT 33.039 2.016 33.041 4.452 ;
  LAYER M1 ;
        RECT 33.119 2.016 33.121 4.452 ;
  LAYER M1 ;
        RECT 33.199 2.016 33.201 4.452 ;
  LAYER M1 ;
        RECT 33.279 2.016 33.281 4.452 ;
  LAYER M1 ;
        RECT 33.359 2.016 33.361 4.452 ;
  LAYER M1 ;
        RECT 33.439 2.016 33.441 4.452 ;
  LAYER M1 ;
        RECT 33.519 2.016 33.521 4.452 ;
  LAYER M1 ;
        RECT 33.599 2.016 33.601 4.452 ;
  LAYER M1 ;
        RECT 33.679 2.016 33.681 4.452 ;
  LAYER M1 ;
        RECT 33.759 2.016 33.761 4.452 ;
  LAYER M1 ;
        RECT 33.839 2.016 33.841 4.452 ;
  LAYER M1 ;
        RECT 33.919 2.016 33.921 4.452 ;
  LAYER M2 ;
        RECT 31.6 4.451 34 4.453 ;
  LAYER M2 ;
        RECT 31.6 4.367 34 4.369 ;
  LAYER M2 ;
        RECT 31.6 4.283 34 4.285 ;
  LAYER M2 ;
        RECT 31.6 4.199 34 4.201 ;
  LAYER M2 ;
        RECT 31.6 4.115 34 4.117 ;
  LAYER M2 ;
        RECT 31.6 4.031 34 4.033 ;
  LAYER M2 ;
        RECT 31.6 3.947 34 3.949 ;
  LAYER M2 ;
        RECT 31.6 3.863 34 3.865 ;
  LAYER M2 ;
        RECT 31.6 3.779 34 3.781 ;
  LAYER M2 ;
        RECT 31.6 3.695 34 3.697 ;
  LAYER M2 ;
        RECT 31.6 3.611 34 3.613 ;
  LAYER M2 ;
        RECT 31.6 3.527 34 3.529 ;
  LAYER M2 ;
        RECT 31.6 3.4435 34 3.4455 ;
  LAYER M2 ;
        RECT 31.6 3.359 34 3.361 ;
  LAYER M2 ;
        RECT 31.6 3.275 34 3.277 ;
  LAYER M2 ;
        RECT 31.6 3.191 34 3.193 ;
  LAYER M2 ;
        RECT 31.6 3.107 34 3.109 ;
  LAYER M2 ;
        RECT 31.6 3.023 34 3.025 ;
  LAYER M2 ;
        RECT 31.6 2.939 34 2.941 ;
  LAYER M2 ;
        RECT 31.6 2.855 34 2.857 ;
  LAYER M2 ;
        RECT 31.6 2.771 34 2.773 ;
  LAYER M2 ;
        RECT 31.6 2.687 34 2.689 ;
  LAYER M2 ;
        RECT 31.6 2.603 34 2.605 ;
  LAYER M2 ;
        RECT 31.6 2.519 34 2.521 ;
  LAYER M2 ;
        RECT 31.6 2.435 34 2.437 ;
  LAYER M2 ;
        RECT 31.6 2.351 34 2.353 ;
  LAYER M2 ;
        RECT 31.6 2.267 34 2.269 ;
  LAYER M2 ;
        RECT 31.6 2.183 34 2.185 ;
  LAYER M2 ;
        RECT 31.6 2.099 34 2.101 ;
  LAYER M1 ;
        RECT 34.464 13.74 34.496 16.248 ;
  LAYER M1 ;
        RECT 34.528 13.74 34.56 16.248 ;
  LAYER M1 ;
        RECT 34.592 13.74 34.624 16.248 ;
  LAYER M1 ;
        RECT 34.656 13.74 34.688 16.248 ;
  LAYER M1 ;
        RECT 34.72 13.74 34.752 16.248 ;
  LAYER M1 ;
        RECT 34.784 13.74 34.816 16.248 ;
  LAYER M1 ;
        RECT 34.848 13.74 34.88 16.248 ;
  LAYER M1 ;
        RECT 34.912 13.74 34.944 16.248 ;
  LAYER M1 ;
        RECT 34.976 13.74 35.008 16.248 ;
  LAYER M1 ;
        RECT 35.04 13.74 35.072 16.248 ;
  LAYER M1 ;
        RECT 35.104 13.74 35.136 16.248 ;
  LAYER M1 ;
        RECT 35.168 13.74 35.2 16.248 ;
  LAYER M1 ;
        RECT 35.232 13.74 35.264 16.248 ;
  LAYER M1 ;
        RECT 35.296 13.74 35.328 16.248 ;
  LAYER M1 ;
        RECT 35.36 13.74 35.392 16.248 ;
  LAYER M1 ;
        RECT 35.424 13.74 35.456 16.248 ;
  LAYER M1 ;
        RECT 35.488 13.74 35.52 16.248 ;
  LAYER M1 ;
        RECT 35.552 13.74 35.584 16.248 ;
  LAYER M1 ;
        RECT 35.616 13.74 35.648 16.248 ;
  LAYER M1 ;
        RECT 35.68 13.74 35.712 16.248 ;
  LAYER M1 ;
        RECT 35.744 13.74 35.776 16.248 ;
  LAYER M1 ;
        RECT 35.808 13.74 35.84 16.248 ;
  LAYER M1 ;
        RECT 35.872 13.74 35.904 16.248 ;
  LAYER M1 ;
        RECT 35.936 13.74 35.968 16.248 ;
  LAYER M1 ;
        RECT 36 13.74 36.032 16.248 ;
  LAYER M1 ;
        RECT 36.064 13.74 36.096 16.248 ;
  LAYER M1 ;
        RECT 36.128 13.74 36.16 16.248 ;
  LAYER M1 ;
        RECT 36.192 13.74 36.224 16.248 ;
  LAYER M1 ;
        RECT 36.256 13.74 36.288 16.248 ;
  LAYER M1 ;
        RECT 36.32 13.74 36.352 16.248 ;
  LAYER M1 ;
        RECT 36.384 13.74 36.416 16.248 ;
  LAYER M1 ;
        RECT 36.448 13.74 36.48 16.248 ;
  LAYER M1 ;
        RECT 36.512 13.74 36.544 16.248 ;
  LAYER M1 ;
        RECT 36.576 13.74 36.608 16.248 ;
  LAYER M1 ;
        RECT 36.64 13.74 36.672 16.248 ;
  LAYER M1 ;
        RECT 36.704 13.74 36.736 16.248 ;
  LAYER M1 ;
        RECT 36.768 13.74 36.8 16.248 ;
  LAYER M2 ;
        RECT 34.444 16.132 36.916 16.164 ;
  LAYER M2 ;
        RECT 34.444 16.068 36.916 16.1 ;
  LAYER M2 ;
        RECT 34.444 16.004 36.916 16.036 ;
  LAYER M2 ;
        RECT 34.444 15.94 36.916 15.972 ;
  LAYER M2 ;
        RECT 34.444 15.876 36.916 15.908 ;
  LAYER M2 ;
        RECT 34.444 15.812 36.916 15.844 ;
  LAYER M2 ;
        RECT 34.444 15.748 36.916 15.78 ;
  LAYER M2 ;
        RECT 34.444 15.684 36.916 15.716 ;
  LAYER M2 ;
        RECT 34.444 15.62 36.916 15.652 ;
  LAYER M2 ;
        RECT 34.444 15.556 36.916 15.588 ;
  LAYER M2 ;
        RECT 34.444 15.492 36.916 15.524 ;
  LAYER M2 ;
        RECT 34.444 15.428 36.916 15.46 ;
  LAYER M2 ;
        RECT 34.444 15.364 36.916 15.396 ;
  LAYER M2 ;
        RECT 34.444 15.3 36.916 15.332 ;
  LAYER M2 ;
        RECT 34.444 15.236 36.916 15.268 ;
  LAYER M2 ;
        RECT 34.444 15.172 36.916 15.204 ;
  LAYER M2 ;
        RECT 34.444 15.108 36.916 15.14 ;
  LAYER M2 ;
        RECT 34.444 15.044 36.916 15.076 ;
  LAYER M2 ;
        RECT 34.444 14.98 36.916 15.012 ;
  LAYER M2 ;
        RECT 34.444 14.916 36.916 14.948 ;
  LAYER M2 ;
        RECT 34.444 14.852 36.916 14.884 ;
  LAYER M2 ;
        RECT 34.444 14.788 36.916 14.82 ;
  LAYER M2 ;
        RECT 34.444 14.724 36.916 14.756 ;
  LAYER M2 ;
        RECT 34.444 14.66 36.916 14.692 ;
  LAYER M2 ;
        RECT 34.444 14.596 36.916 14.628 ;
  LAYER M2 ;
        RECT 34.444 14.532 36.916 14.564 ;
  LAYER M2 ;
        RECT 34.444 14.468 36.916 14.5 ;
  LAYER M2 ;
        RECT 34.444 14.404 36.916 14.436 ;
  LAYER M2 ;
        RECT 34.444 14.34 36.916 14.372 ;
  LAYER M2 ;
        RECT 34.444 14.276 36.916 14.308 ;
  LAYER M2 ;
        RECT 34.444 14.212 36.916 14.244 ;
  LAYER M2 ;
        RECT 34.444 14.148 36.916 14.18 ;
  LAYER M2 ;
        RECT 34.444 14.084 36.916 14.116 ;
  LAYER M2 ;
        RECT 34.444 14.02 36.916 14.052 ;
  LAYER M2 ;
        RECT 34.444 13.956 36.916 13.988 ;
  LAYER M2 ;
        RECT 34.444 13.892 36.916 13.924 ;
  LAYER M3 ;
        RECT 34.464 13.74 34.496 16.248 ;
  LAYER M3 ;
        RECT 34.528 13.74 34.56 16.248 ;
  LAYER M3 ;
        RECT 34.592 13.74 34.624 16.248 ;
  LAYER M3 ;
        RECT 34.656 13.74 34.688 16.248 ;
  LAYER M3 ;
        RECT 34.72 13.74 34.752 16.248 ;
  LAYER M3 ;
        RECT 34.784 13.74 34.816 16.248 ;
  LAYER M3 ;
        RECT 34.848 13.74 34.88 16.248 ;
  LAYER M3 ;
        RECT 34.912 13.74 34.944 16.248 ;
  LAYER M3 ;
        RECT 34.976 13.74 35.008 16.248 ;
  LAYER M3 ;
        RECT 35.04 13.74 35.072 16.248 ;
  LAYER M3 ;
        RECT 35.104 13.74 35.136 16.248 ;
  LAYER M3 ;
        RECT 35.168 13.74 35.2 16.248 ;
  LAYER M3 ;
        RECT 35.232 13.74 35.264 16.248 ;
  LAYER M3 ;
        RECT 35.296 13.74 35.328 16.248 ;
  LAYER M3 ;
        RECT 35.36 13.74 35.392 16.248 ;
  LAYER M3 ;
        RECT 35.424 13.74 35.456 16.248 ;
  LAYER M3 ;
        RECT 35.488 13.74 35.52 16.248 ;
  LAYER M3 ;
        RECT 35.552 13.74 35.584 16.248 ;
  LAYER M3 ;
        RECT 35.616 13.74 35.648 16.248 ;
  LAYER M3 ;
        RECT 35.68 13.74 35.712 16.248 ;
  LAYER M3 ;
        RECT 35.744 13.74 35.776 16.248 ;
  LAYER M3 ;
        RECT 35.808 13.74 35.84 16.248 ;
  LAYER M3 ;
        RECT 35.872 13.74 35.904 16.248 ;
  LAYER M3 ;
        RECT 35.936 13.74 35.968 16.248 ;
  LAYER M3 ;
        RECT 36 13.74 36.032 16.248 ;
  LAYER M3 ;
        RECT 36.064 13.74 36.096 16.248 ;
  LAYER M3 ;
        RECT 36.128 13.74 36.16 16.248 ;
  LAYER M3 ;
        RECT 36.192 13.74 36.224 16.248 ;
  LAYER M3 ;
        RECT 36.256 13.74 36.288 16.248 ;
  LAYER M3 ;
        RECT 36.32 13.74 36.352 16.248 ;
  LAYER M3 ;
        RECT 36.384 13.74 36.416 16.248 ;
  LAYER M3 ;
        RECT 36.448 13.74 36.48 16.248 ;
  LAYER M3 ;
        RECT 36.512 13.74 36.544 16.248 ;
  LAYER M3 ;
        RECT 36.576 13.74 36.608 16.248 ;
  LAYER M3 ;
        RECT 36.64 13.74 36.672 16.248 ;
  LAYER M3 ;
        RECT 36.704 13.74 36.736 16.248 ;
  LAYER M3 ;
        RECT 36.768 13.74 36.8 16.248 ;
  LAYER M3 ;
        RECT 36.864 13.74 36.896 16.248 ;
  LAYER M1 ;
        RECT 34.479 13.776 34.481 16.212 ;
  LAYER M1 ;
        RECT 34.559 13.776 34.561 16.212 ;
  LAYER M1 ;
        RECT 34.639 13.776 34.641 16.212 ;
  LAYER M1 ;
        RECT 34.719 13.776 34.721 16.212 ;
  LAYER M1 ;
        RECT 34.799 13.776 34.801 16.212 ;
  LAYER M1 ;
        RECT 34.879 13.776 34.881 16.212 ;
  LAYER M1 ;
        RECT 34.959 13.776 34.961 16.212 ;
  LAYER M1 ;
        RECT 35.039 13.776 35.041 16.212 ;
  LAYER M1 ;
        RECT 35.119 13.776 35.121 16.212 ;
  LAYER M1 ;
        RECT 35.199 13.776 35.201 16.212 ;
  LAYER M1 ;
        RECT 35.279 13.776 35.281 16.212 ;
  LAYER M1 ;
        RECT 35.359 13.776 35.361 16.212 ;
  LAYER M1 ;
        RECT 35.439 13.776 35.441 16.212 ;
  LAYER M1 ;
        RECT 35.519 13.776 35.521 16.212 ;
  LAYER M1 ;
        RECT 35.599 13.776 35.601 16.212 ;
  LAYER M1 ;
        RECT 35.679 13.776 35.681 16.212 ;
  LAYER M1 ;
        RECT 35.759 13.776 35.761 16.212 ;
  LAYER M1 ;
        RECT 35.839 13.776 35.841 16.212 ;
  LAYER M1 ;
        RECT 35.919 13.776 35.921 16.212 ;
  LAYER M1 ;
        RECT 35.999 13.776 36.001 16.212 ;
  LAYER M1 ;
        RECT 36.079 13.776 36.081 16.212 ;
  LAYER M1 ;
        RECT 36.159 13.776 36.161 16.212 ;
  LAYER M1 ;
        RECT 36.239 13.776 36.241 16.212 ;
  LAYER M1 ;
        RECT 36.319 13.776 36.321 16.212 ;
  LAYER M1 ;
        RECT 36.399 13.776 36.401 16.212 ;
  LAYER M1 ;
        RECT 36.479 13.776 36.481 16.212 ;
  LAYER M1 ;
        RECT 36.559 13.776 36.561 16.212 ;
  LAYER M1 ;
        RECT 36.639 13.776 36.641 16.212 ;
  LAYER M1 ;
        RECT 36.719 13.776 36.721 16.212 ;
  LAYER M1 ;
        RECT 36.799 13.776 36.801 16.212 ;
  LAYER M2 ;
        RECT 34.48 16.211 36.88 16.213 ;
  LAYER M2 ;
        RECT 34.48 16.127 36.88 16.129 ;
  LAYER M2 ;
        RECT 34.48 16.043 36.88 16.045 ;
  LAYER M2 ;
        RECT 34.48 15.959 36.88 15.961 ;
  LAYER M2 ;
        RECT 34.48 15.875 36.88 15.877 ;
  LAYER M2 ;
        RECT 34.48 15.791 36.88 15.793 ;
  LAYER M2 ;
        RECT 34.48 15.707 36.88 15.709 ;
  LAYER M2 ;
        RECT 34.48 15.623 36.88 15.625 ;
  LAYER M2 ;
        RECT 34.48 15.539 36.88 15.541 ;
  LAYER M2 ;
        RECT 34.48 15.455 36.88 15.457 ;
  LAYER M2 ;
        RECT 34.48 15.371 36.88 15.373 ;
  LAYER M2 ;
        RECT 34.48 15.287 36.88 15.289 ;
  LAYER M2 ;
        RECT 34.48 15.2035 36.88 15.2055 ;
  LAYER M2 ;
        RECT 34.48 15.119 36.88 15.121 ;
  LAYER M2 ;
        RECT 34.48 15.035 36.88 15.037 ;
  LAYER M2 ;
        RECT 34.48 14.951 36.88 14.953 ;
  LAYER M2 ;
        RECT 34.48 14.867 36.88 14.869 ;
  LAYER M2 ;
        RECT 34.48 14.783 36.88 14.785 ;
  LAYER M2 ;
        RECT 34.48 14.699 36.88 14.701 ;
  LAYER M2 ;
        RECT 34.48 14.615 36.88 14.617 ;
  LAYER M2 ;
        RECT 34.48 14.531 36.88 14.533 ;
  LAYER M2 ;
        RECT 34.48 14.447 36.88 14.449 ;
  LAYER M2 ;
        RECT 34.48 14.363 36.88 14.365 ;
  LAYER M2 ;
        RECT 34.48 14.279 36.88 14.281 ;
  LAYER M2 ;
        RECT 34.48 14.195 36.88 14.197 ;
  LAYER M2 ;
        RECT 34.48 14.111 36.88 14.113 ;
  LAYER M2 ;
        RECT 34.48 14.027 36.88 14.029 ;
  LAYER M2 ;
        RECT 34.48 13.943 36.88 13.945 ;
  LAYER M2 ;
        RECT 34.48 13.859 36.88 13.861 ;
  LAYER M1 ;
        RECT 34.464 10.8 34.496 13.308 ;
  LAYER M1 ;
        RECT 34.528 10.8 34.56 13.308 ;
  LAYER M1 ;
        RECT 34.592 10.8 34.624 13.308 ;
  LAYER M1 ;
        RECT 34.656 10.8 34.688 13.308 ;
  LAYER M1 ;
        RECT 34.72 10.8 34.752 13.308 ;
  LAYER M1 ;
        RECT 34.784 10.8 34.816 13.308 ;
  LAYER M1 ;
        RECT 34.848 10.8 34.88 13.308 ;
  LAYER M1 ;
        RECT 34.912 10.8 34.944 13.308 ;
  LAYER M1 ;
        RECT 34.976 10.8 35.008 13.308 ;
  LAYER M1 ;
        RECT 35.04 10.8 35.072 13.308 ;
  LAYER M1 ;
        RECT 35.104 10.8 35.136 13.308 ;
  LAYER M1 ;
        RECT 35.168 10.8 35.2 13.308 ;
  LAYER M1 ;
        RECT 35.232 10.8 35.264 13.308 ;
  LAYER M1 ;
        RECT 35.296 10.8 35.328 13.308 ;
  LAYER M1 ;
        RECT 35.36 10.8 35.392 13.308 ;
  LAYER M1 ;
        RECT 35.424 10.8 35.456 13.308 ;
  LAYER M1 ;
        RECT 35.488 10.8 35.52 13.308 ;
  LAYER M1 ;
        RECT 35.552 10.8 35.584 13.308 ;
  LAYER M1 ;
        RECT 35.616 10.8 35.648 13.308 ;
  LAYER M1 ;
        RECT 35.68 10.8 35.712 13.308 ;
  LAYER M1 ;
        RECT 35.744 10.8 35.776 13.308 ;
  LAYER M1 ;
        RECT 35.808 10.8 35.84 13.308 ;
  LAYER M1 ;
        RECT 35.872 10.8 35.904 13.308 ;
  LAYER M1 ;
        RECT 35.936 10.8 35.968 13.308 ;
  LAYER M1 ;
        RECT 36 10.8 36.032 13.308 ;
  LAYER M1 ;
        RECT 36.064 10.8 36.096 13.308 ;
  LAYER M1 ;
        RECT 36.128 10.8 36.16 13.308 ;
  LAYER M1 ;
        RECT 36.192 10.8 36.224 13.308 ;
  LAYER M1 ;
        RECT 36.256 10.8 36.288 13.308 ;
  LAYER M1 ;
        RECT 36.32 10.8 36.352 13.308 ;
  LAYER M1 ;
        RECT 36.384 10.8 36.416 13.308 ;
  LAYER M1 ;
        RECT 36.448 10.8 36.48 13.308 ;
  LAYER M1 ;
        RECT 36.512 10.8 36.544 13.308 ;
  LAYER M1 ;
        RECT 36.576 10.8 36.608 13.308 ;
  LAYER M1 ;
        RECT 36.64 10.8 36.672 13.308 ;
  LAYER M1 ;
        RECT 36.704 10.8 36.736 13.308 ;
  LAYER M1 ;
        RECT 36.768 10.8 36.8 13.308 ;
  LAYER M2 ;
        RECT 34.444 13.192 36.916 13.224 ;
  LAYER M2 ;
        RECT 34.444 13.128 36.916 13.16 ;
  LAYER M2 ;
        RECT 34.444 13.064 36.916 13.096 ;
  LAYER M2 ;
        RECT 34.444 13 36.916 13.032 ;
  LAYER M2 ;
        RECT 34.444 12.936 36.916 12.968 ;
  LAYER M2 ;
        RECT 34.444 12.872 36.916 12.904 ;
  LAYER M2 ;
        RECT 34.444 12.808 36.916 12.84 ;
  LAYER M2 ;
        RECT 34.444 12.744 36.916 12.776 ;
  LAYER M2 ;
        RECT 34.444 12.68 36.916 12.712 ;
  LAYER M2 ;
        RECT 34.444 12.616 36.916 12.648 ;
  LAYER M2 ;
        RECT 34.444 12.552 36.916 12.584 ;
  LAYER M2 ;
        RECT 34.444 12.488 36.916 12.52 ;
  LAYER M2 ;
        RECT 34.444 12.424 36.916 12.456 ;
  LAYER M2 ;
        RECT 34.444 12.36 36.916 12.392 ;
  LAYER M2 ;
        RECT 34.444 12.296 36.916 12.328 ;
  LAYER M2 ;
        RECT 34.444 12.232 36.916 12.264 ;
  LAYER M2 ;
        RECT 34.444 12.168 36.916 12.2 ;
  LAYER M2 ;
        RECT 34.444 12.104 36.916 12.136 ;
  LAYER M2 ;
        RECT 34.444 12.04 36.916 12.072 ;
  LAYER M2 ;
        RECT 34.444 11.976 36.916 12.008 ;
  LAYER M2 ;
        RECT 34.444 11.912 36.916 11.944 ;
  LAYER M2 ;
        RECT 34.444 11.848 36.916 11.88 ;
  LAYER M2 ;
        RECT 34.444 11.784 36.916 11.816 ;
  LAYER M2 ;
        RECT 34.444 11.72 36.916 11.752 ;
  LAYER M2 ;
        RECT 34.444 11.656 36.916 11.688 ;
  LAYER M2 ;
        RECT 34.444 11.592 36.916 11.624 ;
  LAYER M2 ;
        RECT 34.444 11.528 36.916 11.56 ;
  LAYER M2 ;
        RECT 34.444 11.464 36.916 11.496 ;
  LAYER M2 ;
        RECT 34.444 11.4 36.916 11.432 ;
  LAYER M2 ;
        RECT 34.444 11.336 36.916 11.368 ;
  LAYER M2 ;
        RECT 34.444 11.272 36.916 11.304 ;
  LAYER M2 ;
        RECT 34.444 11.208 36.916 11.24 ;
  LAYER M2 ;
        RECT 34.444 11.144 36.916 11.176 ;
  LAYER M2 ;
        RECT 34.444 11.08 36.916 11.112 ;
  LAYER M2 ;
        RECT 34.444 11.016 36.916 11.048 ;
  LAYER M2 ;
        RECT 34.444 10.952 36.916 10.984 ;
  LAYER M3 ;
        RECT 34.464 10.8 34.496 13.308 ;
  LAYER M3 ;
        RECT 34.528 10.8 34.56 13.308 ;
  LAYER M3 ;
        RECT 34.592 10.8 34.624 13.308 ;
  LAYER M3 ;
        RECT 34.656 10.8 34.688 13.308 ;
  LAYER M3 ;
        RECT 34.72 10.8 34.752 13.308 ;
  LAYER M3 ;
        RECT 34.784 10.8 34.816 13.308 ;
  LAYER M3 ;
        RECT 34.848 10.8 34.88 13.308 ;
  LAYER M3 ;
        RECT 34.912 10.8 34.944 13.308 ;
  LAYER M3 ;
        RECT 34.976 10.8 35.008 13.308 ;
  LAYER M3 ;
        RECT 35.04 10.8 35.072 13.308 ;
  LAYER M3 ;
        RECT 35.104 10.8 35.136 13.308 ;
  LAYER M3 ;
        RECT 35.168 10.8 35.2 13.308 ;
  LAYER M3 ;
        RECT 35.232 10.8 35.264 13.308 ;
  LAYER M3 ;
        RECT 35.296 10.8 35.328 13.308 ;
  LAYER M3 ;
        RECT 35.36 10.8 35.392 13.308 ;
  LAYER M3 ;
        RECT 35.424 10.8 35.456 13.308 ;
  LAYER M3 ;
        RECT 35.488 10.8 35.52 13.308 ;
  LAYER M3 ;
        RECT 35.552 10.8 35.584 13.308 ;
  LAYER M3 ;
        RECT 35.616 10.8 35.648 13.308 ;
  LAYER M3 ;
        RECT 35.68 10.8 35.712 13.308 ;
  LAYER M3 ;
        RECT 35.744 10.8 35.776 13.308 ;
  LAYER M3 ;
        RECT 35.808 10.8 35.84 13.308 ;
  LAYER M3 ;
        RECT 35.872 10.8 35.904 13.308 ;
  LAYER M3 ;
        RECT 35.936 10.8 35.968 13.308 ;
  LAYER M3 ;
        RECT 36 10.8 36.032 13.308 ;
  LAYER M3 ;
        RECT 36.064 10.8 36.096 13.308 ;
  LAYER M3 ;
        RECT 36.128 10.8 36.16 13.308 ;
  LAYER M3 ;
        RECT 36.192 10.8 36.224 13.308 ;
  LAYER M3 ;
        RECT 36.256 10.8 36.288 13.308 ;
  LAYER M3 ;
        RECT 36.32 10.8 36.352 13.308 ;
  LAYER M3 ;
        RECT 36.384 10.8 36.416 13.308 ;
  LAYER M3 ;
        RECT 36.448 10.8 36.48 13.308 ;
  LAYER M3 ;
        RECT 36.512 10.8 36.544 13.308 ;
  LAYER M3 ;
        RECT 36.576 10.8 36.608 13.308 ;
  LAYER M3 ;
        RECT 36.64 10.8 36.672 13.308 ;
  LAYER M3 ;
        RECT 36.704 10.8 36.736 13.308 ;
  LAYER M3 ;
        RECT 36.768 10.8 36.8 13.308 ;
  LAYER M3 ;
        RECT 36.864 10.8 36.896 13.308 ;
  LAYER M1 ;
        RECT 34.479 10.836 34.481 13.272 ;
  LAYER M1 ;
        RECT 34.559 10.836 34.561 13.272 ;
  LAYER M1 ;
        RECT 34.639 10.836 34.641 13.272 ;
  LAYER M1 ;
        RECT 34.719 10.836 34.721 13.272 ;
  LAYER M1 ;
        RECT 34.799 10.836 34.801 13.272 ;
  LAYER M1 ;
        RECT 34.879 10.836 34.881 13.272 ;
  LAYER M1 ;
        RECT 34.959 10.836 34.961 13.272 ;
  LAYER M1 ;
        RECT 35.039 10.836 35.041 13.272 ;
  LAYER M1 ;
        RECT 35.119 10.836 35.121 13.272 ;
  LAYER M1 ;
        RECT 35.199 10.836 35.201 13.272 ;
  LAYER M1 ;
        RECT 35.279 10.836 35.281 13.272 ;
  LAYER M1 ;
        RECT 35.359 10.836 35.361 13.272 ;
  LAYER M1 ;
        RECT 35.439 10.836 35.441 13.272 ;
  LAYER M1 ;
        RECT 35.519 10.836 35.521 13.272 ;
  LAYER M1 ;
        RECT 35.599 10.836 35.601 13.272 ;
  LAYER M1 ;
        RECT 35.679 10.836 35.681 13.272 ;
  LAYER M1 ;
        RECT 35.759 10.836 35.761 13.272 ;
  LAYER M1 ;
        RECT 35.839 10.836 35.841 13.272 ;
  LAYER M1 ;
        RECT 35.919 10.836 35.921 13.272 ;
  LAYER M1 ;
        RECT 35.999 10.836 36.001 13.272 ;
  LAYER M1 ;
        RECT 36.079 10.836 36.081 13.272 ;
  LAYER M1 ;
        RECT 36.159 10.836 36.161 13.272 ;
  LAYER M1 ;
        RECT 36.239 10.836 36.241 13.272 ;
  LAYER M1 ;
        RECT 36.319 10.836 36.321 13.272 ;
  LAYER M1 ;
        RECT 36.399 10.836 36.401 13.272 ;
  LAYER M1 ;
        RECT 36.479 10.836 36.481 13.272 ;
  LAYER M1 ;
        RECT 36.559 10.836 36.561 13.272 ;
  LAYER M1 ;
        RECT 36.639 10.836 36.641 13.272 ;
  LAYER M1 ;
        RECT 36.719 10.836 36.721 13.272 ;
  LAYER M1 ;
        RECT 36.799 10.836 36.801 13.272 ;
  LAYER M2 ;
        RECT 34.48 13.271 36.88 13.273 ;
  LAYER M2 ;
        RECT 34.48 13.187 36.88 13.189 ;
  LAYER M2 ;
        RECT 34.48 13.103 36.88 13.105 ;
  LAYER M2 ;
        RECT 34.48 13.019 36.88 13.021 ;
  LAYER M2 ;
        RECT 34.48 12.935 36.88 12.937 ;
  LAYER M2 ;
        RECT 34.48 12.851 36.88 12.853 ;
  LAYER M2 ;
        RECT 34.48 12.767 36.88 12.769 ;
  LAYER M2 ;
        RECT 34.48 12.683 36.88 12.685 ;
  LAYER M2 ;
        RECT 34.48 12.599 36.88 12.601 ;
  LAYER M2 ;
        RECT 34.48 12.515 36.88 12.517 ;
  LAYER M2 ;
        RECT 34.48 12.431 36.88 12.433 ;
  LAYER M2 ;
        RECT 34.48 12.347 36.88 12.349 ;
  LAYER M2 ;
        RECT 34.48 12.2635 36.88 12.2655 ;
  LAYER M2 ;
        RECT 34.48 12.179 36.88 12.181 ;
  LAYER M2 ;
        RECT 34.48 12.095 36.88 12.097 ;
  LAYER M2 ;
        RECT 34.48 12.011 36.88 12.013 ;
  LAYER M2 ;
        RECT 34.48 11.927 36.88 11.929 ;
  LAYER M2 ;
        RECT 34.48 11.843 36.88 11.845 ;
  LAYER M2 ;
        RECT 34.48 11.759 36.88 11.761 ;
  LAYER M2 ;
        RECT 34.48 11.675 36.88 11.677 ;
  LAYER M2 ;
        RECT 34.48 11.591 36.88 11.593 ;
  LAYER M2 ;
        RECT 34.48 11.507 36.88 11.509 ;
  LAYER M2 ;
        RECT 34.48 11.423 36.88 11.425 ;
  LAYER M2 ;
        RECT 34.48 11.339 36.88 11.341 ;
  LAYER M2 ;
        RECT 34.48 11.255 36.88 11.257 ;
  LAYER M2 ;
        RECT 34.48 11.171 36.88 11.173 ;
  LAYER M2 ;
        RECT 34.48 11.087 36.88 11.089 ;
  LAYER M2 ;
        RECT 34.48 11.003 36.88 11.005 ;
  LAYER M2 ;
        RECT 34.48 10.919 36.88 10.921 ;
  LAYER M1 ;
        RECT 34.464 7.86 34.496 10.368 ;
  LAYER M1 ;
        RECT 34.528 7.86 34.56 10.368 ;
  LAYER M1 ;
        RECT 34.592 7.86 34.624 10.368 ;
  LAYER M1 ;
        RECT 34.656 7.86 34.688 10.368 ;
  LAYER M1 ;
        RECT 34.72 7.86 34.752 10.368 ;
  LAYER M1 ;
        RECT 34.784 7.86 34.816 10.368 ;
  LAYER M1 ;
        RECT 34.848 7.86 34.88 10.368 ;
  LAYER M1 ;
        RECT 34.912 7.86 34.944 10.368 ;
  LAYER M1 ;
        RECT 34.976 7.86 35.008 10.368 ;
  LAYER M1 ;
        RECT 35.04 7.86 35.072 10.368 ;
  LAYER M1 ;
        RECT 35.104 7.86 35.136 10.368 ;
  LAYER M1 ;
        RECT 35.168 7.86 35.2 10.368 ;
  LAYER M1 ;
        RECT 35.232 7.86 35.264 10.368 ;
  LAYER M1 ;
        RECT 35.296 7.86 35.328 10.368 ;
  LAYER M1 ;
        RECT 35.36 7.86 35.392 10.368 ;
  LAYER M1 ;
        RECT 35.424 7.86 35.456 10.368 ;
  LAYER M1 ;
        RECT 35.488 7.86 35.52 10.368 ;
  LAYER M1 ;
        RECT 35.552 7.86 35.584 10.368 ;
  LAYER M1 ;
        RECT 35.616 7.86 35.648 10.368 ;
  LAYER M1 ;
        RECT 35.68 7.86 35.712 10.368 ;
  LAYER M1 ;
        RECT 35.744 7.86 35.776 10.368 ;
  LAYER M1 ;
        RECT 35.808 7.86 35.84 10.368 ;
  LAYER M1 ;
        RECT 35.872 7.86 35.904 10.368 ;
  LAYER M1 ;
        RECT 35.936 7.86 35.968 10.368 ;
  LAYER M1 ;
        RECT 36 7.86 36.032 10.368 ;
  LAYER M1 ;
        RECT 36.064 7.86 36.096 10.368 ;
  LAYER M1 ;
        RECT 36.128 7.86 36.16 10.368 ;
  LAYER M1 ;
        RECT 36.192 7.86 36.224 10.368 ;
  LAYER M1 ;
        RECT 36.256 7.86 36.288 10.368 ;
  LAYER M1 ;
        RECT 36.32 7.86 36.352 10.368 ;
  LAYER M1 ;
        RECT 36.384 7.86 36.416 10.368 ;
  LAYER M1 ;
        RECT 36.448 7.86 36.48 10.368 ;
  LAYER M1 ;
        RECT 36.512 7.86 36.544 10.368 ;
  LAYER M1 ;
        RECT 36.576 7.86 36.608 10.368 ;
  LAYER M1 ;
        RECT 36.64 7.86 36.672 10.368 ;
  LAYER M1 ;
        RECT 36.704 7.86 36.736 10.368 ;
  LAYER M1 ;
        RECT 36.768 7.86 36.8 10.368 ;
  LAYER M2 ;
        RECT 34.444 10.252 36.916 10.284 ;
  LAYER M2 ;
        RECT 34.444 10.188 36.916 10.22 ;
  LAYER M2 ;
        RECT 34.444 10.124 36.916 10.156 ;
  LAYER M2 ;
        RECT 34.444 10.06 36.916 10.092 ;
  LAYER M2 ;
        RECT 34.444 9.996 36.916 10.028 ;
  LAYER M2 ;
        RECT 34.444 9.932 36.916 9.964 ;
  LAYER M2 ;
        RECT 34.444 9.868 36.916 9.9 ;
  LAYER M2 ;
        RECT 34.444 9.804 36.916 9.836 ;
  LAYER M2 ;
        RECT 34.444 9.74 36.916 9.772 ;
  LAYER M2 ;
        RECT 34.444 9.676 36.916 9.708 ;
  LAYER M2 ;
        RECT 34.444 9.612 36.916 9.644 ;
  LAYER M2 ;
        RECT 34.444 9.548 36.916 9.58 ;
  LAYER M2 ;
        RECT 34.444 9.484 36.916 9.516 ;
  LAYER M2 ;
        RECT 34.444 9.42 36.916 9.452 ;
  LAYER M2 ;
        RECT 34.444 9.356 36.916 9.388 ;
  LAYER M2 ;
        RECT 34.444 9.292 36.916 9.324 ;
  LAYER M2 ;
        RECT 34.444 9.228 36.916 9.26 ;
  LAYER M2 ;
        RECT 34.444 9.164 36.916 9.196 ;
  LAYER M2 ;
        RECT 34.444 9.1 36.916 9.132 ;
  LAYER M2 ;
        RECT 34.444 9.036 36.916 9.068 ;
  LAYER M2 ;
        RECT 34.444 8.972 36.916 9.004 ;
  LAYER M2 ;
        RECT 34.444 8.908 36.916 8.94 ;
  LAYER M2 ;
        RECT 34.444 8.844 36.916 8.876 ;
  LAYER M2 ;
        RECT 34.444 8.78 36.916 8.812 ;
  LAYER M2 ;
        RECT 34.444 8.716 36.916 8.748 ;
  LAYER M2 ;
        RECT 34.444 8.652 36.916 8.684 ;
  LAYER M2 ;
        RECT 34.444 8.588 36.916 8.62 ;
  LAYER M2 ;
        RECT 34.444 8.524 36.916 8.556 ;
  LAYER M2 ;
        RECT 34.444 8.46 36.916 8.492 ;
  LAYER M2 ;
        RECT 34.444 8.396 36.916 8.428 ;
  LAYER M2 ;
        RECT 34.444 8.332 36.916 8.364 ;
  LAYER M2 ;
        RECT 34.444 8.268 36.916 8.3 ;
  LAYER M2 ;
        RECT 34.444 8.204 36.916 8.236 ;
  LAYER M2 ;
        RECT 34.444 8.14 36.916 8.172 ;
  LAYER M2 ;
        RECT 34.444 8.076 36.916 8.108 ;
  LAYER M2 ;
        RECT 34.444 8.012 36.916 8.044 ;
  LAYER M3 ;
        RECT 34.464 7.86 34.496 10.368 ;
  LAYER M3 ;
        RECT 34.528 7.86 34.56 10.368 ;
  LAYER M3 ;
        RECT 34.592 7.86 34.624 10.368 ;
  LAYER M3 ;
        RECT 34.656 7.86 34.688 10.368 ;
  LAYER M3 ;
        RECT 34.72 7.86 34.752 10.368 ;
  LAYER M3 ;
        RECT 34.784 7.86 34.816 10.368 ;
  LAYER M3 ;
        RECT 34.848 7.86 34.88 10.368 ;
  LAYER M3 ;
        RECT 34.912 7.86 34.944 10.368 ;
  LAYER M3 ;
        RECT 34.976 7.86 35.008 10.368 ;
  LAYER M3 ;
        RECT 35.04 7.86 35.072 10.368 ;
  LAYER M3 ;
        RECT 35.104 7.86 35.136 10.368 ;
  LAYER M3 ;
        RECT 35.168 7.86 35.2 10.368 ;
  LAYER M3 ;
        RECT 35.232 7.86 35.264 10.368 ;
  LAYER M3 ;
        RECT 35.296 7.86 35.328 10.368 ;
  LAYER M3 ;
        RECT 35.36 7.86 35.392 10.368 ;
  LAYER M3 ;
        RECT 35.424 7.86 35.456 10.368 ;
  LAYER M3 ;
        RECT 35.488 7.86 35.52 10.368 ;
  LAYER M3 ;
        RECT 35.552 7.86 35.584 10.368 ;
  LAYER M3 ;
        RECT 35.616 7.86 35.648 10.368 ;
  LAYER M3 ;
        RECT 35.68 7.86 35.712 10.368 ;
  LAYER M3 ;
        RECT 35.744 7.86 35.776 10.368 ;
  LAYER M3 ;
        RECT 35.808 7.86 35.84 10.368 ;
  LAYER M3 ;
        RECT 35.872 7.86 35.904 10.368 ;
  LAYER M3 ;
        RECT 35.936 7.86 35.968 10.368 ;
  LAYER M3 ;
        RECT 36 7.86 36.032 10.368 ;
  LAYER M3 ;
        RECT 36.064 7.86 36.096 10.368 ;
  LAYER M3 ;
        RECT 36.128 7.86 36.16 10.368 ;
  LAYER M3 ;
        RECT 36.192 7.86 36.224 10.368 ;
  LAYER M3 ;
        RECT 36.256 7.86 36.288 10.368 ;
  LAYER M3 ;
        RECT 36.32 7.86 36.352 10.368 ;
  LAYER M3 ;
        RECT 36.384 7.86 36.416 10.368 ;
  LAYER M3 ;
        RECT 36.448 7.86 36.48 10.368 ;
  LAYER M3 ;
        RECT 36.512 7.86 36.544 10.368 ;
  LAYER M3 ;
        RECT 36.576 7.86 36.608 10.368 ;
  LAYER M3 ;
        RECT 36.64 7.86 36.672 10.368 ;
  LAYER M3 ;
        RECT 36.704 7.86 36.736 10.368 ;
  LAYER M3 ;
        RECT 36.768 7.86 36.8 10.368 ;
  LAYER M3 ;
        RECT 36.864 7.86 36.896 10.368 ;
  LAYER M1 ;
        RECT 34.479 7.896 34.481 10.332 ;
  LAYER M1 ;
        RECT 34.559 7.896 34.561 10.332 ;
  LAYER M1 ;
        RECT 34.639 7.896 34.641 10.332 ;
  LAYER M1 ;
        RECT 34.719 7.896 34.721 10.332 ;
  LAYER M1 ;
        RECT 34.799 7.896 34.801 10.332 ;
  LAYER M1 ;
        RECT 34.879 7.896 34.881 10.332 ;
  LAYER M1 ;
        RECT 34.959 7.896 34.961 10.332 ;
  LAYER M1 ;
        RECT 35.039 7.896 35.041 10.332 ;
  LAYER M1 ;
        RECT 35.119 7.896 35.121 10.332 ;
  LAYER M1 ;
        RECT 35.199 7.896 35.201 10.332 ;
  LAYER M1 ;
        RECT 35.279 7.896 35.281 10.332 ;
  LAYER M1 ;
        RECT 35.359 7.896 35.361 10.332 ;
  LAYER M1 ;
        RECT 35.439 7.896 35.441 10.332 ;
  LAYER M1 ;
        RECT 35.519 7.896 35.521 10.332 ;
  LAYER M1 ;
        RECT 35.599 7.896 35.601 10.332 ;
  LAYER M1 ;
        RECT 35.679 7.896 35.681 10.332 ;
  LAYER M1 ;
        RECT 35.759 7.896 35.761 10.332 ;
  LAYER M1 ;
        RECT 35.839 7.896 35.841 10.332 ;
  LAYER M1 ;
        RECT 35.919 7.896 35.921 10.332 ;
  LAYER M1 ;
        RECT 35.999 7.896 36.001 10.332 ;
  LAYER M1 ;
        RECT 36.079 7.896 36.081 10.332 ;
  LAYER M1 ;
        RECT 36.159 7.896 36.161 10.332 ;
  LAYER M1 ;
        RECT 36.239 7.896 36.241 10.332 ;
  LAYER M1 ;
        RECT 36.319 7.896 36.321 10.332 ;
  LAYER M1 ;
        RECT 36.399 7.896 36.401 10.332 ;
  LAYER M1 ;
        RECT 36.479 7.896 36.481 10.332 ;
  LAYER M1 ;
        RECT 36.559 7.896 36.561 10.332 ;
  LAYER M1 ;
        RECT 36.639 7.896 36.641 10.332 ;
  LAYER M1 ;
        RECT 36.719 7.896 36.721 10.332 ;
  LAYER M1 ;
        RECT 36.799 7.896 36.801 10.332 ;
  LAYER M2 ;
        RECT 34.48 10.331 36.88 10.333 ;
  LAYER M2 ;
        RECT 34.48 10.247 36.88 10.249 ;
  LAYER M2 ;
        RECT 34.48 10.163 36.88 10.165 ;
  LAYER M2 ;
        RECT 34.48 10.079 36.88 10.081 ;
  LAYER M2 ;
        RECT 34.48 9.995 36.88 9.997 ;
  LAYER M2 ;
        RECT 34.48 9.911 36.88 9.913 ;
  LAYER M2 ;
        RECT 34.48 9.827 36.88 9.829 ;
  LAYER M2 ;
        RECT 34.48 9.743 36.88 9.745 ;
  LAYER M2 ;
        RECT 34.48 9.659 36.88 9.661 ;
  LAYER M2 ;
        RECT 34.48 9.575 36.88 9.577 ;
  LAYER M2 ;
        RECT 34.48 9.491 36.88 9.493 ;
  LAYER M2 ;
        RECT 34.48 9.407 36.88 9.409 ;
  LAYER M2 ;
        RECT 34.48 9.3235 36.88 9.3255 ;
  LAYER M2 ;
        RECT 34.48 9.239 36.88 9.241 ;
  LAYER M2 ;
        RECT 34.48 9.155 36.88 9.157 ;
  LAYER M2 ;
        RECT 34.48 9.071 36.88 9.073 ;
  LAYER M2 ;
        RECT 34.48 8.987 36.88 8.989 ;
  LAYER M2 ;
        RECT 34.48 8.903 36.88 8.905 ;
  LAYER M2 ;
        RECT 34.48 8.819 36.88 8.821 ;
  LAYER M2 ;
        RECT 34.48 8.735 36.88 8.737 ;
  LAYER M2 ;
        RECT 34.48 8.651 36.88 8.653 ;
  LAYER M2 ;
        RECT 34.48 8.567 36.88 8.569 ;
  LAYER M2 ;
        RECT 34.48 8.483 36.88 8.485 ;
  LAYER M2 ;
        RECT 34.48 8.399 36.88 8.401 ;
  LAYER M2 ;
        RECT 34.48 8.315 36.88 8.317 ;
  LAYER M2 ;
        RECT 34.48 8.231 36.88 8.233 ;
  LAYER M2 ;
        RECT 34.48 8.147 36.88 8.149 ;
  LAYER M2 ;
        RECT 34.48 8.063 36.88 8.065 ;
  LAYER M2 ;
        RECT 34.48 7.979 36.88 7.981 ;
  LAYER M1 ;
        RECT 34.464 4.92 34.496 7.428 ;
  LAYER M1 ;
        RECT 34.528 4.92 34.56 7.428 ;
  LAYER M1 ;
        RECT 34.592 4.92 34.624 7.428 ;
  LAYER M1 ;
        RECT 34.656 4.92 34.688 7.428 ;
  LAYER M1 ;
        RECT 34.72 4.92 34.752 7.428 ;
  LAYER M1 ;
        RECT 34.784 4.92 34.816 7.428 ;
  LAYER M1 ;
        RECT 34.848 4.92 34.88 7.428 ;
  LAYER M1 ;
        RECT 34.912 4.92 34.944 7.428 ;
  LAYER M1 ;
        RECT 34.976 4.92 35.008 7.428 ;
  LAYER M1 ;
        RECT 35.04 4.92 35.072 7.428 ;
  LAYER M1 ;
        RECT 35.104 4.92 35.136 7.428 ;
  LAYER M1 ;
        RECT 35.168 4.92 35.2 7.428 ;
  LAYER M1 ;
        RECT 35.232 4.92 35.264 7.428 ;
  LAYER M1 ;
        RECT 35.296 4.92 35.328 7.428 ;
  LAYER M1 ;
        RECT 35.36 4.92 35.392 7.428 ;
  LAYER M1 ;
        RECT 35.424 4.92 35.456 7.428 ;
  LAYER M1 ;
        RECT 35.488 4.92 35.52 7.428 ;
  LAYER M1 ;
        RECT 35.552 4.92 35.584 7.428 ;
  LAYER M1 ;
        RECT 35.616 4.92 35.648 7.428 ;
  LAYER M1 ;
        RECT 35.68 4.92 35.712 7.428 ;
  LAYER M1 ;
        RECT 35.744 4.92 35.776 7.428 ;
  LAYER M1 ;
        RECT 35.808 4.92 35.84 7.428 ;
  LAYER M1 ;
        RECT 35.872 4.92 35.904 7.428 ;
  LAYER M1 ;
        RECT 35.936 4.92 35.968 7.428 ;
  LAYER M1 ;
        RECT 36 4.92 36.032 7.428 ;
  LAYER M1 ;
        RECT 36.064 4.92 36.096 7.428 ;
  LAYER M1 ;
        RECT 36.128 4.92 36.16 7.428 ;
  LAYER M1 ;
        RECT 36.192 4.92 36.224 7.428 ;
  LAYER M1 ;
        RECT 36.256 4.92 36.288 7.428 ;
  LAYER M1 ;
        RECT 36.32 4.92 36.352 7.428 ;
  LAYER M1 ;
        RECT 36.384 4.92 36.416 7.428 ;
  LAYER M1 ;
        RECT 36.448 4.92 36.48 7.428 ;
  LAYER M1 ;
        RECT 36.512 4.92 36.544 7.428 ;
  LAYER M1 ;
        RECT 36.576 4.92 36.608 7.428 ;
  LAYER M1 ;
        RECT 36.64 4.92 36.672 7.428 ;
  LAYER M1 ;
        RECT 36.704 4.92 36.736 7.428 ;
  LAYER M1 ;
        RECT 36.768 4.92 36.8 7.428 ;
  LAYER M2 ;
        RECT 34.444 7.312 36.916 7.344 ;
  LAYER M2 ;
        RECT 34.444 7.248 36.916 7.28 ;
  LAYER M2 ;
        RECT 34.444 7.184 36.916 7.216 ;
  LAYER M2 ;
        RECT 34.444 7.12 36.916 7.152 ;
  LAYER M2 ;
        RECT 34.444 7.056 36.916 7.088 ;
  LAYER M2 ;
        RECT 34.444 6.992 36.916 7.024 ;
  LAYER M2 ;
        RECT 34.444 6.928 36.916 6.96 ;
  LAYER M2 ;
        RECT 34.444 6.864 36.916 6.896 ;
  LAYER M2 ;
        RECT 34.444 6.8 36.916 6.832 ;
  LAYER M2 ;
        RECT 34.444 6.736 36.916 6.768 ;
  LAYER M2 ;
        RECT 34.444 6.672 36.916 6.704 ;
  LAYER M2 ;
        RECT 34.444 6.608 36.916 6.64 ;
  LAYER M2 ;
        RECT 34.444 6.544 36.916 6.576 ;
  LAYER M2 ;
        RECT 34.444 6.48 36.916 6.512 ;
  LAYER M2 ;
        RECT 34.444 6.416 36.916 6.448 ;
  LAYER M2 ;
        RECT 34.444 6.352 36.916 6.384 ;
  LAYER M2 ;
        RECT 34.444 6.288 36.916 6.32 ;
  LAYER M2 ;
        RECT 34.444 6.224 36.916 6.256 ;
  LAYER M2 ;
        RECT 34.444 6.16 36.916 6.192 ;
  LAYER M2 ;
        RECT 34.444 6.096 36.916 6.128 ;
  LAYER M2 ;
        RECT 34.444 6.032 36.916 6.064 ;
  LAYER M2 ;
        RECT 34.444 5.968 36.916 6 ;
  LAYER M2 ;
        RECT 34.444 5.904 36.916 5.936 ;
  LAYER M2 ;
        RECT 34.444 5.84 36.916 5.872 ;
  LAYER M2 ;
        RECT 34.444 5.776 36.916 5.808 ;
  LAYER M2 ;
        RECT 34.444 5.712 36.916 5.744 ;
  LAYER M2 ;
        RECT 34.444 5.648 36.916 5.68 ;
  LAYER M2 ;
        RECT 34.444 5.584 36.916 5.616 ;
  LAYER M2 ;
        RECT 34.444 5.52 36.916 5.552 ;
  LAYER M2 ;
        RECT 34.444 5.456 36.916 5.488 ;
  LAYER M2 ;
        RECT 34.444 5.392 36.916 5.424 ;
  LAYER M2 ;
        RECT 34.444 5.328 36.916 5.36 ;
  LAYER M2 ;
        RECT 34.444 5.264 36.916 5.296 ;
  LAYER M2 ;
        RECT 34.444 5.2 36.916 5.232 ;
  LAYER M2 ;
        RECT 34.444 5.136 36.916 5.168 ;
  LAYER M2 ;
        RECT 34.444 5.072 36.916 5.104 ;
  LAYER M3 ;
        RECT 34.464 4.92 34.496 7.428 ;
  LAYER M3 ;
        RECT 34.528 4.92 34.56 7.428 ;
  LAYER M3 ;
        RECT 34.592 4.92 34.624 7.428 ;
  LAYER M3 ;
        RECT 34.656 4.92 34.688 7.428 ;
  LAYER M3 ;
        RECT 34.72 4.92 34.752 7.428 ;
  LAYER M3 ;
        RECT 34.784 4.92 34.816 7.428 ;
  LAYER M3 ;
        RECT 34.848 4.92 34.88 7.428 ;
  LAYER M3 ;
        RECT 34.912 4.92 34.944 7.428 ;
  LAYER M3 ;
        RECT 34.976 4.92 35.008 7.428 ;
  LAYER M3 ;
        RECT 35.04 4.92 35.072 7.428 ;
  LAYER M3 ;
        RECT 35.104 4.92 35.136 7.428 ;
  LAYER M3 ;
        RECT 35.168 4.92 35.2 7.428 ;
  LAYER M3 ;
        RECT 35.232 4.92 35.264 7.428 ;
  LAYER M3 ;
        RECT 35.296 4.92 35.328 7.428 ;
  LAYER M3 ;
        RECT 35.36 4.92 35.392 7.428 ;
  LAYER M3 ;
        RECT 35.424 4.92 35.456 7.428 ;
  LAYER M3 ;
        RECT 35.488 4.92 35.52 7.428 ;
  LAYER M3 ;
        RECT 35.552 4.92 35.584 7.428 ;
  LAYER M3 ;
        RECT 35.616 4.92 35.648 7.428 ;
  LAYER M3 ;
        RECT 35.68 4.92 35.712 7.428 ;
  LAYER M3 ;
        RECT 35.744 4.92 35.776 7.428 ;
  LAYER M3 ;
        RECT 35.808 4.92 35.84 7.428 ;
  LAYER M3 ;
        RECT 35.872 4.92 35.904 7.428 ;
  LAYER M3 ;
        RECT 35.936 4.92 35.968 7.428 ;
  LAYER M3 ;
        RECT 36 4.92 36.032 7.428 ;
  LAYER M3 ;
        RECT 36.064 4.92 36.096 7.428 ;
  LAYER M3 ;
        RECT 36.128 4.92 36.16 7.428 ;
  LAYER M3 ;
        RECT 36.192 4.92 36.224 7.428 ;
  LAYER M3 ;
        RECT 36.256 4.92 36.288 7.428 ;
  LAYER M3 ;
        RECT 36.32 4.92 36.352 7.428 ;
  LAYER M3 ;
        RECT 36.384 4.92 36.416 7.428 ;
  LAYER M3 ;
        RECT 36.448 4.92 36.48 7.428 ;
  LAYER M3 ;
        RECT 36.512 4.92 36.544 7.428 ;
  LAYER M3 ;
        RECT 36.576 4.92 36.608 7.428 ;
  LAYER M3 ;
        RECT 36.64 4.92 36.672 7.428 ;
  LAYER M3 ;
        RECT 36.704 4.92 36.736 7.428 ;
  LAYER M3 ;
        RECT 36.768 4.92 36.8 7.428 ;
  LAYER M3 ;
        RECT 36.864 4.92 36.896 7.428 ;
  LAYER M1 ;
        RECT 34.479 4.956 34.481 7.392 ;
  LAYER M1 ;
        RECT 34.559 4.956 34.561 7.392 ;
  LAYER M1 ;
        RECT 34.639 4.956 34.641 7.392 ;
  LAYER M1 ;
        RECT 34.719 4.956 34.721 7.392 ;
  LAYER M1 ;
        RECT 34.799 4.956 34.801 7.392 ;
  LAYER M1 ;
        RECT 34.879 4.956 34.881 7.392 ;
  LAYER M1 ;
        RECT 34.959 4.956 34.961 7.392 ;
  LAYER M1 ;
        RECT 35.039 4.956 35.041 7.392 ;
  LAYER M1 ;
        RECT 35.119 4.956 35.121 7.392 ;
  LAYER M1 ;
        RECT 35.199 4.956 35.201 7.392 ;
  LAYER M1 ;
        RECT 35.279 4.956 35.281 7.392 ;
  LAYER M1 ;
        RECT 35.359 4.956 35.361 7.392 ;
  LAYER M1 ;
        RECT 35.439 4.956 35.441 7.392 ;
  LAYER M1 ;
        RECT 35.519 4.956 35.521 7.392 ;
  LAYER M1 ;
        RECT 35.599 4.956 35.601 7.392 ;
  LAYER M1 ;
        RECT 35.679 4.956 35.681 7.392 ;
  LAYER M1 ;
        RECT 35.759 4.956 35.761 7.392 ;
  LAYER M1 ;
        RECT 35.839 4.956 35.841 7.392 ;
  LAYER M1 ;
        RECT 35.919 4.956 35.921 7.392 ;
  LAYER M1 ;
        RECT 35.999 4.956 36.001 7.392 ;
  LAYER M1 ;
        RECT 36.079 4.956 36.081 7.392 ;
  LAYER M1 ;
        RECT 36.159 4.956 36.161 7.392 ;
  LAYER M1 ;
        RECT 36.239 4.956 36.241 7.392 ;
  LAYER M1 ;
        RECT 36.319 4.956 36.321 7.392 ;
  LAYER M1 ;
        RECT 36.399 4.956 36.401 7.392 ;
  LAYER M1 ;
        RECT 36.479 4.956 36.481 7.392 ;
  LAYER M1 ;
        RECT 36.559 4.956 36.561 7.392 ;
  LAYER M1 ;
        RECT 36.639 4.956 36.641 7.392 ;
  LAYER M1 ;
        RECT 36.719 4.956 36.721 7.392 ;
  LAYER M1 ;
        RECT 36.799 4.956 36.801 7.392 ;
  LAYER M2 ;
        RECT 34.48 7.391 36.88 7.393 ;
  LAYER M2 ;
        RECT 34.48 7.307 36.88 7.309 ;
  LAYER M2 ;
        RECT 34.48 7.223 36.88 7.225 ;
  LAYER M2 ;
        RECT 34.48 7.139 36.88 7.141 ;
  LAYER M2 ;
        RECT 34.48 7.055 36.88 7.057 ;
  LAYER M2 ;
        RECT 34.48 6.971 36.88 6.973 ;
  LAYER M2 ;
        RECT 34.48 6.887 36.88 6.889 ;
  LAYER M2 ;
        RECT 34.48 6.803 36.88 6.805 ;
  LAYER M2 ;
        RECT 34.48 6.719 36.88 6.721 ;
  LAYER M2 ;
        RECT 34.48 6.635 36.88 6.637 ;
  LAYER M2 ;
        RECT 34.48 6.551 36.88 6.553 ;
  LAYER M2 ;
        RECT 34.48 6.467 36.88 6.469 ;
  LAYER M2 ;
        RECT 34.48 6.3835 36.88 6.3855 ;
  LAYER M2 ;
        RECT 34.48 6.299 36.88 6.301 ;
  LAYER M2 ;
        RECT 34.48 6.215 36.88 6.217 ;
  LAYER M2 ;
        RECT 34.48 6.131 36.88 6.133 ;
  LAYER M2 ;
        RECT 34.48 6.047 36.88 6.049 ;
  LAYER M2 ;
        RECT 34.48 5.963 36.88 5.965 ;
  LAYER M2 ;
        RECT 34.48 5.879 36.88 5.881 ;
  LAYER M2 ;
        RECT 34.48 5.795 36.88 5.797 ;
  LAYER M2 ;
        RECT 34.48 5.711 36.88 5.713 ;
  LAYER M2 ;
        RECT 34.48 5.627 36.88 5.629 ;
  LAYER M2 ;
        RECT 34.48 5.543 36.88 5.545 ;
  LAYER M2 ;
        RECT 34.48 5.459 36.88 5.461 ;
  LAYER M2 ;
        RECT 34.48 5.375 36.88 5.377 ;
  LAYER M2 ;
        RECT 34.48 5.291 36.88 5.293 ;
  LAYER M2 ;
        RECT 34.48 5.207 36.88 5.209 ;
  LAYER M2 ;
        RECT 34.48 5.123 36.88 5.125 ;
  LAYER M2 ;
        RECT 34.48 5.039 36.88 5.041 ;
  LAYER M1 ;
        RECT 34.464 1.98 34.496 4.488 ;
  LAYER M1 ;
        RECT 34.528 1.98 34.56 4.488 ;
  LAYER M1 ;
        RECT 34.592 1.98 34.624 4.488 ;
  LAYER M1 ;
        RECT 34.656 1.98 34.688 4.488 ;
  LAYER M1 ;
        RECT 34.72 1.98 34.752 4.488 ;
  LAYER M1 ;
        RECT 34.784 1.98 34.816 4.488 ;
  LAYER M1 ;
        RECT 34.848 1.98 34.88 4.488 ;
  LAYER M1 ;
        RECT 34.912 1.98 34.944 4.488 ;
  LAYER M1 ;
        RECT 34.976 1.98 35.008 4.488 ;
  LAYER M1 ;
        RECT 35.04 1.98 35.072 4.488 ;
  LAYER M1 ;
        RECT 35.104 1.98 35.136 4.488 ;
  LAYER M1 ;
        RECT 35.168 1.98 35.2 4.488 ;
  LAYER M1 ;
        RECT 35.232 1.98 35.264 4.488 ;
  LAYER M1 ;
        RECT 35.296 1.98 35.328 4.488 ;
  LAYER M1 ;
        RECT 35.36 1.98 35.392 4.488 ;
  LAYER M1 ;
        RECT 35.424 1.98 35.456 4.488 ;
  LAYER M1 ;
        RECT 35.488 1.98 35.52 4.488 ;
  LAYER M1 ;
        RECT 35.552 1.98 35.584 4.488 ;
  LAYER M1 ;
        RECT 35.616 1.98 35.648 4.488 ;
  LAYER M1 ;
        RECT 35.68 1.98 35.712 4.488 ;
  LAYER M1 ;
        RECT 35.744 1.98 35.776 4.488 ;
  LAYER M1 ;
        RECT 35.808 1.98 35.84 4.488 ;
  LAYER M1 ;
        RECT 35.872 1.98 35.904 4.488 ;
  LAYER M1 ;
        RECT 35.936 1.98 35.968 4.488 ;
  LAYER M1 ;
        RECT 36 1.98 36.032 4.488 ;
  LAYER M1 ;
        RECT 36.064 1.98 36.096 4.488 ;
  LAYER M1 ;
        RECT 36.128 1.98 36.16 4.488 ;
  LAYER M1 ;
        RECT 36.192 1.98 36.224 4.488 ;
  LAYER M1 ;
        RECT 36.256 1.98 36.288 4.488 ;
  LAYER M1 ;
        RECT 36.32 1.98 36.352 4.488 ;
  LAYER M1 ;
        RECT 36.384 1.98 36.416 4.488 ;
  LAYER M1 ;
        RECT 36.448 1.98 36.48 4.488 ;
  LAYER M1 ;
        RECT 36.512 1.98 36.544 4.488 ;
  LAYER M1 ;
        RECT 36.576 1.98 36.608 4.488 ;
  LAYER M1 ;
        RECT 36.64 1.98 36.672 4.488 ;
  LAYER M1 ;
        RECT 36.704 1.98 36.736 4.488 ;
  LAYER M1 ;
        RECT 36.768 1.98 36.8 4.488 ;
  LAYER M2 ;
        RECT 34.444 4.372 36.916 4.404 ;
  LAYER M2 ;
        RECT 34.444 4.308 36.916 4.34 ;
  LAYER M2 ;
        RECT 34.444 4.244 36.916 4.276 ;
  LAYER M2 ;
        RECT 34.444 4.18 36.916 4.212 ;
  LAYER M2 ;
        RECT 34.444 4.116 36.916 4.148 ;
  LAYER M2 ;
        RECT 34.444 4.052 36.916 4.084 ;
  LAYER M2 ;
        RECT 34.444 3.988 36.916 4.02 ;
  LAYER M2 ;
        RECT 34.444 3.924 36.916 3.956 ;
  LAYER M2 ;
        RECT 34.444 3.86 36.916 3.892 ;
  LAYER M2 ;
        RECT 34.444 3.796 36.916 3.828 ;
  LAYER M2 ;
        RECT 34.444 3.732 36.916 3.764 ;
  LAYER M2 ;
        RECT 34.444 3.668 36.916 3.7 ;
  LAYER M2 ;
        RECT 34.444 3.604 36.916 3.636 ;
  LAYER M2 ;
        RECT 34.444 3.54 36.916 3.572 ;
  LAYER M2 ;
        RECT 34.444 3.476 36.916 3.508 ;
  LAYER M2 ;
        RECT 34.444 3.412 36.916 3.444 ;
  LAYER M2 ;
        RECT 34.444 3.348 36.916 3.38 ;
  LAYER M2 ;
        RECT 34.444 3.284 36.916 3.316 ;
  LAYER M2 ;
        RECT 34.444 3.22 36.916 3.252 ;
  LAYER M2 ;
        RECT 34.444 3.156 36.916 3.188 ;
  LAYER M2 ;
        RECT 34.444 3.092 36.916 3.124 ;
  LAYER M2 ;
        RECT 34.444 3.028 36.916 3.06 ;
  LAYER M2 ;
        RECT 34.444 2.964 36.916 2.996 ;
  LAYER M2 ;
        RECT 34.444 2.9 36.916 2.932 ;
  LAYER M2 ;
        RECT 34.444 2.836 36.916 2.868 ;
  LAYER M2 ;
        RECT 34.444 2.772 36.916 2.804 ;
  LAYER M2 ;
        RECT 34.444 2.708 36.916 2.74 ;
  LAYER M2 ;
        RECT 34.444 2.644 36.916 2.676 ;
  LAYER M2 ;
        RECT 34.444 2.58 36.916 2.612 ;
  LAYER M2 ;
        RECT 34.444 2.516 36.916 2.548 ;
  LAYER M2 ;
        RECT 34.444 2.452 36.916 2.484 ;
  LAYER M2 ;
        RECT 34.444 2.388 36.916 2.42 ;
  LAYER M2 ;
        RECT 34.444 2.324 36.916 2.356 ;
  LAYER M2 ;
        RECT 34.444 2.26 36.916 2.292 ;
  LAYER M2 ;
        RECT 34.444 2.196 36.916 2.228 ;
  LAYER M2 ;
        RECT 34.444 2.132 36.916 2.164 ;
  LAYER M3 ;
        RECT 34.464 1.98 34.496 4.488 ;
  LAYER M3 ;
        RECT 34.528 1.98 34.56 4.488 ;
  LAYER M3 ;
        RECT 34.592 1.98 34.624 4.488 ;
  LAYER M3 ;
        RECT 34.656 1.98 34.688 4.488 ;
  LAYER M3 ;
        RECT 34.72 1.98 34.752 4.488 ;
  LAYER M3 ;
        RECT 34.784 1.98 34.816 4.488 ;
  LAYER M3 ;
        RECT 34.848 1.98 34.88 4.488 ;
  LAYER M3 ;
        RECT 34.912 1.98 34.944 4.488 ;
  LAYER M3 ;
        RECT 34.976 1.98 35.008 4.488 ;
  LAYER M3 ;
        RECT 35.04 1.98 35.072 4.488 ;
  LAYER M3 ;
        RECT 35.104 1.98 35.136 4.488 ;
  LAYER M3 ;
        RECT 35.168 1.98 35.2 4.488 ;
  LAYER M3 ;
        RECT 35.232 1.98 35.264 4.488 ;
  LAYER M3 ;
        RECT 35.296 1.98 35.328 4.488 ;
  LAYER M3 ;
        RECT 35.36 1.98 35.392 4.488 ;
  LAYER M3 ;
        RECT 35.424 1.98 35.456 4.488 ;
  LAYER M3 ;
        RECT 35.488 1.98 35.52 4.488 ;
  LAYER M3 ;
        RECT 35.552 1.98 35.584 4.488 ;
  LAYER M3 ;
        RECT 35.616 1.98 35.648 4.488 ;
  LAYER M3 ;
        RECT 35.68 1.98 35.712 4.488 ;
  LAYER M3 ;
        RECT 35.744 1.98 35.776 4.488 ;
  LAYER M3 ;
        RECT 35.808 1.98 35.84 4.488 ;
  LAYER M3 ;
        RECT 35.872 1.98 35.904 4.488 ;
  LAYER M3 ;
        RECT 35.936 1.98 35.968 4.488 ;
  LAYER M3 ;
        RECT 36 1.98 36.032 4.488 ;
  LAYER M3 ;
        RECT 36.064 1.98 36.096 4.488 ;
  LAYER M3 ;
        RECT 36.128 1.98 36.16 4.488 ;
  LAYER M3 ;
        RECT 36.192 1.98 36.224 4.488 ;
  LAYER M3 ;
        RECT 36.256 1.98 36.288 4.488 ;
  LAYER M3 ;
        RECT 36.32 1.98 36.352 4.488 ;
  LAYER M3 ;
        RECT 36.384 1.98 36.416 4.488 ;
  LAYER M3 ;
        RECT 36.448 1.98 36.48 4.488 ;
  LAYER M3 ;
        RECT 36.512 1.98 36.544 4.488 ;
  LAYER M3 ;
        RECT 36.576 1.98 36.608 4.488 ;
  LAYER M3 ;
        RECT 36.64 1.98 36.672 4.488 ;
  LAYER M3 ;
        RECT 36.704 1.98 36.736 4.488 ;
  LAYER M3 ;
        RECT 36.768 1.98 36.8 4.488 ;
  LAYER M3 ;
        RECT 36.864 1.98 36.896 4.488 ;
  LAYER M1 ;
        RECT 34.479 2.016 34.481 4.452 ;
  LAYER M1 ;
        RECT 34.559 2.016 34.561 4.452 ;
  LAYER M1 ;
        RECT 34.639 2.016 34.641 4.452 ;
  LAYER M1 ;
        RECT 34.719 2.016 34.721 4.452 ;
  LAYER M1 ;
        RECT 34.799 2.016 34.801 4.452 ;
  LAYER M1 ;
        RECT 34.879 2.016 34.881 4.452 ;
  LAYER M1 ;
        RECT 34.959 2.016 34.961 4.452 ;
  LAYER M1 ;
        RECT 35.039 2.016 35.041 4.452 ;
  LAYER M1 ;
        RECT 35.119 2.016 35.121 4.452 ;
  LAYER M1 ;
        RECT 35.199 2.016 35.201 4.452 ;
  LAYER M1 ;
        RECT 35.279 2.016 35.281 4.452 ;
  LAYER M1 ;
        RECT 35.359 2.016 35.361 4.452 ;
  LAYER M1 ;
        RECT 35.439 2.016 35.441 4.452 ;
  LAYER M1 ;
        RECT 35.519 2.016 35.521 4.452 ;
  LAYER M1 ;
        RECT 35.599 2.016 35.601 4.452 ;
  LAYER M1 ;
        RECT 35.679 2.016 35.681 4.452 ;
  LAYER M1 ;
        RECT 35.759 2.016 35.761 4.452 ;
  LAYER M1 ;
        RECT 35.839 2.016 35.841 4.452 ;
  LAYER M1 ;
        RECT 35.919 2.016 35.921 4.452 ;
  LAYER M1 ;
        RECT 35.999 2.016 36.001 4.452 ;
  LAYER M1 ;
        RECT 36.079 2.016 36.081 4.452 ;
  LAYER M1 ;
        RECT 36.159 2.016 36.161 4.452 ;
  LAYER M1 ;
        RECT 36.239 2.016 36.241 4.452 ;
  LAYER M1 ;
        RECT 36.319 2.016 36.321 4.452 ;
  LAYER M1 ;
        RECT 36.399 2.016 36.401 4.452 ;
  LAYER M1 ;
        RECT 36.479 2.016 36.481 4.452 ;
  LAYER M1 ;
        RECT 36.559 2.016 36.561 4.452 ;
  LAYER M1 ;
        RECT 36.639 2.016 36.641 4.452 ;
  LAYER M1 ;
        RECT 36.719 2.016 36.721 4.452 ;
  LAYER M1 ;
        RECT 36.799 2.016 36.801 4.452 ;
  LAYER M2 ;
        RECT 34.48 4.451 36.88 4.453 ;
  LAYER M2 ;
        RECT 34.48 4.367 36.88 4.369 ;
  LAYER M2 ;
        RECT 34.48 4.283 36.88 4.285 ;
  LAYER M2 ;
        RECT 34.48 4.199 36.88 4.201 ;
  LAYER M2 ;
        RECT 34.48 4.115 36.88 4.117 ;
  LAYER M2 ;
        RECT 34.48 4.031 36.88 4.033 ;
  LAYER M2 ;
        RECT 34.48 3.947 36.88 3.949 ;
  LAYER M2 ;
        RECT 34.48 3.863 36.88 3.865 ;
  LAYER M2 ;
        RECT 34.48 3.779 36.88 3.781 ;
  LAYER M2 ;
        RECT 34.48 3.695 36.88 3.697 ;
  LAYER M2 ;
        RECT 34.48 3.611 36.88 3.613 ;
  LAYER M2 ;
        RECT 34.48 3.527 36.88 3.529 ;
  LAYER M2 ;
        RECT 34.48 3.4435 36.88 3.4455 ;
  LAYER M2 ;
        RECT 34.48 3.359 36.88 3.361 ;
  LAYER M2 ;
        RECT 34.48 3.275 36.88 3.277 ;
  LAYER M2 ;
        RECT 34.48 3.191 36.88 3.193 ;
  LAYER M2 ;
        RECT 34.48 3.107 36.88 3.109 ;
  LAYER M2 ;
        RECT 34.48 3.023 36.88 3.025 ;
  LAYER M2 ;
        RECT 34.48 2.939 36.88 2.941 ;
  LAYER M2 ;
        RECT 34.48 2.855 36.88 2.857 ;
  LAYER M2 ;
        RECT 34.48 2.771 36.88 2.773 ;
  LAYER M2 ;
        RECT 34.48 2.687 36.88 2.689 ;
  LAYER M2 ;
        RECT 34.48 2.603 36.88 2.605 ;
  LAYER M2 ;
        RECT 34.48 2.519 36.88 2.521 ;
  LAYER M2 ;
        RECT 34.48 2.435 36.88 2.437 ;
  LAYER M2 ;
        RECT 34.48 2.351 36.88 2.353 ;
  LAYER M2 ;
        RECT 34.48 2.267 36.88 2.269 ;
  LAYER M2 ;
        RECT 34.48 2.183 36.88 2.185 ;
  LAYER M2 ;
        RECT 34.48 2.099 36.88 2.101 ;
  LAYER M1 ;
        RECT 37.344 13.74 37.376 16.248 ;
  LAYER M1 ;
        RECT 37.408 13.74 37.44 16.248 ;
  LAYER M1 ;
        RECT 37.472 13.74 37.504 16.248 ;
  LAYER M1 ;
        RECT 37.536 13.74 37.568 16.248 ;
  LAYER M1 ;
        RECT 37.6 13.74 37.632 16.248 ;
  LAYER M1 ;
        RECT 37.664 13.74 37.696 16.248 ;
  LAYER M1 ;
        RECT 37.728 13.74 37.76 16.248 ;
  LAYER M1 ;
        RECT 37.792 13.74 37.824 16.248 ;
  LAYER M1 ;
        RECT 37.856 13.74 37.888 16.248 ;
  LAYER M1 ;
        RECT 37.92 13.74 37.952 16.248 ;
  LAYER M1 ;
        RECT 37.984 13.74 38.016 16.248 ;
  LAYER M1 ;
        RECT 38.048 13.74 38.08 16.248 ;
  LAYER M1 ;
        RECT 38.112 13.74 38.144 16.248 ;
  LAYER M1 ;
        RECT 38.176 13.74 38.208 16.248 ;
  LAYER M1 ;
        RECT 38.24 13.74 38.272 16.248 ;
  LAYER M1 ;
        RECT 38.304 13.74 38.336 16.248 ;
  LAYER M1 ;
        RECT 38.368 13.74 38.4 16.248 ;
  LAYER M1 ;
        RECT 38.432 13.74 38.464 16.248 ;
  LAYER M1 ;
        RECT 38.496 13.74 38.528 16.248 ;
  LAYER M1 ;
        RECT 38.56 13.74 38.592 16.248 ;
  LAYER M1 ;
        RECT 38.624 13.74 38.656 16.248 ;
  LAYER M1 ;
        RECT 38.688 13.74 38.72 16.248 ;
  LAYER M1 ;
        RECT 38.752 13.74 38.784 16.248 ;
  LAYER M1 ;
        RECT 38.816 13.74 38.848 16.248 ;
  LAYER M1 ;
        RECT 38.88 13.74 38.912 16.248 ;
  LAYER M1 ;
        RECT 38.944 13.74 38.976 16.248 ;
  LAYER M1 ;
        RECT 39.008 13.74 39.04 16.248 ;
  LAYER M1 ;
        RECT 39.072 13.74 39.104 16.248 ;
  LAYER M1 ;
        RECT 39.136 13.74 39.168 16.248 ;
  LAYER M1 ;
        RECT 39.2 13.74 39.232 16.248 ;
  LAYER M1 ;
        RECT 39.264 13.74 39.296 16.248 ;
  LAYER M1 ;
        RECT 39.328 13.74 39.36 16.248 ;
  LAYER M1 ;
        RECT 39.392 13.74 39.424 16.248 ;
  LAYER M1 ;
        RECT 39.456 13.74 39.488 16.248 ;
  LAYER M1 ;
        RECT 39.52 13.74 39.552 16.248 ;
  LAYER M1 ;
        RECT 39.584 13.74 39.616 16.248 ;
  LAYER M1 ;
        RECT 39.648 13.74 39.68 16.248 ;
  LAYER M2 ;
        RECT 37.324 16.132 39.796 16.164 ;
  LAYER M2 ;
        RECT 37.324 16.068 39.796 16.1 ;
  LAYER M2 ;
        RECT 37.324 16.004 39.796 16.036 ;
  LAYER M2 ;
        RECT 37.324 15.94 39.796 15.972 ;
  LAYER M2 ;
        RECT 37.324 15.876 39.796 15.908 ;
  LAYER M2 ;
        RECT 37.324 15.812 39.796 15.844 ;
  LAYER M2 ;
        RECT 37.324 15.748 39.796 15.78 ;
  LAYER M2 ;
        RECT 37.324 15.684 39.796 15.716 ;
  LAYER M2 ;
        RECT 37.324 15.62 39.796 15.652 ;
  LAYER M2 ;
        RECT 37.324 15.556 39.796 15.588 ;
  LAYER M2 ;
        RECT 37.324 15.492 39.796 15.524 ;
  LAYER M2 ;
        RECT 37.324 15.428 39.796 15.46 ;
  LAYER M2 ;
        RECT 37.324 15.364 39.796 15.396 ;
  LAYER M2 ;
        RECT 37.324 15.3 39.796 15.332 ;
  LAYER M2 ;
        RECT 37.324 15.236 39.796 15.268 ;
  LAYER M2 ;
        RECT 37.324 15.172 39.796 15.204 ;
  LAYER M2 ;
        RECT 37.324 15.108 39.796 15.14 ;
  LAYER M2 ;
        RECT 37.324 15.044 39.796 15.076 ;
  LAYER M2 ;
        RECT 37.324 14.98 39.796 15.012 ;
  LAYER M2 ;
        RECT 37.324 14.916 39.796 14.948 ;
  LAYER M2 ;
        RECT 37.324 14.852 39.796 14.884 ;
  LAYER M2 ;
        RECT 37.324 14.788 39.796 14.82 ;
  LAYER M2 ;
        RECT 37.324 14.724 39.796 14.756 ;
  LAYER M2 ;
        RECT 37.324 14.66 39.796 14.692 ;
  LAYER M2 ;
        RECT 37.324 14.596 39.796 14.628 ;
  LAYER M2 ;
        RECT 37.324 14.532 39.796 14.564 ;
  LAYER M2 ;
        RECT 37.324 14.468 39.796 14.5 ;
  LAYER M2 ;
        RECT 37.324 14.404 39.796 14.436 ;
  LAYER M2 ;
        RECT 37.324 14.34 39.796 14.372 ;
  LAYER M2 ;
        RECT 37.324 14.276 39.796 14.308 ;
  LAYER M2 ;
        RECT 37.324 14.212 39.796 14.244 ;
  LAYER M2 ;
        RECT 37.324 14.148 39.796 14.18 ;
  LAYER M2 ;
        RECT 37.324 14.084 39.796 14.116 ;
  LAYER M2 ;
        RECT 37.324 14.02 39.796 14.052 ;
  LAYER M2 ;
        RECT 37.324 13.956 39.796 13.988 ;
  LAYER M2 ;
        RECT 37.324 13.892 39.796 13.924 ;
  LAYER M3 ;
        RECT 37.344 13.74 37.376 16.248 ;
  LAYER M3 ;
        RECT 37.408 13.74 37.44 16.248 ;
  LAYER M3 ;
        RECT 37.472 13.74 37.504 16.248 ;
  LAYER M3 ;
        RECT 37.536 13.74 37.568 16.248 ;
  LAYER M3 ;
        RECT 37.6 13.74 37.632 16.248 ;
  LAYER M3 ;
        RECT 37.664 13.74 37.696 16.248 ;
  LAYER M3 ;
        RECT 37.728 13.74 37.76 16.248 ;
  LAYER M3 ;
        RECT 37.792 13.74 37.824 16.248 ;
  LAYER M3 ;
        RECT 37.856 13.74 37.888 16.248 ;
  LAYER M3 ;
        RECT 37.92 13.74 37.952 16.248 ;
  LAYER M3 ;
        RECT 37.984 13.74 38.016 16.248 ;
  LAYER M3 ;
        RECT 38.048 13.74 38.08 16.248 ;
  LAYER M3 ;
        RECT 38.112 13.74 38.144 16.248 ;
  LAYER M3 ;
        RECT 38.176 13.74 38.208 16.248 ;
  LAYER M3 ;
        RECT 38.24 13.74 38.272 16.248 ;
  LAYER M3 ;
        RECT 38.304 13.74 38.336 16.248 ;
  LAYER M3 ;
        RECT 38.368 13.74 38.4 16.248 ;
  LAYER M3 ;
        RECT 38.432 13.74 38.464 16.248 ;
  LAYER M3 ;
        RECT 38.496 13.74 38.528 16.248 ;
  LAYER M3 ;
        RECT 38.56 13.74 38.592 16.248 ;
  LAYER M3 ;
        RECT 38.624 13.74 38.656 16.248 ;
  LAYER M3 ;
        RECT 38.688 13.74 38.72 16.248 ;
  LAYER M3 ;
        RECT 38.752 13.74 38.784 16.248 ;
  LAYER M3 ;
        RECT 38.816 13.74 38.848 16.248 ;
  LAYER M3 ;
        RECT 38.88 13.74 38.912 16.248 ;
  LAYER M3 ;
        RECT 38.944 13.74 38.976 16.248 ;
  LAYER M3 ;
        RECT 39.008 13.74 39.04 16.248 ;
  LAYER M3 ;
        RECT 39.072 13.74 39.104 16.248 ;
  LAYER M3 ;
        RECT 39.136 13.74 39.168 16.248 ;
  LAYER M3 ;
        RECT 39.2 13.74 39.232 16.248 ;
  LAYER M3 ;
        RECT 39.264 13.74 39.296 16.248 ;
  LAYER M3 ;
        RECT 39.328 13.74 39.36 16.248 ;
  LAYER M3 ;
        RECT 39.392 13.74 39.424 16.248 ;
  LAYER M3 ;
        RECT 39.456 13.74 39.488 16.248 ;
  LAYER M3 ;
        RECT 39.52 13.74 39.552 16.248 ;
  LAYER M3 ;
        RECT 39.584 13.74 39.616 16.248 ;
  LAYER M3 ;
        RECT 39.648 13.74 39.68 16.248 ;
  LAYER M3 ;
        RECT 39.744 13.74 39.776 16.248 ;
  LAYER M1 ;
        RECT 37.359 13.776 37.361 16.212 ;
  LAYER M1 ;
        RECT 37.439 13.776 37.441 16.212 ;
  LAYER M1 ;
        RECT 37.519 13.776 37.521 16.212 ;
  LAYER M1 ;
        RECT 37.599 13.776 37.601 16.212 ;
  LAYER M1 ;
        RECT 37.679 13.776 37.681 16.212 ;
  LAYER M1 ;
        RECT 37.759 13.776 37.761 16.212 ;
  LAYER M1 ;
        RECT 37.839 13.776 37.841 16.212 ;
  LAYER M1 ;
        RECT 37.919 13.776 37.921 16.212 ;
  LAYER M1 ;
        RECT 37.999 13.776 38.001 16.212 ;
  LAYER M1 ;
        RECT 38.079 13.776 38.081 16.212 ;
  LAYER M1 ;
        RECT 38.159 13.776 38.161 16.212 ;
  LAYER M1 ;
        RECT 38.239 13.776 38.241 16.212 ;
  LAYER M1 ;
        RECT 38.319 13.776 38.321 16.212 ;
  LAYER M1 ;
        RECT 38.399 13.776 38.401 16.212 ;
  LAYER M1 ;
        RECT 38.479 13.776 38.481 16.212 ;
  LAYER M1 ;
        RECT 38.559 13.776 38.561 16.212 ;
  LAYER M1 ;
        RECT 38.639 13.776 38.641 16.212 ;
  LAYER M1 ;
        RECT 38.719 13.776 38.721 16.212 ;
  LAYER M1 ;
        RECT 38.799 13.776 38.801 16.212 ;
  LAYER M1 ;
        RECT 38.879 13.776 38.881 16.212 ;
  LAYER M1 ;
        RECT 38.959 13.776 38.961 16.212 ;
  LAYER M1 ;
        RECT 39.039 13.776 39.041 16.212 ;
  LAYER M1 ;
        RECT 39.119 13.776 39.121 16.212 ;
  LAYER M1 ;
        RECT 39.199 13.776 39.201 16.212 ;
  LAYER M1 ;
        RECT 39.279 13.776 39.281 16.212 ;
  LAYER M1 ;
        RECT 39.359 13.776 39.361 16.212 ;
  LAYER M1 ;
        RECT 39.439 13.776 39.441 16.212 ;
  LAYER M1 ;
        RECT 39.519 13.776 39.521 16.212 ;
  LAYER M1 ;
        RECT 39.599 13.776 39.601 16.212 ;
  LAYER M1 ;
        RECT 39.679 13.776 39.681 16.212 ;
  LAYER M2 ;
        RECT 37.36 16.211 39.76 16.213 ;
  LAYER M2 ;
        RECT 37.36 16.127 39.76 16.129 ;
  LAYER M2 ;
        RECT 37.36 16.043 39.76 16.045 ;
  LAYER M2 ;
        RECT 37.36 15.959 39.76 15.961 ;
  LAYER M2 ;
        RECT 37.36 15.875 39.76 15.877 ;
  LAYER M2 ;
        RECT 37.36 15.791 39.76 15.793 ;
  LAYER M2 ;
        RECT 37.36 15.707 39.76 15.709 ;
  LAYER M2 ;
        RECT 37.36 15.623 39.76 15.625 ;
  LAYER M2 ;
        RECT 37.36 15.539 39.76 15.541 ;
  LAYER M2 ;
        RECT 37.36 15.455 39.76 15.457 ;
  LAYER M2 ;
        RECT 37.36 15.371 39.76 15.373 ;
  LAYER M2 ;
        RECT 37.36 15.287 39.76 15.289 ;
  LAYER M2 ;
        RECT 37.36 15.2035 39.76 15.2055 ;
  LAYER M2 ;
        RECT 37.36 15.119 39.76 15.121 ;
  LAYER M2 ;
        RECT 37.36 15.035 39.76 15.037 ;
  LAYER M2 ;
        RECT 37.36 14.951 39.76 14.953 ;
  LAYER M2 ;
        RECT 37.36 14.867 39.76 14.869 ;
  LAYER M2 ;
        RECT 37.36 14.783 39.76 14.785 ;
  LAYER M2 ;
        RECT 37.36 14.699 39.76 14.701 ;
  LAYER M2 ;
        RECT 37.36 14.615 39.76 14.617 ;
  LAYER M2 ;
        RECT 37.36 14.531 39.76 14.533 ;
  LAYER M2 ;
        RECT 37.36 14.447 39.76 14.449 ;
  LAYER M2 ;
        RECT 37.36 14.363 39.76 14.365 ;
  LAYER M2 ;
        RECT 37.36 14.279 39.76 14.281 ;
  LAYER M2 ;
        RECT 37.36 14.195 39.76 14.197 ;
  LAYER M2 ;
        RECT 37.36 14.111 39.76 14.113 ;
  LAYER M2 ;
        RECT 37.36 14.027 39.76 14.029 ;
  LAYER M2 ;
        RECT 37.36 13.943 39.76 13.945 ;
  LAYER M2 ;
        RECT 37.36 13.859 39.76 13.861 ;
  LAYER M1 ;
        RECT 37.344 10.8 37.376 13.308 ;
  LAYER M1 ;
        RECT 37.408 10.8 37.44 13.308 ;
  LAYER M1 ;
        RECT 37.472 10.8 37.504 13.308 ;
  LAYER M1 ;
        RECT 37.536 10.8 37.568 13.308 ;
  LAYER M1 ;
        RECT 37.6 10.8 37.632 13.308 ;
  LAYER M1 ;
        RECT 37.664 10.8 37.696 13.308 ;
  LAYER M1 ;
        RECT 37.728 10.8 37.76 13.308 ;
  LAYER M1 ;
        RECT 37.792 10.8 37.824 13.308 ;
  LAYER M1 ;
        RECT 37.856 10.8 37.888 13.308 ;
  LAYER M1 ;
        RECT 37.92 10.8 37.952 13.308 ;
  LAYER M1 ;
        RECT 37.984 10.8 38.016 13.308 ;
  LAYER M1 ;
        RECT 38.048 10.8 38.08 13.308 ;
  LAYER M1 ;
        RECT 38.112 10.8 38.144 13.308 ;
  LAYER M1 ;
        RECT 38.176 10.8 38.208 13.308 ;
  LAYER M1 ;
        RECT 38.24 10.8 38.272 13.308 ;
  LAYER M1 ;
        RECT 38.304 10.8 38.336 13.308 ;
  LAYER M1 ;
        RECT 38.368 10.8 38.4 13.308 ;
  LAYER M1 ;
        RECT 38.432 10.8 38.464 13.308 ;
  LAYER M1 ;
        RECT 38.496 10.8 38.528 13.308 ;
  LAYER M1 ;
        RECT 38.56 10.8 38.592 13.308 ;
  LAYER M1 ;
        RECT 38.624 10.8 38.656 13.308 ;
  LAYER M1 ;
        RECT 38.688 10.8 38.72 13.308 ;
  LAYER M1 ;
        RECT 38.752 10.8 38.784 13.308 ;
  LAYER M1 ;
        RECT 38.816 10.8 38.848 13.308 ;
  LAYER M1 ;
        RECT 38.88 10.8 38.912 13.308 ;
  LAYER M1 ;
        RECT 38.944 10.8 38.976 13.308 ;
  LAYER M1 ;
        RECT 39.008 10.8 39.04 13.308 ;
  LAYER M1 ;
        RECT 39.072 10.8 39.104 13.308 ;
  LAYER M1 ;
        RECT 39.136 10.8 39.168 13.308 ;
  LAYER M1 ;
        RECT 39.2 10.8 39.232 13.308 ;
  LAYER M1 ;
        RECT 39.264 10.8 39.296 13.308 ;
  LAYER M1 ;
        RECT 39.328 10.8 39.36 13.308 ;
  LAYER M1 ;
        RECT 39.392 10.8 39.424 13.308 ;
  LAYER M1 ;
        RECT 39.456 10.8 39.488 13.308 ;
  LAYER M1 ;
        RECT 39.52 10.8 39.552 13.308 ;
  LAYER M1 ;
        RECT 39.584 10.8 39.616 13.308 ;
  LAYER M1 ;
        RECT 39.648 10.8 39.68 13.308 ;
  LAYER M2 ;
        RECT 37.324 13.192 39.796 13.224 ;
  LAYER M2 ;
        RECT 37.324 13.128 39.796 13.16 ;
  LAYER M2 ;
        RECT 37.324 13.064 39.796 13.096 ;
  LAYER M2 ;
        RECT 37.324 13 39.796 13.032 ;
  LAYER M2 ;
        RECT 37.324 12.936 39.796 12.968 ;
  LAYER M2 ;
        RECT 37.324 12.872 39.796 12.904 ;
  LAYER M2 ;
        RECT 37.324 12.808 39.796 12.84 ;
  LAYER M2 ;
        RECT 37.324 12.744 39.796 12.776 ;
  LAYER M2 ;
        RECT 37.324 12.68 39.796 12.712 ;
  LAYER M2 ;
        RECT 37.324 12.616 39.796 12.648 ;
  LAYER M2 ;
        RECT 37.324 12.552 39.796 12.584 ;
  LAYER M2 ;
        RECT 37.324 12.488 39.796 12.52 ;
  LAYER M2 ;
        RECT 37.324 12.424 39.796 12.456 ;
  LAYER M2 ;
        RECT 37.324 12.36 39.796 12.392 ;
  LAYER M2 ;
        RECT 37.324 12.296 39.796 12.328 ;
  LAYER M2 ;
        RECT 37.324 12.232 39.796 12.264 ;
  LAYER M2 ;
        RECT 37.324 12.168 39.796 12.2 ;
  LAYER M2 ;
        RECT 37.324 12.104 39.796 12.136 ;
  LAYER M2 ;
        RECT 37.324 12.04 39.796 12.072 ;
  LAYER M2 ;
        RECT 37.324 11.976 39.796 12.008 ;
  LAYER M2 ;
        RECT 37.324 11.912 39.796 11.944 ;
  LAYER M2 ;
        RECT 37.324 11.848 39.796 11.88 ;
  LAYER M2 ;
        RECT 37.324 11.784 39.796 11.816 ;
  LAYER M2 ;
        RECT 37.324 11.72 39.796 11.752 ;
  LAYER M2 ;
        RECT 37.324 11.656 39.796 11.688 ;
  LAYER M2 ;
        RECT 37.324 11.592 39.796 11.624 ;
  LAYER M2 ;
        RECT 37.324 11.528 39.796 11.56 ;
  LAYER M2 ;
        RECT 37.324 11.464 39.796 11.496 ;
  LAYER M2 ;
        RECT 37.324 11.4 39.796 11.432 ;
  LAYER M2 ;
        RECT 37.324 11.336 39.796 11.368 ;
  LAYER M2 ;
        RECT 37.324 11.272 39.796 11.304 ;
  LAYER M2 ;
        RECT 37.324 11.208 39.796 11.24 ;
  LAYER M2 ;
        RECT 37.324 11.144 39.796 11.176 ;
  LAYER M2 ;
        RECT 37.324 11.08 39.796 11.112 ;
  LAYER M2 ;
        RECT 37.324 11.016 39.796 11.048 ;
  LAYER M2 ;
        RECT 37.324 10.952 39.796 10.984 ;
  LAYER M3 ;
        RECT 37.344 10.8 37.376 13.308 ;
  LAYER M3 ;
        RECT 37.408 10.8 37.44 13.308 ;
  LAYER M3 ;
        RECT 37.472 10.8 37.504 13.308 ;
  LAYER M3 ;
        RECT 37.536 10.8 37.568 13.308 ;
  LAYER M3 ;
        RECT 37.6 10.8 37.632 13.308 ;
  LAYER M3 ;
        RECT 37.664 10.8 37.696 13.308 ;
  LAYER M3 ;
        RECT 37.728 10.8 37.76 13.308 ;
  LAYER M3 ;
        RECT 37.792 10.8 37.824 13.308 ;
  LAYER M3 ;
        RECT 37.856 10.8 37.888 13.308 ;
  LAYER M3 ;
        RECT 37.92 10.8 37.952 13.308 ;
  LAYER M3 ;
        RECT 37.984 10.8 38.016 13.308 ;
  LAYER M3 ;
        RECT 38.048 10.8 38.08 13.308 ;
  LAYER M3 ;
        RECT 38.112 10.8 38.144 13.308 ;
  LAYER M3 ;
        RECT 38.176 10.8 38.208 13.308 ;
  LAYER M3 ;
        RECT 38.24 10.8 38.272 13.308 ;
  LAYER M3 ;
        RECT 38.304 10.8 38.336 13.308 ;
  LAYER M3 ;
        RECT 38.368 10.8 38.4 13.308 ;
  LAYER M3 ;
        RECT 38.432 10.8 38.464 13.308 ;
  LAYER M3 ;
        RECT 38.496 10.8 38.528 13.308 ;
  LAYER M3 ;
        RECT 38.56 10.8 38.592 13.308 ;
  LAYER M3 ;
        RECT 38.624 10.8 38.656 13.308 ;
  LAYER M3 ;
        RECT 38.688 10.8 38.72 13.308 ;
  LAYER M3 ;
        RECT 38.752 10.8 38.784 13.308 ;
  LAYER M3 ;
        RECT 38.816 10.8 38.848 13.308 ;
  LAYER M3 ;
        RECT 38.88 10.8 38.912 13.308 ;
  LAYER M3 ;
        RECT 38.944 10.8 38.976 13.308 ;
  LAYER M3 ;
        RECT 39.008 10.8 39.04 13.308 ;
  LAYER M3 ;
        RECT 39.072 10.8 39.104 13.308 ;
  LAYER M3 ;
        RECT 39.136 10.8 39.168 13.308 ;
  LAYER M3 ;
        RECT 39.2 10.8 39.232 13.308 ;
  LAYER M3 ;
        RECT 39.264 10.8 39.296 13.308 ;
  LAYER M3 ;
        RECT 39.328 10.8 39.36 13.308 ;
  LAYER M3 ;
        RECT 39.392 10.8 39.424 13.308 ;
  LAYER M3 ;
        RECT 39.456 10.8 39.488 13.308 ;
  LAYER M3 ;
        RECT 39.52 10.8 39.552 13.308 ;
  LAYER M3 ;
        RECT 39.584 10.8 39.616 13.308 ;
  LAYER M3 ;
        RECT 39.648 10.8 39.68 13.308 ;
  LAYER M3 ;
        RECT 39.744 10.8 39.776 13.308 ;
  LAYER M1 ;
        RECT 37.359 10.836 37.361 13.272 ;
  LAYER M1 ;
        RECT 37.439 10.836 37.441 13.272 ;
  LAYER M1 ;
        RECT 37.519 10.836 37.521 13.272 ;
  LAYER M1 ;
        RECT 37.599 10.836 37.601 13.272 ;
  LAYER M1 ;
        RECT 37.679 10.836 37.681 13.272 ;
  LAYER M1 ;
        RECT 37.759 10.836 37.761 13.272 ;
  LAYER M1 ;
        RECT 37.839 10.836 37.841 13.272 ;
  LAYER M1 ;
        RECT 37.919 10.836 37.921 13.272 ;
  LAYER M1 ;
        RECT 37.999 10.836 38.001 13.272 ;
  LAYER M1 ;
        RECT 38.079 10.836 38.081 13.272 ;
  LAYER M1 ;
        RECT 38.159 10.836 38.161 13.272 ;
  LAYER M1 ;
        RECT 38.239 10.836 38.241 13.272 ;
  LAYER M1 ;
        RECT 38.319 10.836 38.321 13.272 ;
  LAYER M1 ;
        RECT 38.399 10.836 38.401 13.272 ;
  LAYER M1 ;
        RECT 38.479 10.836 38.481 13.272 ;
  LAYER M1 ;
        RECT 38.559 10.836 38.561 13.272 ;
  LAYER M1 ;
        RECT 38.639 10.836 38.641 13.272 ;
  LAYER M1 ;
        RECT 38.719 10.836 38.721 13.272 ;
  LAYER M1 ;
        RECT 38.799 10.836 38.801 13.272 ;
  LAYER M1 ;
        RECT 38.879 10.836 38.881 13.272 ;
  LAYER M1 ;
        RECT 38.959 10.836 38.961 13.272 ;
  LAYER M1 ;
        RECT 39.039 10.836 39.041 13.272 ;
  LAYER M1 ;
        RECT 39.119 10.836 39.121 13.272 ;
  LAYER M1 ;
        RECT 39.199 10.836 39.201 13.272 ;
  LAYER M1 ;
        RECT 39.279 10.836 39.281 13.272 ;
  LAYER M1 ;
        RECT 39.359 10.836 39.361 13.272 ;
  LAYER M1 ;
        RECT 39.439 10.836 39.441 13.272 ;
  LAYER M1 ;
        RECT 39.519 10.836 39.521 13.272 ;
  LAYER M1 ;
        RECT 39.599 10.836 39.601 13.272 ;
  LAYER M1 ;
        RECT 39.679 10.836 39.681 13.272 ;
  LAYER M2 ;
        RECT 37.36 13.271 39.76 13.273 ;
  LAYER M2 ;
        RECT 37.36 13.187 39.76 13.189 ;
  LAYER M2 ;
        RECT 37.36 13.103 39.76 13.105 ;
  LAYER M2 ;
        RECT 37.36 13.019 39.76 13.021 ;
  LAYER M2 ;
        RECT 37.36 12.935 39.76 12.937 ;
  LAYER M2 ;
        RECT 37.36 12.851 39.76 12.853 ;
  LAYER M2 ;
        RECT 37.36 12.767 39.76 12.769 ;
  LAYER M2 ;
        RECT 37.36 12.683 39.76 12.685 ;
  LAYER M2 ;
        RECT 37.36 12.599 39.76 12.601 ;
  LAYER M2 ;
        RECT 37.36 12.515 39.76 12.517 ;
  LAYER M2 ;
        RECT 37.36 12.431 39.76 12.433 ;
  LAYER M2 ;
        RECT 37.36 12.347 39.76 12.349 ;
  LAYER M2 ;
        RECT 37.36 12.2635 39.76 12.2655 ;
  LAYER M2 ;
        RECT 37.36 12.179 39.76 12.181 ;
  LAYER M2 ;
        RECT 37.36 12.095 39.76 12.097 ;
  LAYER M2 ;
        RECT 37.36 12.011 39.76 12.013 ;
  LAYER M2 ;
        RECT 37.36 11.927 39.76 11.929 ;
  LAYER M2 ;
        RECT 37.36 11.843 39.76 11.845 ;
  LAYER M2 ;
        RECT 37.36 11.759 39.76 11.761 ;
  LAYER M2 ;
        RECT 37.36 11.675 39.76 11.677 ;
  LAYER M2 ;
        RECT 37.36 11.591 39.76 11.593 ;
  LAYER M2 ;
        RECT 37.36 11.507 39.76 11.509 ;
  LAYER M2 ;
        RECT 37.36 11.423 39.76 11.425 ;
  LAYER M2 ;
        RECT 37.36 11.339 39.76 11.341 ;
  LAYER M2 ;
        RECT 37.36 11.255 39.76 11.257 ;
  LAYER M2 ;
        RECT 37.36 11.171 39.76 11.173 ;
  LAYER M2 ;
        RECT 37.36 11.087 39.76 11.089 ;
  LAYER M2 ;
        RECT 37.36 11.003 39.76 11.005 ;
  LAYER M2 ;
        RECT 37.36 10.919 39.76 10.921 ;
  LAYER M1 ;
        RECT 37.344 7.86 37.376 10.368 ;
  LAYER M1 ;
        RECT 37.408 7.86 37.44 10.368 ;
  LAYER M1 ;
        RECT 37.472 7.86 37.504 10.368 ;
  LAYER M1 ;
        RECT 37.536 7.86 37.568 10.368 ;
  LAYER M1 ;
        RECT 37.6 7.86 37.632 10.368 ;
  LAYER M1 ;
        RECT 37.664 7.86 37.696 10.368 ;
  LAYER M1 ;
        RECT 37.728 7.86 37.76 10.368 ;
  LAYER M1 ;
        RECT 37.792 7.86 37.824 10.368 ;
  LAYER M1 ;
        RECT 37.856 7.86 37.888 10.368 ;
  LAYER M1 ;
        RECT 37.92 7.86 37.952 10.368 ;
  LAYER M1 ;
        RECT 37.984 7.86 38.016 10.368 ;
  LAYER M1 ;
        RECT 38.048 7.86 38.08 10.368 ;
  LAYER M1 ;
        RECT 38.112 7.86 38.144 10.368 ;
  LAYER M1 ;
        RECT 38.176 7.86 38.208 10.368 ;
  LAYER M1 ;
        RECT 38.24 7.86 38.272 10.368 ;
  LAYER M1 ;
        RECT 38.304 7.86 38.336 10.368 ;
  LAYER M1 ;
        RECT 38.368 7.86 38.4 10.368 ;
  LAYER M1 ;
        RECT 38.432 7.86 38.464 10.368 ;
  LAYER M1 ;
        RECT 38.496 7.86 38.528 10.368 ;
  LAYER M1 ;
        RECT 38.56 7.86 38.592 10.368 ;
  LAYER M1 ;
        RECT 38.624 7.86 38.656 10.368 ;
  LAYER M1 ;
        RECT 38.688 7.86 38.72 10.368 ;
  LAYER M1 ;
        RECT 38.752 7.86 38.784 10.368 ;
  LAYER M1 ;
        RECT 38.816 7.86 38.848 10.368 ;
  LAYER M1 ;
        RECT 38.88 7.86 38.912 10.368 ;
  LAYER M1 ;
        RECT 38.944 7.86 38.976 10.368 ;
  LAYER M1 ;
        RECT 39.008 7.86 39.04 10.368 ;
  LAYER M1 ;
        RECT 39.072 7.86 39.104 10.368 ;
  LAYER M1 ;
        RECT 39.136 7.86 39.168 10.368 ;
  LAYER M1 ;
        RECT 39.2 7.86 39.232 10.368 ;
  LAYER M1 ;
        RECT 39.264 7.86 39.296 10.368 ;
  LAYER M1 ;
        RECT 39.328 7.86 39.36 10.368 ;
  LAYER M1 ;
        RECT 39.392 7.86 39.424 10.368 ;
  LAYER M1 ;
        RECT 39.456 7.86 39.488 10.368 ;
  LAYER M1 ;
        RECT 39.52 7.86 39.552 10.368 ;
  LAYER M1 ;
        RECT 39.584 7.86 39.616 10.368 ;
  LAYER M1 ;
        RECT 39.648 7.86 39.68 10.368 ;
  LAYER M2 ;
        RECT 37.324 10.252 39.796 10.284 ;
  LAYER M2 ;
        RECT 37.324 10.188 39.796 10.22 ;
  LAYER M2 ;
        RECT 37.324 10.124 39.796 10.156 ;
  LAYER M2 ;
        RECT 37.324 10.06 39.796 10.092 ;
  LAYER M2 ;
        RECT 37.324 9.996 39.796 10.028 ;
  LAYER M2 ;
        RECT 37.324 9.932 39.796 9.964 ;
  LAYER M2 ;
        RECT 37.324 9.868 39.796 9.9 ;
  LAYER M2 ;
        RECT 37.324 9.804 39.796 9.836 ;
  LAYER M2 ;
        RECT 37.324 9.74 39.796 9.772 ;
  LAYER M2 ;
        RECT 37.324 9.676 39.796 9.708 ;
  LAYER M2 ;
        RECT 37.324 9.612 39.796 9.644 ;
  LAYER M2 ;
        RECT 37.324 9.548 39.796 9.58 ;
  LAYER M2 ;
        RECT 37.324 9.484 39.796 9.516 ;
  LAYER M2 ;
        RECT 37.324 9.42 39.796 9.452 ;
  LAYER M2 ;
        RECT 37.324 9.356 39.796 9.388 ;
  LAYER M2 ;
        RECT 37.324 9.292 39.796 9.324 ;
  LAYER M2 ;
        RECT 37.324 9.228 39.796 9.26 ;
  LAYER M2 ;
        RECT 37.324 9.164 39.796 9.196 ;
  LAYER M2 ;
        RECT 37.324 9.1 39.796 9.132 ;
  LAYER M2 ;
        RECT 37.324 9.036 39.796 9.068 ;
  LAYER M2 ;
        RECT 37.324 8.972 39.796 9.004 ;
  LAYER M2 ;
        RECT 37.324 8.908 39.796 8.94 ;
  LAYER M2 ;
        RECT 37.324 8.844 39.796 8.876 ;
  LAYER M2 ;
        RECT 37.324 8.78 39.796 8.812 ;
  LAYER M2 ;
        RECT 37.324 8.716 39.796 8.748 ;
  LAYER M2 ;
        RECT 37.324 8.652 39.796 8.684 ;
  LAYER M2 ;
        RECT 37.324 8.588 39.796 8.62 ;
  LAYER M2 ;
        RECT 37.324 8.524 39.796 8.556 ;
  LAYER M2 ;
        RECT 37.324 8.46 39.796 8.492 ;
  LAYER M2 ;
        RECT 37.324 8.396 39.796 8.428 ;
  LAYER M2 ;
        RECT 37.324 8.332 39.796 8.364 ;
  LAYER M2 ;
        RECT 37.324 8.268 39.796 8.3 ;
  LAYER M2 ;
        RECT 37.324 8.204 39.796 8.236 ;
  LAYER M2 ;
        RECT 37.324 8.14 39.796 8.172 ;
  LAYER M2 ;
        RECT 37.324 8.076 39.796 8.108 ;
  LAYER M2 ;
        RECT 37.324 8.012 39.796 8.044 ;
  LAYER M3 ;
        RECT 37.344 7.86 37.376 10.368 ;
  LAYER M3 ;
        RECT 37.408 7.86 37.44 10.368 ;
  LAYER M3 ;
        RECT 37.472 7.86 37.504 10.368 ;
  LAYER M3 ;
        RECT 37.536 7.86 37.568 10.368 ;
  LAYER M3 ;
        RECT 37.6 7.86 37.632 10.368 ;
  LAYER M3 ;
        RECT 37.664 7.86 37.696 10.368 ;
  LAYER M3 ;
        RECT 37.728 7.86 37.76 10.368 ;
  LAYER M3 ;
        RECT 37.792 7.86 37.824 10.368 ;
  LAYER M3 ;
        RECT 37.856 7.86 37.888 10.368 ;
  LAYER M3 ;
        RECT 37.92 7.86 37.952 10.368 ;
  LAYER M3 ;
        RECT 37.984 7.86 38.016 10.368 ;
  LAYER M3 ;
        RECT 38.048 7.86 38.08 10.368 ;
  LAYER M3 ;
        RECT 38.112 7.86 38.144 10.368 ;
  LAYER M3 ;
        RECT 38.176 7.86 38.208 10.368 ;
  LAYER M3 ;
        RECT 38.24 7.86 38.272 10.368 ;
  LAYER M3 ;
        RECT 38.304 7.86 38.336 10.368 ;
  LAYER M3 ;
        RECT 38.368 7.86 38.4 10.368 ;
  LAYER M3 ;
        RECT 38.432 7.86 38.464 10.368 ;
  LAYER M3 ;
        RECT 38.496 7.86 38.528 10.368 ;
  LAYER M3 ;
        RECT 38.56 7.86 38.592 10.368 ;
  LAYER M3 ;
        RECT 38.624 7.86 38.656 10.368 ;
  LAYER M3 ;
        RECT 38.688 7.86 38.72 10.368 ;
  LAYER M3 ;
        RECT 38.752 7.86 38.784 10.368 ;
  LAYER M3 ;
        RECT 38.816 7.86 38.848 10.368 ;
  LAYER M3 ;
        RECT 38.88 7.86 38.912 10.368 ;
  LAYER M3 ;
        RECT 38.944 7.86 38.976 10.368 ;
  LAYER M3 ;
        RECT 39.008 7.86 39.04 10.368 ;
  LAYER M3 ;
        RECT 39.072 7.86 39.104 10.368 ;
  LAYER M3 ;
        RECT 39.136 7.86 39.168 10.368 ;
  LAYER M3 ;
        RECT 39.2 7.86 39.232 10.368 ;
  LAYER M3 ;
        RECT 39.264 7.86 39.296 10.368 ;
  LAYER M3 ;
        RECT 39.328 7.86 39.36 10.368 ;
  LAYER M3 ;
        RECT 39.392 7.86 39.424 10.368 ;
  LAYER M3 ;
        RECT 39.456 7.86 39.488 10.368 ;
  LAYER M3 ;
        RECT 39.52 7.86 39.552 10.368 ;
  LAYER M3 ;
        RECT 39.584 7.86 39.616 10.368 ;
  LAYER M3 ;
        RECT 39.648 7.86 39.68 10.368 ;
  LAYER M3 ;
        RECT 39.744 7.86 39.776 10.368 ;
  LAYER M1 ;
        RECT 37.359 7.896 37.361 10.332 ;
  LAYER M1 ;
        RECT 37.439 7.896 37.441 10.332 ;
  LAYER M1 ;
        RECT 37.519 7.896 37.521 10.332 ;
  LAYER M1 ;
        RECT 37.599 7.896 37.601 10.332 ;
  LAYER M1 ;
        RECT 37.679 7.896 37.681 10.332 ;
  LAYER M1 ;
        RECT 37.759 7.896 37.761 10.332 ;
  LAYER M1 ;
        RECT 37.839 7.896 37.841 10.332 ;
  LAYER M1 ;
        RECT 37.919 7.896 37.921 10.332 ;
  LAYER M1 ;
        RECT 37.999 7.896 38.001 10.332 ;
  LAYER M1 ;
        RECT 38.079 7.896 38.081 10.332 ;
  LAYER M1 ;
        RECT 38.159 7.896 38.161 10.332 ;
  LAYER M1 ;
        RECT 38.239 7.896 38.241 10.332 ;
  LAYER M1 ;
        RECT 38.319 7.896 38.321 10.332 ;
  LAYER M1 ;
        RECT 38.399 7.896 38.401 10.332 ;
  LAYER M1 ;
        RECT 38.479 7.896 38.481 10.332 ;
  LAYER M1 ;
        RECT 38.559 7.896 38.561 10.332 ;
  LAYER M1 ;
        RECT 38.639 7.896 38.641 10.332 ;
  LAYER M1 ;
        RECT 38.719 7.896 38.721 10.332 ;
  LAYER M1 ;
        RECT 38.799 7.896 38.801 10.332 ;
  LAYER M1 ;
        RECT 38.879 7.896 38.881 10.332 ;
  LAYER M1 ;
        RECT 38.959 7.896 38.961 10.332 ;
  LAYER M1 ;
        RECT 39.039 7.896 39.041 10.332 ;
  LAYER M1 ;
        RECT 39.119 7.896 39.121 10.332 ;
  LAYER M1 ;
        RECT 39.199 7.896 39.201 10.332 ;
  LAYER M1 ;
        RECT 39.279 7.896 39.281 10.332 ;
  LAYER M1 ;
        RECT 39.359 7.896 39.361 10.332 ;
  LAYER M1 ;
        RECT 39.439 7.896 39.441 10.332 ;
  LAYER M1 ;
        RECT 39.519 7.896 39.521 10.332 ;
  LAYER M1 ;
        RECT 39.599 7.896 39.601 10.332 ;
  LAYER M1 ;
        RECT 39.679 7.896 39.681 10.332 ;
  LAYER M2 ;
        RECT 37.36 10.331 39.76 10.333 ;
  LAYER M2 ;
        RECT 37.36 10.247 39.76 10.249 ;
  LAYER M2 ;
        RECT 37.36 10.163 39.76 10.165 ;
  LAYER M2 ;
        RECT 37.36 10.079 39.76 10.081 ;
  LAYER M2 ;
        RECT 37.36 9.995 39.76 9.997 ;
  LAYER M2 ;
        RECT 37.36 9.911 39.76 9.913 ;
  LAYER M2 ;
        RECT 37.36 9.827 39.76 9.829 ;
  LAYER M2 ;
        RECT 37.36 9.743 39.76 9.745 ;
  LAYER M2 ;
        RECT 37.36 9.659 39.76 9.661 ;
  LAYER M2 ;
        RECT 37.36 9.575 39.76 9.577 ;
  LAYER M2 ;
        RECT 37.36 9.491 39.76 9.493 ;
  LAYER M2 ;
        RECT 37.36 9.407 39.76 9.409 ;
  LAYER M2 ;
        RECT 37.36 9.3235 39.76 9.3255 ;
  LAYER M2 ;
        RECT 37.36 9.239 39.76 9.241 ;
  LAYER M2 ;
        RECT 37.36 9.155 39.76 9.157 ;
  LAYER M2 ;
        RECT 37.36 9.071 39.76 9.073 ;
  LAYER M2 ;
        RECT 37.36 8.987 39.76 8.989 ;
  LAYER M2 ;
        RECT 37.36 8.903 39.76 8.905 ;
  LAYER M2 ;
        RECT 37.36 8.819 39.76 8.821 ;
  LAYER M2 ;
        RECT 37.36 8.735 39.76 8.737 ;
  LAYER M2 ;
        RECT 37.36 8.651 39.76 8.653 ;
  LAYER M2 ;
        RECT 37.36 8.567 39.76 8.569 ;
  LAYER M2 ;
        RECT 37.36 8.483 39.76 8.485 ;
  LAYER M2 ;
        RECT 37.36 8.399 39.76 8.401 ;
  LAYER M2 ;
        RECT 37.36 8.315 39.76 8.317 ;
  LAYER M2 ;
        RECT 37.36 8.231 39.76 8.233 ;
  LAYER M2 ;
        RECT 37.36 8.147 39.76 8.149 ;
  LAYER M2 ;
        RECT 37.36 8.063 39.76 8.065 ;
  LAYER M2 ;
        RECT 37.36 7.979 39.76 7.981 ;
  LAYER M1 ;
        RECT 37.344 4.92 37.376 7.428 ;
  LAYER M1 ;
        RECT 37.408 4.92 37.44 7.428 ;
  LAYER M1 ;
        RECT 37.472 4.92 37.504 7.428 ;
  LAYER M1 ;
        RECT 37.536 4.92 37.568 7.428 ;
  LAYER M1 ;
        RECT 37.6 4.92 37.632 7.428 ;
  LAYER M1 ;
        RECT 37.664 4.92 37.696 7.428 ;
  LAYER M1 ;
        RECT 37.728 4.92 37.76 7.428 ;
  LAYER M1 ;
        RECT 37.792 4.92 37.824 7.428 ;
  LAYER M1 ;
        RECT 37.856 4.92 37.888 7.428 ;
  LAYER M1 ;
        RECT 37.92 4.92 37.952 7.428 ;
  LAYER M1 ;
        RECT 37.984 4.92 38.016 7.428 ;
  LAYER M1 ;
        RECT 38.048 4.92 38.08 7.428 ;
  LAYER M1 ;
        RECT 38.112 4.92 38.144 7.428 ;
  LAYER M1 ;
        RECT 38.176 4.92 38.208 7.428 ;
  LAYER M1 ;
        RECT 38.24 4.92 38.272 7.428 ;
  LAYER M1 ;
        RECT 38.304 4.92 38.336 7.428 ;
  LAYER M1 ;
        RECT 38.368 4.92 38.4 7.428 ;
  LAYER M1 ;
        RECT 38.432 4.92 38.464 7.428 ;
  LAYER M1 ;
        RECT 38.496 4.92 38.528 7.428 ;
  LAYER M1 ;
        RECT 38.56 4.92 38.592 7.428 ;
  LAYER M1 ;
        RECT 38.624 4.92 38.656 7.428 ;
  LAYER M1 ;
        RECT 38.688 4.92 38.72 7.428 ;
  LAYER M1 ;
        RECT 38.752 4.92 38.784 7.428 ;
  LAYER M1 ;
        RECT 38.816 4.92 38.848 7.428 ;
  LAYER M1 ;
        RECT 38.88 4.92 38.912 7.428 ;
  LAYER M1 ;
        RECT 38.944 4.92 38.976 7.428 ;
  LAYER M1 ;
        RECT 39.008 4.92 39.04 7.428 ;
  LAYER M1 ;
        RECT 39.072 4.92 39.104 7.428 ;
  LAYER M1 ;
        RECT 39.136 4.92 39.168 7.428 ;
  LAYER M1 ;
        RECT 39.2 4.92 39.232 7.428 ;
  LAYER M1 ;
        RECT 39.264 4.92 39.296 7.428 ;
  LAYER M1 ;
        RECT 39.328 4.92 39.36 7.428 ;
  LAYER M1 ;
        RECT 39.392 4.92 39.424 7.428 ;
  LAYER M1 ;
        RECT 39.456 4.92 39.488 7.428 ;
  LAYER M1 ;
        RECT 39.52 4.92 39.552 7.428 ;
  LAYER M1 ;
        RECT 39.584 4.92 39.616 7.428 ;
  LAYER M1 ;
        RECT 39.648 4.92 39.68 7.428 ;
  LAYER M2 ;
        RECT 37.324 7.312 39.796 7.344 ;
  LAYER M2 ;
        RECT 37.324 7.248 39.796 7.28 ;
  LAYER M2 ;
        RECT 37.324 7.184 39.796 7.216 ;
  LAYER M2 ;
        RECT 37.324 7.12 39.796 7.152 ;
  LAYER M2 ;
        RECT 37.324 7.056 39.796 7.088 ;
  LAYER M2 ;
        RECT 37.324 6.992 39.796 7.024 ;
  LAYER M2 ;
        RECT 37.324 6.928 39.796 6.96 ;
  LAYER M2 ;
        RECT 37.324 6.864 39.796 6.896 ;
  LAYER M2 ;
        RECT 37.324 6.8 39.796 6.832 ;
  LAYER M2 ;
        RECT 37.324 6.736 39.796 6.768 ;
  LAYER M2 ;
        RECT 37.324 6.672 39.796 6.704 ;
  LAYER M2 ;
        RECT 37.324 6.608 39.796 6.64 ;
  LAYER M2 ;
        RECT 37.324 6.544 39.796 6.576 ;
  LAYER M2 ;
        RECT 37.324 6.48 39.796 6.512 ;
  LAYER M2 ;
        RECT 37.324 6.416 39.796 6.448 ;
  LAYER M2 ;
        RECT 37.324 6.352 39.796 6.384 ;
  LAYER M2 ;
        RECT 37.324 6.288 39.796 6.32 ;
  LAYER M2 ;
        RECT 37.324 6.224 39.796 6.256 ;
  LAYER M2 ;
        RECT 37.324 6.16 39.796 6.192 ;
  LAYER M2 ;
        RECT 37.324 6.096 39.796 6.128 ;
  LAYER M2 ;
        RECT 37.324 6.032 39.796 6.064 ;
  LAYER M2 ;
        RECT 37.324 5.968 39.796 6 ;
  LAYER M2 ;
        RECT 37.324 5.904 39.796 5.936 ;
  LAYER M2 ;
        RECT 37.324 5.84 39.796 5.872 ;
  LAYER M2 ;
        RECT 37.324 5.776 39.796 5.808 ;
  LAYER M2 ;
        RECT 37.324 5.712 39.796 5.744 ;
  LAYER M2 ;
        RECT 37.324 5.648 39.796 5.68 ;
  LAYER M2 ;
        RECT 37.324 5.584 39.796 5.616 ;
  LAYER M2 ;
        RECT 37.324 5.52 39.796 5.552 ;
  LAYER M2 ;
        RECT 37.324 5.456 39.796 5.488 ;
  LAYER M2 ;
        RECT 37.324 5.392 39.796 5.424 ;
  LAYER M2 ;
        RECT 37.324 5.328 39.796 5.36 ;
  LAYER M2 ;
        RECT 37.324 5.264 39.796 5.296 ;
  LAYER M2 ;
        RECT 37.324 5.2 39.796 5.232 ;
  LAYER M2 ;
        RECT 37.324 5.136 39.796 5.168 ;
  LAYER M2 ;
        RECT 37.324 5.072 39.796 5.104 ;
  LAYER M3 ;
        RECT 37.344 4.92 37.376 7.428 ;
  LAYER M3 ;
        RECT 37.408 4.92 37.44 7.428 ;
  LAYER M3 ;
        RECT 37.472 4.92 37.504 7.428 ;
  LAYER M3 ;
        RECT 37.536 4.92 37.568 7.428 ;
  LAYER M3 ;
        RECT 37.6 4.92 37.632 7.428 ;
  LAYER M3 ;
        RECT 37.664 4.92 37.696 7.428 ;
  LAYER M3 ;
        RECT 37.728 4.92 37.76 7.428 ;
  LAYER M3 ;
        RECT 37.792 4.92 37.824 7.428 ;
  LAYER M3 ;
        RECT 37.856 4.92 37.888 7.428 ;
  LAYER M3 ;
        RECT 37.92 4.92 37.952 7.428 ;
  LAYER M3 ;
        RECT 37.984 4.92 38.016 7.428 ;
  LAYER M3 ;
        RECT 38.048 4.92 38.08 7.428 ;
  LAYER M3 ;
        RECT 38.112 4.92 38.144 7.428 ;
  LAYER M3 ;
        RECT 38.176 4.92 38.208 7.428 ;
  LAYER M3 ;
        RECT 38.24 4.92 38.272 7.428 ;
  LAYER M3 ;
        RECT 38.304 4.92 38.336 7.428 ;
  LAYER M3 ;
        RECT 38.368 4.92 38.4 7.428 ;
  LAYER M3 ;
        RECT 38.432 4.92 38.464 7.428 ;
  LAYER M3 ;
        RECT 38.496 4.92 38.528 7.428 ;
  LAYER M3 ;
        RECT 38.56 4.92 38.592 7.428 ;
  LAYER M3 ;
        RECT 38.624 4.92 38.656 7.428 ;
  LAYER M3 ;
        RECT 38.688 4.92 38.72 7.428 ;
  LAYER M3 ;
        RECT 38.752 4.92 38.784 7.428 ;
  LAYER M3 ;
        RECT 38.816 4.92 38.848 7.428 ;
  LAYER M3 ;
        RECT 38.88 4.92 38.912 7.428 ;
  LAYER M3 ;
        RECT 38.944 4.92 38.976 7.428 ;
  LAYER M3 ;
        RECT 39.008 4.92 39.04 7.428 ;
  LAYER M3 ;
        RECT 39.072 4.92 39.104 7.428 ;
  LAYER M3 ;
        RECT 39.136 4.92 39.168 7.428 ;
  LAYER M3 ;
        RECT 39.2 4.92 39.232 7.428 ;
  LAYER M3 ;
        RECT 39.264 4.92 39.296 7.428 ;
  LAYER M3 ;
        RECT 39.328 4.92 39.36 7.428 ;
  LAYER M3 ;
        RECT 39.392 4.92 39.424 7.428 ;
  LAYER M3 ;
        RECT 39.456 4.92 39.488 7.428 ;
  LAYER M3 ;
        RECT 39.52 4.92 39.552 7.428 ;
  LAYER M3 ;
        RECT 39.584 4.92 39.616 7.428 ;
  LAYER M3 ;
        RECT 39.648 4.92 39.68 7.428 ;
  LAYER M3 ;
        RECT 39.744 4.92 39.776 7.428 ;
  LAYER M1 ;
        RECT 37.359 4.956 37.361 7.392 ;
  LAYER M1 ;
        RECT 37.439 4.956 37.441 7.392 ;
  LAYER M1 ;
        RECT 37.519 4.956 37.521 7.392 ;
  LAYER M1 ;
        RECT 37.599 4.956 37.601 7.392 ;
  LAYER M1 ;
        RECT 37.679 4.956 37.681 7.392 ;
  LAYER M1 ;
        RECT 37.759 4.956 37.761 7.392 ;
  LAYER M1 ;
        RECT 37.839 4.956 37.841 7.392 ;
  LAYER M1 ;
        RECT 37.919 4.956 37.921 7.392 ;
  LAYER M1 ;
        RECT 37.999 4.956 38.001 7.392 ;
  LAYER M1 ;
        RECT 38.079 4.956 38.081 7.392 ;
  LAYER M1 ;
        RECT 38.159 4.956 38.161 7.392 ;
  LAYER M1 ;
        RECT 38.239 4.956 38.241 7.392 ;
  LAYER M1 ;
        RECT 38.319 4.956 38.321 7.392 ;
  LAYER M1 ;
        RECT 38.399 4.956 38.401 7.392 ;
  LAYER M1 ;
        RECT 38.479 4.956 38.481 7.392 ;
  LAYER M1 ;
        RECT 38.559 4.956 38.561 7.392 ;
  LAYER M1 ;
        RECT 38.639 4.956 38.641 7.392 ;
  LAYER M1 ;
        RECT 38.719 4.956 38.721 7.392 ;
  LAYER M1 ;
        RECT 38.799 4.956 38.801 7.392 ;
  LAYER M1 ;
        RECT 38.879 4.956 38.881 7.392 ;
  LAYER M1 ;
        RECT 38.959 4.956 38.961 7.392 ;
  LAYER M1 ;
        RECT 39.039 4.956 39.041 7.392 ;
  LAYER M1 ;
        RECT 39.119 4.956 39.121 7.392 ;
  LAYER M1 ;
        RECT 39.199 4.956 39.201 7.392 ;
  LAYER M1 ;
        RECT 39.279 4.956 39.281 7.392 ;
  LAYER M1 ;
        RECT 39.359 4.956 39.361 7.392 ;
  LAYER M1 ;
        RECT 39.439 4.956 39.441 7.392 ;
  LAYER M1 ;
        RECT 39.519 4.956 39.521 7.392 ;
  LAYER M1 ;
        RECT 39.599 4.956 39.601 7.392 ;
  LAYER M1 ;
        RECT 39.679 4.956 39.681 7.392 ;
  LAYER M2 ;
        RECT 37.36 7.391 39.76 7.393 ;
  LAYER M2 ;
        RECT 37.36 7.307 39.76 7.309 ;
  LAYER M2 ;
        RECT 37.36 7.223 39.76 7.225 ;
  LAYER M2 ;
        RECT 37.36 7.139 39.76 7.141 ;
  LAYER M2 ;
        RECT 37.36 7.055 39.76 7.057 ;
  LAYER M2 ;
        RECT 37.36 6.971 39.76 6.973 ;
  LAYER M2 ;
        RECT 37.36 6.887 39.76 6.889 ;
  LAYER M2 ;
        RECT 37.36 6.803 39.76 6.805 ;
  LAYER M2 ;
        RECT 37.36 6.719 39.76 6.721 ;
  LAYER M2 ;
        RECT 37.36 6.635 39.76 6.637 ;
  LAYER M2 ;
        RECT 37.36 6.551 39.76 6.553 ;
  LAYER M2 ;
        RECT 37.36 6.467 39.76 6.469 ;
  LAYER M2 ;
        RECT 37.36 6.3835 39.76 6.3855 ;
  LAYER M2 ;
        RECT 37.36 6.299 39.76 6.301 ;
  LAYER M2 ;
        RECT 37.36 6.215 39.76 6.217 ;
  LAYER M2 ;
        RECT 37.36 6.131 39.76 6.133 ;
  LAYER M2 ;
        RECT 37.36 6.047 39.76 6.049 ;
  LAYER M2 ;
        RECT 37.36 5.963 39.76 5.965 ;
  LAYER M2 ;
        RECT 37.36 5.879 39.76 5.881 ;
  LAYER M2 ;
        RECT 37.36 5.795 39.76 5.797 ;
  LAYER M2 ;
        RECT 37.36 5.711 39.76 5.713 ;
  LAYER M2 ;
        RECT 37.36 5.627 39.76 5.629 ;
  LAYER M2 ;
        RECT 37.36 5.543 39.76 5.545 ;
  LAYER M2 ;
        RECT 37.36 5.459 39.76 5.461 ;
  LAYER M2 ;
        RECT 37.36 5.375 39.76 5.377 ;
  LAYER M2 ;
        RECT 37.36 5.291 39.76 5.293 ;
  LAYER M2 ;
        RECT 37.36 5.207 39.76 5.209 ;
  LAYER M2 ;
        RECT 37.36 5.123 39.76 5.125 ;
  LAYER M2 ;
        RECT 37.36 5.039 39.76 5.041 ;
  LAYER M1 ;
        RECT 37.344 1.98 37.376 4.488 ;
  LAYER M1 ;
        RECT 37.408 1.98 37.44 4.488 ;
  LAYER M1 ;
        RECT 37.472 1.98 37.504 4.488 ;
  LAYER M1 ;
        RECT 37.536 1.98 37.568 4.488 ;
  LAYER M1 ;
        RECT 37.6 1.98 37.632 4.488 ;
  LAYER M1 ;
        RECT 37.664 1.98 37.696 4.488 ;
  LAYER M1 ;
        RECT 37.728 1.98 37.76 4.488 ;
  LAYER M1 ;
        RECT 37.792 1.98 37.824 4.488 ;
  LAYER M1 ;
        RECT 37.856 1.98 37.888 4.488 ;
  LAYER M1 ;
        RECT 37.92 1.98 37.952 4.488 ;
  LAYER M1 ;
        RECT 37.984 1.98 38.016 4.488 ;
  LAYER M1 ;
        RECT 38.048 1.98 38.08 4.488 ;
  LAYER M1 ;
        RECT 38.112 1.98 38.144 4.488 ;
  LAYER M1 ;
        RECT 38.176 1.98 38.208 4.488 ;
  LAYER M1 ;
        RECT 38.24 1.98 38.272 4.488 ;
  LAYER M1 ;
        RECT 38.304 1.98 38.336 4.488 ;
  LAYER M1 ;
        RECT 38.368 1.98 38.4 4.488 ;
  LAYER M1 ;
        RECT 38.432 1.98 38.464 4.488 ;
  LAYER M1 ;
        RECT 38.496 1.98 38.528 4.488 ;
  LAYER M1 ;
        RECT 38.56 1.98 38.592 4.488 ;
  LAYER M1 ;
        RECT 38.624 1.98 38.656 4.488 ;
  LAYER M1 ;
        RECT 38.688 1.98 38.72 4.488 ;
  LAYER M1 ;
        RECT 38.752 1.98 38.784 4.488 ;
  LAYER M1 ;
        RECT 38.816 1.98 38.848 4.488 ;
  LAYER M1 ;
        RECT 38.88 1.98 38.912 4.488 ;
  LAYER M1 ;
        RECT 38.944 1.98 38.976 4.488 ;
  LAYER M1 ;
        RECT 39.008 1.98 39.04 4.488 ;
  LAYER M1 ;
        RECT 39.072 1.98 39.104 4.488 ;
  LAYER M1 ;
        RECT 39.136 1.98 39.168 4.488 ;
  LAYER M1 ;
        RECT 39.2 1.98 39.232 4.488 ;
  LAYER M1 ;
        RECT 39.264 1.98 39.296 4.488 ;
  LAYER M1 ;
        RECT 39.328 1.98 39.36 4.488 ;
  LAYER M1 ;
        RECT 39.392 1.98 39.424 4.488 ;
  LAYER M1 ;
        RECT 39.456 1.98 39.488 4.488 ;
  LAYER M1 ;
        RECT 39.52 1.98 39.552 4.488 ;
  LAYER M1 ;
        RECT 39.584 1.98 39.616 4.488 ;
  LAYER M1 ;
        RECT 39.648 1.98 39.68 4.488 ;
  LAYER M2 ;
        RECT 37.324 4.372 39.796 4.404 ;
  LAYER M2 ;
        RECT 37.324 4.308 39.796 4.34 ;
  LAYER M2 ;
        RECT 37.324 4.244 39.796 4.276 ;
  LAYER M2 ;
        RECT 37.324 4.18 39.796 4.212 ;
  LAYER M2 ;
        RECT 37.324 4.116 39.796 4.148 ;
  LAYER M2 ;
        RECT 37.324 4.052 39.796 4.084 ;
  LAYER M2 ;
        RECT 37.324 3.988 39.796 4.02 ;
  LAYER M2 ;
        RECT 37.324 3.924 39.796 3.956 ;
  LAYER M2 ;
        RECT 37.324 3.86 39.796 3.892 ;
  LAYER M2 ;
        RECT 37.324 3.796 39.796 3.828 ;
  LAYER M2 ;
        RECT 37.324 3.732 39.796 3.764 ;
  LAYER M2 ;
        RECT 37.324 3.668 39.796 3.7 ;
  LAYER M2 ;
        RECT 37.324 3.604 39.796 3.636 ;
  LAYER M2 ;
        RECT 37.324 3.54 39.796 3.572 ;
  LAYER M2 ;
        RECT 37.324 3.476 39.796 3.508 ;
  LAYER M2 ;
        RECT 37.324 3.412 39.796 3.444 ;
  LAYER M2 ;
        RECT 37.324 3.348 39.796 3.38 ;
  LAYER M2 ;
        RECT 37.324 3.284 39.796 3.316 ;
  LAYER M2 ;
        RECT 37.324 3.22 39.796 3.252 ;
  LAYER M2 ;
        RECT 37.324 3.156 39.796 3.188 ;
  LAYER M2 ;
        RECT 37.324 3.092 39.796 3.124 ;
  LAYER M2 ;
        RECT 37.324 3.028 39.796 3.06 ;
  LAYER M2 ;
        RECT 37.324 2.964 39.796 2.996 ;
  LAYER M2 ;
        RECT 37.324 2.9 39.796 2.932 ;
  LAYER M2 ;
        RECT 37.324 2.836 39.796 2.868 ;
  LAYER M2 ;
        RECT 37.324 2.772 39.796 2.804 ;
  LAYER M2 ;
        RECT 37.324 2.708 39.796 2.74 ;
  LAYER M2 ;
        RECT 37.324 2.644 39.796 2.676 ;
  LAYER M2 ;
        RECT 37.324 2.58 39.796 2.612 ;
  LAYER M2 ;
        RECT 37.324 2.516 39.796 2.548 ;
  LAYER M2 ;
        RECT 37.324 2.452 39.796 2.484 ;
  LAYER M2 ;
        RECT 37.324 2.388 39.796 2.42 ;
  LAYER M2 ;
        RECT 37.324 2.324 39.796 2.356 ;
  LAYER M2 ;
        RECT 37.324 2.26 39.796 2.292 ;
  LAYER M2 ;
        RECT 37.324 2.196 39.796 2.228 ;
  LAYER M2 ;
        RECT 37.324 2.132 39.796 2.164 ;
  LAYER M3 ;
        RECT 37.344 1.98 37.376 4.488 ;
  LAYER M3 ;
        RECT 37.408 1.98 37.44 4.488 ;
  LAYER M3 ;
        RECT 37.472 1.98 37.504 4.488 ;
  LAYER M3 ;
        RECT 37.536 1.98 37.568 4.488 ;
  LAYER M3 ;
        RECT 37.6 1.98 37.632 4.488 ;
  LAYER M3 ;
        RECT 37.664 1.98 37.696 4.488 ;
  LAYER M3 ;
        RECT 37.728 1.98 37.76 4.488 ;
  LAYER M3 ;
        RECT 37.792 1.98 37.824 4.488 ;
  LAYER M3 ;
        RECT 37.856 1.98 37.888 4.488 ;
  LAYER M3 ;
        RECT 37.92 1.98 37.952 4.488 ;
  LAYER M3 ;
        RECT 37.984 1.98 38.016 4.488 ;
  LAYER M3 ;
        RECT 38.048 1.98 38.08 4.488 ;
  LAYER M3 ;
        RECT 38.112 1.98 38.144 4.488 ;
  LAYER M3 ;
        RECT 38.176 1.98 38.208 4.488 ;
  LAYER M3 ;
        RECT 38.24 1.98 38.272 4.488 ;
  LAYER M3 ;
        RECT 38.304 1.98 38.336 4.488 ;
  LAYER M3 ;
        RECT 38.368 1.98 38.4 4.488 ;
  LAYER M3 ;
        RECT 38.432 1.98 38.464 4.488 ;
  LAYER M3 ;
        RECT 38.496 1.98 38.528 4.488 ;
  LAYER M3 ;
        RECT 38.56 1.98 38.592 4.488 ;
  LAYER M3 ;
        RECT 38.624 1.98 38.656 4.488 ;
  LAYER M3 ;
        RECT 38.688 1.98 38.72 4.488 ;
  LAYER M3 ;
        RECT 38.752 1.98 38.784 4.488 ;
  LAYER M3 ;
        RECT 38.816 1.98 38.848 4.488 ;
  LAYER M3 ;
        RECT 38.88 1.98 38.912 4.488 ;
  LAYER M3 ;
        RECT 38.944 1.98 38.976 4.488 ;
  LAYER M3 ;
        RECT 39.008 1.98 39.04 4.488 ;
  LAYER M3 ;
        RECT 39.072 1.98 39.104 4.488 ;
  LAYER M3 ;
        RECT 39.136 1.98 39.168 4.488 ;
  LAYER M3 ;
        RECT 39.2 1.98 39.232 4.488 ;
  LAYER M3 ;
        RECT 39.264 1.98 39.296 4.488 ;
  LAYER M3 ;
        RECT 39.328 1.98 39.36 4.488 ;
  LAYER M3 ;
        RECT 39.392 1.98 39.424 4.488 ;
  LAYER M3 ;
        RECT 39.456 1.98 39.488 4.488 ;
  LAYER M3 ;
        RECT 39.52 1.98 39.552 4.488 ;
  LAYER M3 ;
        RECT 39.584 1.98 39.616 4.488 ;
  LAYER M3 ;
        RECT 39.648 1.98 39.68 4.488 ;
  LAYER M3 ;
        RECT 39.744 1.98 39.776 4.488 ;
  LAYER M1 ;
        RECT 37.359 2.016 37.361 4.452 ;
  LAYER M1 ;
        RECT 37.439 2.016 37.441 4.452 ;
  LAYER M1 ;
        RECT 37.519 2.016 37.521 4.452 ;
  LAYER M1 ;
        RECT 37.599 2.016 37.601 4.452 ;
  LAYER M1 ;
        RECT 37.679 2.016 37.681 4.452 ;
  LAYER M1 ;
        RECT 37.759 2.016 37.761 4.452 ;
  LAYER M1 ;
        RECT 37.839 2.016 37.841 4.452 ;
  LAYER M1 ;
        RECT 37.919 2.016 37.921 4.452 ;
  LAYER M1 ;
        RECT 37.999 2.016 38.001 4.452 ;
  LAYER M1 ;
        RECT 38.079 2.016 38.081 4.452 ;
  LAYER M1 ;
        RECT 38.159 2.016 38.161 4.452 ;
  LAYER M1 ;
        RECT 38.239 2.016 38.241 4.452 ;
  LAYER M1 ;
        RECT 38.319 2.016 38.321 4.452 ;
  LAYER M1 ;
        RECT 38.399 2.016 38.401 4.452 ;
  LAYER M1 ;
        RECT 38.479 2.016 38.481 4.452 ;
  LAYER M1 ;
        RECT 38.559 2.016 38.561 4.452 ;
  LAYER M1 ;
        RECT 38.639 2.016 38.641 4.452 ;
  LAYER M1 ;
        RECT 38.719 2.016 38.721 4.452 ;
  LAYER M1 ;
        RECT 38.799 2.016 38.801 4.452 ;
  LAYER M1 ;
        RECT 38.879 2.016 38.881 4.452 ;
  LAYER M1 ;
        RECT 38.959 2.016 38.961 4.452 ;
  LAYER M1 ;
        RECT 39.039 2.016 39.041 4.452 ;
  LAYER M1 ;
        RECT 39.119 2.016 39.121 4.452 ;
  LAYER M1 ;
        RECT 39.199 2.016 39.201 4.452 ;
  LAYER M1 ;
        RECT 39.279 2.016 39.281 4.452 ;
  LAYER M1 ;
        RECT 39.359 2.016 39.361 4.452 ;
  LAYER M1 ;
        RECT 39.439 2.016 39.441 4.452 ;
  LAYER M1 ;
        RECT 39.519 2.016 39.521 4.452 ;
  LAYER M1 ;
        RECT 39.599 2.016 39.601 4.452 ;
  LAYER M1 ;
        RECT 39.679 2.016 39.681 4.452 ;
  LAYER M2 ;
        RECT 37.36 4.451 39.76 4.453 ;
  LAYER M2 ;
        RECT 37.36 4.367 39.76 4.369 ;
  LAYER M2 ;
        RECT 37.36 4.283 39.76 4.285 ;
  LAYER M2 ;
        RECT 37.36 4.199 39.76 4.201 ;
  LAYER M2 ;
        RECT 37.36 4.115 39.76 4.117 ;
  LAYER M2 ;
        RECT 37.36 4.031 39.76 4.033 ;
  LAYER M2 ;
        RECT 37.36 3.947 39.76 3.949 ;
  LAYER M2 ;
        RECT 37.36 3.863 39.76 3.865 ;
  LAYER M2 ;
        RECT 37.36 3.779 39.76 3.781 ;
  LAYER M2 ;
        RECT 37.36 3.695 39.76 3.697 ;
  LAYER M2 ;
        RECT 37.36 3.611 39.76 3.613 ;
  LAYER M2 ;
        RECT 37.36 3.527 39.76 3.529 ;
  LAYER M2 ;
        RECT 37.36 3.4435 39.76 3.4455 ;
  LAYER M2 ;
        RECT 37.36 3.359 39.76 3.361 ;
  LAYER M2 ;
        RECT 37.36 3.275 39.76 3.277 ;
  LAYER M2 ;
        RECT 37.36 3.191 39.76 3.193 ;
  LAYER M2 ;
        RECT 37.36 3.107 39.76 3.109 ;
  LAYER M2 ;
        RECT 37.36 3.023 39.76 3.025 ;
  LAYER M2 ;
        RECT 37.36 2.939 39.76 2.941 ;
  LAYER M2 ;
        RECT 37.36 2.855 39.76 2.857 ;
  LAYER M2 ;
        RECT 37.36 2.771 39.76 2.773 ;
  LAYER M2 ;
        RECT 37.36 2.687 39.76 2.689 ;
  LAYER M2 ;
        RECT 37.36 2.603 39.76 2.605 ;
  LAYER M2 ;
        RECT 37.36 2.519 39.76 2.521 ;
  LAYER M2 ;
        RECT 37.36 2.435 39.76 2.437 ;
  LAYER M2 ;
        RECT 37.36 2.351 39.76 2.353 ;
  LAYER M2 ;
        RECT 37.36 2.267 39.76 2.269 ;
  LAYER M2 ;
        RECT 37.36 2.183 39.76 2.185 ;
  LAYER M2 ;
        RECT 37.36 2.099 39.76 2.101 ;
  LAYER M1 ;
        RECT 40.224 13.74 40.256 16.248 ;
  LAYER M1 ;
        RECT 40.288 13.74 40.32 16.248 ;
  LAYER M1 ;
        RECT 40.352 13.74 40.384 16.248 ;
  LAYER M1 ;
        RECT 40.416 13.74 40.448 16.248 ;
  LAYER M1 ;
        RECT 40.48 13.74 40.512 16.248 ;
  LAYER M1 ;
        RECT 40.544 13.74 40.576 16.248 ;
  LAYER M1 ;
        RECT 40.608 13.74 40.64 16.248 ;
  LAYER M1 ;
        RECT 40.672 13.74 40.704 16.248 ;
  LAYER M1 ;
        RECT 40.736 13.74 40.768 16.248 ;
  LAYER M1 ;
        RECT 40.8 13.74 40.832 16.248 ;
  LAYER M1 ;
        RECT 40.864 13.74 40.896 16.248 ;
  LAYER M1 ;
        RECT 40.928 13.74 40.96 16.248 ;
  LAYER M1 ;
        RECT 40.992 13.74 41.024 16.248 ;
  LAYER M1 ;
        RECT 41.056 13.74 41.088 16.248 ;
  LAYER M1 ;
        RECT 41.12 13.74 41.152 16.248 ;
  LAYER M1 ;
        RECT 41.184 13.74 41.216 16.248 ;
  LAYER M1 ;
        RECT 41.248 13.74 41.28 16.248 ;
  LAYER M1 ;
        RECT 41.312 13.74 41.344 16.248 ;
  LAYER M1 ;
        RECT 41.376 13.74 41.408 16.248 ;
  LAYER M1 ;
        RECT 41.44 13.74 41.472 16.248 ;
  LAYER M1 ;
        RECT 41.504 13.74 41.536 16.248 ;
  LAYER M1 ;
        RECT 41.568 13.74 41.6 16.248 ;
  LAYER M1 ;
        RECT 41.632 13.74 41.664 16.248 ;
  LAYER M1 ;
        RECT 41.696 13.74 41.728 16.248 ;
  LAYER M1 ;
        RECT 41.76 13.74 41.792 16.248 ;
  LAYER M1 ;
        RECT 41.824 13.74 41.856 16.248 ;
  LAYER M1 ;
        RECT 41.888 13.74 41.92 16.248 ;
  LAYER M1 ;
        RECT 41.952 13.74 41.984 16.248 ;
  LAYER M1 ;
        RECT 42.016 13.74 42.048 16.248 ;
  LAYER M1 ;
        RECT 42.08 13.74 42.112 16.248 ;
  LAYER M1 ;
        RECT 42.144 13.74 42.176 16.248 ;
  LAYER M1 ;
        RECT 42.208 13.74 42.24 16.248 ;
  LAYER M1 ;
        RECT 42.272 13.74 42.304 16.248 ;
  LAYER M1 ;
        RECT 42.336 13.74 42.368 16.248 ;
  LAYER M1 ;
        RECT 42.4 13.74 42.432 16.248 ;
  LAYER M1 ;
        RECT 42.464 13.74 42.496 16.248 ;
  LAYER M1 ;
        RECT 42.528 13.74 42.56 16.248 ;
  LAYER M2 ;
        RECT 40.204 16.132 42.676 16.164 ;
  LAYER M2 ;
        RECT 40.204 16.068 42.676 16.1 ;
  LAYER M2 ;
        RECT 40.204 16.004 42.676 16.036 ;
  LAYER M2 ;
        RECT 40.204 15.94 42.676 15.972 ;
  LAYER M2 ;
        RECT 40.204 15.876 42.676 15.908 ;
  LAYER M2 ;
        RECT 40.204 15.812 42.676 15.844 ;
  LAYER M2 ;
        RECT 40.204 15.748 42.676 15.78 ;
  LAYER M2 ;
        RECT 40.204 15.684 42.676 15.716 ;
  LAYER M2 ;
        RECT 40.204 15.62 42.676 15.652 ;
  LAYER M2 ;
        RECT 40.204 15.556 42.676 15.588 ;
  LAYER M2 ;
        RECT 40.204 15.492 42.676 15.524 ;
  LAYER M2 ;
        RECT 40.204 15.428 42.676 15.46 ;
  LAYER M2 ;
        RECT 40.204 15.364 42.676 15.396 ;
  LAYER M2 ;
        RECT 40.204 15.3 42.676 15.332 ;
  LAYER M2 ;
        RECT 40.204 15.236 42.676 15.268 ;
  LAYER M2 ;
        RECT 40.204 15.172 42.676 15.204 ;
  LAYER M2 ;
        RECT 40.204 15.108 42.676 15.14 ;
  LAYER M2 ;
        RECT 40.204 15.044 42.676 15.076 ;
  LAYER M2 ;
        RECT 40.204 14.98 42.676 15.012 ;
  LAYER M2 ;
        RECT 40.204 14.916 42.676 14.948 ;
  LAYER M2 ;
        RECT 40.204 14.852 42.676 14.884 ;
  LAYER M2 ;
        RECT 40.204 14.788 42.676 14.82 ;
  LAYER M2 ;
        RECT 40.204 14.724 42.676 14.756 ;
  LAYER M2 ;
        RECT 40.204 14.66 42.676 14.692 ;
  LAYER M2 ;
        RECT 40.204 14.596 42.676 14.628 ;
  LAYER M2 ;
        RECT 40.204 14.532 42.676 14.564 ;
  LAYER M2 ;
        RECT 40.204 14.468 42.676 14.5 ;
  LAYER M2 ;
        RECT 40.204 14.404 42.676 14.436 ;
  LAYER M2 ;
        RECT 40.204 14.34 42.676 14.372 ;
  LAYER M2 ;
        RECT 40.204 14.276 42.676 14.308 ;
  LAYER M2 ;
        RECT 40.204 14.212 42.676 14.244 ;
  LAYER M2 ;
        RECT 40.204 14.148 42.676 14.18 ;
  LAYER M2 ;
        RECT 40.204 14.084 42.676 14.116 ;
  LAYER M2 ;
        RECT 40.204 14.02 42.676 14.052 ;
  LAYER M2 ;
        RECT 40.204 13.956 42.676 13.988 ;
  LAYER M2 ;
        RECT 40.204 13.892 42.676 13.924 ;
  LAYER M3 ;
        RECT 40.224 13.74 40.256 16.248 ;
  LAYER M3 ;
        RECT 40.288 13.74 40.32 16.248 ;
  LAYER M3 ;
        RECT 40.352 13.74 40.384 16.248 ;
  LAYER M3 ;
        RECT 40.416 13.74 40.448 16.248 ;
  LAYER M3 ;
        RECT 40.48 13.74 40.512 16.248 ;
  LAYER M3 ;
        RECT 40.544 13.74 40.576 16.248 ;
  LAYER M3 ;
        RECT 40.608 13.74 40.64 16.248 ;
  LAYER M3 ;
        RECT 40.672 13.74 40.704 16.248 ;
  LAYER M3 ;
        RECT 40.736 13.74 40.768 16.248 ;
  LAYER M3 ;
        RECT 40.8 13.74 40.832 16.248 ;
  LAYER M3 ;
        RECT 40.864 13.74 40.896 16.248 ;
  LAYER M3 ;
        RECT 40.928 13.74 40.96 16.248 ;
  LAYER M3 ;
        RECT 40.992 13.74 41.024 16.248 ;
  LAYER M3 ;
        RECT 41.056 13.74 41.088 16.248 ;
  LAYER M3 ;
        RECT 41.12 13.74 41.152 16.248 ;
  LAYER M3 ;
        RECT 41.184 13.74 41.216 16.248 ;
  LAYER M3 ;
        RECT 41.248 13.74 41.28 16.248 ;
  LAYER M3 ;
        RECT 41.312 13.74 41.344 16.248 ;
  LAYER M3 ;
        RECT 41.376 13.74 41.408 16.248 ;
  LAYER M3 ;
        RECT 41.44 13.74 41.472 16.248 ;
  LAYER M3 ;
        RECT 41.504 13.74 41.536 16.248 ;
  LAYER M3 ;
        RECT 41.568 13.74 41.6 16.248 ;
  LAYER M3 ;
        RECT 41.632 13.74 41.664 16.248 ;
  LAYER M3 ;
        RECT 41.696 13.74 41.728 16.248 ;
  LAYER M3 ;
        RECT 41.76 13.74 41.792 16.248 ;
  LAYER M3 ;
        RECT 41.824 13.74 41.856 16.248 ;
  LAYER M3 ;
        RECT 41.888 13.74 41.92 16.248 ;
  LAYER M3 ;
        RECT 41.952 13.74 41.984 16.248 ;
  LAYER M3 ;
        RECT 42.016 13.74 42.048 16.248 ;
  LAYER M3 ;
        RECT 42.08 13.74 42.112 16.248 ;
  LAYER M3 ;
        RECT 42.144 13.74 42.176 16.248 ;
  LAYER M3 ;
        RECT 42.208 13.74 42.24 16.248 ;
  LAYER M3 ;
        RECT 42.272 13.74 42.304 16.248 ;
  LAYER M3 ;
        RECT 42.336 13.74 42.368 16.248 ;
  LAYER M3 ;
        RECT 42.4 13.74 42.432 16.248 ;
  LAYER M3 ;
        RECT 42.464 13.74 42.496 16.248 ;
  LAYER M3 ;
        RECT 42.528 13.74 42.56 16.248 ;
  LAYER M3 ;
        RECT 42.624 13.74 42.656 16.248 ;
  LAYER M1 ;
        RECT 40.239 13.776 40.241 16.212 ;
  LAYER M1 ;
        RECT 40.319 13.776 40.321 16.212 ;
  LAYER M1 ;
        RECT 40.399 13.776 40.401 16.212 ;
  LAYER M1 ;
        RECT 40.479 13.776 40.481 16.212 ;
  LAYER M1 ;
        RECT 40.559 13.776 40.561 16.212 ;
  LAYER M1 ;
        RECT 40.639 13.776 40.641 16.212 ;
  LAYER M1 ;
        RECT 40.719 13.776 40.721 16.212 ;
  LAYER M1 ;
        RECT 40.799 13.776 40.801 16.212 ;
  LAYER M1 ;
        RECT 40.879 13.776 40.881 16.212 ;
  LAYER M1 ;
        RECT 40.959 13.776 40.961 16.212 ;
  LAYER M1 ;
        RECT 41.039 13.776 41.041 16.212 ;
  LAYER M1 ;
        RECT 41.119 13.776 41.121 16.212 ;
  LAYER M1 ;
        RECT 41.199 13.776 41.201 16.212 ;
  LAYER M1 ;
        RECT 41.279 13.776 41.281 16.212 ;
  LAYER M1 ;
        RECT 41.359 13.776 41.361 16.212 ;
  LAYER M1 ;
        RECT 41.439 13.776 41.441 16.212 ;
  LAYER M1 ;
        RECT 41.519 13.776 41.521 16.212 ;
  LAYER M1 ;
        RECT 41.599 13.776 41.601 16.212 ;
  LAYER M1 ;
        RECT 41.679 13.776 41.681 16.212 ;
  LAYER M1 ;
        RECT 41.759 13.776 41.761 16.212 ;
  LAYER M1 ;
        RECT 41.839 13.776 41.841 16.212 ;
  LAYER M1 ;
        RECT 41.919 13.776 41.921 16.212 ;
  LAYER M1 ;
        RECT 41.999 13.776 42.001 16.212 ;
  LAYER M1 ;
        RECT 42.079 13.776 42.081 16.212 ;
  LAYER M1 ;
        RECT 42.159 13.776 42.161 16.212 ;
  LAYER M1 ;
        RECT 42.239 13.776 42.241 16.212 ;
  LAYER M1 ;
        RECT 42.319 13.776 42.321 16.212 ;
  LAYER M1 ;
        RECT 42.399 13.776 42.401 16.212 ;
  LAYER M1 ;
        RECT 42.479 13.776 42.481 16.212 ;
  LAYER M1 ;
        RECT 42.559 13.776 42.561 16.212 ;
  LAYER M2 ;
        RECT 40.24 16.211 42.64 16.213 ;
  LAYER M2 ;
        RECT 40.24 16.127 42.64 16.129 ;
  LAYER M2 ;
        RECT 40.24 16.043 42.64 16.045 ;
  LAYER M2 ;
        RECT 40.24 15.959 42.64 15.961 ;
  LAYER M2 ;
        RECT 40.24 15.875 42.64 15.877 ;
  LAYER M2 ;
        RECT 40.24 15.791 42.64 15.793 ;
  LAYER M2 ;
        RECT 40.24 15.707 42.64 15.709 ;
  LAYER M2 ;
        RECT 40.24 15.623 42.64 15.625 ;
  LAYER M2 ;
        RECT 40.24 15.539 42.64 15.541 ;
  LAYER M2 ;
        RECT 40.24 15.455 42.64 15.457 ;
  LAYER M2 ;
        RECT 40.24 15.371 42.64 15.373 ;
  LAYER M2 ;
        RECT 40.24 15.287 42.64 15.289 ;
  LAYER M2 ;
        RECT 40.24 15.2035 42.64 15.2055 ;
  LAYER M2 ;
        RECT 40.24 15.119 42.64 15.121 ;
  LAYER M2 ;
        RECT 40.24 15.035 42.64 15.037 ;
  LAYER M2 ;
        RECT 40.24 14.951 42.64 14.953 ;
  LAYER M2 ;
        RECT 40.24 14.867 42.64 14.869 ;
  LAYER M2 ;
        RECT 40.24 14.783 42.64 14.785 ;
  LAYER M2 ;
        RECT 40.24 14.699 42.64 14.701 ;
  LAYER M2 ;
        RECT 40.24 14.615 42.64 14.617 ;
  LAYER M2 ;
        RECT 40.24 14.531 42.64 14.533 ;
  LAYER M2 ;
        RECT 40.24 14.447 42.64 14.449 ;
  LAYER M2 ;
        RECT 40.24 14.363 42.64 14.365 ;
  LAYER M2 ;
        RECT 40.24 14.279 42.64 14.281 ;
  LAYER M2 ;
        RECT 40.24 14.195 42.64 14.197 ;
  LAYER M2 ;
        RECT 40.24 14.111 42.64 14.113 ;
  LAYER M2 ;
        RECT 40.24 14.027 42.64 14.029 ;
  LAYER M2 ;
        RECT 40.24 13.943 42.64 13.945 ;
  LAYER M2 ;
        RECT 40.24 13.859 42.64 13.861 ;
  LAYER M1 ;
        RECT 40.224 10.8 40.256 13.308 ;
  LAYER M1 ;
        RECT 40.288 10.8 40.32 13.308 ;
  LAYER M1 ;
        RECT 40.352 10.8 40.384 13.308 ;
  LAYER M1 ;
        RECT 40.416 10.8 40.448 13.308 ;
  LAYER M1 ;
        RECT 40.48 10.8 40.512 13.308 ;
  LAYER M1 ;
        RECT 40.544 10.8 40.576 13.308 ;
  LAYER M1 ;
        RECT 40.608 10.8 40.64 13.308 ;
  LAYER M1 ;
        RECT 40.672 10.8 40.704 13.308 ;
  LAYER M1 ;
        RECT 40.736 10.8 40.768 13.308 ;
  LAYER M1 ;
        RECT 40.8 10.8 40.832 13.308 ;
  LAYER M1 ;
        RECT 40.864 10.8 40.896 13.308 ;
  LAYER M1 ;
        RECT 40.928 10.8 40.96 13.308 ;
  LAYER M1 ;
        RECT 40.992 10.8 41.024 13.308 ;
  LAYER M1 ;
        RECT 41.056 10.8 41.088 13.308 ;
  LAYER M1 ;
        RECT 41.12 10.8 41.152 13.308 ;
  LAYER M1 ;
        RECT 41.184 10.8 41.216 13.308 ;
  LAYER M1 ;
        RECT 41.248 10.8 41.28 13.308 ;
  LAYER M1 ;
        RECT 41.312 10.8 41.344 13.308 ;
  LAYER M1 ;
        RECT 41.376 10.8 41.408 13.308 ;
  LAYER M1 ;
        RECT 41.44 10.8 41.472 13.308 ;
  LAYER M1 ;
        RECT 41.504 10.8 41.536 13.308 ;
  LAYER M1 ;
        RECT 41.568 10.8 41.6 13.308 ;
  LAYER M1 ;
        RECT 41.632 10.8 41.664 13.308 ;
  LAYER M1 ;
        RECT 41.696 10.8 41.728 13.308 ;
  LAYER M1 ;
        RECT 41.76 10.8 41.792 13.308 ;
  LAYER M1 ;
        RECT 41.824 10.8 41.856 13.308 ;
  LAYER M1 ;
        RECT 41.888 10.8 41.92 13.308 ;
  LAYER M1 ;
        RECT 41.952 10.8 41.984 13.308 ;
  LAYER M1 ;
        RECT 42.016 10.8 42.048 13.308 ;
  LAYER M1 ;
        RECT 42.08 10.8 42.112 13.308 ;
  LAYER M1 ;
        RECT 42.144 10.8 42.176 13.308 ;
  LAYER M1 ;
        RECT 42.208 10.8 42.24 13.308 ;
  LAYER M1 ;
        RECT 42.272 10.8 42.304 13.308 ;
  LAYER M1 ;
        RECT 42.336 10.8 42.368 13.308 ;
  LAYER M1 ;
        RECT 42.4 10.8 42.432 13.308 ;
  LAYER M1 ;
        RECT 42.464 10.8 42.496 13.308 ;
  LAYER M1 ;
        RECT 42.528 10.8 42.56 13.308 ;
  LAYER M2 ;
        RECT 40.204 13.192 42.676 13.224 ;
  LAYER M2 ;
        RECT 40.204 13.128 42.676 13.16 ;
  LAYER M2 ;
        RECT 40.204 13.064 42.676 13.096 ;
  LAYER M2 ;
        RECT 40.204 13 42.676 13.032 ;
  LAYER M2 ;
        RECT 40.204 12.936 42.676 12.968 ;
  LAYER M2 ;
        RECT 40.204 12.872 42.676 12.904 ;
  LAYER M2 ;
        RECT 40.204 12.808 42.676 12.84 ;
  LAYER M2 ;
        RECT 40.204 12.744 42.676 12.776 ;
  LAYER M2 ;
        RECT 40.204 12.68 42.676 12.712 ;
  LAYER M2 ;
        RECT 40.204 12.616 42.676 12.648 ;
  LAYER M2 ;
        RECT 40.204 12.552 42.676 12.584 ;
  LAYER M2 ;
        RECT 40.204 12.488 42.676 12.52 ;
  LAYER M2 ;
        RECT 40.204 12.424 42.676 12.456 ;
  LAYER M2 ;
        RECT 40.204 12.36 42.676 12.392 ;
  LAYER M2 ;
        RECT 40.204 12.296 42.676 12.328 ;
  LAYER M2 ;
        RECT 40.204 12.232 42.676 12.264 ;
  LAYER M2 ;
        RECT 40.204 12.168 42.676 12.2 ;
  LAYER M2 ;
        RECT 40.204 12.104 42.676 12.136 ;
  LAYER M2 ;
        RECT 40.204 12.04 42.676 12.072 ;
  LAYER M2 ;
        RECT 40.204 11.976 42.676 12.008 ;
  LAYER M2 ;
        RECT 40.204 11.912 42.676 11.944 ;
  LAYER M2 ;
        RECT 40.204 11.848 42.676 11.88 ;
  LAYER M2 ;
        RECT 40.204 11.784 42.676 11.816 ;
  LAYER M2 ;
        RECT 40.204 11.72 42.676 11.752 ;
  LAYER M2 ;
        RECT 40.204 11.656 42.676 11.688 ;
  LAYER M2 ;
        RECT 40.204 11.592 42.676 11.624 ;
  LAYER M2 ;
        RECT 40.204 11.528 42.676 11.56 ;
  LAYER M2 ;
        RECT 40.204 11.464 42.676 11.496 ;
  LAYER M2 ;
        RECT 40.204 11.4 42.676 11.432 ;
  LAYER M2 ;
        RECT 40.204 11.336 42.676 11.368 ;
  LAYER M2 ;
        RECT 40.204 11.272 42.676 11.304 ;
  LAYER M2 ;
        RECT 40.204 11.208 42.676 11.24 ;
  LAYER M2 ;
        RECT 40.204 11.144 42.676 11.176 ;
  LAYER M2 ;
        RECT 40.204 11.08 42.676 11.112 ;
  LAYER M2 ;
        RECT 40.204 11.016 42.676 11.048 ;
  LAYER M2 ;
        RECT 40.204 10.952 42.676 10.984 ;
  LAYER M3 ;
        RECT 40.224 10.8 40.256 13.308 ;
  LAYER M3 ;
        RECT 40.288 10.8 40.32 13.308 ;
  LAYER M3 ;
        RECT 40.352 10.8 40.384 13.308 ;
  LAYER M3 ;
        RECT 40.416 10.8 40.448 13.308 ;
  LAYER M3 ;
        RECT 40.48 10.8 40.512 13.308 ;
  LAYER M3 ;
        RECT 40.544 10.8 40.576 13.308 ;
  LAYER M3 ;
        RECT 40.608 10.8 40.64 13.308 ;
  LAYER M3 ;
        RECT 40.672 10.8 40.704 13.308 ;
  LAYER M3 ;
        RECT 40.736 10.8 40.768 13.308 ;
  LAYER M3 ;
        RECT 40.8 10.8 40.832 13.308 ;
  LAYER M3 ;
        RECT 40.864 10.8 40.896 13.308 ;
  LAYER M3 ;
        RECT 40.928 10.8 40.96 13.308 ;
  LAYER M3 ;
        RECT 40.992 10.8 41.024 13.308 ;
  LAYER M3 ;
        RECT 41.056 10.8 41.088 13.308 ;
  LAYER M3 ;
        RECT 41.12 10.8 41.152 13.308 ;
  LAYER M3 ;
        RECT 41.184 10.8 41.216 13.308 ;
  LAYER M3 ;
        RECT 41.248 10.8 41.28 13.308 ;
  LAYER M3 ;
        RECT 41.312 10.8 41.344 13.308 ;
  LAYER M3 ;
        RECT 41.376 10.8 41.408 13.308 ;
  LAYER M3 ;
        RECT 41.44 10.8 41.472 13.308 ;
  LAYER M3 ;
        RECT 41.504 10.8 41.536 13.308 ;
  LAYER M3 ;
        RECT 41.568 10.8 41.6 13.308 ;
  LAYER M3 ;
        RECT 41.632 10.8 41.664 13.308 ;
  LAYER M3 ;
        RECT 41.696 10.8 41.728 13.308 ;
  LAYER M3 ;
        RECT 41.76 10.8 41.792 13.308 ;
  LAYER M3 ;
        RECT 41.824 10.8 41.856 13.308 ;
  LAYER M3 ;
        RECT 41.888 10.8 41.92 13.308 ;
  LAYER M3 ;
        RECT 41.952 10.8 41.984 13.308 ;
  LAYER M3 ;
        RECT 42.016 10.8 42.048 13.308 ;
  LAYER M3 ;
        RECT 42.08 10.8 42.112 13.308 ;
  LAYER M3 ;
        RECT 42.144 10.8 42.176 13.308 ;
  LAYER M3 ;
        RECT 42.208 10.8 42.24 13.308 ;
  LAYER M3 ;
        RECT 42.272 10.8 42.304 13.308 ;
  LAYER M3 ;
        RECT 42.336 10.8 42.368 13.308 ;
  LAYER M3 ;
        RECT 42.4 10.8 42.432 13.308 ;
  LAYER M3 ;
        RECT 42.464 10.8 42.496 13.308 ;
  LAYER M3 ;
        RECT 42.528 10.8 42.56 13.308 ;
  LAYER M3 ;
        RECT 42.624 10.8 42.656 13.308 ;
  LAYER M1 ;
        RECT 40.239 10.836 40.241 13.272 ;
  LAYER M1 ;
        RECT 40.319 10.836 40.321 13.272 ;
  LAYER M1 ;
        RECT 40.399 10.836 40.401 13.272 ;
  LAYER M1 ;
        RECT 40.479 10.836 40.481 13.272 ;
  LAYER M1 ;
        RECT 40.559 10.836 40.561 13.272 ;
  LAYER M1 ;
        RECT 40.639 10.836 40.641 13.272 ;
  LAYER M1 ;
        RECT 40.719 10.836 40.721 13.272 ;
  LAYER M1 ;
        RECT 40.799 10.836 40.801 13.272 ;
  LAYER M1 ;
        RECT 40.879 10.836 40.881 13.272 ;
  LAYER M1 ;
        RECT 40.959 10.836 40.961 13.272 ;
  LAYER M1 ;
        RECT 41.039 10.836 41.041 13.272 ;
  LAYER M1 ;
        RECT 41.119 10.836 41.121 13.272 ;
  LAYER M1 ;
        RECT 41.199 10.836 41.201 13.272 ;
  LAYER M1 ;
        RECT 41.279 10.836 41.281 13.272 ;
  LAYER M1 ;
        RECT 41.359 10.836 41.361 13.272 ;
  LAYER M1 ;
        RECT 41.439 10.836 41.441 13.272 ;
  LAYER M1 ;
        RECT 41.519 10.836 41.521 13.272 ;
  LAYER M1 ;
        RECT 41.599 10.836 41.601 13.272 ;
  LAYER M1 ;
        RECT 41.679 10.836 41.681 13.272 ;
  LAYER M1 ;
        RECT 41.759 10.836 41.761 13.272 ;
  LAYER M1 ;
        RECT 41.839 10.836 41.841 13.272 ;
  LAYER M1 ;
        RECT 41.919 10.836 41.921 13.272 ;
  LAYER M1 ;
        RECT 41.999 10.836 42.001 13.272 ;
  LAYER M1 ;
        RECT 42.079 10.836 42.081 13.272 ;
  LAYER M1 ;
        RECT 42.159 10.836 42.161 13.272 ;
  LAYER M1 ;
        RECT 42.239 10.836 42.241 13.272 ;
  LAYER M1 ;
        RECT 42.319 10.836 42.321 13.272 ;
  LAYER M1 ;
        RECT 42.399 10.836 42.401 13.272 ;
  LAYER M1 ;
        RECT 42.479 10.836 42.481 13.272 ;
  LAYER M1 ;
        RECT 42.559 10.836 42.561 13.272 ;
  LAYER M2 ;
        RECT 40.24 13.271 42.64 13.273 ;
  LAYER M2 ;
        RECT 40.24 13.187 42.64 13.189 ;
  LAYER M2 ;
        RECT 40.24 13.103 42.64 13.105 ;
  LAYER M2 ;
        RECT 40.24 13.019 42.64 13.021 ;
  LAYER M2 ;
        RECT 40.24 12.935 42.64 12.937 ;
  LAYER M2 ;
        RECT 40.24 12.851 42.64 12.853 ;
  LAYER M2 ;
        RECT 40.24 12.767 42.64 12.769 ;
  LAYER M2 ;
        RECT 40.24 12.683 42.64 12.685 ;
  LAYER M2 ;
        RECT 40.24 12.599 42.64 12.601 ;
  LAYER M2 ;
        RECT 40.24 12.515 42.64 12.517 ;
  LAYER M2 ;
        RECT 40.24 12.431 42.64 12.433 ;
  LAYER M2 ;
        RECT 40.24 12.347 42.64 12.349 ;
  LAYER M2 ;
        RECT 40.24 12.2635 42.64 12.2655 ;
  LAYER M2 ;
        RECT 40.24 12.179 42.64 12.181 ;
  LAYER M2 ;
        RECT 40.24 12.095 42.64 12.097 ;
  LAYER M2 ;
        RECT 40.24 12.011 42.64 12.013 ;
  LAYER M2 ;
        RECT 40.24 11.927 42.64 11.929 ;
  LAYER M2 ;
        RECT 40.24 11.843 42.64 11.845 ;
  LAYER M2 ;
        RECT 40.24 11.759 42.64 11.761 ;
  LAYER M2 ;
        RECT 40.24 11.675 42.64 11.677 ;
  LAYER M2 ;
        RECT 40.24 11.591 42.64 11.593 ;
  LAYER M2 ;
        RECT 40.24 11.507 42.64 11.509 ;
  LAYER M2 ;
        RECT 40.24 11.423 42.64 11.425 ;
  LAYER M2 ;
        RECT 40.24 11.339 42.64 11.341 ;
  LAYER M2 ;
        RECT 40.24 11.255 42.64 11.257 ;
  LAYER M2 ;
        RECT 40.24 11.171 42.64 11.173 ;
  LAYER M2 ;
        RECT 40.24 11.087 42.64 11.089 ;
  LAYER M2 ;
        RECT 40.24 11.003 42.64 11.005 ;
  LAYER M2 ;
        RECT 40.24 10.919 42.64 10.921 ;
  LAYER M1 ;
        RECT 40.224 7.86 40.256 10.368 ;
  LAYER M1 ;
        RECT 40.288 7.86 40.32 10.368 ;
  LAYER M1 ;
        RECT 40.352 7.86 40.384 10.368 ;
  LAYER M1 ;
        RECT 40.416 7.86 40.448 10.368 ;
  LAYER M1 ;
        RECT 40.48 7.86 40.512 10.368 ;
  LAYER M1 ;
        RECT 40.544 7.86 40.576 10.368 ;
  LAYER M1 ;
        RECT 40.608 7.86 40.64 10.368 ;
  LAYER M1 ;
        RECT 40.672 7.86 40.704 10.368 ;
  LAYER M1 ;
        RECT 40.736 7.86 40.768 10.368 ;
  LAYER M1 ;
        RECT 40.8 7.86 40.832 10.368 ;
  LAYER M1 ;
        RECT 40.864 7.86 40.896 10.368 ;
  LAYER M1 ;
        RECT 40.928 7.86 40.96 10.368 ;
  LAYER M1 ;
        RECT 40.992 7.86 41.024 10.368 ;
  LAYER M1 ;
        RECT 41.056 7.86 41.088 10.368 ;
  LAYER M1 ;
        RECT 41.12 7.86 41.152 10.368 ;
  LAYER M1 ;
        RECT 41.184 7.86 41.216 10.368 ;
  LAYER M1 ;
        RECT 41.248 7.86 41.28 10.368 ;
  LAYER M1 ;
        RECT 41.312 7.86 41.344 10.368 ;
  LAYER M1 ;
        RECT 41.376 7.86 41.408 10.368 ;
  LAYER M1 ;
        RECT 41.44 7.86 41.472 10.368 ;
  LAYER M1 ;
        RECT 41.504 7.86 41.536 10.368 ;
  LAYER M1 ;
        RECT 41.568 7.86 41.6 10.368 ;
  LAYER M1 ;
        RECT 41.632 7.86 41.664 10.368 ;
  LAYER M1 ;
        RECT 41.696 7.86 41.728 10.368 ;
  LAYER M1 ;
        RECT 41.76 7.86 41.792 10.368 ;
  LAYER M1 ;
        RECT 41.824 7.86 41.856 10.368 ;
  LAYER M1 ;
        RECT 41.888 7.86 41.92 10.368 ;
  LAYER M1 ;
        RECT 41.952 7.86 41.984 10.368 ;
  LAYER M1 ;
        RECT 42.016 7.86 42.048 10.368 ;
  LAYER M1 ;
        RECT 42.08 7.86 42.112 10.368 ;
  LAYER M1 ;
        RECT 42.144 7.86 42.176 10.368 ;
  LAYER M1 ;
        RECT 42.208 7.86 42.24 10.368 ;
  LAYER M1 ;
        RECT 42.272 7.86 42.304 10.368 ;
  LAYER M1 ;
        RECT 42.336 7.86 42.368 10.368 ;
  LAYER M1 ;
        RECT 42.4 7.86 42.432 10.368 ;
  LAYER M1 ;
        RECT 42.464 7.86 42.496 10.368 ;
  LAYER M1 ;
        RECT 42.528 7.86 42.56 10.368 ;
  LAYER M2 ;
        RECT 40.204 10.252 42.676 10.284 ;
  LAYER M2 ;
        RECT 40.204 10.188 42.676 10.22 ;
  LAYER M2 ;
        RECT 40.204 10.124 42.676 10.156 ;
  LAYER M2 ;
        RECT 40.204 10.06 42.676 10.092 ;
  LAYER M2 ;
        RECT 40.204 9.996 42.676 10.028 ;
  LAYER M2 ;
        RECT 40.204 9.932 42.676 9.964 ;
  LAYER M2 ;
        RECT 40.204 9.868 42.676 9.9 ;
  LAYER M2 ;
        RECT 40.204 9.804 42.676 9.836 ;
  LAYER M2 ;
        RECT 40.204 9.74 42.676 9.772 ;
  LAYER M2 ;
        RECT 40.204 9.676 42.676 9.708 ;
  LAYER M2 ;
        RECT 40.204 9.612 42.676 9.644 ;
  LAYER M2 ;
        RECT 40.204 9.548 42.676 9.58 ;
  LAYER M2 ;
        RECT 40.204 9.484 42.676 9.516 ;
  LAYER M2 ;
        RECT 40.204 9.42 42.676 9.452 ;
  LAYER M2 ;
        RECT 40.204 9.356 42.676 9.388 ;
  LAYER M2 ;
        RECT 40.204 9.292 42.676 9.324 ;
  LAYER M2 ;
        RECT 40.204 9.228 42.676 9.26 ;
  LAYER M2 ;
        RECT 40.204 9.164 42.676 9.196 ;
  LAYER M2 ;
        RECT 40.204 9.1 42.676 9.132 ;
  LAYER M2 ;
        RECT 40.204 9.036 42.676 9.068 ;
  LAYER M2 ;
        RECT 40.204 8.972 42.676 9.004 ;
  LAYER M2 ;
        RECT 40.204 8.908 42.676 8.94 ;
  LAYER M2 ;
        RECT 40.204 8.844 42.676 8.876 ;
  LAYER M2 ;
        RECT 40.204 8.78 42.676 8.812 ;
  LAYER M2 ;
        RECT 40.204 8.716 42.676 8.748 ;
  LAYER M2 ;
        RECT 40.204 8.652 42.676 8.684 ;
  LAYER M2 ;
        RECT 40.204 8.588 42.676 8.62 ;
  LAYER M2 ;
        RECT 40.204 8.524 42.676 8.556 ;
  LAYER M2 ;
        RECT 40.204 8.46 42.676 8.492 ;
  LAYER M2 ;
        RECT 40.204 8.396 42.676 8.428 ;
  LAYER M2 ;
        RECT 40.204 8.332 42.676 8.364 ;
  LAYER M2 ;
        RECT 40.204 8.268 42.676 8.3 ;
  LAYER M2 ;
        RECT 40.204 8.204 42.676 8.236 ;
  LAYER M2 ;
        RECT 40.204 8.14 42.676 8.172 ;
  LAYER M2 ;
        RECT 40.204 8.076 42.676 8.108 ;
  LAYER M2 ;
        RECT 40.204 8.012 42.676 8.044 ;
  LAYER M3 ;
        RECT 40.224 7.86 40.256 10.368 ;
  LAYER M3 ;
        RECT 40.288 7.86 40.32 10.368 ;
  LAYER M3 ;
        RECT 40.352 7.86 40.384 10.368 ;
  LAYER M3 ;
        RECT 40.416 7.86 40.448 10.368 ;
  LAYER M3 ;
        RECT 40.48 7.86 40.512 10.368 ;
  LAYER M3 ;
        RECT 40.544 7.86 40.576 10.368 ;
  LAYER M3 ;
        RECT 40.608 7.86 40.64 10.368 ;
  LAYER M3 ;
        RECT 40.672 7.86 40.704 10.368 ;
  LAYER M3 ;
        RECT 40.736 7.86 40.768 10.368 ;
  LAYER M3 ;
        RECT 40.8 7.86 40.832 10.368 ;
  LAYER M3 ;
        RECT 40.864 7.86 40.896 10.368 ;
  LAYER M3 ;
        RECT 40.928 7.86 40.96 10.368 ;
  LAYER M3 ;
        RECT 40.992 7.86 41.024 10.368 ;
  LAYER M3 ;
        RECT 41.056 7.86 41.088 10.368 ;
  LAYER M3 ;
        RECT 41.12 7.86 41.152 10.368 ;
  LAYER M3 ;
        RECT 41.184 7.86 41.216 10.368 ;
  LAYER M3 ;
        RECT 41.248 7.86 41.28 10.368 ;
  LAYER M3 ;
        RECT 41.312 7.86 41.344 10.368 ;
  LAYER M3 ;
        RECT 41.376 7.86 41.408 10.368 ;
  LAYER M3 ;
        RECT 41.44 7.86 41.472 10.368 ;
  LAYER M3 ;
        RECT 41.504 7.86 41.536 10.368 ;
  LAYER M3 ;
        RECT 41.568 7.86 41.6 10.368 ;
  LAYER M3 ;
        RECT 41.632 7.86 41.664 10.368 ;
  LAYER M3 ;
        RECT 41.696 7.86 41.728 10.368 ;
  LAYER M3 ;
        RECT 41.76 7.86 41.792 10.368 ;
  LAYER M3 ;
        RECT 41.824 7.86 41.856 10.368 ;
  LAYER M3 ;
        RECT 41.888 7.86 41.92 10.368 ;
  LAYER M3 ;
        RECT 41.952 7.86 41.984 10.368 ;
  LAYER M3 ;
        RECT 42.016 7.86 42.048 10.368 ;
  LAYER M3 ;
        RECT 42.08 7.86 42.112 10.368 ;
  LAYER M3 ;
        RECT 42.144 7.86 42.176 10.368 ;
  LAYER M3 ;
        RECT 42.208 7.86 42.24 10.368 ;
  LAYER M3 ;
        RECT 42.272 7.86 42.304 10.368 ;
  LAYER M3 ;
        RECT 42.336 7.86 42.368 10.368 ;
  LAYER M3 ;
        RECT 42.4 7.86 42.432 10.368 ;
  LAYER M3 ;
        RECT 42.464 7.86 42.496 10.368 ;
  LAYER M3 ;
        RECT 42.528 7.86 42.56 10.368 ;
  LAYER M3 ;
        RECT 42.624 7.86 42.656 10.368 ;
  LAYER M1 ;
        RECT 40.239 7.896 40.241 10.332 ;
  LAYER M1 ;
        RECT 40.319 7.896 40.321 10.332 ;
  LAYER M1 ;
        RECT 40.399 7.896 40.401 10.332 ;
  LAYER M1 ;
        RECT 40.479 7.896 40.481 10.332 ;
  LAYER M1 ;
        RECT 40.559 7.896 40.561 10.332 ;
  LAYER M1 ;
        RECT 40.639 7.896 40.641 10.332 ;
  LAYER M1 ;
        RECT 40.719 7.896 40.721 10.332 ;
  LAYER M1 ;
        RECT 40.799 7.896 40.801 10.332 ;
  LAYER M1 ;
        RECT 40.879 7.896 40.881 10.332 ;
  LAYER M1 ;
        RECT 40.959 7.896 40.961 10.332 ;
  LAYER M1 ;
        RECT 41.039 7.896 41.041 10.332 ;
  LAYER M1 ;
        RECT 41.119 7.896 41.121 10.332 ;
  LAYER M1 ;
        RECT 41.199 7.896 41.201 10.332 ;
  LAYER M1 ;
        RECT 41.279 7.896 41.281 10.332 ;
  LAYER M1 ;
        RECT 41.359 7.896 41.361 10.332 ;
  LAYER M1 ;
        RECT 41.439 7.896 41.441 10.332 ;
  LAYER M1 ;
        RECT 41.519 7.896 41.521 10.332 ;
  LAYER M1 ;
        RECT 41.599 7.896 41.601 10.332 ;
  LAYER M1 ;
        RECT 41.679 7.896 41.681 10.332 ;
  LAYER M1 ;
        RECT 41.759 7.896 41.761 10.332 ;
  LAYER M1 ;
        RECT 41.839 7.896 41.841 10.332 ;
  LAYER M1 ;
        RECT 41.919 7.896 41.921 10.332 ;
  LAYER M1 ;
        RECT 41.999 7.896 42.001 10.332 ;
  LAYER M1 ;
        RECT 42.079 7.896 42.081 10.332 ;
  LAYER M1 ;
        RECT 42.159 7.896 42.161 10.332 ;
  LAYER M1 ;
        RECT 42.239 7.896 42.241 10.332 ;
  LAYER M1 ;
        RECT 42.319 7.896 42.321 10.332 ;
  LAYER M1 ;
        RECT 42.399 7.896 42.401 10.332 ;
  LAYER M1 ;
        RECT 42.479 7.896 42.481 10.332 ;
  LAYER M1 ;
        RECT 42.559 7.896 42.561 10.332 ;
  LAYER M2 ;
        RECT 40.24 10.331 42.64 10.333 ;
  LAYER M2 ;
        RECT 40.24 10.247 42.64 10.249 ;
  LAYER M2 ;
        RECT 40.24 10.163 42.64 10.165 ;
  LAYER M2 ;
        RECT 40.24 10.079 42.64 10.081 ;
  LAYER M2 ;
        RECT 40.24 9.995 42.64 9.997 ;
  LAYER M2 ;
        RECT 40.24 9.911 42.64 9.913 ;
  LAYER M2 ;
        RECT 40.24 9.827 42.64 9.829 ;
  LAYER M2 ;
        RECT 40.24 9.743 42.64 9.745 ;
  LAYER M2 ;
        RECT 40.24 9.659 42.64 9.661 ;
  LAYER M2 ;
        RECT 40.24 9.575 42.64 9.577 ;
  LAYER M2 ;
        RECT 40.24 9.491 42.64 9.493 ;
  LAYER M2 ;
        RECT 40.24 9.407 42.64 9.409 ;
  LAYER M2 ;
        RECT 40.24 9.3235 42.64 9.3255 ;
  LAYER M2 ;
        RECT 40.24 9.239 42.64 9.241 ;
  LAYER M2 ;
        RECT 40.24 9.155 42.64 9.157 ;
  LAYER M2 ;
        RECT 40.24 9.071 42.64 9.073 ;
  LAYER M2 ;
        RECT 40.24 8.987 42.64 8.989 ;
  LAYER M2 ;
        RECT 40.24 8.903 42.64 8.905 ;
  LAYER M2 ;
        RECT 40.24 8.819 42.64 8.821 ;
  LAYER M2 ;
        RECT 40.24 8.735 42.64 8.737 ;
  LAYER M2 ;
        RECT 40.24 8.651 42.64 8.653 ;
  LAYER M2 ;
        RECT 40.24 8.567 42.64 8.569 ;
  LAYER M2 ;
        RECT 40.24 8.483 42.64 8.485 ;
  LAYER M2 ;
        RECT 40.24 8.399 42.64 8.401 ;
  LAYER M2 ;
        RECT 40.24 8.315 42.64 8.317 ;
  LAYER M2 ;
        RECT 40.24 8.231 42.64 8.233 ;
  LAYER M2 ;
        RECT 40.24 8.147 42.64 8.149 ;
  LAYER M2 ;
        RECT 40.24 8.063 42.64 8.065 ;
  LAYER M2 ;
        RECT 40.24 7.979 42.64 7.981 ;
  LAYER M1 ;
        RECT 40.224 4.92 40.256 7.428 ;
  LAYER M1 ;
        RECT 40.288 4.92 40.32 7.428 ;
  LAYER M1 ;
        RECT 40.352 4.92 40.384 7.428 ;
  LAYER M1 ;
        RECT 40.416 4.92 40.448 7.428 ;
  LAYER M1 ;
        RECT 40.48 4.92 40.512 7.428 ;
  LAYER M1 ;
        RECT 40.544 4.92 40.576 7.428 ;
  LAYER M1 ;
        RECT 40.608 4.92 40.64 7.428 ;
  LAYER M1 ;
        RECT 40.672 4.92 40.704 7.428 ;
  LAYER M1 ;
        RECT 40.736 4.92 40.768 7.428 ;
  LAYER M1 ;
        RECT 40.8 4.92 40.832 7.428 ;
  LAYER M1 ;
        RECT 40.864 4.92 40.896 7.428 ;
  LAYER M1 ;
        RECT 40.928 4.92 40.96 7.428 ;
  LAYER M1 ;
        RECT 40.992 4.92 41.024 7.428 ;
  LAYER M1 ;
        RECT 41.056 4.92 41.088 7.428 ;
  LAYER M1 ;
        RECT 41.12 4.92 41.152 7.428 ;
  LAYER M1 ;
        RECT 41.184 4.92 41.216 7.428 ;
  LAYER M1 ;
        RECT 41.248 4.92 41.28 7.428 ;
  LAYER M1 ;
        RECT 41.312 4.92 41.344 7.428 ;
  LAYER M1 ;
        RECT 41.376 4.92 41.408 7.428 ;
  LAYER M1 ;
        RECT 41.44 4.92 41.472 7.428 ;
  LAYER M1 ;
        RECT 41.504 4.92 41.536 7.428 ;
  LAYER M1 ;
        RECT 41.568 4.92 41.6 7.428 ;
  LAYER M1 ;
        RECT 41.632 4.92 41.664 7.428 ;
  LAYER M1 ;
        RECT 41.696 4.92 41.728 7.428 ;
  LAYER M1 ;
        RECT 41.76 4.92 41.792 7.428 ;
  LAYER M1 ;
        RECT 41.824 4.92 41.856 7.428 ;
  LAYER M1 ;
        RECT 41.888 4.92 41.92 7.428 ;
  LAYER M1 ;
        RECT 41.952 4.92 41.984 7.428 ;
  LAYER M1 ;
        RECT 42.016 4.92 42.048 7.428 ;
  LAYER M1 ;
        RECT 42.08 4.92 42.112 7.428 ;
  LAYER M1 ;
        RECT 42.144 4.92 42.176 7.428 ;
  LAYER M1 ;
        RECT 42.208 4.92 42.24 7.428 ;
  LAYER M1 ;
        RECT 42.272 4.92 42.304 7.428 ;
  LAYER M1 ;
        RECT 42.336 4.92 42.368 7.428 ;
  LAYER M1 ;
        RECT 42.4 4.92 42.432 7.428 ;
  LAYER M1 ;
        RECT 42.464 4.92 42.496 7.428 ;
  LAYER M1 ;
        RECT 42.528 4.92 42.56 7.428 ;
  LAYER M2 ;
        RECT 40.204 7.312 42.676 7.344 ;
  LAYER M2 ;
        RECT 40.204 7.248 42.676 7.28 ;
  LAYER M2 ;
        RECT 40.204 7.184 42.676 7.216 ;
  LAYER M2 ;
        RECT 40.204 7.12 42.676 7.152 ;
  LAYER M2 ;
        RECT 40.204 7.056 42.676 7.088 ;
  LAYER M2 ;
        RECT 40.204 6.992 42.676 7.024 ;
  LAYER M2 ;
        RECT 40.204 6.928 42.676 6.96 ;
  LAYER M2 ;
        RECT 40.204 6.864 42.676 6.896 ;
  LAYER M2 ;
        RECT 40.204 6.8 42.676 6.832 ;
  LAYER M2 ;
        RECT 40.204 6.736 42.676 6.768 ;
  LAYER M2 ;
        RECT 40.204 6.672 42.676 6.704 ;
  LAYER M2 ;
        RECT 40.204 6.608 42.676 6.64 ;
  LAYER M2 ;
        RECT 40.204 6.544 42.676 6.576 ;
  LAYER M2 ;
        RECT 40.204 6.48 42.676 6.512 ;
  LAYER M2 ;
        RECT 40.204 6.416 42.676 6.448 ;
  LAYER M2 ;
        RECT 40.204 6.352 42.676 6.384 ;
  LAYER M2 ;
        RECT 40.204 6.288 42.676 6.32 ;
  LAYER M2 ;
        RECT 40.204 6.224 42.676 6.256 ;
  LAYER M2 ;
        RECT 40.204 6.16 42.676 6.192 ;
  LAYER M2 ;
        RECT 40.204 6.096 42.676 6.128 ;
  LAYER M2 ;
        RECT 40.204 6.032 42.676 6.064 ;
  LAYER M2 ;
        RECT 40.204 5.968 42.676 6 ;
  LAYER M2 ;
        RECT 40.204 5.904 42.676 5.936 ;
  LAYER M2 ;
        RECT 40.204 5.84 42.676 5.872 ;
  LAYER M2 ;
        RECT 40.204 5.776 42.676 5.808 ;
  LAYER M2 ;
        RECT 40.204 5.712 42.676 5.744 ;
  LAYER M2 ;
        RECT 40.204 5.648 42.676 5.68 ;
  LAYER M2 ;
        RECT 40.204 5.584 42.676 5.616 ;
  LAYER M2 ;
        RECT 40.204 5.52 42.676 5.552 ;
  LAYER M2 ;
        RECT 40.204 5.456 42.676 5.488 ;
  LAYER M2 ;
        RECT 40.204 5.392 42.676 5.424 ;
  LAYER M2 ;
        RECT 40.204 5.328 42.676 5.36 ;
  LAYER M2 ;
        RECT 40.204 5.264 42.676 5.296 ;
  LAYER M2 ;
        RECT 40.204 5.2 42.676 5.232 ;
  LAYER M2 ;
        RECT 40.204 5.136 42.676 5.168 ;
  LAYER M2 ;
        RECT 40.204 5.072 42.676 5.104 ;
  LAYER M3 ;
        RECT 40.224 4.92 40.256 7.428 ;
  LAYER M3 ;
        RECT 40.288 4.92 40.32 7.428 ;
  LAYER M3 ;
        RECT 40.352 4.92 40.384 7.428 ;
  LAYER M3 ;
        RECT 40.416 4.92 40.448 7.428 ;
  LAYER M3 ;
        RECT 40.48 4.92 40.512 7.428 ;
  LAYER M3 ;
        RECT 40.544 4.92 40.576 7.428 ;
  LAYER M3 ;
        RECT 40.608 4.92 40.64 7.428 ;
  LAYER M3 ;
        RECT 40.672 4.92 40.704 7.428 ;
  LAYER M3 ;
        RECT 40.736 4.92 40.768 7.428 ;
  LAYER M3 ;
        RECT 40.8 4.92 40.832 7.428 ;
  LAYER M3 ;
        RECT 40.864 4.92 40.896 7.428 ;
  LAYER M3 ;
        RECT 40.928 4.92 40.96 7.428 ;
  LAYER M3 ;
        RECT 40.992 4.92 41.024 7.428 ;
  LAYER M3 ;
        RECT 41.056 4.92 41.088 7.428 ;
  LAYER M3 ;
        RECT 41.12 4.92 41.152 7.428 ;
  LAYER M3 ;
        RECT 41.184 4.92 41.216 7.428 ;
  LAYER M3 ;
        RECT 41.248 4.92 41.28 7.428 ;
  LAYER M3 ;
        RECT 41.312 4.92 41.344 7.428 ;
  LAYER M3 ;
        RECT 41.376 4.92 41.408 7.428 ;
  LAYER M3 ;
        RECT 41.44 4.92 41.472 7.428 ;
  LAYER M3 ;
        RECT 41.504 4.92 41.536 7.428 ;
  LAYER M3 ;
        RECT 41.568 4.92 41.6 7.428 ;
  LAYER M3 ;
        RECT 41.632 4.92 41.664 7.428 ;
  LAYER M3 ;
        RECT 41.696 4.92 41.728 7.428 ;
  LAYER M3 ;
        RECT 41.76 4.92 41.792 7.428 ;
  LAYER M3 ;
        RECT 41.824 4.92 41.856 7.428 ;
  LAYER M3 ;
        RECT 41.888 4.92 41.92 7.428 ;
  LAYER M3 ;
        RECT 41.952 4.92 41.984 7.428 ;
  LAYER M3 ;
        RECT 42.016 4.92 42.048 7.428 ;
  LAYER M3 ;
        RECT 42.08 4.92 42.112 7.428 ;
  LAYER M3 ;
        RECT 42.144 4.92 42.176 7.428 ;
  LAYER M3 ;
        RECT 42.208 4.92 42.24 7.428 ;
  LAYER M3 ;
        RECT 42.272 4.92 42.304 7.428 ;
  LAYER M3 ;
        RECT 42.336 4.92 42.368 7.428 ;
  LAYER M3 ;
        RECT 42.4 4.92 42.432 7.428 ;
  LAYER M3 ;
        RECT 42.464 4.92 42.496 7.428 ;
  LAYER M3 ;
        RECT 42.528 4.92 42.56 7.428 ;
  LAYER M3 ;
        RECT 42.624 4.92 42.656 7.428 ;
  LAYER M1 ;
        RECT 40.239 4.956 40.241 7.392 ;
  LAYER M1 ;
        RECT 40.319 4.956 40.321 7.392 ;
  LAYER M1 ;
        RECT 40.399 4.956 40.401 7.392 ;
  LAYER M1 ;
        RECT 40.479 4.956 40.481 7.392 ;
  LAYER M1 ;
        RECT 40.559 4.956 40.561 7.392 ;
  LAYER M1 ;
        RECT 40.639 4.956 40.641 7.392 ;
  LAYER M1 ;
        RECT 40.719 4.956 40.721 7.392 ;
  LAYER M1 ;
        RECT 40.799 4.956 40.801 7.392 ;
  LAYER M1 ;
        RECT 40.879 4.956 40.881 7.392 ;
  LAYER M1 ;
        RECT 40.959 4.956 40.961 7.392 ;
  LAYER M1 ;
        RECT 41.039 4.956 41.041 7.392 ;
  LAYER M1 ;
        RECT 41.119 4.956 41.121 7.392 ;
  LAYER M1 ;
        RECT 41.199 4.956 41.201 7.392 ;
  LAYER M1 ;
        RECT 41.279 4.956 41.281 7.392 ;
  LAYER M1 ;
        RECT 41.359 4.956 41.361 7.392 ;
  LAYER M1 ;
        RECT 41.439 4.956 41.441 7.392 ;
  LAYER M1 ;
        RECT 41.519 4.956 41.521 7.392 ;
  LAYER M1 ;
        RECT 41.599 4.956 41.601 7.392 ;
  LAYER M1 ;
        RECT 41.679 4.956 41.681 7.392 ;
  LAYER M1 ;
        RECT 41.759 4.956 41.761 7.392 ;
  LAYER M1 ;
        RECT 41.839 4.956 41.841 7.392 ;
  LAYER M1 ;
        RECT 41.919 4.956 41.921 7.392 ;
  LAYER M1 ;
        RECT 41.999 4.956 42.001 7.392 ;
  LAYER M1 ;
        RECT 42.079 4.956 42.081 7.392 ;
  LAYER M1 ;
        RECT 42.159 4.956 42.161 7.392 ;
  LAYER M1 ;
        RECT 42.239 4.956 42.241 7.392 ;
  LAYER M1 ;
        RECT 42.319 4.956 42.321 7.392 ;
  LAYER M1 ;
        RECT 42.399 4.956 42.401 7.392 ;
  LAYER M1 ;
        RECT 42.479 4.956 42.481 7.392 ;
  LAYER M1 ;
        RECT 42.559 4.956 42.561 7.392 ;
  LAYER M2 ;
        RECT 40.24 7.391 42.64 7.393 ;
  LAYER M2 ;
        RECT 40.24 7.307 42.64 7.309 ;
  LAYER M2 ;
        RECT 40.24 7.223 42.64 7.225 ;
  LAYER M2 ;
        RECT 40.24 7.139 42.64 7.141 ;
  LAYER M2 ;
        RECT 40.24 7.055 42.64 7.057 ;
  LAYER M2 ;
        RECT 40.24 6.971 42.64 6.973 ;
  LAYER M2 ;
        RECT 40.24 6.887 42.64 6.889 ;
  LAYER M2 ;
        RECT 40.24 6.803 42.64 6.805 ;
  LAYER M2 ;
        RECT 40.24 6.719 42.64 6.721 ;
  LAYER M2 ;
        RECT 40.24 6.635 42.64 6.637 ;
  LAYER M2 ;
        RECT 40.24 6.551 42.64 6.553 ;
  LAYER M2 ;
        RECT 40.24 6.467 42.64 6.469 ;
  LAYER M2 ;
        RECT 40.24 6.3835 42.64 6.3855 ;
  LAYER M2 ;
        RECT 40.24 6.299 42.64 6.301 ;
  LAYER M2 ;
        RECT 40.24 6.215 42.64 6.217 ;
  LAYER M2 ;
        RECT 40.24 6.131 42.64 6.133 ;
  LAYER M2 ;
        RECT 40.24 6.047 42.64 6.049 ;
  LAYER M2 ;
        RECT 40.24 5.963 42.64 5.965 ;
  LAYER M2 ;
        RECT 40.24 5.879 42.64 5.881 ;
  LAYER M2 ;
        RECT 40.24 5.795 42.64 5.797 ;
  LAYER M2 ;
        RECT 40.24 5.711 42.64 5.713 ;
  LAYER M2 ;
        RECT 40.24 5.627 42.64 5.629 ;
  LAYER M2 ;
        RECT 40.24 5.543 42.64 5.545 ;
  LAYER M2 ;
        RECT 40.24 5.459 42.64 5.461 ;
  LAYER M2 ;
        RECT 40.24 5.375 42.64 5.377 ;
  LAYER M2 ;
        RECT 40.24 5.291 42.64 5.293 ;
  LAYER M2 ;
        RECT 40.24 5.207 42.64 5.209 ;
  LAYER M2 ;
        RECT 40.24 5.123 42.64 5.125 ;
  LAYER M2 ;
        RECT 40.24 5.039 42.64 5.041 ;
  LAYER M1 ;
        RECT 40.224 1.98 40.256 4.488 ;
  LAYER M1 ;
        RECT 40.288 1.98 40.32 4.488 ;
  LAYER M1 ;
        RECT 40.352 1.98 40.384 4.488 ;
  LAYER M1 ;
        RECT 40.416 1.98 40.448 4.488 ;
  LAYER M1 ;
        RECT 40.48 1.98 40.512 4.488 ;
  LAYER M1 ;
        RECT 40.544 1.98 40.576 4.488 ;
  LAYER M1 ;
        RECT 40.608 1.98 40.64 4.488 ;
  LAYER M1 ;
        RECT 40.672 1.98 40.704 4.488 ;
  LAYER M1 ;
        RECT 40.736 1.98 40.768 4.488 ;
  LAYER M1 ;
        RECT 40.8 1.98 40.832 4.488 ;
  LAYER M1 ;
        RECT 40.864 1.98 40.896 4.488 ;
  LAYER M1 ;
        RECT 40.928 1.98 40.96 4.488 ;
  LAYER M1 ;
        RECT 40.992 1.98 41.024 4.488 ;
  LAYER M1 ;
        RECT 41.056 1.98 41.088 4.488 ;
  LAYER M1 ;
        RECT 41.12 1.98 41.152 4.488 ;
  LAYER M1 ;
        RECT 41.184 1.98 41.216 4.488 ;
  LAYER M1 ;
        RECT 41.248 1.98 41.28 4.488 ;
  LAYER M1 ;
        RECT 41.312 1.98 41.344 4.488 ;
  LAYER M1 ;
        RECT 41.376 1.98 41.408 4.488 ;
  LAYER M1 ;
        RECT 41.44 1.98 41.472 4.488 ;
  LAYER M1 ;
        RECT 41.504 1.98 41.536 4.488 ;
  LAYER M1 ;
        RECT 41.568 1.98 41.6 4.488 ;
  LAYER M1 ;
        RECT 41.632 1.98 41.664 4.488 ;
  LAYER M1 ;
        RECT 41.696 1.98 41.728 4.488 ;
  LAYER M1 ;
        RECT 41.76 1.98 41.792 4.488 ;
  LAYER M1 ;
        RECT 41.824 1.98 41.856 4.488 ;
  LAYER M1 ;
        RECT 41.888 1.98 41.92 4.488 ;
  LAYER M1 ;
        RECT 41.952 1.98 41.984 4.488 ;
  LAYER M1 ;
        RECT 42.016 1.98 42.048 4.488 ;
  LAYER M1 ;
        RECT 42.08 1.98 42.112 4.488 ;
  LAYER M1 ;
        RECT 42.144 1.98 42.176 4.488 ;
  LAYER M1 ;
        RECT 42.208 1.98 42.24 4.488 ;
  LAYER M1 ;
        RECT 42.272 1.98 42.304 4.488 ;
  LAYER M1 ;
        RECT 42.336 1.98 42.368 4.488 ;
  LAYER M1 ;
        RECT 42.4 1.98 42.432 4.488 ;
  LAYER M1 ;
        RECT 42.464 1.98 42.496 4.488 ;
  LAYER M1 ;
        RECT 42.528 1.98 42.56 4.488 ;
  LAYER M2 ;
        RECT 40.204 4.372 42.676 4.404 ;
  LAYER M2 ;
        RECT 40.204 4.308 42.676 4.34 ;
  LAYER M2 ;
        RECT 40.204 4.244 42.676 4.276 ;
  LAYER M2 ;
        RECT 40.204 4.18 42.676 4.212 ;
  LAYER M2 ;
        RECT 40.204 4.116 42.676 4.148 ;
  LAYER M2 ;
        RECT 40.204 4.052 42.676 4.084 ;
  LAYER M2 ;
        RECT 40.204 3.988 42.676 4.02 ;
  LAYER M2 ;
        RECT 40.204 3.924 42.676 3.956 ;
  LAYER M2 ;
        RECT 40.204 3.86 42.676 3.892 ;
  LAYER M2 ;
        RECT 40.204 3.796 42.676 3.828 ;
  LAYER M2 ;
        RECT 40.204 3.732 42.676 3.764 ;
  LAYER M2 ;
        RECT 40.204 3.668 42.676 3.7 ;
  LAYER M2 ;
        RECT 40.204 3.604 42.676 3.636 ;
  LAYER M2 ;
        RECT 40.204 3.54 42.676 3.572 ;
  LAYER M2 ;
        RECT 40.204 3.476 42.676 3.508 ;
  LAYER M2 ;
        RECT 40.204 3.412 42.676 3.444 ;
  LAYER M2 ;
        RECT 40.204 3.348 42.676 3.38 ;
  LAYER M2 ;
        RECT 40.204 3.284 42.676 3.316 ;
  LAYER M2 ;
        RECT 40.204 3.22 42.676 3.252 ;
  LAYER M2 ;
        RECT 40.204 3.156 42.676 3.188 ;
  LAYER M2 ;
        RECT 40.204 3.092 42.676 3.124 ;
  LAYER M2 ;
        RECT 40.204 3.028 42.676 3.06 ;
  LAYER M2 ;
        RECT 40.204 2.964 42.676 2.996 ;
  LAYER M2 ;
        RECT 40.204 2.9 42.676 2.932 ;
  LAYER M2 ;
        RECT 40.204 2.836 42.676 2.868 ;
  LAYER M2 ;
        RECT 40.204 2.772 42.676 2.804 ;
  LAYER M2 ;
        RECT 40.204 2.708 42.676 2.74 ;
  LAYER M2 ;
        RECT 40.204 2.644 42.676 2.676 ;
  LAYER M2 ;
        RECT 40.204 2.58 42.676 2.612 ;
  LAYER M2 ;
        RECT 40.204 2.516 42.676 2.548 ;
  LAYER M2 ;
        RECT 40.204 2.452 42.676 2.484 ;
  LAYER M2 ;
        RECT 40.204 2.388 42.676 2.42 ;
  LAYER M2 ;
        RECT 40.204 2.324 42.676 2.356 ;
  LAYER M2 ;
        RECT 40.204 2.26 42.676 2.292 ;
  LAYER M2 ;
        RECT 40.204 2.196 42.676 2.228 ;
  LAYER M2 ;
        RECT 40.204 2.132 42.676 2.164 ;
  LAYER M3 ;
        RECT 40.224 1.98 40.256 4.488 ;
  LAYER M3 ;
        RECT 40.288 1.98 40.32 4.488 ;
  LAYER M3 ;
        RECT 40.352 1.98 40.384 4.488 ;
  LAYER M3 ;
        RECT 40.416 1.98 40.448 4.488 ;
  LAYER M3 ;
        RECT 40.48 1.98 40.512 4.488 ;
  LAYER M3 ;
        RECT 40.544 1.98 40.576 4.488 ;
  LAYER M3 ;
        RECT 40.608 1.98 40.64 4.488 ;
  LAYER M3 ;
        RECT 40.672 1.98 40.704 4.488 ;
  LAYER M3 ;
        RECT 40.736 1.98 40.768 4.488 ;
  LAYER M3 ;
        RECT 40.8 1.98 40.832 4.488 ;
  LAYER M3 ;
        RECT 40.864 1.98 40.896 4.488 ;
  LAYER M3 ;
        RECT 40.928 1.98 40.96 4.488 ;
  LAYER M3 ;
        RECT 40.992 1.98 41.024 4.488 ;
  LAYER M3 ;
        RECT 41.056 1.98 41.088 4.488 ;
  LAYER M3 ;
        RECT 41.12 1.98 41.152 4.488 ;
  LAYER M3 ;
        RECT 41.184 1.98 41.216 4.488 ;
  LAYER M3 ;
        RECT 41.248 1.98 41.28 4.488 ;
  LAYER M3 ;
        RECT 41.312 1.98 41.344 4.488 ;
  LAYER M3 ;
        RECT 41.376 1.98 41.408 4.488 ;
  LAYER M3 ;
        RECT 41.44 1.98 41.472 4.488 ;
  LAYER M3 ;
        RECT 41.504 1.98 41.536 4.488 ;
  LAYER M3 ;
        RECT 41.568 1.98 41.6 4.488 ;
  LAYER M3 ;
        RECT 41.632 1.98 41.664 4.488 ;
  LAYER M3 ;
        RECT 41.696 1.98 41.728 4.488 ;
  LAYER M3 ;
        RECT 41.76 1.98 41.792 4.488 ;
  LAYER M3 ;
        RECT 41.824 1.98 41.856 4.488 ;
  LAYER M3 ;
        RECT 41.888 1.98 41.92 4.488 ;
  LAYER M3 ;
        RECT 41.952 1.98 41.984 4.488 ;
  LAYER M3 ;
        RECT 42.016 1.98 42.048 4.488 ;
  LAYER M3 ;
        RECT 42.08 1.98 42.112 4.488 ;
  LAYER M3 ;
        RECT 42.144 1.98 42.176 4.488 ;
  LAYER M3 ;
        RECT 42.208 1.98 42.24 4.488 ;
  LAYER M3 ;
        RECT 42.272 1.98 42.304 4.488 ;
  LAYER M3 ;
        RECT 42.336 1.98 42.368 4.488 ;
  LAYER M3 ;
        RECT 42.4 1.98 42.432 4.488 ;
  LAYER M3 ;
        RECT 42.464 1.98 42.496 4.488 ;
  LAYER M3 ;
        RECT 42.528 1.98 42.56 4.488 ;
  LAYER M3 ;
        RECT 42.624 1.98 42.656 4.488 ;
  LAYER M1 ;
        RECT 40.239 2.016 40.241 4.452 ;
  LAYER M1 ;
        RECT 40.319 2.016 40.321 4.452 ;
  LAYER M1 ;
        RECT 40.399 2.016 40.401 4.452 ;
  LAYER M1 ;
        RECT 40.479 2.016 40.481 4.452 ;
  LAYER M1 ;
        RECT 40.559 2.016 40.561 4.452 ;
  LAYER M1 ;
        RECT 40.639 2.016 40.641 4.452 ;
  LAYER M1 ;
        RECT 40.719 2.016 40.721 4.452 ;
  LAYER M1 ;
        RECT 40.799 2.016 40.801 4.452 ;
  LAYER M1 ;
        RECT 40.879 2.016 40.881 4.452 ;
  LAYER M1 ;
        RECT 40.959 2.016 40.961 4.452 ;
  LAYER M1 ;
        RECT 41.039 2.016 41.041 4.452 ;
  LAYER M1 ;
        RECT 41.119 2.016 41.121 4.452 ;
  LAYER M1 ;
        RECT 41.199 2.016 41.201 4.452 ;
  LAYER M1 ;
        RECT 41.279 2.016 41.281 4.452 ;
  LAYER M1 ;
        RECT 41.359 2.016 41.361 4.452 ;
  LAYER M1 ;
        RECT 41.439 2.016 41.441 4.452 ;
  LAYER M1 ;
        RECT 41.519 2.016 41.521 4.452 ;
  LAYER M1 ;
        RECT 41.599 2.016 41.601 4.452 ;
  LAYER M1 ;
        RECT 41.679 2.016 41.681 4.452 ;
  LAYER M1 ;
        RECT 41.759 2.016 41.761 4.452 ;
  LAYER M1 ;
        RECT 41.839 2.016 41.841 4.452 ;
  LAYER M1 ;
        RECT 41.919 2.016 41.921 4.452 ;
  LAYER M1 ;
        RECT 41.999 2.016 42.001 4.452 ;
  LAYER M1 ;
        RECT 42.079 2.016 42.081 4.452 ;
  LAYER M1 ;
        RECT 42.159 2.016 42.161 4.452 ;
  LAYER M1 ;
        RECT 42.239 2.016 42.241 4.452 ;
  LAYER M1 ;
        RECT 42.319 2.016 42.321 4.452 ;
  LAYER M1 ;
        RECT 42.399 2.016 42.401 4.452 ;
  LAYER M1 ;
        RECT 42.479 2.016 42.481 4.452 ;
  LAYER M1 ;
        RECT 42.559 2.016 42.561 4.452 ;
  LAYER M2 ;
        RECT 40.24 4.451 42.64 4.453 ;
  LAYER M2 ;
        RECT 40.24 4.367 42.64 4.369 ;
  LAYER M2 ;
        RECT 40.24 4.283 42.64 4.285 ;
  LAYER M2 ;
        RECT 40.24 4.199 42.64 4.201 ;
  LAYER M2 ;
        RECT 40.24 4.115 42.64 4.117 ;
  LAYER M2 ;
        RECT 40.24 4.031 42.64 4.033 ;
  LAYER M2 ;
        RECT 40.24 3.947 42.64 3.949 ;
  LAYER M2 ;
        RECT 40.24 3.863 42.64 3.865 ;
  LAYER M2 ;
        RECT 40.24 3.779 42.64 3.781 ;
  LAYER M2 ;
        RECT 40.24 3.695 42.64 3.697 ;
  LAYER M2 ;
        RECT 40.24 3.611 42.64 3.613 ;
  LAYER M2 ;
        RECT 40.24 3.527 42.64 3.529 ;
  LAYER M2 ;
        RECT 40.24 3.4435 42.64 3.4455 ;
  LAYER M2 ;
        RECT 40.24 3.359 42.64 3.361 ;
  LAYER M2 ;
        RECT 40.24 3.275 42.64 3.277 ;
  LAYER M2 ;
        RECT 40.24 3.191 42.64 3.193 ;
  LAYER M2 ;
        RECT 40.24 3.107 42.64 3.109 ;
  LAYER M2 ;
        RECT 40.24 3.023 42.64 3.025 ;
  LAYER M2 ;
        RECT 40.24 2.939 42.64 2.941 ;
  LAYER M2 ;
        RECT 40.24 2.855 42.64 2.857 ;
  LAYER M2 ;
        RECT 40.24 2.771 42.64 2.773 ;
  LAYER M2 ;
        RECT 40.24 2.687 42.64 2.689 ;
  LAYER M2 ;
        RECT 40.24 2.603 42.64 2.605 ;
  LAYER M2 ;
        RECT 40.24 2.519 42.64 2.521 ;
  LAYER M2 ;
        RECT 40.24 2.435 42.64 2.437 ;
  LAYER M2 ;
        RECT 40.24 2.351 42.64 2.353 ;
  LAYER M2 ;
        RECT 40.24 2.267 42.64 2.269 ;
  LAYER M2 ;
        RECT 40.24 2.183 42.64 2.185 ;
  LAYER M2 ;
        RECT 40.24 2.099 42.64 2.101 ;
  LAYER M1 ;
        RECT 43.104 13.74 43.136 16.248 ;
  LAYER M1 ;
        RECT 43.168 13.74 43.2 16.248 ;
  LAYER M1 ;
        RECT 43.232 13.74 43.264 16.248 ;
  LAYER M1 ;
        RECT 43.296 13.74 43.328 16.248 ;
  LAYER M1 ;
        RECT 43.36 13.74 43.392 16.248 ;
  LAYER M1 ;
        RECT 43.424 13.74 43.456 16.248 ;
  LAYER M1 ;
        RECT 43.488 13.74 43.52 16.248 ;
  LAYER M1 ;
        RECT 43.552 13.74 43.584 16.248 ;
  LAYER M1 ;
        RECT 43.616 13.74 43.648 16.248 ;
  LAYER M1 ;
        RECT 43.68 13.74 43.712 16.248 ;
  LAYER M1 ;
        RECT 43.744 13.74 43.776 16.248 ;
  LAYER M1 ;
        RECT 43.808 13.74 43.84 16.248 ;
  LAYER M1 ;
        RECT 43.872 13.74 43.904 16.248 ;
  LAYER M1 ;
        RECT 43.936 13.74 43.968 16.248 ;
  LAYER M1 ;
        RECT 44 13.74 44.032 16.248 ;
  LAYER M1 ;
        RECT 44.064 13.74 44.096 16.248 ;
  LAYER M1 ;
        RECT 44.128 13.74 44.16 16.248 ;
  LAYER M1 ;
        RECT 44.192 13.74 44.224 16.248 ;
  LAYER M1 ;
        RECT 44.256 13.74 44.288 16.248 ;
  LAYER M1 ;
        RECT 44.32 13.74 44.352 16.248 ;
  LAYER M1 ;
        RECT 44.384 13.74 44.416 16.248 ;
  LAYER M1 ;
        RECT 44.448 13.74 44.48 16.248 ;
  LAYER M1 ;
        RECT 44.512 13.74 44.544 16.248 ;
  LAYER M1 ;
        RECT 44.576 13.74 44.608 16.248 ;
  LAYER M1 ;
        RECT 44.64 13.74 44.672 16.248 ;
  LAYER M1 ;
        RECT 44.704 13.74 44.736 16.248 ;
  LAYER M1 ;
        RECT 44.768 13.74 44.8 16.248 ;
  LAYER M1 ;
        RECT 44.832 13.74 44.864 16.248 ;
  LAYER M1 ;
        RECT 44.896 13.74 44.928 16.248 ;
  LAYER M1 ;
        RECT 44.96 13.74 44.992 16.248 ;
  LAYER M1 ;
        RECT 45.024 13.74 45.056 16.248 ;
  LAYER M1 ;
        RECT 45.088 13.74 45.12 16.248 ;
  LAYER M1 ;
        RECT 45.152 13.74 45.184 16.248 ;
  LAYER M1 ;
        RECT 45.216 13.74 45.248 16.248 ;
  LAYER M1 ;
        RECT 45.28 13.74 45.312 16.248 ;
  LAYER M1 ;
        RECT 45.344 13.74 45.376 16.248 ;
  LAYER M1 ;
        RECT 45.408 13.74 45.44 16.248 ;
  LAYER M2 ;
        RECT 43.084 16.132 45.556 16.164 ;
  LAYER M2 ;
        RECT 43.084 16.068 45.556 16.1 ;
  LAYER M2 ;
        RECT 43.084 16.004 45.556 16.036 ;
  LAYER M2 ;
        RECT 43.084 15.94 45.556 15.972 ;
  LAYER M2 ;
        RECT 43.084 15.876 45.556 15.908 ;
  LAYER M2 ;
        RECT 43.084 15.812 45.556 15.844 ;
  LAYER M2 ;
        RECT 43.084 15.748 45.556 15.78 ;
  LAYER M2 ;
        RECT 43.084 15.684 45.556 15.716 ;
  LAYER M2 ;
        RECT 43.084 15.62 45.556 15.652 ;
  LAYER M2 ;
        RECT 43.084 15.556 45.556 15.588 ;
  LAYER M2 ;
        RECT 43.084 15.492 45.556 15.524 ;
  LAYER M2 ;
        RECT 43.084 15.428 45.556 15.46 ;
  LAYER M2 ;
        RECT 43.084 15.364 45.556 15.396 ;
  LAYER M2 ;
        RECT 43.084 15.3 45.556 15.332 ;
  LAYER M2 ;
        RECT 43.084 15.236 45.556 15.268 ;
  LAYER M2 ;
        RECT 43.084 15.172 45.556 15.204 ;
  LAYER M2 ;
        RECT 43.084 15.108 45.556 15.14 ;
  LAYER M2 ;
        RECT 43.084 15.044 45.556 15.076 ;
  LAYER M2 ;
        RECT 43.084 14.98 45.556 15.012 ;
  LAYER M2 ;
        RECT 43.084 14.916 45.556 14.948 ;
  LAYER M2 ;
        RECT 43.084 14.852 45.556 14.884 ;
  LAYER M2 ;
        RECT 43.084 14.788 45.556 14.82 ;
  LAYER M2 ;
        RECT 43.084 14.724 45.556 14.756 ;
  LAYER M2 ;
        RECT 43.084 14.66 45.556 14.692 ;
  LAYER M2 ;
        RECT 43.084 14.596 45.556 14.628 ;
  LAYER M2 ;
        RECT 43.084 14.532 45.556 14.564 ;
  LAYER M2 ;
        RECT 43.084 14.468 45.556 14.5 ;
  LAYER M2 ;
        RECT 43.084 14.404 45.556 14.436 ;
  LAYER M2 ;
        RECT 43.084 14.34 45.556 14.372 ;
  LAYER M2 ;
        RECT 43.084 14.276 45.556 14.308 ;
  LAYER M2 ;
        RECT 43.084 14.212 45.556 14.244 ;
  LAYER M2 ;
        RECT 43.084 14.148 45.556 14.18 ;
  LAYER M2 ;
        RECT 43.084 14.084 45.556 14.116 ;
  LAYER M2 ;
        RECT 43.084 14.02 45.556 14.052 ;
  LAYER M2 ;
        RECT 43.084 13.956 45.556 13.988 ;
  LAYER M2 ;
        RECT 43.084 13.892 45.556 13.924 ;
  LAYER M3 ;
        RECT 43.104 13.74 43.136 16.248 ;
  LAYER M3 ;
        RECT 43.168 13.74 43.2 16.248 ;
  LAYER M3 ;
        RECT 43.232 13.74 43.264 16.248 ;
  LAYER M3 ;
        RECT 43.296 13.74 43.328 16.248 ;
  LAYER M3 ;
        RECT 43.36 13.74 43.392 16.248 ;
  LAYER M3 ;
        RECT 43.424 13.74 43.456 16.248 ;
  LAYER M3 ;
        RECT 43.488 13.74 43.52 16.248 ;
  LAYER M3 ;
        RECT 43.552 13.74 43.584 16.248 ;
  LAYER M3 ;
        RECT 43.616 13.74 43.648 16.248 ;
  LAYER M3 ;
        RECT 43.68 13.74 43.712 16.248 ;
  LAYER M3 ;
        RECT 43.744 13.74 43.776 16.248 ;
  LAYER M3 ;
        RECT 43.808 13.74 43.84 16.248 ;
  LAYER M3 ;
        RECT 43.872 13.74 43.904 16.248 ;
  LAYER M3 ;
        RECT 43.936 13.74 43.968 16.248 ;
  LAYER M3 ;
        RECT 44 13.74 44.032 16.248 ;
  LAYER M3 ;
        RECT 44.064 13.74 44.096 16.248 ;
  LAYER M3 ;
        RECT 44.128 13.74 44.16 16.248 ;
  LAYER M3 ;
        RECT 44.192 13.74 44.224 16.248 ;
  LAYER M3 ;
        RECT 44.256 13.74 44.288 16.248 ;
  LAYER M3 ;
        RECT 44.32 13.74 44.352 16.248 ;
  LAYER M3 ;
        RECT 44.384 13.74 44.416 16.248 ;
  LAYER M3 ;
        RECT 44.448 13.74 44.48 16.248 ;
  LAYER M3 ;
        RECT 44.512 13.74 44.544 16.248 ;
  LAYER M3 ;
        RECT 44.576 13.74 44.608 16.248 ;
  LAYER M3 ;
        RECT 44.64 13.74 44.672 16.248 ;
  LAYER M3 ;
        RECT 44.704 13.74 44.736 16.248 ;
  LAYER M3 ;
        RECT 44.768 13.74 44.8 16.248 ;
  LAYER M3 ;
        RECT 44.832 13.74 44.864 16.248 ;
  LAYER M3 ;
        RECT 44.896 13.74 44.928 16.248 ;
  LAYER M3 ;
        RECT 44.96 13.74 44.992 16.248 ;
  LAYER M3 ;
        RECT 45.024 13.74 45.056 16.248 ;
  LAYER M3 ;
        RECT 45.088 13.74 45.12 16.248 ;
  LAYER M3 ;
        RECT 45.152 13.74 45.184 16.248 ;
  LAYER M3 ;
        RECT 45.216 13.74 45.248 16.248 ;
  LAYER M3 ;
        RECT 45.28 13.74 45.312 16.248 ;
  LAYER M3 ;
        RECT 45.344 13.74 45.376 16.248 ;
  LAYER M3 ;
        RECT 45.408 13.74 45.44 16.248 ;
  LAYER M3 ;
        RECT 45.504 13.74 45.536 16.248 ;
  LAYER M1 ;
        RECT 43.119 13.776 43.121 16.212 ;
  LAYER M1 ;
        RECT 43.199 13.776 43.201 16.212 ;
  LAYER M1 ;
        RECT 43.279 13.776 43.281 16.212 ;
  LAYER M1 ;
        RECT 43.359 13.776 43.361 16.212 ;
  LAYER M1 ;
        RECT 43.439 13.776 43.441 16.212 ;
  LAYER M1 ;
        RECT 43.519 13.776 43.521 16.212 ;
  LAYER M1 ;
        RECT 43.599 13.776 43.601 16.212 ;
  LAYER M1 ;
        RECT 43.679 13.776 43.681 16.212 ;
  LAYER M1 ;
        RECT 43.759 13.776 43.761 16.212 ;
  LAYER M1 ;
        RECT 43.839 13.776 43.841 16.212 ;
  LAYER M1 ;
        RECT 43.919 13.776 43.921 16.212 ;
  LAYER M1 ;
        RECT 43.999 13.776 44.001 16.212 ;
  LAYER M1 ;
        RECT 44.079 13.776 44.081 16.212 ;
  LAYER M1 ;
        RECT 44.159 13.776 44.161 16.212 ;
  LAYER M1 ;
        RECT 44.239 13.776 44.241 16.212 ;
  LAYER M1 ;
        RECT 44.319 13.776 44.321 16.212 ;
  LAYER M1 ;
        RECT 44.399 13.776 44.401 16.212 ;
  LAYER M1 ;
        RECT 44.479 13.776 44.481 16.212 ;
  LAYER M1 ;
        RECT 44.559 13.776 44.561 16.212 ;
  LAYER M1 ;
        RECT 44.639 13.776 44.641 16.212 ;
  LAYER M1 ;
        RECT 44.719 13.776 44.721 16.212 ;
  LAYER M1 ;
        RECT 44.799 13.776 44.801 16.212 ;
  LAYER M1 ;
        RECT 44.879 13.776 44.881 16.212 ;
  LAYER M1 ;
        RECT 44.959 13.776 44.961 16.212 ;
  LAYER M1 ;
        RECT 45.039 13.776 45.041 16.212 ;
  LAYER M1 ;
        RECT 45.119 13.776 45.121 16.212 ;
  LAYER M1 ;
        RECT 45.199 13.776 45.201 16.212 ;
  LAYER M1 ;
        RECT 45.279 13.776 45.281 16.212 ;
  LAYER M1 ;
        RECT 45.359 13.776 45.361 16.212 ;
  LAYER M1 ;
        RECT 45.439 13.776 45.441 16.212 ;
  LAYER M2 ;
        RECT 43.12 16.211 45.52 16.213 ;
  LAYER M2 ;
        RECT 43.12 16.127 45.52 16.129 ;
  LAYER M2 ;
        RECT 43.12 16.043 45.52 16.045 ;
  LAYER M2 ;
        RECT 43.12 15.959 45.52 15.961 ;
  LAYER M2 ;
        RECT 43.12 15.875 45.52 15.877 ;
  LAYER M2 ;
        RECT 43.12 15.791 45.52 15.793 ;
  LAYER M2 ;
        RECT 43.12 15.707 45.52 15.709 ;
  LAYER M2 ;
        RECT 43.12 15.623 45.52 15.625 ;
  LAYER M2 ;
        RECT 43.12 15.539 45.52 15.541 ;
  LAYER M2 ;
        RECT 43.12 15.455 45.52 15.457 ;
  LAYER M2 ;
        RECT 43.12 15.371 45.52 15.373 ;
  LAYER M2 ;
        RECT 43.12 15.287 45.52 15.289 ;
  LAYER M2 ;
        RECT 43.12 15.2035 45.52 15.2055 ;
  LAYER M2 ;
        RECT 43.12 15.119 45.52 15.121 ;
  LAYER M2 ;
        RECT 43.12 15.035 45.52 15.037 ;
  LAYER M2 ;
        RECT 43.12 14.951 45.52 14.953 ;
  LAYER M2 ;
        RECT 43.12 14.867 45.52 14.869 ;
  LAYER M2 ;
        RECT 43.12 14.783 45.52 14.785 ;
  LAYER M2 ;
        RECT 43.12 14.699 45.52 14.701 ;
  LAYER M2 ;
        RECT 43.12 14.615 45.52 14.617 ;
  LAYER M2 ;
        RECT 43.12 14.531 45.52 14.533 ;
  LAYER M2 ;
        RECT 43.12 14.447 45.52 14.449 ;
  LAYER M2 ;
        RECT 43.12 14.363 45.52 14.365 ;
  LAYER M2 ;
        RECT 43.12 14.279 45.52 14.281 ;
  LAYER M2 ;
        RECT 43.12 14.195 45.52 14.197 ;
  LAYER M2 ;
        RECT 43.12 14.111 45.52 14.113 ;
  LAYER M2 ;
        RECT 43.12 14.027 45.52 14.029 ;
  LAYER M2 ;
        RECT 43.12 13.943 45.52 13.945 ;
  LAYER M2 ;
        RECT 43.12 13.859 45.52 13.861 ;
  LAYER M1 ;
        RECT 43.104 10.8 43.136 13.308 ;
  LAYER M1 ;
        RECT 43.168 10.8 43.2 13.308 ;
  LAYER M1 ;
        RECT 43.232 10.8 43.264 13.308 ;
  LAYER M1 ;
        RECT 43.296 10.8 43.328 13.308 ;
  LAYER M1 ;
        RECT 43.36 10.8 43.392 13.308 ;
  LAYER M1 ;
        RECT 43.424 10.8 43.456 13.308 ;
  LAYER M1 ;
        RECT 43.488 10.8 43.52 13.308 ;
  LAYER M1 ;
        RECT 43.552 10.8 43.584 13.308 ;
  LAYER M1 ;
        RECT 43.616 10.8 43.648 13.308 ;
  LAYER M1 ;
        RECT 43.68 10.8 43.712 13.308 ;
  LAYER M1 ;
        RECT 43.744 10.8 43.776 13.308 ;
  LAYER M1 ;
        RECT 43.808 10.8 43.84 13.308 ;
  LAYER M1 ;
        RECT 43.872 10.8 43.904 13.308 ;
  LAYER M1 ;
        RECT 43.936 10.8 43.968 13.308 ;
  LAYER M1 ;
        RECT 44 10.8 44.032 13.308 ;
  LAYER M1 ;
        RECT 44.064 10.8 44.096 13.308 ;
  LAYER M1 ;
        RECT 44.128 10.8 44.16 13.308 ;
  LAYER M1 ;
        RECT 44.192 10.8 44.224 13.308 ;
  LAYER M1 ;
        RECT 44.256 10.8 44.288 13.308 ;
  LAYER M1 ;
        RECT 44.32 10.8 44.352 13.308 ;
  LAYER M1 ;
        RECT 44.384 10.8 44.416 13.308 ;
  LAYER M1 ;
        RECT 44.448 10.8 44.48 13.308 ;
  LAYER M1 ;
        RECT 44.512 10.8 44.544 13.308 ;
  LAYER M1 ;
        RECT 44.576 10.8 44.608 13.308 ;
  LAYER M1 ;
        RECT 44.64 10.8 44.672 13.308 ;
  LAYER M1 ;
        RECT 44.704 10.8 44.736 13.308 ;
  LAYER M1 ;
        RECT 44.768 10.8 44.8 13.308 ;
  LAYER M1 ;
        RECT 44.832 10.8 44.864 13.308 ;
  LAYER M1 ;
        RECT 44.896 10.8 44.928 13.308 ;
  LAYER M1 ;
        RECT 44.96 10.8 44.992 13.308 ;
  LAYER M1 ;
        RECT 45.024 10.8 45.056 13.308 ;
  LAYER M1 ;
        RECT 45.088 10.8 45.12 13.308 ;
  LAYER M1 ;
        RECT 45.152 10.8 45.184 13.308 ;
  LAYER M1 ;
        RECT 45.216 10.8 45.248 13.308 ;
  LAYER M1 ;
        RECT 45.28 10.8 45.312 13.308 ;
  LAYER M1 ;
        RECT 45.344 10.8 45.376 13.308 ;
  LAYER M1 ;
        RECT 45.408 10.8 45.44 13.308 ;
  LAYER M2 ;
        RECT 43.084 13.192 45.556 13.224 ;
  LAYER M2 ;
        RECT 43.084 13.128 45.556 13.16 ;
  LAYER M2 ;
        RECT 43.084 13.064 45.556 13.096 ;
  LAYER M2 ;
        RECT 43.084 13 45.556 13.032 ;
  LAYER M2 ;
        RECT 43.084 12.936 45.556 12.968 ;
  LAYER M2 ;
        RECT 43.084 12.872 45.556 12.904 ;
  LAYER M2 ;
        RECT 43.084 12.808 45.556 12.84 ;
  LAYER M2 ;
        RECT 43.084 12.744 45.556 12.776 ;
  LAYER M2 ;
        RECT 43.084 12.68 45.556 12.712 ;
  LAYER M2 ;
        RECT 43.084 12.616 45.556 12.648 ;
  LAYER M2 ;
        RECT 43.084 12.552 45.556 12.584 ;
  LAYER M2 ;
        RECT 43.084 12.488 45.556 12.52 ;
  LAYER M2 ;
        RECT 43.084 12.424 45.556 12.456 ;
  LAYER M2 ;
        RECT 43.084 12.36 45.556 12.392 ;
  LAYER M2 ;
        RECT 43.084 12.296 45.556 12.328 ;
  LAYER M2 ;
        RECT 43.084 12.232 45.556 12.264 ;
  LAYER M2 ;
        RECT 43.084 12.168 45.556 12.2 ;
  LAYER M2 ;
        RECT 43.084 12.104 45.556 12.136 ;
  LAYER M2 ;
        RECT 43.084 12.04 45.556 12.072 ;
  LAYER M2 ;
        RECT 43.084 11.976 45.556 12.008 ;
  LAYER M2 ;
        RECT 43.084 11.912 45.556 11.944 ;
  LAYER M2 ;
        RECT 43.084 11.848 45.556 11.88 ;
  LAYER M2 ;
        RECT 43.084 11.784 45.556 11.816 ;
  LAYER M2 ;
        RECT 43.084 11.72 45.556 11.752 ;
  LAYER M2 ;
        RECT 43.084 11.656 45.556 11.688 ;
  LAYER M2 ;
        RECT 43.084 11.592 45.556 11.624 ;
  LAYER M2 ;
        RECT 43.084 11.528 45.556 11.56 ;
  LAYER M2 ;
        RECT 43.084 11.464 45.556 11.496 ;
  LAYER M2 ;
        RECT 43.084 11.4 45.556 11.432 ;
  LAYER M2 ;
        RECT 43.084 11.336 45.556 11.368 ;
  LAYER M2 ;
        RECT 43.084 11.272 45.556 11.304 ;
  LAYER M2 ;
        RECT 43.084 11.208 45.556 11.24 ;
  LAYER M2 ;
        RECT 43.084 11.144 45.556 11.176 ;
  LAYER M2 ;
        RECT 43.084 11.08 45.556 11.112 ;
  LAYER M2 ;
        RECT 43.084 11.016 45.556 11.048 ;
  LAYER M2 ;
        RECT 43.084 10.952 45.556 10.984 ;
  LAYER M3 ;
        RECT 43.104 10.8 43.136 13.308 ;
  LAYER M3 ;
        RECT 43.168 10.8 43.2 13.308 ;
  LAYER M3 ;
        RECT 43.232 10.8 43.264 13.308 ;
  LAYER M3 ;
        RECT 43.296 10.8 43.328 13.308 ;
  LAYER M3 ;
        RECT 43.36 10.8 43.392 13.308 ;
  LAYER M3 ;
        RECT 43.424 10.8 43.456 13.308 ;
  LAYER M3 ;
        RECT 43.488 10.8 43.52 13.308 ;
  LAYER M3 ;
        RECT 43.552 10.8 43.584 13.308 ;
  LAYER M3 ;
        RECT 43.616 10.8 43.648 13.308 ;
  LAYER M3 ;
        RECT 43.68 10.8 43.712 13.308 ;
  LAYER M3 ;
        RECT 43.744 10.8 43.776 13.308 ;
  LAYER M3 ;
        RECT 43.808 10.8 43.84 13.308 ;
  LAYER M3 ;
        RECT 43.872 10.8 43.904 13.308 ;
  LAYER M3 ;
        RECT 43.936 10.8 43.968 13.308 ;
  LAYER M3 ;
        RECT 44 10.8 44.032 13.308 ;
  LAYER M3 ;
        RECT 44.064 10.8 44.096 13.308 ;
  LAYER M3 ;
        RECT 44.128 10.8 44.16 13.308 ;
  LAYER M3 ;
        RECT 44.192 10.8 44.224 13.308 ;
  LAYER M3 ;
        RECT 44.256 10.8 44.288 13.308 ;
  LAYER M3 ;
        RECT 44.32 10.8 44.352 13.308 ;
  LAYER M3 ;
        RECT 44.384 10.8 44.416 13.308 ;
  LAYER M3 ;
        RECT 44.448 10.8 44.48 13.308 ;
  LAYER M3 ;
        RECT 44.512 10.8 44.544 13.308 ;
  LAYER M3 ;
        RECT 44.576 10.8 44.608 13.308 ;
  LAYER M3 ;
        RECT 44.64 10.8 44.672 13.308 ;
  LAYER M3 ;
        RECT 44.704 10.8 44.736 13.308 ;
  LAYER M3 ;
        RECT 44.768 10.8 44.8 13.308 ;
  LAYER M3 ;
        RECT 44.832 10.8 44.864 13.308 ;
  LAYER M3 ;
        RECT 44.896 10.8 44.928 13.308 ;
  LAYER M3 ;
        RECT 44.96 10.8 44.992 13.308 ;
  LAYER M3 ;
        RECT 45.024 10.8 45.056 13.308 ;
  LAYER M3 ;
        RECT 45.088 10.8 45.12 13.308 ;
  LAYER M3 ;
        RECT 45.152 10.8 45.184 13.308 ;
  LAYER M3 ;
        RECT 45.216 10.8 45.248 13.308 ;
  LAYER M3 ;
        RECT 45.28 10.8 45.312 13.308 ;
  LAYER M3 ;
        RECT 45.344 10.8 45.376 13.308 ;
  LAYER M3 ;
        RECT 45.408 10.8 45.44 13.308 ;
  LAYER M3 ;
        RECT 45.504 10.8 45.536 13.308 ;
  LAYER M1 ;
        RECT 43.119 10.836 43.121 13.272 ;
  LAYER M1 ;
        RECT 43.199 10.836 43.201 13.272 ;
  LAYER M1 ;
        RECT 43.279 10.836 43.281 13.272 ;
  LAYER M1 ;
        RECT 43.359 10.836 43.361 13.272 ;
  LAYER M1 ;
        RECT 43.439 10.836 43.441 13.272 ;
  LAYER M1 ;
        RECT 43.519 10.836 43.521 13.272 ;
  LAYER M1 ;
        RECT 43.599 10.836 43.601 13.272 ;
  LAYER M1 ;
        RECT 43.679 10.836 43.681 13.272 ;
  LAYER M1 ;
        RECT 43.759 10.836 43.761 13.272 ;
  LAYER M1 ;
        RECT 43.839 10.836 43.841 13.272 ;
  LAYER M1 ;
        RECT 43.919 10.836 43.921 13.272 ;
  LAYER M1 ;
        RECT 43.999 10.836 44.001 13.272 ;
  LAYER M1 ;
        RECT 44.079 10.836 44.081 13.272 ;
  LAYER M1 ;
        RECT 44.159 10.836 44.161 13.272 ;
  LAYER M1 ;
        RECT 44.239 10.836 44.241 13.272 ;
  LAYER M1 ;
        RECT 44.319 10.836 44.321 13.272 ;
  LAYER M1 ;
        RECT 44.399 10.836 44.401 13.272 ;
  LAYER M1 ;
        RECT 44.479 10.836 44.481 13.272 ;
  LAYER M1 ;
        RECT 44.559 10.836 44.561 13.272 ;
  LAYER M1 ;
        RECT 44.639 10.836 44.641 13.272 ;
  LAYER M1 ;
        RECT 44.719 10.836 44.721 13.272 ;
  LAYER M1 ;
        RECT 44.799 10.836 44.801 13.272 ;
  LAYER M1 ;
        RECT 44.879 10.836 44.881 13.272 ;
  LAYER M1 ;
        RECT 44.959 10.836 44.961 13.272 ;
  LAYER M1 ;
        RECT 45.039 10.836 45.041 13.272 ;
  LAYER M1 ;
        RECT 45.119 10.836 45.121 13.272 ;
  LAYER M1 ;
        RECT 45.199 10.836 45.201 13.272 ;
  LAYER M1 ;
        RECT 45.279 10.836 45.281 13.272 ;
  LAYER M1 ;
        RECT 45.359 10.836 45.361 13.272 ;
  LAYER M1 ;
        RECT 45.439 10.836 45.441 13.272 ;
  LAYER M2 ;
        RECT 43.12 13.271 45.52 13.273 ;
  LAYER M2 ;
        RECT 43.12 13.187 45.52 13.189 ;
  LAYER M2 ;
        RECT 43.12 13.103 45.52 13.105 ;
  LAYER M2 ;
        RECT 43.12 13.019 45.52 13.021 ;
  LAYER M2 ;
        RECT 43.12 12.935 45.52 12.937 ;
  LAYER M2 ;
        RECT 43.12 12.851 45.52 12.853 ;
  LAYER M2 ;
        RECT 43.12 12.767 45.52 12.769 ;
  LAYER M2 ;
        RECT 43.12 12.683 45.52 12.685 ;
  LAYER M2 ;
        RECT 43.12 12.599 45.52 12.601 ;
  LAYER M2 ;
        RECT 43.12 12.515 45.52 12.517 ;
  LAYER M2 ;
        RECT 43.12 12.431 45.52 12.433 ;
  LAYER M2 ;
        RECT 43.12 12.347 45.52 12.349 ;
  LAYER M2 ;
        RECT 43.12 12.2635 45.52 12.2655 ;
  LAYER M2 ;
        RECT 43.12 12.179 45.52 12.181 ;
  LAYER M2 ;
        RECT 43.12 12.095 45.52 12.097 ;
  LAYER M2 ;
        RECT 43.12 12.011 45.52 12.013 ;
  LAYER M2 ;
        RECT 43.12 11.927 45.52 11.929 ;
  LAYER M2 ;
        RECT 43.12 11.843 45.52 11.845 ;
  LAYER M2 ;
        RECT 43.12 11.759 45.52 11.761 ;
  LAYER M2 ;
        RECT 43.12 11.675 45.52 11.677 ;
  LAYER M2 ;
        RECT 43.12 11.591 45.52 11.593 ;
  LAYER M2 ;
        RECT 43.12 11.507 45.52 11.509 ;
  LAYER M2 ;
        RECT 43.12 11.423 45.52 11.425 ;
  LAYER M2 ;
        RECT 43.12 11.339 45.52 11.341 ;
  LAYER M2 ;
        RECT 43.12 11.255 45.52 11.257 ;
  LAYER M2 ;
        RECT 43.12 11.171 45.52 11.173 ;
  LAYER M2 ;
        RECT 43.12 11.087 45.52 11.089 ;
  LAYER M2 ;
        RECT 43.12 11.003 45.52 11.005 ;
  LAYER M2 ;
        RECT 43.12 10.919 45.52 10.921 ;
  LAYER M1 ;
        RECT 43.104 7.86 43.136 10.368 ;
  LAYER M1 ;
        RECT 43.168 7.86 43.2 10.368 ;
  LAYER M1 ;
        RECT 43.232 7.86 43.264 10.368 ;
  LAYER M1 ;
        RECT 43.296 7.86 43.328 10.368 ;
  LAYER M1 ;
        RECT 43.36 7.86 43.392 10.368 ;
  LAYER M1 ;
        RECT 43.424 7.86 43.456 10.368 ;
  LAYER M1 ;
        RECT 43.488 7.86 43.52 10.368 ;
  LAYER M1 ;
        RECT 43.552 7.86 43.584 10.368 ;
  LAYER M1 ;
        RECT 43.616 7.86 43.648 10.368 ;
  LAYER M1 ;
        RECT 43.68 7.86 43.712 10.368 ;
  LAYER M1 ;
        RECT 43.744 7.86 43.776 10.368 ;
  LAYER M1 ;
        RECT 43.808 7.86 43.84 10.368 ;
  LAYER M1 ;
        RECT 43.872 7.86 43.904 10.368 ;
  LAYER M1 ;
        RECT 43.936 7.86 43.968 10.368 ;
  LAYER M1 ;
        RECT 44 7.86 44.032 10.368 ;
  LAYER M1 ;
        RECT 44.064 7.86 44.096 10.368 ;
  LAYER M1 ;
        RECT 44.128 7.86 44.16 10.368 ;
  LAYER M1 ;
        RECT 44.192 7.86 44.224 10.368 ;
  LAYER M1 ;
        RECT 44.256 7.86 44.288 10.368 ;
  LAYER M1 ;
        RECT 44.32 7.86 44.352 10.368 ;
  LAYER M1 ;
        RECT 44.384 7.86 44.416 10.368 ;
  LAYER M1 ;
        RECT 44.448 7.86 44.48 10.368 ;
  LAYER M1 ;
        RECT 44.512 7.86 44.544 10.368 ;
  LAYER M1 ;
        RECT 44.576 7.86 44.608 10.368 ;
  LAYER M1 ;
        RECT 44.64 7.86 44.672 10.368 ;
  LAYER M1 ;
        RECT 44.704 7.86 44.736 10.368 ;
  LAYER M1 ;
        RECT 44.768 7.86 44.8 10.368 ;
  LAYER M1 ;
        RECT 44.832 7.86 44.864 10.368 ;
  LAYER M1 ;
        RECT 44.896 7.86 44.928 10.368 ;
  LAYER M1 ;
        RECT 44.96 7.86 44.992 10.368 ;
  LAYER M1 ;
        RECT 45.024 7.86 45.056 10.368 ;
  LAYER M1 ;
        RECT 45.088 7.86 45.12 10.368 ;
  LAYER M1 ;
        RECT 45.152 7.86 45.184 10.368 ;
  LAYER M1 ;
        RECT 45.216 7.86 45.248 10.368 ;
  LAYER M1 ;
        RECT 45.28 7.86 45.312 10.368 ;
  LAYER M1 ;
        RECT 45.344 7.86 45.376 10.368 ;
  LAYER M1 ;
        RECT 45.408 7.86 45.44 10.368 ;
  LAYER M2 ;
        RECT 43.084 10.252 45.556 10.284 ;
  LAYER M2 ;
        RECT 43.084 10.188 45.556 10.22 ;
  LAYER M2 ;
        RECT 43.084 10.124 45.556 10.156 ;
  LAYER M2 ;
        RECT 43.084 10.06 45.556 10.092 ;
  LAYER M2 ;
        RECT 43.084 9.996 45.556 10.028 ;
  LAYER M2 ;
        RECT 43.084 9.932 45.556 9.964 ;
  LAYER M2 ;
        RECT 43.084 9.868 45.556 9.9 ;
  LAYER M2 ;
        RECT 43.084 9.804 45.556 9.836 ;
  LAYER M2 ;
        RECT 43.084 9.74 45.556 9.772 ;
  LAYER M2 ;
        RECT 43.084 9.676 45.556 9.708 ;
  LAYER M2 ;
        RECT 43.084 9.612 45.556 9.644 ;
  LAYER M2 ;
        RECT 43.084 9.548 45.556 9.58 ;
  LAYER M2 ;
        RECT 43.084 9.484 45.556 9.516 ;
  LAYER M2 ;
        RECT 43.084 9.42 45.556 9.452 ;
  LAYER M2 ;
        RECT 43.084 9.356 45.556 9.388 ;
  LAYER M2 ;
        RECT 43.084 9.292 45.556 9.324 ;
  LAYER M2 ;
        RECT 43.084 9.228 45.556 9.26 ;
  LAYER M2 ;
        RECT 43.084 9.164 45.556 9.196 ;
  LAYER M2 ;
        RECT 43.084 9.1 45.556 9.132 ;
  LAYER M2 ;
        RECT 43.084 9.036 45.556 9.068 ;
  LAYER M2 ;
        RECT 43.084 8.972 45.556 9.004 ;
  LAYER M2 ;
        RECT 43.084 8.908 45.556 8.94 ;
  LAYER M2 ;
        RECT 43.084 8.844 45.556 8.876 ;
  LAYER M2 ;
        RECT 43.084 8.78 45.556 8.812 ;
  LAYER M2 ;
        RECT 43.084 8.716 45.556 8.748 ;
  LAYER M2 ;
        RECT 43.084 8.652 45.556 8.684 ;
  LAYER M2 ;
        RECT 43.084 8.588 45.556 8.62 ;
  LAYER M2 ;
        RECT 43.084 8.524 45.556 8.556 ;
  LAYER M2 ;
        RECT 43.084 8.46 45.556 8.492 ;
  LAYER M2 ;
        RECT 43.084 8.396 45.556 8.428 ;
  LAYER M2 ;
        RECT 43.084 8.332 45.556 8.364 ;
  LAYER M2 ;
        RECT 43.084 8.268 45.556 8.3 ;
  LAYER M2 ;
        RECT 43.084 8.204 45.556 8.236 ;
  LAYER M2 ;
        RECT 43.084 8.14 45.556 8.172 ;
  LAYER M2 ;
        RECT 43.084 8.076 45.556 8.108 ;
  LAYER M2 ;
        RECT 43.084 8.012 45.556 8.044 ;
  LAYER M3 ;
        RECT 43.104 7.86 43.136 10.368 ;
  LAYER M3 ;
        RECT 43.168 7.86 43.2 10.368 ;
  LAYER M3 ;
        RECT 43.232 7.86 43.264 10.368 ;
  LAYER M3 ;
        RECT 43.296 7.86 43.328 10.368 ;
  LAYER M3 ;
        RECT 43.36 7.86 43.392 10.368 ;
  LAYER M3 ;
        RECT 43.424 7.86 43.456 10.368 ;
  LAYER M3 ;
        RECT 43.488 7.86 43.52 10.368 ;
  LAYER M3 ;
        RECT 43.552 7.86 43.584 10.368 ;
  LAYER M3 ;
        RECT 43.616 7.86 43.648 10.368 ;
  LAYER M3 ;
        RECT 43.68 7.86 43.712 10.368 ;
  LAYER M3 ;
        RECT 43.744 7.86 43.776 10.368 ;
  LAYER M3 ;
        RECT 43.808 7.86 43.84 10.368 ;
  LAYER M3 ;
        RECT 43.872 7.86 43.904 10.368 ;
  LAYER M3 ;
        RECT 43.936 7.86 43.968 10.368 ;
  LAYER M3 ;
        RECT 44 7.86 44.032 10.368 ;
  LAYER M3 ;
        RECT 44.064 7.86 44.096 10.368 ;
  LAYER M3 ;
        RECT 44.128 7.86 44.16 10.368 ;
  LAYER M3 ;
        RECT 44.192 7.86 44.224 10.368 ;
  LAYER M3 ;
        RECT 44.256 7.86 44.288 10.368 ;
  LAYER M3 ;
        RECT 44.32 7.86 44.352 10.368 ;
  LAYER M3 ;
        RECT 44.384 7.86 44.416 10.368 ;
  LAYER M3 ;
        RECT 44.448 7.86 44.48 10.368 ;
  LAYER M3 ;
        RECT 44.512 7.86 44.544 10.368 ;
  LAYER M3 ;
        RECT 44.576 7.86 44.608 10.368 ;
  LAYER M3 ;
        RECT 44.64 7.86 44.672 10.368 ;
  LAYER M3 ;
        RECT 44.704 7.86 44.736 10.368 ;
  LAYER M3 ;
        RECT 44.768 7.86 44.8 10.368 ;
  LAYER M3 ;
        RECT 44.832 7.86 44.864 10.368 ;
  LAYER M3 ;
        RECT 44.896 7.86 44.928 10.368 ;
  LAYER M3 ;
        RECT 44.96 7.86 44.992 10.368 ;
  LAYER M3 ;
        RECT 45.024 7.86 45.056 10.368 ;
  LAYER M3 ;
        RECT 45.088 7.86 45.12 10.368 ;
  LAYER M3 ;
        RECT 45.152 7.86 45.184 10.368 ;
  LAYER M3 ;
        RECT 45.216 7.86 45.248 10.368 ;
  LAYER M3 ;
        RECT 45.28 7.86 45.312 10.368 ;
  LAYER M3 ;
        RECT 45.344 7.86 45.376 10.368 ;
  LAYER M3 ;
        RECT 45.408 7.86 45.44 10.368 ;
  LAYER M3 ;
        RECT 45.504 7.86 45.536 10.368 ;
  LAYER M1 ;
        RECT 43.119 7.896 43.121 10.332 ;
  LAYER M1 ;
        RECT 43.199 7.896 43.201 10.332 ;
  LAYER M1 ;
        RECT 43.279 7.896 43.281 10.332 ;
  LAYER M1 ;
        RECT 43.359 7.896 43.361 10.332 ;
  LAYER M1 ;
        RECT 43.439 7.896 43.441 10.332 ;
  LAYER M1 ;
        RECT 43.519 7.896 43.521 10.332 ;
  LAYER M1 ;
        RECT 43.599 7.896 43.601 10.332 ;
  LAYER M1 ;
        RECT 43.679 7.896 43.681 10.332 ;
  LAYER M1 ;
        RECT 43.759 7.896 43.761 10.332 ;
  LAYER M1 ;
        RECT 43.839 7.896 43.841 10.332 ;
  LAYER M1 ;
        RECT 43.919 7.896 43.921 10.332 ;
  LAYER M1 ;
        RECT 43.999 7.896 44.001 10.332 ;
  LAYER M1 ;
        RECT 44.079 7.896 44.081 10.332 ;
  LAYER M1 ;
        RECT 44.159 7.896 44.161 10.332 ;
  LAYER M1 ;
        RECT 44.239 7.896 44.241 10.332 ;
  LAYER M1 ;
        RECT 44.319 7.896 44.321 10.332 ;
  LAYER M1 ;
        RECT 44.399 7.896 44.401 10.332 ;
  LAYER M1 ;
        RECT 44.479 7.896 44.481 10.332 ;
  LAYER M1 ;
        RECT 44.559 7.896 44.561 10.332 ;
  LAYER M1 ;
        RECT 44.639 7.896 44.641 10.332 ;
  LAYER M1 ;
        RECT 44.719 7.896 44.721 10.332 ;
  LAYER M1 ;
        RECT 44.799 7.896 44.801 10.332 ;
  LAYER M1 ;
        RECT 44.879 7.896 44.881 10.332 ;
  LAYER M1 ;
        RECT 44.959 7.896 44.961 10.332 ;
  LAYER M1 ;
        RECT 45.039 7.896 45.041 10.332 ;
  LAYER M1 ;
        RECT 45.119 7.896 45.121 10.332 ;
  LAYER M1 ;
        RECT 45.199 7.896 45.201 10.332 ;
  LAYER M1 ;
        RECT 45.279 7.896 45.281 10.332 ;
  LAYER M1 ;
        RECT 45.359 7.896 45.361 10.332 ;
  LAYER M1 ;
        RECT 45.439 7.896 45.441 10.332 ;
  LAYER M2 ;
        RECT 43.12 10.331 45.52 10.333 ;
  LAYER M2 ;
        RECT 43.12 10.247 45.52 10.249 ;
  LAYER M2 ;
        RECT 43.12 10.163 45.52 10.165 ;
  LAYER M2 ;
        RECT 43.12 10.079 45.52 10.081 ;
  LAYER M2 ;
        RECT 43.12 9.995 45.52 9.997 ;
  LAYER M2 ;
        RECT 43.12 9.911 45.52 9.913 ;
  LAYER M2 ;
        RECT 43.12 9.827 45.52 9.829 ;
  LAYER M2 ;
        RECT 43.12 9.743 45.52 9.745 ;
  LAYER M2 ;
        RECT 43.12 9.659 45.52 9.661 ;
  LAYER M2 ;
        RECT 43.12 9.575 45.52 9.577 ;
  LAYER M2 ;
        RECT 43.12 9.491 45.52 9.493 ;
  LAYER M2 ;
        RECT 43.12 9.407 45.52 9.409 ;
  LAYER M2 ;
        RECT 43.12 9.3235 45.52 9.3255 ;
  LAYER M2 ;
        RECT 43.12 9.239 45.52 9.241 ;
  LAYER M2 ;
        RECT 43.12 9.155 45.52 9.157 ;
  LAYER M2 ;
        RECT 43.12 9.071 45.52 9.073 ;
  LAYER M2 ;
        RECT 43.12 8.987 45.52 8.989 ;
  LAYER M2 ;
        RECT 43.12 8.903 45.52 8.905 ;
  LAYER M2 ;
        RECT 43.12 8.819 45.52 8.821 ;
  LAYER M2 ;
        RECT 43.12 8.735 45.52 8.737 ;
  LAYER M2 ;
        RECT 43.12 8.651 45.52 8.653 ;
  LAYER M2 ;
        RECT 43.12 8.567 45.52 8.569 ;
  LAYER M2 ;
        RECT 43.12 8.483 45.52 8.485 ;
  LAYER M2 ;
        RECT 43.12 8.399 45.52 8.401 ;
  LAYER M2 ;
        RECT 43.12 8.315 45.52 8.317 ;
  LAYER M2 ;
        RECT 43.12 8.231 45.52 8.233 ;
  LAYER M2 ;
        RECT 43.12 8.147 45.52 8.149 ;
  LAYER M2 ;
        RECT 43.12 8.063 45.52 8.065 ;
  LAYER M2 ;
        RECT 43.12 7.979 45.52 7.981 ;
  LAYER M1 ;
        RECT 43.104 4.92 43.136 7.428 ;
  LAYER M1 ;
        RECT 43.168 4.92 43.2 7.428 ;
  LAYER M1 ;
        RECT 43.232 4.92 43.264 7.428 ;
  LAYER M1 ;
        RECT 43.296 4.92 43.328 7.428 ;
  LAYER M1 ;
        RECT 43.36 4.92 43.392 7.428 ;
  LAYER M1 ;
        RECT 43.424 4.92 43.456 7.428 ;
  LAYER M1 ;
        RECT 43.488 4.92 43.52 7.428 ;
  LAYER M1 ;
        RECT 43.552 4.92 43.584 7.428 ;
  LAYER M1 ;
        RECT 43.616 4.92 43.648 7.428 ;
  LAYER M1 ;
        RECT 43.68 4.92 43.712 7.428 ;
  LAYER M1 ;
        RECT 43.744 4.92 43.776 7.428 ;
  LAYER M1 ;
        RECT 43.808 4.92 43.84 7.428 ;
  LAYER M1 ;
        RECT 43.872 4.92 43.904 7.428 ;
  LAYER M1 ;
        RECT 43.936 4.92 43.968 7.428 ;
  LAYER M1 ;
        RECT 44 4.92 44.032 7.428 ;
  LAYER M1 ;
        RECT 44.064 4.92 44.096 7.428 ;
  LAYER M1 ;
        RECT 44.128 4.92 44.16 7.428 ;
  LAYER M1 ;
        RECT 44.192 4.92 44.224 7.428 ;
  LAYER M1 ;
        RECT 44.256 4.92 44.288 7.428 ;
  LAYER M1 ;
        RECT 44.32 4.92 44.352 7.428 ;
  LAYER M1 ;
        RECT 44.384 4.92 44.416 7.428 ;
  LAYER M1 ;
        RECT 44.448 4.92 44.48 7.428 ;
  LAYER M1 ;
        RECT 44.512 4.92 44.544 7.428 ;
  LAYER M1 ;
        RECT 44.576 4.92 44.608 7.428 ;
  LAYER M1 ;
        RECT 44.64 4.92 44.672 7.428 ;
  LAYER M1 ;
        RECT 44.704 4.92 44.736 7.428 ;
  LAYER M1 ;
        RECT 44.768 4.92 44.8 7.428 ;
  LAYER M1 ;
        RECT 44.832 4.92 44.864 7.428 ;
  LAYER M1 ;
        RECT 44.896 4.92 44.928 7.428 ;
  LAYER M1 ;
        RECT 44.96 4.92 44.992 7.428 ;
  LAYER M1 ;
        RECT 45.024 4.92 45.056 7.428 ;
  LAYER M1 ;
        RECT 45.088 4.92 45.12 7.428 ;
  LAYER M1 ;
        RECT 45.152 4.92 45.184 7.428 ;
  LAYER M1 ;
        RECT 45.216 4.92 45.248 7.428 ;
  LAYER M1 ;
        RECT 45.28 4.92 45.312 7.428 ;
  LAYER M1 ;
        RECT 45.344 4.92 45.376 7.428 ;
  LAYER M1 ;
        RECT 45.408 4.92 45.44 7.428 ;
  LAYER M2 ;
        RECT 43.084 7.312 45.556 7.344 ;
  LAYER M2 ;
        RECT 43.084 7.248 45.556 7.28 ;
  LAYER M2 ;
        RECT 43.084 7.184 45.556 7.216 ;
  LAYER M2 ;
        RECT 43.084 7.12 45.556 7.152 ;
  LAYER M2 ;
        RECT 43.084 7.056 45.556 7.088 ;
  LAYER M2 ;
        RECT 43.084 6.992 45.556 7.024 ;
  LAYER M2 ;
        RECT 43.084 6.928 45.556 6.96 ;
  LAYER M2 ;
        RECT 43.084 6.864 45.556 6.896 ;
  LAYER M2 ;
        RECT 43.084 6.8 45.556 6.832 ;
  LAYER M2 ;
        RECT 43.084 6.736 45.556 6.768 ;
  LAYER M2 ;
        RECT 43.084 6.672 45.556 6.704 ;
  LAYER M2 ;
        RECT 43.084 6.608 45.556 6.64 ;
  LAYER M2 ;
        RECT 43.084 6.544 45.556 6.576 ;
  LAYER M2 ;
        RECT 43.084 6.48 45.556 6.512 ;
  LAYER M2 ;
        RECT 43.084 6.416 45.556 6.448 ;
  LAYER M2 ;
        RECT 43.084 6.352 45.556 6.384 ;
  LAYER M2 ;
        RECT 43.084 6.288 45.556 6.32 ;
  LAYER M2 ;
        RECT 43.084 6.224 45.556 6.256 ;
  LAYER M2 ;
        RECT 43.084 6.16 45.556 6.192 ;
  LAYER M2 ;
        RECT 43.084 6.096 45.556 6.128 ;
  LAYER M2 ;
        RECT 43.084 6.032 45.556 6.064 ;
  LAYER M2 ;
        RECT 43.084 5.968 45.556 6 ;
  LAYER M2 ;
        RECT 43.084 5.904 45.556 5.936 ;
  LAYER M2 ;
        RECT 43.084 5.84 45.556 5.872 ;
  LAYER M2 ;
        RECT 43.084 5.776 45.556 5.808 ;
  LAYER M2 ;
        RECT 43.084 5.712 45.556 5.744 ;
  LAYER M2 ;
        RECT 43.084 5.648 45.556 5.68 ;
  LAYER M2 ;
        RECT 43.084 5.584 45.556 5.616 ;
  LAYER M2 ;
        RECT 43.084 5.52 45.556 5.552 ;
  LAYER M2 ;
        RECT 43.084 5.456 45.556 5.488 ;
  LAYER M2 ;
        RECT 43.084 5.392 45.556 5.424 ;
  LAYER M2 ;
        RECT 43.084 5.328 45.556 5.36 ;
  LAYER M2 ;
        RECT 43.084 5.264 45.556 5.296 ;
  LAYER M2 ;
        RECT 43.084 5.2 45.556 5.232 ;
  LAYER M2 ;
        RECT 43.084 5.136 45.556 5.168 ;
  LAYER M2 ;
        RECT 43.084 5.072 45.556 5.104 ;
  LAYER M3 ;
        RECT 43.104 4.92 43.136 7.428 ;
  LAYER M3 ;
        RECT 43.168 4.92 43.2 7.428 ;
  LAYER M3 ;
        RECT 43.232 4.92 43.264 7.428 ;
  LAYER M3 ;
        RECT 43.296 4.92 43.328 7.428 ;
  LAYER M3 ;
        RECT 43.36 4.92 43.392 7.428 ;
  LAYER M3 ;
        RECT 43.424 4.92 43.456 7.428 ;
  LAYER M3 ;
        RECT 43.488 4.92 43.52 7.428 ;
  LAYER M3 ;
        RECT 43.552 4.92 43.584 7.428 ;
  LAYER M3 ;
        RECT 43.616 4.92 43.648 7.428 ;
  LAYER M3 ;
        RECT 43.68 4.92 43.712 7.428 ;
  LAYER M3 ;
        RECT 43.744 4.92 43.776 7.428 ;
  LAYER M3 ;
        RECT 43.808 4.92 43.84 7.428 ;
  LAYER M3 ;
        RECT 43.872 4.92 43.904 7.428 ;
  LAYER M3 ;
        RECT 43.936 4.92 43.968 7.428 ;
  LAYER M3 ;
        RECT 44 4.92 44.032 7.428 ;
  LAYER M3 ;
        RECT 44.064 4.92 44.096 7.428 ;
  LAYER M3 ;
        RECT 44.128 4.92 44.16 7.428 ;
  LAYER M3 ;
        RECT 44.192 4.92 44.224 7.428 ;
  LAYER M3 ;
        RECT 44.256 4.92 44.288 7.428 ;
  LAYER M3 ;
        RECT 44.32 4.92 44.352 7.428 ;
  LAYER M3 ;
        RECT 44.384 4.92 44.416 7.428 ;
  LAYER M3 ;
        RECT 44.448 4.92 44.48 7.428 ;
  LAYER M3 ;
        RECT 44.512 4.92 44.544 7.428 ;
  LAYER M3 ;
        RECT 44.576 4.92 44.608 7.428 ;
  LAYER M3 ;
        RECT 44.64 4.92 44.672 7.428 ;
  LAYER M3 ;
        RECT 44.704 4.92 44.736 7.428 ;
  LAYER M3 ;
        RECT 44.768 4.92 44.8 7.428 ;
  LAYER M3 ;
        RECT 44.832 4.92 44.864 7.428 ;
  LAYER M3 ;
        RECT 44.896 4.92 44.928 7.428 ;
  LAYER M3 ;
        RECT 44.96 4.92 44.992 7.428 ;
  LAYER M3 ;
        RECT 45.024 4.92 45.056 7.428 ;
  LAYER M3 ;
        RECT 45.088 4.92 45.12 7.428 ;
  LAYER M3 ;
        RECT 45.152 4.92 45.184 7.428 ;
  LAYER M3 ;
        RECT 45.216 4.92 45.248 7.428 ;
  LAYER M3 ;
        RECT 45.28 4.92 45.312 7.428 ;
  LAYER M3 ;
        RECT 45.344 4.92 45.376 7.428 ;
  LAYER M3 ;
        RECT 45.408 4.92 45.44 7.428 ;
  LAYER M3 ;
        RECT 45.504 4.92 45.536 7.428 ;
  LAYER M1 ;
        RECT 43.119 4.956 43.121 7.392 ;
  LAYER M1 ;
        RECT 43.199 4.956 43.201 7.392 ;
  LAYER M1 ;
        RECT 43.279 4.956 43.281 7.392 ;
  LAYER M1 ;
        RECT 43.359 4.956 43.361 7.392 ;
  LAYER M1 ;
        RECT 43.439 4.956 43.441 7.392 ;
  LAYER M1 ;
        RECT 43.519 4.956 43.521 7.392 ;
  LAYER M1 ;
        RECT 43.599 4.956 43.601 7.392 ;
  LAYER M1 ;
        RECT 43.679 4.956 43.681 7.392 ;
  LAYER M1 ;
        RECT 43.759 4.956 43.761 7.392 ;
  LAYER M1 ;
        RECT 43.839 4.956 43.841 7.392 ;
  LAYER M1 ;
        RECT 43.919 4.956 43.921 7.392 ;
  LAYER M1 ;
        RECT 43.999 4.956 44.001 7.392 ;
  LAYER M1 ;
        RECT 44.079 4.956 44.081 7.392 ;
  LAYER M1 ;
        RECT 44.159 4.956 44.161 7.392 ;
  LAYER M1 ;
        RECT 44.239 4.956 44.241 7.392 ;
  LAYER M1 ;
        RECT 44.319 4.956 44.321 7.392 ;
  LAYER M1 ;
        RECT 44.399 4.956 44.401 7.392 ;
  LAYER M1 ;
        RECT 44.479 4.956 44.481 7.392 ;
  LAYER M1 ;
        RECT 44.559 4.956 44.561 7.392 ;
  LAYER M1 ;
        RECT 44.639 4.956 44.641 7.392 ;
  LAYER M1 ;
        RECT 44.719 4.956 44.721 7.392 ;
  LAYER M1 ;
        RECT 44.799 4.956 44.801 7.392 ;
  LAYER M1 ;
        RECT 44.879 4.956 44.881 7.392 ;
  LAYER M1 ;
        RECT 44.959 4.956 44.961 7.392 ;
  LAYER M1 ;
        RECT 45.039 4.956 45.041 7.392 ;
  LAYER M1 ;
        RECT 45.119 4.956 45.121 7.392 ;
  LAYER M1 ;
        RECT 45.199 4.956 45.201 7.392 ;
  LAYER M1 ;
        RECT 45.279 4.956 45.281 7.392 ;
  LAYER M1 ;
        RECT 45.359 4.956 45.361 7.392 ;
  LAYER M1 ;
        RECT 45.439 4.956 45.441 7.392 ;
  LAYER M2 ;
        RECT 43.12 7.391 45.52 7.393 ;
  LAYER M2 ;
        RECT 43.12 7.307 45.52 7.309 ;
  LAYER M2 ;
        RECT 43.12 7.223 45.52 7.225 ;
  LAYER M2 ;
        RECT 43.12 7.139 45.52 7.141 ;
  LAYER M2 ;
        RECT 43.12 7.055 45.52 7.057 ;
  LAYER M2 ;
        RECT 43.12 6.971 45.52 6.973 ;
  LAYER M2 ;
        RECT 43.12 6.887 45.52 6.889 ;
  LAYER M2 ;
        RECT 43.12 6.803 45.52 6.805 ;
  LAYER M2 ;
        RECT 43.12 6.719 45.52 6.721 ;
  LAYER M2 ;
        RECT 43.12 6.635 45.52 6.637 ;
  LAYER M2 ;
        RECT 43.12 6.551 45.52 6.553 ;
  LAYER M2 ;
        RECT 43.12 6.467 45.52 6.469 ;
  LAYER M2 ;
        RECT 43.12 6.3835 45.52 6.3855 ;
  LAYER M2 ;
        RECT 43.12 6.299 45.52 6.301 ;
  LAYER M2 ;
        RECT 43.12 6.215 45.52 6.217 ;
  LAYER M2 ;
        RECT 43.12 6.131 45.52 6.133 ;
  LAYER M2 ;
        RECT 43.12 6.047 45.52 6.049 ;
  LAYER M2 ;
        RECT 43.12 5.963 45.52 5.965 ;
  LAYER M2 ;
        RECT 43.12 5.879 45.52 5.881 ;
  LAYER M2 ;
        RECT 43.12 5.795 45.52 5.797 ;
  LAYER M2 ;
        RECT 43.12 5.711 45.52 5.713 ;
  LAYER M2 ;
        RECT 43.12 5.627 45.52 5.629 ;
  LAYER M2 ;
        RECT 43.12 5.543 45.52 5.545 ;
  LAYER M2 ;
        RECT 43.12 5.459 45.52 5.461 ;
  LAYER M2 ;
        RECT 43.12 5.375 45.52 5.377 ;
  LAYER M2 ;
        RECT 43.12 5.291 45.52 5.293 ;
  LAYER M2 ;
        RECT 43.12 5.207 45.52 5.209 ;
  LAYER M2 ;
        RECT 43.12 5.123 45.52 5.125 ;
  LAYER M2 ;
        RECT 43.12 5.039 45.52 5.041 ;
  LAYER M1 ;
        RECT 43.104 1.98 43.136 4.488 ;
  LAYER M1 ;
        RECT 43.168 1.98 43.2 4.488 ;
  LAYER M1 ;
        RECT 43.232 1.98 43.264 4.488 ;
  LAYER M1 ;
        RECT 43.296 1.98 43.328 4.488 ;
  LAYER M1 ;
        RECT 43.36 1.98 43.392 4.488 ;
  LAYER M1 ;
        RECT 43.424 1.98 43.456 4.488 ;
  LAYER M1 ;
        RECT 43.488 1.98 43.52 4.488 ;
  LAYER M1 ;
        RECT 43.552 1.98 43.584 4.488 ;
  LAYER M1 ;
        RECT 43.616 1.98 43.648 4.488 ;
  LAYER M1 ;
        RECT 43.68 1.98 43.712 4.488 ;
  LAYER M1 ;
        RECT 43.744 1.98 43.776 4.488 ;
  LAYER M1 ;
        RECT 43.808 1.98 43.84 4.488 ;
  LAYER M1 ;
        RECT 43.872 1.98 43.904 4.488 ;
  LAYER M1 ;
        RECT 43.936 1.98 43.968 4.488 ;
  LAYER M1 ;
        RECT 44 1.98 44.032 4.488 ;
  LAYER M1 ;
        RECT 44.064 1.98 44.096 4.488 ;
  LAYER M1 ;
        RECT 44.128 1.98 44.16 4.488 ;
  LAYER M1 ;
        RECT 44.192 1.98 44.224 4.488 ;
  LAYER M1 ;
        RECT 44.256 1.98 44.288 4.488 ;
  LAYER M1 ;
        RECT 44.32 1.98 44.352 4.488 ;
  LAYER M1 ;
        RECT 44.384 1.98 44.416 4.488 ;
  LAYER M1 ;
        RECT 44.448 1.98 44.48 4.488 ;
  LAYER M1 ;
        RECT 44.512 1.98 44.544 4.488 ;
  LAYER M1 ;
        RECT 44.576 1.98 44.608 4.488 ;
  LAYER M1 ;
        RECT 44.64 1.98 44.672 4.488 ;
  LAYER M1 ;
        RECT 44.704 1.98 44.736 4.488 ;
  LAYER M1 ;
        RECT 44.768 1.98 44.8 4.488 ;
  LAYER M1 ;
        RECT 44.832 1.98 44.864 4.488 ;
  LAYER M1 ;
        RECT 44.896 1.98 44.928 4.488 ;
  LAYER M1 ;
        RECT 44.96 1.98 44.992 4.488 ;
  LAYER M1 ;
        RECT 45.024 1.98 45.056 4.488 ;
  LAYER M1 ;
        RECT 45.088 1.98 45.12 4.488 ;
  LAYER M1 ;
        RECT 45.152 1.98 45.184 4.488 ;
  LAYER M1 ;
        RECT 45.216 1.98 45.248 4.488 ;
  LAYER M1 ;
        RECT 45.28 1.98 45.312 4.488 ;
  LAYER M1 ;
        RECT 45.344 1.98 45.376 4.488 ;
  LAYER M1 ;
        RECT 45.408 1.98 45.44 4.488 ;
  LAYER M2 ;
        RECT 43.084 4.372 45.556 4.404 ;
  LAYER M2 ;
        RECT 43.084 4.308 45.556 4.34 ;
  LAYER M2 ;
        RECT 43.084 4.244 45.556 4.276 ;
  LAYER M2 ;
        RECT 43.084 4.18 45.556 4.212 ;
  LAYER M2 ;
        RECT 43.084 4.116 45.556 4.148 ;
  LAYER M2 ;
        RECT 43.084 4.052 45.556 4.084 ;
  LAYER M2 ;
        RECT 43.084 3.988 45.556 4.02 ;
  LAYER M2 ;
        RECT 43.084 3.924 45.556 3.956 ;
  LAYER M2 ;
        RECT 43.084 3.86 45.556 3.892 ;
  LAYER M2 ;
        RECT 43.084 3.796 45.556 3.828 ;
  LAYER M2 ;
        RECT 43.084 3.732 45.556 3.764 ;
  LAYER M2 ;
        RECT 43.084 3.668 45.556 3.7 ;
  LAYER M2 ;
        RECT 43.084 3.604 45.556 3.636 ;
  LAYER M2 ;
        RECT 43.084 3.54 45.556 3.572 ;
  LAYER M2 ;
        RECT 43.084 3.476 45.556 3.508 ;
  LAYER M2 ;
        RECT 43.084 3.412 45.556 3.444 ;
  LAYER M2 ;
        RECT 43.084 3.348 45.556 3.38 ;
  LAYER M2 ;
        RECT 43.084 3.284 45.556 3.316 ;
  LAYER M2 ;
        RECT 43.084 3.22 45.556 3.252 ;
  LAYER M2 ;
        RECT 43.084 3.156 45.556 3.188 ;
  LAYER M2 ;
        RECT 43.084 3.092 45.556 3.124 ;
  LAYER M2 ;
        RECT 43.084 3.028 45.556 3.06 ;
  LAYER M2 ;
        RECT 43.084 2.964 45.556 2.996 ;
  LAYER M2 ;
        RECT 43.084 2.9 45.556 2.932 ;
  LAYER M2 ;
        RECT 43.084 2.836 45.556 2.868 ;
  LAYER M2 ;
        RECT 43.084 2.772 45.556 2.804 ;
  LAYER M2 ;
        RECT 43.084 2.708 45.556 2.74 ;
  LAYER M2 ;
        RECT 43.084 2.644 45.556 2.676 ;
  LAYER M2 ;
        RECT 43.084 2.58 45.556 2.612 ;
  LAYER M2 ;
        RECT 43.084 2.516 45.556 2.548 ;
  LAYER M2 ;
        RECT 43.084 2.452 45.556 2.484 ;
  LAYER M2 ;
        RECT 43.084 2.388 45.556 2.42 ;
  LAYER M2 ;
        RECT 43.084 2.324 45.556 2.356 ;
  LAYER M2 ;
        RECT 43.084 2.26 45.556 2.292 ;
  LAYER M2 ;
        RECT 43.084 2.196 45.556 2.228 ;
  LAYER M2 ;
        RECT 43.084 2.132 45.556 2.164 ;
  LAYER M3 ;
        RECT 43.104 1.98 43.136 4.488 ;
  LAYER M3 ;
        RECT 43.168 1.98 43.2 4.488 ;
  LAYER M3 ;
        RECT 43.232 1.98 43.264 4.488 ;
  LAYER M3 ;
        RECT 43.296 1.98 43.328 4.488 ;
  LAYER M3 ;
        RECT 43.36 1.98 43.392 4.488 ;
  LAYER M3 ;
        RECT 43.424 1.98 43.456 4.488 ;
  LAYER M3 ;
        RECT 43.488 1.98 43.52 4.488 ;
  LAYER M3 ;
        RECT 43.552 1.98 43.584 4.488 ;
  LAYER M3 ;
        RECT 43.616 1.98 43.648 4.488 ;
  LAYER M3 ;
        RECT 43.68 1.98 43.712 4.488 ;
  LAYER M3 ;
        RECT 43.744 1.98 43.776 4.488 ;
  LAYER M3 ;
        RECT 43.808 1.98 43.84 4.488 ;
  LAYER M3 ;
        RECT 43.872 1.98 43.904 4.488 ;
  LAYER M3 ;
        RECT 43.936 1.98 43.968 4.488 ;
  LAYER M3 ;
        RECT 44 1.98 44.032 4.488 ;
  LAYER M3 ;
        RECT 44.064 1.98 44.096 4.488 ;
  LAYER M3 ;
        RECT 44.128 1.98 44.16 4.488 ;
  LAYER M3 ;
        RECT 44.192 1.98 44.224 4.488 ;
  LAYER M3 ;
        RECT 44.256 1.98 44.288 4.488 ;
  LAYER M3 ;
        RECT 44.32 1.98 44.352 4.488 ;
  LAYER M3 ;
        RECT 44.384 1.98 44.416 4.488 ;
  LAYER M3 ;
        RECT 44.448 1.98 44.48 4.488 ;
  LAYER M3 ;
        RECT 44.512 1.98 44.544 4.488 ;
  LAYER M3 ;
        RECT 44.576 1.98 44.608 4.488 ;
  LAYER M3 ;
        RECT 44.64 1.98 44.672 4.488 ;
  LAYER M3 ;
        RECT 44.704 1.98 44.736 4.488 ;
  LAYER M3 ;
        RECT 44.768 1.98 44.8 4.488 ;
  LAYER M3 ;
        RECT 44.832 1.98 44.864 4.488 ;
  LAYER M3 ;
        RECT 44.896 1.98 44.928 4.488 ;
  LAYER M3 ;
        RECT 44.96 1.98 44.992 4.488 ;
  LAYER M3 ;
        RECT 45.024 1.98 45.056 4.488 ;
  LAYER M3 ;
        RECT 45.088 1.98 45.12 4.488 ;
  LAYER M3 ;
        RECT 45.152 1.98 45.184 4.488 ;
  LAYER M3 ;
        RECT 45.216 1.98 45.248 4.488 ;
  LAYER M3 ;
        RECT 45.28 1.98 45.312 4.488 ;
  LAYER M3 ;
        RECT 45.344 1.98 45.376 4.488 ;
  LAYER M3 ;
        RECT 45.408 1.98 45.44 4.488 ;
  LAYER M3 ;
        RECT 45.504 1.98 45.536 4.488 ;
  LAYER M1 ;
        RECT 43.119 2.016 43.121 4.452 ;
  LAYER M1 ;
        RECT 43.199 2.016 43.201 4.452 ;
  LAYER M1 ;
        RECT 43.279 2.016 43.281 4.452 ;
  LAYER M1 ;
        RECT 43.359 2.016 43.361 4.452 ;
  LAYER M1 ;
        RECT 43.439 2.016 43.441 4.452 ;
  LAYER M1 ;
        RECT 43.519 2.016 43.521 4.452 ;
  LAYER M1 ;
        RECT 43.599 2.016 43.601 4.452 ;
  LAYER M1 ;
        RECT 43.679 2.016 43.681 4.452 ;
  LAYER M1 ;
        RECT 43.759 2.016 43.761 4.452 ;
  LAYER M1 ;
        RECT 43.839 2.016 43.841 4.452 ;
  LAYER M1 ;
        RECT 43.919 2.016 43.921 4.452 ;
  LAYER M1 ;
        RECT 43.999 2.016 44.001 4.452 ;
  LAYER M1 ;
        RECT 44.079 2.016 44.081 4.452 ;
  LAYER M1 ;
        RECT 44.159 2.016 44.161 4.452 ;
  LAYER M1 ;
        RECT 44.239 2.016 44.241 4.452 ;
  LAYER M1 ;
        RECT 44.319 2.016 44.321 4.452 ;
  LAYER M1 ;
        RECT 44.399 2.016 44.401 4.452 ;
  LAYER M1 ;
        RECT 44.479 2.016 44.481 4.452 ;
  LAYER M1 ;
        RECT 44.559 2.016 44.561 4.452 ;
  LAYER M1 ;
        RECT 44.639 2.016 44.641 4.452 ;
  LAYER M1 ;
        RECT 44.719 2.016 44.721 4.452 ;
  LAYER M1 ;
        RECT 44.799 2.016 44.801 4.452 ;
  LAYER M1 ;
        RECT 44.879 2.016 44.881 4.452 ;
  LAYER M1 ;
        RECT 44.959 2.016 44.961 4.452 ;
  LAYER M1 ;
        RECT 45.039 2.016 45.041 4.452 ;
  LAYER M1 ;
        RECT 45.119 2.016 45.121 4.452 ;
  LAYER M1 ;
        RECT 45.199 2.016 45.201 4.452 ;
  LAYER M1 ;
        RECT 45.279 2.016 45.281 4.452 ;
  LAYER M1 ;
        RECT 45.359 2.016 45.361 4.452 ;
  LAYER M1 ;
        RECT 45.439 2.016 45.441 4.452 ;
  LAYER M2 ;
        RECT 43.12 4.451 45.52 4.453 ;
  LAYER M2 ;
        RECT 43.12 4.367 45.52 4.369 ;
  LAYER M2 ;
        RECT 43.12 4.283 45.52 4.285 ;
  LAYER M2 ;
        RECT 43.12 4.199 45.52 4.201 ;
  LAYER M2 ;
        RECT 43.12 4.115 45.52 4.117 ;
  LAYER M2 ;
        RECT 43.12 4.031 45.52 4.033 ;
  LAYER M2 ;
        RECT 43.12 3.947 45.52 3.949 ;
  LAYER M2 ;
        RECT 43.12 3.863 45.52 3.865 ;
  LAYER M2 ;
        RECT 43.12 3.779 45.52 3.781 ;
  LAYER M2 ;
        RECT 43.12 3.695 45.52 3.697 ;
  LAYER M2 ;
        RECT 43.12 3.611 45.52 3.613 ;
  LAYER M2 ;
        RECT 43.12 3.527 45.52 3.529 ;
  LAYER M2 ;
        RECT 43.12 3.4435 45.52 3.4455 ;
  LAYER M2 ;
        RECT 43.12 3.359 45.52 3.361 ;
  LAYER M2 ;
        RECT 43.12 3.275 45.52 3.277 ;
  LAYER M2 ;
        RECT 43.12 3.191 45.52 3.193 ;
  LAYER M2 ;
        RECT 43.12 3.107 45.52 3.109 ;
  LAYER M2 ;
        RECT 43.12 3.023 45.52 3.025 ;
  LAYER M2 ;
        RECT 43.12 2.939 45.52 2.941 ;
  LAYER M2 ;
        RECT 43.12 2.855 45.52 2.857 ;
  LAYER M2 ;
        RECT 43.12 2.771 45.52 2.773 ;
  LAYER M2 ;
        RECT 43.12 2.687 45.52 2.689 ;
  LAYER M2 ;
        RECT 43.12 2.603 45.52 2.605 ;
  LAYER M2 ;
        RECT 43.12 2.519 45.52 2.521 ;
  LAYER M2 ;
        RECT 43.12 2.435 45.52 2.437 ;
  LAYER M2 ;
        RECT 43.12 2.351 45.52 2.353 ;
  LAYER M2 ;
        RECT 43.12 2.267 45.52 2.269 ;
  LAYER M2 ;
        RECT 43.12 2.183 45.52 2.185 ;
  LAYER M2 ;
        RECT 43.12 2.099 45.52 2.101 ;
  LAYER M1 ;
        RECT 24.224 11.892 24.256 11.964 ;
  LAYER M2 ;
        RECT 24.204 11.912 24.276 11.944 ;
  LAYER M2 ;
        RECT 24.24 11.912 24.56 11.944 ;
  LAYER M1 ;
        RECT 24.544 11.892 24.576 11.964 ;
  LAYER M2 ;
        RECT 24.524 11.912 24.596 11.944 ;
  LAYER M1 ;
        RECT 27.104 14.832 27.136 14.904 ;
  LAYER M2 ;
        RECT 27.084 14.852 27.156 14.884 ;
  LAYER M1 ;
        RECT 27.104 14.868 27.136 15.036 ;
  LAYER M1 ;
        RECT 27.104 15 27.136 15.072 ;
  LAYER M2 ;
        RECT 27.084 15.02 27.156 15.052 ;
  LAYER M2 ;
        RECT 24.56 15.02 27.12 15.052 ;
  LAYER M1 ;
        RECT 24.544 15 24.576 15.072 ;
  LAYER M2 ;
        RECT 24.524 15.02 24.596 15.052 ;
  LAYER M1 ;
        RECT 24.544 18.276 24.576 18.348 ;
  LAYER M2 ;
        RECT 24.524 18.296 24.596 18.328 ;
  LAYER M1 ;
        RECT 24.544 18.144 24.576 18.312 ;
  LAYER M1 ;
        RECT 24.544 11.928 24.576 18.144 ;
  LAYER M1 ;
        RECT 21.344 11.892 21.376 11.964 ;
  LAYER M2 ;
        RECT 21.324 11.912 21.396 11.944 ;
  LAYER M2 ;
        RECT 21.36 11.912 21.68 11.944 ;
  LAYER M1 ;
        RECT 21.664 11.892 21.696 11.964 ;
  LAYER M2 ;
        RECT 21.644 11.912 21.716 11.944 ;
  LAYER M1 ;
        RECT 21.664 18.276 21.696 18.348 ;
  LAYER M2 ;
        RECT 21.644 18.296 21.716 18.328 ;
  LAYER M1 ;
        RECT 21.664 18.144 21.696 18.312 ;
  LAYER M1 ;
        RECT 21.664 11.928 21.696 18.144 ;
  LAYER M2 ;
        RECT 21.68 18.296 24.56 18.328 ;
  LAYER M1 ;
        RECT 27.104 11.892 27.136 11.964 ;
  LAYER M2 ;
        RECT 27.084 11.912 27.156 11.944 ;
  LAYER M2 ;
        RECT 27.12 11.912 27.44 11.944 ;
  LAYER M1 ;
        RECT 27.424 11.892 27.456 11.964 ;
  LAYER M2 ;
        RECT 27.404 11.912 27.476 11.944 ;
  LAYER M1 ;
        RECT 27.424 18.444 27.456 18.516 ;
  LAYER M2 ;
        RECT 27.404 18.464 27.476 18.496 ;
  LAYER M1 ;
        RECT 27.424 18.144 27.456 18.48 ;
  LAYER M1 ;
        RECT 27.424 11.928 27.456 18.144 ;
  LAYER M1 ;
        RECT 21.344 14.832 21.376 14.904 ;
  LAYER M2 ;
        RECT 21.324 14.852 21.396 14.884 ;
  LAYER M1 ;
        RECT 21.344 14.868 21.376 15.036 ;
  LAYER M1 ;
        RECT 21.344 15 21.376 15.072 ;
  LAYER M2 ;
        RECT 21.324 15.02 21.396 15.052 ;
  LAYER M2 ;
        RECT 18.8 15.02 21.36 15.052 ;
  LAYER M1 ;
        RECT 18.784 15 18.816 15.072 ;
  LAYER M2 ;
        RECT 18.764 15.02 18.836 15.052 ;
  LAYER M1 ;
        RECT 18.784 18.444 18.816 18.516 ;
  LAYER M2 ;
        RECT 18.764 18.464 18.836 18.496 ;
  LAYER M1 ;
        RECT 18.784 18.144 18.816 18.48 ;
  LAYER M1 ;
        RECT 18.784 15.036 18.816 18.144 ;
  LAYER M2 ;
        RECT 18.8 18.464 27.44 18.496 ;
  LAYER M1 ;
        RECT 24.224 14.832 24.256 14.904 ;
  LAYER M2 ;
        RECT 24.204 14.852 24.276 14.884 ;
  LAYER M2 ;
        RECT 21.36 14.852 24.24 14.884 ;
  LAYER M1 ;
        RECT 21.344 14.832 21.376 14.904 ;
  LAYER M2 ;
        RECT 21.324 14.852 21.396 14.884 ;
  LAYER M1 ;
        RECT 29.984 17.772 30.016 17.844 ;
  LAYER M2 ;
        RECT 29.964 17.792 30.036 17.824 ;
  LAYER M2 ;
        RECT 30 17.792 30.32 17.824 ;
  LAYER M1 ;
        RECT 30.304 17.772 30.336 17.844 ;
  LAYER M2 ;
        RECT 30.284 17.792 30.356 17.824 ;
  LAYER M1 ;
        RECT 29.984 14.832 30.016 14.904 ;
  LAYER M2 ;
        RECT 29.964 14.852 30.036 14.884 ;
  LAYER M2 ;
        RECT 30 14.852 30.32 14.884 ;
  LAYER M1 ;
        RECT 30.304 14.832 30.336 14.904 ;
  LAYER M2 ;
        RECT 30.284 14.852 30.356 14.884 ;
  LAYER M1 ;
        RECT 29.984 11.892 30.016 11.964 ;
  LAYER M2 ;
        RECT 29.964 11.912 30.036 11.944 ;
  LAYER M2 ;
        RECT 30 11.912 30.32 11.944 ;
  LAYER M1 ;
        RECT 30.304 11.892 30.336 11.964 ;
  LAYER M2 ;
        RECT 30.284 11.912 30.356 11.944 ;
  LAYER M1 ;
        RECT 29.984 8.952 30.016 9.024 ;
  LAYER M2 ;
        RECT 29.964 8.972 30.036 9.004 ;
  LAYER M2 ;
        RECT 30 8.972 30.32 9.004 ;
  LAYER M1 ;
        RECT 30.304 8.952 30.336 9.024 ;
  LAYER M2 ;
        RECT 30.284 8.972 30.356 9.004 ;
  LAYER M1 ;
        RECT 30.304 18.612 30.336 18.684 ;
  LAYER M2 ;
        RECT 30.284 18.632 30.356 18.664 ;
  LAYER M1 ;
        RECT 30.304 18.144 30.336 18.648 ;
  LAYER M1 ;
        RECT 30.304 8.988 30.336 18.144 ;
  LAYER M1 ;
        RECT 18.464 17.772 18.496 17.844 ;
  LAYER M2 ;
        RECT 18.444 17.792 18.516 17.824 ;
  LAYER M1 ;
        RECT 18.464 17.808 18.496 17.976 ;
  LAYER M1 ;
        RECT 18.464 17.94 18.496 18.012 ;
  LAYER M2 ;
        RECT 18.444 17.96 18.516 17.992 ;
  LAYER M2 ;
        RECT 15.92 17.96 18.48 17.992 ;
  LAYER M1 ;
        RECT 15.904 17.94 15.936 18.012 ;
  LAYER M2 ;
        RECT 15.884 17.96 15.956 17.992 ;
  LAYER M1 ;
        RECT 18.464 14.832 18.496 14.904 ;
  LAYER M2 ;
        RECT 18.444 14.852 18.516 14.884 ;
  LAYER M1 ;
        RECT 18.464 14.868 18.496 15.036 ;
  LAYER M1 ;
        RECT 18.464 15 18.496 15.072 ;
  LAYER M2 ;
        RECT 18.444 15.02 18.516 15.052 ;
  LAYER M2 ;
        RECT 15.92 15.02 18.48 15.052 ;
  LAYER M1 ;
        RECT 15.904 15 15.936 15.072 ;
  LAYER M2 ;
        RECT 15.884 15.02 15.956 15.052 ;
  LAYER M1 ;
        RECT 18.464 11.892 18.496 11.964 ;
  LAYER M2 ;
        RECT 18.444 11.912 18.516 11.944 ;
  LAYER M1 ;
        RECT 18.464 11.928 18.496 12.096 ;
  LAYER M1 ;
        RECT 18.464 12.06 18.496 12.132 ;
  LAYER M2 ;
        RECT 18.444 12.08 18.516 12.112 ;
  LAYER M2 ;
        RECT 15.92 12.08 18.48 12.112 ;
  LAYER M1 ;
        RECT 15.904 12.06 15.936 12.132 ;
  LAYER M2 ;
        RECT 15.884 12.08 15.956 12.112 ;
  LAYER M1 ;
        RECT 18.464 8.952 18.496 9.024 ;
  LAYER M2 ;
        RECT 18.444 8.972 18.516 9.004 ;
  LAYER M1 ;
        RECT 18.464 8.988 18.496 9.156 ;
  LAYER M1 ;
        RECT 18.464 9.12 18.496 9.192 ;
  LAYER M2 ;
        RECT 18.444 9.14 18.516 9.172 ;
  LAYER M2 ;
        RECT 15.92 9.14 18.48 9.172 ;
  LAYER M1 ;
        RECT 15.904 9.12 15.936 9.192 ;
  LAYER M2 ;
        RECT 15.884 9.14 15.956 9.172 ;
  LAYER M1 ;
        RECT 15.904 18.612 15.936 18.684 ;
  LAYER M2 ;
        RECT 15.884 18.632 15.956 18.664 ;
  LAYER M1 ;
        RECT 15.904 18.144 15.936 18.648 ;
  LAYER M1 ;
        RECT 15.904 9.156 15.936 18.144 ;
  LAYER M2 ;
        RECT 15.92 18.632 30.32 18.664 ;
  LAYER M1 ;
        RECT 27.104 17.772 27.136 17.844 ;
  LAYER M2 ;
        RECT 27.084 17.792 27.156 17.824 ;
  LAYER M2 ;
        RECT 27.12 17.792 30 17.824 ;
  LAYER M1 ;
        RECT 29.984 17.772 30.016 17.844 ;
  LAYER M2 ;
        RECT 29.964 17.792 30.036 17.824 ;
  LAYER M1 ;
        RECT 27.104 8.952 27.136 9.024 ;
  LAYER M2 ;
        RECT 27.084 8.972 27.156 9.004 ;
  LAYER M2 ;
        RECT 27.12 8.972 30 9.004 ;
  LAYER M1 ;
        RECT 29.984 8.952 30.016 9.024 ;
  LAYER M2 ;
        RECT 29.964 8.972 30.036 9.004 ;
  LAYER M1 ;
        RECT 24.224 8.952 24.256 9.024 ;
  LAYER M2 ;
        RECT 24.204 8.972 24.276 9.004 ;
  LAYER M2 ;
        RECT 24.24 8.972 27.12 9.004 ;
  LAYER M1 ;
        RECT 27.104 8.952 27.136 9.024 ;
  LAYER M2 ;
        RECT 27.084 8.972 27.156 9.004 ;
  LAYER M1 ;
        RECT 21.344 8.952 21.376 9.024 ;
  LAYER M2 ;
        RECT 21.324 8.972 21.396 9.004 ;
  LAYER M2 ;
        RECT 21.36 8.972 24.24 9.004 ;
  LAYER M1 ;
        RECT 24.224 8.952 24.256 9.024 ;
  LAYER M2 ;
        RECT 24.204 8.972 24.276 9.004 ;
  LAYER M1 ;
        RECT 21.344 17.772 21.376 17.844 ;
  LAYER M2 ;
        RECT 21.324 17.792 21.396 17.824 ;
  LAYER M2 ;
        RECT 18.48 17.792 21.36 17.824 ;
  LAYER M1 ;
        RECT 18.464 17.772 18.496 17.844 ;
  LAYER M2 ;
        RECT 18.444 17.792 18.516 17.824 ;
  LAYER M1 ;
        RECT 24.224 17.772 24.256 17.844 ;
  LAYER M2 ;
        RECT 24.204 17.792 24.276 17.824 ;
  LAYER M2 ;
        RECT 21.36 17.792 24.24 17.824 ;
  LAYER M1 ;
        RECT 21.344 17.772 21.376 17.844 ;
  LAYER M2 ;
        RECT 21.324 17.792 21.396 17.824 ;
  LAYER M1 ;
        RECT 21.824 9.456 21.856 9.528 ;
  LAYER M2 ;
        RECT 21.804 9.476 21.876 9.508 ;
  LAYER M2 ;
        RECT 21.84 9.476 24.4 9.508 ;
  LAYER M1 ;
        RECT 24.384 9.456 24.416 9.528 ;
  LAYER M2 ;
        RECT 24.364 9.476 24.436 9.508 ;
  LAYER M1 ;
        RECT 24.704 12.396 24.736 12.468 ;
  LAYER M2 ;
        RECT 24.684 12.416 24.756 12.448 ;
  LAYER M1 ;
        RECT 24.704 12.264 24.736 12.432 ;
  LAYER M1 ;
        RECT 24.704 12.228 24.736 12.3 ;
  LAYER M2 ;
        RECT 24.684 12.248 24.756 12.28 ;
  LAYER M2 ;
        RECT 24.4 12.248 24.72 12.28 ;
  LAYER M1 ;
        RECT 24.384 12.228 24.416 12.3 ;
  LAYER M2 ;
        RECT 24.364 12.248 24.436 12.28 ;
  LAYER M1 ;
        RECT 24.384 6.012 24.416 6.084 ;
  LAYER M2 ;
        RECT 24.364 6.032 24.436 6.064 ;
  LAYER M1 ;
        RECT 24.384 6.048 24.416 6.216 ;
  LAYER M1 ;
        RECT 24.384 6.216 24.416 12.264 ;
  LAYER M1 ;
        RECT 18.944 9.456 18.976 9.528 ;
  LAYER M2 ;
        RECT 18.924 9.476 18.996 9.508 ;
  LAYER M2 ;
        RECT 18.96 9.476 21.52 9.508 ;
  LAYER M1 ;
        RECT 21.504 9.456 21.536 9.528 ;
  LAYER M2 ;
        RECT 21.484 9.476 21.556 9.508 ;
  LAYER M1 ;
        RECT 21.504 6.012 21.536 6.084 ;
  LAYER M2 ;
        RECT 21.484 6.032 21.556 6.064 ;
  LAYER M1 ;
        RECT 21.504 6.048 21.536 6.216 ;
  LAYER M1 ;
        RECT 21.504 6.216 21.536 9.492 ;
  LAYER M2 ;
        RECT 21.52 6.032 24.4 6.064 ;
  LAYER M1 ;
        RECT 24.704 9.456 24.736 9.528 ;
  LAYER M2 ;
        RECT 24.684 9.476 24.756 9.508 ;
  LAYER M2 ;
        RECT 24.72 9.476 27.28 9.508 ;
  LAYER M1 ;
        RECT 27.264 9.456 27.296 9.528 ;
  LAYER M2 ;
        RECT 27.244 9.476 27.316 9.508 ;
  LAYER M1 ;
        RECT 27.264 5.844 27.296 5.916 ;
  LAYER M2 ;
        RECT 27.244 5.864 27.316 5.896 ;
  LAYER M1 ;
        RECT 27.264 5.88 27.296 6.216 ;
  LAYER M1 ;
        RECT 27.264 6.216 27.296 9.492 ;
  LAYER M1 ;
        RECT 18.944 12.396 18.976 12.468 ;
  LAYER M2 ;
        RECT 18.924 12.416 18.996 12.448 ;
  LAYER M1 ;
        RECT 18.944 12.264 18.976 12.432 ;
  LAYER M1 ;
        RECT 18.944 12.228 18.976 12.3 ;
  LAYER M2 ;
        RECT 18.924 12.248 18.996 12.28 ;
  LAYER M2 ;
        RECT 18.64 12.248 18.96 12.28 ;
  LAYER M1 ;
        RECT 18.624 12.228 18.656 12.3 ;
  LAYER M2 ;
        RECT 18.604 12.248 18.676 12.28 ;
  LAYER M1 ;
        RECT 18.624 5.844 18.656 5.916 ;
  LAYER M2 ;
        RECT 18.604 5.864 18.676 5.896 ;
  LAYER M1 ;
        RECT 18.624 5.88 18.656 6.216 ;
  LAYER M1 ;
        RECT 18.624 6.216 18.656 12.264 ;
  LAYER M2 ;
        RECT 18.64 5.864 27.28 5.896 ;
  LAYER M1 ;
        RECT 21.824 12.396 21.856 12.468 ;
  LAYER M2 ;
        RECT 21.804 12.416 21.876 12.448 ;
  LAYER M2 ;
        RECT 18.96 12.416 21.84 12.448 ;
  LAYER M1 ;
        RECT 18.944 12.396 18.976 12.468 ;
  LAYER M2 ;
        RECT 18.924 12.416 18.996 12.448 ;
  LAYER M1 ;
        RECT 27.584 15.336 27.616 15.408 ;
  LAYER M2 ;
        RECT 27.564 15.356 27.636 15.388 ;
  LAYER M2 ;
        RECT 27.6 15.356 30.16 15.388 ;
  LAYER M1 ;
        RECT 30.144 15.336 30.176 15.408 ;
  LAYER M2 ;
        RECT 30.124 15.356 30.196 15.388 ;
  LAYER M1 ;
        RECT 27.584 12.396 27.616 12.468 ;
  LAYER M2 ;
        RECT 27.564 12.416 27.636 12.448 ;
  LAYER M2 ;
        RECT 27.6 12.416 30.16 12.448 ;
  LAYER M1 ;
        RECT 30.144 12.396 30.176 12.468 ;
  LAYER M2 ;
        RECT 30.124 12.416 30.196 12.448 ;
  LAYER M1 ;
        RECT 27.584 9.456 27.616 9.528 ;
  LAYER M2 ;
        RECT 27.564 9.476 27.636 9.508 ;
  LAYER M2 ;
        RECT 27.6 9.476 30.16 9.508 ;
  LAYER M1 ;
        RECT 30.144 9.456 30.176 9.528 ;
  LAYER M2 ;
        RECT 30.124 9.476 30.196 9.508 ;
  LAYER M1 ;
        RECT 27.584 6.516 27.616 6.588 ;
  LAYER M2 ;
        RECT 27.564 6.536 27.636 6.568 ;
  LAYER M2 ;
        RECT 27.6 6.536 30.16 6.568 ;
  LAYER M1 ;
        RECT 30.144 6.516 30.176 6.588 ;
  LAYER M2 ;
        RECT 30.124 6.536 30.196 6.568 ;
  LAYER M1 ;
        RECT 30.144 5.676 30.176 5.748 ;
  LAYER M2 ;
        RECT 30.124 5.696 30.196 5.728 ;
  LAYER M1 ;
        RECT 30.144 5.712 30.176 6.216 ;
  LAYER M1 ;
        RECT 30.144 6.216 30.176 15.372 ;
  LAYER M1 ;
        RECT 16.064 15.336 16.096 15.408 ;
  LAYER M2 ;
        RECT 16.044 15.356 16.116 15.388 ;
  LAYER M1 ;
        RECT 16.064 15.204 16.096 15.372 ;
  LAYER M1 ;
        RECT 16.064 15.168 16.096 15.24 ;
  LAYER M2 ;
        RECT 16.044 15.188 16.116 15.22 ;
  LAYER M2 ;
        RECT 15.76 15.188 16.08 15.22 ;
  LAYER M1 ;
        RECT 15.744 15.168 15.776 15.24 ;
  LAYER M2 ;
        RECT 15.724 15.188 15.796 15.22 ;
  LAYER M1 ;
        RECT 16.064 12.396 16.096 12.468 ;
  LAYER M2 ;
        RECT 16.044 12.416 16.116 12.448 ;
  LAYER M1 ;
        RECT 16.064 12.264 16.096 12.432 ;
  LAYER M1 ;
        RECT 16.064 12.228 16.096 12.3 ;
  LAYER M2 ;
        RECT 16.044 12.248 16.116 12.28 ;
  LAYER M2 ;
        RECT 15.76 12.248 16.08 12.28 ;
  LAYER M1 ;
        RECT 15.744 12.228 15.776 12.3 ;
  LAYER M2 ;
        RECT 15.724 12.248 15.796 12.28 ;
  LAYER M1 ;
        RECT 16.064 9.456 16.096 9.528 ;
  LAYER M2 ;
        RECT 16.044 9.476 16.116 9.508 ;
  LAYER M1 ;
        RECT 16.064 9.324 16.096 9.492 ;
  LAYER M1 ;
        RECT 16.064 9.288 16.096 9.36 ;
  LAYER M2 ;
        RECT 16.044 9.308 16.116 9.34 ;
  LAYER M2 ;
        RECT 15.76 9.308 16.08 9.34 ;
  LAYER M1 ;
        RECT 15.744 9.288 15.776 9.36 ;
  LAYER M2 ;
        RECT 15.724 9.308 15.796 9.34 ;
  LAYER M1 ;
        RECT 16.064 6.516 16.096 6.588 ;
  LAYER M2 ;
        RECT 16.044 6.536 16.116 6.568 ;
  LAYER M1 ;
        RECT 16.064 6.384 16.096 6.552 ;
  LAYER M1 ;
        RECT 16.064 6.348 16.096 6.42 ;
  LAYER M2 ;
        RECT 16.044 6.368 16.116 6.4 ;
  LAYER M2 ;
        RECT 15.76 6.368 16.08 6.4 ;
  LAYER M1 ;
        RECT 15.744 6.348 15.776 6.42 ;
  LAYER M2 ;
        RECT 15.724 6.368 15.796 6.4 ;
  LAYER M1 ;
        RECT 15.744 5.676 15.776 5.748 ;
  LAYER M2 ;
        RECT 15.724 5.696 15.796 5.728 ;
  LAYER M1 ;
        RECT 15.744 5.712 15.776 6.216 ;
  LAYER M1 ;
        RECT 15.744 6.216 15.776 15.204 ;
  LAYER M2 ;
        RECT 15.76 5.696 30.16 5.728 ;
  LAYER M1 ;
        RECT 24.704 15.336 24.736 15.408 ;
  LAYER M2 ;
        RECT 24.684 15.356 24.756 15.388 ;
  LAYER M2 ;
        RECT 24.72 15.356 27.6 15.388 ;
  LAYER M1 ;
        RECT 27.584 15.336 27.616 15.408 ;
  LAYER M2 ;
        RECT 27.564 15.356 27.636 15.388 ;
  LAYER M1 ;
        RECT 24.704 6.516 24.736 6.588 ;
  LAYER M2 ;
        RECT 24.684 6.536 24.756 6.568 ;
  LAYER M2 ;
        RECT 24.72 6.536 27.6 6.568 ;
  LAYER M1 ;
        RECT 27.584 6.516 27.616 6.588 ;
  LAYER M2 ;
        RECT 27.564 6.536 27.636 6.568 ;
  LAYER M1 ;
        RECT 21.824 6.516 21.856 6.588 ;
  LAYER M2 ;
        RECT 21.804 6.536 21.876 6.568 ;
  LAYER M2 ;
        RECT 21.84 6.536 24.72 6.568 ;
  LAYER M1 ;
        RECT 24.704 6.516 24.736 6.588 ;
  LAYER M2 ;
        RECT 24.684 6.536 24.756 6.568 ;
  LAYER M1 ;
        RECT 18.944 6.516 18.976 6.588 ;
  LAYER M2 ;
        RECT 18.924 6.536 18.996 6.568 ;
  LAYER M2 ;
        RECT 18.96 6.536 21.84 6.568 ;
  LAYER M1 ;
        RECT 21.824 6.516 21.856 6.588 ;
  LAYER M2 ;
        RECT 21.804 6.536 21.876 6.568 ;
  LAYER M1 ;
        RECT 18.944 15.336 18.976 15.408 ;
  LAYER M2 ;
        RECT 18.924 15.356 18.996 15.388 ;
  LAYER M2 ;
        RECT 16.08 15.356 18.96 15.388 ;
  LAYER M1 ;
        RECT 16.064 15.336 16.096 15.408 ;
  LAYER M2 ;
        RECT 16.044 15.356 16.116 15.388 ;
  LAYER M1 ;
        RECT 21.824 15.336 21.856 15.408 ;
  LAYER M2 ;
        RECT 21.804 15.356 21.876 15.388 ;
  LAYER M2 ;
        RECT 18.96 15.356 21.84 15.388 ;
  LAYER M1 ;
        RECT 18.944 15.336 18.976 15.408 ;
  LAYER M2 ;
        RECT 18.924 15.356 18.996 15.388 ;
  LAYER M1 ;
        RECT 29.984 15.336 30.016 17.844 ;
  LAYER M1 ;
        RECT 29.92 15.336 29.952 17.844 ;
  LAYER M1 ;
        RECT 29.856 15.336 29.888 17.844 ;
  LAYER M1 ;
        RECT 29.792 15.336 29.824 17.844 ;
  LAYER M1 ;
        RECT 29.728 15.336 29.76 17.844 ;
  LAYER M1 ;
        RECT 29.664 15.336 29.696 17.844 ;
  LAYER M1 ;
        RECT 29.6 15.336 29.632 17.844 ;
  LAYER M1 ;
        RECT 29.536 15.336 29.568 17.844 ;
  LAYER M1 ;
        RECT 29.472 15.336 29.504 17.844 ;
  LAYER M1 ;
        RECT 29.408 15.336 29.44 17.844 ;
  LAYER M1 ;
        RECT 29.344 15.336 29.376 17.844 ;
  LAYER M1 ;
        RECT 29.28 15.336 29.312 17.844 ;
  LAYER M1 ;
        RECT 29.216 15.336 29.248 17.844 ;
  LAYER M1 ;
        RECT 29.152 15.336 29.184 17.844 ;
  LAYER M1 ;
        RECT 29.088 15.336 29.12 17.844 ;
  LAYER M1 ;
        RECT 29.024 15.336 29.056 17.844 ;
  LAYER M1 ;
        RECT 28.96 15.336 28.992 17.844 ;
  LAYER M1 ;
        RECT 28.896 15.336 28.928 17.844 ;
  LAYER M1 ;
        RECT 28.832 15.336 28.864 17.844 ;
  LAYER M1 ;
        RECT 28.768 15.336 28.8 17.844 ;
  LAYER M1 ;
        RECT 28.704 15.336 28.736 17.844 ;
  LAYER M1 ;
        RECT 28.64 15.336 28.672 17.844 ;
  LAYER M1 ;
        RECT 28.576 15.336 28.608 17.844 ;
  LAYER M1 ;
        RECT 28.512 15.336 28.544 17.844 ;
  LAYER M1 ;
        RECT 28.448 15.336 28.48 17.844 ;
  LAYER M1 ;
        RECT 28.384 15.336 28.416 17.844 ;
  LAYER M1 ;
        RECT 28.32 15.336 28.352 17.844 ;
  LAYER M1 ;
        RECT 28.256 15.336 28.288 17.844 ;
  LAYER M1 ;
        RECT 28.192 15.336 28.224 17.844 ;
  LAYER M1 ;
        RECT 28.128 15.336 28.16 17.844 ;
  LAYER M1 ;
        RECT 28.064 15.336 28.096 17.844 ;
  LAYER M1 ;
        RECT 28 15.336 28.032 17.844 ;
  LAYER M1 ;
        RECT 27.936 15.336 27.968 17.844 ;
  LAYER M1 ;
        RECT 27.872 15.336 27.904 17.844 ;
  LAYER M1 ;
        RECT 27.808 15.336 27.84 17.844 ;
  LAYER M1 ;
        RECT 27.744 15.336 27.776 17.844 ;
  LAYER M1 ;
        RECT 27.68 15.336 27.712 17.844 ;
  LAYER M2 ;
        RECT 27.564 17.728 30.036 17.76 ;
  LAYER M2 ;
        RECT 27.564 17.664 30.036 17.696 ;
  LAYER M2 ;
        RECT 27.564 17.6 30.036 17.632 ;
  LAYER M2 ;
        RECT 27.564 17.536 30.036 17.568 ;
  LAYER M2 ;
        RECT 27.564 17.472 30.036 17.504 ;
  LAYER M2 ;
        RECT 27.564 17.408 30.036 17.44 ;
  LAYER M2 ;
        RECT 27.564 17.344 30.036 17.376 ;
  LAYER M2 ;
        RECT 27.564 17.28 30.036 17.312 ;
  LAYER M2 ;
        RECT 27.564 17.216 30.036 17.248 ;
  LAYER M2 ;
        RECT 27.564 17.152 30.036 17.184 ;
  LAYER M2 ;
        RECT 27.564 17.088 30.036 17.12 ;
  LAYER M2 ;
        RECT 27.564 17.024 30.036 17.056 ;
  LAYER M2 ;
        RECT 27.564 16.96 30.036 16.992 ;
  LAYER M2 ;
        RECT 27.564 16.896 30.036 16.928 ;
  LAYER M2 ;
        RECT 27.564 16.832 30.036 16.864 ;
  LAYER M2 ;
        RECT 27.564 16.768 30.036 16.8 ;
  LAYER M2 ;
        RECT 27.564 16.704 30.036 16.736 ;
  LAYER M2 ;
        RECT 27.564 16.64 30.036 16.672 ;
  LAYER M2 ;
        RECT 27.564 16.576 30.036 16.608 ;
  LAYER M2 ;
        RECT 27.564 16.512 30.036 16.544 ;
  LAYER M2 ;
        RECT 27.564 16.448 30.036 16.48 ;
  LAYER M2 ;
        RECT 27.564 16.384 30.036 16.416 ;
  LAYER M2 ;
        RECT 27.564 16.32 30.036 16.352 ;
  LAYER M2 ;
        RECT 27.564 16.256 30.036 16.288 ;
  LAYER M2 ;
        RECT 27.564 16.192 30.036 16.224 ;
  LAYER M2 ;
        RECT 27.564 16.128 30.036 16.16 ;
  LAYER M2 ;
        RECT 27.564 16.064 30.036 16.096 ;
  LAYER M2 ;
        RECT 27.564 16 30.036 16.032 ;
  LAYER M2 ;
        RECT 27.564 15.936 30.036 15.968 ;
  LAYER M2 ;
        RECT 27.564 15.872 30.036 15.904 ;
  LAYER M2 ;
        RECT 27.564 15.808 30.036 15.84 ;
  LAYER M2 ;
        RECT 27.564 15.744 30.036 15.776 ;
  LAYER M2 ;
        RECT 27.564 15.68 30.036 15.712 ;
  LAYER M2 ;
        RECT 27.564 15.616 30.036 15.648 ;
  LAYER M2 ;
        RECT 27.564 15.552 30.036 15.584 ;
  LAYER M2 ;
        RECT 27.564 15.488 30.036 15.52 ;
  LAYER M3 ;
        RECT 29.984 15.336 30.016 17.844 ;
  LAYER M3 ;
        RECT 29.92 15.336 29.952 17.844 ;
  LAYER M3 ;
        RECT 29.856 15.336 29.888 17.844 ;
  LAYER M3 ;
        RECT 29.792 15.336 29.824 17.844 ;
  LAYER M3 ;
        RECT 29.728 15.336 29.76 17.844 ;
  LAYER M3 ;
        RECT 29.664 15.336 29.696 17.844 ;
  LAYER M3 ;
        RECT 29.6 15.336 29.632 17.844 ;
  LAYER M3 ;
        RECT 29.536 15.336 29.568 17.844 ;
  LAYER M3 ;
        RECT 29.472 15.336 29.504 17.844 ;
  LAYER M3 ;
        RECT 29.408 15.336 29.44 17.844 ;
  LAYER M3 ;
        RECT 29.344 15.336 29.376 17.844 ;
  LAYER M3 ;
        RECT 29.28 15.336 29.312 17.844 ;
  LAYER M3 ;
        RECT 29.216 15.336 29.248 17.844 ;
  LAYER M3 ;
        RECT 29.152 15.336 29.184 17.844 ;
  LAYER M3 ;
        RECT 29.088 15.336 29.12 17.844 ;
  LAYER M3 ;
        RECT 29.024 15.336 29.056 17.844 ;
  LAYER M3 ;
        RECT 28.96 15.336 28.992 17.844 ;
  LAYER M3 ;
        RECT 28.896 15.336 28.928 17.844 ;
  LAYER M3 ;
        RECT 28.832 15.336 28.864 17.844 ;
  LAYER M3 ;
        RECT 28.768 15.336 28.8 17.844 ;
  LAYER M3 ;
        RECT 28.704 15.336 28.736 17.844 ;
  LAYER M3 ;
        RECT 28.64 15.336 28.672 17.844 ;
  LAYER M3 ;
        RECT 28.576 15.336 28.608 17.844 ;
  LAYER M3 ;
        RECT 28.512 15.336 28.544 17.844 ;
  LAYER M3 ;
        RECT 28.448 15.336 28.48 17.844 ;
  LAYER M3 ;
        RECT 28.384 15.336 28.416 17.844 ;
  LAYER M3 ;
        RECT 28.32 15.336 28.352 17.844 ;
  LAYER M3 ;
        RECT 28.256 15.336 28.288 17.844 ;
  LAYER M3 ;
        RECT 28.192 15.336 28.224 17.844 ;
  LAYER M3 ;
        RECT 28.128 15.336 28.16 17.844 ;
  LAYER M3 ;
        RECT 28.064 15.336 28.096 17.844 ;
  LAYER M3 ;
        RECT 28 15.336 28.032 17.844 ;
  LAYER M3 ;
        RECT 27.936 15.336 27.968 17.844 ;
  LAYER M3 ;
        RECT 27.872 15.336 27.904 17.844 ;
  LAYER M3 ;
        RECT 27.808 15.336 27.84 17.844 ;
  LAYER M3 ;
        RECT 27.744 15.336 27.776 17.844 ;
  LAYER M3 ;
        RECT 27.68 15.336 27.712 17.844 ;
  LAYER M3 ;
        RECT 27.584 15.336 27.616 17.844 ;
  LAYER M1 ;
        RECT 29.999 15.372 30.001 17.808 ;
  LAYER M1 ;
        RECT 29.919 15.372 29.921 17.808 ;
  LAYER M1 ;
        RECT 29.839 15.372 29.841 17.808 ;
  LAYER M1 ;
        RECT 29.759 15.372 29.761 17.808 ;
  LAYER M1 ;
        RECT 29.679 15.372 29.681 17.808 ;
  LAYER M1 ;
        RECT 29.599 15.372 29.601 17.808 ;
  LAYER M1 ;
        RECT 29.519 15.372 29.521 17.808 ;
  LAYER M1 ;
        RECT 29.439 15.372 29.441 17.808 ;
  LAYER M1 ;
        RECT 29.359 15.372 29.361 17.808 ;
  LAYER M1 ;
        RECT 29.279 15.372 29.281 17.808 ;
  LAYER M1 ;
        RECT 29.199 15.372 29.201 17.808 ;
  LAYER M1 ;
        RECT 29.119 15.372 29.121 17.808 ;
  LAYER M1 ;
        RECT 29.039 15.372 29.041 17.808 ;
  LAYER M1 ;
        RECT 28.959 15.372 28.961 17.808 ;
  LAYER M1 ;
        RECT 28.879 15.372 28.881 17.808 ;
  LAYER M1 ;
        RECT 28.799 15.372 28.801 17.808 ;
  LAYER M1 ;
        RECT 28.719 15.372 28.721 17.808 ;
  LAYER M1 ;
        RECT 28.639 15.372 28.641 17.808 ;
  LAYER M1 ;
        RECT 28.559 15.372 28.561 17.808 ;
  LAYER M1 ;
        RECT 28.479 15.372 28.481 17.808 ;
  LAYER M1 ;
        RECT 28.399 15.372 28.401 17.808 ;
  LAYER M1 ;
        RECT 28.319 15.372 28.321 17.808 ;
  LAYER M1 ;
        RECT 28.239 15.372 28.241 17.808 ;
  LAYER M1 ;
        RECT 28.159 15.372 28.161 17.808 ;
  LAYER M1 ;
        RECT 28.079 15.372 28.081 17.808 ;
  LAYER M1 ;
        RECT 27.999 15.372 28.001 17.808 ;
  LAYER M1 ;
        RECT 27.919 15.372 27.921 17.808 ;
  LAYER M1 ;
        RECT 27.839 15.372 27.841 17.808 ;
  LAYER M1 ;
        RECT 27.759 15.372 27.761 17.808 ;
  LAYER M1 ;
        RECT 27.679 15.372 27.681 17.808 ;
  LAYER M2 ;
        RECT 27.6 17.807 30 17.809 ;
  LAYER M2 ;
        RECT 27.6 17.723 30 17.725 ;
  LAYER M2 ;
        RECT 27.6 17.639 30 17.641 ;
  LAYER M2 ;
        RECT 27.6 17.555 30 17.557 ;
  LAYER M2 ;
        RECT 27.6 17.471 30 17.473 ;
  LAYER M2 ;
        RECT 27.6 17.387 30 17.389 ;
  LAYER M2 ;
        RECT 27.6 17.303 30 17.305 ;
  LAYER M2 ;
        RECT 27.6 17.219 30 17.221 ;
  LAYER M2 ;
        RECT 27.6 17.135 30 17.137 ;
  LAYER M2 ;
        RECT 27.6 17.051 30 17.053 ;
  LAYER M2 ;
        RECT 27.6 16.967 30 16.969 ;
  LAYER M2 ;
        RECT 27.6 16.883 30 16.885 ;
  LAYER M2 ;
        RECT 27.6 16.7995 30 16.8015 ;
  LAYER M2 ;
        RECT 27.6 16.715 30 16.717 ;
  LAYER M2 ;
        RECT 27.6 16.631 30 16.633 ;
  LAYER M2 ;
        RECT 27.6 16.547 30 16.549 ;
  LAYER M2 ;
        RECT 27.6 16.463 30 16.465 ;
  LAYER M2 ;
        RECT 27.6 16.379 30 16.381 ;
  LAYER M2 ;
        RECT 27.6 16.295 30 16.297 ;
  LAYER M2 ;
        RECT 27.6 16.211 30 16.213 ;
  LAYER M2 ;
        RECT 27.6 16.127 30 16.129 ;
  LAYER M2 ;
        RECT 27.6 16.043 30 16.045 ;
  LAYER M2 ;
        RECT 27.6 15.959 30 15.961 ;
  LAYER M2 ;
        RECT 27.6 15.875 30 15.877 ;
  LAYER M2 ;
        RECT 27.6 15.791 30 15.793 ;
  LAYER M2 ;
        RECT 27.6 15.707 30 15.709 ;
  LAYER M2 ;
        RECT 27.6 15.623 30 15.625 ;
  LAYER M2 ;
        RECT 27.6 15.539 30 15.541 ;
  LAYER M2 ;
        RECT 27.6 15.455 30 15.457 ;
  LAYER M1 ;
        RECT 29.984 12.396 30.016 14.904 ;
  LAYER M1 ;
        RECT 29.92 12.396 29.952 14.904 ;
  LAYER M1 ;
        RECT 29.856 12.396 29.888 14.904 ;
  LAYER M1 ;
        RECT 29.792 12.396 29.824 14.904 ;
  LAYER M1 ;
        RECT 29.728 12.396 29.76 14.904 ;
  LAYER M1 ;
        RECT 29.664 12.396 29.696 14.904 ;
  LAYER M1 ;
        RECT 29.6 12.396 29.632 14.904 ;
  LAYER M1 ;
        RECT 29.536 12.396 29.568 14.904 ;
  LAYER M1 ;
        RECT 29.472 12.396 29.504 14.904 ;
  LAYER M1 ;
        RECT 29.408 12.396 29.44 14.904 ;
  LAYER M1 ;
        RECT 29.344 12.396 29.376 14.904 ;
  LAYER M1 ;
        RECT 29.28 12.396 29.312 14.904 ;
  LAYER M1 ;
        RECT 29.216 12.396 29.248 14.904 ;
  LAYER M1 ;
        RECT 29.152 12.396 29.184 14.904 ;
  LAYER M1 ;
        RECT 29.088 12.396 29.12 14.904 ;
  LAYER M1 ;
        RECT 29.024 12.396 29.056 14.904 ;
  LAYER M1 ;
        RECT 28.96 12.396 28.992 14.904 ;
  LAYER M1 ;
        RECT 28.896 12.396 28.928 14.904 ;
  LAYER M1 ;
        RECT 28.832 12.396 28.864 14.904 ;
  LAYER M1 ;
        RECT 28.768 12.396 28.8 14.904 ;
  LAYER M1 ;
        RECT 28.704 12.396 28.736 14.904 ;
  LAYER M1 ;
        RECT 28.64 12.396 28.672 14.904 ;
  LAYER M1 ;
        RECT 28.576 12.396 28.608 14.904 ;
  LAYER M1 ;
        RECT 28.512 12.396 28.544 14.904 ;
  LAYER M1 ;
        RECT 28.448 12.396 28.48 14.904 ;
  LAYER M1 ;
        RECT 28.384 12.396 28.416 14.904 ;
  LAYER M1 ;
        RECT 28.32 12.396 28.352 14.904 ;
  LAYER M1 ;
        RECT 28.256 12.396 28.288 14.904 ;
  LAYER M1 ;
        RECT 28.192 12.396 28.224 14.904 ;
  LAYER M1 ;
        RECT 28.128 12.396 28.16 14.904 ;
  LAYER M1 ;
        RECT 28.064 12.396 28.096 14.904 ;
  LAYER M1 ;
        RECT 28 12.396 28.032 14.904 ;
  LAYER M1 ;
        RECT 27.936 12.396 27.968 14.904 ;
  LAYER M1 ;
        RECT 27.872 12.396 27.904 14.904 ;
  LAYER M1 ;
        RECT 27.808 12.396 27.84 14.904 ;
  LAYER M1 ;
        RECT 27.744 12.396 27.776 14.904 ;
  LAYER M1 ;
        RECT 27.68 12.396 27.712 14.904 ;
  LAYER M2 ;
        RECT 27.564 14.788 30.036 14.82 ;
  LAYER M2 ;
        RECT 27.564 14.724 30.036 14.756 ;
  LAYER M2 ;
        RECT 27.564 14.66 30.036 14.692 ;
  LAYER M2 ;
        RECT 27.564 14.596 30.036 14.628 ;
  LAYER M2 ;
        RECT 27.564 14.532 30.036 14.564 ;
  LAYER M2 ;
        RECT 27.564 14.468 30.036 14.5 ;
  LAYER M2 ;
        RECT 27.564 14.404 30.036 14.436 ;
  LAYER M2 ;
        RECT 27.564 14.34 30.036 14.372 ;
  LAYER M2 ;
        RECT 27.564 14.276 30.036 14.308 ;
  LAYER M2 ;
        RECT 27.564 14.212 30.036 14.244 ;
  LAYER M2 ;
        RECT 27.564 14.148 30.036 14.18 ;
  LAYER M2 ;
        RECT 27.564 14.084 30.036 14.116 ;
  LAYER M2 ;
        RECT 27.564 14.02 30.036 14.052 ;
  LAYER M2 ;
        RECT 27.564 13.956 30.036 13.988 ;
  LAYER M2 ;
        RECT 27.564 13.892 30.036 13.924 ;
  LAYER M2 ;
        RECT 27.564 13.828 30.036 13.86 ;
  LAYER M2 ;
        RECT 27.564 13.764 30.036 13.796 ;
  LAYER M2 ;
        RECT 27.564 13.7 30.036 13.732 ;
  LAYER M2 ;
        RECT 27.564 13.636 30.036 13.668 ;
  LAYER M2 ;
        RECT 27.564 13.572 30.036 13.604 ;
  LAYER M2 ;
        RECT 27.564 13.508 30.036 13.54 ;
  LAYER M2 ;
        RECT 27.564 13.444 30.036 13.476 ;
  LAYER M2 ;
        RECT 27.564 13.38 30.036 13.412 ;
  LAYER M2 ;
        RECT 27.564 13.316 30.036 13.348 ;
  LAYER M2 ;
        RECT 27.564 13.252 30.036 13.284 ;
  LAYER M2 ;
        RECT 27.564 13.188 30.036 13.22 ;
  LAYER M2 ;
        RECT 27.564 13.124 30.036 13.156 ;
  LAYER M2 ;
        RECT 27.564 13.06 30.036 13.092 ;
  LAYER M2 ;
        RECT 27.564 12.996 30.036 13.028 ;
  LAYER M2 ;
        RECT 27.564 12.932 30.036 12.964 ;
  LAYER M2 ;
        RECT 27.564 12.868 30.036 12.9 ;
  LAYER M2 ;
        RECT 27.564 12.804 30.036 12.836 ;
  LAYER M2 ;
        RECT 27.564 12.74 30.036 12.772 ;
  LAYER M2 ;
        RECT 27.564 12.676 30.036 12.708 ;
  LAYER M2 ;
        RECT 27.564 12.612 30.036 12.644 ;
  LAYER M2 ;
        RECT 27.564 12.548 30.036 12.58 ;
  LAYER M3 ;
        RECT 29.984 12.396 30.016 14.904 ;
  LAYER M3 ;
        RECT 29.92 12.396 29.952 14.904 ;
  LAYER M3 ;
        RECT 29.856 12.396 29.888 14.904 ;
  LAYER M3 ;
        RECT 29.792 12.396 29.824 14.904 ;
  LAYER M3 ;
        RECT 29.728 12.396 29.76 14.904 ;
  LAYER M3 ;
        RECT 29.664 12.396 29.696 14.904 ;
  LAYER M3 ;
        RECT 29.6 12.396 29.632 14.904 ;
  LAYER M3 ;
        RECT 29.536 12.396 29.568 14.904 ;
  LAYER M3 ;
        RECT 29.472 12.396 29.504 14.904 ;
  LAYER M3 ;
        RECT 29.408 12.396 29.44 14.904 ;
  LAYER M3 ;
        RECT 29.344 12.396 29.376 14.904 ;
  LAYER M3 ;
        RECT 29.28 12.396 29.312 14.904 ;
  LAYER M3 ;
        RECT 29.216 12.396 29.248 14.904 ;
  LAYER M3 ;
        RECT 29.152 12.396 29.184 14.904 ;
  LAYER M3 ;
        RECT 29.088 12.396 29.12 14.904 ;
  LAYER M3 ;
        RECT 29.024 12.396 29.056 14.904 ;
  LAYER M3 ;
        RECT 28.96 12.396 28.992 14.904 ;
  LAYER M3 ;
        RECT 28.896 12.396 28.928 14.904 ;
  LAYER M3 ;
        RECT 28.832 12.396 28.864 14.904 ;
  LAYER M3 ;
        RECT 28.768 12.396 28.8 14.904 ;
  LAYER M3 ;
        RECT 28.704 12.396 28.736 14.904 ;
  LAYER M3 ;
        RECT 28.64 12.396 28.672 14.904 ;
  LAYER M3 ;
        RECT 28.576 12.396 28.608 14.904 ;
  LAYER M3 ;
        RECT 28.512 12.396 28.544 14.904 ;
  LAYER M3 ;
        RECT 28.448 12.396 28.48 14.904 ;
  LAYER M3 ;
        RECT 28.384 12.396 28.416 14.904 ;
  LAYER M3 ;
        RECT 28.32 12.396 28.352 14.904 ;
  LAYER M3 ;
        RECT 28.256 12.396 28.288 14.904 ;
  LAYER M3 ;
        RECT 28.192 12.396 28.224 14.904 ;
  LAYER M3 ;
        RECT 28.128 12.396 28.16 14.904 ;
  LAYER M3 ;
        RECT 28.064 12.396 28.096 14.904 ;
  LAYER M3 ;
        RECT 28 12.396 28.032 14.904 ;
  LAYER M3 ;
        RECT 27.936 12.396 27.968 14.904 ;
  LAYER M3 ;
        RECT 27.872 12.396 27.904 14.904 ;
  LAYER M3 ;
        RECT 27.808 12.396 27.84 14.904 ;
  LAYER M3 ;
        RECT 27.744 12.396 27.776 14.904 ;
  LAYER M3 ;
        RECT 27.68 12.396 27.712 14.904 ;
  LAYER M3 ;
        RECT 27.584 12.396 27.616 14.904 ;
  LAYER M1 ;
        RECT 29.999 12.432 30.001 14.868 ;
  LAYER M1 ;
        RECT 29.919 12.432 29.921 14.868 ;
  LAYER M1 ;
        RECT 29.839 12.432 29.841 14.868 ;
  LAYER M1 ;
        RECT 29.759 12.432 29.761 14.868 ;
  LAYER M1 ;
        RECT 29.679 12.432 29.681 14.868 ;
  LAYER M1 ;
        RECT 29.599 12.432 29.601 14.868 ;
  LAYER M1 ;
        RECT 29.519 12.432 29.521 14.868 ;
  LAYER M1 ;
        RECT 29.439 12.432 29.441 14.868 ;
  LAYER M1 ;
        RECT 29.359 12.432 29.361 14.868 ;
  LAYER M1 ;
        RECT 29.279 12.432 29.281 14.868 ;
  LAYER M1 ;
        RECT 29.199 12.432 29.201 14.868 ;
  LAYER M1 ;
        RECT 29.119 12.432 29.121 14.868 ;
  LAYER M1 ;
        RECT 29.039 12.432 29.041 14.868 ;
  LAYER M1 ;
        RECT 28.959 12.432 28.961 14.868 ;
  LAYER M1 ;
        RECT 28.879 12.432 28.881 14.868 ;
  LAYER M1 ;
        RECT 28.799 12.432 28.801 14.868 ;
  LAYER M1 ;
        RECT 28.719 12.432 28.721 14.868 ;
  LAYER M1 ;
        RECT 28.639 12.432 28.641 14.868 ;
  LAYER M1 ;
        RECT 28.559 12.432 28.561 14.868 ;
  LAYER M1 ;
        RECT 28.479 12.432 28.481 14.868 ;
  LAYER M1 ;
        RECT 28.399 12.432 28.401 14.868 ;
  LAYER M1 ;
        RECT 28.319 12.432 28.321 14.868 ;
  LAYER M1 ;
        RECT 28.239 12.432 28.241 14.868 ;
  LAYER M1 ;
        RECT 28.159 12.432 28.161 14.868 ;
  LAYER M1 ;
        RECT 28.079 12.432 28.081 14.868 ;
  LAYER M1 ;
        RECT 27.999 12.432 28.001 14.868 ;
  LAYER M1 ;
        RECT 27.919 12.432 27.921 14.868 ;
  LAYER M1 ;
        RECT 27.839 12.432 27.841 14.868 ;
  LAYER M1 ;
        RECT 27.759 12.432 27.761 14.868 ;
  LAYER M1 ;
        RECT 27.679 12.432 27.681 14.868 ;
  LAYER M2 ;
        RECT 27.6 14.867 30 14.869 ;
  LAYER M2 ;
        RECT 27.6 14.783 30 14.785 ;
  LAYER M2 ;
        RECT 27.6 14.699 30 14.701 ;
  LAYER M2 ;
        RECT 27.6 14.615 30 14.617 ;
  LAYER M2 ;
        RECT 27.6 14.531 30 14.533 ;
  LAYER M2 ;
        RECT 27.6 14.447 30 14.449 ;
  LAYER M2 ;
        RECT 27.6 14.363 30 14.365 ;
  LAYER M2 ;
        RECT 27.6 14.279 30 14.281 ;
  LAYER M2 ;
        RECT 27.6 14.195 30 14.197 ;
  LAYER M2 ;
        RECT 27.6 14.111 30 14.113 ;
  LAYER M2 ;
        RECT 27.6 14.027 30 14.029 ;
  LAYER M2 ;
        RECT 27.6 13.943 30 13.945 ;
  LAYER M2 ;
        RECT 27.6 13.8595 30 13.8615 ;
  LAYER M2 ;
        RECT 27.6 13.775 30 13.777 ;
  LAYER M2 ;
        RECT 27.6 13.691 30 13.693 ;
  LAYER M2 ;
        RECT 27.6 13.607 30 13.609 ;
  LAYER M2 ;
        RECT 27.6 13.523 30 13.525 ;
  LAYER M2 ;
        RECT 27.6 13.439 30 13.441 ;
  LAYER M2 ;
        RECT 27.6 13.355 30 13.357 ;
  LAYER M2 ;
        RECT 27.6 13.271 30 13.273 ;
  LAYER M2 ;
        RECT 27.6 13.187 30 13.189 ;
  LAYER M2 ;
        RECT 27.6 13.103 30 13.105 ;
  LAYER M2 ;
        RECT 27.6 13.019 30 13.021 ;
  LAYER M2 ;
        RECT 27.6 12.935 30 12.937 ;
  LAYER M2 ;
        RECT 27.6 12.851 30 12.853 ;
  LAYER M2 ;
        RECT 27.6 12.767 30 12.769 ;
  LAYER M2 ;
        RECT 27.6 12.683 30 12.685 ;
  LAYER M2 ;
        RECT 27.6 12.599 30 12.601 ;
  LAYER M2 ;
        RECT 27.6 12.515 30 12.517 ;
  LAYER M1 ;
        RECT 29.984 9.456 30.016 11.964 ;
  LAYER M1 ;
        RECT 29.92 9.456 29.952 11.964 ;
  LAYER M1 ;
        RECT 29.856 9.456 29.888 11.964 ;
  LAYER M1 ;
        RECT 29.792 9.456 29.824 11.964 ;
  LAYER M1 ;
        RECT 29.728 9.456 29.76 11.964 ;
  LAYER M1 ;
        RECT 29.664 9.456 29.696 11.964 ;
  LAYER M1 ;
        RECT 29.6 9.456 29.632 11.964 ;
  LAYER M1 ;
        RECT 29.536 9.456 29.568 11.964 ;
  LAYER M1 ;
        RECT 29.472 9.456 29.504 11.964 ;
  LAYER M1 ;
        RECT 29.408 9.456 29.44 11.964 ;
  LAYER M1 ;
        RECT 29.344 9.456 29.376 11.964 ;
  LAYER M1 ;
        RECT 29.28 9.456 29.312 11.964 ;
  LAYER M1 ;
        RECT 29.216 9.456 29.248 11.964 ;
  LAYER M1 ;
        RECT 29.152 9.456 29.184 11.964 ;
  LAYER M1 ;
        RECT 29.088 9.456 29.12 11.964 ;
  LAYER M1 ;
        RECT 29.024 9.456 29.056 11.964 ;
  LAYER M1 ;
        RECT 28.96 9.456 28.992 11.964 ;
  LAYER M1 ;
        RECT 28.896 9.456 28.928 11.964 ;
  LAYER M1 ;
        RECT 28.832 9.456 28.864 11.964 ;
  LAYER M1 ;
        RECT 28.768 9.456 28.8 11.964 ;
  LAYER M1 ;
        RECT 28.704 9.456 28.736 11.964 ;
  LAYER M1 ;
        RECT 28.64 9.456 28.672 11.964 ;
  LAYER M1 ;
        RECT 28.576 9.456 28.608 11.964 ;
  LAYER M1 ;
        RECT 28.512 9.456 28.544 11.964 ;
  LAYER M1 ;
        RECT 28.448 9.456 28.48 11.964 ;
  LAYER M1 ;
        RECT 28.384 9.456 28.416 11.964 ;
  LAYER M1 ;
        RECT 28.32 9.456 28.352 11.964 ;
  LAYER M1 ;
        RECT 28.256 9.456 28.288 11.964 ;
  LAYER M1 ;
        RECT 28.192 9.456 28.224 11.964 ;
  LAYER M1 ;
        RECT 28.128 9.456 28.16 11.964 ;
  LAYER M1 ;
        RECT 28.064 9.456 28.096 11.964 ;
  LAYER M1 ;
        RECT 28 9.456 28.032 11.964 ;
  LAYER M1 ;
        RECT 27.936 9.456 27.968 11.964 ;
  LAYER M1 ;
        RECT 27.872 9.456 27.904 11.964 ;
  LAYER M1 ;
        RECT 27.808 9.456 27.84 11.964 ;
  LAYER M1 ;
        RECT 27.744 9.456 27.776 11.964 ;
  LAYER M1 ;
        RECT 27.68 9.456 27.712 11.964 ;
  LAYER M2 ;
        RECT 27.564 11.848 30.036 11.88 ;
  LAYER M2 ;
        RECT 27.564 11.784 30.036 11.816 ;
  LAYER M2 ;
        RECT 27.564 11.72 30.036 11.752 ;
  LAYER M2 ;
        RECT 27.564 11.656 30.036 11.688 ;
  LAYER M2 ;
        RECT 27.564 11.592 30.036 11.624 ;
  LAYER M2 ;
        RECT 27.564 11.528 30.036 11.56 ;
  LAYER M2 ;
        RECT 27.564 11.464 30.036 11.496 ;
  LAYER M2 ;
        RECT 27.564 11.4 30.036 11.432 ;
  LAYER M2 ;
        RECT 27.564 11.336 30.036 11.368 ;
  LAYER M2 ;
        RECT 27.564 11.272 30.036 11.304 ;
  LAYER M2 ;
        RECT 27.564 11.208 30.036 11.24 ;
  LAYER M2 ;
        RECT 27.564 11.144 30.036 11.176 ;
  LAYER M2 ;
        RECT 27.564 11.08 30.036 11.112 ;
  LAYER M2 ;
        RECT 27.564 11.016 30.036 11.048 ;
  LAYER M2 ;
        RECT 27.564 10.952 30.036 10.984 ;
  LAYER M2 ;
        RECT 27.564 10.888 30.036 10.92 ;
  LAYER M2 ;
        RECT 27.564 10.824 30.036 10.856 ;
  LAYER M2 ;
        RECT 27.564 10.76 30.036 10.792 ;
  LAYER M2 ;
        RECT 27.564 10.696 30.036 10.728 ;
  LAYER M2 ;
        RECT 27.564 10.632 30.036 10.664 ;
  LAYER M2 ;
        RECT 27.564 10.568 30.036 10.6 ;
  LAYER M2 ;
        RECT 27.564 10.504 30.036 10.536 ;
  LAYER M2 ;
        RECT 27.564 10.44 30.036 10.472 ;
  LAYER M2 ;
        RECT 27.564 10.376 30.036 10.408 ;
  LAYER M2 ;
        RECT 27.564 10.312 30.036 10.344 ;
  LAYER M2 ;
        RECT 27.564 10.248 30.036 10.28 ;
  LAYER M2 ;
        RECT 27.564 10.184 30.036 10.216 ;
  LAYER M2 ;
        RECT 27.564 10.12 30.036 10.152 ;
  LAYER M2 ;
        RECT 27.564 10.056 30.036 10.088 ;
  LAYER M2 ;
        RECT 27.564 9.992 30.036 10.024 ;
  LAYER M2 ;
        RECT 27.564 9.928 30.036 9.96 ;
  LAYER M2 ;
        RECT 27.564 9.864 30.036 9.896 ;
  LAYER M2 ;
        RECT 27.564 9.8 30.036 9.832 ;
  LAYER M2 ;
        RECT 27.564 9.736 30.036 9.768 ;
  LAYER M2 ;
        RECT 27.564 9.672 30.036 9.704 ;
  LAYER M2 ;
        RECT 27.564 9.608 30.036 9.64 ;
  LAYER M3 ;
        RECT 29.984 9.456 30.016 11.964 ;
  LAYER M3 ;
        RECT 29.92 9.456 29.952 11.964 ;
  LAYER M3 ;
        RECT 29.856 9.456 29.888 11.964 ;
  LAYER M3 ;
        RECT 29.792 9.456 29.824 11.964 ;
  LAYER M3 ;
        RECT 29.728 9.456 29.76 11.964 ;
  LAYER M3 ;
        RECT 29.664 9.456 29.696 11.964 ;
  LAYER M3 ;
        RECT 29.6 9.456 29.632 11.964 ;
  LAYER M3 ;
        RECT 29.536 9.456 29.568 11.964 ;
  LAYER M3 ;
        RECT 29.472 9.456 29.504 11.964 ;
  LAYER M3 ;
        RECT 29.408 9.456 29.44 11.964 ;
  LAYER M3 ;
        RECT 29.344 9.456 29.376 11.964 ;
  LAYER M3 ;
        RECT 29.28 9.456 29.312 11.964 ;
  LAYER M3 ;
        RECT 29.216 9.456 29.248 11.964 ;
  LAYER M3 ;
        RECT 29.152 9.456 29.184 11.964 ;
  LAYER M3 ;
        RECT 29.088 9.456 29.12 11.964 ;
  LAYER M3 ;
        RECT 29.024 9.456 29.056 11.964 ;
  LAYER M3 ;
        RECT 28.96 9.456 28.992 11.964 ;
  LAYER M3 ;
        RECT 28.896 9.456 28.928 11.964 ;
  LAYER M3 ;
        RECT 28.832 9.456 28.864 11.964 ;
  LAYER M3 ;
        RECT 28.768 9.456 28.8 11.964 ;
  LAYER M3 ;
        RECT 28.704 9.456 28.736 11.964 ;
  LAYER M3 ;
        RECT 28.64 9.456 28.672 11.964 ;
  LAYER M3 ;
        RECT 28.576 9.456 28.608 11.964 ;
  LAYER M3 ;
        RECT 28.512 9.456 28.544 11.964 ;
  LAYER M3 ;
        RECT 28.448 9.456 28.48 11.964 ;
  LAYER M3 ;
        RECT 28.384 9.456 28.416 11.964 ;
  LAYER M3 ;
        RECT 28.32 9.456 28.352 11.964 ;
  LAYER M3 ;
        RECT 28.256 9.456 28.288 11.964 ;
  LAYER M3 ;
        RECT 28.192 9.456 28.224 11.964 ;
  LAYER M3 ;
        RECT 28.128 9.456 28.16 11.964 ;
  LAYER M3 ;
        RECT 28.064 9.456 28.096 11.964 ;
  LAYER M3 ;
        RECT 28 9.456 28.032 11.964 ;
  LAYER M3 ;
        RECT 27.936 9.456 27.968 11.964 ;
  LAYER M3 ;
        RECT 27.872 9.456 27.904 11.964 ;
  LAYER M3 ;
        RECT 27.808 9.456 27.84 11.964 ;
  LAYER M3 ;
        RECT 27.744 9.456 27.776 11.964 ;
  LAYER M3 ;
        RECT 27.68 9.456 27.712 11.964 ;
  LAYER M3 ;
        RECT 27.584 9.456 27.616 11.964 ;
  LAYER M1 ;
        RECT 29.999 9.492 30.001 11.928 ;
  LAYER M1 ;
        RECT 29.919 9.492 29.921 11.928 ;
  LAYER M1 ;
        RECT 29.839 9.492 29.841 11.928 ;
  LAYER M1 ;
        RECT 29.759 9.492 29.761 11.928 ;
  LAYER M1 ;
        RECT 29.679 9.492 29.681 11.928 ;
  LAYER M1 ;
        RECT 29.599 9.492 29.601 11.928 ;
  LAYER M1 ;
        RECT 29.519 9.492 29.521 11.928 ;
  LAYER M1 ;
        RECT 29.439 9.492 29.441 11.928 ;
  LAYER M1 ;
        RECT 29.359 9.492 29.361 11.928 ;
  LAYER M1 ;
        RECT 29.279 9.492 29.281 11.928 ;
  LAYER M1 ;
        RECT 29.199 9.492 29.201 11.928 ;
  LAYER M1 ;
        RECT 29.119 9.492 29.121 11.928 ;
  LAYER M1 ;
        RECT 29.039 9.492 29.041 11.928 ;
  LAYER M1 ;
        RECT 28.959 9.492 28.961 11.928 ;
  LAYER M1 ;
        RECT 28.879 9.492 28.881 11.928 ;
  LAYER M1 ;
        RECT 28.799 9.492 28.801 11.928 ;
  LAYER M1 ;
        RECT 28.719 9.492 28.721 11.928 ;
  LAYER M1 ;
        RECT 28.639 9.492 28.641 11.928 ;
  LAYER M1 ;
        RECT 28.559 9.492 28.561 11.928 ;
  LAYER M1 ;
        RECT 28.479 9.492 28.481 11.928 ;
  LAYER M1 ;
        RECT 28.399 9.492 28.401 11.928 ;
  LAYER M1 ;
        RECT 28.319 9.492 28.321 11.928 ;
  LAYER M1 ;
        RECT 28.239 9.492 28.241 11.928 ;
  LAYER M1 ;
        RECT 28.159 9.492 28.161 11.928 ;
  LAYER M1 ;
        RECT 28.079 9.492 28.081 11.928 ;
  LAYER M1 ;
        RECT 27.999 9.492 28.001 11.928 ;
  LAYER M1 ;
        RECT 27.919 9.492 27.921 11.928 ;
  LAYER M1 ;
        RECT 27.839 9.492 27.841 11.928 ;
  LAYER M1 ;
        RECT 27.759 9.492 27.761 11.928 ;
  LAYER M1 ;
        RECT 27.679 9.492 27.681 11.928 ;
  LAYER M2 ;
        RECT 27.6 11.927 30 11.929 ;
  LAYER M2 ;
        RECT 27.6 11.843 30 11.845 ;
  LAYER M2 ;
        RECT 27.6 11.759 30 11.761 ;
  LAYER M2 ;
        RECT 27.6 11.675 30 11.677 ;
  LAYER M2 ;
        RECT 27.6 11.591 30 11.593 ;
  LAYER M2 ;
        RECT 27.6 11.507 30 11.509 ;
  LAYER M2 ;
        RECT 27.6 11.423 30 11.425 ;
  LAYER M2 ;
        RECT 27.6 11.339 30 11.341 ;
  LAYER M2 ;
        RECT 27.6 11.255 30 11.257 ;
  LAYER M2 ;
        RECT 27.6 11.171 30 11.173 ;
  LAYER M2 ;
        RECT 27.6 11.087 30 11.089 ;
  LAYER M2 ;
        RECT 27.6 11.003 30 11.005 ;
  LAYER M2 ;
        RECT 27.6 10.9195 30 10.9215 ;
  LAYER M2 ;
        RECT 27.6 10.835 30 10.837 ;
  LAYER M2 ;
        RECT 27.6 10.751 30 10.753 ;
  LAYER M2 ;
        RECT 27.6 10.667 30 10.669 ;
  LAYER M2 ;
        RECT 27.6 10.583 30 10.585 ;
  LAYER M2 ;
        RECT 27.6 10.499 30 10.501 ;
  LAYER M2 ;
        RECT 27.6 10.415 30 10.417 ;
  LAYER M2 ;
        RECT 27.6 10.331 30 10.333 ;
  LAYER M2 ;
        RECT 27.6 10.247 30 10.249 ;
  LAYER M2 ;
        RECT 27.6 10.163 30 10.165 ;
  LAYER M2 ;
        RECT 27.6 10.079 30 10.081 ;
  LAYER M2 ;
        RECT 27.6 9.995 30 9.997 ;
  LAYER M2 ;
        RECT 27.6 9.911 30 9.913 ;
  LAYER M2 ;
        RECT 27.6 9.827 30 9.829 ;
  LAYER M2 ;
        RECT 27.6 9.743 30 9.745 ;
  LAYER M2 ;
        RECT 27.6 9.659 30 9.661 ;
  LAYER M2 ;
        RECT 27.6 9.575 30 9.577 ;
  LAYER M1 ;
        RECT 29.984 6.516 30.016 9.024 ;
  LAYER M1 ;
        RECT 29.92 6.516 29.952 9.024 ;
  LAYER M1 ;
        RECT 29.856 6.516 29.888 9.024 ;
  LAYER M1 ;
        RECT 29.792 6.516 29.824 9.024 ;
  LAYER M1 ;
        RECT 29.728 6.516 29.76 9.024 ;
  LAYER M1 ;
        RECT 29.664 6.516 29.696 9.024 ;
  LAYER M1 ;
        RECT 29.6 6.516 29.632 9.024 ;
  LAYER M1 ;
        RECT 29.536 6.516 29.568 9.024 ;
  LAYER M1 ;
        RECT 29.472 6.516 29.504 9.024 ;
  LAYER M1 ;
        RECT 29.408 6.516 29.44 9.024 ;
  LAYER M1 ;
        RECT 29.344 6.516 29.376 9.024 ;
  LAYER M1 ;
        RECT 29.28 6.516 29.312 9.024 ;
  LAYER M1 ;
        RECT 29.216 6.516 29.248 9.024 ;
  LAYER M1 ;
        RECT 29.152 6.516 29.184 9.024 ;
  LAYER M1 ;
        RECT 29.088 6.516 29.12 9.024 ;
  LAYER M1 ;
        RECT 29.024 6.516 29.056 9.024 ;
  LAYER M1 ;
        RECT 28.96 6.516 28.992 9.024 ;
  LAYER M1 ;
        RECT 28.896 6.516 28.928 9.024 ;
  LAYER M1 ;
        RECT 28.832 6.516 28.864 9.024 ;
  LAYER M1 ;
        RECT 28.768 6.516 28.8 9.024 ;
  LAYER M1 ;
        RECT 28.704 6.516 28.736 9.024 ;
  LAYER M1 ;
        RECT 28.64 6.516 28.672 9.024 ;
  LAYER M1 ;
        RECT 28.576 6.516 28.608 9.024 ;
  LAYER M1 ;
        RECT 28.512 6.516 28.544 9.024 ;
  LAYER M1 ;
        RECT 28.448 6.516 28.48 9.024 ;
  LAYER M1 ;
        RECT 28.384 6.516 28.416 9.024 ;
  LAYER M1 ;
        RECT 28.32 6.516 28.352 9.024 ;
  LAYER M1 ;
        RECT 28.256 6.516 28.288 9.024 ;
  LAYER M1 ;
        RECT 28.192 6.516 28.224 9.024 ;
  LAYER M1 ;
        RECT 28.128 6.516 28.16 9.024 ;
  LAYER M1 ;
        RECT 28.064 6.516 28.096 9.024 ;
  LAYER M1 ;
        RECT 28 6.516 28.032 9.024 ;
  LAYER M1 ;
        RECT 27.936 6.516 27.968 9.024 ;
  LAYER M1 ;
        RECT 27.872 6.516 27.904 9.024 ;
  LAYER M1 ;
        RECT 27.808 6.516 27.84 9.024 ;
  LAYER M1 ;
        RECT 27.744 6.516 27.776 9.024 ;
  LAYER M1 ;
        RECT 27.68 6.516 27.712 9.024 ;
  LAYER M2 ;
        RECT 27.564 8.908 30.036 8.94 ;
  LAYER M2 ;
        RECT 27.564 8.844 30.036 8.876 ;
  LAYER M2 ;
        RECT 27.564 8.78 30.036 8.812 ;
  LAYER M2 ;
        RECT 27.564 8.716 30.036 8.748 ;
  LAYER M2 ;
        RECT 27.564 8.652 30.036 8.684 ;
  LAYER M2 ;
        RECT 27.564 8.588 30.036 8.62 ;
  LAYER M2 ;
        RECT 27.564 8.524 30.036 8.556 ;
  LAYER M2 ;
        RECT 27.564 8.46 30.036 8.492 ;
  LAYER M2 ;
        RECT 27.564 8.396 30.036 8.428 ;
  LAYER M2 ;
        RECT 27.564 8.332 30.036 8.364 ;
  LAYER M2 ;
        RECT 27.564 8.268 30.036 8.3 ;
  LAYER M2 ;
        RECT 27.564 8.204 30.036 8.236 ;
  LAYER M2 ;
        RECT 27.564 8.14 30.036 8.172 ;
  LAYER M2 ;
        RECT 27.564 8.076 30.036 8.108 ;
  LAYER M2 ;
        RECT 27.564 8.012 30.036 8.044 ;
  LAYER M2 ;
        RECT 27.564 7.948 30.036 7.98 ;
  LAYER M2 ;
        RECT 27.564 7.884 30.036 7.916 ;
  LAYER M2 ;
        RECT 27.564 7.82 30.036 7.852 ;
  LAYER M2 ;
        RECT 27.564 7.756 30.036 7.788 ;
  LAYER M2 ;
        RECT 27.564 7.692 30.036 7.724 ;
  LAYER M2 ;
        RECT 27.564 7.628 30.036 7.66 ;
  LAYER M2 ;
        RECT 27.564 7.564 30.036 7.596 ;
  LAYER M2 ;
        RECT 27.564 7.5 30.036 7.532 ;
  LAYER M2 ;
        RECT 27.564 7.436 30.036 7.468 ;
  LAYER M2 ;
        RECT 27.564 7.372 30.036 7.404 ;
  LAYER M2 ;
        RECT 27.564 7.308 30.036 7.34 ;
  LAYER M2 ;
        RECT 27.564 7.244 30.036 7.276 ;
  LAYER M2 ;
        RECT 27.564 7.18 30.036 7.212 ;
  LAYER M2 ;
        RECT 27.564 7.116 30.036 7.148 ;
  LAYER M2 ;
        RECT 27.564 7.052 30.036 7.084 ;
  LAYER M2 ;
        RECT 27.564 6.988 30.036 7.02 ;
  LAYER M2 ;
        RECT 27.564 6.924 30.036 6.956 ;
  LAYER M2 ;
        RECT 27.564 6.86 30.036 6.892 ;
  LAYER M2 ;
        RECT 27.564 6.796 30.036 6.828 ;
  LAYER M2 ;
        RECT 27.564 6.732 30.036 6.764 ;
  LAYER M2 ;
        RECT 27.564 6.668 30.036 6.7 ;
  LAYER M3 ;
        RECT 29.984 6.516 30.016 9.024 ;
  LAYER M3 ;
        RECT 29.92 6.516 29.952 9.024 ;
  LAYER M3 ;
        RECT 29.856 6.516 29.888 9.024 ;
  LAYER M3 ;
        RECT 29.792 6.516 29.824 9.024 ;
  LAYER M3 ;
        RECT 29.728 6.516 29.76 9.024 ;
  LAYER M3 ;
        RECT 29.664 6.516 29.696 9.024 ;
  LAYER M3 ;
        RECT 29.6 6.516 29.632 9.024 ;
  LAYER M3 ;
        RECT 29.536 6.516 29.568 9.024 ;
  LAYER M3 ;
        RECT 29.472 6.516 29.504 9.024 ;
  LAYER M3 ;
        RECT 29.408 6.516 29.44 9.024 ;
  LAYER M3 ;
        RECT 29.344 6.516 29.376 9.024 ;
  LAYER M3 ;
        RECT 29.28 6.516 29.312 9.024 ;
  LAYER M3 ;
        RECT 29.216 6.516 29.248 9.024 ;
  LAYER M3 ;
        RECT 29.152 6.516 29.184 9.024 ;
  LAYER M3 ;
        RECT 29.088 6.516 29.12 9.024 ;
  LAYER M3 ;
        RECT 29.024 6.516 29.056 9.024 ;
  LAYER M3 ;
        RECT 28.96 6.516 28.992 9.024 ;
  LAYER M3 ;
        RECT 28.896 6.516 28.928 9.024 ;
  LAYER M3 ;
        RECT 28.832 6.516 28.864 9.024 ;
  LAYER M3 ;
        RECT 28.768 6.516 28.8 9.024 ;
  LAYER M3 ;
        RECT 28.704 6.516 28.736 9.024 ;
  LAYER M3 ;
        RECT 28.64 6.516 28.672 9.024 ;
  LAYER M3 ;
        RECT 28.576 6.516 28.608 9.024 ;
  LAYER M3 ;
        RECT 28.512 6.516 28.544 9.024 ;
  LAYER M3 ;
        RECT 28.448 6.516 28.48 9.024 ;
  LAYER M3 ;
        RECT 28.384 6.516 28.416 9.024 ;
  LAYER M3 ;
        RECT 28.32 6.516 28.352 9.024 ;
  LAYER M3 ;
        RECT 28.256 6.516 28.288 9.024 ;
  LAYER M3 ;
        RECT 28.192 6.516 28.224 9.024 ;
  LAYER M3 ;
        RECT 28.128 6.516 28.16 9.024 ;
  LAYER M3 ;
        RECT 28.064 6.516 28.096 9.024 ;
  LAYER M3 ;
        RECT 28 6.516 28.032 9.024 ;
  LAYER M3 ;
        RECT 27.936 6.516 27.968 9.024 ;
  LAYER M3 ;
        RECT 27.872 6.516 27.904 9.024 ;
  LAYER M3 ;
        RECT 27.808 6.516 27.84 9.024 ;
  LAYER M3 ;
        RECT 27.744 6.516 27.776 9.024 ;
  LAYER M3 ;
        RECT 27.68 6.516 27.712 9.024 ;
  LAYER M3 ;
        RECT 27.584 6.516 27.616 9.024 ;
  LAYER M1 ;
        RECT 29.999 6.552 30.001 8.988 ;
  LAYER M1 ;
        RECT 29.919 6.552 29.921 8.988 ;
  LAYER M1 ;
        RECT 29.839 6.552 29.841 8.988 ;
  LAYER M1 ;
        RECT 29.759 6.552 29.761 8.988 ;
  LAYER M1 ;
        RECT 29.679 6.552 29.681 8.988 ;
  LAYER M1 ;
        RECT 29.599 6.552 29.601 8.988 ;
  LAYER M1 ;
        RECT 29.519 6.552 29.521 8.988 ;
  LAYER M1 ;
        RECT 29.439 6.552 29.441 8.988 ;
  LAYER M1 ;
        RECT 29.359 6.552 29.361 8.988 ;
  LAYER M1 ;
        RECT 29.279 6.552 29.281 8.988 ;
  LAYER M1 ;
        RECT 29.199 6.552 29.201 8.988 ;
  LAYER M1 ;
        RECT 29.119 6.552 29.121 8.988 ;
  LAYER M1 ;
        RECT 29.039 6.552 29.041 8.988 ;
  LAYER M1 ;
        RECT 28.959 6.552 28.961 8.988 ;
  LAYER M1 ;
        RECT 28.879 6.552 28.881 8.988 ;
  LAYER M1 ;
        RECT 28.799 6.552 28.801 8.988 ;
  LAYER M1 ;
        RECT 28.719 6.552 28.721 8.988 ;
  LAYER M1 ;
        RECT 28.639 6.552 28.641 8.988 ;
  LAYER M1 ;
        RECT 28.559 6.552 28.561 8.988 ;
  LAYER M1 ;
        RECT 28.479 6.552 28.481 8.988 ;
  LAYER M1 ;
        RECT 28.399 6.552 28.401 8.988 ;
  LAYER M1 ;
        RECT 28.319 6.552 28.321 8.988 ;
  LAYER M1 ;
        RECT 28.239 6.552 28.241 8.988 ;
  LAYER M1 ;
        RECT 28.159 6.552 28.161 8.988 ;
  LAYER M1 ;
        RECT 28.079 6.552 28.081 8.988 ;
  LAYER M1 ;
        RECT 27.999 6.552 28.001 8.988 ;
  LAYER M1 ;
        RECT 27.919 6.552 27.921 8.988 ;
  LAYER M1 ;
        RECT 27.839 6.552 27.841 8.988 ;
  LAYER M1 ;
        RECT 27.759 6.552 27.761 8.988 ;
  LAYER M1 ;
        RECT 27.679 6.552 27.681 8.988 ;
  LAYER M2 ;
        RECT 27.6 8.987 30 8.989 ;
  LAYER M2 ;
        RECT 27.6 8.903 30 8.905 ;
  LAYER M2 ;
        RECT 27.6 8.819 30 8.821 ;
  LAYER M2 ;
        RECT 27.6 8.735 30 8.737 ;
  LAYER M2 ;
        RECT 27.6 8.651 30 8.653 ;
  LAYER M2 ;
        RECT 27.6 8.567 30 8.569 ;
  LAYER M2 ;
        RECT 27.6 8.483 30 8.485 ;
  LAYER M2 ;
        RECT 27.6 8.399 30 8.401 ;
  LAYER M2 ;
        RECT 27.6 8.315 30 8.317 ;
  LAYER M2 ;
        RECT 27.6 8.231 30 8.233 ;
  LAYER M2 ;
        RECT 27.6 8.147 30 8.149 ;
  LAYER M2 ;
        RECT 27.6 8.063 30 8.065 ;
  LAYER M2 ;
        RECT 27.6 7.9795 30 7.9815 ;
  LAYER M2 ;
        RECT 27.6 7.895 30 7.897 ;
  LAYER M2 ;
        RECT 27.6 7.811 30 7.813 ;
  LAYER M2 ;
        RECT 27.6 7.727 30 7.729 ;
  LAYER M2 ;
        RECT 27.6 7.643 30 7.645 ;
  LAYER M2 ;
        RECT 27.6 7.559 30 7.561 ;
  LAYER M2 ;
        RECT 27.6 7.475 30 7.477 ;
  LAYER M2 ;
        RECT 27.6 7.391 30 7.393 ;
  LAYER M2 ;
        RECT 27.6 7.307 30 7.309 ;
  LAYER M2 ;
        RECT 27.6 7.223 30 7.225 ;
  LAYER M2 ;
        RECT 27.6 7.139 30 7.141 ;
  LAYER M2 ;
        RECT 27.6 7.055 30 7.057 ;
  LAYER M2 ;
        RECT 27.6 6.971 30 6.973 ;
  LAYER M2 ;
        RECT 27.6 6.887 30 6.889 ;
  LAYER M2 ;
        RECT 27.6 6.803 30 6.805 ;
  LAYER M2 ;
        RECT 27.6 6.719 30 6.721 ;
  LAYER M2 ;
        RECT 27.6 6.635 30 6.637 ;
  LAYER M1 ;
        RECT 27.104 15.336 27.136 17.844 ;
  LAYER M1 ;
        RECT 27.04 15.336 27.072 17.844 ;
  LAYER M1 ;
        RECT 26.976 15.336 27.008 17.844 ;
  LAYER M1 ;
        RECT 26.912 15.336 26.944 17.844 ;
  LAYER M1 ;
        RECT 26.848 15.336 26.88 17.844 ;
  LAYER M1 ;
        RECT 26.784 15.336 26.816 17.844 ;
  LAYER M1 ;
        RECT 26.72 15.336 26.752 17.844 ;
  LAYER M1 ;
        RECT 26.656 15.336 26.688 17.844 ;
  LAYER M1 ;
        RECT 26.592 15.336 26.624 17.844 ;
  LAYER M1 ;
        RECT 26.528 15.336 26.56 17.844 ;
  LAYER M1 ;
        RECT 26.464 15.336 26.496 17.844 ;
  LAYER M1 ;
        RECT 26.4 15.336 26.432 17.844 ;
  LAYER M1 ;
        RECT 26.336 15.336 26.368 17.844 ;
  LAYER M1 ;
        RECT 26.272 15.336 26.304 17.844 ;
  LAYER M1 ;
        RECT 26.208 15.336 26.24 17.844 ;
  LAYER M1 ;
        RECT 26.144 15.336 26.176 17.844 ;
  LAYER M1 ;
        RECT 26.08 15.336 26.112 17.844 ;
  LAYER M1 ;
        RECT 26.016 15.336 26.048 17.844 ;
  LAYER M1 ;
        RECT 25.952 15.336 25.984 17.844 ;
  LAYER M1 ;
        RECT 25.888 15.336 25.92 17.844 ;
  LAYER M1 ;
        RECT 25.824 15.336 25.856 17.844 ;
  LAYER M1 ;
        RECT 25.76 15.336 25.792 17.844 ;
  LAYER M1 ;
        RECT 25.696 15.336 25.728 17.844 ;
  LAYER M1 ;
        RECT 25.632 15.336 25.664 17.844 ;
  LAYER M1 ;
        RECT 25.568 15.336 25.6 17.844 ;
  LAYER M1 ;
        RECT 25.504 15.336 25.536 17.844 ;
  LAYER M1 ;
        RECT 25.44 15.336 25.472 17.844 ;
  LAYER M1 ;
        RECT 25.376 15.336 25.408 17.844 ;
  LAYER M1 ;
        RECT 25.312 15.336 25.344 17.844 ;
  LAYER M1 ;
        RECT 25.248 15.336 25.28 17.844 ;
  LAYER M1 ;
        RECT 25.184 15.336 25.216 17.844 ;
  LAYER M1 ;
        RECT 25.12 15.336 25.152 17.844 ;
  LAYER M1 ;
        RECT 25.056 15.336 25.088 17.844 ;
  LAYER M1 ;
        RECT 24.992 15.336 25.024 17.844 ;
  LAYER M1 ;
        RECT 24.928 15.336 24.96 17.844 ;
  LAYER M1 ;
        RECT 24.864 15.336 24.896 17.844 ;
  LAYER M1 ;
        RECT 24.8 15.336 24.832 17.844 ;
  LAYER M2 ;
        RECT 24.684 17.728 27.156 17.76 ;
  LAYER M2 ;
        RECT 24.684 17.664 27.156 17.696 ;
  LAYER M2 ;
        RECT 24.684 17.6 27.156 17.632 ;
  LAYER M2 ;
        RECT 24.684 17.536 27.156 17.568 ;
  LAYER M2 ;
        RECT 24.684 17.472 27.156 17.504 ;
  LAYER M2 ;
        RECT 24.684 17.408 27.156 17.44 ;
  LAYER M2 ;
        RECT 24.684 17.344 27.156 17.376 ;
  LAYER M2 ;
        RECT 24.684 17.28 27.156 17.312 ;
  LAYER M2 ;
        RECT 24.684 17.216 27.156 17.248 ;
  LAYER M2 ;
        RECT 24.684 17.152 27.156 17.184 ;
  LAYER M2 ;
        RECT 24.684 17.088 27.156 17.12 ;
  LAYER M2 ;
        RECT 24.684 17.024 27.156 17.056 ;
  LAYER M2 ;
        RECT 24.684 16.96 27.156 16.992 ;
  LAYER M2 ;
        RECT 24.684 16.896 27.156 16.928 ;
  LAYER M2 ;
        RECT 24.684 16.832 27.156 16.864 ;
  LAYER M2 ;
        RECT 24.684 16.768 27.156 16.8 ;
  LAYER M2 ;
        RECT 24.684 16.704 27.156 16.736 ;
  LAYER M2 ;
        RECT 24.684 16.64 27.156 16.672 ;
  LAYER M2 ;
        RECT 24.684 16.576 27.156 16.608 ;
  LAYER M2 ;
        RECT 24.684 16.512 27.156 16.544 ;
  LAYER M2 ;
        RECT 24.684 16.448 27.156 16.48 ;
  LAYER M2 ;
        RECT 24.684 16.384 27.156 16.416 ;
  LAYER M2 ;
        RECT 24.684 16.32 27.156 16.352 ;
  LAYER M2 ;
        RECT 24.684 16.256 27.156 16.288 ;
  LAYER M2 ;
        RECT 24.684 16.192 27.156 16.224 ;
  LAYER M2 ;
        RECT 24.684 16.128 27.156 16.16 ;
  LAYER M2 ;
        RECT 24.684 16.064 27.156 16.096 ;
  LAYER M2 ;
        RECT 24.684 16 27.156 16.032 ;
  LAYER M2 ;
        RECT 24.684 15.936 27.156 15.968 ;
  LAYER M2 ;
        RECT 24.684 15.872 27.156 15.904 ;
  LAYER M2 ;
        RECT 24.684 15.808 27.156 15.84 ;
  LAYER M2 ;
        RECT 24.684 15.744 27.156 15.776 ;
  LAYER M2 ;
        RECT 24.684 15.68 27.156 15.712 ;
  LAYER M2 ;
        RECT 24.684 15.616 27.156 15.648 ;
  LAYER M2 ;
        RECT 24.684 15.552 27.156 15.584 ;
  LAYER M2 ;
        RECT 24.684 15.488 27.156 15.52 ;
  LAYER M3 ;
        RECT 27.104 15.336 27.136 17.844 ;
  LAYER M3 ;
        RECT 27.04 15.336 27.072 17.844 ;
  LAYER M3 ;
        RECT 26.976 15.336 27.008 17.844 ;
  LAYER M3 ;
        RECT 26.912 15.336 26.944 17.844 ;
  LAYER M3 ;
        RECT 26.848 15.336 26.88 17.844 ;
  LAYER M3 ;
        RECT 26.784 15.336 26.816 17.844 ;
  LAYER M3 ;
        RECT 26.72 15.336 26.752 17.844 ;
  LAYER M3 ;
        RECT 26.656 15.336 26.688 17.844 ;
  LAYER M3 ;
        RECT 26.592 15.336 26.624 17.844 ;
  LAYER M3 ;
        RECT 26.528 15.336 26.56 17.844 ;
  LAYER M3 ;
        RECT 26.464 15.336 26.496 17.844 ;
  LAYER M3 ;
        RECT 26.4 15.336 26.432 17.844 ;
  LAYER M3 ;
        RECT 26.336 15.336 26.368 17.844 ;
  LAYER M3 ;
        RECT 26.272 15.336 26.304 17.844 ;
  LAYER M3 ;
        RECT 26.208 15.336 26.24 17.844 ;
  LAYER M3 ;
        RECT 26.144 15.336 26.176 17.844 ;
  LAYER M3 ;
        RECT 26.08 15.336 26.112 17.844 ;
  LAYER M3 ;
        RECT 26.016 15.336 26.048 17.844 ;
  LAYER M3 ;
        RECT 25.952 15.336 25.984 17.844 ;
  LAYER M3 ;
        RECT 25.888 15.336 25.92 17.844 ;
  LAYER M3 ;
        RECT 25.824 15.336 25.856 17.844 ;
  LAYER M3 ;
        RECT 25.76 15.336 25.792 17.844 ;
  LAYER M3 ;
        RECT 25.696 15.336 25.728 17.844 ;
  LAYER M3 ;
        RECT 25.632 15.336 25.664 17.844 ;
  LAYER M3 ;
        RECT 25.568 15.336 25.6 17.844 ;
  LAYER M3 ;
        RECT 25.504 15.336 25.536 17.844 ;
  LAYER M3 ;
        RECT 25.44 15.336 25.472 17.844 ;
  LAYER M3 ;
        RECT 25.376 15.336 25.408 17.844 ;
  LAYER M3 ;
        RECT 25.312 15.336 25.344 17.844 ;
  LAYER M3 ;
        RECT 25.248 15.336 25.28 17.844 ;
  LAYER M3 ;
        RECT 25.184 15.336 25.216 17.844 ;
  LAYER M3 ;
        RECT 25.12 15.336 25.152 17.844 ;
  LAYER M3 ;
        RECT 25.056 15.336 25.088 17.844 ;
  LAYER M3 ;
        RECT 24.992 15.336 25.024 17.844 ;
  LAYER M3 ;
        RECT 24.928 15.336 24.96 17.844 ;
  LAYER M3 ;
        RECT 24.864 15.336 24.896 17.844 ;
  LAYER M3 ;
        RECT 24.8 15.336 24.832 17.844 ;
  LAYER M3 ;
        RECT 24.704 15.336 24.736 17.844 ;
  LAYER M1 ;
        RECT 27.119 15.372 27.121 17.808 ;
  LAYER M1 ;
        RECT 27.039 15.372 27.041 17.808 ;
  LAYER M1 ;
        RECT 26.959 15.372 26.961 17.808 ;
  LAYER M1 ;
        RECT 26.879 15.372 26.881 17.808 ;
  LAYER M1 ;
        RECT 26.799 15.372 26.801 17.808 ;
  LAYER M1 ;
        RECT 26.719 15.372 26.721 17.808 ;
  LAYER M1 ;
        RECT 26.639 15.372 26.641 17.808 ;
  LAYER M1 ;
        RECT 26.559 15.372 26.561 17.808 ;
  LAYER M1 ;
        RECT 26.479 15.372 26.481 17.808 ;
  LAYER M1 ;
        RECT 26.399 15.372 26.401 17.808 ;
  LAYER M1 ;
        RECT 26.319 15.372 26.321 17.808 ;
  LAYER M1 ;
        RECT 26.239 15.372 26.241 17.808 ;
  LAYER M1 ;
        RECT 26.159 15.372 26.161 17.808 ;
  LAYER M1 ;
        RECT 26.079 15.372 26.081 17.808 ;
  LAYER M1 ;
        RECT 25.999 15.372 26.001 17.808 ;
  LAYER M1 ;
        RECT 25.919 15.372 25.921 17.808 ;
  LAYER M1 ;
        RECT 25.839 15.372 25.841 17.808 ;
  LAYER M1 ;
        RECT 25.759 15.372 25.761 17.808 ;
  LAYER M1 ;
        RECT 25.679 15.372 25.681 17.808 ;
  LAYER M1 ;
        RECT 25.599 15.372 25.601 17.808 ;
  LAYER M1 ;
        RECT 25.519 15.372 25.521 17.808 ;
  LAYER M1 ;
        RECT 25.439 15.372 25.441 17.808 ;
  LAYER M1 ;
        RECT 25.359 15.372 25.361 17.808 ;
  LAYER M1 ;
        RECT 25.279 15.372 25.281 17.808 ;
  LAYER M1 ;
        RECT 25.199 15.372 25.201 17.808 ;
  LAYER M1 ;
        RECT 25.119 15.372 25.121 17.808 ;
  LAYER M1 ;
        RECT 25.039 15.372 25.041 17.808 ;
  LAYER M1 ;
        RECT 24.959 15.372 24.961 17.808 ;
  LAYER M1 ;
        RECT 24.879 15.372 24.881 17.808 ;
  LAYER M1 ;
        RECT 24.799 15.372 24.801 17.808 ;
  LAYER M2 ;
        RECT 24.72 17.807 27.12 17.809 ;
  LAYER M2 ;
        RECT 24.72 17.723 27.12 17.725 ;
  LAYER M2 ;
        RECT 24.72 17.639 27.12 17.641 ;
  LAYER M2 ;
        RECT 24.72 17.555 27.12 17.557 ;
  LAYER M2 ;
        RECT 24.72 17.471 27.12 17.473 ;
  LAYER M2 ;
        RECT 24.72 17.387 27.12 17.389 ;
  LAYER M2 ;
        RECT 24.72 17.303 27.12 17.305 ;
  LAYER M2 ;
        RECT 24.72 17.219 27.12 17.221 ;
  LAYER M2 ;
        RECT 24.72 17.135 27.12 17.137 ;
  LAYER M2 ;
        RECT 24.72 17.051 27.12 17.053 ;
  LAYER M2 ;
        RECT 24.72 16.967 27.12 16.969 ;
  LAYER M2 ;
        RECT 24.72 16.883 27.12 16.885 ;
  LAYER M2 ;
        RECT 24.72 16.7995 27.12 16.8015 ;
  LAYER M2 ;
        RECT 24.72 16.715 27.12 16.717 ;
  LAYER M2 ;
        RECT 24.72 16.631 27.12 16.633 ;
  LAYER M2 ;
        RECT 24.72 16.547 27.12 16.549 ;
  LAYER M2 ;
        RECT 24.72 16.463 27.12 16.465 ;
  LAYER M2 ;
        RECT 24.72 16.379 27.12 16.381 ;
  LAYER M2 ;
        RECT 24.72 16.295 27.12 16.297 ;
  LAYER M2 ;
        RECT 24.72 16.211 27.12 16.213 ;
  LAYER M2 ;
        RECT 24.72 16.127 27.12 16.129 ;
  LAYER M2 ;
        RECT 24.72 16.043 27.12 16.045 ;
  LAYER M2 ;
        RECT 24.72 15.959 27.12 15.961 ;
  LAYER M2 ;
        RECT 24.72 15.875 27.12 15.877 ;
  LAYER M2 ;
        RECT 24.72 15.791 27.12 15.793 ;
  LAYER M2 ;
        RECT 24.72 15.707 27.12 15.709 ;
  LAYER M2 ;
        RECT 24.72 15.623 27.12 15.625 ;
  LAYER M2 ;
        RECT 24.72 15.539 27.12 15.541 ;
  LAYER M2 ;
        RECT 24.72 15.455 27.12 15.457 ;
  LAYER M1 ;
        RECT 27.104 12.396 27.136 14.904 ;
  LAYER M1 ;
        RECT 27.04 12.396 27.072 14.904 ;
  LAYER M1 ;
        RECT 26.976 12.396 27.008 14.904 ;
  LAYER M1 ;
        RECT 26.912 12.396 26.944 14.904 ;
  LAYER M1 ;
        RECT 26.848 12.396 26.88 14.904 ;
  LAYER M1 ;
        RECT 26.784 12.396 26.816 14.904 ;
  LAYER M1 ;
        RECT 26.72 12.396 26.752 14.904 ;
  LAYER M1 ;
        RECT 26.656 12.396 26.688 14.904 ;
  LAYER M1 ;
        RECT 26.592 12.396 26.624 14.904 ;
  LAYER M1 ;
        RECT 26.528 12.396 26.56 14.904 ;
  LAYER M1 ;
        RECT 26.464 12.396 26.496 14.904 ;
  LAYER M1 ;
        RECT 26.4 12.396 26.432 14.904 ;
  LAYER M1 ;
        RECT 26.336 12.396 26.368 14.904 ;
  LAYER M1 ;
        RECT 26.272 12.396 26.304 14.904 ;
  LAYER M1 ;
        RECT 26.208 12.396 26.24 14.904 ;
  LAYER M1 ;
        RECT 26.144 12.396 26.176 14.904 ;
  LAYER M1 ;
        RECT 26.08 12.396 26.112 14.904 ;
  LAYER M1 ;
        RECT 26.016 12.396 26.048 14.904 ;
  LAYER M1 ;
        RECT 25.952 12.396 25.984 14.904 ;
  LAYER M1 ;
        RECT 25.888 12.396 25.92 14.904 ;
  LAYER M1 ;
        RECT 25.824 12.396 25.856 14.904 ;
  LAYER M1 ;
        RECT 25.76 12.396 25.792 14.904 ;
  LAYER M1 ;
        RECT 25.696 12.396 25.728 14.904 ;
  LAYER M1 ;
        RECT 25.632 12.396 25.664 14.904 ;
  LAYER M1 ;
        RECT 25.568 12.396 25.6 14.904 ;
  LAYER M1 ;
        RECT 25.504 12.396 25.536 14.904 ;
  LAYER M1 ;
        RECT 25.44 12.396 25.472 14.904 ;
  LAYER M1 ;
        RECT 25.376 12.396 25.408 14.904 ;
  LAYER M1 ;
        RECT 25.312 12.396 25.344 14.904 ;
  LAYER M1 ;
        RECT 25.248 12.396 25.28 14.904 ;
  LAYER M1 ;
        RECT 25.184 12.396 25.216 14.904 ;
  LAYER M1 ;
        RECT 25.12 12.396 25.152 14.904 ;
  LAYER M1 ;
        RECT 25.056 12.396 25.088 14.904 ;
  LAYER M1 ;
        RECT 24.992 12.396 25.024 14.904 ;
  LAYER M1 ;
        RECT 24.928 12.396 24.96 14.904 ;
  LAYER M1 ;
        RECT 24.864 12.396 24.896 14.904 ;
  LAYER M1 ;
        RECT 24.8 12.396 24.832 14.904 ;
  LAYER M2 ;
        RECT 24.684 14.788 27.156 14.82 ;
  LAYER M2 ;
        RECT 24.684 14.724 27.156 14.756 ;
  LAYER M2 ;
        RECT 24.684 14.66 27.156 14.692 ;
  LAYER M2 ;
        RECT 24.684 14.596 27.156 14.628 ;
  LAYER M2 ;
        RECT 24.684 14.532 27.156 14.564 ;
  LAYER M2 ;
        RECT 24.684 14.468 27.156 14.5 ;
  LAYER M2 ;
        RECT 24.684 14.404 27.156 14.436 ;
  LAYER M2 ;
        RECT 24.684 14.34 27.156 14.372 ;
  LAYER M2 ;
        RECT 24.684 14.276 27.156 14.308 ;
  LAYER M2 ;
        RECT 24.684 14.212 27.156 14.244 ;
  LAYER M2 ;
        RECT 24.684 14.148 27.156 14.18 ;
  LAYER M2 ;
        RECT 24.684 14.084 27.156 14.116 ;
  LAYER M2 ;
        RECT 24.684 14.02 27.156 14.052 ;
  LAYER M2 ;
        RECT 24.684 13.956 27.156 13.988 ;
  LAYER M2 ;
        RECT 24.684 13.892 27.156 13.924 ;
  LAYER M2 ;
        RECT 24.684 13.828 27.156 13.86 ;
  LAYER M2 ;
        RECT 24.684 13.764 27.156 13.796 ;
  LAYER M2 ;
        RECT 24.684 13.7 27.156 13.732 ;
  LAYER M2 ;
        RECT 24.684 13.636 27.156 13.668 ;
  LAYER M2 ;
        RECT 24.684 13.572 27.156 13.604 ;
  LAYER M2 ;
        RECT 24.684 13.508 27.156 13.54 ;
  LAYER M2 ;
        RECT 24.684 13.444 27.156 13.476 ;
  LAYER M2 ;
        RECT 24.684 13.38 27.156 13.412 ;
  LAYER M2 ;
        RECT 24.684 13.316 27.156 13.348 ;
  LAYER M2 ;
        RECT 24.684 13.252 27.156 13.284 ;
  LAYER M2 ;
        RECT 24.684 13.188 27.156 13.22 ;
  LAYER M2 ;
        RECT 24.684 13.124 27.156 13.156 ;
  LAYER M2 ;
        RECT 24.684 13.06 27.156 13.092 ;
  LAYER M2 ;
        RECT 24.684 12.996 27.156 13.028 ;
  LAYER M2 ;
        RECT 24.684 12.932 27.156 12.964 ;
  LAYER M2 ;
        RECT 24.684 12.868 27.156 12.9 ;
  LAYER M2 ;
        RECT 24.684 12.804 27.156 12.836 ;
  LAYER M2 ;
        RECT 24.684 12.74 27.156 12.772 ;
  LAYER M2 ;
        RECT 24.684 12.676 27.156 12.708 ;
  LAYER M2 ;
        RECT 24.684 12.612 27.156 12.644 ;
  LAYER M2 ;
        RECT 24.684 12.548 27.156 12.58 ;
  LAYER M3 ;
        RECT 27.104 12.396 27.136 14.904 ;
  LAYER M3 ;
        RECT 27.04 12.396 27.072 14.904 ;
  LAYER M3 ;
        RECT 26.976 12.396 27.008 14.904 ;
  LAYER M3 ;
        RECT 26.912 12.396 26.944 14.904 ;
  LAYER M3 ;
        RECT 26.848 12.396 26.88 14.904 ;
  LAYER M3 ;
        RECT 26.784 12.396 26.816 14.904 ;
  LAYER M3 ;
        RECT 26.72 12.396 26.752 14.904 ;
  LAYER M3 ;
        RECT 26.656 12.396 26.688 14.904 ;
  LAYER M3 ;
        RECT 26.592 12.396 26.624 14.904 ;
  LAYER M3 ;
        RECT 26.528 12.396 26.56 14.904 ;
  LAYER M3 ;
        RECT 26.464 12.396 26.496 14.904 ;
  LAYER M3 ;
        RECT 26.4 12.396 26.432 14.904 ;
  LAYER M3 ;
        RECT 26.336 12.396 26.368 14.904 ;
  LAYER M3 ;
        RECT 26.272 12.396 26.304 14.904 ;
  LAYER M3 ;
        RECT 26.208 12.396 26.24 14.904 ;
  LAYER M3 ;
        RECT 26.144 12.396 26.176 14.904 ;
  LAYER M3 ;
        RECT 26.08 12.396 26.112 14.904 ;
  LAYER M3 ;
        RECT 26.016 12.396 26.048 14.904 ;
  LAYER M3 ;
        RECT 25.952 12.396 25.984 14.904 ;
  LAYER M3 ;
        RECT 25.888 12.396 25.92 14.904 ;
  LAYER M3 ;
        RECT 25.824 12.396 25.856 14.904 ;
  LAYER M3 ;
        RECT 25.76 12.396 25.792 14.904 ;
  LAYER M3 ;
        RECT 25.696 12.396 25.728 14.904 ;
  LAYER M3 ;
        RECT 25.632 12.396 25.664 14.904 ;
  LAYER M3 ;
        RECT 25.568 12.396 25.6 14.904 ;
  LAYER M3 ;
        RECT 25.504 12.396 25.536 14.904 ;
  LAYER M3 ;
        RECT 25.44 12.396 25.472 14.904 ;
  LAYER M3 ;
        RECT 25.376 12.396 25.408 14.904 ;
  LAYER M3 ;
        RECT 25.312 12.396 25.344 14.904 ;
  LAYER M3 ;
        RECT 25.248 12.396 25.28 14.904 ;
  LAYER M3 ;
        RECT 25.184 12.396 25.216 14.904 ;
  LAYER M3 ;
        RECT 25.12 12.396 25.152 14.904 ;
  LAYER M3 ;
        RECT 25.056 12.396 25.088 14.904 ;
  LAYER M3 ;
        RECT 24.992 12.396 25.024 14.904 ;
  LAYER M3 ;
        RECT 24.928 12.396 24.96 14.904 ;
  LAYER M3 ;
        RECT 24.864 12.396 24.896 14.904 ;
  LAYER M3 ;
        RECT 24.8 12.396 24.832 14.904 ;
  LAYER M3 ;
        RECT 24.704 12.396 24.736 14.904 ;
  LAYER M1 ;
        RECT 27.119 12.432 27.121 14.868 ;
  LAYER M1 ;
        RECT 27.039 12.432 27.041 14.868 ;
  LAYER M1 ;
        RECT 26.959 12.432 26.961 14.868 ;
  LAYER M1 ;
        RECT 26.879 12.432 26.881 14.868 ;
  LAYER M1 ;
        RECT 26.799 12.432 26.801 14.868 ;
  LAYER M1 ;
        RECT 26.719 12.432 26.721 14.868 ;
  LAYER M1 ;
        RECT 26.639 12.432 26.641 14.868 ;
  LAYER M1 ;
        RECT 26.559 12.432 26.561 14.868 ;
  LAYER M1 ;
        RECT 26.479 12.432 26.481 14.868 ;
  LAYER M1 ;
        RECT 26.399 12.432 26.401 14.868 ;
  LAYER M1 ;
        RECT 26.319 12.432 26.321 14.868 ;
  LAYER M1 ;
        RECT 26.239 12.432 26.241 14.868 ;
  LAYER M1 ;
        RECT 26.159 12.432 26.161 14.868 ;
  LAYER M1 ;
        RECT 26.079 12.432 26.081 14.868 ;
  LAYER M1 ;
        RECT 25.999 12.432 26.001 14.868 ;
  LAYER M1 ;
        RECT 25.919 12.432 25.921 14.868 ;
  LAYER M1 ;
        RECT 25.839 12.432 25.841 14.868 ;
  LAYER M1 ;
        RECT 25.759 12.432 25.761 14.868 ;
  LAYER M1 ;
        RECT 25.679 12.432 25.681 14.868 ;
  LAYER M1 ;
        RECT 25.599 12.432 25.601 14.868 ;
  LAYER M1 ;
        RECT 25.519 12.432 25.521 14.868 ;
  LAYER M1 ;
        RECT 25.439 12.432 25.441 14.868 ;
  LAYER M1 ;
        RECT 25.359 12.432 25.361 14.868 ;
  LAYER M1 ;
        RECT 25.279 12.432 25.281 14.868 ;
  LAYER M1 ;
        RECT 25.199 12.432 25.201 14.868 ;
  LAYER M1 ;
        RECT 25.119 12.432 25.121 14.868 ;
  LAYER M1 ;
        RECT 25.039 12.432 25.041 14.868 ;
  LAYER M1 ;
        RECT 24.959 12.432 24.961 14.868 ;
  LAYER M1 ;
        RECT 24.879 12.432 24.881 14.868 ;
  LAYER M1 ;
        RECT 24.799 12.432 24.801 14.868 ;
  LAYER M2 ;
        RECT 24.72 14.867 27.12 14.869 ;
  LAYER M2 ;
        RECT 24.72 14.783 27.12 14.785 ;
  LAYER M2 ;
        RECT 24.72 14.699 27.12 14.701 ;
  LAYER M2 ;
        RECT 24.72 14.615 27.12 14.617 ;
  LAYER M2 ;
        RECT 24.72 14.531 27.12 14.533 ;
  LAYER M2 ;
        RECT 24.72 14.447 27.12 14.449 ;
  LAYER M2 ;
        RECT 24.72 14.363 27.12 14.365 ;
  LAYER M2 ;
        RECT 24.72 14.279 27.12 14.281 ;
  LAYER M2 ;
        RECT 24.72 14.195 27.12 14.197 ;
  LAYER M2 ;
        RECT 24.72 14.111 27.12 14.113 ;
  LAYER M2 ;
        RECT 24.72 14.027 27.12 14.029 ;
  LAYER M2 ;
        RECT 24.72 13.943 27.12 13.945 ;
  LAYER M2 ;
        RECT 24.72 13.8595 27.12 13.8615 ;
  LAYER M2 ;
        RECT 24.72 13.775 27.12 13.777 ;
  LAYER M2 ;
        RECT 24.72 13.691 27.12 13.693 ;
  LAYER M2 ;
        RECT 24.72 13.607 27.12 13.609 ;
  LAYER M2 ;
        RECT 24.72 13.523 27.12 13.525 ;
  LAYER M2 ;
        RECT 24.72 13.439 27.12 13.441 ;
  LAYER M2 ;
        RECT 24.72 13.355 27.12 13.357 ;
  LAYER M2 ;
        RECT 24.72 13.271 27.12 13.273 ;
  LAYER M2 ;
        RECT 24.72 13.187 27.12 13.189 ;
  LAYER M2 ;
        RECT 24.72 13.103 27.12 13.105 ;
  LAYER M2 ;
        RECT 24.72 13.019 27.12 13.021 ;
  LAYER M2 ;
        RECT 24.72 12.935 27.12 12.937 ;
  LAYER M2 ;
        RECT 24.72 12.851 27.12 12.853 ;
  LAYER M2 ;
        RECT 24.72 12.767 27.12 12.769 ;
  LAYER M2 ;
        RECT 24.72 12.683 27.12 12.685 ;
  LAYER M2 ;
        RECT 24.72 12.599 27.12 12.601 ;
  LAYER M2 ;
        RECT 24.72 12.515 27.12 12.517 ;
  LAYER M1 ;
        RECT 27.104 9.456 27.136 11.964 ;
  LAYER M1 ;
        RECT 27.04 9.456 27.072 11.964 ;
  LAYER M1 ;
        RECT 26.976 9.456 27.008 11.964 ;
  LAYER M1 ;
        RECT 26.912 9.456 26.944 11.964 ;
  LAYER M1 ;
        RECT 26.848 9.456 26.88 11.964 ;
  LAYER M1 ;
        RECT 26.784 9.456 26.816 11.964 ;
  LAYER M1 ;
        RECT 26.72 9.456 26.752 11.964 ;
  LAYER M1 ;
        RECT 26.656 9.456 26.688 11.964 ;
  LAYER M1 ;
        RECT 26.592 9.456 26.624 11.964 ;
  LAYER M1 ;
        RECT 26.528 9.456 26.56 11.964 ;
  LAYER M1 ;
        RECT 26.464 9.456 26.496 11.964 ;
  LAYER M1 ;
        RECT 26.4 9.456 26.432 11.964 ;
  LAYER M1 ;
        RECT 26.336 9.456 26.368 11.964 ;
  LAYER M1 ;
        RECT 26.272 9.456 26.304 11.964 ;
  LAYER M1 ;
        RECT 26.208 9.456 26.24 11.964 ;
  LAYER M1 ;
        RECT 26.144 9.456 26.176 11.964 ;
  LAYER M1 ;
        RECT 26.08 9.456 26.112 11.964 ;
  LAYER M1 ;
        RECT 26.016 9.456 26.048 11.964 ;
  LAYER M1 ;
        RECT 25.952 9.456 25.984 11.964 ;
  LAYER M1 ;
        RECT 25.888 9.456 25.92 11.964 ;
  LAYER M1 ;
        RECT 25.824 9.456 25.856 11.964 ;
  LAYER M1 ;
        RECT 25.76 9.456 25.792 11.964 ;
  LAYER M1 ;
        RECT 25.696 9.456 25.728 11.964 ;
  LAYER M1 ;
        RECT 25.632 9.456 25.664 11.964 ;
  LAYER M1 ;
        RECT 25.568 9.456 25.6 11.964 ;
  LAYER M1 ;
        RECT 25.504 9.456 25.536 11.964 ;
  LAYER M1 ;
        RECT 25.44 9.456 25.472 11.964 ;
  LAYER M1 ;
        RECT 25.376 9.456 25.408 11.964 ;
  LAYER M1 ;
        RECT 25.312 9.456 25.344 11.964 ;
  LAYER M1 ;
        RECT 25.248 9.456 25.28 11.964 ;
  LAYER M1 ;
        RECT 25.184 9.456 25.216 11.964 ;
  LAYER M1 ;
        RECT 25.12 9.456 25.152 11.964 ;
  LAYER M1 ;
        RECT 25.056 9.456 25.088 11.964 ;
  LAYER M1 ;
        RECT 24.992 9.456 25.024 11.964 ;
  LAYER M1 ;
        RECT 24.928 9.456 24.96 11.964 ;
  LAYER M1 ;
        RECT 24.864 9.456 24.896 11.964 ;
  LAYER M1 ;
        RECT 24.8 9.456 24.832 11.964 ;
  LAYER M2 ;
        RECT 24.684 11.848 27.156 11.88 ;
  LAYER M2 ;
        RECT 24.684 11.784 27.156 11.816 ;
  LAYER M2 ;
        RECT 24.684 11.72 27.156 11.752 ;
  LAYER M2 ;
        RECT 24.684 11.656 27.156 11.688 ;
  LAYER M2 ;
        RECT 24.684 11.592 27.156 11.624 ;
  LAYER M2 ;
        RECT 24.684 11.528 27.156 11.56 ;
  LAYER M2 ;
        RECT 24.684 11.464 27.156 11.496 ;
  LAYER M2 ;
        RECT 24.684 11.4 27.156 11.432 ;
  LAYER M2 ;
        RECT 24.684 11.336 27.156 11.368 ;
  LAYER M2 ;
        RECT 24.684 11.272 27.156 11.304 ;
  LAYER M2 ;
        RECT 24.684 11.208 27.156 11.24 ;
  LAYER M2 ;
        RECT 24.684 11.144 27.156 11.176 ;
  LAYER M2 ;
        RECT 24.684 11.08 27.156 11.112 ;
  LAYER M2 ;
        RECT 24.684 11.016 27.156 11.048 ;
  LAYER M2 ;
        RECT 24.684 10.952 27.156 10.984 ;
  LAYER M2 ;
        RECT 24.684 10.888 27.156 10.92 ;
  LAYER M2 ;
        RECT 24.684 10.824 27.156 10.856 ;
  LAYER M2 ;
        RECT 24.684 10.76 27.156 10.792 ;
  LAYER M2 ;
        RECT 24.684 10.696 27.156 10.728 ;
  LAYER M2 ;
        RECT 24.684 10.632 27.156 10.664 ;
  LAYER M2 ;
        RECT 24.684 10.568 27.156 10.6 ;
  LAYER M2 ;
        RECT 24.684 10.504 27.156 10.536 ;
  LAYER M2 ;
        RECT 24.684 10.44 27.156 10.472 ;
  LAYER M2 ;
        RECT 24.684 10.376 27.156 10.408 ;
  LAYER M2 ;
        RECT 24.684 10.312 27.156 10.344 ;
  LAYER M2 ;
        RECT 24.684 10.248 27.156 10.28 ;
  LAYER M2 ;
        RECT 24.684 10.184 27.156 10.216 ;
  LAYER M2 ;
        RECT 24.684 10.12 27.156 10.152 ;
  LAYER M2 ;
        RECT 24.684 10.056 27.156 10.088 ;
  LAYER M2 ;
        RECT 24.684 9.992 27.156 10.024 ;
  LAYER M2 ;
        RECT 24.684 9.928 27.156 9.96 ;
  LAYER M2 ;
        RECT 24.684 9.864 27.156 9.896 ;
  LAYER M2 ;
        RECT 24.684 9.8 27.156 9.832 ;
  LAYER M2 ;
        RECT 24.684 9.736 27.156 9.768 ;
  LAYER M2 ;
        RECT 24.684 9.672 27.156 9.704 ;
  LAYER M2 ;
        RECT 24.684 9.608 27.156 9.64 ;
  LAYER M3 ;
        RECT 27.104 9.456 27.136 11.964 ;
  LAYER M3 ;
        RECT 27.04 9.456 27.072 11.964 ;
  LAYER M3 ;
        RECT 26.976 9.456 27.008 11.964 ;
  LAYER M3 ;
        RECT 26.912 9.456 26.944 11.964 ;
  LAYER M3 ;
        RECT 26.848 9.456 26.88 11.964 ;
  LAYER M3 ;
        RECT 26.784 9.456 26.816 11.964 ;
  LAYER M3 ;
        RECT 26.72 9.456 26.752 11.964 ;
  LAYER M3 ;
        RECT 26.656 9.456 26.688 11.964 ;
  LAYER M3 ;
        RECT 26.592 9.456 26.624 11.964 ;
  LAYER M3 ;
        RECT 26.528 9.456 26.56 11.964 ;
  LAYER M3 ;
        RECT 26.464 9.456 26.496 11.964 ;
  LAYER M3 ;
        RECT 26.4 9.456 26.432 11.964 ;
  LAYER M3 ;
        RECT 26.336 9.456 26.368 11.964 ;
  LAYER M3 ;
        RECT 26.272 9.456 26.304 11.964 ;
  LAYER M3 ;
        RECT 26.208 9.456 26.24 11.964 ;
  LAYER M3 ;
        RECT 26.144 9.456 26.176 11.964 ;
  LAYER M3 ;
        RECT 26.08 9.456 26.112 11.964 ;
  LAYER M3 ;
        RECT 26.016 9.456 26.048 11.964 ;
  LAYER M3 ;
        RECT 25.952 9.456 25.984 11.964 ;
  LAYER M3 ;
        RECT 25.888 9.456 25.92 11.964 ;
  LAYER M3 ;
        RECT 25.824 9.456 25.856 11.964 ;
  LAYER M3 ;
        RECT 25.76 9.456 25.792 11.964 ;
  LAYER M3 ;
        RECT 25.696 9.456 25.728 11.964 ;
  LAYER M3 ;
        RECT 25.632 9.456 25.664 11.964 ;
  LAYER M3 ;
        RECT 25.568 9.456 25.6 11.964 ;
  LAYER M3 ;
        RECT 25.504 9.456 25.536 11.964 ;
  LAYER M3 ;
        RECT 25.44 9.456 25.472 11.964 ;
  LAYER M3 ;
        RECT 25.376 9.456 25.408 11.964 ;
  LAYER M3 ;
        RECT 25.312 9.456 25.344 11.964 ;
  LAYER M3 ;
        RECT 25.248 9.456 25.28 11.964 ;
  LAYER M3 ;
        RECT 25.184 9.456 25.216 11.964 ;
  LAYER M3 ;
        RECT 25.12 9.456 25.152 11.964 ;
  LAYER M3 ;
        RECT 25.056 9.456 25.088 11.964 ;
  LAYER M3 ;
        RECT 24.992 9.456 25.024 11.964 ;
  LAYER M3 ;
        RECT 24.928 9.456 24.96 11.964 ;
  LAYER M3 ;
        RECT 24.864 9.456 24.896 11.964 ;
  LAYER M3 ;
        RECT 24.8 9.456 24.832 11.964 ;
  LAYER M3 ;
        RECT 24.704 9.456 24.736 11.964 ;
  LAYER M1 ;
        RECT 27.119 9.492 27.121 11.928 ;
  LAYER M1 ;
        RECT 27.039 9.492 27.041 11.928 ;
  LAYER M1 ;
        RECT 26.959 9.492 26.961 11.928 ;
  LAYER M1 ;
        RECT 26.879 9.492 26.881 11.928 ;
  LAYER M1 ;
        RECT 26.799 9.492 26.801 11.928 ;
  LAYER M1 ;
        RECT 26.719 9.492 26.721 11.928 ;
  LAYER M1 ;
        RECT 26.639 9.492 26.641 11.928 ;
  LAYER M1 ;
        RECT 26.559 9.492 26.561 11.928 ;
  LAYER M1 ;
        RECT 26.479 9.492 26.481 11.928 ;
  LAYER M1 ;
        RECT 26.399 9.492 26.401 11.928 ;
  LAYER M1 ;
        RECT 26.319 9.492 26.321 11.928 ;
  LAYER M1 ;
        RECT 26.239 9.492 26.241 11.928 ;
  LAYER M1 ;
        RECT 26.159 9.492 26.161 11.928 ;
  LAYER M1 ;
        RECT 26.079 9.492 26.081 11.928 ;
  LAYER M1 ;
        RECT 25.999 9.492 26.001 11.928 ;
  LAYER M1 ;
        RECT 25.919 9.492 25.921 11.928 ;
  LAYER M1 ;
        RECT 25.839 9.492 25.841 11.928 ;
  LAYER M1 ;
        RECT 25.759 9.492 25.761 11.928 ;
  LAYER M1 ;
        RECT 25.679 9.492 25.681 11.928 ;
  LAYER M1 ;
        RECT 25.599 9.492 25.601 11.928 ;
  LAYER M1 ;
        RECT 25.519 9.492 25.521 11.928 ;
  LAYER M1 ;
        RECT 25.439 9.492 25.441 11.928 ;
  LAYER M1 ;
        RECT 25.359 9.492 25.361 11.928 ;
  LAYER M1 ;
        RECT 25.279 9.492 25.281 11.928 ;
  LAYER M1 ;
        RECT 25.199 9.492 25.201 11.928 ;
  LAYER M1 ;
        RECT 25.119 9.492 25.121 11.928 ;
  LAYER M1 ;
        RECT 25.039 9.492 25.041 11.928 ;
  LAYER M1 ;
        RECT 24.959 9.492 24.961 11.928 ;
  LAYER M1 ;
        RECT 24.879 9.492 24.881 11.928 ;
  LAYER M1 ;
        RECT 24.799 9.492 24.801 11.928 ;
  LAYER M2 ;
        RECT 24.72 11.927 27.12 11.929 ;
  LAYER M2 ;
        RECT 24.72 11.843 27.12 11.845 ;
  LAYER M2 ;
        RECT 24.72 11.759 27.12 11.761 ;
  LAYER M2 ;
        RECT 24.72 11.675 27.12 11.677 ;
  LAYER M2 ;
        RECT 24.72 11.591 27.12 11.593 ;
  LAYER M2 ;
        RECT 24.72 11.507 27.12 11.509 ;
  LAYER M2 ;
        RECT 24.72 11.423 27.12 11.425 ;
  LAYER M2 ;
        RECT 24.72 11.339 27.12 11.341 ;
  LAYER M2 ;
        RECT 24.72 11.255 27.12 11.257 ;
  LAYER M2 ;
        RECT 24.72 11.171 27.12 11.173 ;
  LAYER M2 ;
        RECT 24.72 11.087 27.12 11.089 ;
  LAYER M2 ;
        RECT 24.72 11.003 27.12 11.005 ;
  LAYER M2 ;
        RECT 24.72 10.9195 27.12 10.9215 ;
  LAYER M2 ;
        RECT 24.72 10.835 27.12 10.837 ;
  LAYER M2 ;
        RECT 24.72 10.751 27.12 10.753 ;
  LAYER M2 ;
        RECT 24.72 10.667 27.12 10.669 ;
  LAYER M2 ;
        RECT 24.72 10.583 27.12 10.585 ;
  LAYER M2 ;
        RECT 24.72 10.499 27.12 10.501 ;
  LAYER M2 ;
        RECT 24.72 10.415 27.12 10.417 ;
  LAYER M2 ;
        RECT 24.72 10.331 27.12 10.333 ;
  LAYER M2 ;
        RECT 24.72 10.247 27.12 10.249 ;
  LAYER M2 ;
        RECT 24.72 10.163 27.12 10.165 ;
  LAYER M2 ;
        RECT 24.72 10.079 27.12 10.081 ;
  LAYER M2 ;
        RECT 24.72 9.995 27.12 9.997 ;
  LAYER M2 ;
        RECT 24.72 9.911 27.12 9.913 ;
  LAYER M2 ;
        RECT 24.72 9.827 27.12 9.829 ;
  LAYER M2 ;
        RECT 24.72 9.743 27.12 9.745 ;
  LAYER M2 ;
        RECT 24.72 9.659 27.12 9.661 ;
  LAYER M2 ;
        RECT 24.72 9.575 27.12 9.577 ;
  LAYER M1 ;
        RECT 27.104 6.516 27.136 9.024 ;
  LAYER M1 ;
        RECT 27.04 6.516 27.072 9.024 ;
  LAYER M1 ;
        RECT 26.976 6.516 27.008 9.024 ;
  LAYER M1 ;
        RECT 26.912 6.516 26.944 9.024 ;
  LAYER M1 ;
        RECT 26.848 6.516 26.88 9.024 ;
  LAYER M1 ;
        RECT 26.784 6.516 26.816 9.024 ;
  LAYER M1 ;
        RECT 26.72 6.516 26.752 9.024 ;
  LAYER M1 ;
        RECT 26.656 6.516 26.688 9.024 ;
  LAYER M1 ;
        RECT 26.592 6.516 26.624 9.024 ;
  LAYER M1 ;
        RECT 26.528 6.516 26.56 9.024 ;
  LAYER M1 ;
        RECT 26.464 6.516 26.496 9.024 ;
  LAYER M1 ;
        RECT 26.4 6.516 26.432 9.024 ;
  LAYER M1 ;
        RECT 26.336 6.516 26.368 9.024 ;
  LAYER M1 ;
        RECT 26.272 6.516 26.304 9.024 ;
  LAYER M1 ;
        RECT 26.208 6.516 26.24 9.024 ;
  LAYER M1 ;
        RECT 26.144 6.516 26.176 9.024 ;
  LAYER M1 ;
        RECT 26.08 6.516 26.112 9.024 ;
  LAYER M1 ;
        RECT 26.016 6.516 26.048 9.024 ;
  LAYER M1 ;
        RECT 25.952 6.516 25.984 9.024 ;
  LAYER M1 ;
        RECT 25.888 6.516 25.92 9.024 ;
  LAYER M1 ;
        RECT 25.824 6.516 25.856 9.024 ;
  LAYER M1 ;
        RECT 25.76 6.516 25.792 9.024 ;
  LAYER M1 ;
        RECT 25.696 6.516 25.728 9.024 ;
  LAYER M1 ;
        RECT 25.632 6.516 25.664 9.024 ;
  LAYER M1 ;
        RECT 25.568 6.516 25.6 9.024 ;
  LAYER M1 ;
        RECT 25.504 6.516 25.536 9.024 ;
  LAYER M1 ;
        RECT 25.44 6.516 25.472 9.024 ;
  LAYER M1 ;
        RECT 25.376 6.516 25.408 9.024 ;
  LAYER M1 ;
        RECT 25.312 6.516 25.344 9.024 ;
  LAYER M1 ;
        RECT 25.248 6.516 25.28 9.024 ;
  LAYER M1 ;
        RECT 25.184 6.516 25.216 9.024 ;
  LAYER M1 ;
        RECT 25.12 6.516 25.152 9.024 ;
  LAYER M1 ;
        RECT 25.056 6.516 25.088 9.024 ;
  LAYER M1 ;
        RECT 24.992 6.516 25.024 9.024 ;
  LAYER M1 ;
        RECT 24.928 6.516 24.96 9.024 ;
  LAYER M1 ;
        RECT 24.864 6.516 24.896 9.024 ;
  LAYER M1 ;
        RECT 24.8 6.516 24.832 9.024 ;
  LAYER M2 ;
        RECT 24.684 8.908 27.156 8.94 ;
  LAYER M2 ;
        RECT 24.684 8.844 27.156 8.876 ;
  LAYER M2 ;
        RECT 24.684 8.78 27.156 8.812 ;
  LAYER M2 ;
        RECT 24.684 8.716 27.156 8.748 ;
  LAYER M2 ;
        RECT 24.684 8.652 27.156 8.684 ;
  LAYER M2 ;
        RECT 24.684 8.588 27.156 8.62 ;
  LAYER M2 ;
        RECT 24.684 8.524 27.156 8.556 ;
  LAYER M2 ;
        RECT 24.684 8.46 27.156 8.492 ;
  LAYER M2 ;
        RECT 24.684 8.396 27.156 8.428 ;
  LAYER M2 ;
        RECT 24.684 8.332 27.156 8.364 ;
  LAYER M2 ;
        RECT 24.684 8.268 27.156 8.3 ;
  LAYER M2 ;
        RECT 24.684 8.204 27.156 8.236 ;
  LAYER M2 ;
        RECT 24.684 8.14 27.156 8.172 ;
  LAYER M2 ;
        RECT 24.684 8.076 27.156 8.108 ;
  LAYER M2 ;
        RECT 24.684 8.012 27.156 8.044 ;
  LAYER M2 ;
        RECT 24.684 7.948 27.156 7.98 ;
  LAYER M2 ;
        RECT 24.684 7.884 27.156 7.916 ;
  LAYER M2 ;
        RECT 24.684 7.82 27.156 7.852 ;
  LAYER M2 ;
        RECT 24.684 7.756 27.156 7.788 ;
  LAYER M2 ;
        RECT 24.684 7.692 27.156 7.724 ;
  LAYER M2 ;
        RECT 24.684 7.628 27.156 7.66 ;
  LAYER M2 ;
        RECT 24.684 7.564 27.156 7.596 ;
  LAYER M2 ;
        RECT 24.684 7.5 27.156 7.532 ;
  LAYER M2 ;
        RECT 24.684 7.436 27.156 7.468 ;
  LAYER M2 ;
        RECT 24.684 7.372 27.156 7.404 ;
  LAYER M2 ;
        RECT 24.684 7.308 27.156 7.34 ;
  LAYER M2 ;
        RECT 24.684 7.244 27.156 7.276 ;
  LAYER M2 ;
        RECT 24.684 7.18 27.156 7.212 ;
  LAYER M2 ;
        RECT 24.684 7.116 27.156 7.148 ;
  LAYER M2 ;
        RECT 24.684 7.052 27.156 7.084 ;
  LAYER M2 ;
        RECT 24.684 6.988 27.156 7.02 ;
  LAYER M2 ;
        RECT 24.684 6.924 27.156 6.956 ;
  LAYER M2 ;
        RECT 24.684 6.86 27.156 6.892 ;
  LAYER M2 ;
        RECT 24.684 6.796 27.156 6.828 ;
  LAYER M2 ;
        RECT 24.684 6.732 27.156 6.764 ;
  LAYER M2 ;
        RECT 24.684 6.668 27.156 6.7 ;
  LAYER M3 ;
        RECT 27.104 6.516 27.136 9.024 ;
  LAYER M3 ;
        RECT 27.04 6.516 27.072 9.024 ;
  LAYER M3 ;
        RECT 26.976 6.516 27.008 9.024 ;
  LAYER M3 ;
        RECT 26.912 6.516 26.944 9.024 ;
  LAYER M3 ;
        RECT 26.848 6.516 26.88 9.024 ;
  LAYER M3 ;
        RECT 26.784 6.516 26.816 9.024 ;
  LAYER M3 ;
        RECT 26.72 6.516 26.752 9.024 ;
  LAYER M3 ;
        RECT 26.656 6.516 26.688 9.024 ;
  LAYER M3 ;
        RECT 26.592 6.516 26.624 9.024 ;
  LAYER M3 ;
        RECT 26.528 6.516 26.56 9.024 ;
  LAYER M3 ;
        RECT 26.464 6.516 26.496 9.024 ;
  LAYER M3 ;
        RECT 26.4 6.516 26.432 9.024 ;
  LAYER M3 ;
        RECT 26.336 6.516 26.368 9.024 ;
  LAYER M3 ;
        RECT 26.272 6.516 26.304 9.024 ;
  LAYER M3 ;
        RECT 26.208 6.516 26.24 9.024 ;
  LAYER M3 ;
        RECT 26.144 6.516 26.176 9.024 ;
  LAYER M3 ;
        RECT 26.08 6.516 26.112 9.024 ;
  LAYER M3 ;
        RECT 26.016 6.516 26.048 9.024 ;
  LAYER M3 ;
        RECT 25.952 6.516 25.984 9.024 ;
  LAYER M3 ;
        RECT 25.888 6.516 25.92 9.024 ;
  LAYER M3 ;
        RECT 25.824 6.516 25.856 9.024 ;
  LAYER M3 ;
        RECT 25.76 6.516 25.792 9.024 ;
  LAYER M3 ;
        RECT 25.696 6.516 25.728 9.024 ;
  LAYER M3 ;
        RECT 25.632 6.516 25.664 9.024 ;
  LAYER M3 ;
        RECT 25.568 6.516 25.6 9.024 ;
  LAYER M3 ;
        RECT 25.504 6.516 25.536 9.024 ;
  LAYER M3 ;
        RECT 25.44 6.516 25.472 9.024 ;
  LAYER M3 ;
        RECT 25.376 6.516 25.408 9.024 ;
  LAYER M3 ;
        RECT 25.312 6.516 25.344 9.024 ;
  LAYER M3 ;
        RECT 25.248 6.516 25.28 9.024 ;
  LAYER M3 ;
        RECT 25.184 6.516 25.216 9.024 ;
  LAYER M3 ;
        RECT 25.12 6.516 25.152 9.024 ;
  LAYER M3 ;
        RECT 25.056 6.516 25.088 9.024 ;
  LAYER M3 ;
        RECT 24.992 6.516 25.024 9.024 ;
  LAYER M3 ;
        RECT 24.928 6.516 24.96 9.024 ;
  LAYER M3 ;
        RECT 24.864 6.516 24.896 9.024 ;
  LAYER M3 ;
        RECT 24.8 6.516 24.832 9.024 ;
  LAYER M3 ;
        RECT 24.704 6.516 24.736 9.024 ;
  LAYER M1 ;
        RECT 27.119 6.552 27.121 8.988 ;
  LAYER M1 ;
        RECT 27.039 6.552 27.041 8.988 ;
  LAYER M1 ;
        RECT 26.959 6.552 26.961 8.988 ;
  LAYER M1 ;
        RECT 26.879 6.552 26.881 8.988 ;
  LAYER M1 ;
        RECT 26.799 6.552 26.801 8.988 ;
  LAYER M1 ;
        RECT 26.719 6.552 26.721 8.988 ;
  LAYER M1 ;
        RECT 26.639 6.552 26.641 8.988 ;
  LAYER M1 ;
        RECT 26.559 6.552 26.561 8.988 ;
  LAYER M1 ;
        RECT 26.479 6.552 26.481 8.988 ;
  LAYER M1 ;
        RECT 26.399 6.552 26.401 8.988 ;
  LAYER M1 ;
        RECT 26.319 6.552 26.321 8.988 ;
  LAYER M1 ;
        RECT 26.239 6.552 26.241 8.988 ;
  LAYER M1 ;
        RECT 26.159 6.552 26.161 8.988 ;
  LAYER M1 ;
        RECT 26.079 6.552 26.081 8.988 ;
  LAYER M1 ;
        RECT 25.999 6.552 26.001 8.988 ;
  LAYER M1 ;
        RECT 25.919 6.552 25.921 8.988 ;
  LAYER M1 ;
        RECT 25.839 6.552 25.841 8.988 ;
  LAYER M1 ;
        RECT 25.759 6.552 25.761 8.988 ;
  LAYER M1 ;
        RECT 25.679 6.552 25.681 8.988 ;
  LAYER M1 ;
        RECT 25.599 6.552 25.601 8.988 ;
  LAYER M1 ;
        RECT 25.519 6.552 25.521 8.988 ;
  LAYER M1 ;
        RECT 25.439 6.552 25.441 8.988 ;
  LAYER M1 ;
        RECT 25.359 6.552 25.361 8.988 ;
  LAYER M1 ;
        RECT 25.279 6.552 25.281 8.988 ;
  LAYER M1 ;
        RECT 25.199 6.552 25.201 8.988 ;
  LAYER M1 ;
        RECT 25.119 6.552 25.121 8.988 ;
  LAYER M1 ;
        RECT 25.039 6.552 25.041 8.988 ;
  LAYER M1 ;
        RECT 24.959 6.552 24.961 8.988 ;
  LAYER M1 ;
        RECT 24.879 6.552 24.881 8.988 ;
  LAYER M1 ;
        RECT 24.799 6.552 24.801 8.988 ;
  LAYER M2 ;
        RECT 24.72 8.987 27.12 8.989 ;
  LAYER M2 ;
        RECT 24.72 8.903 27.12 8.905 ;
  LAYER M2 ;
        RECT 24.72 8.819 27.12 8.821 ;
  LAYER M2 ;
        RECT 24.72 8.735 27.12 8.737 ;
  LAYER M2 ;
        RECT 24.72 8.651 27.12 8.653 ;
  LAYER M2 ;
        RECT 24.72 8.567 27.12 8.569 ;
  LAYER M2 ;
        RECT 24.72 8.483 27.12 8.485 ;
  LAYER M2 ;
        RECT 24.72 8.399 27.12 8.401 ;
  LAYER M2 ;
        RECT 24.72 8.315 27.12 8.317 ;
  LAYER M2 ;
        RECT 24.72 8.231 27.12 8.233 ;
  LAYER M2 ;
        RECT 24.72 8.147 27.12 8.149 ;
  LAYER M2 ;
        RECT 24.72 8.063 27.12 8.065 ;
  LAYER M2 ;
        RECT 24.72 7.9795 27.12 7.9815 ;
  LAYER M2 ;
        RECT 24.72 7.895 27.12 7.897 ;
  LAYER M2 ;
        RECT 24.72 7.811 27.12 7.813 ;
  LAYER M2 ;
        RECT 24.72 7.727 27.12 7.729 ;
  LAYER M2 ;
        RECT 24.72 7.643 27.12 7.645 ;
  LAYER M2 ;
        RECT 24.72 7.559 27.12 7.561 ;
  LAYER M2 ;
        RECT 24.72 7.475 27.12 7.477 ;
  LAYER M2 ;
        RECT 24.72 7.391 27.12 7.393 ;
  LAYER M2 ;
        RECT 24.72 7.307 27.12 7.309 ;
  LAYER M2 ;
        RECT 24.72 7.223 27.12 7.225 ;
  LAYER M2 ;
        RECT 24.72 7.139 27.12 7.141 ;
  LAYER M2 ;
        RECT 24.72 7.055 27.12 7.057 ;
  LAYER M2 ;
        RECT 24.72 6.971 27.12 6.973 ;
  LAYER M2 ;
        RECT 24.72 6.887 27.12 6.889 ;
  LAYER M2 ;
        RECT 24.72 6.803 27.12 6.805 ;
  LAYER M2 ;
        RECT 24.72 6.719 27.12 6.721 ;
  LAYER M2 ;
        RECT 24.72 6.635 27.12 6.637 ;
  LAYER M1 ;
        RECT 24.224 15.336 24.256 17.844 ;
  LAYER M1 ;
        RECT 24.16 15.336 24.192 17.844 ;
  LAYER M1 ;
        RECT 24.096 15.336 24.128 17.844 ;
  LAYER M1 ;
        RECT 24.032 15.336 24.064 17.844 ;
  LAYER M1 ;
        RECT 23.968 15.336 24 17.844 ;
  LAYER M1 ;
        RECT 23.904 15.336 23.936 17.844 ;
  LAYER M1 ;
        RECT 23.84 15.336 23.872 17.844 ;
  LAYER M1 ;
        RECT 23.776 15.336 23.808 17.844 ;
  LAYER M1 ;
        RECT 23.712 15.336 23.744 17.844 ;
  LAYER M1 ;
        RECT 23.648 15.336 23.68 17.844 ;
  LAYER M1 ;
        RECT 23.584 15.336 23.616 17.844 ;
  LAYER M1 ;
        RECT 23.52 15.336 23.552 17.844 ;
  LAYER M1 ;
        RECT 23.456 15.336 23.488 17.844 ;
  LAYER M1 ;
        RECT 23.392 15.336 23.424 17.844 ;
  LAYER M1 ;
        RECT 23.328 15.336 23.36 17.844 ;
  LAYER M1 ;
        RECT 23.264 15.336 23.296 17.844 ;
  LAYER M1 ;
        RECT 23.2 15.336 23.232 17.844 ;
  LAYER M1 ;
        RECT 23.136 15.336 23.168 17.844 ;
  LAYER M1 ;
        RECT 23.072 15.336 23.104 17.844 ;
  LAYER M1 ;
        RECT 23.008 15.336 23.04 17.844 ;
  LAYER M1 ;
        RECT 22.944 15.336 22.976 17.844 ;
  LAYER M1 ;
        RECT 22.88 15.336 22.912 17.844 ;
  LAYER M1 ;
        RECT 22.816 15.336 22.848 17.844 ;
  LAYER M1 ;
        RECT 22.752 15.336 22.784 17.844 ;
  LAYER M1 ;
        RECT 22.688 15.336 22.72 17.844 ;
  LAYER M1 ;
        RECT 22.624 15.336 22.656 17.844 ;
  LAYER M1 ;
        RECT 22.56 15.336 22.592 17.844 ;
  LAYER M1 ;
        RECT 22.496 15.336 22.528 17.844 ;
  LAYER M1 ;
        RECT 22.432 15.336 22.464 17.844 ;
  LAYER M1 ;
        RECT 22.368 15.336 22.4 17.844 ;
  LAYER M1 ;
        RECT 22.304 15.336 22.336 17.844 ;
  LAYER M1 ;
        RECT 22.24 15.336 22.272 17.844 ;
  LAYER M1 ;
        RECT 22.176 15.336 22.208 17.844 ;
  LAYER M1 ;
        RECT 22.112 15.336 22.144 17.844 ;
  LAYER M1 ;
        RECT 22.048 15.336 22.08 17.844 ;
  LAYER M1 ;
        RECT 21.984 15.336 22.016 17.844 ;
  LAYER M1 ;
        RECT 21.92 15.336 21.952 17.844 ;
  LAYER M2 ;
        RECT 21.804 17.728 24.276 17.76 ;
  LAYER M2 ;
        RECT 21.804 17.664 24.276 17.696 ;
  LAYER M2 ;
        RECT 21.804 17.6 24.276 17.632 ;
  LAYER M2 ;
        RECT 21.804 17.536 24.276 17.568 ;
  LAYER M2 ;
        RECT 21.804 17.472 24.276 17.504 ;
  LAYER M2 ;
        RECT 21.804 17.408 24.276 17.44 ;
  LAYER M2 ;
        RECT 21.804 17.344 24.276 17.376 ;
  LAYER M2 ;
        RECT 21.804 17.28 24.276 17.312 ;
  LAYER M2 ;
        RECT 21.804 17.216 24.276 17.248 ;
  LAYER M2 ;
        RECT 21.804 17.152 24.276 17.184 ;
  LAYER M2 ;
        RECT 21.804 17.088 24.276 17.12 ;
  LAYER M2 ;
        RECT 21.804 17.024 24.276 17.056 ;
  LAYER M2 ;
        RECT 21.804 16.96 24.276 16.992 ;
  LAYER M2 ;
        RECT 21.804 16.896 24.276 16.928 ;
  LAYER M2 ;
        RECT 21.804 16.832 24.276 16.864 ;
  LAYER M2 ;
        RECT 21.804 16.768 24.276 16.8 ;
  LAYER M2 ;
        RECT 21.804 16.704 24.276 16.736 ;
  LAYER M2 ;
        RECT 21.804 16.64 24.276 16.672 ;
  LAYER M2 ;
        RECT 21.804 16.576 24.276 16.608 ;
  LAYER M2 ;
        RECT 21.804 16.512 24.276 16.544 ;
  LAYER M2 ;
        RECT 21.804 16.448 24.276 16.48 ;
  LAYER M2 ;
        RECT 21.804 16.384 24.276 16.416 ;
  LAYER M2 ;
        RECT 21.804 16.32 24.276 16.352 ;
  LAYER M2 ;
        RECT 21.804 16.256 24.276 16.288 ;
  LAYER M2 ;
        RECT 21.804 16.192 24.276 16.224 ;
  LAYER M2 ;
        RECT 21.804 16.128 24.276 16.16 ;
  LAYER M2 ;
        RECT 21.804 16.064 24.276 16.096 ;
  LAYER M2 ;
        RECT 21.804 16 24.276 16.032 ;
  LAYER M2 ;
        RECT 21.804 15.936 24.276 15.968 ;
  LAYER M2 ;
        RECT 21.804 15.872 24.276 15.904 ;
  LAYER M2 ;
        RECT 21.804 15.808 24.276 15.84 ;
  LAYER M2 ;
        RECT 21.804 15.744 24.276 15.776 ;
  LAYER M2 ;
        RECT 21.804 15.68 24.276 15.712 ;
  LAYER M2 ;
        RECT 21.804 15.616 24.276 15.648 ;
  LAYER M2 ;
        RECT 21.804 15.552 24.276 15.584 ;
  LAYER M2 ;
        RECT 21.804 15.488 24.276 15.52 ;
  LAYER M3 ;
        RECT 24.224 15.336 24.256 17.844 ;
  LAYER M3 ;
        RECT 24.16 15.336 24.192 17.844 ;
  LAYER M3 ;
        RECT 24.096 15.336 24.128 17.844 ;
  LAYER M3 ;
        RECT 24.032 15.336 24.064 17.844 ;
  LAYER M3 ;
        RECT 23.968 15.336 24 17.844 ;
  LAYER M3 ;
        RECT 23.904 15.336 23.936 17.844 ;
  LAYER M3 ;
        RECT 23.84 15.336 23.872 17.844 ;
  LAYER M3 ;
        RECT 23.776 15.336 23.808 17.844 ;
  LAYER M3 ;
        RECT 23.712 15.336 23.744 17.844 ;
  LAYER M3 ;
        RECT 23.648 15.336 23.68 17.844 ;
  LAYER M3 ;
        RECT 23.584 15.336 23.616 17.844 ;
  LAYER M3 ;
        RECT 23.52 15.336 23.552 17.844 ;
  LAYER M3 ;
        RECT 23.456 15.336 23.488 17.844 ;
  LAYER M3 ;
        RECT 23.392 15.336 23.424 17.844 ;
  LAYER M3 ;
        RECT 23.328 15.336 23.36 17.844 ;
  LAYER M3 ;
        RECT 23.264 15.336 23.296 17.844 ;
  LAYER M3 ;
        RECT 23.2 15.336 23.232 17.844 ;
  LAYER M3 ;
        RECT 23.136 15.336 23.168 17.844 ;
  LAYER M3 ;
        RECT 23.072 15.336 23.104 17.844 ;
  LAYER M3 ;
        RECT 23.008 15.336 23.04 17.844 ;
  LAYER M3 ;
        RECT 22.944 15.336 22.976 17.844 ;
  LAYER M3 ;
        RECT 22.88 15.336 22.912 17.844 ;
  LAYER M3 ;
        RECT 22.816 15.336 22.848 17.844 ;
  LAYER M3 ;
        RECT 22.752 15.336 22.784 17.844 ;
  LAYER M3 ;
        RECT 22.688 15.336 22.72 17.844 ;
  LAYER M3 ;
        RECT 22.624 15.336 22.656 17.844 ;
  LAYER M3 ;
        RECT 22.56 15.336 22.592 17.844 ;
  LAYER M3 ;
        RECT 22.496 15.336 22.528 17.844 ;
  LAYER M3 ;
        RECT 22.432 15.336 22.464 17.844 ;
  LAYER M3 ;
        RECT 22.368 15.336 22.4 17.844 ;
  LAYER M3 ;
        RECT 22.304 15.336 22.336 17.844 ;
  LAYER M3 ;
        RECT 22.24 15.336 22.272 17.844 ;
  LAYER M3 ;
        RECT 22.176 15.336 22.208 17.844 ;
  LAYER M3 ;
        RECT 22.112 15.336 22.144 17.844 ;
  LAYER M3 ;
        RECT 22.048 15.336 22.08 17.844 ;
  LAYER M3 ;
        RECT 21.984 15.336 22.016 17.844 ;
  LAYER M3 ;
        RECT 21.92 15.336 21.952 17.844 ;
  LAYER M3 ;
        RECT 21.824 15.336 21.856 17.844 ;
  LAYER M1 ;
        RECT 24.239 15.372 24.241 17.808 ;
  LAYER M1 ;
        RECT 24.159 15.372 24.161 17.808 ;
  LAYER M1 ;
        RECT 24.079 15.372 24.081 17.808 ;
  LAYER M1 ;
        RECT 23.999 15.372 24.001 17.808 ;
  LAYER M1 ;
        RECT 23.919 15.372 23.921 17.808 ;
  LAYER M1 ;
        RECT 23.839 15.372 23.841 17.808 ;
  LAYER M1 ;
        RECT 23.759 15.372 23.761 17.808 ;
  LAYER M1 ;
        RECT 23.679 15.372 23.681 17.808 ;
  LAYER M1 ;
        RECT 23.599 15.372 23.601 17.808 ;
  LAYER M1 ;
        RECT 23.519 15.372 23.521 17.808 ;
  LAYER M1 ;
        RECT 23.439 15.372 23.441 17.808 ;
  LAYER M1 ;
        RECT 23.359 15.372 23.361 17.808 ;
  LAYER M1 ;
        RECT 23.279 15.372 23.281 17.808 ;
  LAYER M1 ;
        RECT 23.199 15.372 23.201 17.808 ;
  LAYER M1 ;
        RECT 23.119 15.372 23.121 17.808 ;
  LAYER M1 ;
        RECT 23.039 15.372 23.041 17.808 ;
  LAYER M1 ;
        RECT 22.959 15.372 22.961 17.808 ;
  LAYER M1 ;
        RECT 22.879 15.372 22.881 17.808 ;
  LAYER M1 ;
        RECT 22.799 15.372 22.801 17.808 ;
  LAYER M1 ;
        RECT 22.719 15.372 22.721 17.808 ;
  LAYER M1 ;
        RECT 22.639 15.372 22.641 17.808 ;
  LAYER M1 ;
        RECT 22.559 15.372 22.561 17.808 ;
  LAYER M1 ;
        RECT 22.479 15.372 22.481 17.808 ;
  LAYER M1 ;
        RECT 22.399 15.372 22.401 17.808 ;
  LAYER M1 ;
        RECT 22.319 15.372 22.321 17.808 ;
  LAYER M1 ;
        RECT 22.239 15.372 22.241 17.808 ;
  LAYER M1 ;
        RECT 22.159 15.372 22.161 17.808 ;
  LAYER M1 ;
        RECT 22.079 15.372 22.081 17.808 ;
  LAYER M1 ;
        RECT 21.999 15.372 22.001 17.808 ;
  LAYER M1 ;
        RECT 21.919 15.372 21.921 17.808 ;
  LAYER M2 ;
        RECT 21.84 17.807 24.24 17.809 ;
  LAYER M2 ;
        RECT 21.84 17.723 24.24 17.725 ;
  LAYER M2 ;
        RECT 21.84 17.639 24.24 17.641 ;
  LAYER M2 ;
        RECT 21.84 17.555 24.24 17.557 ;
  LAYER M2 ;
        RECT 21.84 17.471 24.24 17.473 ;
  LAYER M2 ;
        RECT 21.84 17.387 24.24 17.389 ;
  LAYER M2 ;
        RECT 21.84 17.303 24.24 17.305 ;
  LAYER M2 ;
        RECT 21.84 17.219 24.24 17.221 ;
  LAYER M2 ;
        RECT 21.84 17.135 24.24 17.137 ;
  LAYER M2 ;
        RECT 21.84 17.051 24.24 17.053 ;
  LAYER M2 ;
        RECT 21.84 16.967 24.24 16.969 ;
  LAYER M2 ;
        RECT 21.84 16.883 24.24 16.885 ;
  LAYER M2 ;
        RECT 21.84 16.7995 24.24 16.8015 ;
  LAYER M2 ;
        RECT 21.84 16.715 24.24 16.717 ;
  LAYER M2 ;
        RECT 21.84 16.631 24.24 16.633 ;
  LAYER M2 ;
        RECT 21.84 16.547 24.24 16.549 ;
  LAYER M2 ;
        RECT 21.84 16.463 24.24 16.465 ;
  LAYER M2 ;
        RECT 21.84 16.379 24.24 16.381 ;
  LAYER M2 ;
        RECT 21.84 16.295 24.24 16.297 ;
  LAYER M2 ;
        RECT 21.84 16.211 24.24 16.213 ;
  LAYER M2 ;
        RECT 21.84 16.127 24.24 16.129 ;
  LAYER M2 ;
        RECT 21.84 16.043 24.24 16.045 ;
  LAYER M2 ;
        RECT 21.84 15.959 24.24 15.961 ;
  LAYER M2 ;
        RECT 21.84 15.875 24.24 15.877 ;
  LAYER M2 ;
        RECT 21.84 15.791 24.24 15.793 ;
  LAYER M2 ;
        RECT 21.84 15.707 24.24 15.709 ;
  LAYER M2 ;
        RECT 21.84 15.623 24.24 15.625 ;
  LAYER M2 ;
        RECT 21.84 15.539 24.24 15.541 ;
  LAYER M2 ;
        RECT 21.84 15.455 24.24 15.457 ;
  LAYER M1 ;
        RECT 24.224 12.396 24.256 14.904 ;
  LAYER M1 ;
        RECT 24.16 12.396 24.192 14.904 ;
  LAYER M1 ;
        RECT 24.096 12.396 24.128 14.904 ;
  LAYER M1 ;
        RECT 24.032 12.396 24.064 14.904 ;
  LAYER M1 ;
        RECT 23.968 12.396 24 14.904 ;
  LAYER M1 ;
        RECT 23.904 12.396 23.936 14.904 ;
  LAYER M1 ;
        RECT 23.84 12.396 23.872 14.904 ;
  LAYER M1 ;
        RECT 23.776 12.396 23.808 14.904 ;
  LAYER M1 ;
        RECT 23.712 12.396 23.744 14.904 ;
  LAYER M1 ;
        RECT 23.648 12.396 23.68 14.904 ;
  LAYER M1 ;
        RECT 23.584 12.396 23.616 14.904 ;
  LAYER M1 ;
        RECT 23.52 12.396 23.552 14.904 ;
  LAYER M1 ;
        RECT 23.456 12.396 23.488 14.904 ;
  LAYER M1 ;
        RECT 23.392 12.396 23.424 14.904 ;
  LAYER M1 ;
        RECT 23.328 12.396 23.36 14.904 ;
  LAYER M1 ;
        RECT 23.264 12.396 23.296 14.904 ;
  LAYER M1 ;
        RECT 23.2 12.396 23.232 14.904 ;
  LAYER M1 ;
        RECT 23.136 12.396 23.168 14.904 ;
  LAYER M1 ;
        RECT 23.072 12.396 23.104 14.904 ;
  LAYER M1 ;
        RECT 23.008 12.396 23.04 14.904 ;
  LAYER M1 ;
        RECT 22.944 12.396 22.976 14.904 ;
  LAYER M1 ;
        RECT 22.88 12.396 22.912 14.904 ;
  LAYER M1 ;
        RECT 22.816 12.396 22.848 14.904 ;
  LAYER M1 ;
        RECT 22.752 12.396 22.784 14.904 ;
  LAYER M1 ;
        RECT 22.688 12.396 22.72 14.904 ;
  LAYER M1 ;
        RECT 22.624 12.396 22.656 14.904 ;
  LAYER M1 ;
        RECT 22.56 12.396 22.592 14.904 ;
  LAYER M1 ;
        RECT 22.496 12.396 22.528 14.904 ;
  LAYER M1 ;
        RECT 22.432 12.396 22.464 14.904 ;
  LAYER M1 ;
        RECT 22.368 12.396 22.4 14.904 ;
  LAYER M1 ;
        RECT 22.304 12.396 22.336 14.904 ;
  LAYER M1 ;
        RECT 22.24 12.396 22.272 14.904 ;
  LAYER M1 ;
        RECT 22.176 12.396 22.208 14.904 ;
  LAYER M1 ;
        RECT 22.112 12.396 22.144 14.904 ;
  LAYER M1 ;
        RECT 22.048 12.396 22.08 14.904 ;
  LAYER M1 ;
        RECT 21.984 12.396 22.016 14.904 ;
  LAYER M1 ;
        RECT 21.92 12.396 21.952 14.904 ;
  LAYER M2 ;
        RECT 21.804 14.788 24.276 14.82 ;
  LAYER M2 ;
        RECT 21.804 14.724 24.276 14.756 ;
  LAYER M2 ;
        RECT 21.804 14.66 24.276 14.692 ;
  LAYER M2 ;
        RECT 21.804 14.596 24.276 14.628 ;
  LAYER M2 ;
        RECT 21.804 14.532 24.276 14.564 ;
  LAYER M2 ;
        RECT 21.804 14.468 24.276 14.5 ;
  LAYER M2 ;
        RECT 21.804 14.404 24.276 14.436 ;
  LAYER M2 ;
        RECT 21.804 14.34 24.276 14.372 ;
  LAYER M2 ;
        RECT 21.804 14.276 24.276 14.308 ;
  LAYER M2 ;
        RECT 21.804 14.212 24.276 14.244 ;
  LAYER M2 ;
        RECT 21.804 14.148 24.276 14.18 ;
  LAYER M2 ;
        RECT 21.804 14.084 24.276 14.116 ;
  LAYER M2 ;
        RECT 21.804 14.02 24.276 14.052 ;
  LAYER M2 ;
        RECT 21.804 13.956 24.276 13.988 ;
  LAYER M2 ;
        RECT 21.804 13.892 24.276 13.924 ;
  LAYER M2 ;
        RECT 21.804 13.828 24.276 13.86 ;
  LAYER M2 ;
        RECT 21.804 13.764 24.276 13.796 ;
  LAYER M2 ;
        RECT 21.804 13.7 24.276 13.732 ;
  LAYER M2 ;
        RECT 21.804 13.636 24.276 13.668 ;
  LAYER M2 ;
        RECT 21.804 13.572 24.276 13.604 ;
  LAYER M2 ;
        RECT 21.804 13.508 24.276 13.54 ;
  LAYER M2 ;
        RECT 21.804 13.444 24.276 13.476 ;
  LAYER M2 ;
        RECT 21.804 13.38 24.276 13.412 ;
  LAYER M2 ;
        RECT 21.804 13.316 24.276 13.348 ;
  LAYER M2 ;
        RECT 21.804 13.252 24.276 13.284 ;
  LAYER M2 ;
        RECT 21.804 13.188 24.276 13.22 ;
  LAYER M2 ;
        RECT 21.804 13.124 24.276 13.156 ;
  LAYER M2 ;
        RECT 21.804 13.06 24.276 13.092 ;
  LAYER M2 ;
        RECT 21.804 12.996 24.276 13.028 ;
  LAYER M2 ;
        RECT 21.804 12.932 24.276 12.964 ;
  LAYER M2 ;
        RECT 21.804 12.868 24.276 12.9 ;
  LAYER M2 ;
        RECT 21.804 12.804 24.276 12.836 ;
  LAYER M2 ;
        RECT 21.804 12.74 24.276 12.772 ;
  LAYER M2 ;
        RECT 21.804 12.676 24.276 12.708 ;
  LAYER M2 ;
        RECT 21.804 12.612 24.276 12.644 ;
  LAYER M2 ;
        RECT 21.804 12.548 24.276 12.58 ;
  LAYER M3 ;
        RECT 24.224 12.396 24.256 14.904 ;
  LAYER M3 ;
        RECT 24.16 12.396 24.192 14.904 ;
  LAYER M3 ;
        RECT 24.096 12.396 24.128 14.904 ;
  LAYER M3 ;
        RECT 24.032 12.396 24.064 14.904 ;
  LAYER M3 ;
        RECT 23.968 12.396 24 14.904 ;
  LAYER M3 ;
        RECT 23.904 12.396 23.936 14.904 ;
  LAYER M3 ;
        RECT 23.84 12.396 23.872 14.904 ;
  LAYER M3 ;
        RECT 23.776 12.396 23.808 14.904 ;
  LAYER M3 ;
        RECT 23.712 12.396 23.744 14.904 ;
  LAYER M3 ;
        RECT 23.648 12.396 23.68 14.904 ;
  LAYER M3 ;
        RECT 23.584 12.396 23.616 14.904 ;
  LAYER M3 ;
        RECT 23.52 12.396 23.552 14.904 ;
  LAYER M3 ;
        RECT 23.456 12.396 23.488 14.904 ;
  LAYER M3 ;
        RECT 23.392 12.396 23.424 14.904 ;
  LAYER M3 ;
        RECT 23.328 12.396 23.36 14.904 ;
  LAYER M3 ;
        RECT 23.264 12.396 23.296 14.904 ;
  LAYER M3 ;
        RECT 23.2 12.396 23.232 14.904 ;
  LAYER M3 ;
        RECT 23.136 12.396 23.168 14.904 ;
  LAYER M3 ;
        RECT 23.072 12.396 23.104 14.904 ;
  LAYER M3 ;
        RECT 23.008 12.396 23.04 14.904 ;
  LAYER M3 ;
        RECT 22.944 12.396 22.976 14.904 ;
  LAYER M3 ;
        RECT 22.88 12.396 22.912 14.904 ;
  LAYER M3 ;
        RECT 22.816 12.396 22.848 14.904 ;
  LAYER M3 ;
        RECT 22.752 12.396 22.784 14.904 ;
  LAYER M3 ;
        RECT 22.688 12.396 22.72 14.904 ;
  LAYER M3 ;
        RECT 22.624 12.396 22.656 14.904 ;
  LAYER M3 ;
        RECT 22.56 12.396 22.592 14.904 ;
  LAYER M3 ;
        RECT 22.496 12.396 22.528 14.904 ;
  LAYER M3 ;
        RECT 22.432 12.396 22.464 14.904 ;
  LAYER M3 ;
        RECT 22.368 12.396 22.4 14.904 ;
  LAYER M3 ;
        RECT 22.304 12.396 22.336 14.904 ;
  LAYER M3 ;
        RECT 22.24 12.396 22.272 14.904 ;
  LAYER M3 ;
        RECT 22.176 12.396 22.208 14.904 ;
  LAYER M3 ;
        RECT 22.112 12.396 22.144 14.904 ;
  LAYER M3 ;
        RECT 22.048 12.396 22.08 14.904 ;
  LAYER M3 ;
        RECT 21.984 12.396 22.016 14.904 ;
  LAYER M3 ;
        RECT 21.92 12.396 21.952 14.904 ;
  LAYER M3 ;
        RECT 21.824 12.396 21.856 14.904 ;
  LAYER M1 ;
        RECT 24.239 12.432 24.241 14.868 ;
  LAYER M1 ;
        RECT 24.159 12.432 24.161 14.868 ;
  LAYER M1 ;
        RECT 24.079 12.432 24.081 14.868 ;
  LAYER M1 ;
        RECT 23.999 12.432 24.001 14.868 ;
  LAYER M1 ;
        RECT 23.919 12.432 23.921 14.868 ;
  LAYER M1 ;
        RECT 23.839 12.432 23.841 14.868 ;
  LAYER M1 ;
        RECT 23.759 12.432 23.761 14.868 ;
  LAYER M1 ;
        RECT 23.679 12.432 23.681 14.868 ;
  LAYER M1 ;
        RECT 23.599 12.432 23.601 14.868 ;
  LAYER M1 ;
        RECT 23.519 12.432 23.521 14.868 ;
  LAYER M1 ;
        RECT 23.439 12.432 23.441 14.868 ;
  LAYER M1 ;
        RECT 23.359 12.432 23.361 14.868 ;
  LAYER M1 ;
        RECT 23.279 12.432 23.281 14.868 ;
  LAYER M1 ;
        RECT 23.199 12.432 23.201 14.868 ;
  LAYER M1 ;
        RECT 23.119 12.432 23.121 14.868 ;
  LAYER M1 ;
        RECT 23.039 12.432 23.041 14.868 ;
  LAYER M1 ;
        RECT 22.959 12.432 22.961 14.868 ;
  LAYER M1 ;
        RECT 22.879 12.432 22.881 14.868 ;
  LAYER M1 ;
        RECT 22.799 12.432 22.801 14.868 ;
  LAYER M1 ;
        RECT 22.719 12.432 22.721 14.868 ;
  LAYER M1 ;
        RECT 22.639 12.432 22.641 14.868 ;
  LAYER M1 ;
        RECT 22.559 12.432 22.561 14.868 ;
  LAYER M1 ;
        RECT 22.479 12.432 22.481 14.868 ;
  LAYER M1 ;
        RECT 22.399 12.432 22.401 14.868 ;
  LAYER M1 ;
        RECT 22.319 12.432 22.321 14.868 ;
  LAYER M1 ;
        RECT 22.239 12.432 22.241 14.868 ;
  LAYER M1 ;
        RECT 22.159 12.432 22.161 14.868 ;
  LAYER M1 ;
        RECT 22.079 12.432 22.081 14.868 ;
  LAYER M1 ;
        RECT 21.999 12.432 22.001 14.868 ;
  LAYER M1 ;
        RECT 21.919 12.432 21.921 14.868 ;
  LAYER M2 ;
        RECT 21.84 14.867 24.24 14.869 ;
  LAYER M2 ;
        RECT 21.84 14.783 24.24 14.785 ;
  LAYER M2 ;
        RECT 21.84 14.699 24.24 14.701 ;
  LAYER M2 ;
        RECT 21.84 14.615 24.24 14.617 ;
  LAYER M2 ;
        RECT 21.84 14.531 24.24 14.533 ;
  LAYER M2 ;
        RECT 21.84 14.447 24.24 14.449 ;
  LAYER M2 ;
        RECT 21.84 14.363 24.24 14.365 ;
  LAYER M2 ;
        RECT 21.84 14.279 24.24 14.281 ;
  LAYER M2 ;
        RECT 21.84 14.195 24.24 14.197 ;
  LAYER M2 ;
        RECT 21.84 14.111 24.24 14.113 ;
  LAYER M2 ;
        RECT 21.84 14.027 24.24 14.029 ;
  LAYER M2 ;
        RECT 21.84 13.943 24.24 13.945 ;
  LAYER M2 ;
        RECT 21.84 13.8595 24.24 13.8615 ;
  LAYER M2 ;
        RECT 21.84 13.775 24.24 13.777 ;
  LAYER M2 ;
        RECT 21.84 13.691 24.24 13.693 ;
  LAYER M2 ;
        RECT 21.84 13.607 24.24 13.609 ;
  LAYER M2 ;
        RECT 21.84 13.523 24.24 13.525 ;
  LAYER M2 ;
        RECT 21.84 13.439 24.24 13.441 ;
  LAYER M2 ;
        RECT 21.84 13.355 24.24 13.357 ;
  LAYER M2 ;
        RECT 21.84 13.271 24.24 13.273 ;
  LAYER M2 ;
        RECT 21.84 13.187 24.24 13.189 ;
  LAYER M2 ;
        RECT 21.84 13.103 24.24 13.105 ;
  LAYER M2 ;
        RECT 21.84 13.019 24.24 13.021 ;
  LAYER M2 ;
        RECT 21.84 12.935 24.24 12.937 ;
  LAYER M2 ;
        RECT 21.84 12.851 24.24 12.853 ;
  LAYER M2 ;
        RECT 21.84 12.767 24.24 12.769 ;
  LAYER M2 ;
        RECT 21.84 12.683 24.24 12.685 ;
  LAYER M2 ;
        RECT 21.84 12.599 24.24 12.601 ;
  LAYER M2 ;
        RECT 21.84 12.515 24.24 12.517 ;
  LAYER M1 ;
        RECT 24.224 9.456 24.256 11.964 ;
  LAYER M1 ;
        RECT 24.16 9.456 24.192 11.964 ;
  LAYER M1 ;
        RECT 24.096 9.456 24.128 11.964 ;
  LAYER M1 ;
        RECT 24.032 9.456 24.064 11.964 ;
  LAYER M1 ;
        RECT 23.968 9.456 24 11.964 ;
  LAYER M1 ;
        RECT 23.904 9.456 23.936 11.964 ;
  LAYER M1 ;
        RECT 23.84 9.456 23.872 11.964 ;
  LAYER M1 ;
        RECT 23.776 9.456 23.808 11.964 ;
  LAYER M1 ;
        RECT 23.712 9.456 23.744 11.964 ;
  LAYER M1 ;
        RECT 23.648 9.456 23.68 11.964 ;
  LAYER M1 ;
        RECT 23.584 9.456 23.616 11.964 ;
  LAYER M1 ;
        RECT 23.52 9.456 23.552 11.964 ;
  LAYER M1 ;
        RECT 23.456 9.456 23.488 11.964 ;
  LAYER M1 ;
        RECT 23.392 9.456 23.424 11.964 ;
  LAYER M1 ;
        RECT 23.328 9.456 23.36 11.964 ;
  LAYER M1 ;
        RECT 23.264 9.456 23.296 11.964 ;
  LAYER M1 ;
        RECT 23.2 9.456 23.232 11.964 ;
  LAYER M1 ;
        RECT 23.136 9.456 23.168 11.964 ;
  LAYER M1 ;
        RECT 23.072 9.456 23.104 11.964 ;
  LAYER M1 ;
        RECT 23.008 9.456 23.04 11.964 ;
  LAYER M1 ;
        RECT 22.944 9.456 22.976 11.964 ;
  LAYER M1 ;
        RECT 22.88 9.456 22.912 11.964 ;
  LAYER M1 ;
        RECT 22.816 9.456 22.848 11.964 ;
  LAYER M1 ;
        RECT 22.752 9.456 22.784 11.964 ;
  LAYER M1 ;
        RECT 22.688 9.456 22.72 11.964 ;
  LAYER M1 ;
        RECT 22.624 9.456 22.656 11.964 ;
  LAYER M1 ;
        RECT 22.56 9.456 22.592 11.964 ;
  LAYER M1 ;
        RECT 22.496 9.456 22.528 11.964 ;
  LAYER M1 ;
        RECT 22.432 9.456 22.464 11.964 ;
  LAYER M1 ;
        RECT 22.368 9.456 22.4 11.964 ;
  LAYER M1 ;
        RECT 22.304 9.456 22.336 11.964 ;
  LAYER M1 ;
        RECT 22.24 9.456 22.272 11.964 ;
  LAYER M1 ;
        RECT 22.176 9.456 22.208 11.964 ;
  LAYER M1 ;
        RECT 22.112 9.456 22.144 11.964 ;
  LAYER M1 ;
        RECT 22.048 9.456 22.08 11.964 ;
  LAYER M1 ;
        RECT 21.984 9.456 22.016 11.964 ;
  LAYER M1 ;
        RECT 21.92 9.456 21.952 11.964 ;
  LAYER M2 ;
        RECT 21.804 11.848 24.276 11.88 ;
  LAYER M2 ;
        RECT 21.804 11.784 24.276 11.816 ;
  LAYER M2 ;
        RECT 21.804 11.72 24.276 11.752 ;
  LAYER M2 ;
        RECT 21.804 11.656 24.276 11.688 ;
  LAYER M2 ;
        RECT 21.804 11.592 24.276 11.624 ;
  LAYER M2 ;
        RECT 21.804 11.528 24.276 11.56 ;
  LAYER M2 ;
        RECT 21.804 11.464 24.276 11.496 ;
  LAYER M2 ;
        RECT 21.804 11.4 24.276 11.432 ;
  LAYER M2 ;
        RECT 21.804 11.336 24.276 11.368 ;
  LAYER M2 ;
        RECT 21.804 11.272 24.276 11.304 ;
  LAYER M2 ;
        RECT 21.804 11.208 24.276 11.24 ;
  LAYER M2 ;
        RECT 21.804 11.144 24.276 11.176 ;
  LAYER M2 ;
        RECT 21.804 11.08 24.276 11.112 ;
  LAYER M2 ;
        RECT 21.804 11.016 24.276 11.048 ;
  LAYER M2 ;
        RECT 21.804 10.952 24.276 10.984 ;
  LAYER M2 ;
        RECT 21.804 10.888 24.276 10.92 ;
  LAYER M2 ;
        RECT 21.804 10.824 24.276 10.856 ;
  LAYER M2 ;
        RECT 21.804 10.76 24.276 10.792 ;
  LAYER M2 ;
        RECT 21.804 10.696 24.276 10.728 ;
  LAYER M2 ;
        RECT 21.804 10.632 24.276 10.664 ;
  LAYER M2 ;
        RECT 21.804 10.568 24.276 10.6 ;
  LAYER M2 ;
        RECT 21.804 10.504 24.276 10.536 ;
  LAYER M2 ;
        RECT 21.804 10.44 24.276 10.472 ;
  LAYER M2 ;
        RECT 21.804 10.376 24.276 10.408 ;
  LAYER M2 ;
        RECT 21.804 10.312 24.276 10.344 ;
  LAYER M2 ;
        RECT 21.804 10.248 24.276 10.28 ;
  LAYER M2 ;
        RECT 21.804 10.184 24.276 10.216 ;
  LAYER M2 ;
        RECT 21.804 10.12 24.276 10.152 ;
  LAYER M2 ;
        RECT 21.804 10.056 24.276 10.088 ;
  LAYER M2 ;
        RECT 21.804 9.992 24.276 10.024 ;
  LAYER M2 ;
        RECT 21.804 9.928 24.276 9.96 ;
  LAYER M2 ;
        RECT 21.804 9.864 24.276 9.896 ;
  LAYER M2 ;
        RECT 21.804 9.8 24.276 9.832 ;
  LAYER M2 ;
        RECT 21.804 9.736 24.276 9.768 ;
  LAYER M2 ;
        RECT 21.804 9.672 24.276 9.704 ;
  LAYER M2 ;
        RECT 21.804 9.608 24.276 9.64 ;
  LAYER M3 ;
        RECT 24.224 9.456 24.256 11.964 ;
  LAYER M3 ;
        RECT 24.16 9.456 24.192 11.964 ;
  LAYER M3 ;
        RECT 24.096 9.456 24.128 11.964 ;
  LAYER M3 ;
        RECT 24.032 9.456 24.064 11.964 ;
  LAYER M3 ;
        RECT 23.968 9.456 24 11.964 ;
  LAYER M3 ;
        RECT 23.904 9.456 23.936 11.964 ;
  LAYER M3 ;
        RECT 23.84 9.456 23.872 11.964 ;
  LAYER M3 ;
        RECT 23.776 9.456 23.808 11.964 ;
  LAYER M3 ;
        RECT 23.712 9.456 23.744 11.964 ;
  LAYER M3 ;
        RECT 23.648 9.456 23.68 11.964 ;
  LAYER M3 ;
        RECT 23.584 9.456 23.616 11.964 ;
  LAYER M3 ;
        RECT 23.52 9.456 23.552 11.964 ;
  LAYER M3 ;
        RECT 23.456 9.456 23.488 11.964 ;
  LAYER M3 ;
        RECT 23.392 9.456 23.424 11.964 ;
  LAYER M3 ;
        RECT 23.328 9.456 23.36 11.964 ;
  LAYER M3 ;
        RECT 23.264 9.456 23.296 11.964 ;
  LAYER M3 ;
        RECT 23.2 9.456 23.232 11.964 ;
  LAYER M3 ;
        RECT 23.136 9.456 23.168 11.964 ;
  LAYER M3 ;
        RECT 23.072 9.456 23.104 11.964 ;
  LAYER M3 ;
        RECT 23.008 9.456 23.04 11.964 ;
  LAYER M3 ;
        RECT 22.944 9.456 22.976 11.964 ;
  LAYER M3 ;
        RECT 22.88 9.456 22.912 11.964 ;
  LAYER M3 ;
        RECT 22.816 9.456 22.848 11.964 ;
  LAYER M3 ;
        RECT 22.752 9.456 22.784 11.964 ;
  LAYER M3 ;
        RECT 22.688 9.456 22.72 11.964 ;
  LAYER M3 ;
        RECT 22.624 9.456 22.656 11.964 ;
  LAYER M3 ;
        RECT 22.56 9.456 22.592 11.964 ;
  LAYER M3 ;
        RECT 22.496 9.456 22.528 11.964 ;
  LAYER M3 ;
        RECT 22.432 9.456 22.464 11.964 ;
  LAYER M3 ;
        RECT 22.368 9.456 22.4 11.964 ;
  LAYER M3 ;
        RECT 22.304 9.456 22.336 11.964 ;
  LAYER M3 ;
        RECT 22.24 9.456 22.272 11.964 ;
  LAYER M3 ;
        RECT 22.176 9.456 22.208 11.964 ;
  LAYER M3 ;
        RECT 22.112 9.456 22.144 11.964 ;
  LAYER M3 ;
        RECT 22.048 9.456 22.08 11.964 ;
  LAYER M3 ;
        RECT 21.984 9.456 22.016 11.964 ;
  LAYER M3 ;
        RECT 21.92 9.456 21.952 11.964 ;
  LAYER M3 ;
        RECT 21.824 9.456 21.856 11.964 ;
  LAYER M1 ;
        RECT 24.239 9.492 24.241 11.928 ;
  LAYER M1 ;
        RECT 24.159 9.492 24.161 11.928 ;
  LAYER M1 ;
        RECT 24.079 9.492 24.081 11.928 ;
  LAYER M1 ;
        RECT 23.999 9.492 24.001 11.928 ;
  LAYER M1 ;
        RECT 23.919 9.492 23.921 11.928 ;
  LAYER M1 ;
        RECT 23.839 9.492 23.841 11.928 ;
  LAYER M1 ;
        RECT 23.759 9.492 23.761 11.928 ;
  LAYER M1 ;
        RECT 23.679 9.492 23.681 11.928 ;
  LAYER M1 ;
        RECT 23.599 9.492 23.601 11.928 ;
  LAYER M1 ;
        RECT 23.519 9.492 23.521 11.928 ;
  LAYER M1 ;
        RECT 23.439 9.492 23.441 11.928 ;
  LAYER M1 ;
        RECT 23.359 9.492 23.361 11.928 ;
  LAYER M1 ;
        RECT 23.279 9.492 23.281 11.928 ;
  LAYER M1 ;
        RECT 23.199 9.492 23.201 11.928 ;
  LAYER M1 ;
        RECT 23.119 9.492 23.121 11.928 ;
  LAYER M1 ;
        RECT 23.039 9.492 23.041 11.928 ;
  LAYER M1 ;
        RECT 22.959 9.492 22.961 11.928 ;
  LAYER M1 ;
        RECT 22.879 9.492 22.881 11.928 ;
  LAYER M1 ;
        RECT 22.799 9.492 22.801 11.928 ;
  LAYER M1 ;
        RECT 22.719 9.492 22.721 11.928 ;
  LAYER M1 ;
        RECT 22.639 9.492 22.641 11.928 ;
  LAYER M1 ;
        RECT 22.559 9.492 22.561 11.928 ;
  LAYER M1 ;
        RECT 22.479 9.492 22.481 11.928 ;
  LAYER M1 ;
        RECT 22.399 9.492 22.401 11.928 ;
  LAYER M1 ;
        RECT 22.319 9.492 22.321 11.928 ;
  LAYER M1 ;
        RECT 22.239 9.492 22.241 11.928 ;
  LAYER M1 ;
        RECT 22.159 9.492 22.161 11.928 ;
  LAYER M1 ;
        RECT 22.079 9.492 22.081 11.928 ;
  LAYER M1 ;
        RECT 21.999 9.492 22.001 11.928 ;
  LAYER M1 ;
        RECT 21.919 9.492 21.921 11.928 ;
  LAYER M2 ;
        RECT 21.84 11.927 24.24 11.929 ;
  LAYER M2 ;
        RECT 21.84 11.843 24.24 11.845 ;
  LAYER M2 ;
        RECT 21.84 11.759 24.24 11.761 ;
  LAYER M2 ;
        RECT 21.84 11.675 24.24 11.677 ;
  LAYER M2 ;
        RECT 21.84 11.591 24.24 11.593 ;
  LAYER M2 ;
        RECT 21.84 11.507 24.24 11.509 ;
  LAYER M2 ;
        RECT 21.84 11.423 24.24 11.425 ;
  LAYER M2 ;
        RECT 21.84 11.339 24.24 11.341 ;
  LAYER M2 ;
        RECT 21.84 11.255 24.24 11.257 ;
  LAYER M2 ;
        RECT 21.84 11.171 24.24 11.173 ;
  LAYER M2 ;
        RECT 21.84 11.087 24.24 11.089 ;
  LAYER M2 ;
        RECT 21.84 11.003 24.24 11.005 ;
  LAYER M2 ;
        RECT 21.84 10.9195 24.24 10.9215 ;
  LAYER M2 ;
        RECT 21.84 10.835 24.24 10.837 ;
  LAYER M2 ;
        RECT 21.84 10.751 24.24 10.753 ;
  LAYER M2 ;
        RECT 21.84 10.667 24.24 10.669 ;
  LAYER M2 ;
        RECT 21.84 10.583 24.24 10.585 ;
  LAYER M2 ;
        RECT 21.84 10.499 24.24 10.501 ;
  LAYER M2 ;
        RECT 21.84 10.415 24.24 10.417 ;
  LAYER M2 ;
        RECT 21.84 10.331 24.24 10.333 ;
  LAYER M2 ;
        RECT 21.84 10.247 24.24 10.249 ;
  LAYER M2 ;
        RECT 21.84 10.163 24.24 10.165 ;
  LAYER M2 ;
        RECT 21.84 10.079 24.24 10.081 ;
  LAYER M2 ;
        RECT 21.84 9.995 24.24 9.997 ;
  LAYER M2 ;
        RECT 21.84 9.911 24.24 9.913 ;
  LAYER M2 ;
        RECT 21.84 9.827 24.24 9.829 ;
  LAYER M2 ;
        RECT 21.84 9.743 24.24 9.745 ;
  LAYER M2 ;
        RECT 21.84 9.659 24.24 9.661 ;
  LAYER M2 ;
        RECT 21.84 9.575 24.24 9.577 ;
  LAYER M1 ;
        RECT 24.224 6.516 24.256 9.024 ;
  LAYER M1 ;
        RECT 24.16 6.516 24.192 9.024 ;
  LAYER M1 ;
        RECT 24.096 6.516 24.128 9.024 ;
  LAYER M1 ;
        RECT 24.032 6.516 24.064 9.024 ;
  LAYER M1 ;
        RECT 23.968 6.516 24 9.024 ;
  LAYER M1 ;
        RECT 23.904 6.516 23.936 9.024 ;
  LAYER M1 ;
        RECT 23.84 6.516 23.872 9.024 ;
  LAYER M1 ;
        RECT 23.776 6.516 23.808 9.024 ;
  LAYER M1 ;
        RECT 23.712 6.516 23.744 9.024 ;
  LAYER M1 ;
        RECT 23.648 6.516 23.68 9.024 ;
  LAYER M1 ;
        RECT 23.584 6.516 23.616 9.024 ;
  LAYER M1 ;
        RECT 23.52 6.516 23.552 9.024 ;
  LAYER M1 ;
        RECT 23.456 6.516 23.488 9.024 ;
  LAYER M1 ;
        RECT 23.392 6.516 23.424 9.024 ;
  LAYER M1 ;
        RECT 23.328 6.516 23.36 9.024 ;
  LAYER M1 ;
        RECT 23.264 6.516 23.296 9.024 ;
  LAYER M1 ;
        RECT 23.2 6.516 23.232 9.024 ;
  LAYER M1 ;
        RECT 23.136 6.516 23.168 9.024 ;
  LAYER M1 ;
        RECT 23.072 6.516 23.104 9.024 ;
  LAYER M1 ;
        RECT 23.008 6.516 23.04 9.024 ;
  LAYER M1 ;
        RECT 22.944 6.516 22.976 9.024 ;
  LAYER M1 ;
        RECT 22.88 6.516 22.912 9.024 ;
  LAYER M1 ;
        RECT 22.816 6.516 22.848 9.024 ;
  LAYER M1 ;
        RECT 22.752 6.516 22.784 9.024 ;
  LAYER M1 ;
        RECT 22.688 6.516 22.72 9.024 ;
  LAYER M1 ;
        RECT 22.624 6.516 22.656 9.024 ;
  LAYER M1 ;
        RECT 22.56 6.516 22.592 9.024 ;
  LAYER M1 ;
        RECT 22.496 6.516 22.528 9.024 ;
  LAYER M1 ;
        RECT 22.432 6.516 22.464 9.024 ;
  LAYER M1 ;
        RECT 22.368 6.516 22.4 9.024 ;
  LAYER M1 ;
        RECT 22.304 6.516 22.336 9.024 ;
  LAYER M1 ;
        RECT 22.24 6.516 22.272 9.024 ;
  LAYER M1 ;
        RECT 22.176 6.516 22.208 9.024 ;
  LAYER M1 ;
        RECT 22.112 6.516 22.144 9.024 ;
  LAYER M1 ;
        RECT 22.048 6.516 22.08 9.024 ;
  LAYER M1 ;
        RECT 21.984 6.516 22.016 9.024 ;
  LAYER M1 ;
        RECT 21.92 6.516 21.952 9.024 ;
  LAYER M2 ;
        RECT 21.804 8.908 24.276 8.94 ;
  LAYER M2 ;
        RECT 21.804 8.844 24.276 8.876 ;
  LAYER M2 ;
        RECT 21.804 8.78 24.276 8.812 ;
  LAYER M2 ;
        RECT 21.804 8.716 24.276 8.748 ;
  LAYER M2 ;
        RECT 21.804 8.652 24.276 8.684 ;
  LAYER M2 ;
        RECT 21.804 8.588 24.276 8.62 ;
  LAYER M2 ;
        RECT 21.804 8.524 24.276 8.556 ;
  LAYER M2 ;
        RECT 21.804 8.46 24.276 8.492 ;
  LAYER M2 ;
        RECT 21.804 8.396 24.276 8.428 ;
  LAYER M2 ;
        RECT 21.804 8.332 24.276 8.364 ;
  LAYER M2 ;
        RECT 21.804 8.268 24.276 8.3 ;
  LAYER M2 ;
        RECT 21.804 8.204 24.276 8.236 ;
  LAYER M2 ;
        RECT 21.804 8.14 24.276 8.172 ;
  LAYER M2 ;
        RECT 21.804 8.076 24.276 8.108 ;
  LAYER M2 ;
        RECT 21.804 8.012 24.276 8.044 ;
  LAYER M2 ;
        RECT 21.804 7.948 24.276 7.98 ;
  LAYER M2 ;
        RECT 21.804 7.884 24.276 7.916 ;
  LAYER M2 ;
        RECT 21.804 7.82 24.276 7.852 ;
  LAYER M2 ;
        RECT 21.804 7.756 24.276 7.788 ;
  LAYER M2 ;
        RECT 21.804 7.692 24.276 7.724 ;
  LAYER M2 ;
        RECT 21.804 7.628 24.276 7.66 ;
  LAYER M2 ;
        RECT 21.804 7.564 24.276 7.596 ;
  LAYER M2 ;
        RECT 21.804 7.5 24.276 7.532 ;
  LAYER M2 ;
        RECT 21.804 7.436 24.276 7.468 ;
  LAYER M2 ;
        RECT 21.804 7.372 24.276 7.404 ;
  LAYER M2 ;
        RECT 21.804 7.308 24.276 7.34 ;
  LAYER M2 ;
        RECT 21.804 7.244 24.276 7.276 ;
  LAYER M2 ;
        RECT 21.804 7.18 24.276 7.212 ;
  LAYER M2 ;
        RECT 21.804 7.116 24.276 7.148 ;
  LAYER M2 ;
        RECT 21.804 7.052 24.276 7.084 ;
  LAYER M2 ;
        RECT 21.804 6.988 24.276 7.02 ;
  LAYER M2 ;
        RECT 21.804 6.924 24.276 6.956 ;
  LAYER M2 ;
        RECT 21.804 6.86 24.276 6.892 ;
  LAYER M2 ;
        RECT 21.804 6.796 24.276 6.828 ;
  LAYER M2 ;
        RECT 21.804 6.732 24.276 6.764 ;
  LAYER M2 ;
        RECT 21.804 6.668 24.276 6.7 ;
  LAYER M3 ;
        RECT 24.224 6.516 24.256 9.024 ;
  LAYER M3 ;
        RECT 24.16 6.516 24.192 9.024 ;
  LAYER M3 ;
        RECT 24.096 6.516 24.128 9.024 ;
  LAYER M3 ;
        RECT 24.032 6.516 24.064 9.024 ;
  LAYER M3 ;
        RECT 23.968 6.516 24 9.024 ;
  LAYER M3 ;
        RECT 23.904 6.516 23.936 9.024 ;
  LAYER M3 ;
        RECT 23.84 6.516 23.872 9.024 ;
  LAYER M3 ;
        RECT 23.776 6.516 23.808 9.024 ;
  LAYER M3 ;
        RECT 23.712 6.516 23.744 9.024 ;
  LAYER M3 ;
        RECT 23.648 6.516 23.68 9.024 ;
  LAYER M3 ;
        RECT 23.584 6.516 23.616 9.024 ;
  LAYER M3 ;
        RECT 23.52 6.516 23.552 9.024 ;
  LAYER M3 ;
        RECT 23.456 6.516 23.488 9.024 ;
  LAYER M3 ;
        RECT 23.392 6.516 23.424 9.024 ;
  LAYER M3 ;
        RECT 23.328 6.516 23.36 9.024 ;
  LAYER M3 ;
        RECT 23.264 6.516 23.296 9.024 ;
  LAYER M3 ;
        RECT 23.2 6.516 23.232 9.024 ;
  LAYER M3 ;
        RECT 23.136 6.516 23.168 9.024 ;
  LAYER M3 ;
        RECT 23.072 6.516 23.104 9.024 ;
  LAYER M3 ;
        RECT 23.008 6.516 23.04 9.024 ;
  LAYER M3 ;
        RECT 22.944 6.516 22.976 9.024 ;
  LAYER M3 ;
        RECT 22.88 6.516 22.912 9.024 ;
  LAYER M3 ;
        RECT 22.816 6.516 22.848 9.024 ;
  LAYER M3 ;
        RECT 22.752 6.516 22.784 9.024 ;
  LAYER M3 ;
        RECT 22.688 6.516 22.72 9.024 ;
  LAYER M3 ;
        RECT 22.624 6.516 22.656 9.024 ;
  LAYER M3 ;
        RECT 22.56 6.516 22.592 9.024 ;
  LAYER M3 ;
        RECT 22.496 6.516 22.528 9.024 ;
  LAYER M3 ;
        RECT 22.432 6.516 22.464 9.024 ;
  LAYER M3 ;
        RECT 22.368 6.516 22.4 9.024 ;
  LAYER M3 ;
        RECT 22.304 6.516 22.336 9.024 ;
  LAYER M3 ;
        RECT 22.24 6.516 22.272 9.024 ;
  LAYER M3 ;
        RECT 22.176 6.516 22.208 9.024 ;
  LAYER M3 ;
        RECT 22.112 6.516 22.144 9.024 ;
  LAYER M3 ;
        RECT 22.048 6.516 22.08 9.024 ;
  LAYER M3 ;
        RECT 21.984 6.516 22.016 9.024 ;
  LAYER M3 ;
        RECT 21.92 6.516 21.952 9.024 ;
  LAYER M3 ;
        RECT 21.824 6.516 21.856 9.024 ;
  LAYER M1 ;
        RECT 24.239 6.552 24.241 8.988 ;
  LAYER M1 ;
        RECT 24.159 6.552 24.161 8.988 ;
  LAYER M1 ;
        RECT 24.079 6.552 24.081 8.988 ;
  LAYER M1 ;
        RECT 23.999 6.552 24.001 8.988 ;
  LAYER M1 ;
        RECT 23.919 6.552 23.921 8.988 ;
  LAYER M1 ;
        RECT 23.839 6.552 23.841 8.988 ;
  LAYER M1 ;
        RECT 23.759 6.552 23.761 8.988 ;
  LAYER M1 ;
        RECT 23.679 6.552 23.681 8.988 ;
  LAYER M1 ;
        RECT 23.599 6.552 23.601 8.988 ;
  LAYER M1 ;
        RECT 23.519 6.552 23.521 8.988 ;
  LAYER M1 ;
        RECT 23.439 6.552 23.441 8.988 ;
  LAYER M1 ;
        RECT 23.359 6.552 23.361 8.988 ;
  LAYER M1 ;
        RECT 23.279 6.552 23.281 8.988 ;
  LAYER M1 ;
        RECT 23.199 6.552 23.201 8.988 ;
  LAYER M1 ;
        RECT 23.119 6.552 23.121 8.988 ;
  LAYER M1 ;
        RECT 23.039 6.552 23.041 8.988 ;
  LAYER M1 ;
        RECT 22.959 6.552 22.961 8.988 ;
  LAYER M1 ;
        RECT 22.879 6.552 22.881 8.988 ;
  LAYER M1 ;
        RECT 22.799 6.552 22.801 8.988 ;
  LAYER M1 ;
        RECT 22.719 6.552 22.721 8.988 ;
  LAYER M1 ;
        RECT 22.639 6.552 22.641 8.988 ;
  LAYER M1 ;
        RECT 22.559 6.552 22.561 8.988 ;
  LAYER M1 ;
        RECT 22.479 6.552 22.481 8.988 ;
  LAYER M1 ;
        RECT 22.399 6.552 22.401 8.988 ;
  LAYER M1 ;
        RECT 22.319 6.552 22.321 8.988 ;
  LAYER M1 ;
        RECT 22.239 6.552 22.241 8.988 ;
  LAYER M1 ;
        RECT 22.159 6.552 22.161 8.988 ;
  LAYER M1 ;
        RECT 22.079 6.552 22.081 8.988 ;
  LAYER M1 ;
        RECT 21.999 6.552 22.001 8.988 ;
  LAYER M1 ;
        RECT 21.919 6.552 21.921 8.988 ;
  LAYER M2 ;
        RECT 21.84 8.987 24.24 8.989 ;
  LAYER M2 ;
        RECT 21.84 8.903 24.24 8.905 ;
  LAYER M2 ;
        RECT 21.84 8.819 24.24 8.821 ;
  LAYER M2 ;
        RECT 21.84 8.735 24.24 8.737 ;
  LAYER M2 ;
        RECT 21.84 8.651 24.24 8.653 ;
  LAYER M2 ;
        RECT 21.84 8.567 24.24 8.569 ;
  LAYER M2 ;
        RECT 21.84 8.483 24.24 8.485 ;
  LAYER M2 ;
        RECT 21.84 8.399 24.24 8.401 ;
  LAYER M2 ;
        RECT 21.84 8.315 24.24 8.317 ;
  LAYER M2 ;
        RECT 21.84 8.231 24.24 8.233 ;
  LAYER M2 ;
        RECT 21.84 8.147 24.24 8.149 ;
  LAYER M2 ;
        RECT 21.84 8.063 24.24 8.065 ;
  LAYER M2 ;
        RECT 21.84 7.9795 24.24 7.9815 ;
  LAYER M2 ;
        RECT 21.84 7.895 24.24 7.897 ;
  LAYER M2 ;
        RECT 21.84 7.811 24.24 7.813 ;
  LAYER M2 ;
        RECT 21.84 7.727 24.24 7.729 ;
  LAYER M2 ;
        RECT 21.84 7.643 24.24 7.645 ;
  LAYER M2 ;
        RECT 21.84 7.559 24.24 7.561 ;
  LAYER M2 ;
        RECT 21.84 7.475 24.24 7.477 ;
  LAYER M2 ;
        RECT 21.84 7.391 24.24 7.393 ;
  LAYER M2 ;
        RECT 21.84 7.307 24.24 7.309 ;
  LAYER M2 ;
        RECT 21.84 7.223 24.24 7.225 ;
  LAYER M2 ;
        RECT 21.84 7.139 24.24 7.141 ;
  LAYER M2 ;
        RECT 21.84 7.055 24.24 7.057 ;
  LAYER M2 ;
        RECT 21.84 6.971 24.24 6.973 ;
  LAYER M2 ;
        RECT 21.84 6.887 24.24 6.889 ;
  LAYER M2 ;
        RECT 21.84 6.803 24.24 6.805 ;
  LAYER M2 ;
        RECT 21.84 6.719 24.24 6.721 ;
  LAYER M2 ;
        RECT 21.84 6.635 24.24 6.637 ;
  LAYER M1 ;
        RECT 21.344 15.336 21.376 17.844 ;
  LAYER M1 ;
        RECT 21.28 15.336 21.312 17.844 ;
  LAYER M1 ;
        RECT 21.216 15.336 21.248 17.844 ;
  LAYER M1 ;
        RECT 21.152 15.336 21.184 17.844 ;
  LAYER M1 ;
        RECT 21.088 15.336 21.12 17.844 ;
  LAYER M1 ;
        RECT 21.024 15.336 21.056 17.844 ;
  LAYER M1 ;
        RECT 20.96 15.336 20.992 17.844 ;
  LAYER M1 ;
        RECT 20.896 15.336 20.928 17.844 ;
  LAYER M1 ;
        RECT 20.832 15.336 20.864 17.844 ;
  LAYER M1 ;
        RECT 20.768 15.336 20.8 17.844 ;
  LAYER M1 ;
        RECT 20.704 15.336 20.736 17.844 ;
  LAYER M1 ;
        RECT 20.64 15.336 20.672 17.844 ;
  LAYER M1 ;
        RECT 20.576 15.336 20.608 17.844 ;
  LAYER M1 ;
        RECT 20.512 15.336 20.544 17.844 ;
  LAYER M1 ;
        RECT 20.448 15.336 20.48 17.844 ;
  LAYER M1 ;
        RECT 20.384 15.336 20.416 17.844 ;
  LAYER M1 ;
        RECT 20.32 15.336 20.352 17.844 ;
  LAYER M1 ;
        RECT 20.256 15.336 20.288 17.844 ;
  LAYER M1 ;
        RECT 20.192 15.336 20.224 17.844 ;
  LAYER M1 ;
        RECT 20.128 15.336 20.16 17.844 ;
  LAYER M1 ;
        RECT 20.064 15.336 20.096 17.844 ;
  LAYER M1 ;
        RECT 20 15.336 20.032 17.844 ;
  LAYER M1 ;
        RECT 19.936 15.336 19.968 17.844 ;
  LAYER M1 ;
        RECT 19.872 15.336 19.904 17.844 ;
  LAYER M1 ;
        RECT 19.808 15.336 19.84 17.844 ;
  LAYER M1 ;
        RECT 19.744 15.336 19.776 17.844 ;
  LAYER M1 ;
        RECT 19.68 15.336 19.712 17.844 ;
  LAYER M1 ;
        RECT 19.616 15.336 19.648 17.844 ;
  LAYER M1 ;
        RECT 19.552 15.336 19.584 17.844 ;
  LAYER M1 ;
        RECT 19.488 15.336 19.52 17.844 ;
  LAYER M1 ;
        RECT 19.424 15.336 19.456 17.844 ;
  LAYER M1 ;
        RECT 19.36 15.336 19.392 17.844 ;
  LAYER M1 ;
        RECT 19.296 15.336 19.328 17.844 ;
  LAYER M1 ;
        RECT 19.232 15.336 19.264 17.844 ;
  LAYER M1 ;
        RECT 19.168 15.336 19.2 17.844 ;
  LAYER M1 ;
        RECT 19.104 15.336 19.136 17.844 ;
  LAYER M1 ;
        RECT 19.04 15.336 19.072 17.844 ;
  LAYER M2 ;
        RECT 18.924 17.728 21.396 17.76 ;
  LAYER M2 ;
        RECT 18.924 17.664 21.396 17.696 ;
  LAYER M2 ;
        RECT 18.924 17.6 21.396 17.632 ;
  LAYER M2 ;
        RECT 18.924 17.536 21.396 17.568 ;
  LAYER M2 ;
        RECT 18.924 17.472 21.396 17.504 ;
  LAYER M2 ;
        RECT 18.924 17.408 21.396 17.44 ;
  LAYER M2 ;
        RECT 18.924 17.344 21.396 17.376 ;
  LAYER M2 ;
        RECT 18.924 17.28 21.396 17.312 ;
  LAYER M2 ;
        RECT 18.924 17.216 21.396 17.248 ;
  LAYER M2 ;
        RECT 18.924 17.152 21.396 17.184 ;
  LAYER M2 ;
        RECT 18.924 17.088 21.396 17.12 ;
  LAYER M2 ;
        RECT 18.924 17.024 21.396 17.056 ;
  LAYER M2 ;
        RECT 18.924 16.96 21.396 16.992 ;
  LAYER M2 ;
        RECT 18.924 16.896 21.396 16.928 ;
  LAYER M2 ;
        RECT 18.924 16.832 21.396 16.864 ;
  LAYER M2 ;
        RECT 18.924 16.768 21.396 16.8 ;
  LAYER M2 ;
        RECT 18.924 16.704 21.396 16.736 ;
  LAYER M2 ;
        RECT 18.924 16.64 21.396 16.672 ;
  LAYER M2 ;
        RECT 18.924 16.576 21.396 16.608 ;
  LAYER M2 ;
        RECT 18.924 16.512 21.396 16.544 ;
  LAYER M2 ;
        RECT 18.924 16.448 21.396 16.48 ;
  LAYER M2 ;
        RECT 18.924 16.384 21.396 16.416 ;
  LAYER M2 ;
        RECT 18.924 16.32 21.396 16.352 ;
  LAYER M2 ;
        RECT 18.924 16.256 21.396 16.288 ;
  LAYER M2 ;
        RECT 18.924 16.192 21.396 16.224 ;
  LAYER M2 ;
        RECT 18.924 16.128 21.396 16.16 ;
  LAYER M2 ;
        RECT 18.924 16.064 21.396 16.096 ;
  LAYER M2 ;
        RECT 18.924 16 21.396 16.032 ;
  LAYER M2 ;
        RECT 18.924 15.936 21.396 15.968 ;
  LAYER M2 ;
        RECT 18.924 15.872 21.396 15.904 ;
  LAYER M2 ;
        RECT 18.924 15.808 21.396 15.84 ;
  LAYER M2 ;
        RECT 18.924 15.744 21.396 15.776 ;
  LAYER M2 ;
        RECT 18.924 15.68 21.396 15.712 ;
  LAYER M2 ;
        RECT 18.924 15.616 21.396 15.648 ;
  LAYER M2 ;
        RECT 18.924 15.552 21.396 15.584 ;
  LAYER M2 ;
        RECT 18.924 15.488 21.396 15.52 ;
  LAYER M3 ;
        RECT 21.344 15.336 21.376 17.844 ;
  LAYER M3 ;
        RECT 21.28 15.336 21.312 17.844 ;
  LAYER M3 ;
        RECT 21.216 15.336 21.248 17.844 ;
  LAYER M3 ;
        RECT 21.152 15.336 21.184 17.844 ;
  LAYER M3 ;
        RECT 21.088 15.336 21.12 17.844 ;
  LAYER M3 ;
        RECT 21.024 15.336 21.056 17.844 ;
  LAYER M3 ;
        RECT 20.96 15.336 20.992 17.844 ;
  LAYER M3 ;
        RECT 20.896 15.336 20.928 17.844 ;
  LAYER M3 ;
        RECT 20.832 15.336 20.864 17.844 ;
  LAYER M3 ;
        RECT 20.768 15.336 20.8 17.844 ;
  LAYER M3 ;
        RECT 20.704 15.336 20.736 17.844 ;
  LAYER M3 ;
        RECT 20.64 15.336 20.672 17.844 ;
  LAYER M3 ;
        RECT 20.576 15.336 20.608 17.844 ;
  LAYER M3 ;
        RECT 20.512 15.336 20.544 17.844 ;
  LAYER M3 ;
        RECT 20.448 15.336 20.48 17.844 ;
  LAYER M3 ;
        RECT 20.384 15.336 20.416 17.844 ;
  LAYER M3 ;
        RECT 20.32 15.336 20.352 17.844 ;
  LAYER M3 ;
        RECT 20.256 15.336 20.288 17.844 ;
  LAYER M3 ;
        RECT 20.192 15.336 20.224 17.844 ;
  LAYER M3 ;
        RECT 20.128 15.336 20.16 17.844 ;
  LAYER M3 ;
        RECT 20.064 15.336 20.096 17.844 ;
  LAYER M3 ;
        RECT 20 15.336 20.032 17.844 ;
  LAYER M3 ;
        RECT 19.936 15.336 19.968 17.844 ;
  LAYER M3 ;
        RECT 19.872 15.336 19.904 17.844 ;
  LAYER M3 ;
        RECT 19.808 15.336 19.84 17.844 ;
  LAYER M3 ;
        RECT 19.744 15.336 19.776 17.844 ;
  LAYER M3 ;
        RECT 19.68 15.336 19.712 17.844 ;
  LAYER M3 ;
        RECT 19.616 15.336 19.648 17.844 ;
  LAYER M3 ;
        RECT 19.552 15.336 19.584 17.844 ;
  LAYER M3 ;
        RECT 19.488 15.336 19.52 17.844 ;
  LAYER M3 ;
        RECT 19.424 15.336 19.456 17.844 ;
  LAYER M3 ;
        RECT 19.36 15.336 19.392 17.844 ;
  LAYER M3 ;
        RECT 19.296 15.336 19.328 17.844 ;
  LAYER M3 ;
        RECT 19.232 15.336 19.264 17.844 ;
  LAYER M3 ;
        RECT 19.168 15.336 19.2 17.844 ;
  LAYER M3 ;
        RECT 19.104 15.336 19.136 17.844 ;
  LAYER M3 ;
        RECT 19.04 15.336 19.072 17.844 ;
  LAYER M3 ;
        RECT 18.944 15.336 18.976 17.844 ;
  LAYER M1 ;
        RECT 21.359 15.372 21.361 17.808 ;
  LAYER M1 ;
        RECT 21.279 15.372 21.281 17.808 ;
  LAYER M1 ;
        RECT 21.199 15.372 21.201 17.808 ;
  LAYER M1 ;
        RECT 21.119 15.372 21.121 17.808 ;
  LAYER M1 ;
        RECT 21.039 15.372 21.041 17.808 ;
  LAYER M1 ;
        RECT 20.959 15.372 20.961 17.808 ;
  LAYER M1 ;
        RECT 20.879 15.372 20.881 17.808 ;
  LAYER M1 ;
        RECT 20.799 15.372 20.801 17.808 ;
  LAYER M1 ;
        RECT 20.719 15.372 20.721 17.808 ;
  LAYER M1 ;
        RECT 20.639 15.372 20.641 17.808 ;
  LAYER M1 ;
        RECT 20.559 15.372 20.561 17.808 ;
  LAYER M1 ;
        RECT 20.479 15.372 20.481 17.808 ;
  LAYER M1 ;
        RECT 20.399 15.372 20.401 17.808 ;
  LAYER M1 ;
        RECT 20.319 15.372 20.321 17.808 ;
  LAYER M1 ;
        RECT 20.239 15.372 20.241 17.808 ;
  LAYER M1 ;
        RECT 20.159 15.372 20.161 17.808 ;
  LAYER M1 ;
        RECT 20.079 15.372 20.081 17.808 ;
  LAYER M1 ;
        RECT 19.999 15.372 20.001 17.808 ;
  LAYER M1 ;
        RECT 19.919 15.372 19.921 17.808 ;
  LAYER M1 ;
        RECT 19.839 15.372 19.841 17.808 ;
  LAYER M1 ;
        RECT 19.759 15.372 19.761 17.808 ;
  LAYER M1 ;
        RECT 19.679 15.372 19.681 17.808 ;
  LAYER M1 ;
        RECT 19.599 15.372 19.601 17.808 ;
  LAYER M1 ;
        RECT 19.519 15.372 19.521 17.808 ;
  LAYER M1 ;
        RECT 19.439 15.372 19.441 17.808 ;
  LAYER M1 ;
        RECT 19.359 15.372 19.361 17.808 ;
  LAYER M1 ;
        RECT 19.279 15.372 19.281 17.808 ;
  LAYER M1 ;
        RECT 19.199 15.372 19.201 17.808 ;
  LAYER M1 ;
        RECT 19.119 15.372 19.121 17.808 ;
  LAYER M1 ;
        RECT 19.039 15.372 19.041 17.808 ;
  LAYER M2 ;
        RECT 18.96 17.807 21.36 17.809 ;
  LAYER M2 ;
        RECT 18.96 17.723 21.36 17.725 ;
  LAYER M2 ;
        RECT 18.96 17.639 21.36 17.641 ;
  LAYER M2 ;
        RECT 18.96 17.555 21.36 17.557 ;
  LAYER M2 ;
        RECT 18.96 17.471 21.36 17.473 ;
  LAYER M2 ;
        RECT 18.96 17.387 21.36 17.389 ;
  LAYER M2 ;
        RECT 18.96 17.303 21.36 17.305 ;
  LAYER M2 ;
        RECT 18.96 17.219 21.36 17.221 ;
  LAYER M2 ;
        RECT 18.96 17.135 21.36 17.137 ;
  LAYER M2 ;
        RECT 18.96 17.051 21.36 17.053 ;
  LAYER M2 ;
        RECT 18.96 16.967 21.36 16.969 ;
  LAYER M2 ;
        RECT 18.96 16.883 21.36 16.885 ;
  LAYER M2 ;
        RECT 18.96 16.7995 21.36 16.8015 ;
  LAYER M2 ;
        RECT 18.96 16.715 21.36 16.717 ;
  LAYER M2 ;
        RECT 18.96 16.631 21.36 16.633 ;
  LAYER M2 ;
        RECT 18.96 16.547 21.36 16.549 ;
  LAYER M2 ;
        RECT 18.96 16.463 21.36 16.465 ;
  LAYER M2 ;
        RECT 18.96 16.379 21.36 16.381 ;
  LAYER M2 ;
        RECT 18.96 16.295 21.36 16.297 ;
  LAYER M2 ;
        RECT 18.96 16.211 21.36 16.213 ;
  LAYER M2 ;
        RECT 18.96 16.127 21.36 16.129 ;
  LAYER M2 ;
        RECT 18.96 16.043 21.36 16.045 ;
  LAYER M2 ;
        RECT 18.96 15.959 21.36 15.961 ;
  LAYER M2 ;
        RECT 18.96 15.875 21.36 15.877 ;
  LAYER M2 ;
        RECT 18.96 15.791 21.36 15.793 ;
  LAYER M2 ;
        RECT 18.96 15.707 21.36 15.709 ;
  LAYER M2 ;
        RECT 18.96 15.623 21.36 15.625 ;
  LAYER M2 ;
        RECT 18.96 15.539 21.36 15.541 ;
  LAYER M2 ;
        RECT 18.96 15.455 21.36 15.457 ;
  LAYER M1 ;
        RECT 21.344 12.396 21.376 14.904 ;
  LAYER M1 ;
        RECT 21.28 12.396 21.312 14.904 ;
  LAYER M1 ;
        RECT 21.216 12.396 21.248 14.904 ;
  LAYER M1 ;
        RECT 21.152 12.396 21.184 14.904 ;
  LAYER M1 ;
        RECT 21.088 12.396 21.12 14.904 ;
  LAYER M1 ;
        RECT 21.024 12.396 21.056 14.904 ;
  LAYER M1 ;
        RECT 20.96 12.396 20.992 14.904 ;
  LAYER M1 ;
        RECT 20.896 12.396 20.928 14.904 ;
  LAYER M1 ;
        RECT 20.832 12.396 20.864 14.904 ;
  LAYER M1 ;
        RECT 20.768 12.396 20.8 14.904 ;
  LAYER M1 ;
        RECT 20.704 12.396 20.736 14.904 ;
  LAYER M1 ;
        RECT 20.64 12.396 20.672 14.904 ;
  LAYER M1 ;
        RECT 20.576 12.396 20.608 14.904 ;
  LAYER M1 ;
        RECT 20.512 12.396 20.544 14.904 ;
  LAYER M1 ;
        RECT 20.448 12.396 20.48 14.904 ;
  LAYER M1 ;
        RECT 20.384 12.396 20.416 14.904 ;
  LAYER M1 ;
        RECT 20.32 12.396 20.352 14.904 ;
  LAYER M1 ;
        RECT 20.256 12.396 20.288 14.904 ;
  LAYER M1 ;
        RECT 20.192 12.396 20.224 14.904 ;
  LAYER M1 ;
        RECT 20.128 12.396 20.16 14.904 ;
  LAYER M1 ;
        RECT 20.064 12.396 20.096 14.904 ;
  LAYER M1 ;
        RECT 20 12.396 20.032 14.904 ;
  LAYER M1 ;
        RECT 19.936 12.396 19.968 14.904 ;
  LAYER M1 ;
        RECT 19.872 12.396 19.904 14.904 ;
  LAYER M1 ;
        RECT 19.808 12.396 19.84 14.904 ;
  LAYER M1 ;
        RECT 19.744 12.396 19.776 14.904 ;
  LAYER M1 ;
        RECT 19.68 12.396 19.712 14.904 ;
  LAYER M1 ;
        RECT 19.616 12.396 19.648 14.904 ;
  LAYER M1 ;
        RECT 19.552 12.396 19.584 14.904 ;
  LAYER M1 ;
        RECT 19.488 12.396 19.52 14.904 ;
  LAYER M1 ;
        RECT 19.424 12.396 19.456 14.904 ;
  LAYER M1 ;
        RECT 19.36 12.396 19.392 14.904 ;
  LAYER M1 ;
        RECT 19.296 12.396 19.328 14.904 ;
  LAYER M1 ;
        RECT 19.232 12.396 19.264 14.904 ;
  LAYER M1 ;
        RECT 19.168 12.396 19.2 14.904 ;
  LAYER M1 ;
        RECT 19.104 12.396 19.136 14.904 ;
  LAYER M1 ;
        RECT 19.04 12.396 19.072 14.904 ;
  LAYER M2 ;
        RECT 18.924 14.788 21.396 14.82 ;
  LAYER M2 ;
        RECT 18.924 14.724 21.396 14.756 ;
  LAYER M2 ;
        RECT 18.924 14.66 21.396 14.692 ;
  LAYER M2 ;
        RECT 18.924 14.596 21.396 14.628 ;
  LAYER M2 ;
        RECT 18.924 14.532 21.396 14.564 ;
  LAYER M2 ;
        RECT 18.924 14.468 21.396 14.5 ;
  LAYER M2 ;
        RECT 18.924 14.404 21.396 14.436 ;
  LAYER M2 ;
        RECT 18.924 14.34 21.396 14.372 ;
  LAYER M2 ;
        RECT 18.924 14.276 21.396 14.308 ;
  LAYER M2 ;
        RECT 18.924 14.212 21.396 14.244 ;
  LAYER M2 ;
        RECT 18.924 14.148 21.396 14.18 ;
  LAYER M2 ;
        RECT 18.924 14.084 21.396 14.116 ;
  LAYER M2 ;
        RECT 18.924 14.02 21.396 14.052 ;
  LAYER M2 ;
        RECT 18.924 13.956 21.396 13.988 ;
  LAYER M2 ;
        RECT 18.924 13.892 21.396 13.924 ;
  LAYER M2 ;
        RECT 18.924 13.828 21.396 13.86 ;
  LAYER M2 ;
        RECT 18.924 13.764 21.396 13.796 ;
  LAYER M2 ;
        RECT 18.924 13.7 21.396 13.732 ;
  LAYER M2 ;
        RECT 18.924 13.636 21.396 13.668 ;
  LAYER M2 ;
        RECT 18.924 13.572 21.396 13.604 ;
  LAYER M2 ;
        RECT 18.924 13.508 21.396 13.54 ;
  LAYER M2 ;
        RECT 18.924 13.444 21.396 13.476 ;
  LAYER M2 ;
        RECT 18.924 13.38 21.396 13.412 ;
  LAYER M2 ;
        RECT 18.924 13.316 21.396 13.348 ;
  LAYER M2 ;
        RECT 18.924 13.252 21.396 13.284 ;
  LAYER M2 ;
        RECT 18.924 13.188 21.396 13.22 ;
  LAYER M2 ;
        RECT 18.924 13.124 21.396 13.156 ;
  LAYER M2 ;
        RECT 18.924 13.06 21.396 13.092 ;
  LAYER M2 ;
        RECT 18.924 12.996 21.396 13.028 ;
  LAYER M2 ;
        RECT 18.924 12.932 21.396 12.964 ;
  LAYER M2 ;
        RECT 18.924 12.868 21.396 12.9 ;
  LAYER M2 ;
        RECT 18.924 12.804 21.396 12.836 ;
  LAYER M2 ;
        RECT 18.924 12.74 21.396 12.772 ;
  LAYER M2 ;
        RECT 18.924 12.676 21.396 12.708 ;
  LAYER M2 ;
        RECT 18.924 12.612 21.396 12.644 ;
  LAYER M2 ;
        RECT 18.924 12.548 21.396 12.58 ;
  LAYER M3 ;
        RECT 21.344 12.396 21.376 14.904 ;
  LAYER M3 ;
        RECT 21.28 12.396 21.312 14.904 ;
  LAYER M3 ;
        RECT 21.216 12.396 21.248 14.904 ;
  LAYER M3 ;
        RECT 21.152 12.396 21.184 14.904 ;
  LAYER M3 ;
        RECT 21.088 12.396 21.12 14.904 ;
  LAYER M3 ;
        RECT 21.024 12.396 21.056 14.904 ;
  LAYER M3 ;
        RECT 20.96 12.396 20.992 14.904 ;
  LAYER M3 ;
        RECT 20.896 12.396 20.928 14.904 ;
  LAYER M3 ;
        RECT 20.832 12.396 20.864 14.904 ;
  LAYER M3 ;
        RECT 20.768 12.396 20.8 14.904 ;
  LAYER M3 ;
        RECT 20.704 12.396 20.736 14.904 ;
  LAYER M3 ;
        RECT 20.64 12.396 20.672 14.904 ;
  LAYER M3 ;
        RECT 20.576 12.396 20.608 14.904 ;
  LAYER M3 ;
        RECT 20.512 12.396 20.544 14.904 ;
  LAYER M3 ;
        RECT 20.448 12.396 20.48 14.904 ;
  LAYER M3 ;
        RECT 20.384 12.396 20.416 14.904 ;
  LAYER M3 ;
        RECT 20.32 12.396 20.352 14.904 ;
  LAYER M3 ;
        RECT 20.256 12.396 20.288 14.904 ;
  LAYER M3 ;
        RECT 20.192 12.396 20.224 14.904 ;
  LAYER M3 ;
        RECT 20.128 12.396 20.16 14.904 ;
  LAYER M3 ;
        RECT 20.064 12.396 20.096 14.904 ;
  LAYER M3 ;
        RECT 20 12.396 20.032 14.904 ;
  LAYER M3 ;
        RECT 19.936 12.396 19.968 14.904 ;
  LAYER M3 ;
        RECT 19.872 12.396 19.904 14.904 ;
  LAYER M3 ;
        RECT 19.808 12.396 19.84 14.904 ;
  LAYER M3 ;
        RECT 19.744 12.396 19.776 14.904 ;
  LAYER M3 ;
        RECT 19.68 12.396 19.712 14.904 ;
  LAYER M3 ;
        RECT 19.616 12.396 19.648 14.904 ;
  LAYER M3 ;
        RECT 19.552 12.396 19.584 14.904 ;
  LAYER M3 ;
        RECT 19.488 12.396 19.52 14.904 ;
  LAYER M3 ;
        RECT 19.424 12.396 19.456 14.904 ;
  LAYER M3 ;
        RECT 19.36 12.396 19.392 14.904 ;
  LAYER M3 ;
        RECT 19.296 12.396 19.328 14.904 ;
  LAYER M3 ;
        RECT 19.232 12.396 19.264 14.904 ;
  LAYER M3 ;
        RECT 19.168 12.396 19.2 14.904 ;
  LAYER M3 ;
        RECT 19.104 12.396 19.136 14.904 ;
  LAYER M3 ;
        RECT 19.04 12.396 19.072 14.904 ;
  LAYER M3 ;
        RECT 18.944 12.396 18.976 14.904 ;
  LAYER M1 ;
        RECT 21.359 12.432 21.361 14.868 ;
  LAYER M1 ;
        RECT 21.279 12.432 21.281 14.868 ;
  LAYER M1 ;
        RECT 21.199 12.432 21.201 14.868 ;
  LAYER M1 ;
        RECT 21.119 12.432 21.121 14.868 ;
  LAYER M1 ;
        RECT 21.039 12.432 21.041 14.868 ;
  LAYER M1 ;
        RECT 20.959 12.432 20.961 14.868 ;
  LAYER M1 ;
        RECT 20.879 12.432 20.881 14.868 ;
  LAYER M1 ;
        RECT 20.799 12.432 20.801 14.868 ;
  LAYER M1 ;
        RECT 20.719 12.432 20.721 14.868 ;
  LAYER M1 ;
        RECT 20.639 12.432 20.641 14.868 ;
  LAYER M1 ;
        RECT 20.559 12.432 20.561 14.868 ;
  LAYER M1 ;
        RECT 20.479 12.432 20.481 14.868 ;
  LAYER M1 ;
        RECT 20.399 12.432 20.401 14.868 ;
  LAYER M1 ;
        RECT 20.319 12.432 20.321 14.868 ;
  LAYER M1 ;
        RECT 20.239 12.432 20.241 14.868 ;
  LAYER M1 ;
        RECT 20.159 12.432 20.161 14.868 ;
  LAYER M1 ;
        RECT 20.079 12.432 20.081 14.868 ;
  LAYER M1 ;
        RECT 19.999 12.432 20.001 14.868 ;
  LAYER M1 ;
        RECT 19.919 12.432 19.921 14.868 ;
  LAYER M1 ;
        RECT 19.839 12.432 19.841 14.868 ;
  LAYER M1 ;
        RECT 19.759 12.432 19.761 14.868 ;
  LAYER M1 ;
        RECT 19.679 12.432 19.681 14.868 ;
  LAYER M1 ;
        RECT 19.599 12.432 19.601 14.868 ;
  LAYER M1 ;
        RECT 19.519 12.432 19.521 14.868 ;
  LAYER M1 ;
        RECT 19.439 12.432 19.441 14.868 ;
  LAYER M1 ;
        RECT 19.359 12.432 19.361 14.868 ;
  LAYER M1 ;
        RECT 19.279 12.432 19.281 14.868 ;
  LAYER M1 ;
        RECT 19.199 12.432 19.201 14.868 ;
  LAYER M1 ;
        RECT 19.119 12.432 19.121 14.868 ;
  LAYER M1 ;
        RECT 19.039 12.432 19.041 14.868 ;
  LAYER M2 ;
        RECT 18.96 14.867 21.36 14.869 ;
  LAYER M2 ;
        RECT 18.96 14.783 21.36 14.785 ;
  LAYER M2 ;
        RECT 18.96 14.699 21.36 14.701 ;
  LAYER M2 ;
        RECT 18.96 14.615 21.36 14.617 ;
  LAYER M2 ;
        RECT 18.96 14.531 21.36 14.533 ;
  LAYER M2 ;
        RECT 18.96 14.447 21.36 14.449 ;
  LAYER M2 ;
        RECT 18.96 14.363 21.36 14.365 ;
  LAYER M2 ;
        RECT 18.96 14.279 21.36 14.281 ;
  LAYER M2 ;
        RECT 18.96 14.195 21.36 14.197 ;
  LAYER M2 ;
        RECT 18.96 14.111 21.36 14.113 ;
  LAYER M2 ;
        RECT 18.96 14.027 21.36 14.029 ;
  LAYER M2 ;
        RECT 18.96 13.943 21.36 13.945 ;
  LAYER M2 ;
        RECT 18.96 13.8595 21.36 13.8615 ;
  LAYER M2 ;
        RECT 18.96 13.775 21.36 13.777 ;
  LAYER M2 ;
        RECT 18.96 13.691 21.36 13.693 ;
  LAYER M2 ;
        RECT 18.96 13.607 21.36 13.609 ;
  LAYER M2 ;
        RECT 18.96 13.523 21.36 13.525 ;
  LAYER M2 ;
        RECT 18.96 13.439 21.36 13.441 ;
  LAYER M2 ;
        RECT 18.96 13.355 21.36 13.357 ;
  LAYER M2 ;
        RECT 18.96 13.271 21.36 13.273 ;
  LAYER M2 ;
        RECT 18.96 13.187 21.36 13.189 ;
  LAYER M2 ;
        RECT 18.96 13.103 21.36 13.105 ;
  LAYER M2 ;
        RECT 18.96 13.019 21.36 13.021 ;
  LAYER M2 ;
        RECT 18.96 12.935 21.36 12.937 ;
  LAYER M2 ;
        RECT 18.96 12.851 21.36 12.853 ;
  LAYER M2 ;
        RECT 18.96 12.767 21.36 12.769 ;
  LAYER M2 ;
        RECT 18.96 12.683 21.36 12.685 ;
  LAYER M2 ;
        RECT 18.96 12.599 21.36 12.601 ;
  LAYER M2 ;
        RECT 18.96 12.515 21.36 12.517 ;
  LAYER M1 ;
        RECT 21.344 9.456 21.376 11.964 ;
  LAYER M1 ;
        RECT 21.28 9.456 21.312 11.964 ;
  LAYER M1 ;
        RECT 21.216 9.456 21.248 11.964 ;
  LAYER M1 ;
        RECT 21.152 9.456 21.184 11.964 ;
  LAYER M1 ;
        RECT 21.088 9.456 21.12 11.964 ;
  LAYER M1 ;
        RECT 21.024 9.456 21.056 11.964 ;
  LAYER M1 ;
        RECT 20.96 9.456 20.992 11.964 ;
  LAYER M1 ;
        RECT 20.896 9.456 20.928 11.964 ;
  LAYER M1 ;
        RECT 20.832 9.456 20.864 11.964 ;
  LAYER M1 ;
        RECT 20.768 9.456 20.8 11.964 ;
  LAYER M1 ;
        RECT 20.704 9.456 20.736 11.964 ;
  LAYER M1 ;
        RECT 20.64 9.456 20.672 11.964 ;
  LAYER M1 ;
        RECT 20.576 9.456 20.608 11.964 ;
  LAYER M1 ;
        RECT 20.512 9.456 20.544 11.964 ;
  LAYER M1 ;
        RECT 20.448 9.456 20.48 11.964 ;
  LAYER M1 ;
        RECT 20.384 9.456 20.416 11.964 ;
  LAYER M1 ;
        RECT 20.32 9.456 20.352 11.964 ;
  LAYER M1 ;
        RECT 20.256 9.456 20.288 11.964 ;
  LAYER M1 ;
        RECT 20.192 9.456 20.224 11.964 ;
  LAYER M1 ;
        RECT 20.128 9.456 20.16 11.964 ;
  LAYER M1 ;
        RECT 20.064 9.456 20.096 11.964 ;
  LAYER M1 ;
        RECT 20 9.456 20.032 11.964 ;
  LAYER M1 ;
        RECT 19.936 9.456 19.968 11.964 ;
  LAYER M1 ;
        RECT 19.872 9.456 19.904 11.964 ;
  LAYER M1 ;
        RECT 19.808 9.456 19.84 11.964 ;
  LAYER M1 ;
        RECT 19.744 9.456 19.776 11.964 ;
  LAYER M1 ;
        RECT 19.68 9.456 19.712 11.964 ;
  LAYER M1 ;
        RECT 19.616 9.456 19.648 11.964 ;
  LAYER M1 ;
        RECT 19.552 9.456 19.584 11.964 ;
  LAYER M1 ;
        RECT 19.488 9.456 19.52 11.964 ;
  LAYER M1 ;
        RECT 19.424 9.456 19.456 11.964 ;
  LAYER M1 ;
        RECT 19.36 9.456 19.392 11.964 ;
  LAYER M1 ;
        RECT 19.296 9.456 19.328 11.964 ;
  LAYER M1 ;
        RECT 19.232 9.456 19.264 11.964 ;
  LAYER M1 ;
        RECT 19.168 9.456 19.2 11.964 ;
  LAYER M1 ;
        RECT 19.104 9.456 19.136 11.964 ;
  LAYER M1 ;
        RECT 19.04 9.456 19.072 11.964 ;
  LAYER M2 ;
        RECT 18.924 11.848 21.396 11.88 ;
  LAYER M2 ;
        RECT 18.924 11.784 21.396 11.816 ;
  LAYER M2 ;
        RECT 18.924 11.72 21.396 11.752 ;
  LAYER M2 ;
        RECT 18.924 11.656 21.396 11.688 ;
  LAYER M2 ;
        RECT 18.924 11.592 21.396 11.624 ;
  LAYER M2 ;
        RECT 18.924 11.528 21.396 11.56 ;
  LAYER M2 ;
        RECT 18.924 11.464 21.396 11.496 ;
  LAYER M2 ;
        RECT 18.924 11.4 21.396 11.432 ;
  LAYER M2 ;
        RECT 18.924 11.336 21.396 11.368 ;
  LAYER M2 ;
        RECT 18.924 11.272 21.396 11.304 ;
  LAYER M2 ;
        RECT 18.924 11.208 21.396 11.24 ;
  LAYER M2 ;
        RECT 18.924 11.144 21.396 11.176 ;
  LAYER M2 ;
        RECT 18.924 11.08 21.396 11.112 ;
  LAYER M2 ;
        RECT 18.924 11.016 21.396 11.048 ;
  LAYER M2 ;
        RECT 18.924 10.952 21.396 10.984 ;
  LAYER M2 ;
        RECT 18.924 10.888 21.396 10.92 ;
  LAYER M2 ;
        RECT 18.924 10.824 21.396 10.856 ;
  LAYER M2 ;
        RECT 18.924 10.76 21.396 10.792 ;
  LAYER M2 ;
        RECT 18.924 10.696 21.396 10.728 ;
  LAYER M2 ;
        RECT 18.924 10.632 21.396 10.664 ;
  LAYER M2 ;
        RECT 18.924 10.568 21.396 10.6 ;
  LAYER M2 ;
        RECT 18.924 10.504 21.396 10.536 ;
  LAYER M2 ;
        RECT 18.924 10.44 21.396 10.472 ;
  LAYER M2 ;
        RECT 18.924 10.376 21.396 10.408 ;
  LAYER M2 ;
        RECT 18.924 10.312 21.396 10.344 ;
  LAYER M2 ;
        RECT 18.924 10.248 21.396 10.28 ;
  LAYER M2 ;
        RECT 18.924 10.184 21.396 10.216 ;
  LAYER M2 ;
        RECT 18.924 10.12 21.396 10.152 ;
  LAYER M2 ;
        RECT 18.924 10.056 21.396 10.088 ;
  LAYER M2 ;
        RECT 18.924 9.992 21.396 10.024 ;
  LAYER M2 ;
        RECT 18.924 9.928 21.396 9.96 ;
  LAYER M2 ;
        RECT 18.924 9.864 21.396 9.896 ;
  LAYER M2 ;
        RECT 18.924 9.8 21.396 9.832 ;
  LAYER M2 ;
        RECT 18.924 9.736 21.396 9.768 ;
  LAYER M2 ;
        RECT 18.924 9.672 21.396 9.704 ;
  LAYER M2 ;
        RECT 18.924 9.608 21.396 9.64 ;
  LAYER M3 ;
        RECT 21.344 9.456 21.376 11.964 ;
  LAYER M3 ;
        RECT 21.28 9.456 21.312 11.964 ;
  LAYER M3 ;
        RECT 21.216 9.456 21.248 11.964 ;
  LAYER M3 ;
        RECT 21.152 9.456 21.184 11.964 ;
  LAYER M3 ;
        RECT 21.088 9.456 21.12 11.964 ;
  LAYER M3 ;
        RECT 21.024 9.456 21.056 11.964 ;
  LAYER M3 ;
        RECT 20.96 9.456 20.992 11.964 ;
  LAYER M3 ;
        RECT 20.896 9.456 20.928 11.964 ;
  LAYER M3 ;
        RECT 20.832 9.456 20.864 11.964 ;
  LAYER M3 ;
        RECT 20.768 9.456 20.8 11.964 ;
  LAYER M3 ;
        RECT 20.704 9.456 20.736 11.964 ;
  LAYER M3 ;
        RECT 20.64 9.456 20.672 11.964 ;
  LAYER M3 ;
        RECT 20.576 9.456 20.608 11.964 ;
  LAYER M3 ;
        RECT 20.512 9.456 20.544 11.964 ;
  LAYER M3 ;
        RECT 20.448 9.456 20.48 11.964 ;
  LAYER M3 ;
        RECT 20.384 9.456 20.416 11.964 ;
  LAYER M3 ;
        RECT 20.32 9.456 20.352 11.964 ;
  LAYER M3 ;
        RECT 20.256 9.456 20.288 11.964 ;
  LAYER M3 ;
        RECT 20.192 9.456 20.224 11.964 ;
  LAYER M3 ;
        RECT 20.128 9.456 20.16 11.964 ;
  LAYER M3 ;
        RECT 20.064 9.456 20.096 11.964 ;
  LAYER M3 ;
        RECT 20 9.456 20.032 11.964 ;
  LAYER M3 ;
        RECT 19.936 9.456 19.968 11.964 ;
  LAYER M3 ;
        RECT 19.872 9.456 19.904 11.964 ;
  LAYER M3 ;
        RECT 19.808 9.456 19.84 11.964 ;
  LAYER M3 ;
        RECT 19.744 9.456 19.776 11.964 ;
  LAYER M3 ;
        RECT 19.68 9.456 19.712 11.964 ;
  LAYER M3 ;
        RECT 19.616 9.456 19.648 11.964 ;
  LAYER M3 ;
        RECT 19.552 9.456 19.584 11.964 ;
  LAYER M3 ;
        RECT 19.488 9.456 19.52 11.964 ;
  LAYER M3 ;
        RECT 19.424 9.456 19.456 11.964 ;
  LAYER M3 ;
        RECT 19.36 9.456 19.392 11.964 ;
  LAYER M3 ;
        RECT 19.296 9.456 19.328 11.964 ;
  LAYER M3 ;
        RECT 19.232 9.456 19.264 11.964 ;
  LAYER M3 ;
        RECT 19.168 9.456 19.2 11.964 ;
  LAYER M3 ;
        RECT 19.104 9.456 19.136 11.964 ;
  LAYER M3 ;
        RECT 19.04 9.456 19.072 11.964 ;
  LAYER M3 ;
        RECT 18.944 9.456 18.976 11.964 ;
  LAYER M1 ;
        RECT 21.359 9.492 21.361 11.928 ;
  LAYER M1 ;
        RECT 21.279 9.492 21.281 11.928 ;
  LAYER M1 ;
        RECT 21.199 9.492 21.201 11.928 ;
  LAYER M1 ;
        RECT 21.119 9.492 21.121 11.928 ;
  LAYER M1 ;
        RECT 21.039 9.492 21.041 11.928 ;
  LAYER M1 ;
        RECT 20.959 9.492 20.961 11.928 ;
  LAYER M1 ;
        RECT 20.879 9.492 20.881 11.928 ;
  LAYER M1 ;
        RECT 20.799 9.492 20.801 11.928 ;
  LAYER M1 ;
        RECT 20.719 9.492 20.721 11.928 ;
  LAYER M1 ;
        RECT 20.639 9.492 20.641 11.928 ;
  LAYER M1 ;
        RECT 20.559 9.492 20.561 11.928 ;
  LAYER M1 ;
        RECT 20.479 9.492 20.481 11.928 ;
  LAYER M1 ;
        RECT 20.399 9.492 20.401 11.928 ;
  LAYER M1 ;
        RECT 20.319 9.492 20.321 11.928 ;
  LAYER M1 ;
        RECT 20.239 9.492 20.241 11.928 ;
  LAYER M1 ;
        RECT 20.159 9.492 20.161 11.928 ;
  LAYER M1 ;
        RECT 20.079 9.492 20.081 11.928 ;
  LAYER M1 ;
        RECT 19.999 9.492 20.001 11.928 ;
  LAYER M1 ;
        RECT 19.919 9.492 19.921 11.928 ;
  LAYER M1 ;
        RECT 19.839 9.492 19.841 11.928 ;
  LAYER M1 ;
        RECT 19.759 9.492 19.761 11.928 ;
  LAYER M1 ;
        RECT 19.679 9.492 19.681 11.928 ;
  LAYER M1 ;
        RECT 19.599 9.492 19.601 11.928 ;
  LAYER M1 ;
        RECT 19.519 9.492 19.521 11.928 ;
  LAYER M1 ;
        RECT 19.439 9.492 19.441 11.928 ;
  LAYER M1 ;
        RECT 19.359 9.492 19.361 11.928 ;
  LAYER M1 ;
        RECT 19.279 9.492 19.281 11.928 ;
  LAYER M1 ;
        RECT 19.199 9.492 19.201 11.928 ;
  LAYER M1 ;
        RECT 19.119 9.492 19.121 11.928 ;
  LAYER M1 ;
        RECT 19.039 9.492 19.041 11.928 ;
  LAYER M2 ;
        RECT 18.96 11.927 21.36 11.929 ;
  LAYER M2 ;
        RECT 18.96 11.843 21.36 11.845 ;
  LAYER M2 ;
        RECT 18.96 11.759 21.36 11.761 ;
  LAYER M2 ;
        RECT 18.96 11.675 21.36 11.677 ;
  LAYER M2 ;
        RECT 18.96 11.591 21.36 11.593 ;
  LAYER M2 ;
        RECT 18.96 11.507 21.36 11.509 ;
  LAYER M2 ;
        RECT 18.96 11.423 21.36 11.425 ;
  LAYER M2 ;
        RECT 18.96 11.339 21.36 11.341 ;
  LAYER M2 ;
        RECT 18.96 11.255 21.36 11.257 ;
  LAYER M2 ;
        RECT 18.96 11.171 21.36 11.173 ;
  LAYER M2 ;
        RECT 18.96 11.087 21.36 11.089 ;
  LAYER M2 ;
        RECT 18.96 11.003 21.36 11.005 ;
  LAYER M2 ;
        RECT 18.96 10.9195 21.36 10.9215 ;
  LAYER M2 ;
        RECT 18.96 10.835 21.36 10.837 ;
  LAYER M2 ;
        RECT 18.96 10.751 21.36 10.753 ;
  LAYER M2 ;
        RECT 18.96 10.667 21.36 10.669 ;
  LAYER M2 ;
        RECT 18.96 10.583 21.36 10.585 ;
  LAYER M2 ;
        RECT 18.96 10.499 21.36 10.501 ;
  LAYER M2 ;
        RECT 18.96 10.415 21.36 10.417 ;
  LAYER M2 ;
        RECT 18.96 10.331 21.36 10.333 ;
  LAYER M2 ;
        RECT 18.96 10.247 21.36 10.249 ;
  LAYER M2 ;
        RECT 18.96 10.163 21.36 10.165 ;
  LAYER M2 ;
        RECT 18.96 10.079 21.36 10.081 ;
  LAYER M2 ;
        RECT 18.96 9.995 21.36 9.997 ;
  LAYER M2 ;
        RECT 18.96 9.911 21.36 9.913 ;
  LAYER M2 ;
        RECT 18.96 9.827 21.36 9.829 ;
  LAYER M2 ;
        RECT 18.96 9.743 21.36 9.745 ;
  LAYER M2 ;
        RECT 18.96 9.659 21.36 9.661 ;
  LAYER M2 ;
        RECT 18.96 9.575 21.36 9.577 ;
  LAYER M1 ;
        RECT 21.344 6.516 21.376 9.024 ;
  LAYER M1 ;
        RECT 21.28 6.516 21.312 9.024 ;
  LAYER M1 ;
        RECT 21.216 6.516 21.248 9.024 ;
  LAYER M1 ;
        RECT 21.152 6.516 21.184 9.024 ;
  LAYER M1 ;
        RECT 21.088 6.516 21.12 9.024 ;
  LAYER M1 ;
        RECT 21.024 6.516 21.056 9.024 ;
  LAYER M1 ;
        RECT 20.96 6.516 20.992 9.024 ;
  LAYER M1 ;
        RECT 20.896 6.516 20.928 9.024 ;
  LAYER M1 ;
        RECT 20.832 6.516 20.864 9.024 ;
  LAYER M1 ;
        RECT 20.768 6.516 20.8 9.024 ;
  LAYER M1 ;
        RECT 20.704 6.516 20.736 9.024 ;
  LAYER M1 ;
        RECT 20.64 6.516 20.672 9.024 ;
  LAYER M1 ;
        RECT 20.576 6.516 20.608 9.024 ;
  LAYER M1 ;
        RECT 20.512 6.516 20.544 9.024 ;
  LAYER M1 ;
        RECT 20.448 6.516 20.48 9.024 ;
  LAYER M1 ;
        RECT 20.384 6.516 20.416 9.024 ;
  LAYER M1 ;
        RECT 20.32 6.516 20.352 9.024 ;
  LAYER M1 ;
        RECT 20.256 6.516 20.288 9.024 ;
  LAYER M1 ;
        RECT 20.192 6.516 20.224 9.024 ;
  LAYER M1 ;
        RECT 20.128 6.516 20.16 9.024 ;
  LAYER M1 ;
        RECT 20.064 6.516 20.096 9.024 ;
  LAYER M1 ;
        RECT 20 6.516 20.032 9.024 ;
  LAYER M1 ;
        RECT 19.936 6.516 19.968 9.024 ;
  LAYER M1 ;
        RECT 19.872 6.516 19.904 9.024 ;
  LAYER M1 ;
        RECT 19.808 6.516 19.84 9.024 ;
  LAYER M1 ;
        RECT 19.744 6.516 19.776 9.024 ;
  LAYER M1 ;
        RECT 19.68 6.516 19.712 9.024 ;
  LAYER M1 ;
        RECT 19.616 6.516 19.648 9.024 ;
  LAYER M1 ;
        RECT 19.552 6.516 19.584 9.024 ;
  LAYER M1 ;
        RECT 19.488 6.516 19.52 9.024 ;
  LAYER M1 ;
        RECT 19.424 6.516 19.456 9.024 ;
  LAYER M1 ;
        RECT 19.36 6.516 19.392 9.024 ;
  LAYER M1 ;
        RECT 19.296 6.516 19.328 9.024 ;
  LAYER M1 ;
        RECT 19.232 6.516 19.264 9.024 ;
  LAYER M1 ;
        RECT 19.168 6.516 19.2 9.024 ;
  LAYER M1 ;
        RECT 19.104 6.516 19.136 9.024 ;
  LAYER M1 ;
        RECT 19.04 6.516 19.072 9.024 ;
  LAYER M2 ;
        RECT 18.924 8.908 21.396 8.94 ;
  LAYER M2 ;
        RECT 18.924 8.844 21.396 8.876 ;
  LAYER M2 ;
        RECT 18.924 8.78 21.396 8.812 ;
  LAYER M2 ;
        RECT 18.924 8.716 21.396 8.748 ;
  LAYER M2 ;
        RECT 18.924 8.652 21.396 8.684 ;
  LAYER M2 ;
        RECT 18.924 8.588 21.396 8.62 ;
  LAYER M2 ;
        RECT 18.924 8.524 21.396 8.556 ;
  LAYER M2 ;
        RECT 18.924 8.46 21.396 8.492 ;
  LAYER M2 ;
        RECT 18.924 8.396 21.396 8.428 ;
  LAYER M2 ;
        RECT 18.924 8.332 21.396 8.364 ;
  LAYER M2 ;
        RECT 18.924 8.268 21.396 8.3 ;
  LAYER M2 ;
        RECT 18.924 8.204 21.396 8.236 ;
  LAYER M2 ;
        RECT 18.924 8.14 21.396 8.172 ;
  LAYER M2 ;
        RECT 18.924 8.076 21.396 8.108 ;
  LAYER M2 ;
        RECT 18.924 8.012 21.396 8.044 ;
  LAYER M2 ;
        RECT 18.924 7.948 21.396 7.98 ;
  LAYER M2 ;
        RECT 18.924 7.884 21.396 7.916 ;
  LAYER M2 ;
        RECT 18.924 7.82 21.396 7.852 ;
  LAYER M2 ;
        RECT 18.924 7.756 21.396 7.788 ;
  LAYER M2 ;
        RECT 18.924 7.692 21.396 7.724 ;
  LAYER M2 ;
        RECT 18.924 7.628 21.396 7.66 ;
  LAYER M2 ;
        RECT 18.924 7.564 21.396 7.596 ;
  LAYER M2 ;
        RECT 18.924 7.5 21.396 7.532 ;
  LAYER M2 ;
        RECT 18.924 7.436 21.396 7.468 ;
  LAYER M2 ;
        RECT 18.924 7.372 21.396 7.404 ;
  LAYER M2 ;
        RECT 18.924 7.308 21.396 7.34 ;
  LAYER M2 ;
        RECT 18.924 7.244 21.396 7.276 ;
  LAYER M2 ;
        RECT 18.924 7.18 21.396 7.212 ;
  LAYER M2 ;
        RECT 18.924 7.116 21.396 7.148 ;
  LAYER M2 ;
        RECT 18.924 7.052 21.396 7.084 ;
  LAYER M2 ;
        RECT 18.924 6.988 21.396 7.02 ;
  LAYER M2 ;
        RECT 18.924 6.924 21.396 6.956 ;
  LAYER M2 ;
        RECT 18.924 6.86 21.396 6.892 ;
  LAYER M2 ;
        RECT 18.924 6.796 21.396 6.828 ;
  LAYER M2 ;
        RECT 18.924 6.732 21.396 6.764 ;
  LAYER M2 ;
        RECT 18.924 6.668 21.396 6.7 ;
  LAYER M3 ;
        RECT 21.344 6.516 21.376 9.024 ;
  LAYER M3 ;
        RECT 21.28 6.516 21.312 9.024 ;
  LAYER M3 ;
        RECT 21.216 6.516 21.248 9.024 ;
  LAYER M3 ;
        RECT 21.152 6.516 21.184 9.024 ;
  LAYER M3 ;
        RECT 21.088 6.516 21.12 9.024 ;
  LAYER M3 ;
        RECT 21.024 6.516 21.056 9.024 ;
  LAYER M3 ;
        RECT 20.96 6.516 20.992 9.024 ;
  LAYER M3 ;
        RECT 20.896 6.516 20.928 9.024 ;
  LAYER M3 ;
        RECT 20.832 6.516 20.864 9.024 ;
  LAYER M3 ;
        RECT 20.768 6.516 20.8 9.024 ;
  LAYER M3 ;
        RECT 20.704 6.516 20.736 9.024 ;
  LAYER M3 ;
        RECT 20.64 6.516 20.672 9.024 ;
  LAYER M3 ;
        RECT 20.576 6.516 20.608 9.024 ;
  LAYER M3 ;
        RECT 20.512 6.516 20.544 9.024 ;
  LAYER M3 ;
        RECT 20.448 6.516 20.48 9.024 ;
  LAYER M3 ;
        RECT 20.384 6.516 20.416 9.024 ;
  LAYER M3 ;
        RECT 20.32 6.516 20.352 9.024 ;
  LAYER M3 ;
        RECT 20.256 6.516 20.288 9.024 ;
  LAYER M3 ;
        RECT 20.192 6.516 20.224 9.024 ;
  LAYER M3 ;
        RECT 20.128 6.516 20.16 9.024 ;
  LAYER M3 ;
        RECT 20.064 6.516 20.096 9.024 ;
  LAYER M3 ;
        RECT 20 6.516 20.032 9.024 ;
  LAYER M3 ;
        RECT 19.936 6.516 19.968 9.024 ;
  LAYER M3 ;
        RECT 19.872 6.516 19.904 9.024 ;
  LAYER M3 ;
        RECT 19.808 6.516 19.84 9.024 ;
  LAYER M3 ;
        RECT 19.744 6.516 19.776 9.024 ;
  LAYER M3 ;
        RECT 19.68 6.516 19.712 9.024 ;
  LAYER M3 ;
        RECT 19.616 6.516 19.648 9.024 ;
  LAYER M3 ;
        RECT 19.552 6.516 19.584 9.024 ;
  LAYER M3 ;
        RECT 19.488 6.516 19.52 9.024 ;
  LAYER M3 ;
        RECT 19.424 6.516 19.456 9.024 ;
  LAYER M3 ;
        RECT 19.36 6.516 19.392 9.024 ;
  LAYER M3 ;
        RECT 19.296 6.516 19.328 9.024 ;
  LAYER M3 ;
        RECT 19.232 6.516 19.264 9.024 ;
  LAYER M3 ;
        RECT 19.168 6.516 19.2 9.024 ;
  LAYER M3 ;
        RECT 19.104 6.516 19.136 9.024 ;
  LAYER M3 ;
        RECT 19.04 6.516 19.072 9.024 ;
  LAYER M3 ;
        RECT 18.944 6.516 18.976 9.024 ;
  LAYER M1 ;
        RECT 21.359 6.552 21.361 8.988 ;
  LAYER M1 ;
        RECT 21.279 6.552 21.281 8.988 ;
  LAYER M1 ;
        RECT 21.199 6.552 21.201 8.988 ;
  LAYER M1 ;
        RECT 21.119 6.552 21.121 8.988 ;
  LAYER M1 ;
        RECT 21.039 6.552 21.041 8.988 ;
  LAYER M1 ;
        RECT 20.959 6.552 20.961 8.988 ;
  LAYER M1 ;
        RECT 20.879 6.552 20.881 8.988 ;
  LAYER M1 ;
        RECT 20.799 6.552 20.801 8.988 ;
  LAYER M1 ;
        RECT 20.719 6.552 20.721 8.988 ;
  LAYER M1 ;
        RECT 20.639 6.552 20.641 8.988 ;
  LAYER M1 ;
        RECT 20.559 6.552 20.561 8.988 ;
  LAYER M1 ;
        RECT 20.479 6.552 20.481 8.988 ;
  LAYER M1 ;
        RECT 20.399 6.552 20.401 8.988 ;
  LAYER M1 ;
        RECT 20.319 6.552 20.321 8.988 ;
  LAYER M1 ;
        RECT 20.239 6.552 20.241 8.988 ;
  LAYER M1 ;
        RECT 20.159 6.552 20.161 8.988 ;
  LAYER M1 ;
        RECT 20.079 6.552 20.081 8.988 ;
  LAYER M1 ;
        RECT 19.999 6.552 20.001 8.988 ;
  LAYER M1 ;
        RECT 19.919 6.552 19.921 8.988 ;
  LAYER M1 ;
        RECT 19.839 6.552 19.841 8.988 ;
  LAYER M1 ;
        RECT 19.759 6.552 19.761 8.988 ;
  LAYER M1 ;
        RECT 19.679 6.552 19.681 8.988 ;
  LAYER M1 ;
        RECT 19.599 6.552 19.601 8.988 ;
  LAYER M1 ;
        RECT 19.519 6.552 19.521 8.988 ;
  LAYER M1 ;
        RECT 19.439 6.552 19.441 8.988 ;
  LAYER M1 ;
        RECT 19.359 6.552 19.361 8.988 ;
  LAYER M1 ;
        RECT 19.279 6.552 19.281 8.988 ;
  LAYER M1 ;
        RECT 19.199 6.552 19.201 8.988 ;
  LAYER M1 ;
        RECT 19.119 6.552 19.121 8.988 ;
  LAYER M1 ;
        RECT 19.039 6.552 19.041 8.988 ;
  LAYER M2 ;
        RECT 18.96 8.987 21.36 8.989 ;
  LAYER M2 ;
        RECT 18.96 8.903 21.36 8.905 ;
  LAYER M2 ;
        RECT 18.96 8.819 21.36 8.821 ;
  LAYER M2 ;
        RECT 18.96 8.735 21.36 8.737 ;
  LAYER M2 ;
        RECT 18.96 8.651 21.36 8.653 ;
  LAYER M2 ;
        RECT 18.96 8.567 21.36 8.569 ;
  LAYER M2 ;
        RECT 18.96 8.483 21.36 8.485 ;
  LAYER M2 ;
        RECT 18.96 8.399 21.36 8.401 ;
  LAYER M2 ;
        RECT 18.96 8.315 21.36 8.317 ;
  LAYER M2 ;
        RECT 18.96 8.231 21.36 8.233 ;
  LAYER M2 ;
        RECT 18.96 8.147 21.36 8.149 ;
  LAYER M2 ;
        RECT 18.96 8.063 21.36 8.065 ;
  LAYER M2 ;
        RECT 18.96 7.9795 21.36 7.9815 ;
  LAYER M2 ;
        RECT 18.96 7.895 21.36 7.897 ;
  LAYER M2 ;
        RECT 18.96 7.811 21.36 7.813 ;
  LAYER M2 ;
        RECT 18.96 7.727 21.36 7.729 ;
  LAYER M2 ;
        RECT 18.96 7.643 21.36 7.645 ;
  LAYER M2 ;
        RECT 18.96 7.559 21.36 7.561 ;
  LAYER M2 ;
        RECT 18.96 7.475 21.36 7.477 ;
  LAYER M2 ;
        RECT 18.96 7.391 21.36 7.393 ;
  LAYER M2 ;
        RECT 18.96 7.307 21.36 7.309 ;
  LAYER M2 ;
        RECT 18.96 7.223 21.36 7.225 ;
  LAYER M2 ;
        RECT 18.96 7.139 21.36 7.141 ;
  LAYER M2 ;
        RECT 18.96 7.055 21.36 7.057 ;
  LAYER M2 ;
        RECT 18.96 6.971 21.36 6.973 ;
  LAYER M2 ;
        RECT 18.96 6.887 21.36 6.889 ;
  LAYER M2 ;
        RECT 18.96 6.803 21.36 6.805 ;
  LAYER M2 ;
        RECT 18.96 6.719 21.36 6.721 ;
  LAYER M2 ;
        RECT 18.96 6.635 21.36 6.637 ;
  LAYER M1 ;
        RECT 18.464 15.336 18.496 17.844 ;
  LAYER M1 ;
        RECT 18.4 15.336 18.432 17.844 ;
  LAYER M1 ;
        RECT 18.336 15.336 18.368 17.844 ;
  LAYER M1 ;
        RECT 18.272 15.336 18.304 17.844 ;
  LAYER M1 ;
        RECT 18.208 15.336 18.24 17.844 ;
  LAYER M1 ;
        RECT 18.144 15.336 18.176 17.844 ;
  LAYER M1 ;
        RECT 18.08 15.336 18.112 17.844 ;
  LAYER M1 ;
        RECT 18.016 15.336 18.048 17.844 ;
  LAYER M1 ;
        RECT 17.952 15.336 17.984 17.844 ;
  LAYER M1 ;
        RECT 17.888 15.336 17.92 17.844 ;
  LAYER M1 ;
        RECT 17.824 15.336 17.856 17.844 ;
  LAYER M1 ;
        RECT 17.76 15.336 17.792 17.844 ;
  LAYER M1 ;
        RECT 17.696 15.336 17.728 17.844 ;
  LAYER M1 ;
        RECT 17.632 15.336 17.664 17.844 ;
  LAYER M1 ;
        RECT 17.568 15.336 17.6 17.844 ;
  LAYER M1 ;
        RECT 17.504 15.336 17.536 17.844 ;
  LAYER M1 ;
        RECT 17.44 15.336 17.472 17.844 ;
  LAYER M1 ;
        RECT 17.376 15.336 17.408 17.844 ;
  LAYER M1 ;
        RECT 17.312 15.336 17.344 17.844 ;
  LAYER M1 ;
        RECT 17.248 15.336 17.28 17.844 ;
  LAYER M1 ;
        RECT 17.184 15.336 17.216 17.844 ;
  LAYER M1 ;
        RECT 17.12 15.336 17.152 17.844 ;
  LAYER M1 ;
        RECT 17.056 15.336 17.088 17.844 ;
  LAYER M1 ;
        RECT 16.992 15.336 17.024 17.844 ;
  LAYER M1 ;
        RECT 16.928 15.336 16.96 17.844 ;
  LAYER M1 ;
        RECT 16.864 15.336 16.896 17.844 ;
  LAYER M1 ;
        RECT 16.8 15.336 16.832 17.844 ;
  LAYER M1 ;
        RECT 16.736 15.336 16.768 17.844 ;
  LAYER M1 ;
        RECT 16.672 15.336 16.704 17.844 ;
  LAYER M1 ;
        RECT 16.608 15.336 16.64 17.844 ;
  LAYER M1 ;
        RECT 16.544 15.336 16.576 17.844 ;
  LAYER M1 ;
        RECT 16.48 15.336 16.512 17.844 ;
  LAYER M1 ;
        RECT 16.416 15.336 16.448 17.844 ;
  LAYER M1 ;
        RECT 16.352 15.336 16.384 17.844 ;
  LAYER M1 ;
        RECT 16.288 15.336 16.32 17.844 ;
  LAYER M1 ;
        RECT 16.224 15.336 16.256 17.844 ;
  LAYER M1 ;
        RECT 16.16 15.336 16.192 17.844 ;
  LAYER M2 ;
        RECT 16.044 17.728 18.516 17.76 ;
  LAYER M2 ;
        RECT 16.044 17.664 18.516 17.696 ;
  LAYER M2 ;
        RECT 16.044 17.6 18.516 17.632 ;
  LAYER M2 ;
        RECT 16.044 17.536 18.516 17.568 ;
  LAYER M2 ;
        RECT 16.044 17.472 18.516 17.504 ;
  LAYER M2 ;
        RECT 16.044 17.408 18.516 17.44 ;
  LAYER M2 ;
        RECT 16.044 17.344 18.516 17.376 ;
  LAYER M2 ;
        RECT 16.044 17.28 18.516 17.312 ;
  LAYER M2 ;
        RECT 16.044 17.216 18.516 17.248 ;
  LAYER M2 ;
        RECT 16.044 17.152 18.516 17.184 ;
  LAYER M2 ;
        RECT 16.044 17.088 18.516 17.12 ;
  LAYER M2 ;
        RECT 16.044 17.024 18.516 17.056 ;
  LAYER M2 ;
        RECT 16.044 16.96 18.516 16.992 ;
  LAYER M2 ;
        RECT 16.044 16.896 18.516 16.928 ;
  LAYER M2 ;
        RECT 16.044 16.832 18.516 16.864 ;
  LAYER M2 ;
        RECT 16.044 16.768 18.516 16.8 ;
  LAYER M2 ;
        RECT 16.044 16.704 18.516 16.736 ;
  LAYER M2 ;
        RECT 16.044 16.64 18.516 16.672 ;
  LAYER M2 ;
        RECT 16.044 16.576 18.516 16.608 ;
  LAYER M2 ;
        RECT 16.044 16.512 18.516 16.544 ;
  LAYER M2 ;
        RECT 16.044 16.448 18.516 16.48 ;
  LAYER M2 ;
        RECT 16.044 16.384 18.516 16.416 ;
  LAYER M2 ;
        RECT 16.044 16.32 18.516 16.352 ;
  LAYER M2 ;
        RECT 16.044 16.256 18.516 16.288 ;
  LAYER M2 ;
        RECT 16.044 16.192 18.516 16.224 ;
  LAYER M2 ;
        RECT 16.044 16.128 18.516 16.16 ;
  LAYER M2 ;
        RECT 16.044 16.064 18.516 16.096 ;
  LAYER M2 ;
        RECT 16.044 16 18.516 16.032 ;
  LAYER M2 ;
        RECT 16.044 15.936 18.516 15.968 ;
  LAYER M2 ;
        RECT 16.044 15.872 18.516 15.904 ;
  LAYER M2 ;
        RECT 16.044 15.808 18.516 15.84 ;
  LAYER M2 ;
        RECT 16.044 15.744 18.516 15.776 ;
  LAYER M2 ;
        RECT 16.044 15.68 18.516 15.712 ;
  LAYER M2 ;
        RECT 16.044 15.616 18.516 15.648 ;
  LAYER M2 ;
        RECT 16.044 15.552 18.516 15.584 ;
  LAYER M2 ;
        RECT 16.044 15.488 18.516 15.52 ;
  LAYER M3 ;
        RECT 18.464 15.336 18.496 17.844 ;
  LAYER M3 ;
        RECT 18.4 15.336 18.432 17.844 ;
  LAYER M3 ;
        RECT 18.336 15.336 18.368 17.844 ;
  LAYER M3 ;
        RECT 18.272 15.336 18.304 17.844 ;
  LAYER M3 ;
        RECT 18.208 15.336 18.24 17.844 ;
  LAYER M3 ;
        RECT 18.144 15.336 18.176 17.844 ;
  LAYER M3 ;
        RECT 18.08 15.336 18.112 17.844 ;
  LAYER M3 ;
        RECT 18.016 15.336 18.048 17.844 ;
  LAYER M3 ;
        RECT 17.952 15.336 17.984 17.844 ;
  LAYER M3 ;
        RECT 17.888 15.336 17.92 17.844 ;
  LAYER M3 ;
        RECT 17.824 15.336 17.856 17.844 ;
  LAYER M3 ;
        RECT 17.76 15.336 17.792 17.844 ;
  LAYER M3 ;
        RECT 17.696 15.336 17.728 17.844 ;
  LAYER M3 ;
        RECT 17.632 15.336 17.664 17.844 ;
  LAYER M3 ;
        RECT 17.568 15.336 17.6 17.844 ;
  LAYER M3 ;
        RECT 17.504 15.336 17.536 17.844 ;
  LAYER M3 ;
        RECT 17.44 15.336 17.472 17.844 ;
  LAYER M3 ;
        RECT 17.376 15.336 17.408 17.844 ;
  LAYER M3 ;
        RECT 17.312 15.336 17.344 17.844 ;
  LAYER M3 ;
        RECT 17.248 15.336 17.28 17.844 ;
  LAYER M3 ;
        RECT 17.184 15.336 17.216 17.844 ;
  LAYER M3 ;
        RECT 17.12 15.336 17.152 17.844 ;
  LAYER M3 ;
        RECT 17.056 15.336 17.088 17.844 ;
  LAYER M3 ;
        RECT 16.992 15.336 17.024 17.844 ;
  LAYER M3 ;
        RECT 16.928 15.336 16.96 17.844 ;
  LAYER M3 ;
        RECT 16.864 15.336 16.896 17.844 ;
  LAYER M3 ;
        RECT 16.8 15.336 16.832 17.844 ;
  LAYER M3 ;
        RECT 16.736 15.336 16.768 17.844 ;
  LAYER M3 ;
        RECT 16.672 15.336 16.704 17.844 ;
  LAYER M3 ;
        RECT 16.608 15.336 16.64 17.844 ;
  LAYER M3 ;
        RECT 16.544 15.336 16.576 17.844 ;
  LAYER M3 ;
        RECT 16.48 15.336 16.512 17.844 ;
  LAYER M3 ;
        RECT 16.416 15.336 16.448 17.844 ;
  LAYER M3 ;
        RECT 16.352 15.336 16.384 17.844 ;
  LAYER M3 ;
        RECT 16.288 15.336 16.32 17.844 ;
  LAYER M3 ;
        RECT 16.224 15.336 16.256 17.844 ;
  LAYER M3 ;
        RECT 16.16 15.336 16.192 17.844 ;
  LAYER M3 ;
        RECT 16.064 15.336 16.096 17.844 ;
  LAYER M1 ;
        RECT 18.479 15.372 18.481 17.808 ;
  LAYER M1 ;
        RECT 18.399 15.372 18.401 17.808 ;
  LAYER M1 ;
        RECT 18.319 15.372 18.321 17.808 ;
  LAYER M1 ;
        RECT 18.239 15.372 18.241 17.808 ;
  LAYER M1 ;
        RECT 18.159 15.372 18.161 17.808 ;
  LAYER M1 ;
        RECT 18.079 15.372 18.081 17.808 ;
  LAYER M1 ;
        RECT 17.999 15.372 18.001 17.808 ;
  LAYER M1 ;
        RECT 17.919 15.372 17.921 17.808 ;
  LAYER M1 ;
        RECT 17.839 15.372 17.841 17.808 ;
  LAYER M1 ;
        RECT 17.759 15.372 17.761 17.808 ;
  LAYER M1 ;
        RECT 17.679 15.372 17.681 17.808 ;
  LAYER M1 ;
        RECT 17.599 15.372 17.601 17.808 ;
  LAYER M1 ;
        RECT 17.519 15.372 17.521 17.808 ;
  LAYER M1 ;
        RECT 17.439 15.372 17.441 17.808 ;
  LAYER M1 ;
        RECT 17.359 15.372 17.361 17.808 ;
  LAYER M1 ;
        RECT 17.279 15.372 17.281 17.808 ;
  LAYER M1 ;
        RECT 17.199 15.372 17.201 17.808 ;
  LAYER M1 ;
        RECT 17.119 15.372 17.121 17.808 ;
  LAYER M1 ;
        RECT 17.039 15.372 17.041 17.808 ;
  LAYER M1 ;
        RECT 16.959 15.372 16.961 17.808 ;
  LAYER M1 ;
        RECT 16.879 15.372 16.881 17.808 ;
  LAYER M1 ;
        RECT 16.799 15.372 16.801 17.808 ;
  LAYER M1 ;
        RECT 16.719 15.372 16.721 17.808 ;
  LAYER M1 ;
        RECT 16.639 15.372 16.641 17.808 ;
  LAYER M1 ;
        RECT 16.559 15.372 16.561 17.808 ;
  LAYER M1 ;
        RECT 16.479 15.372 16.481 17.808 ;
  LAYER M1 ;
        RECT 16.399 15.372 16.401 17.808 ;
  LAYER M1 ;
        RECT 16.319 15.372 16.321 17.808 ;
  LAYER M1 ;
        RECT 16.239 15.372 16.241 17.808 ;
  LAYER M1 ;
        RECT 16.159 15.372 16.161 17.808 ;
  LAYER M2 ;
        RECT 16.08 17.807 18.48 17.809 ;
  LAYER M2 ;
        RECT 16.08 17.723 18.48 17.725 ;
  LAYER M2 ;
        RECT 16.08 17.639 18.48 17.641 ;
  LAYER M2 ;
        RECT 16.08 17.555 18.48 17.557 ;
  LAYER M2 ;
        RECT 16.08 17.471 18.48 17.473 ;
  LAYER M2 ;
        RECT 16.08 17.387 18.48 17.389 ;
  LAYER M2 ;
        RECT 16.08 17.303 18.48 17.305 ;
  LAYER M2 ;
        RECT 16.08 17.219 18.48 17.221 ;
  LAYER M2 ;
        RECT 16.08 17.135 18.48 17.137 ;
  LAYER M2 ;
        RECT 16.08 17.051 18.48 17.053 ;
  LAYER M2 ;
        RECT 16.08 16.967 18.48 16.969 ;
  LAYER M2 ;
        RECT 16.08 16.883 18.48 16.885 ;
  LAYER M2 ;
        RECT 16.08 16.7995 18.48 16.8015 ;
  LAYER M2 ;
        RECT 16.08 16.715 18.48 16.717 ;
  LAYER M2 ;
        RECT 16.08 16.631 18.48 16.633 ;
  LAYER M2 ;
        RECT 16.08 16.547 18.48 16.549 ;
  LAYER M2 ;
        RECT 16.08 16.463 18.48 16.465 ;
  LAYER M2 ;
        RECT 16.08 16.379 18.48 16.381 ;
  LAYER M2 ;
        RECT 16.08 16.295 18.48 16.297 ;
  LAYER M2 ;
        RECT 16.08 16.211 18.48 16.213 ;
  LAYER M2 ;
        RECT 16.08 16.127 18.48 16.129 ;
  LAYER M2 ;
        RECT 16.08 16.043 18.48 16.045 ;
  LAYER M2 ;
        RECT 16.08 15.959 18.48 15.961 ;
  LAYER M2 ;
        RECT 16.08 15.875 18.48 15.877 ;
  LAYER M2 ;
        RECT 16.08 15.791 18.48 15.793 ;
  LAYER M2 ;
        RECT 16.08 15.707 18.48 15.709 ;
  LAYER M2 ;
        RECT 16.08 15.623 18.48 15.625 ;
  LAYER M2 ;
        RECT 16.08 15.539 18.48 15.541 ;
  LAYER M2 ;
        RECT 16.08 15.455 18.48 15.457 ;
  LAYER M1 ;
        RECT 18.464 12.396 18.496 14.904 ;
  LAYER M1 ;
        RECT 18.4 12.396 18.432 14.904 ;
  LAYER M1 ;
        RECT 18.336 12.396 18.368 14.904 ;
  LAYER M1 ;
        RECT 18.272 12.396 18.304 14.904 ;
  LAYER M1 ;
        RECT 18.208 12.396 18.24 14.904 ;
  LAYER M1 ;
        RECT 18.144 12.396 18.176 14.904 ;
  LAYER M1 ;
        RECT 18.08 12.396 18.112 14.904 ;
  LAYER M1 ;
        RECT 18.016 12.396 18.048 14.904 ;
  LAYER M1 ;
        RECT 17.952 12.396 17.984 14.904 ;
  LAYER M1 ;
        RECT 17.888 12.396 17.92 14.904 ;
  LAYER M1 ;
        RECT 17.824 12.396 17.856 14.904 ;
  LAYER M1 ;
        RECT 17.76 12.396 17.792 14.904 ;
  LAYER M1 ;
        RECT 17.696 12.396 17.728 14.904 ;
  LAYER M1 ;
        RECT 17.632 12.396 17.664 14.904 ;
  LAYER M1 ;
        RECT 17.568 12.396 17.6 14.904 ;
  LAYER M1 ;
        RECT 17.504 12.396 17.536 14.904 ;
  LAYER M1 ;
        RECT 17.44 12.396 17.472 14.904 ;
  LAYER M1 ;
        RECT 17.376 12.396 17.408 14.904 ;
  LAYER M1 ;
        RECT 17.312 12.396 17.344 14.904 ;
  LAYER M1 ;
        RECT 17.248 12.396 17.28 14.904 ;
  LAYER M1 ;
        RECT 17.184 12.396 17.216 14.904 ;
  LAYER M1 ;
        RECT 17.12 12.396 17.152 14.904 ;
  LAYER M1 ;
        RECT 17.056 12.396 17.088 14.904 ;
  LAYER M1 ;
        RECT 16.992 12.396 17.024 14.904 ;
  LAYER M1 ;
        RECT 16.928 12.396 16.96 14.904 ;
  LAYER M1 ;
        RECT 16.864 12.396 16.896 14.904 ;
  LAYER M1 ;
        RECT 16.8 12.396 16.832 14.904 ;
  LAYER M1 ;
        RECT 16.736 12.396 16.768 14.904 ;
  LAYER M1 ;
        RECT 16.672 12.396 16.704 14.904 ;
  LAYER M1 ;
        RECT 16.608 12.396 16.64 14.904 ;
  LAYER M1 ;
        RECT 16.544 12.396 16.576 14.904 ;
  LAYER M1 ;
        RECT 16.48 12.396 16.512 14.904 ;
  LAYER M1 ;
        RECT 16.416 12.396 16.448 14.904 ;
  LAYER M1 ;
        RECT 16.352 12.396 16.384 14.904 ;
  LAYER M1 ;
        RECT 16.288 12.396 16.32 14.904 ;
  LAYER M1 ;
        RECT 16.224 12.396 16.256 14.904 ;
  LAYER M1 ;
        RECT 16.16 12.396 16.192 14.904 ;
  LAYER M2 ;
        RECT 16.044 14.788 18.516 14.82 ;
  LAYER M2 ;
        RECT 16.044 14.724 18.516 14.756 ;
  LAYER M2 ;
        RECT 16.044 14.66 18.516 14.692 ;
  LAYER M2 ;
        RECT 16.044 14.596 18.516 14.628 ;
  LAYER M2 ;
        RECT 16.044 14.532 18.516 14.564 ;
  LAYER M2 ;
        RECT 16.044 14.468 18.516 14.5 ;
  LAYER M2 ;
        RECT 16.044 14.404 18.516 14.436 ;
  LAYER M2 ;
        RECT 16.044 14.34 18.516 14.372 ;
  LAYER M2 ;
        RECT 16.044 14.276 18.516 14.308 ;
  LAYER M2 ;
        RECT 16.044 14.212 18.516 14.244 ;
  LAYER M2 ;
        RECT 16.044 14.148 18.516 14.18 ;
  LAYER M2 ;
        RECT 16.044 14.084 18.516 14.116 ;
  LAYER M2 ;
        RECT 16.044 14.02 18.516 14.052 ;
  LAYER M2 ;
        RECT 16.044 13.956 18.516 13.988 ;
  LAYER M2 ;
        RECT 16.044 13.892 18.516 13.924 ;
  LAYER M2 ;
        RECT 16.044 13.828 18.516 13.86 ;
  LAYER M2 ;
        RECT 16.044 13.764 18.516 13.796 ;
  LAYER M2 ;
        RECT 16.044 13.7 18.516 13.732 ;
  LAYER M2 ;
        RECT 16.044 13.636 18.516 13.668 ;
  LAYER M2 ;
        RECT 16.044 13.572 18.516 13.604 ;
  LAYER M2 ;
        RECT 16.044 13.508 18.516 13.54 ;
  LAYER M2 ;
        RECT 16.044 13.444 18.516 13.476 ;
  LAYER M2 ;
        RECT 16.044 13.38 18.516 13.412 ;
  LAYER M2 ;
        RECT 16.044 13.316 18.516 13.348 ;
  LAYER M2 ;
        RECT 16.044 13.252 18.516 13.284 ;
  LAYER M2 ;
        RECT 16.044 13.188 18.516 13.22 ;
  LAYER M2 ;
        RECT 16.044 13.124 18.516 13.156 ;
  LAYER M2 ;
        RECT 16.044 13.06 18.516 13.092 ;
  LAYER M2 ;
        RECT 16.044 12.996 18.516 13.028 ;
  LAYER M2 ;
        RECT 16.044 12.932 18.516 12.964 ;
  LAYER M2 ;
        RECT 16.044 12.868 18.516 12.9 ;
  LAYER M2 ;
        RECT 16.044 12.804 18.516 12.836 ;
  LAYER M2 ;
        RECT 16.044 12.74 18.516 12.772 ;
  LAYER M2 ;
        RECT 16.044 12.676 18.516 12.708 ;
  LAYER M2 ;
        RECT 16.044 12.612 18.516 12.644 ;
  LAYER M2 ;
        RECT 16.044 12.548 18.516 12.58 ;
  LAYER M3 ;
        RECT 18.464 12.396 18.496 14.904 ;
  LAYER M3 ;
        RECT 18.4 12.396 18.432 14.904 ;
  LAYER M3 ;
        RECT 18.336 12.396 18.368 14.904 ;
  LAYER M3 ;
        RECT 18.272 12.396 18.304 14.904 ;
  LAYER M3 ;
        RECT 18.208 12.396 18.24 14.904 ;
  LAYER M3 ;
        RECT 18.144 12.396 18.176 14.904 ;
  LAYER M3 ;
        RECT 18.08 12.396 18.112 14.904 ;
  LAYER M3 ;
        RECT 18.016 12.396 18.048 14.904 ;
  LAYER M3 ;
        RECT 17.952 12.396 17.984 14.904 ;
  LAYER M3 ;
        RECT 17.888 12.396 17.92 14.904 ;
  LAYER M3 ;
        RECT 17.824 12.396 17.856 14.904 ;
  LAYER M3 ;
        RECT 17.76 12.396 17.792 14.904 ;
  LAYER M3 ;
        RECT 17.696 12.396 17.728 14.904 ;
  LAYER M3 ;
        RECT 17.632 12.396 17.664 14.904 ;
  LAYER M3 ;
        RECT 17.568 12.396 17.6 14.904 ;
  LAYER M3 ;
        RECT 17.504 12.396 17.536 14.904 ;
  LAYER M3 ;
        RECT 17.44 12.396 17.472 14.904 ;
  LAYER M3 ;
        RECT 17.376 12.396 17.408 14.904 ;
  LAYER M3 ;
        RECT 17.312 12.396 17.344 14.904 ;
  LAYER M3 ;
        RECT 17.248 12.396 17.28 14.904 ;
  LAYER M3 ;
        RECT 17.184 12.396 17.216 14.904 ;
  LAYER M3 ;
        RECT 17.12 12.396 17.152 14.904 ;
  LAYER M3 ;
        RECT 17.056 12.396 17.088 14.904 ;
  LAYER M3 ;
        RECT 16.992 12.396 17.024 14.904 ;
  LAYER M3 ;
        RECT 16.928 12.396 16.96 14.904 ;
  LAYER M3 ;
        RECT 16.864 12.396 16.896 14.904 ;
  LAYER M3 ;
        RECT 16.8 12.396 16.832 14.904 ;
  LAYER M3 ;
        RECT 16.736 12.396 16.768 14.904 ;
  LAYER M3 ;
        RECT 16.672 12.396 16.704 14.904 ;
  LAYER M3 ;
        RECT 16.608 12.396 16.64 14.904 ;
  LAYER M3 ;
        RECT 16.544 12.396 16.576 14.904 ;
  LAYER M3 ;
        RECT 16.48 12.396 16.512 14.904 ;
  LAYER M3 ;
        RECT 16.416 12.396 16.448 14.904 ;
  LAYER M3 ;
        RECT 16.352 12.396 16.384 14.904 ;
  LAYER M3 ;
        RECT 16.288 12.396 16.32 14.904 ;
  LAYER M3 ;
        RECT 16.224 12.396 16.256 14.904 ;
  LAYER M3 ;
        RECT 16.16 12.396 16.192 14.904 ;
  LAYER M3 ;
        RECT 16.064 12.396 16.096 14.904 ;
  LAYER M1 ;
        RECT 18.479 12.432 18.481 14.868 ;
  LAYER M1 ;
        RECT 18.399 12.432 18.401 14.868 ;
  LAYER M1 ;
        RECT 18.319 12.432 18.321 14.868 ;
  LAYER M1 ;
        RECT 18.239 12.432 18.241 14.868 ;
  LAYER M1 ;
        RECT 18.159 12.432 18.161 14.868 ;
  LAYER M1 ;
        RECT 18.079 12.432 18.081 14.868 ;
  LAYER M1 ;
        RECT 17.999 12.432 18.001 14.868 ;
  LAYER M1 ;
        RECT 17.919 12.432 17.921 14.868 ;
  LAYER M1 ;
        RECT 17.839 12.432 17.841 14.868 ;
  LAYER M1 ;
        RECT 17.759 12.432 17.761 14.868 ;
  LAYER M1 ;
        RECT 17.679 12.432 17.681 14.868 ;
  LAYER M1 ;
        RECT 17.599 12.432 17.601 14.868 ;
  LAYER M1 ;
        RECT 17.519 12.432 17.521 14.868 ;
  LAYER M1 ;
        RECT 17.439 12.432 17.441 14.868 ;
  LAYER M1 ;
        RECT 17.359 12.432 17.361 14.868 ;
  LAYER M1 ;
        RECT 17.279 12.432 17.281 14.868 ;
  LAYER M1 ;
        RECT 17.199 12.432 17.201 14.868 ;
  LAYER M1 ;
        RECT 17.119 12.432 17.121 14.868 ;
  LAYER M1 ;
        RECT 17.039 12.432 17.041 14.868 ;
  LAYER M1 ;
        RECT 16.959 12.432 16.961 14.868 ;
  LAYER M1 ;
        RECT 16.879 12.432 16.881 14.868 ;
  LAYER M1 ;
        RECT 16.799 12.432 16.801 14.868 ;
  LAYER M1 ;
        RECT 16.719 12.432 16.721 14.868 ;
  LAYER M1 ;
        RECT 16.639 12.432 16.641 14.868 ;
  LAYER M1 ;
        RECT 16.559 12.432 16.561 14.868 ;
  LAYER M1 ;
        RECT 16.479 12.432 16.481 14.868 ;
  LAYER M1 ;
        RECT 16.399 12.432 16.401 14.868 ;
  LAYER M1 ;
        RECT 16.319 12.432 16.321 14.868 ;
  LAYER M1 ;
        RECT 16.239 12.432 16.241 14.868 ;
  LAYER M1 ;
        RECT 16.159 12.432 16.161 14.868 ;
  LAYER M2 ;
        RECT 16.08 14.867 18.48 14.869 ;
  LAYER M2 ;
        RECT 16.08 14.783 18.48 14.785 ;
  LAYER M2 ;
        RECT 16.08 14.699 18.48 14.701 ;
  LAYER M2 ;
        RECT 16.08 14.615 18.48 14.617 ;
  LAYER M2 ;
        RECT 16.08 14.531 18.48 14.533 ;
  LAYER M2 ;
        RECT 16.08 14.447 18.48 14.449 ;
  LAYER M2 ;
        RECT 16.08 14.363 18.48 14.365 ;
  LAYER M2 ;
        RECT 16.08 14.279 18.48 14.281 ;
  LAYER M2 ;
        RECT 16.08 14.195 18.48 14.197 ;
  LAYER M2 ;
        RECT 16.08 14.111 18.48 14.113 ;
  LAYER M2 ;
        RECT 16.08 14.027 18.48 14.029 ;
  LAYER M2 ;
        RECT 16.08 13.943 18.48 13.945 ;
  LAYER M2 ;
        RECT 16.08 13.8595 18.48 13.8615 ;
  LAYER M2 ;
        RECT 16.08 13.775 18.48 13.777 ;
  LAYER M2 ;
        RECT 16.08 13.691 18.48 13.693 ;
  LAYER M2 ;
        RECT 16.08 13.607 18.48 13.609 ;
  LAYER M2 ;
        RECT 16.08 13.523 18.48 13.525 ;
  LAYER M2 ;
        RECT 16.08 13.439 18.48 13.441 ;
  LAYER M2 ;
        RECT 16.08 13.355 18.48 13.357 ;
  LAYER M2 ;
        RECT 16.08 13.271 18.48 13.273 ;
  LAYER M2 ;
        RECT 16.08 13.187 18.48 13.189 ;
  LAYER M2 ;
        RECT 16.08 13.103 18.48 13.105 ;
  LAYER M2 ;
        RECT 16.08 13.019 18.48 13.021 ;
  LAYER M2 ;
        RECT 16.08 12.935 18.48 12.937 ;
  LAYER M2 ;
        RECT 16.08 12.851 18.48 12.853 ;
  LAYER M2 ;
        RECT 16.08 12.767 18.48 12.769 ;
  LAYER M2 ;
        RECT 16.08 12.683 18.48 12.685 ;
  LAYER M2 ;
        RECT 16.08 12.599 18.48 12.601 ;
  LAYER M2 ;
        RECT 16.08 12.515 18.48 12.517 ;
  LAYER M1 ;
        RECT 18.464 9.456 18.496 11.964 ;
  LAYER M1 ;
        RECT 18.4 9.456 18.432 11.964 ;
  LAYER M1 ;
        RECT 18.336 9.456 18.368 11.964 ;
  LAYER M1 ;
        RECT 18.272 9.456 18.304 11.964 ;
  LAYER M1 ;
        RECT 18.208 9.456 18.24 11.964 ;
  LAYER M1 ;
        RECT 18.144 9.456 18.176 11.964 ;
  LAYER M1 ;
        RECT 18.08 9.456 18.112 11.964 ;
  LAYER M1 ;
        RECT 18.016 9.456 18.048 11.964 ;
  LAYER M1 ;
        RECT 17.952 9.456 17.984 11.964 ;
  LAYER M1 ;
        RECT 17.888 9.456 17.92 11.964 ;
  LAYER M1 ;
        RECT 17.824 9.456 17.856 11.964 ;
  LAYER M1 ;
        RECT 17.76 9.456 17.792 11.964 ;
  LAYER M1 ;
        RECT 17.696 9.456 17.728 11.964 ;
  LAYER M1 ;
        RECT 17.632 9.456 17.664 11.964 ;
  LAYER M1 ;
        RECT 17.568 9.456 17.6 11.964 ;
  LAYER M1 ;
        RECT 17.504 9.456 17.536 11.964 ;
  LAYER M1 ;
        RECT 17.44 9.456 17.472 11.964 ;
  LAYER M1 ;
        RECT 17.376 9.456 17.408 11.964 ;
  LAYER M1 ;
        RECT 17.312 9.456 17.344 11.964 ;
  LAYER M1 ;
        RECT 17.248 9.456 17.28 11.964 ;
  LAYER M1 ;
        RECT 17.184 9.456 17.216 11.964 ;
  LAYER M1 ;
        RECT 17.12 9.456 17.152 11.964 ;
  LAYER M1 ;
        RECT 17.056 9.456 17.088 11.964 ;
  LAYER M1 ;
        RECT 16.992 9.456 17.024 11.964 ;
  LAYER M1 ;
        RECT 16.928 9.456 16.96 11.964 ;
  LAYER M1 ;
        RECT 16.864 9.456 16.896 11.964 ;
  LAYER M1 ;
        RECT 16.8 9.456 16.832 11.964 ;
  LAYER M1 ;
        RECT 16.736 9.456 16.768 11.964 ;
  LAYER M1 ;
        RECT 16.672 9.456 16.704 11.964 ;
  LAYER M1 ;
        RECT 16.608 9.456 16.64 11.964 ;
  LAYER M1 ;
        RECT 16.544 9.456 16.576 11.964 ;
  LAYER M1 ;
        RECT 16.48 9.456 16.512 11.964 ;
  LAYER M1 ;
        RECT 16.416 9.456 16.448 11.964 ;
  LAYER M1 ;
        RECT 16.352 9.456 16.384 11.964 ;
  LAYER M1 ;
        RECT 16.288 9.456 16.32 11.964 ;
  LAYER M1 ;
        RECT 16.224 9.456 16.256 11.964 ;
  LAYER M1 ;
        RECT 16.16 9.456 16.192 11.964 ;
  LAYER M2 ;
        RECT 16.044 11.848 18.516 11.88 ;
  LAYER M2 ;
        RECT 16.044 11.784 18.516 11.816 ;
  LAYER M2 ;
        RECT 16.044 11.72 18.516 11.752 ;
  LAYER M2 ;
        RECT 16.044 11.656 18.516 11.688 ;
  LAYER M2 ;
        RECT 16.044 11.592 18.516 11.624 ;
  LAYER M2 ;
        RECT 16.044 11.528 18.516 11.56 ;
  LAYER M2 ;
        RECT 16.044 11.464 18.516 11.496 ;
  LAYER M2 ;
        RECT 16.044 11.4 18.516 11.432 ;
  LAYER M2 ;
        RECT 16.044 11.336 18.516 11.368 ;
  LAYER M2 ;
        RECT 16.044 11.272 18.516 11.304 ;
  LAYER M2 ;
        RECT 16.044 11.208 18.516 11.24 ;
  LAYER M2 ;
        RECT 16.044 11.144 18.516 11.176 ;
  LAYER M2 ;
        RECT 16.044 11.08 18.516 11.112 ;
  LAYER M2 ;
        RECT 16.044 11.016 18.516 11.048 ;
  LAYER M2 ;
        RECT 16.044 10.952 18.516 10.984 ;
  LAYER M2 ;
        RECT 16.044 10.888 18.516 10.92 ;
  LAYER M2 ;
        RECT 16.044 10.824 18.516 10.856 ;
  LAYER M2 ;
        RECT 16.044 10.76 18.516 10.792 ;
  LAYER M2 ;
        RECT 16.044 10.696 18.516 10.728 ;
  LAYER M2 ;
        RECT 16.044 10.632 18.516 10.664 ;
  LAYER M2 ;
        RECT 16.044 10.568 18.516 10.6 ;
  LAYER M2 ;
        RECT 16.044 10.504 18.516 10.536 ;
  LAYER M2 ;
        RECT 16.044 10.44 18.516 10.472 ;
  LAYER M2 ;
        RECT 16.044 10.376 18.516 10.408 ;
  LAYER M2 ;
        RECT 16.044 10.312 18.516 10.344 ;
  LAYER M2 ;
        RECT 16.044 10.248 18.516 10.28 ;
  LAYER M2 ;
        RECT 16.044 10.184 18.516 10.216 ;
  LAYER M2 ;
        RECT 16.044 10.12 18.516 10.152 ;
  LAYER M2 ;
        RECT 16.044 10.056 18.516 10.088 ;
  LAYER M2 ;
        RECT 16.044 9.992 18.516 10.024 ;
  LAYER M2 ;
        RECT 16.044 9.928 18.516 9.96 ;
  LAYER M2 ;
        RECT 16.044 9.864 18.516 9.896 ;
  LAYER M2 ;
        RECT 16.044 9.8 18.516 9.832 ;
  LAYER M2 ;
        RECT 16.044 9.736 18.516 9.768 ;
  LAYER M2 ;
        RECT 16.044 9.672 18.516 9.704 ;
  LAYER M2 ;
        RECT 16.044 9.608 18.516 9.64 ;
  LAYER M3 ;
        RECT 18.464 9.456 18.496 11.964 ;
  LAYER M3 ;
        RECT 18.4 9.456 18.432 11.964 ;
  LAYER M3 ;
        RECT 18.336 9.456 18.368 11.964 ;
  LAYER M3 ;
        RECT 18.272 9.456 18.304 11.964 ;
  LAYER M3 ;
        RECT 18.208 9.456 18.24 11.964 ;
  LAYER M3 ;
        RECT 18.144 9.456 18.176 11.964 ;
  LAYER M3 ;
        RECT 18.08 9.456 18.112 11.964 ;
  LAYER M3 ;
        RECT 18.016 9.456 18.048 11.964 ;
  LAYER M3 ;
        RECT 17.952 9.456 17.984 11.964 ;
  LAYER M3 ;
        RECT 17.888 9.456 17.92 11.964 ;
  LAYER M3 ;
        RECT 17.824 9.456 17.856 11.964 ;
  LAYER M3 ;
        RECT 17.76 9.456 17.792 11.964 ;
  LAYER M3 ;
        RECT 17.696 9.456 17.728 11.964 ;
  LAYER M3 ;
        RECT 17.632 9.456 17.664 11.964 ;
  LAYER M3 ;
        RECT 17.568 9.456 17.6 11.964 ;
  LAYER M3 ;
        RECT 17.504 9.456 17.536 11.964 ;
  LAYER M3 ;
        RECT 17.44 9.456 17.472 11.964 ;
  LAYER M3 ;
        RECT 17.376 9.456 17.408 11.964 ;
  LAYER M3 ;
        RECT 17.312 9.456 17.344 11.964 ;
  LAYER M3 ;
        RECT 17.248 9.456 17.28 11.964 ;
  LAYER M3 ;
        RECT 17.184 9.456 17.216 11.964 ;
  LAYER M3 ;
        RECT 17.12 9.456 17.152 11.964 ;
  LAYER M3 ;
        RECT 17.056 9.456 17.088 11.964 ;
  LAYER M3 ;
        RECT 16.992 9.456 17.024 11.964 ;
  LAYER M3 ;
        RECT 16.928 9.456 16.96 11.964 ;
  LAYER M3 ;
        RECT 16.864 9.456 16.896 11.964 ;
  LAYER M3 ;
        RECT 16.8 9.456 16.832 11.964 ;
  LAYER M3 ;
        RECT 16.736 9.456 16.768 11.964 ;
  LAYER M3 ;
        RECT 16.672 9.456 16.704 11.964 ;
  LAYER M3 ;
        RECT 16.608 9.456 16.64 11.964 ;
  LAYER M3 ;
        RECT 16.544 9.456 16.576 11.964 ;
  LAYER M3 ;
        RECT 16.48 9.456 16.512 11.964 ;
  LAYER M3 ;
        RECT 16.416 9.456 16.448 11.964 ;
  LAYER M3 ;
        RECT 16.352 9.456 16.384 11.964 ;
  LAYER M3 ;
        RECT 16.288 9.456 16.32 11.964 ;
  LAYER M3 ;
        RECT 16.224 9.456 16.256 11.964 ;
  LAYER M3 ;
        RECT 16.16 9.456 16.192 11.964 ;
  LAYER M3 ;
        RECT 16.064 9.456 16.096 11.964 ;
  LAYER M1 ;
        RECT 18.479 9.492 18.481 11.928 ;
  LAYER M1 ;
        RECT 18.399 9.492 18.401 11.928 ;
  LAYER M1 ;
        RECT 18.319 9.492 18.321 11.928 ;
  LAYER M1 ;
        RECT 18.239 9.492 18.241 11.928 ;
  LAYER M1 ;
        RECT 18.159 9.492 18.161 11.928 ;
  LAYER M1 ;
        RECT 18.079 9.492 18.081 11.928 ;
  LAYER M1 ;
        RECT 17.999 9.492 18.001 11.928 ;
  LAYER M1 ;
        RECT 17.919 9.492 17.921 11.928 ;
  LAYER M1 ;
        RECT 17.839 9.492 17.841 11.928 ;
  LAYER M1 ;
        RECT 17.759 9.492 17.761 11.928 ;
  LAYER M1 ;
        RECT 17.679 9.492 17.681 11.928 ;
  LAYER M1 ;
        RECT 17.599 9.492 17.601 11.928 ;
  LAYER M1 ;
        RECT 17.519 9.492 17.521 11.928 ;
  LAYER M1 ;
        RECT 17.439 9.492 17.441 11.928 ;
  LAYER M1 ;
        RECT 17.359 9.492 17.361 11.928 ;
  LAYER M1 ;
        RECT 17.279 9.492 17.281 11.928 ;
  LAYER M1 ;
        RECT 17.199 9.492 17.201 11.928 ;
  LAYER M1 ;
        RECT 17.119 9.492 17.121 11.928 ;
  LAYER M1 ;
        RECT 17.039 9.492 17.041 11.928 ;
  LAYER M1 ;
        RECT 16.959 9.492 16.961 11.928 ;
  LAYER M1 ;
        RECT 16.879 9.492 16.881 11.928 ;
  LAYER M1 ;
        RECT 16.799 9.492 16.801 11.928 ;
  LAYER M1 ;
        RECT 16.719 9.492 16.721 11.928 ;
  LAYER M1 ;
        RECT 16.639 9.492 16.641 11.928 ;
  LAYER M1 ;
        RECT 16.559 9.492 16.561 11.928 ;
  LAYER M1 ;
        RECT 16.479 9.492 16.481 11.928 ;
  LAYER M1 ;
        RECT 16.399 9.492 16.401 11.928 ;
  LAYER M1 ;
        RECT 16.319 9.492 16.321 11.928 ;
  LAYER M1 ;
        RECT 16.239 9.492 16.241 11.928 ;
  LAYER M1 ;
        RECT 16.159 9.492 16.161 11.928 ;
  LAYER M2 ;
        RECT 16.08 11.927 18.48 11.929 ;
  LAYER M2 ;
        RECT 16.08 11.843 18.48 11.845 ;
  LAYER M2 ;
        RECT 16.08 11.759 18.48 11.761 ;
  LAYER M2 ;
        RECT 16.08 11.675 18.48 11.677 ;
  LAYER M2 ;
        RECT 16.08 11.591 18.48 11.593 ;
  LAYER M2 ;
        RECT 16.08 11.507 18.48 11.509 ;
  LAYER M2 ;
        RECT 16.08 11.423 18.48 11.425 ;
  LAYER M2 ;
        RECT 16.08 11.339 18.48 11.341 ;
  LAYER M2 ;
        RECT 16.08 11.255 18.48 11.257 ;
  LAYER M2 ;
        RECT 16.08 11.171 18.48 11.173 ;
  LAYER M2 ;
        RECT 16.08 11.087 18.48 11.089 ;
  LAYER M2 ;
        RECT 16.08 11.003 18.48 11.005 ;
  LAYER M2 ;
        RECT 16.08 10.9195 18.48 10.9215 ;
  LAYER M2 ;
        RECT 16.08 10.835 18.48 10.837 ;
  LAYER M2 ;
        RECT 16.08 10.751 18.48 10.753 ;
  LAYER M2 ;
        RECT 16.08 10.667 18.48 10.669 ;
  LAYER M2 ;
        RECT 16.08 10.583 18.48 10.585 ;
  LAYER M2 ;
        RECT 16.08 10.499 18.48 10.501 ;
  LAYER M2 ;
        RECT 16.08 10.415 18.48 10.417 ;
  LAYER M2 ;
        RECT 16.08 10.331 18.48 10.333 ;
  LAYER M2 ;
        RECT 16.08 10.247 18.48 10.249 ;
  LAYER M2 ;
        RECT 16.08 10.163 18.48 10.165 ;
  LAYER M2 ;
        RECT 16.08 10.079 18.48 10.081 ;
  LAYER M2 ;
        RECT 16.08 9.995 18.48 9.997 ;
  LAYER M2 ;
        RECT 16.08 9.911 18.48 9.913 ;
  LAYER M2 ;
        RECT 16.08 9.827 18.48 9.829 ;
  LAYER M2 ;
        RECT 16.08 9.743 18.48 9.745 ;
  LAYER M2 ;
        RECT 16.08 9.659 18.48 9.661 ;
  LAYER M2 ;
        RECT 16.08 9.575 18.48 9.577 ;
  LAYER M1 ;
        RECT 18.464 6.516 18.496 9.024 ;
  LAYER M1 ;
        RECT 18.4 6.516 18.432 9.024 ;
  LAYER M1 ;
        RECT 18.336 6.516 18.368 9.024 ;
  LAYER M1 ;
        RECT 18.272 6.516 18.304 9.024 ;
  LAYER M1 ;
        RECT 18.208 6.516 18.24 9.024 ;
  LAYER M1 ;
        RECT 18.144 6.516 18.176 9.024 ;
  LAYER M1 ;
        RECT 18.08 6.516 18.112 9.024 ;
  LAYER M1 ;
        RECT 18.016 6.516 18.048 9.024 ;
  LAYER M1 ;
        RECT 17.952 6.516 17.984 9.024 ;
  LAYER M1 ;
        RECT 17.888 6.516 17.92 9.024 ;
  LAYER M1 ;
        RECT 17.824 6.516 17.856 9.024 ;
  LAYER M1 ;
        RECT 17.76 6.516 17.792 9.024 ;
  LAYER M1 ;
        RECT 17.696 6.516 17.728 9.024 ;
  LAYER M1 ;
        RECT 17.632 6.516 17.664 9.024 ;
  LAYER M1 ;
        RECT 17.568 6.516 17.6 9.024 ;
  LAYER M1 ;
        RECT 17.504 6.516 17.536 9.024 ;
  LAYER M1 ;
        RECT 17.44 6.516 17.472 9.024 ;
  LAYER M1 ;
        RECT 17.376 6.516 17.408 9.024 ;
  LAYER M1 ;
        RECT 17.312 6.516 17.344 9.024 ;
  LAYER M1 ;
        RECT 17.248 6.516 17.28 9.024 ;
  LAYER M1 ;
        RECT 17.184 6.516 17.216 9.024 ;
  LAYER M1 ;
        RECT 17.12 6.516 17.152 9.024 ;
  LAYER M1 ;
        RECT 17.056 6.516 17.088 9.024 ;
  LAYER M1 ;
        RECT 16.992 6.516 17.024 9.024 ;
  LAYER M1 ;
        RECT 16.928 6.516 16.96 9.024 ;
  LAYER M1 ;
        RECT 16.864 6.516 16.896 9.024 ;
  LAYER M1 ;
        RECT 16.8 6.516 16.832 9.024 ;
  LAYER M1 ;
        RECT 16.736 6.516 16.768 9.024 ;
  LAYER M1 ;
        RECT 16.672 6.516 16.704 9.024 ;
  LAYER M1 ;
        RECT 16.608 6.516 16.64 9.024 ;
  LAYER M1 ;
        RECT 16.544 6.516 16.576 9.024 ;
  LAYER M1 ;
        RECT 16.48 6.516 16.512 9.024 ;
  LAYER M1 ;
        RECT 16.416 6.516 16.448 9.024 ;
  LAYER M1 ;
        RECT 16.352 6.516 16.384 9.024 ;
  LAYER M1 ;
        RECT 16.288 6.516 16.32 9.024 ;
  LAYER M1 ;
        RECT 16.224 6.516 16.256 9.024 ;
  LAYER M1 ;
        RECT 16.16 6.516 16.192 9.024 ;
  LAYER M2 ;
        RECT 16.044 8.908 18.516 8.94 ;
  LAYER M2 ;
        RECT 16.044 8.844 18.516 8.876 ;
  LAYER M2 ;
        RECT 16.044 8.78 18.516 8.812 ;
  LAYER M2 ;
        RECT 16.044 8.716 18.516 8.748 ;
  LAYER M2 ;
        RECT 16.044 8.652 18.516 8.684 ;
  LAYER M2 ;
        RECT 16.044 8.588 18.516 8.62 ;
  LAYER M2 ;
        RECT 16.044 8.524 18.516 8.556 ;
  LAYER M2 ;
        RECT 16.044 8.46 18.516 8.492 ;
  LAYER M2 ;
        RECT 16.044 8.396 18.516 8.428 ;
  LAYER M2 ;
        RECT 16.044 8.332 18.516 8.364 ;
  LAYER M2 ;
        RECT 16.044 8.268 18.516 8.3 ;
  LAYER M2 ;
        RECT 16.044 8.204 18.516 8.236 ;
  LAYER M2 ;
        RECT 16.044 8.14 18.516 8.172 ;
  LAYER M2 ;
        RECT 16.044 8.076 18.516 8.108 ;
  LAYER M2 ;
        RECT 16.044 8.012 18.516 8.044 ;
  LAYER M2 ;
        RECT 16.044 7.948 18.516 7.98 ;
  LAYER M2 ;
        RECT 16.044 7.884 18.516 7.916 ;
  LAYER M2 ;
        RECT 16.044 7.82 18.516 7.852 ;
  LAYER M2 ;
        RECT 16.044 7.756 18.516 7.788 ;
  LAYER M2 ;
        RECT 16.044 7.692 18.516 7.724 ;
  LAYER M2 ;
        RECT 16.044 7.628 18.516 7.66 ;
  LAYER M2 ;
        RECT 16.044 7.564 18.516 7.596 ;
  LAYER M2 ;
        RECT 16.044 7.5 18.516 7.532 ;
  LAYER M2 ;
        RECT 16.044 7.436 18.516 7.468 ;
  LAYER M2 ;
        RECT 16.044 7.372 18.516 7.404 ;
  LAYER M2 ;
        RECT 16.044 7.308 18.516 7.34 ;
  LAYER M2 ;
        RECT 16.044 7.244 18.516 7.276 ;
  LAYER M2 ;
        RECT 16.044 7.18 18.516 7.212 ;
  LAYER M2 ;
        RECT 16.044 7.116 18.516 7.148 ;
  LAYER M2 ;
        RECT 16.044 7.052 18.516 7.084 ;
  LAYER M2 ;
        RECT 16.044 6.988 18.516 7.02 ;
  LAYER M2 ;
        RECT 16.044 6.924 18.516 6.956 ;
  LAYER M2 ;
        RECT 16.044 6.86 18.516 6.892 ;
  LAYER M2 ;
        RECT 16.044 6.796 18.516 6.828 ;
  LAYER M2 ;
        RECT 16.044 6.732 18.516 6.764 ;
  LAYER M2 ;
        RECT 16.044 6.668 18.516 6.7 ;
  LAYER M3 ;
        RECT 18.464 6.516 18.496 9.024 ;
  LAYER M3 ;
        RECT 18.4 6.516 18.432 9.024 ;
  LAYER M3 ;
        RECT 18.336 6.516 18.368 9.024 ;
  LAYER M3 ;
        RECT 18.272 6.516 18.304 9.024 ;
  LAYER M3 ;
        RECT 18.208 6.516 18.24 9.024 ;
  LAYER M3 ;
        RECT 18.144 6.516 18.176 9.024 ;
  LAYER M3 ;
        RECT 18.08 6.516 18.112 9.024 ;
  LAYER M3 ;
        RECT 18.016 6.516 18.048 9.024 ;
  LAYER M3 ;
        RECT 17.952 6.516 17.984 9.024 ;
  LAYER M3 ;
        RECT 17.888 6.516 17.92 9.024 ;
  LAYER M3 ;
        RECT 17.824 6.516 17.856 9.024 ;
  LAYER M3 ;
        RECT 17.76 6.516 17.792 9.024 ;
  LAYER M3 ;
        RECT 17.696 6.516 17.728 9.024 ;
  LAYER M3 ;
        RECT 17.632 6.516 17.664 9.024 ;
  LAYER M3 ;
        RECT 17.568 6.516 17.6 9.024 ;
  LAYER M3 ;
        RECT 17.504 6.516 17.536 9.024 ;
  LAYER M3 ;
        RECT 17.44 6.516 17.472 9.024 ;
  LAYER M3 ;
        RECT 17.376 6.516 17.408 9.024 ;
  LAYER M3 ;
        RECT 17.312 6.516 17.344 9.024 ;
  LAYER M3 ;
        RECT 17.248 6.516 17.28 9.024 ;
  LAYER M3 ;
        RECT 17.184 6.516 17.216 9.024 ;
  LAYER M3 ;
        RECT 17.12 6.516 17.152 9.024 ;
  LAYER M3 ;
        RECT 17.056 6.516 17.088 9.024 ;
  LAYER M3 ;
        RECT 16.992 6.516 17.024 9.024 ;
  LAYER M3 ;
        RECT 16.928 6.516 16.96 9.024 ;
  LAYER M3 ;
        RECT 16.864 6.516 16.896 9.024 ;
  LAYER M3 ;
        RECT 16.8 6.516 16.832 9.024 ;
  LAYER M3 ;
        RECT 16.736 6.516 16.768 9.024 ;
  LAYER M3 ;
        RECT 16.672 6.516 16.704 9.024 ;
  LAYER M3 ;
        RECT 16.608 6.516 16.64 9.024 ;
  LAYER M3 ;
        RECT 16.544 6.516 16.576 9.024 ;
  LAYER M3 ;
        RECT 16.48 6.516 16.512 9.024 ;
  LAYER M3 ;
        RECT 16.416 6.516 16.448 9.024 ;
  LAYER M3 ;
        RECT 16.352 6.516 16.384 9.024 ;
  LAYER M3 ;
        RECT 16.288 6.516 16.32 9.024 ;
  LAYER M3 ;
        RECT 16.224 6.516 16.256 9.024 ;
  LAYER M3 ;
        RECT 16.16 6.516 16.192 9.024 ;
  LAYER M3 ;
        RECT 16.064 6.516 16.096 9.024 ;
  LAYER M1 ;
        RECT 18.479 6.552 18.481 8.988 ;
  LAYER M1 ;
        RECT 18.399 6.552 18.401 8.988 ;
  LAYER M1 ;
        RECT 18.319 6.552 18.321 8.988 ;
  LAYER M1 ;
        RECT 18.239 6.552 18.241 8.988 ;
  LAYER M1 ;
        RECT 18.159 6.552 18.161 8.988 ;
  LAYER M1 ;
        RECT 18.079 6.552 18.081 8.988 ;
  LAYER M1 ;
        RECT 17.999 6.552 18.001 8.988 ;
  LAYER M1 ;
        RECT 17.919 6.552 17.921 8.988 ;
  LAYER M1 ;
        RECT 17.839 6.552 17.841 8.988 ;
  LAYER M1 ;
        RECT 17.759 6.552 17.761 8.988 ;
  LAYER M1 ;
        RECT 17.679 6.552 17.681 8.988 ;
  LAYER M1 ;
        RECT 17.599 6.552 17.601 8.988 ;
  LAYER M1 ;
        RECT 17.519 6.552 17.521 8.988 ;
  LAYER M1 ;
        RECT 17.439 6.552 17.441 8.988 ;
  LAYER M1 ;
        RECT 17.359 6.552 17.361 8.988 ;
  LAYER M1 ;
        RECT 17.279 6.552 17.281 8.988 ;
  LAYER M1 ;
        RECT 17.199 6.552 17.201 8.988 ;
  LAYER M1 ;
        RECT 17.119 6.552 17.121 8.988 ;
  LAYER M1 ;
        RECT 17.039 6.552 17.041 8.988 ;
  LAYER M1 ;
        RECT 16.959 6.552 16.961 8.988 ;
  LAYER M1 ;
        RECT 16.879 6.552 16.881 8.988 ;
  LAYER M1 ;
        RECT 16.799 6.552 16.801 8.988 ;
  LAYER M1 ;
        RECT 16.719 6.552 16.721 8.988 ;
  LAYER M1 ;
        RECT 16.639 6.552 16.641 8.988 ;
  LAYER M1 ;
        RECT 16.559 6.552 16.561 8.988 ;
  LAYER M1 ;
        RECT 16.479 6.552 16.481 8.988 ;
  LAYER M1 ;
        RECT 16.399 6.552 16.401 8.988 ;
  LAYER M1 ;
        RECT 16.319 6.552 16.321 8.988 ;
  LAYER M1 ;
        RECT 16.239 6.552 16.241 8.988 ;
  LAYER M1 ;
        RECT 16.159 6.552 16.161 8.988 ;
  LAYER M2 ;
        RECT 16.08 8.987 18.48 8.989 ;
  LAYER M2 ;
        RECT 16.08 8.903 18.48 8.905 ;
  LAYER M2 ;
        RECT 16.08 8.819 18.48 8.821 ;
  LAYER M2 ;
        RECT 16.08 8.735 18.48 8.737 ;
  LAYER M2 ;
        RECT 16.08 8.651 18.48 8.653 ;
  LAYER M2 ;
        RECT 16.08 8.567 18.48 8.569 ;
  LAYER M2 ;
        RECT 16.08 8.483 18.48 8.485 ;
  LAYER M2 ;
        RECT 16.08 8.399 18.48 8.401 ;
  LAYER M2 ;
        RECT 16.08 8.315 18.48 8.317 ;
  LAYER M2 ;
        RECT 16.08 8.231 18.48 8.233 ;
  LAYER M2 ;
        RECT 16.08 8.147 18.48 8.149 ;
  LAYER M2 ;
        RECT 16.08 8.063 18.48 8.065 ;
  LAYER M2 ;
        RECT 16.08 7.9795 18.48 7.9815 ;
  LAYER M2 ;
        RECT 16.08 7.895 18.48 7.897 ;
  LAYER M2 ;
        RECT 16.08 7.811 18.48 7.813 ;
  LAYER M2 ;
        RECT 16.08 7.727 18.48 7.729 ;
  LAYER M2 ;
        RECT 16.08 7.643 18.48 7.645 ;
  LAYER M2 ;
        RECT 16.08 7.559 18.48 7.561 ;
  LAYER M2 ;
        RECT 16.08 7.475 18.48 7.477 ;
  LAYER M2 ;
        RECT 16.08 7.391 18.48 7.393 ;
  LAYER M2 ;
        RECT 16.08 7.307 18.48 7.309 ;
  LAYER M2 ;
        RECT 16.08 7.223 18.48 7.225 ;
  LAYER M2 ;
        RECT 16.08 7.139 18.48 7.141 ;
  LAYER M2 ;
        RECT 16.08 7.055 18.48 7.057 ;
  LAYER M2 ;
        RECT 16.08 6.971 18.48 6.973 ;
  LAYER M2 ;
        RECT 16.08 6.887 18.48 6.889 ;
  LAYER M2 ;
        RECT 16.08 6.803 18.48 6.805 ;
  LAYER M2 ;
        RECT 16.08 6.719 18.48 6.721 ;
  LAYER M2 ;
        RECT 16.08 6.635 18.48 6.637 ;
  LAYER M1 ;
        RECT 21.824 30.96 21.856 31.032 ;
  LAYER M2 ;
        RECT 21.804 30.98 21.876 31.012 ;
  LAYER M2 ;
        RECT 21.52 30.98 21.84 31.012 ;
  LAYER M1 ;
        RECT 21.504 30.96 21.536 31.032 ;
  LAYER M2 ;
        RECT 21.484 30.98 21.556 31.012 ;
  LAYER M1 ;
        RECT 21.824 28.02 21.856 28.092 ;
  LAYER M2 ;
        RECT 21.804 28.04 21.876 28.072 ;
  LAYER M2 ;
        RECT 21.52 28.04 21.84 28.072 ;
  LAYER M1 ;
        RECT 21.504 28.02 21.536 28.092 ;
  LAYER M2 ;
        RECT 21.484 28.04 21.556 28.072 ;
  LAYER M1 ;
        RECT 18.944 30.96 18.976 31.032 ;
  LAYER M2 ;
        RECT 18.924 30.98 18.996 31.012 ;
  LAYER M1 ;
        RECT 18.944 30.996 18.976 31.164 ;
  LAYER M1 ;
        RECT 18.944 31.128 18.976 31.2 ;
  LAYER M2 ;
        RECT 18.924 31.148 18.996 31.18 ;
  LAYER M2 ;
        RECT 18.96 31.148 21.52 31.18 ;
  LAYER M1 ;
        RECT 21.504 31.128 21.536 31.2 ;
  LAYER M2 ;
        RECT 21.484 31.148 21.556 31.18 ;
  LAYER M1 ;
        RECT 18.944 28.02 18.976 28.092 ;
  LAYER M2 ;
        RECT 18.924 28.04 18.996 28.072 ;
  LAYER M1 ;
        RECT 18.944 28.056 18.976 28.224 ;
  LAYER M1 ;
        RECT 18.944 28.188 18.976 28.26 ;
  LAYER M2 ;
        RECT 18.924 28.208 18.996 28.24 ;
  LAYER M2 ;
        RECT 18.96 28.208 21.52 28.24 ;
  LAYER M1 ;
        RECT 21.504 28.188 21.536 28.26 ;
  LAYER M2 ;
        RECT 21.484 28.208 21.556 28.24 ;
  LAYER M1 ;
        RECT 21.504 37.344 21.536 37.416 ;
  LAYER M2 ;
        RECT 21.484 37.364 21.556 37.396 ;
  LAYER M1 ;
        RECT 21.504 37.212 21.536 37.38 ;
  LAYER M1 ;
        RECT 21.504 28.056 21.536 37.212 ;
  LAYER M1 ;
        RECT 24.704 28.02 24.736 28.092 ;
  LAYER M2 ;
        RECT 24.684 28.04 24.756 28.072 ;
  LAYER M2 ;
        RECT 24.4 28.04 24.72 28.072 ;
  LAYER M1 ;
        RECT 24.384 28.02 24.416 28.092 ;
  LAYER M2 ;
        RECT 24.364 28.04 24.436 28.072 ;
  LAYER M1 ;
        RECT 24.704 30.96 24.736 31.032 ;
  LAYER M2 ;
        RECT 24.684 30.98 24.756 31.012 ;
  LAYER M2 ;
        RECT 24.4 30.98 24.72 31.012 ;
  LAYER M1 ;
        RECT 24.384 30.96 24.416 31.032 ;
  LAYER M2 ;
        RECT 24.364 30.98 24.436 31.012 ;
  LAYER M1 ;
        RECT 24.384 37.344 24.416 37.416 ;
  LAYER M2 ;
        RECT 24.364 37.364 24.436 37.396 ;
  LAYER M1 ;
        RECT 24.384 37.212 24.416 37.38 ;
  LAYER M1 ;
        RECT 24.384 28.056 24.416 37.212 ;
  LAYER M2 ;
        RECT 21.52 37.364 24.4 37.396 ;
  LAYER M1 ;
        RECT 18.944 25.08 18.976 25.152 ;
  LAYER M2 ;
        RECT 18.924 25.1 18.996 25.132 ;
  LAYER M2 ;
        RECT 18.64 25.1 18.96 25.132 ;
  LAYER M1 ;
        RECT 18.624 25.08 18.656 25.152 ;
  LAYER M2 ;
        RECT 18.604 25.1 18.676 25.132 ;
  LAYER M1 ;
        RECT 18.944 33.9 18.976 33.972 ;
  LAYER M2 ;
        RECT 18.924 33.92 18.996 33.952 ;
  LAYER M2 ;
        RECT 18.64 33.92 18.96 33.952 ;
  LAYER M1 ;
        RECT 18.624 33.9 18.656 33.972 ;
  LAYER M2 ;
        RECT 18.604 33.92 18.676 33.952 ;
  LAYER M1 ;
        RECT 18.624 37.512 18.656 37.584 ;
  LAYER M2 ;
        RECT 18.604 37.532 18.676 37.564 ;
  LAYER M1 ;
        RECT 18.624 37.212 18.656 37.548 ;
  LAYER M1 ;
        RECT 18.624 25.116 18.656 37.212 ;
  LAYER M1 ;
        RECT 24.704 33.9 24.736 33.972 ;
  LAYER M2 ;
        RECT 24.684 33.92 24.756 33.952 ;
  LAYER M1 ;
        RECT 24.704 33.936 24.736 34.104 ;
  LAYER M1 ;
        RECT 24.704 34.068 24.736 34.14 ;
  LAYER M2 ;
        RECT 24.684 34.088 24.756 34.12 ;
  LAYER M2 ;
        RECT 24.72 34.088 27.28 34.12 ;
  LAYER M1 ;
        RECT 27.264 34.068 27.296 34.14 ;
  LAYER M2 ;
        RECT 27.244 34.088 27.316 34.12 ;
  LAYER M1 ;
        RECT 24.704 25.08 24.736 25.152 ;
  LAYER M2 ;
        RECT 24.684 25.1 24.756 25.132 ;
  LAYER M1 ;
        RECT 24.704 25.116 24.736 25.284 ;
  LAYER M1 ;
        RECT 24.704 25.248 24.736 25.32 ;
  LAYER M2 ;
        RECT 24.684 25.268 24.756 25.3 ;
  LAYER M2 ;
        RECT 24.72 25.268 27.28 25.3 ;
  LAYER M1 ;
        RECT 27.264 25.248 27.296 25.32 ;
  LAYER M2 ;
        RECT 27.244 25.268 27.316 25.3 ;
  LAYER M1 ;
        RECT 27.264 37.512 27.296 37.584 ;
  LAYER M2 ;
        RECT 27.244 37.532 27.316 37.564 ;
  LAYER M1 ;
        RECT 27.264 37.212 27.296 37.548 ;
  LAYER M1 ;
        RECT 27.264 25.284 27.296 37.212 ;
  LAYER M2 ;
        RECT 18.64 37.532 27.28 37.564 ;
  LAYER M1 ;
        RECT 21.824 33.9 21.856 33.972 ;
  LAYER M2 ;
        RECT 21.804 33.92 21.876 33.952 ;
  LAYER M2 ;
        RECT 21.84 33.92 24.72 33.952 ;
  LAYER M1 ;
        RECT 24.704 33.9 24.736 33.972 ;
  LAYER M2 ;
        RECT 24.684 33.92 24.756 33.952 ;
  LAYER M1 ;
        RECT 21.824 25.08 21.856 25.152 ;
  LAYER M2 ;
        RECT 21.804 25.1 21.876 25.132 ;
  LAYER M2 ;
        RECT 18.96 25.1 21.84 25.132 ;
  LAYER M1 ;
        RECT 18.944 25.08 18.976 25.152 ;
  LAYER M2 ;
        RECT 18.924 25.1 18.996 25.132 ;
  LAYER M1 ;
        RECT 16.064 36.84 16.096 36.912 ;
  LAYER M2 ;
        RECT 16.044 36.86 16.116 36.892 ;
  LAYER M2 ;
        RECT 15.76 36.86 16.08 36.892 ;
  LAYER M1 ;
        RECT 15.744 36.84 15.776 36.912 ;
  LAYER M2 ;
        RECT 15.724 36.86 15.796 36.892 ;
  LAYER M1 ;
        RECT 16.064 33.9 16.096 33.972 ;
  LAYER M2 ;
        RECT 16.044 33.92 16.116 33.952 ;
  LAYER M2 ;
        RECT 15.76 33.92 16.08 33.952 ;
  LAYER M1 ;
        RECT 15.744 33.9 15.776 33.972 ;
  LAYER M2 ;
        RECT 15.724 33.92 15.796 33.952 ;
  LAYER M1 ;
        RECT 16.064 30.96 16.096 31.032 ;
  LAYER M2 ;
        RECT 16.044 30.98 16.116 31.012 ;
  LAYER M2 ;
        RECT 15.76 30.98 16.08 31.012 ;
  LAYER M1 ;
        RECT 15.744 30.96 15.776 31.032 ;
  LAYER M2 ;
        RECT 15.724 30.98 15.796 31.012 ;
  LAYER M1 ;
        RECT 16.064 28.02 16.096 28.092 ;
  LAYER M2 ;
        RECT 16.044 28.04 16.116 28.072 ;
  LAYER M2 ;
        RECT 15.76 28.04 16.08 28.072 ;
  LAYER M1 ;
        RECT 15.744 28.02 15.776 28.092 ;
  LAYER M2 ;
        RECT 15.724 28.04 15.796 28.072 ;
  LAYER M1 ;
        RECT 16.064 25.08 16.096 25.152 ;
  LAYER M2 ;
        RECT 16.044 25.1 16.116 25.132 ;
  LAYER M2 ;
        RECT 15.76 25.1 16.08 25.132 ;
  LAYER M1 ;
        RECT 15.744 25.08 15.776 25.152 ;
  LAYER M2 ;
        RECT 15.724 25.1 15.796 25.132 ;
  LAYER M1 ;
        RECT 16.064 22.14 16.096 22.212 ;
  LAYER M2 ;
        RECT 16.044 22.16 16.116 22.192 ;
  LAYER M2 ;
        RECT 15.76 22.16 16.08 22.192 ;
  LAYER M1 ;
        RECT 15.744 22.14 15.776 22.212 ;
  LAYER M2 ;
        RECT 15.724 22.16 15.796 22.192 ;
  LAYER M1 ;
        RECT 15.744 37.68 15.776 37.752 ;
  LAYER M2 ;
        RECT 15.724 37.7 15.796 37.732 ;
  LAYER M1 ;
        RECT 15.744 37.212 15.776 37.716 ;
  LAYER M1 ;
        RECT 15.744 22.176 15.776 37.212 ;
  LAYER M1 ;
        RECT 27.584 36.84 27.616 36.912 ;
  LAYER M2 ;
        RECT 27.564 36.86 27.636 36.892 ;
  LAYER M1 ;
        RECT 27.584 36.876 27.616 37.044 ;
  LAYER M1 ;
        RECT 27.584 37.008 27.616 37.08 ;
  LAYER M2 ;
        RECT 27.564 37.028 27.636 37.06 ;
  LAYER M2 ;
        RECT 27.6 37.028 30.16 37.06 ;
  LAYER M1 ;
        RECT 30.144 37.008 30.176 37.08 ;
  LAYER M2 ;
        RECT 30.124 37.028 30.196 37.06 ;
  LAYER M1 ;
        RECT 27.584 33.9 27.616 33.972 ;
  LAYER M2 ;
        RECT 27.564 33.92 27.636 33.952 ;
  LAYER M1 ;
        RECT 27.584 33.936 27.616 34.104 ;
  LAYER M1 ;
        RECT 27.584 34.068 27.616 34.14 ;
  LAYER M2 ;
        RECT 27.564 34.088 27.636 34.12 ;
  LAYER M2 ;
        RECT 27.6 34.088 30.16 34.12 ;
  LAYER M1 ;
        RECT 30.144 34.068 30.176 34.14 ;
  LAYER M2 ;
        RECT 30.124 34.088 30.196 34.12 ;
  LAYER M1 ;
        RECT 27.584 30.96 27.616 31.032 ;
  LAYER M2 ;
        RECT 27.564 30.98 27.636 31.012 ;
  LAYER M1 ;
        RECT 27.584 30.996 27.616 31.164 ;
  LAYER M1 ;
        RECT 27.584 31.128 27.616 31.2 ;
  LAYER M2 ;
        RECT 27.564 31.148 27.636 31.18 ;
  LAYER M2 ;
        RECT 27.6 31.148 30.16 31.18 ;
  LAYER M1 ;
        RECT 30.144 31.128 30.176 31.2 ;
  LAYER M2 ;
        RECT 30.124 31.148 30.196 31.18 ;
  LAYER M1 ;
        RECT 27.584 28.02 27.616 28.092 ;
  LAYER M2 ;
        RECT 27.564 28.04 27.636 28.072 ;
  LAYER M1 ;
        RECT 27.584 28.056 27.616 28.224 ;
  LAYER M1 ;
        RECT 27.584 28.188 27.616 28.26 ;
  LAYER M2 ;
        RECT 27.564 28.208 27.636 28.24 ;
  LAYER M2 ;
        RECT 27.6 28.208 30.16 28.24 ;
  LAYER M1 ;
        RECT 30.144 28.188 30.176 28.26 ;
  LAYER M2 ;
        RECT 30.124 28.208 30.196 28.24 ;
  LAYER M1 ;
        RECT 27.584 25.08 27.616 25.152 ;
  LAYER M2 ;
        RECT 27.564 25.1 27.636 25.132 ;
  LAYER M1 ;
        RECT 27.584 25.116 27.616 25.284 ;
  LAYER M1 ;
        RECT 27.584 25.248 27.616 25.32 ;
  LAYER M2 ;
        RECT 27.564 25.268 27.636 25.3 ;
  LAYER M2 ;
        RECT 27.6 25.268 30.16 25.3 ;
  LAYER M1 ;
        RECT 30.144 25.248 30.176 25.32 ;
  LAYER M2 ;
        RECT 30.124 25.268 30.196 25.3 ;
  LAYER M1 ;
        RECT 27.584 22.14 27.616 22.212 ;
  LAYER M2 ;
        RECT 27.564 22.16 27.636 22.192 ;
  LAYER M1 ;
        RECT 27.584 22.176 27.616 22.344 ;
  LAYER M1 ;
        RECT 27.584 22.308 27.616 22.38 ;
  LAYER M2 ;
        RECT 27.564 22.328 27.636 22.36 ;
  LAYER M2 ;
        RECT 27.6 22.328 30.16 22.36 ;
  LAYER M1 ;
        RECT 30.144 22.308 30.176 22.38 ;
  LAYER M2 ;
        RECT 30.124 22.328 30.196 22.36 ;
  LAYER M1 ;
        RECT 30.144 37.68 30.176 37.752 ;
  LAYER M2 ;
        RECT 30.124 37.7 30.196 37.732 ;
  LAYER M1 ;
        RECT 30.144 37.212 30.176 37.716 ;
  LAYER M1 ;
        RECT 30.144 22.344 30.176 37.212 ;
  LAYER M2 ;
        RECT 15.76 37.7 30.16 37.732 ;
  LAYER M1 ;
        RECT 18.944 36.84 18.976 36.912 ;
  LAYER M2 ;
        RECT 18.924 36.86 18.996 36.892 ;
  LAYER M2 ;
        RECT 16.08 36.86 18.96 36.892 ;
  LAYER M1 ;
        RECT 16.064 36.84 16.096 36.912 ;
  LAYER M2 ;
        RECT 16.044 36.86 16.116 36.892 ;
  LAYER M1 ;
        RECT 18.944 22.14 18.976 22.212 ;
  LAYER M2 ;
        RECT 18.924 22.16 18.996 22.192 ;
  LAYER M2 ;
        RECT 16.08 22.16 18.96 22.192 ;
  LAYER M1 ;
        RECT 16.064 22.14 16.096 22.212 ;
  LAYER M2 ;
        RECT 16.044 22.16 16.116 22.192 ;
  LAYER M1 ;
        RECT 21.824 22.14 21.856 22.212 ;
  LAYER M2 ;
        RECT 21.804 22.16 21.876 22.192 ;
  LAYER M2 ;
        RECT 18.96 22.16 21.84 22.192 ;
  LAYER M1 ;
        RECT 18.944 22.14 18.976 22.212 ;
  LAYER M2 ;
        RECT 18.924 22.16 18.996 22.192 ;
  LAYER M1 ;
        RECT 24.704 22.14 24.736 22.212 ;
  LAYER M2 ;
        RECT 24.684 22.16 24.756 22.192 ;
  LAYER M2 ;
        RECT 21.84 22.16 24.72 22.192 ;
  LAYER M1 ;
        RECT 21.824 22.14 21.856 22.212 ;
  LAYER M2 ;
        RECT 21.804 22.16 21.876 22.192 ;
  LAYER M1 ;
        RECT 24.704 36.84 24.736 36.912 ;
  LAYER M2 ;
        RECT 24.684 36.86 24.756 36.892 ;
  LAYER M2 ;
        RECT 24.72 36.86 27.6 36.892 ;
  LAYER M1 ;
        RECT 27.584 36.84 27.616 36.912 ;
  LAYER M2 ;
        RECT 27.564 36.86 27.636 36.892 ;
  LAYER M1 ;
        RECT 21.824 36.84 21.856 36.912 ;
  LAYER M2 ;
        RECT 21.804 36.86 21.876 36.892 ;
  LAYER M2 ;
        RECT 21.84 36.86 24.72 36.892 ;
  LAYER M1 ;
        RECT 24.704 36.84 24.736 36.912 ;
  LAYER M2 ;
        RECT 24.684 36.86 24.756 36.892 ;
  LAYER M1 ;
        RECT 24.224 28.524 24.256 28.596 ;
  LAYER M2 ;
        RECT 24.204 28.544 24.276 28.576 ;
  LAYER M2 ;
        RECT 21.68 28.544 24.24 28.576 ;
  LAYER M1 ;
        RECT 21.664 28.524 21.696 28.596 ;
  LAYER M2 ;
        RECT 21.644 28.544 21.716 28.576 ;
  LAYER M1 ;
        RECT 24.224 25.584 24.256 25.656 ;
  LAYER M2 ;
        RECT 24.204 25.604 24.276 25.636 ;
  LAYER M2 ;
        RECT 21.68 25.604 24.24 25.636 ;
  LAYER M1 ;
        RECT 21.664 25.584 21.696 25.656 ;
  LAYER M2 ;
        RECT 21.644 25.604 21.716 25.636 ;
  LAYER M1 ;
        RECT 21.344 28.524 21.376 28.596 ;
  LAYER M2 ;
        RECT 21.324 28.544 21.396 28.576 ;
  LAYER M1 ;
        RECT 21.344 28.392 21.376 28.56 ;
  LAYER M1 ;
        RECT 21.344 28.356 21.376 28.428 ;
  LAYER M2 ;
        RECT 21.324 28.376 21.396 28.408 ;
  LAYER M2 ;
        RECT 21.36 28.376 21.68 28.408 ;
  LAYER M1 ;
        RECT 21.664 28.356 21.696 28.428 ;
  LAYER M2 ;
        RECT 21.644 28.376 21.716 28.408 ;
  LAYER M1 ;
        RECT 21.344 25.584 21.376 25.656 ;
  LAYER M2 ;
        RECT 21.324 25.604 21.396 25.636 ;
  LAYER M1 ;
        RECT 21.344 25.452 21.376 25.62 ;
  LAYER M1 ;
        RECT 21.344 25.416 21.376 25.488 ;
  LAYER M2 ;
        RECT 21.324 25.436 21.396 25.468 ;
  LAYER M2 ;
        RECT 21.36 25.436 21.68 25.468 ;
  LAYER M1 ;
        RECT 21.664 25.416 21.696 25.488 ;
  LAYER M2 ;
        RECT 21.644 25.436 21.716 25.468 ;
  LAYER M1 ;
        RECT 21.664 19.2 21.696 19.272 ;
  LAYER M2 ;
        RECT 21.644 19.22 21.716 19.252 ;
  LAYER M1 ;
        RECT 21.664 19.236 21.696 19.404 ;
  LAYER M1 ;
        RECT 21.664 19.404 21.696 28.56 ;
  LAYER M1 ;
        RECT 27.104 25.584 27.136 25.656 ;
  LAYER M2 ;
        RECT 27.084 25.604 27.156 25.636 ;
  LAYER M2 ;
        RECT 24.56 25.604 27.12 25.636 ;
  LAYER M1 ;
        RECT 24.544 25.584 24.576 25.656 ;
  LAYER M2 ;
        RECT 24.524 25.604 24.596 25.636 ;
  LAYER M1 ;
        RECT 27.104 28.524 27.136 28.596 ;
  LAYER M2 ;
        RECT 27.084 28.544 27.156 28.576 ;
  LAYER M2 ;
        RECT 24.56 28.544 27.12 28.576 ;
  LAYER M1 ;
        RECT 24.544 28.524 24.576 28.596 ;
  LAYER M2 ;
        RECT 24.524 28.544 24.596 28.576 ;
  LAYER M1 ;
        RECT 24.544 19.2 24.576 19.272 ;
  LAYER M2 ;
        RECT 24.524 19.22 24.596 19.252 ;
  LAYER M1 ;
        RECT 24.544 19.236 24.576 19.404 ;
  LAYER M1 ;
        RECT 24.544 19.404 24.576 28.56 ;
  LAYER M2 ;
        RECT 21.68 19.22 24.56 19.252 ;
  LAYER M1 ;
        RECT 21.344 22.644 21.376 22.716 ;
  LAYER M2 ;
        RECT 21.324 22.664 21.396 22.696 ;
  LAYER M2 ;
        RECT 18.8 22.664 21.36 22.696 ;
  LAYER M1 ;
        RECT 18.784 22.644 18.816 22.716 ;
  LAYER M2 ;
        RECT 18.764 22.664 18.836 22.696 ;
  LAYER M1 ;
        RECT 21.344 31.464 21.376 31.536 ;
  LAYER M2 ;
        RECT 21.324 31.484 21.396 31.516 ;
  LAYER M2 ;
        RECT 18.8 31.484 21.36 31.516 ;
  LAYER M1 ;
        RECT 18.784 31.464 18.816 31.536 ;
  LAYER M2 ;
        RECT 18.764 31.484 18.836 31.516 ;
  LAYER M1 ;
        RECT 18.784 19.032 18.816 19.104 ;
  LAYER M2 ;
        RECT 18.764 19.052 18.836 19.084 ;
  LAYER M1 ;
        RECT 18.784 19.068 18.816 19.404 ;
  LAYER M1 ;
        RECT 18.784 19.404 18.816 31.5 ;
  LAYER M1 ;
        RECT 27.104 31.464 27.136 31.536 ;
  LAYER M2 ;
        RECT 27.084 31.484 27.156 31.516 ;
  LAYER M1 ;
        RECT 27.104 31.332 27.136 31.5 ;
  LAYER M1 ;
        RECT 27.104 31.296 27.136 31.368 ;
  LAYER M2 ;
        RECT 27.084 31.316 27.156 31.348 ;
  LAYER M2 ;
        RECT 27.12 31.316 27.44 31.348 ;
  LAYER M1 ;
        RECT 27.424 31.296 27.456 31.368 ;
  LAYER M2 ;
        RECT 27.404 31.316 27.476 31.348 ;
  LAYER M1 ;
        RECT 27.104 22.644 27.136 22.716 ;
  LAYER M2 ;
        RECT 27.084 22.664 27.156 22.696 ;
  LAYER M1 ;
        RECT 27.104 22.512 27.136 22.68 ;
  LAYER M1 ;
        RECT 27.104 22.476 27.136 22.548 ;
  LAYER M2 ;
        RECT 27.084 22.496 27.156 22.528 ;
  LAYER M2 ;
        RECT 27.12 22.496 27.44 22.528 ;
  LAYER M1 ;
        RECT 27.424 22.476 27.456 22.548 ;
  LAYER M2 ;
        RECT 27.404 22.496 27.476 22.528 ;
  LAYER M1 ;
        RECT 27.424 19.032 27.456 19.104 ;
  LAYER M2 ;
        RECT 27.404 19.052 27.476 19.084 ;
  LAYER M1 ;
        RECT 27.424 19.068 27.456 19.404 ;
  LAYER M1 ;
        RECT 27.424 19.404 27.456 31.332 ;
  LAYER M2 ;
        RECT 18.8 19.052 27.44 19.084 ;
  LAYER M1 ;
        RECT 24.224 31.464 24.256 31.536 ;
  LAYER M2 ;
        RECT 24.204 31.484 24.276 31.516 ;
  LAYER M2 ;
        RECT 24.24 31.484 27.12 31.516 ;
  LAYER M1 ;
        RECT 27.104 31.464 27.136 31.536 ;
  LAYER M2 ;
        RECT 27.084 31.484 27.156 31.516 ;
  LAYER M1 ;
        RECT 24.224 22.644 24.256 22.716 ;
  LAYER M2 ;
        RECT 24.204 22.664 24.276 22.696 ;
  LAYER M2 ;
        RECT 21.36 22.664 24.24 22.696 ;
  LAYER M1 ;
        RECT 21.344 22.644 21.376 22.716 ;
  LAYER M2 ;
        RECT 21.324 22.664 21.396 22.696 ;
  LAYER M1 ;
        RECT 18.464 34.404 18.496 34.476 ;
  LAYER M2 ;
        RECT 18.444 34.424 18.516 34.456 ;
  LAYER M2 ;
        RECT 15.92 34.424 18.48 34.456 ;
  LAYER M1 ;
        RECT 15.904 34.404 15.936 34.476 ;
  LAYER M2 ;
        RECT 15.884 34.424 15.956 34.456 ;
  LAYER M1 ;
        RECT 18.464 31.464 18.496 31.536 ;
  LAYER M2 ;
        RECT 18.444 31.484 18.516 31.516 ;
  LAYER M2 ;
        RECT 15.92 31.484 18.48 31.516 ;
  LAYER M1 ;
        RECT 15.904 31.464 15.936 31.536 ;
  LAYER M2 ;
        RECT 15.884 31.484 15.956 31.516 ;
  LAYER M1 ;
        RECT 18.464 28.524 18.496 28.596 ;
  LAYER M2 ;
        RECT 18.444 28.544 18.516 28.576 ;
  LAYER M2 ;
        RECT 15.92 28.544 18.48 28.576 ;
  LAYER M1 ;
        RECT 15.904 28.524 15.936 28.596 ;
  LAYER M2 ;
        RECT 15.884 28.544 15.956 28.576 ;
  LAYER M1 ;
        RECT 18.464 25.584 18.496 25.656 ;
  LAYER M2 ;
        RECT 18.444 25.604 18.516 25.636 ;
  LAYER M2 ;
        RECT 15.92 25.604 18.48 25.636 ;
  LAYER M1 ;
        RECT 15.904 25.584 15.936 25.656 ;
  LAYER M2 ;
        RECT 15.884 25.604 15.956 25.636 ;
  LAYER M1 ;
        RECT 18.464 22.644 18.496 22.716 ;
  LAYER M2 ;
        RECT 18.444 22.664 18.516 22.696 ;
  LAYER M2 ;
        RECT 15.92 22.664 18.48 22.696 ;
  LAYER M1 ;
        RECT 15.904 22.644 15.936 22.716 ;
  LAYER M2 ;
        RECT 15.884 22.664 15.956 22.696 ;
  LAYER M1 ;
        RECT 18.464 19.704 18.496 19.776 ;
  LAYER M2 ;
        RECT 18.444 19.724 18.516 19.756 ;
  LAYER M2 ;
        RECT 15.92 19.724 18.48 19.756 ;
  LAYER M1 ;
        RECT 15.904 19.704 15.936 19.776 ;
  LAYER M2 ;
        RECT 15.884 19.724 15.956 19.756 ;
  LAYER M1 ;
        RECT 15.904 18.864 15.936 18.936 ;
  LAYER M2 ;
        RECT 15.884 18.884 15.956 18.916 ;
  LAYER M1 ;
        RECT 15.904 18.9 15.936 19.404 ;
  LAYER M1 ;
        RECT 15.904 19.404 15.936 34.44 ;
  LAYER M1 ;
        RECT 29.984 34.404 30.016 34.476 ;
  LAYER M2 ;
        RECT 29.964 34.424 30.036 34.456 ;
  LAYER M1 ;
        RECT 29.984 34.272 30.016 34.44 ;
  LAYER M1 ;
        RECT 29.984 34.236 30.016 34.308 ;
  LAYER M2 ;
        RECT 29.964 34.256 30.036 34.288 ;
  LAYER M2 ;
        RECT 30 34.256 30.32 34.288 ;
  LAYER M1 ;
        RECT 30.304 34.236 30.336 34.308 ;
  LAYER M2 ;
        RECT 30.284 34.256 30.356 34.288 ;
  LAYER M1 ;
        RECT 29.984 31.464 30.016 31.536 ;
  LAYER M2 ;
        RECT 29.964 31.484 30.036 31.516 ;
  LAYER M1 ;
        RECT 29.984 31.332 30.016 31.5 ;
  LAYER M1 ;
        RECT 29.984 31.296 30.016 31.368 ;
  LAYER M2 ;
        RECT 29.964 31.316 30.036 31.348 ;
  LAYER M2 ;
        RECT 30 31.316 30.32 31.348 ;
  LAYER M1 ;
        RECT 30.304 31.296 30.336 31.368 ;
  LAYER M2 ;
        RECT 30.284 31.316 30.356 31.348 ;
  LAYER M1 ;
        RECT 29.984 28.524 30.016 28.596 ;
  LAYER M2 ;
        RECT 29.964 28.544 30.036 28.576 ;
  LAYER M1 ;
        RECT 29.984 28.392 30.016 28.56 ;
  LAYER M1 ;
        RECT 29.984 28.356 30.016 28.428 ;
  LAYER M2 ;
        RECT 29.964 28.376 30.036 28.408 ;
  LAYER M2 ;
        RECT 30 28.376 30.32 28.408 ;
  LAYER M1 ;
        RECT 30.304 28.356 30.336 28.428 ;
  LAYER M2 ;
        RECT 30.284 28.376 30.356 28.408 ;
  LAYER M1 ;
        RECT 29.984 25.584 30.016 25.656 ;
  LAYER M2 ;
        RECT 29.964 25.604 30.036 25.636 ;
  LAYER M1 ;
        RECT 29.984 25.452 30.016 25.62 ;
  LAYER M1 ;
        RECT 29.984 25.416 30.016 25.488 ;
  LAYER M2 ;
        RECT 29.964 25.436 30.036 25.468 ;
  LAYER M2 ;
        RECT 30 25.436 30.32 25.468 ;
  LAYER M1 ;
        RECT 30.304 25.416 30.336 25.488 ;
  LAYER M2 ;
        RECT 30.284 25.436 30.356 25.468 ;
  LAYER M1 ;
        RECT 29.984 22.644 30.016 22.716 ;
  LAYER M2 ;
        RECT 29.964 22.664 30.036 22.696 ;
  LAYER M1 ;
        RECT 29.984 22.512 30.016 22.68 ;
  LAYER M1 ;
        RECT 29.984 22.476 30.016 22.548 ;
  LAYER M2 ;
        RECT 29.964 22.496 30.036 22.528 ;
  LAYER M2 ;
        RECT 30 22.496 30.32 22.528 ;
  LAYER M1 ;
        RECT 30.304 22.476 30.336 22.548 ;
  LAYER M2 ;
        RECT 30.284 22.496 30.356 22.528 ;
  LAYER M1 ;
        RECT 29.984 19.704 30.016 19.776 ;
  LAYER M2 ;
        RECT 29.964 19.724 30.036 19.756 ;
  LAYER M1 ;
        RECT 29.984 19.572 30.016 19.74 ;
  LAYER M1 ;
        RECT 29.984 19.536 30.016 19.608 ;
  LAYER M2 ;
        RECT 29.964 19.556 30.036 19.588 ;
  LAYER M2 ;
        RECT 30 19.556 30.32 19.588 ;
  LAYER M1 ;
        RECT 30.304 19.536 30.336 19.608 ;
  LAYER M2 ;
        RECT 30.284 19.556 30.356 19.588 ;
  LAYER M1 ;
        RECT 30.304 18.864 30.336 18.936 ;
  LAYER M2 ;
        RECT 30.284 18.884 30.356 18.916 ;
  LAYER M1 ;
        RECT 30.304 18.9 30.336 19.404 ;
  LAYER M1 ;
        RECT 30.304 19.404 30.336 34.272 ;
  LAYER M2 ;
        RECT 15.92 18.884 30.32 18.916 ;
  LAYER M1 ;
        RECT 21.344 34.404 21.376 34.476 ;
  LAYER M2 ;
        RECT 21.324 34.424 21.396 34.456 ;
  LAYER M2 ;
        RECT 18.48 34.424 21.36 34.456 ;
  LAYER M1 ;
        RECT 18.464 34.404 18.496 34.476 ;
  LAYER M2 ;
        RECT 18.444 34.424 18.516 34.456 ;
  LAYER M1 ;
        RECT 21.344 19.704 21.376 19.776 ;
  LAYER M2 ;
        RECT 21.324 19.724 21.396 19.756 ;
  LAYER M2 ;
        RECT 18.48 19.724 21.36 19.756 ;
  LAYER M1 ;
        RECT 18.464 19.704 18.496 19.776 ;
  LAYER M2 ;
        RECT 18.444 19.724 18.516 19.756 ;
  LAYER M1 ;
        RECT 24.224 19.704 24.256 19.776 ;
  LAYER M2 ;
        RECT 24.204 19.724 24.276 19.756 ;
  LAYER M2 ;
        RECT 21.36 19.724 24.24 19.756 ;
  LAYER M1 ;
        RECT 21.344 19.704 21.376 19.776 ;
  LAYER M2 ;
        RECT 21.324 19.724 21.396 19.756 ;
  LAYER M1 ;
        RECT 27.104 19.704 27.136 19.776 ;
  LAYER M2 ;
        RECT 27.084 19.724 27.156 19.756 ;
  LAYER M2 ;
        RECT 24.24 19.724 27.12 19.756 ;
  LAYER M1 ;
        RECT 24.224 19.704 24.256 19.776 ;
  LAYER M2 ;
        RECT 24.204 19.724 24.276 19.756 ;
  LAYER M1 ;
        RECT 27.104 34.404 27.136 34.476 ;
  LAYER M2 ;
        RECT 27.084 34.424 27.156 34.456 ;
  LAYER M2 ;
        RECT 27.12 34.424 30 34.456 ;
  LAYER M1 ;
        RECT 29.984 34.404 30.016 34.476 ;
  LAYER M2 ;
        RECT 29.964 34.424 30.036 34.456 ;
  LAYER M1 ;
        RECT 24.224 34.404 24.256 34.476 ;
  LAYER M2 ;
        RECT 24.204 34.424 24.276 34.456 ;
  LAYER M2 ;
        RECT 24.24 34.424 27.12 34.456 ;
  LAYER M1 ;
        RECT 27.104 34.404 27.136 34.476 ;
  LAYER M2 ;
        RECT 27.084 34.424 27.156 34.456 ;
  LAYER M1 ;
        RECT 16.064 34.404 16.096 36.912 ;
  LAYER M1 ;
        RECT 16.128 34.404 16.16 36.912 ;
  LAYER M1 ;
        RECT 16.192 34.404 16.224 36.912 ;
  LAYER M1 ;
        RECT 16.256 34.404 16.288 36.912 ;
  LAYER M1 ;
        RECT 16.32 34.404 16.352 36.912 ;
  LAYER M1 ;
        RECT 16.384 34.404 16.416 36.912 ;
  LAYER M1 ;
        RECT 16.448 34.404 16.48 36.912 ;
  LAYER M1 ;
        RECT 16.512 34.404 16.544 36.912 ;
  LAYER M1 ;
        RECT 16.576 34.404 16.608 36.912 ;
  LAYER M1 ;
        RECT 16.64 34.404 16.672 36.912 ;
  LAYER M1 ;
        RECT 16.704 34.404 16.736 36.912 ;
  LAYER M1 ;
        RECT 16.768 34.404 16.8 36.912 ;
  LAYER M1 ;
        RECT 16.832 34.404 16.864 36.912 ;
  LAYER M1 ;
        RECT 16.896 34.404 16.928 36.912 ;
  LAYER M1 ;
        RECT 16.96 34.404 16.992 36.912 ;
  LAYER M1 ;
        RECT 17.024 34.404 17.056 36.912 ;
  LAYER M1 ;
        RECT 17.088 34.404 17.12 36.912 ;
  LAYER M1 ;
        RECT 17.152 34.404 17.184 36.912 ;
  LAYER M1 ;
        RECT 17.216 34.404 17.248 36.912 ;
  LAYER M1 ;
        RECT 17.28 34.404 17.312 36.912 ;
  LAYER M1 ;
        RECT 17.344 34.404 17.376 36.912 ;
  LAYER M1 ;
        RECT 17.408 34.404 17.44 36.912 ;
  LAYER M1 ;
        RECT 17.472 34.404 17.504 36.912 ;
  LAYER M1 ;
        RECT 17.536 34.404 17.568 36.912 ;
  LAYER M1 ;
        RECT 17.6 34.404 17.632 36.912 ;
  LAYER M1 ;
        RECT 17.664 34.404 17.696 36.912 ;
  LAYER M1 ;
        RECT 17.728 34.404 17.76 36.912 ;
  LAYER M1 ;
        RECT 17.792 34.404 17.824 36.912 ;
  LAYER M1 ;
        RECT 17.856 34.404 17.888 36.912 ;
  LAYER M1 ;
        RECT 17.92 34.404 17.952 36.912 ;
  LAYER M1 ;
        RECT 17.984 34.404 18.016 36.912 ;
  LAYER M1 ;
        RECT 18.048 34.404 18.08 36.912 ;
  LAYER M1 ;
        RECT 18.112 34.404 18.144 36.912 ;
  LAYER M1 ;
        RECT 18.176 34.404 18.208 36.912 ;
  LAYER M1 ;
        RECT 18.24 34.404 18.272 36.912 ;
  LAYER M1 ;
        RECT 18.304 34.404 18.336 36.912 ;
  LAYER M1 ;
        RECT 18.368 34.404 18.4 36.912 ;
  LAYER M2 ;
        RECT 16.044 36.796 18.516 36.828 ;
  LAYER M2 ;
        RECT 16.044 36.732 18.516 36.764 ;
  LAYER M2 ;
        RECT 16.044 36.668 18.516 36.7 ;
  LAYER M2 ;
        RECT 16.044 36.604 18.516 36.636 ;
  LAYER M2 ;
        RECT 16.044 36.54 18.516 36.572 ;
  LAYER M2 ;
        RECT 16.044 36.476 18.516 36.508 ;
  LAYER M2 ;
        RECT 16.044 36.412 18.516 36.444 ;
  LAYER M2 ;
        RECT 16.044 36.348 18.516 36.38 ;
  LAYER M2 ;
        RECT 16.044 36.284 18.516 36.316 ;
  LAYER M2 ;
        RECT 16.044 36.22 18.516 36.252 ;
  LAYER M2 ;
        RECT 16.044 36.156 18.516 36.188 ;
  LAYER M2 ;
        RECT 16.044 36.092 18.516 36.124 ;
  LAYER M2 ;
        RECT 16.044 36.028 18.516 36.06 ;
  LAYER M2 ;
        RECT 16.044 35.964 18.516 35.996 ;
  LAYER M2 ;
        RECT 16.044 35.9 18.516 35.932 ;
  LAYER M2 ;
        RECT 16.044 35.836 18.516 35.868 ;
  LAYER M2 ;
        RECT 16.044 35.772 18.516 35.804 ;
  LAYER M2 ;
        RECT 16.044 35.708 18.516 35.74 ;
  LAYER M2 ;
        RECT 16.044 35.644 18.516 35.676 ;
  LAYER M2 ;
        RECT 16.044 35.58 18.516 35.612 ;
  LAYER M2 ;
        RECT 16.044 35.516 18.516 35.548 ;
  LAYER M2 ;
        RECT 16.044 35.452 18.516 35.484 ;
  LAYER M2 ;
        RECT 16.044 35.388 18.516 35.42 ;
  LAYER M2 ;
        RECT 16.044 35.324 18.516 35.356 ;
  LAYER M2 ;
        RECT 16.044 35.26 18.516 35.292 ;
  LAYER M2 ;
        RECT 16.044 35.196 18.516 35.228 ;
  LAYER M2 ;
        RECT 16.044 35.132 18.516 35.164 ;
  LAYER M2 ;
        RECT 16.044 35.068 18.516 35.1 ;
  LAYER M2 ;
        RECT 16.044 35.004 18.516 35.036 ;
  LAYER M2 ;
        RECT 16.044 34.94 18.516 34.972 ;
  LAYER M2 ;
        RECT 16.044 34.876 18.516 34.908 ;
  LAYER M2 ;
        RECT 16.044 34.812 18.516 34.844 ;
  LAYER M2 ;
        RECT 16.044 34.748 18.516 34.78 ;
  LAYER M2 ;
        RECT 16.044 34.684 18.516 34.716 ;
  LAYER M2 ;
        RECT 16.044 34.62 18.516 34.652 ;
  LAYER M2 ;
        RECT 16.044 34.556 18.516 34.588 ;
  LAYER M3 ;
        RECT 16.064 34.404 16.096 36.912 ;
  LAYER M3 ;
        RECT 16.128 34.404 16.16 36.912 ;
  LAYER M3 ;
        RECT 16.192 34.404 16.224 36.912 ;
  LAYER M3 ;
        RECT 16.256 34.404 16.288 36.912 ;
  LAYER M3 ;
        RECT 16.32 34.404 16.352 36.912 ;
  LAYER M3 ;
        RECT 16.384 34.404 16.416 36.912 ;
  LAYER M3 ;
        RECT 16.448 34.404 16.48 36.912 ;
  LAYER M3 ;
        RECT 16.512 34.404 16.544 36.912 ;
  LAYER M3 ;
        RECT 16.576 34.404 16.608 36.912 ;
  LAYER M3 ;
        RECT 16.64 34.404 16.672 36.912 ;
  LAYER M3 ;
        RECT 16.704 34.404 16.736 36.912 ;
  LAYER M3 ;
        RECT 16.768 34.404 16.8 36.912 ;
  LAYER M3 ;
        RECT 16.832 34.404 16.864 36.912 ;
  LAYER M3 ;
        RECT 16.896 34.404 16.928 36.912 ;
  LAYER M3 ;
        RECT 16.96 34.404 16.992 36.912 ;
  LAYER M3 ;
        RECT 17.024 34.404 17.056 36.912 ;
  LAYER M3 ;
        RECT 17.088 34.404 17.12 36.912 ;
  LAYER M3 ;
        RECT 17.152 34.404 17.184 36.912 ;
  LAYER M3 ;
        RECT 17.216 34.404 17.248 36.912 ;
  LAYER M3 ;
        RECT 17.28 34.404 17.312 36.912 ;
  LAYER M3 ;
        RECT 17.344 34.404 17.376 36.912 ;
  LAYER M3 ;
        RECT 17.408 34.404 17.44 36.912 ;
  LAYER M3 ;
        RECT 17.472 34.404 17.504 36.912 ;
  LAYER M3 ;
        RECT 17.536 34.404 17.568 36.912 ;
  LAYER M3 ;
        RECT 17.6 34.404 17.632 36.912 ;
  LAYER M3 ;
        RECT 17.664 34.404 17.696 36.912 ;
  LAYER M3 ;
        RECT 17.728 34.404 17.76 36.912 ;
  LAYER M3 ;
        RECT 17.792 34.404 17.824 36.912 ;
  LAYER M3 ;
        RECT 17.856 34.404 17.888 36.912 ;
  LAYER M3 ;
        RECT 17.92 34.404 17.952 36.912 ;
  LAYER M3 ;
        RECT 17.984 34.404 18.016 36.912 ;
  LAYER M3 ;
        RECT 18.048 34.404 18.08 36.912 ;
  LAYER M3 ;
        RECT 18.112 34.404 18.144 36.912 ;
  LAYER M3 ;
        RECT 18.176 34.404 18.208 36.912 ;
  LAYER M3 ;
        RECT 18.24 34.404 18.272 36.912 ;
  LAYER M3 ;
        RECT 18.304 34.404 18.336 36.912 ;
  LAYER M3 ;
        RECT 18.368 34.404 18.4 36.912 ;
  LAYER M3 ;
        RECT 18.464 34.404 18.496 36.912 ;
  LAYER M1 ;
        RECT 16.079 34.44 16.081 36.876 ;
  LAYER M1 ;
        RECT 16.159 34.44 16.161 36.876 ;
  LAYER M1 ;
        RECT 16.239 34.44 16.241 36.876 ;
  LAYER M1 ;
        RECT 16.319 34.44 16.321 36.876 ;
  LAYER M1 ;
        RECT 16.399 34.44 16.401 36.876 ;
  LAYER M1 ;
        RECT 16.479 34.44 16.481 36.876 ;
  LAYER M1 ;
        RECT 16.559 34.44 16.561 36.876 ;
  LAYER M1 ;
        RECT 16.639 34.44 16.641 36.876 ;
  LAYER M1 ;
        RECT 16.719 34.44 16.721 36.876 ;
  LAYER M1 ;
        RECT 16.799 34.44 16.801 36.876 ;
  LAYER M1 ;
        RECT 16.879 34.44 16.881 36.876 ;
  LAYER M1 ;
        RECT 16.959 34.44 16.961 36.876 ;
  LAYER M1 ;
        RECT 17.039 34.44 17.041 36.876 ;
  LAYER M1 ;
        RECT 17.119 34.44 17.121 36.876 ;
  LAYER M1 ;
        RECT 17.199 34.44 17.201 36.876 ;
  LAYER M1 ;
        RECT 17.279 34.44 17.281 36.876 ;
  LAYER M1 ;
        RECT 17.359 34.44 17.361 36.876 ;
  LAYER M1 ;
        RECT 17.439 34.44 17.441 36.876 ;
  LAYER M1 ;
        RECT 17.519 34.44 17.521 36.876 ;
  LAYER M1 ;
        RECT 17.599 34.44 17.601 36.876 ;
  LAYER M1 ;
        RECT 17.679 34.44 17.681 36.876 ;
  LAYER M1 ;
        RECT 17.759 34.44 17.761 36.876 ;
  LAYER M1 ;
        RECT 17.839 34.44 17.841 36.876 ;
  LAYER M1 ;
        RECT 17.919 34.44 17.921 36.876 ;
  LAYER M1 ;
        RECT 17.999 34.44 18.001 36.876 ;
  LAYER M1 ;
        RECT 18.079 34.44 18.081 36.876 ;
  LAYER M1 ;
        RECT 18.159 34.44 18.161 36.876 ;
  LAYER M1 ;
        RECT 18.239 34.44 18.241 36.876 ;
  LAYER M1 ;
        RECT 18.319 34.44 18.321 36.876 ;
  LAYER M1 ;
        RECT 18.399 34.44 18.401 36.876 ;
  LAYER M2 ;
        RECT 16.08 36.875 18.48 36.877 ;
  LAYER M2 ;
        RECT 16.08 36.791 18.48 36.793 ;
  LAYER M2 ;
        RECT 16.08 36.707 18.48 36.709 ;
  LAYER M2 ;
        RECT 16.08 36.623 18.48 36.625 ;
  LAYER M2 ;
        RECT 16.08 36.539 18.48 36.541 ;
  LAYER M2 ;
        RECT 16.08 36.455 18.48 36.457 ;
  LAYER M2 ;
        RECT 16.08 36.371 18.48 36.373 ;
  LAYER M2 ;
        RECT 16.08 36.287 18.48 36.289 ;
  LAYER M2 ;
        RECT 16.08 36.203 18.48 36.205 ;
  LAYER M2 ;
        RECT 16.08 36.119 18.48 36.121 ;
  LAYER M2 ;
        RECT 16.08 36.035 18.48 36.037 ;
  LAYER M2 ;
        RECT 16.08 35.951 18.48 35.953 ;
  LAYER M2 ;
        RECT 16.08 35.8675 18.48 35.8695 ;
  LAYER M2 ;
        RECT 16.08 35.783 18.48 35.785 ;
  LAYER M2 ;
        RECT 16.08 35.699 18.48 35.701 ;
  LAYER M2 ;
        RECT 16.08 35.615 18.48 35.617 ;
  LAYER M2 ;
        RECT 16.08 35.531 18.48 35.533 ;
  LAYER M2 ;
        RECT 16.08 35.447 18.48 35.449 ;
  LAYER M2 ;
        RECT 16.08 35.363 18.48 35.365 ;
  LAYER M2 ;
        RECT 16.08 35.279 18.48 35.281 ;
  LAYER M2 ;
        RECT 16.08 35.195 18.48 35.197 ;
  LAYER M2 ;
        RECT 16.08 35.111 18.48 35.113 ;
  LAYER M2 ;
        RECT 16.08 35.027 18.48 35.029 ;
  LAYER M2 ;
        RECT 16.08 34.943 18.48 34.945 ;
  LAYER M2 ;
        RECT 16.08 34.859 18.48 34.861 ;
  LAYER M2 ;
        RECT 16.08 34.775 18.48 34.777 ;
  LAYER M2 ;
        RECT 16.08 34.691 18.48 34.693 ;
  LAYER M2 ;
        RECT 16.08 34.607 18.48 34.609 ;
  LAYER M2 ;
        RECT 16.08 34.523 18.48 34.525 ;
  LAYER M1 ;
        RECT 16.064 31.464 16.096 33.972 ;
  LAYER M1 ;
        RECT 16.128 31.464 16.16 33.972 ;
  LAYER M1 ;
        RECT 16.192 31.464 16.224 33.972 ;
  LAYER M1 ;
        RECT 16.256 31.464 16.288 33.972 ;
  LAYER M1 ;
        RECT 16.32 31.464 16.352 33.972 ;
  LAYER M1 ;
        RECT 16.384 31.464 16.416 33.972 ;
  LAYER M1 ;
        RECT 16.448 31.464 16.48 33.972 ;
  LAYER M1 ;
        RECT 16.512 31.464 16.544 33.972 ;
  LAYER M1 ;
        RECT 16.576 31.464 16.608 33.972 ;
  LAYER M1 ;
        RECT 16.64 31.464 16.672 33.972 ;
  LAYER M1 ;
        RECT 16.704 31.464 16.736 33.972 ;
  LAYER M1 ;
        RECT 16.768 31.464 16.8 33.972 ;
  LAYER M1 ;
        RECT 16.832 31.464 16.864 33.972 ;
  LAYER M1 ;
        RECT 16.896 31.464 16.928 33.972 ;
  LAYER M1 ;
        RECT 16.96 31.464 16.992 33.972 ;
  LAYER M1 ;
        RECT 17.024 31.464 17.056 33.972 ;
  LAYER M1 ;
        RECT 17.088 31.464 17.12 33.972 ;
  LAYER M1 ;
        RECT 17.152 31.464 17.184 33.972 ;
  LAYER M1 ;
        RECT 17.216 31.464 17.248 33.972 ;
  LAYER M1 ;
        RECT 17.28 31.464 17.312 33.972 ;
  LAYER M1 ;
        RECT 17.344 31.464 17.376 33.972 ;
  LAYER M1 ;
        RECT 17.408 31.464 17.44 33.972 ;
  LAYER M1 ;
        RECT 17.472 31.464 17.504 33.972 ;
  LAYER M1 ;
        RECT 17.536 31.464 17.568 33.972 ;
  LAYER M1 ;
        RECT 17.6 31.464 17.632 33.972 ;
  LAYER M1 ;
        RECT 17.664 31.464 17.696 33.972 ;
  LAYER M1 ;
        RECT 17.728 31.464 17.76 33.972 ;
  LAYER M1 ;
        RECT 17.792 31.464 17.824 33.972 ;
  LAYER M1 ;
        RECT 17.856 31.464 17.888 33.972 ;
  LAYER M1 ;
        RECT 17.92 31.464 17.952 33.972 ;
  LAYER M1 ;
        RECT 17.984 31.464 18.016 33.972 ;
  LAYER M1 ;
        RECT 18.048 31.464 18.08 33.972 ;
  LAYER M1 ;
        RECT 18.112 31.464 18.144 33.972 ;
  LAYER M1 ;
        RECT 18.176 31.464 18.208 33.972 ;
  LAYER M1 ;
        RECT 18.24 31.464 18.272 33.972 ;
  LAYER M1 ;
        RECT 18.304 31.464 18.336 33.972 ;
  LAYER M1 ;
        RECT 18.368 31.464 18.4 33.972 ;
  LAYER M2 ;
        RECT 16.044 33.856 18.516 33.888 ;
  LAYER M2 ;
        RECT 16.044 33.792 18.516 33.824 ;
  LAYER M2 ;
        RECT 16.044 33.728 18.516 33.76 ;
  LAYER M2 ;
        RECT 16.044 33.664 18.516 33.696 ;
  LAYER M2 ;
        RECT 16.044 33.6 18.516 33.632 ;
  LAYER M2 ;
        RECT 16.044 33.536 18.516 33.568 ;
  LAYER M2 ;
        RECT 16.044 33.472 18.516 33.504 ;
  LAYER M2 ;
        RECT 16.044 33.408 18.516 33.44 ;
  LAYER M2 ;
        RECT 16.044 33.344 18.516 33.376 ;
  LAYER M2 ;
        RECT 16.044 33.28 18.516 33.312 ;
  LAYER M2 ;
        RECT 16.044 33.216 18.516 33.248 ;
  LAYER M2 ;
        RECT 16.044 33.152 18.516 33.184 ;
  LAYER M2 ;
        RECT 16.044 33.088 18.516 33.12 ;
  LAYER M2 ;
        RECT 16.044 33.024 18.516 33.056 ;
  LAYER M2 ;
        RECT 16.044 32.96 18.516 32.992 ;
  LAYER M2 ;
        RECT 16.044 32.896 18.516 32.928 ;
  LAYER M2 ;
        RECT 16.044 32.832 18.516 32.864 ;
  LAYER M2 ;
        RECT 16.044 32.768 18.516 32.8 ;
  LAYER M2 ;
        RECT 16.044 32.704 18.516 32.736 ;
  LAYER M2 ;
        RECT 16.044 32.64 18.516 32.672 ;
  LAYER M2 ;
        RECT 16.044 32.576 18.516 32.608 ;
  LAYER M2 ;
        RECT 16.044 32.512 18.516 32.544 ;
  LAYER M2 ;
        RECT 16.044 32.448 18.516 32.48 ;
  LAYER M2 ;
        RECT 16.044 32.384 18.516 32.416 ;
  LAYER M2 ;
        RECT 16.044 32.32 18.516 32.352 ;
  LAYER M2 ;
        RECT 16.044 32.256 18.516 32.288 ;
  LAYER M2 ;
        RECT 16.044 32.192 18.516 32.224 ;
  LAYER M2 ;
        RECT 16.044 32.128 18.516 32.16 ;
  LAYER M2 ;
        RECT 16.044 32.064 18.516 32.096 ;
  LAYER M2 ;
        RECT 16.044 32 18.516 32.032 ;
  LAYER M2 ;
        RECT 16.044 31.936 18.516 31.968 ;
  LAYER M2 ;
        RECT 16.044 31.872 18.516 31.904 ;
  LAYER M2 ;
        RECT 16.044 31.808 18.516 31.84 ;
  LAYER M2 ;
        RECT 16.044 31.744 18.516 31.776 ;
  LAYER M2 ;
        RECT 16.044 31.68 18.516 31.712 ;
  LAYER M2 ;
        RECT 16.044 31.616 18.516 31.648 ;
  LAYER M3 ;
        RECT 16.064 31.464 16.096 33.972 ;
  LAYER M3 ;
        RECT 16.128 31.464 16.16 33.972 ;
  LAYER M3 ;
        RECT 16.192 31.464 16.224 33.972 ;
  LAYER M3 ;
        RECT 16.256 31.464 16.288 33.972 ;
  LAYER M3 ;
        RECT 16.32 31.464 16.352 33.972 ;
  LAYER M3 ;
        RECT 16.384 31.464 16.416 33.972 ;
  LAYER M3 ;
        RECT 16.448 31.464 16.48 33.972 ;
  LAYER M3 ;
        RECT 16.512 31.464 16.544 33.972 ;
  LAYER M3 ;
        RECT 16.576 31.464 16.608 33.972 ;
  LAYER M3 ;
        RECT 16.64 31.464 16.672 33.972 ;
  LAYER M3 ;
        RECT 16.704 31.464 16.736 33.972 ;
  LAYER M3 ;
        RECT 16.768 31.464 16.8 33.972 ;
  LAYER M3 ;
        RECT 16.832 31.464 16.864 33.972 ;
  LAYER M3 ;
        RECT 16.896 31.464 16.928 33.972 ;
  LAYER M3 ;
        RECT 16.96 31.464 16.992 33.972 ;
  LAYER M3 ;
        RECT 17.024 31.464 17.056 33.972 ;
  LAYER M3 ;
        RECT 17.088 31.464 17.12 33.972 ;
  LAYER M3 ;
        RECT 17.152 31.464 17.184 33.972 ;
  LAYER M3 ;
        RECT 17.216 31.464 17.248 33.972 ;
  LAYER M3 ;
        RECT 17.28 31.464 17.312 33.972 ;
  LAYER M3 ;
        RECT 17.344 31.464 17.376 33.972 ;
  LAYER M3 ;
        RECT 17.408 31.464 17.44 33.972 ;
  LAYER M3 ;
        RECT 17.472 31.464 17.504 33.972 ;
  LAYER M3 ;
        RECT 17.536 31.464 17.568 33.972 ;
  LAYER M3 ;
        RECT 17.6 31.464 17.632 33.972 ;
  LAYER M3 ;
        RECT 17.664 31.464 17.696 33.972 ;
  LAYER M3 ;
        RECT 17.728 31.464 17.76 33.972 ;
  LAYER M3 ;
        RECT 17.792 31.464 17.824 33.972 ;
  LAYER M3 ;
        RECT 17.856 31.464 17.888 33.972 ;
  LAYER M3 ;
        RECT 17.92 31.464 17.952 33.972 ;
  LAYER M3 ;
        RECT 17.984 31.464 18.016 33.972 ;
  LAYER M3 ;
        RECT 18.048 31.464 18.08 33.972 ;
  LAYER M3 ;
        RECT 18.112 31.464 18.144 33.972 ;
  LAYER M3 ;
        RECT 18.176 31.464 18.208 33.972 ;
  LAYER M3 ;
        RECT 18.24 31.464 18.272 33.972 ;
  LAYER M3 ;
        RECT 18.304 31.464 18.336 33.972 ;
  LAYER M3 ;
        RECT 18.368 31.464 18.4 33.972 ;
  LAYER M3 ;
        RECT 18.464 31.464 18.496 33.972 ;
  LAYER M1 ;
        RECT 16.079 31.5 16.081 33.936 ;
  LAYER M1 ;
        RECT 16.159 31.5 16.161 33.936 ;
  LAYER M1 ;
        RECT 16.239 31.5 16.241 33.936 ;
  LAYER M1 ;
        RECT 16.319 31.5 16.321 33.936 ;
  LAYER M1 ;
        RECT 16.399 31.5 16.401 33.936 ;
  LAYER M1 ;
        RECT 16.479 31.5 16.481 33.936 ;
  LAYER M1 ;
        RECT 16.559 31.5 16.561 33.936 ;
  LAYER M1 ;
        RECT 16.639 31.5 16.641 33.936 ;
  LAYER M1 ;
        RECT 16.719 31.5 16.721 33.936 ;
  LAYER M1 ;
        RECT 16.799 31.5 16.801 33.936 ;
  LAYER M1 ;
        RECT 16.879 31.5 16.881 33.936 ;
  LAYER M1 ;
        RECT 16.959 31.5 16.961 33.936 ;
  LAYER M1 ;
        RECT 17.039 31.5 17.041 33.936 ;
  LAYER M1 ;
        RECT 17.119 31.5 17.121 33.936 ;
  LAYER M1 ;
        RECT 17.199 31.5 17.201 33.936 ;
  LAYER M1 ;
        RECT 17.279 31.5 17.281 33.936 ;
  LAYER M1 ;
        RECT 17.359 31.5 17.361 33.936 ;
  LAYER M1 ;
        RECT 17.439 31.5 17.441 33.936 ;
  LAYER M1 ;
        RECT 17.519 31.5 17.521 33.936 ;
  LAYER M1 ;
        RECT 17.599 31.5 17.601 33.936 ;
  LAYER M1 ;
        RECT 17.679 31.5 17.681 33.936 ;
  LAYER M1 ;
        RECT 17.759 31.5 17.761 33.936 ;
  LAYER M1 ;
        RECT 17.839 31.5 17.841 33.936 ;
  LAYER M1 ;
        RECT 17.919 31.5 17.921 33.936 ;
  LAYER M1 ;
        RECT 17.999 31.5 18.001 33.936 ;
  LAYER M1 ;
        RECT 18.079 31.5 18.081 33.936 ;
  LAYER M1 ;
        RECT 18.159 31.5 18.161 33.936 ;
  LAYER M1 ;
        RECT 18.239 31.5 18.241 33.936 ;
  LAYER M1 ;
        RECT 18.319 31.5 18.321 33.936 ;
  LAYER M1 ;
        RECT 18.399 31.5 18.401 33.936 ;
  LAYER M2 ;
        RECT 16.08 33.935 18.48 33.937 ;
  LAYER M2 ;
        RECT 16.08 33.851 18.48 33.853 ;
  LAYER M2 ;
        RECT 16.08 33.767 18.48 33.769 ;
  LAYER M2 ;
        RECT 16.08 33.683 18.48 33.685 ;
  LAYER M2 ;
        RECT 16.08 33.599 18.48 33.601 ;
  LAYER M2 ;
        RECT 16.08 33.515 18.48 33.517 ;
  LAYER M2 ;
        RECT 16.08 33.431 18.48 33.433 ;
  LAYER M2 ;
        RECT 16.08 33.347 18.48 33.349 ;
  LAYER M2 ;
        RECT 16.08 33.263 18.48 33.265 ;
  LAYER M2 ;
        RECT 16.08 33.179 18.48 33.181 ;
  LAYER M2 ;
        RECT 16.08 33.095 18.48 33.097 ;
  LAYER M2 ;
        RECT 16.08 33.011 18.48 33.013 ;
  LAYER M2 ;
        RECT 16.08 32.9275 18.48 32.9295 ;
  LAYER M2 ;
        RECT 16.08 32.843 18.48 32.845 ;
  LAYER M2 ;
        RECT 16.08 32.759 18.48 32.761 ;
  LAYER M2 ;
        RECT 16.08 32.675 18.48 32.677 ;
  LAYER M2 ;
        RECT 16.08 32.591 18.48 32.593 ;
  LAYER M2 ;
        RECT 16.08 32.507 18.48 32.509 ;
  LAYER M2 ;
        RECT 16.08 32.423 18.48 32.425 ;
  LAYER M2 ;
        RECT 16.08 32.339 18.48 32.341 ;
  LAYER M2 ;
        RECT 16.08 32.255 18.48 32.257 ;
  LAYER M2 ;
        RECT 16.08 32.171 18.48 32.173 ;
  LAYER M2 ;
        RECT 16.08 32.087 18.48 32.089 ;
  LAYER M2 ;
        RECT 16.08 32.003 18.48 32.005 ;
  LAYER M2 ;
        RECT 16.08 31.919 18.48 31.921 ;
  LAYER M2 ;
        RECT 16.08 31.835 18.48 31.837 ;
  LAYER M2 ;
        RECT 16.08 31.751 18.48 31.753 ;
  LAYER M2 ;
        RECT 16.08 31.667 18.48 31.669 ;
  LAYER M2 ;
        RECT 16.08 31.583 18.48 31.585 ;
  LAYER M1 ;
        RECT 16.064 28.524 16.096 31.032 ;
  LAYER M1 ;
        RECT 16.128 28.524 16.16 31.032 ;
  LAYER M1 ;
        RECT 16.192 28.524 16.224 31.032 ;
  LAYER M1 ;
        RECT 16.256 28.524 16.288 31.032 ;
  LAYER M1 ;
        RECT 16.32 28.524 16.352 31.032 ;
  LAYER M1 ;
        RECT 16.384 28.524 16.416 31.032 ;
  LAYER M1 ;
        RECT 16.448 28.524 16.48 31.032 ;
  LAYER M1 ;
        RECT 16.512 28.524 16.544 31.032 ;
  LAYER M1 ;
        RECT 16.576 28.524 16.608 31.032 ;
  LAYER M1 ;
        RECT 16.64 28.524 16.672 31.032 ;
  LAYER M1 ;
        RECT 16.704 28.524 16.736 31.032 ;
  LAYER M1 ;
        RECT 16.768 28.524 16.8 31.032 ;
  LAYER M1 ;
        RECT 16.832 28.524 16.864 31.032 ;
  LAYER M1 ;
        RECT 16.896 28.524 16.928 31.032 ;
  LAYER M1 ;
        RECT 16.96 28.524 16.992 31.032 ;
  LAYER M1 ;
        RECT 17.024 28.524 17.056 31.032 ;
  LAYER M1 ;
        RECT 17.088 28.524 17.12 31.032 ;
  LAYER M1 ;
        RECT 17.152 28.524 17.184 31.032 ;
  LAYER M1 ;
        RECT 17.216 28.524 17.248 31.032 ;
  LAYER M1 ;
        RECT 17.28 28.524 17.312 31.032 ;
  LAYER M1 ;
        RECT 17.344 28.524 17.376 31.032 ;
  LAYER M1 ;
        RECT 17.408 28.524 17.44 31.032 ;
  LAYER M1 ;
        RECT 17.472 28.524 17.504 31.032 ;
  LAYER M1 ;
        RECT 17.536 28.524 17.568 31.032 ;
  LAYER M1 ;
        RECT 17.6 28.524 17.632 31.032 ;
  LAYER M1 ;
        RECT 17.664 28.524 17.696 31.032 ;
  LAYER M1 ;
        RECT 17.728 28.524 17.76 31.032 ;
  LAYER M1 ;
        RECT 17.792 28.524 17.824 31.032 ;
  LAYER M1 ;
        RECT 17.856 28.524 17.888 31.032 ;
  LAYER M1 ;
        RECT 17.92 28.524 17.952 31.032 ;
  LAYER M1 ;
        RECT 17.984 28.524 18.016 31.032 ;
  LAYER M1 ;
        RECT 18.048 28.524 18.08 31.032 ;
  LAYER M1 ;
        RECT 18.112 28.524 18.144 31.032 ;
  LAYER M1 ;
        RECT 18.176 28.524 18.208 31.032 ;
  LAYER M1 ;
        RECT 18.24 28.524 18.272 31.032 ;
  LAYER M1 ;
        RECT 18.304 28.524 18.336 31.032 ;
  LAYER M1 ;
        RECT 18.368 28.524 18.4 31.032 ;
  LAYER M2 ;
        RECT 16.044 30.916 18.516 30.948 ;
  LAYER M2 ;
        RECT 16.044 30.852 18.516 30.884 ;
  LAYER M2 ;
        RECT 16.044 30.788 18.516 30.82 ;
  LAYER M2 ;
        RECT 16.044 30.724 18.516 30.756 ;
  LAYER M2 ;
        RECT 16.044 30.66 18.516 30.692 ;
  LAYER M2 ;
        RECT 16.044 30.596 18.516 30.628 ;
  LAYER M2 ;
        RECT 16.044 30.532 18.516 30.564 ;
  LAYER M2 ;
        RECT 16.044 30.468 18.516 30.5 ;
  LAYER M2 ;
        RECT 16.044 30.404 18.516 30.436 ;
  LAYER M2 ;
        RECT 16.044 30.34 18.516 30.372 ;
  LAYER M2 ;
        RECT 16.044 30.276 18.516 30.308 ;
  LAYER M2 ;
        RECT 16.044 30.212 18.516 30.244 ;
  LAYER M2 ;
        RECT 16.044 30.148 18.516 30.18 ;
  LAYER M2 ;
        RECT 16.044 30.084 18.516 30.116 ;
  LAYER M2 ;
        RECT 16.044 30.02 18.516 30.052 ;
  LAYER M2 ;
        RECT 16.044 29.956 18.516 29.988 ;
  LAYER M2 ;
        RECT 16.044 29.892 18.516 29.924 ;
  LAYER M2 ;
        RECT 16.044 29.828 18.516 29.86 ;
  LAYER M2 ;
        RECT 16.044 29.764 18.516 29.796 ;
  LAYER M2 ;
        RECT 16.044 29.7 18.516 29.732 ;
  LAYER M2 ;
        RECT 16.044 29.636 18.516 29.668 ;
  LAYER M2 ;
        RECT 16.044 29.572 18.516 29.604 ;
  LAYER M2 ;
        RECT 16.044 29.508 18.516 29.54 ;
  LAYER M2 ;
        RECT 16.044 29.444 18.516 29.476 ;
  LAYER M2 ;
        RECT 16.044 29.38 18.516 29.412 ;
  LAYER M2 ;
        RECT 16.044 29.316 18.516 29.348 ;
  LAYER M2 ;
        RECT 16.044 29.252 18.516 29.284 ;
  LAYER M2 ;
        RECT 16.044 29.188 18.516 29.22 ;
  LAYER M2 ;
        RECT 16.044 29.124 18.516 29.156 ;
  LAYER M2 ;
        RECT 16.044 29.06 18.516 29.092 ;
  LAYER M2 ;
        RECT 16.044 28.996 18.516 29.028 ;
  LAYER M2 ;
        RECT 16.044 28.932 18.516 28.964 ;
  LAYER M2 ;
        RECT 16.044 28.868 18.516 28.9 ;
  LAYER M2 ;
        RECT 16.044 28.804 18.516 28.836 ;
  LAYER M2 ;
        RECT 16.044 28.74 18.516 28.772 ;
  LAYER M2 ;
        RECT 16.044 28.676 18.516 28.708 ;
  LAYER M3 ;
        RECT 16.064 28.524 16.096 31.032 ;
  LAYER M3 ;
        RECT 16.128 28.524 16.16 31.032 ;
  LAYER M3 ;
        RECT 16.192 28.524 16.224 31.032 ;
  LAYER M3 ;
        RECT 16.256 28.524 16.288 31.032 ;
  LAYER M3 ;
        RECT 16.32 28.524 16.352 31.032 ;
  LAYER M3 ;
        RECT 16.384 28.524 16.416 31.032 ;
  LAYER M3 ;
        RECT 16.448 28.524 16.48 31.032 ;
  LAYER M3 ;
        RECT 16.512 28.524 16.544 31.032 ;
  LAYER M3 ;
        RECT 16.576 28.524 16.608 31.032 ;
  LAYER M3 ;
        RECT 16.64 28.524 16.672 31.032 ;
  LAYER M3 ;
        RECT 16.704 28.524 16.736 31.032 ;
  LAYER M3 ;
        RECT 16.768 28.524 16.8 31.032 ;
  LAYER M3 ;
        RECT 16.832 28.524 16.864 31.032 ;
  LAYER M3 ;
        RECT 16.896 28.524 16.928 31.032 ;
  LAYER M3 ;
        RECT 16.96 28.524 16.992 31.032 ;
  LAYER M3 ;
        RECT 17.024 28.524 17.056 31.032 ;
  LAYER M3 ;
        RECT 17.088 28.524 17.12 31.032 ;
  LAYER M3 ;
        RECT 17.152 28.524 17.184 31.032 ;
  LAYER M3 ;
        RECT 17.216 28.524 17.248 31.032 ;
  LAYER M3 ;
        RECT 17.28 28.524 17.312 31.032 ;
  LAYER M3 ;
        RECT 17.344 28.524 17.376 31.032 ;
  LAYER M3 ;
        RECT 17.408 28.524 17.44 31.032 ;
  LAYER M3 ;
        RECT 17.472 28.524 17.504 31.032 ;
  LAYER M3 ;
        RECT 17.536 28.524 17.568 31.032 ;
  LAYER M3 ;
        RECT 17.6 28.524 17.632 31.032 ;
  LAYER M3 ;
        RECT 17.664 28.524 17.696 31.032 ;
  LAYER M3 ;
        RECT 17.728 28.524 17.76 31.032 ;
  LAYER M3 ;
        RECT 17.792 28.524 17.824 31.032 ;
  LAYER M3 ;
        RECT 17.856 28.524 17.888 31.032 ;
  LAYER M3 ;
        RECT 17.92 28.524 17.952 31.032 ;
  LAYER M3 ;
        RECT 17.984 28.524 18.016 31.032 ;
  LAYER M3 ;
        RECT 18.048 28.524 18.08 31.032 ;
  LAYER M3 ;
        RECT 18.112 28.524 18.144 31.032 ;
  LAYER M3 ;
        RECT 18.176 28.524 18.208 31.032 ;
  LAYER M3 ;
        RECT 18.24 28.524 18.272 31.032 ;
  LAYER M3 ;
        RECT 18.304 28.524 18.336 31.032 ;
  LAYER M3 ;
        RECT 18.368 28.524 18.4 31.032 ;
  LAYER M3 ;
        RECT 18.464 28.524 18.496 31.032 ;
  LAYER M1 ;
        RECT 16.079 28.56 16.081 30.996 ;
  LAYER M1 ;
        RECT 16.159 28.56 16.161 30.996 ;
  LAYER M1 ;
        RECT 16.239 28.56 16.241 30.996 ;
  LAYER M1 ;
        RECT 16.319 28.56 16.321 30.996 ;
  LAYER M1 ;
        RECT 16.399 28.56 16.401 30.996 ;
  LAYER M1 ;
        RECT 16.479 28.56 16.481 30.996 ;
  LAYER M1 ;
        RECT 16.559 28.56 16.561 30.996 ;
  LAYER M1 ;
        RECT 16.639 28.56 16.641 30.996 ;
  LAYER M1 ;
        RECT 16.719 28.56 16.721 30.996 ;
  LAYER M1 ;
        RECT 16.799 28.56 16.801 30.996 ;
  LAYER M1 ;
        RECT 16.879 28.56 16.881 30.996 ;
  LAYER M1 ;
        RECT 16.959 28.56 16.961 30.996 ;
  LAYER M1 ;
        RECT 17.039 28.56 17.041 30.996 ;
  LAYER M1 ;
        RECT 17.119 28.56 17.121 30.996 ;
  LAYER M1 ;
        RECT 17.199 28.56 17.201 30.996 ;
  LAYER M1 ;
        RECT 17.279 28.56 17.281 30.996 ;
  LAYER M1 ;
        RECT 17.359 28.56 17.361 30.996 ;
  LAYER M1 ;
        RECT 17.439 28.56 17.441 30.996 ;
  LAYER M1 ;
        RECT 17.519 28.56 17.521 30.996 ;
  LAYER M1 ;
        RECT 17.599 28.56 17.601 30.996 ;
  LAYER M1 ;
        RECT 17.679 28.56 17.681 30.996 ;
  LAYER M1 ;
        RECT 17.759 28.56 17.761 30.996 ;
  LAYER M1 ;
        RECT 17.839 28.56 17.841 30.996 ;
  LAYER M1 ;
        RECT 17.919 28.56 17.921 30.996 ;
  LAYER M1 ;
        RECT 17.999 28.56 18.001 30.996 ;
  LAYER M1 ;
        RECT 18.079 28.56 18.081 30.996 ;
  LAYER M1 ;
        RECT 18.159 28.56 18.161 30.996 ;
  LAYER M1 ;
        RECT 18.239 28.56 18.241 30.996 ;
  LAYER M1 ;
        RECT 18.319 28.56 18.321 30.996 ;
  LAYER M1 ;
        RECT 18.399 28.56 18.401 30.996 ;
  LAYER M2 ;
        RECT 16.08 30.995 18.48 30.997 ;
  LAYER M2 ;
        RECT 16.08 30.911 18.48 30.913 ;
  LAYER M2 ;
        RECT 16.08 30.827 18.48 30.829 ;
  LAYER M2 ;
        RECT 16.08 30.743 18.48 30.745 ;
  LAYER M2 ;
        RECT 16.08 30.659 18.48 30.661 ;
  LAYER M2 ;
        RECT 16.08 30.575 18.48 30.577 ;
  LAYER M2 ;
        RECT 16.08 30.491 18.48 30.493 ;
  LAYER M2 ;
        RECT 16.08 30.407 18.48 30.409 ;
  LAYER M2 ;
        RECT 16.08 30.323 18.48 30.325 ;
  LAYER M2 ;
        RECT 16.08 30.239 18.48 30.241 ;
  LAYER M2 ;
        RECT 16.08 30.155 18.48 30.157 ;
  LAYER M2 ;
        RECT 16.08 30.071 18.48 30.073 ;
  LAYER M2 ;
        RECT 16.08 29.9875 18.48 29.9895 ;
  LAYER M2 ;
        RECT 16.08 29.903 18.48 29.905 ;
  LAYER M2 ;
        RECT 16.08 29.819 18.48 29.821 ;
  LAYER M2 ;
        RECT 16.08 29.735 18.48 29.737 ;
  LAYER M2 ;
        RECT 16.08 29.651 18.48 29.653 ;
  LAYER M2 ;
        RECT 16.08 29.567 18.48 29.569 ;
  LAYER M2 ;
        RECT 16.08 29.483 18.48 29.485 ;
  LAYER M2 ;
        RECT 16.08 29.399 18.48 29.401 ;
  LAYER M2 ;
        RECT 16.08 29.315 18.48 29.317 ;
  LAYER M2 ;
        RECT 16.08 29.231 18.48 29.233 ;
  LAYER M2 ;
        RECT 16.08 29.147 18.48 29.149 ;
  LAYER M2 ;
        RECT 16.08 29.063 18.48 29.065 ;
  LAYER M2 ;
        RECT 16.08 28.979 18.48 28.981 ;
  LAYER M2 ;
        RECT 16.08 28.895 18.48 28.897 ;
  LAYER M2 ;
        RECT 16.08 28.811 18.48 28.813 ;
  LAYER M2 ;
        RECT 16.08 28.727 18.48 28.729 ;
  LAYER M2 ;
        RECT 16.08 28.643 18.48 28.645 ;
  LAYER M1 ;
        RECT 16.064 25.584 16.096 28.092 ;
  LAYER M1 ;
        RECT 16.128 25.584 16.16 28.092 ;
  LAYER M1 ;
        RECT 16.192 25.584 16.224 28.092 ;
  LAYER M1 ;
        RECT 16.256 25.584 16.288 28.092 ;
  LAYER M1 ;
        RECT 16.32 25.584 16.352 28.092 ;
  LAYER M1 ;
        RECT 16.384 25.584 16.416 28.092 ;
  LAYER M1 ;
        RECT 16.448 25.584 16.48 28.092 ;
  LAYER M1 ;
        RECT 16.512 25.584 16.544 28.092 ;
  LAYER M1 ;
        RECT 16.576 25.584 16.608 28.092 ;
  LAYER M1 ;
        RECT 16.64 25.584 16.672 28.092 ;
  LAYER M1 ;
        RECT 16.704 25.584 16.736 28.092 ;
  LAYER M1 ;
        RECT 16.768 25.584 16.8 28.092 ;
  LAYER M1 ;
        RECT 16.832 25.584 16.864 28.092 ;
  LAYER M1 ;
        RECT 16.896 25.584 16.928 28.092 ;
  LAYER M1 ;
        RECT 16.96 25.584 16.992 28.092 ;
  LAYER M1 ;
        RECT 17.024 25.584 17.056 28.092 ;
  LAYER M1 ;
        RECT 17.088 25.584 17.12 28.092 ;
  LAYER M1 ;
        RECT 17.152 25.584 17.184 28.092 ;
  LAYER M1 ;
        RECT 17.216 25.584 17.248 28.092 ;
  LAYER M1 ;
        RECT 17.28 25.584 17.312 28.092 ;
  LAYER M1 ;
        RECT 17.344 25.584 17.376 28.092 ;
  LAYER M1 ;
        RECT 17.408 25.584 17.44 28.092 ;
  LAYER M1 ;
        RECT 17.472 25.584 17.504 28.092 ;
  LAYER M1 ;
        RECT 17.536 25.584 17.568 28.092 ;
  LAYER M1 ;
        RECT 17.6 25.584 17.632 28.092 ;
  LAYER M1 ;
        RECT 17.664 25.584 17.696 28.092 ;
  LAYER M1 ;
        RECT 17.728 25.584 17.76 28.092 ;
  LAYER M1 ;
        RECT 17.792 25.584 17.824 28.092 ;
  LAYER M1 ;
        RECT 17.856 25.584 17.888 28.092 ;
  LAYER M1 ;
        RECT 17.92 25.584 17.952 28.092 ;
  LAYER M1 ;
        RECT 17.984 25.584 18.016 28.092 ;
  LAYER M1 ;
        RECT 18.048 25.584 18.08 28.092 ;
  LAYER M1 ;
        RECT 18.112 25.584 18.144 28.092 ;
  LAYER M1 ;
        RECT 18.176 25.584 18.208 28.092 ;
  LAYER M1 ;
        RECT 18.24 25.584 18.272 28.092 ;
  LAYER M1 ;
        RECT 18.304 25.584 18.336 28.092 ;
  LAYER M1 ;
        RECT 18.368 25.584 18.4 28.092 ;
  LAYER M2 ;
        RECT 16.044 27.976 18.516 28.008 ;
  LAYER M2 ;
        RECT 16.044 27.912 18.516 27.944 ;
  LAYER M2 ;
        RECT 16.044 27.848 18.516 27.88 ;
  LAYER M2 ;
        RECT 16.044 27.784 18.516 27.816 ;
  LAYER M2 ;
        RECT 16.044 27.72 18.516 27.752 ;
  LAYER M2 ;
        RECT 16.044 27.656 18.516 27.688 ;
  LAYER M2 ;
        RECT 16.044 27.592 18.516 27.624 ;
  LAYER M2 ;
        RECT 16.044 27.528 18.516 27.56 ;
  LAYER M2 ;
        RECT 16.044 27.464 18.516 27.496 ;
  LAYER M2 ;
        RECT 16.044 27.4 18.516 27.432 ;
  LAYER M2 ;
        RECT 16.044 27.336 18.516 27.368 ;
  LAYER M2 ;
        RECT 16.044 27.272 18.516 27.304 ;
  LAYER M2 ;
        RECT 16.044 27.208 18.516 27.24 ;
  LAYER M2 ;
        RECT 16.044 27.144 18.516 27.176 ;
  LAYER M2 ;
        RECT 16.044 27.08 18.516 27.112 ;
  LAYER M2 ;
        RECT 16.044 27.016 18.516 27.048 ;
  LAYER M2 ;
        RECT 16.044 26.952 18.516 26.984 ;
  LAYER M2 ;
        RECT 16.044 26.888 18.516 26.92 ;
  LAYER M2 ;
        RECT 16.044 26.824 18.516 26.856 ;
  LAYER M2 ;
        RECT 16.044 26.76 18.516 26.792 ;
  LAYER M2 ;
        RECT 16.044 26.696 18.516 26.728 ;
  LAYER M2 ;
        RECT 16.044 26.632 18.516 26.664 ;
  LAYER M2 ;
        RECT 16.044 26.568 18.516 26.6 ;
  LAYER M2 ;
        RECT 16.044 26.504 18.516 26.536 ;
  LAYER M2 ;
        RECT 16.044 26.44 18.516 26.472 ;
  LAYER M2 ;
        RECT 16.044 26.376 18.516 26.408 ;
  LAYER M2 ;
        RECT 16.044 26.312 18.516 26.344 ;
  LAYER M2 ;
        RECT 16.044 26.248 18.516 26.28 ;
  LAYER M2 ;
        RECT 16.044 26.184 18.516 26.216 ;
  LAYER M2 ;
        RECT 16.044 26.12 18.516 26.152 ;
  LAYER M2 ;
        RECT 16.044 26.056 18.516 26.088 ;
  LAYER M2 ;
        RECT 16.044 25.992 18.516 26.024 ;
  LAYER M2 ;
        RECT 16.044 25.928 18.516 25.96 ;
  LAYER M2 ;
        RECT 16.044 25.864 18.516 25.896 ;
  LAYER M2 ;
        RECT 16.044 25.8 18.516 25.832 ;
  LAYER M2 ;
        RECT 16.044 25.736 18.516 25.768 ;
  LAYER M3 ;
        RECT 16.064 25.584 16.096 28.092 ;
  LAYER M3 ;
        RECT 16.128 25.584 16.16 28.092 ;
  LAYER M3 ;
        RECT 16.192 25.584 16.224 28.092 ;
  LAYER M3 ;
        RECT 16.256 25.584 16.288 28.092 ;
  LAYER M3 ;
        RECT 16.32 25.584 16.352 28.092 ;
  LAYER M3 ;
        RECT 16.384 25.584 16.416 28.092 ;
  LAYER M3 ;
        RECT 16.448 25.584 16.48 28.092 ;
  LAYER M3 ;
        RECT 16.512 25.584 16.544 28.092 ;
  LAYER M3 ;
        RECT 16.576 25.584 16.608 28.092 ;
  LAYER M3 ;
        RECT 16.64 25.584 16.672 28.092 ;
  LAYER M3 ;
        RECT 16.704 25.584 16.736 28.092 ;
  LAYER M3 ;
        RECT 16.768 25.584 16.8 28.092 ;
  LAYER M3 ;
        RECT 16.832 25.584 16.864 28.092 ;
  LAYER M3 ;
        RECT 16.896 25.584 16.928 28.092 ;
  LAYER M3 ;
        RECT 16.96 25.584 16.992 28.092 ;
  LAYER M3 ;
        RECT 17.024 25.584 17.056 28.092 ;
  LAYER M3 ;
        RECT 17.088 25.584 17.12 28.092 ;
  LAYER M3 ;
        RECT 17.152 25.584 17.184 28.092 ;
  LAYER M3 ;
        RECT 17.216 25.584 17.248 28.092 ;
  LAYER M3 ;
        RECT 17.28 25.584 17.312 28.092 ;
  LAYER M3 ;
        RECT 17.344 25.584 17.376 28.092 ;
  LAYER M3 ;
        RECT 17.408 25.584 17.44 28.092 ;
  LAYER M3 ;
        RECT 17.472 25.584 17.504 28.092 ;
  LAYER M3 ;
        RECT 17.536 25.584 17.568 28.092 ;
  LAYER M3 ;
        RECT 17.6 25.584 17.632 28.092 ;
  LAYER M3 ;
        RECT 17.664 25.584 17.696 28.092 ;
  LAYER M3 ;
        RECT 17.728 25.584 17.76 28.092 ;
  LAYER M3 ;
        RECT 17.792 25.584 17.824 28.092 ;
  LAYER M3 ;
        RECT 17.856 25.584 17.888 28.092 ;
  LAYER M3 ;
        RECT 17.92 25.584 17.952 28.092 ;
  LAYER M3 ;
        RECT 17.984 25.584 18.016 28.092 ;
  LAYER M3 ;
        RECT 18.048 25.584 18.08 28.092 ;
  LAYER M3 ;
        RECT 18.112 25.584 18.144 28.092 ;
  LAYER M3 ;
        RECT 18.176 25.584 18.208 28.092 ;
  LAYER M3 ;
        RECT 18.24 25.584 18.272 28.092 ;
  LAYER M3 ;
        RECT 18.304 25.584 18.336 28.092 ;
  LAYER M3 ;
        RECT 18.368 25.584 18.4 28.092 ;
  LAYER M3 ;
        RECT 18.464 25.584 18.496 28.092 ;
  LAYER M1 ;
        RECT 16.079 25.62 16.081 28.056 ;
  LAYER M1 ;
        RECT 16.159 25.62 16.161 28.056 ;
  LAYER M1 ;
        RECT 16.239 25.62 16.241 28.056 ;
  LAYER M1 ;
        RECT 16.319 25.62 16.321 28.056 ;
  LAYER M1 ;
        RECT 16.399 25.62 16.401 28.056 ;
  LAYER M1 ;
        RECT 16.479 25.62 16.481 28.056 ;
  LAYER M1 ;
        RECT 16.559 25.62 16.561 28.056 ;
  LAYER M1 ;
        RECT 16.639 25.62 16.641 28.056 ;
  LAYER M1 ;
        RECT 16.719 25.62 16.721 28.056 ;
  LAYER M1 ;
        RECT 16.799 25.62 16.801 28.056 ;
  LAYER M1 ;
        RECT 16.879 25.62 16.881 28.056 ;
  LAYER M1 ;
        RECT 16.959 25.62 16.961 28.056 ;
  LAYER M1 ;
        RECT 17.039 25.62 17.041 28.056 ;
  LAYER M1 ;
        RECT 17.119 25.62 17.121 28.056 ;
  LAYER M1 ;
        RECT 17.199 25.62 17.201 28.056 ;
  LAYER M1 ;
        RECT 17.279 25.62 17.281 28.056 ;
  LAYER M1 ;
        RECT 17.359 25.62 17.361 28.056 ;
  LAYER M1 ;
        RECT 17.439 25.62 17.441 28.056 ;
  LAYER M1 ;
        RECT 17.519 25.62 17.521 28.056 ;
  LAYER M1 ;
        RECT 17.599 25.62 17.601 28.056 ;
  LAYER M1 ;
        RECT 17.679 25.62 17.681 28.056 ;
  LAYER M1 ;
        RECT 17.759 25.62 17.761 28.056 ;
  LAYER M1 ;
        RECT 17.839 25.62 17.841 28.056 ;
  LAYER M1 ;
        RECT 17.919 25.62 17.921 28.056 ;
  LAYER M1 ;
        RECT 17.999 25.62 18.001 28.056 ;
  LAYER M1 ;
        RECT 18.079 25.62 18.081 28.056 ;
  LAYER M1 ;
        RECT 18.159 25.62 18.161 28.056 ;
  LAYER M1 ;
        RECT 18.239 25.62 18.241 28.056 ;
  LAYER M1 ;
        RECT 18.319 25.62 18.321 28.056 ;
  LAYER M1 ;
        RECT 18.399 25.62 18.401 28.056 ;
  LAYER M2 ;
        RECT 16.08 28.055 18.48 28.057 ;
  LAYER M2 ;
        RECT 16.08 27.971 18.48 27.973 ;
  LAYER M2 ;
        RECT 16.08 27.887 18.48 27.889 ;
  LAYER M2 ;
        RECT 16.08 27.803 18.48 27.805 ;
  LAYER M2 ;
        RECT 16.08 27.719 18.48 27.721 ;
  LAYER M2 ;
        RECT 16.08 27.635 18.48 27.637 ;
  LAYER M2 ;
        RECT 16.08 27.551 18.48 27.553 ;
  LAYER M2 ;
        RECT 16.08 27.467 18.48 27.469 ;
  LAYER M2 ;
        RECT 16.08 27.383 18.48 27.385 ;
  LAYER M2 ;
        RECT 16.08 27.299 18.48 27.301 ;
  LAYER M2 ;
        RECT 16.08 27.215 18.48 27.217 ;
  LAYER M2 ;
        RECT 16.08 27.131 18.48 27.133 ;
  LAYER M2 ;
        RECT 16.08 27.0475 18.48 27.0495 ;
  LAYER M2 ;
        RECT 16.08 26.963 18.48 26.965 ;
  LAYER M2 ;
        RECT 16.08 26.879 18.48 26.881 ;
  LAYER M2 ;
        RECT 16.08 26.795 18.48 26.797 ;
  LAYER M2 ;
        RECT 16.08 26.711 18.48 26.713 ;
  LAYER M2 ;
        RECT 16.08 26.627 18.48 26.629 ;
  LAYER M2 ;
        RECT 16.08 26.543 18.48 26.545 ;
  LAYER M2 ;
        RECT 16.08 26.459 18.48 26.461 ;
  LAYER M2 ;
        RECT 16.08 26.375 18.48 26.377 ;
  LAYER M2 ;
        RECT 16.08 26.291 18.48 26.293 ;
  LAYER M2 ;
        RECT 16.08 26.207 18.48 26.209 ;
  LAYER M2 ;
        RECT 16.08 26.123 18.48 26.125 ;
  LAYER M2 ;
        RECT 16.08 26.039 18.48 26.041 ;
  LAYER M2 ;
        RECT 16.08 25.955 18.48 25.957 ;
  LAYER M2 ;
        RECT 16.08 25.871 18.48 25.873 ;
  LAYER M2 ;
        RECT 16.08 25.787 18.48 25.789 ;
  LAYER M2 ;
        RECT 16.08 25.703 18.48 25.705 ;
  LAYER M1 ;
        RECT 16.064 22.644 16.096 25.152 ;
  LAYER M1 ;
        RECT 16.128 22.644 16.16 25.152 ;
  LAYER M1 ;
        RECT 16.192 22.644 16.224 25.152 ;
  LAYER M1 ;
        RECT 16.256 22.644 16.288 25.152 ;
  LAYER M1 ;
        RECT 16.32 22.644 16.352 25.152 ;
  LAYER M1 ;
        RECT 16.384 22.644 16.416 25.152 ;
  LAYER M1 ;
        RECT 16.448 22.644 16.48 25.152 ;
  LAYER M1 ;
        RECT 16.512 22.644 16.544 25.152 ;
  LAYER M1 ;
        RECT 16.576 22.644 16.608 25.152 ;
  LAYER M1 ;
        RECT 16.64 22.644 16.672 25.152 ;
  LAYER M1 ;
        RECT 16.704 22.644 16.736 25.152 ;
  LAYER M1 ;
        RECT 16.768 22.644 16.8 25.152 ;
  LAYER M1 ;
        RECT 16.832 22.644 16.864 25.152 ;
  LAYER M1 ;
        RECT 16.896 22.644 16.928 25.152 ;
  LAYER M1 ;
        RECT 16.96 22.644 16.992 25.152 ;
  LAYER M1 ;
        RECT 17.024 22.644 17.056 25.152 ;
  LAYER M1 ;
        RECT 17.088 22.644 17.12 25.152 ;
  LAYER M1 ;
        RECT 17.152 22.644 17.184 25.152 ;
  LAYER M1 ;
        RECT 17.216 22.644 17.248 25.152 ;
  LAYER M1 ;
        RECT 17.28 22.644 17.312 25.152 ;
  LAYER M1 ;
        RECT 17.344 22.644 17.376 25.152 ;
  LAYER M1 ;
        RECT 17.408 22.644 17.44 25.152 ;
  LAYER M1 ;
        RECT 17.472 22.644 17.504 25.152 ;
  LAYER M1 ;
        RECT 17.536 22.644 17.568 25.152 ;
  LAYER M1 ;
        RECT 17.6 22.644 17.632 25.152 ;
  LAYER M1 ;
        RECT 17.664 22.644 17.696 25.152 ;
  LAYER M1 ;
        RECT 17.728 22.644 17.76 25.152 ;
  LAYER M1 ;
        RECT 17.792 22.644 17.824 25.152 ;
  LAYER M1 ;
        RECT 17.856 22.644 17.888 25.152 ;
  LAYER M1 ;
        RECT 17.92 22.644 17.952 25.152 ;
  LAYER M1 ;
        RECT 17.984 22.644 18.016 25.152 ;
  LAYER M1 ;
        RECT 18.048 22.644 18.08 25.152 ;
  LAYER M1 ;
        RECT 18.112 22.644 18.144 25.152 ;
  LAYER M1 ;
        RECT 18.176 22.644 18.208 25.152 ;
  LAYER M1 ;
        RECT 18.24 22.644 18.272 25.152 ;
  LAYER M1 ;
        RECT 18.304 22.644 18.336 25.152 ;
  LAYER M1 ;
        RECT 18.368 22.644 18.4 25.152 ;
  LAYER M2 ;
        RECT 16.044 25.036 18.516 25.068 ;
  LAYER M2 ;
        RECT 16.044 24.972 18.516 25.004 ;
  LAYER M2 ;
        RECT 16.044 24.908 18.516 24.94 ;
  LAYER M2 ;
        RECT 16.044 24.844 18.516 24.876 ;
  LAYER M2 ;
        RECT 16.044 24.78 18.516 24.812 ;
  LAYER M2 ;
        RECT 16.044 24.716 18.516 24.748 ;
  LAYER M2 ;
        RECT 16.044 24.652 18.516 24.684 ;
  LAYER M2 ;
        RECT 16.044 24.588 18.516 24.62 ;
  LAYER M2 ;
        RECT 16.044 24.524 18.516 24.556 ;
  LAYER M2 ;
        RECT 16.044 24.46 18.516 24.492 ;
  LAYER M2 ;
        RECT 16.044 24.396 18.516 24.428 ;
  LAYER M2 ;
        RECT 16.044 24.332 18.516 24.364 ;
  LAYER M2 ;
        RECT 16.044 24.268 18.516 24.3 ;
  LAYER M2 ;
        RECT 16.044 24.204 18.516 24.236 ;
  LAYER M2 ;
        RECT 16.044 24.14 18.516 24.172 ;
  LAYER M2 ;
        RECT 16.044 24.076 18.516 24.108 ;
  LAYER M2 ;
        RECT 16.044 24.012 18.516 24.044 ;
  LAYER M2 ;
        RECT 16.044 23.948 18.516 23.98 ;
  LAYER M2 ;
        RECT 16.044 23.884 18.516 23.916 ;
  LAYER M2 ;
        RECT 16.044 23.82 18.516 23.852 ;
  LAYER M2 ;
        RECT 16.044 23.756 18.516 23.788 ;
  LAYER M2 ;
        RECT 16.044 23.692 18.516 23.724 ;
  LAYER M2 ;
        RECT 16.044 23.628 18.516 23.66 ;
  LAYER M2 ;
        RECT 16.044 23.564 18.516 23.596 ;
  LAYER M2 ;
        RECT 16.044 23.5 18.516 23.532 ;
  LAYER M2 ;
        RECT 16.044 23.436 18.516 23.468 ;
  LAYER M2 ;
        RECT 16.044 23.372 18.516 23.404 ;
  LAYER M2 ;
        RECT 16.044 23.308 18.516 23.34 ;
  LAYER M2 ;
        RECT 16.044 23.244 18.516 23.276 ;
  LAYER M2 ;
        RECT 16.044 23.18 18.516 23.212 ;
  LAYER M2 ;
        RECT 16.044 23.116 18.516 23.148 ;
  LAYER M2 ;
        RECT 16.044 23.052 18.516 23.084 ;
  LAYER M2 ;
        RECT 16.044 22.988 18.516 23.02 ;
  LAYER M2 ;
        RECT 16.044 22.924 18.516 22.956 ;
  LAYER M2 ;
        RECT 16.044 22.86 18.516 22.892 ;
  LAYER M2 ;
        RECT 16.044 22.796 18.516 22.828 ;
  LAYER M3 ;
        RECT 16.064 22.644 16.096 25.152 ;
  LAYER M3 ;
        RECT 16.128 22.644 16.16 25.152 ;
  LAYER M3 ;
        RECT 16.192 22.644 16.224 25.152 ;
  LAYER M3 ;
        RECT 16.256 22.644 16.288 25.152 ;
  LAYER M3 ;
        RECT 16.32 22.644 16.352 25.152 ;
  LAYER M3 ;
        RECT 16.384 22.644 16.416 25.152 ;
  LAYER M3 ;
        RECT 16.448 22.644 16.48 25.152 ;
  LAYER M3 ;
        RECT 16.512 22.644 16.544 25.152 ;
  LAYER M3 ;
        RECT 16.576 22.644 16.608 25.152 ;
  LAYER M3 ;
        RECT 16.64 22.644 16.672 25.152 ;
  LAYER M3 ;
        RECT 16.704 22.644 16.736 25.152 ;
  LAYER M3 ;
        RECT 16.768 22.644 16.8 25.152 ;
  LAYER M3 ;
        RECT 16.832 22.644 16.864 25.152 ;
  LAYER M3 ;
        RECT 16.896 22.644 16.928 25.152 ;
  LAYER M3 ;
        RECT 16.96 22.644 16.992 25.152 ;
  LAYER M3 ;
        RECT 17.024 22.644 17.056 25.152 ;
  LAYER M3 ;
        RECT 17.088 22.644 17.12 25.152 ;
  LAYER M3 ;
        RECT 17.152 22.644 17.184 25.152 ;
  LAYER M3 ;
        RECT 17.216 22.644 17.248 25.152 ;
  LAYER M3 ;
        RECT 17.28 22.644 17.312 25.152 ;
  LAYER M3 ;
        RECT 17.344 22.644 17.376 25.152 ;
  LAYER M3 ;
        RECT 17.408 22.644 17.44 25.152 ;
  LAYER M3 ;
        RECT 17.472 22.644 17.504 25.152 ;
  LAYER M3 ;
        RECT 17.536 22.644 17.568 25.152 ;
  LAYER M3 ;
        RECT 17.6 22.644 17.632 25.152 ;
  LAYER M3 ;
        RECT 17.664 22.644 17.696 25.152 ;
  LAYER M3 ;
        RECT 17.728 22.644 17.76 25.152 ;
  LAYER M3 ;
        RECT 17.792 22.644 17.824 25.152 ;
  LAYER M3 ;
        RECT 17.856 22.644 17.888 25.152 ;
  LAYER M3 ;
        RECT 17.92 22.644 17.952 25.152 ;
  LAYER M3 ;
        RECT 17.984 22.644 18.016 25.152 ;
  LAYER M3 ;
        RECT 18.048 22.644 18.08 25.152 ;
  LAYER M3 ;
        RECT 18.112 22.644 18.144 25.152 ;
  LAYER M3 ;
        RECT 18.176 22.644 18.208 25.152 ;
  LAYER M3 ;
        RECT 18.24 22.644 18.272 25.152 ;
  LAYER M3 ;
        RECT 18.304 22.644 18.336 25.152 ;
  LAYER M3 ;
        RECT 18.368 22.644 18.4 25.152 ;
  LAYER M3 ;
        RECT 18.464 22.644 18.496 25.152 ;
  LAYER M1 ;
        RECT 16.079 22.68 16.081 25.116 ;
  LAYER M1 ;
        RECT 16.159 22.68 16.161 25.116 ;
  LAYER M1 ;
        RECT 16.239 22.68 16.241 25.116 ;
  LAYER M1 ;
        RECT 16.319 22.68 16.321 25.116 ;
  LAYER M1 ;
        RECT 16.399 22.68 16.401 25.116 ;
  LAYER M1 ;
        RECT 16.479 22.68 16.481 25.116 ;
  LAYER M1 ;
        RECT 16.559 22.68 16.561 25.116 ;
  LAYER M1 ;
        RECT 16.639 22.68 16.641 25.116 ;
  LAYER M1 ;
        RECT 16.719 22.68 16.721 25.116 ;
  LAYER M1 ;
        RECT 16.799 22.68 16.801 25.116 ;
  LAYER M1 ;
        RECT 16.879 22.68 16.881 25.116 ;
  LAYER M1 ;
        RECT 16.959 22.68 16.961 25.116 ;
  LAYER M1 ;
        RECT 17.039 22.68 17.041 25.116 ;
  LAYER M1 ;
        RECT 17.119 22.68 17.121 25.116 ;
  LAYER M1 ;
        RECT 17.199 22.68 17.201 25.116 ;
  LAYER M1 ;
        RECT 17.279 22.68 17.281 25.116 ;
  LAYER M1 ;
        RECT 17.359 22.68 17.361 25.116 ;
  LAYER M1 ;
        RECT 17.439 22.68 17.441 25.116 ;
  LAYER M1 ;
        RECT 17.519 22.68 17.521 25.116 ;
  LAYER M1 ;
        RECT 17.599 22.68 17.601 25.116 ;
  LAYER M1 ;
        RECT 17.679 22.68 17.681 25.116 ;
  LAYER M1 ;
        RECT 17.759 22.68 17.761 25.116 ;
  LAYER M1 ;
        RECT 17.839 22.68 17.841 25.116 ;
  LAYER M1 ;
        RECT 17.919 22.68 17.921 25.116 ;
  LAYER M1 ;
        RECT 17.999 22.68 18.001 25.116 ;
  LAYER M1 ;
        RECT 18.079 22.68 18.081 25.116 ;
  LAYER M1 ;
        RECT 18.159 22.68 18.161 25.116 ;
  LAYER M1 ;
        RECT 18.239 22.68 18.241 25.116 ;
  LAYER M1 ;
        RECT 18.319 22.68 18.321 25.116 ;
  LAYER M1 ;
        RECT 18.399 22.68 18.401 25.116 ;
  LAYER M2 ;
        RECT 16.08 25.115 18.48 25.117 ;
  LAYER M2 ;
        RECT 16.08 25.031 18.48 25.033 ;
  LAYER M2 ;
        RECT 16.08 24.947 18.48 24.949 ;
  LAYER M2 ;
        RECT 16.08 24.863 18.48 24.865 ;
  LAYER M2 ;
        RECT 16.08 24.779 18.48 24.781 ;
  LAYER M2 ;
        RECT 16.08 24.695 18.48 24.697 ;
  LAYER M2 ;
        RECT 16.08 24.611 18.48 24.613 ;
  LAYER M2 ;
        RECT 16.08 24.527 18.48 24.529 ;
  LAYER M2 ;
        RECT 16.08 24.443 18.48 24.445 ;
  LAYER M2 ;
        RECT 16.08 24.359 18.48 24.361 ;
  LAYER M2 ;
        RECT 16.08 24.275 18.48 24.277 ;
  LAYER M2 ;
        RECT 16.08 24.191 18.48 24.193 ;
  LAYER M2 ;
        RECT 16.08 24.1075 18.48 24.1095 ;
  LAYER M2 ;
        RECT 16.08 24.023 18.48 24.025 ;
  LAYER M2 ;
        RECT 16.08 23.939 18.48 23.941 ;
  LAYER M2 ;
        RECT 16.08 23.855 18.48 23.857 ;
  LAYER M2 ;
        RECT 16.08 23.771 18.48 23.773 ;
  LAYER M2 ;
        RECT 16.08 23.687 18.48 23.689 ;
  LAYER M2 ;
        RECT 16.08 23.603 18.48 23.605 ;
  LAYER M2 ;
        RECT 16.08 23.519 18.48 23.521 ;
  LAYER M2 ;
        RECT 16.08 23.435 18.48 23.437 ;
  LAYER M2 ;
        RECT 16.08 23.351 18.48 23.353 ;
  LAYER M2 ;
        RECT 16.08 23.267 18.48 23.269 ;
  LAYER M2 ;
        RECT 16.08 23.183 18.48 23.185 ;
  LAYER M2 ;
        RECT 16.08 23.099 18.48 23.101 ;
  LAYER M2 ;
        RECT 16.08 23.015 18.48 23.017 ;
  LAYER M2 ;
        RECT 16.08 22.931 18.48 22.933 ;
  LAYER M2 ;
        RECT 16.08 22.847 18.48 22.849 ;
  LAYER M2 ;
        RECT 16.08 22.763 18.48 22.765 ;
  LAYER M1 ;
        RECT 16.064 19.704 16.096 22.212 ;
  LAYER M1 ;
        RECT 16.128 19.704 16.16 22.212 ;
  LAYER M1 ;
        RECT 16.192 19.704 16.224 22.212 ;
  LAYER M1 ;
        RECT 16.256 19.704 16.288 22.212 ;
  LAYER M1 ;
        RECT 16.32 19.704 16.352 22.212 ;
  LAYER M1 ;
        RECT 16.384 19.704 16.416 22.212 ;
  LAYER M1 ;
        RECT 16.448 19.704 16.48 22.212 ;
  LAYER M1 ;
        RECT 16.512 19.704 16.544 22.212 ;
  LAYER M1 ;
        RECT 16.576 19.704 16.608 22.212 ;
  LAYER M1 ;
        RECT 16.64 19.704 16.672 22.212 ;
  LAYER M1 ;
        RECT 16.704 19.704 16.736 22.212 ;
  LAYER M1 ;
        RECT 16.768 19.704 16.8 22.212 ;
  LAYER M1 ;
        RECT 16.832 19.704 16.864 22.212 ;
  LAYER M1 ;
        RECT 16.896 19.704 16.928 22.212 ;
  LAYER M1 ;
        RECT 16.96 19.704 16.992 22.212 ;
  LAYER M1 ;
        RECT 17.024 19.704 17.056 22.212 ;
  LAYER M1 ;
        RECT 17.088 19.704 17.12 22.212 ;
  LAYER M1 ;
        RECT 17.152 19.704 17.184 22.212 ;
  LAYER M1 ;
        RECT 17.216 19.704 17.248 22.212 ;
  LAYER M1 ;
        RECT 17.28 19.704 17.312 22.212 ;
  LAYER M1 ;
        RECT 17.344 19.704 17.376 22.212 ;
  LAYER M1 ;
        RECT 17.408 19.704 17.44 22.212 ;
  LAYER M1 ;
        RECT 17.472 19.704 17.504 22.212 ;
  LAYER M1 ;
        RECT 17.536 19.704 17.568 22.212 ;
  LAYER M1 ;
        RECT 17.6 19.704 17.632 22.212 ;
  LAYER M1 ;
        RECT 17.664 19.704 17.696 22.212 ;
  LAYER M1 ;
        RECT 17.728 19.704 17.76 22.212 ;
  LAYER M1 ;
        RECT 17.792 19.704 17.824 22.212 ;
  LAYER M1 ;
        RECT 17.856 19.704 17.888 22.212 ;
  LAYER M1 ;
        RECT 17.92 19.704 17.952 22.212 ;
  LAYER M1 ;
        RECT 17.984 19.704 18.016 22.212 ;
  LAYER M1 ;
        RECT 18.048 19.704 18.08 22.212 ;
  LAYER M1 ;
        RECT 18.112 19.704 18.144 22.212 ;
  LAYER M1 ;
        RECT 18.176 19.704 18.208 22.212 ;
  LAYER M1 ;
        RECT 18.24 19.704 18.272 22.212 ;
  LAYER M1 ;
        RECT 18.304 19.704 18.336 22.212 ;
  LAYER M1 ;
        RECT 18.368 19.704 18.4 22.212 ;
  LAYER M2 ;
        RECT 16.044 22.096 18.516 22.128 ;
  LAYER M2 ;
        RECT 16.044 22.032 18.516 22.064 ;
  LAYER M2 ;
        RECT 16.044 21.968 18.516 22 ;
  LAYER M2 ;
        RECT 16.044 21.904 18.516 21.936 ;
  LAYER M2 ;
        RECT 16.044 21.84 18.516 21.872 ;
  LAYER M2 ;
        RECT 16.044 21.776 18.516 21.808 ;
  LAYER M2 ;
        RECT 16.044 21.712 18.516 21.744 ;
  LAYER M2 ;
        RECT 16.044 21.648 18.516 21.68 ;
  LAYER M2 ;
        RECT 16.044 21.584 18.516 21.616 ;
  LAYER M2 ;
        RECT 16.044 21.52 18.516 21.552 ;
  LAYER M2 ;
        RECT 16.044 21.456 18.516 21.488 ;
  LAYER M2 ;
        RECT 16.044 21.392 18.516 21.424 ;
  LAYER M2 ;
        RECT 16.044 21.328 18.516 21.36 ;
  LAYER M2 ;
        RECT 16.044 21.264 18.516 21.296 ;
  LAYER M2 ;
        RECT 16.044 21.2 18.516 21.232 ;
  LAYER M2 ;
        RECT 16.044 21.136 18.516 21.168 ;
  LAYER M2 ;
        RECT 16.044 21.072 18.516 21.104 ;
  LAYER M2 ;
        RECT 16.044 21.008 18.516 21.04 ;
  LAYER M2 ;
        RECT 16.044 20.944 18.516 20.976 ;
  LAYER M2 ;
        RECT 16.044 20.88 18.516 20.912 ;
  LAYER M2 ;
        RECT 16.044 20.816 18.516 20.848 ;
  LAYER M2 ;
        RECT 16.044 20.752 18.516 20.784 ;
  LAYER M2 ;
        RECT 16.044 20.688 18.516 20.72 ;
  LAYER M2 ;
        RECT 16.044 20.624 18.516 20.656 ;
  LAYER M2 ;
        RECT 16.044 20.56 18.516 20.592 ;
  LAYER M2 ;
        RECT 16.044 20.496 18.516 20.528 ;
  LAYER M2 ;
        RECT 16.044 20.432 18.516 20.464 ;
  LAYER M2 ;
        RECT 16.044 20.368 18.516 20.4 ;
  LAYER M2 ;
        RECT 16.044 20.304 18.516 20.336 ;
  LAYER M2 ;
        RECT 16.044 20.24 18.516 20.272 ;
  LAYER M2 ;
        RECT 16.044 20.176 18.516 20.208 ;
  LAYER M2 ;
        RECT 16.044 20.112 18.516 20.144 ;
  LAYER M2 ;
        RECT 16.044 20.048 18.516 20.08 ;
  LAYER M2 ;
        RECT 16.044 19.984 18.516 20.016 ;
  LAYER M2 ;
        RECT 16.044 19.92 18.516 19.952 ;
  LAYER M2 ;
        RECT 16.044 19.856 18.516 19.888 ;
  LAYER M3 ;
        RECT 16.064 19.704 16.096 22.212 ;
  LAYER M3 ;
        RECT 16.128 19.704 16.16 22.212 ;
  LAYER M3 ;
        RECT 16.192 19.704 16.224 22.212 ;
  LAYER M3 ;
        RECT 16.256 19.704 16.288 22.212 ;
  LAYER M3 ;
        RECT 16.32 19.704 16.352 22.212 ;
  LAYER M3 ;
        RECT 16.384 19.704 16.416 22.212 ;
  LAYER M3 ;
        RECT 16.448 19.704 16.48 22.212 ;
  LAYER M3 ;
        RECT 16.512 19.704 16.544 22.212 ;
  LAYER M3 ;
        RECT 16.576 19.704 16.608 22.212 ;
  LAYER M3 ;
        RECT 16.64 19.704 16.672 22.212 ;
  LAYER M3 ;
        RECT 16.704 19.704 16.736 22.212 ;
  LAYER M3 ;
        RECT 16.768 19.704 16.8 22.212 ;
  LAYER M3 ;
        RECT 16.832 19.704 16.864 22.212 ;
  LAYER M3 ;
        RECT 16.896 19.704 16.928 22.212 ;
  LAYER M3 ;
        RECT 16.96 19.704 16.992 22.212 ;
  LAYER M3 ;
        RECT 17.024 19.704 17.056 22.212 ;
  LAYER M3 ;
        RECT 17.088 19.704 17.12 22.212 ;
  LAYER M3 ;
        RECT 17.152 19.704 17.184 22.212 ;
  LAYER M3 ;
        RECT 17.216 19.704 17.248 22.212 ;
  LAYER M3 ;
        RECT 17.28 19.704 17.312 22.212 ;
  LAYER M3 ;
        RECT 17.344 19.704 17.376 22.212 ;
  LAYER M3 ;
        RECT 17.408 19.704 17.44 22.212 ;
  LAYER M3 ;
        RECT 17.472 19.704 17.504 22.212 ;
  LAYER M3 ;
        RECT 17.536 19.704 17.568 22.212 ;
  LAYER M3 ;
        RECT 17.6 19.704 17.632 22.212 ;
  LAYER M3 ;
        RECT 17.664 19.704 17.696 22.212 ;
  LAYER M3 ;
        RECT 17.728 19.704 17.76 22.212 ;
  LAYER M3 ;
        RECT 17.792 19.704 17.824 22.212 ;
  LAYER M3 ;
        RECT 17.856 19.704 17.888 22.212 ;
  LAYER M3 ;
        RECT 17.92 19.704 17.952 22.212 ;
  LAYER M3 ;
        RECT 17.984 19.704 18.016 22.212 ;
  LAYER M3 ;
        RECT 18.048 19.704 18.08 22.212 ;
  LAYER M3 ;
        RECT 18.112 19.704 18.144 22.212 ;
  LAYER M3 ;
        RECT 18.176 19.704 18.208 22.212 ;
  LAYER M3 ;
        RECT 18.24 19.704 18.272 22.212 ;
  LAYER M3 ;
        RECT 18.304 19.704 18.336 22.212 ;
  LAYER M3 ;
        RECT 18.368 19.704 18.4 22.212 ;
  LAYER M3 ;
        RECT 18.464 19.704 18.496 22.212 ;
  LAYER M1 ;
        RECT 16.079 19.74 16.081 22.176 ;
  LAYER M1 ;
        RECT 16.159 19.74 16.161 22.176 ;
  LAYER M1 ;
        RECT 16.239 19.74 16.241 22.176 ;
  LAYER M1 ;
        RECT 16.319 19.74 16.321 22.176 ;
  LAYER M1 ;
        RECT 16.399 19.74 16.401 22.176 ;
  LAYER M1 ;
        RECT 16.479 19.74 16.481 22.176 ;
  LAYER M1 ;
        RECT 16.559 19.74 16.561 22.176 ;
  LAYER M1 ;
        RECT 16.639 19.74 16.641 22.176 ;
  LAYER M1 ;
        RECT 16.719 19.74 16.721 22.176 ;
  LAYER M1 ;
        RECT 16.799 19.74 16.801 22.176 ;
  LAYER M1 ;
        RECT 16.879 19.74 16.881 22.176 ;
  LAYER M1 ;
        RECT 16.959 19.74 16.961 22.176 ;
  LAYER M1 ;
        RECT 17.039 19.74 17.041 22.176 ;
  LAYER M1 ;
        RECT 17.119 19.74 17.121 22.176 ;
  LAYER M1 ;
        RECT 17.199 19.74 17.201 22.176 ;
  LAYER M1 ;
        RECT 17.279 19.74 17.281 22.176 ;
  LAYER M1 ;
        RECT 17.359 19.74 17.361 22.176 ;
  LAYER M1 ;
        RECT 17.439 19.74 17.441 22.176 ;
  LAYER M1 ;
        RECT 17.519 19.74 17.521 22.176 ;
  LAYER M1 ;
        RECT 17.599 19.74 17.601 22.176 ;
  LAYER M1 ;
        RECT 17.679 19.74 17.681 22.176 ;
  LAYER M1 ;
        RECT 17.759 19.74 17.761 22.176 ;
  LAYER M1 ;
        RECT 17.839 19.74 17.841 22.176 ;
  LAYER M1 ;
        RECT 17.919 19.74 17.921 22.176 ;
  LAYER M1 ;
        RECT 17.999 19.74 18.001 22.176 ;
  LAYER M1 ;
        RECT 18.079 19.74 18.081 22.176 ;
  LAYER M1 ;
        RECT 18.159 19.74 18.161 22.176 ;
  LAYER M1 ;
        RECT 18.239 19.74 18.241 22.176 ;
  LAYER M1 ;
        RECT 18.319 19.74 18.321 22.176 ;
  LAYER M1 ;
        RECT 18.399 19.74 18.401 22.176 ;
  LAYER M2 ;
        RECT 16.08 22.175 18.48 22.177 ;
  LAYER M2 ;
        RECT 16.08 22.091 18.48 22.093 ;
  LAYER M2 ;
        RECT 16.08 22.007 18.48 22.009 ;
  LAYER M2 ;
        RECT 16.08 21.923 18.48 21.925 ;
  LAYER M2 ;
        RECT 16.08 21.839 18.48 21.841 ;
  LAYER M2 ;
        RECT 16.08 21.755 18.48 21.757 ;
  LAYER M2 ;
        RECT 16.08 21.671 18.48 21.673 ;
  LAYER M2 ;
        RECT 16.08 21.587 18.48 21.589 ;
  LAYER M2 ;
        RECT 16.08 21.503 18.48 21.505 ;
  LAYER M2 ;
        RECT 16.08 21.419 18.48 21.421 ;
  LAYER M2 ;
        RECT 16.08 21.335 18.48 21.337 ;
  LAYER M2 ;
        RECT 16.08 21.251 18.48 21.253 ;
  LAYER M2 ;
        RECT 16.08 21.1675 18.48 21.1695 ;
  LAYER M2 ;
        RECT 16.08 21.083 18.48 21.085 ;
  LAYER M2 ;
        RECT 16.08 20.999 18.48 21.001 ;
  LAYER M2 ;
        RECT 16.08 20.915 18.48 20.917 ;
  LAYER M2 ;
        RECT 16.08 20.831 18.48 20.833 ;
  LAYER M2 ;
        RECT 16.08 20.747 18.48 20.749 ;
  LAYER M2 ;
        RECT 16.08 20.663 18.48 20.665 ;
  LAYER M2 ;
        RECT 16.08 20.579 18.48 20.581 ;
  LAYER M2 ;
        RECT 16.08 20.495 18.48 20.497 ;
  LAYER M2 ;
        RECT 16.08 20.411 18.48 20.413 ;
  LAYER M2 ;
        RECT 16.08 20.327 18.48 20.329 ;
  LAYER M2 ;
        RECT 16.08 20.243 18.48 20.245 ;
  LAYER M2 ;
        RECT 16.08 20.159 18.48 20.161 ;
  LAYER M2 ;
        RECT 16.08 20.075 18.48 20.077 ;
  LAYER M2 ;
        RECT 16.08 19.991 18.48 19.993 ;
  LAYER M2 ;
        RECT 16.08 19.907 18.48 19.909 ;
  LAYER M2 ;
        RECT 16.08 19.823 18.48 19.825 ;
  LAYER M1 ;
        RECT 18.944 34.404 18.976 36.912 ;
  LAYER M1 ;
        RECT 19.008 34.404 19.04 36.912 ;
  LAYER M1 ;
        RECT 19.072 34.404 19.104 36.912 ;
  LAYER M1 ;
        RECT 19.136 34.404 19.168 36.912 ;
  LAYER M1 ;
        RECT 19.2 34.404 19.232 36.912 ;
  LAYER M1 ;
        RECT 19.264 34.404 19.296 36.912 ;
  LAYER M1 ;
        RECT 19.328 34.404 19.36 36.912 ;
  LAYER M1 ;
        RECT 19.392 34.404 19.424 36.912 ;
  LAYER M1 ;
        RECT 19.456 34.404 19.488 36.912 ;
  LAYER M1 ;
        RECT 19.52 34.404 19.552 36.912 ;
  LAYER M1 ;
        RECT 19.584 34.404 19.616 36.912 ;
  LAYER M1 ;
        RECT 19.648 34.404 19.68 36.912 ;
  LAYER M1 ;
        RECT 19.712 34.404 19.744 36.912 ;
  LAYER M1 ;
        RECT 19.776 34.404 19.808 36.912 ;
  LAYER M1 ;
        RECT 19.84 34.404 19.872 36.912 ;
  LAYER M1 ;
        RECT 19.904 34.404 19.936 36.912 ;
  LAYER M1 ;
        RECT 19.968 34.404 20 36.912 ;
  LAYER M1 ;
        RECT 20.032 34.404 20.064 36.912 ;
  LAYER M1 ;
        RECT 20.096 34.404 20.128 36.912 ;
  LAYER M1 ;
        RECT 20.16 34.404 20.192 36.912 ;
  LAYER M1 ;
        RECT 20.224 34.404 20.256 36.912 ;
  LAYER M1 ;
        RECT 20.288 34.404 20.32 36.912 ;
  LAYER M1 ;
        RECT 20.352 34.404 20.384 36.912 ;
  LAYER M1 ;
        RECT 20.416 34.404 20.448 36.912 ;
  LAYER M1 ;
        RECT 20.48 34.404 20.512 36.912 ;
  LAYER M1 ;
        RECT 20.544 34.404 20.576 36.912 ;
  LAYER M1 ;
        RECT 20.608 34.404 20.64 36.912 ;
  LAYER M1 ;
        RECT 20.672 34.404 20.704 36.912 ;
  LAYER M1 ;
        RECT 20.736 34.404 20.768 36.912 ;
  LAYER M1 ;
        RECT 20.8 34.404 20.832 36.912 ;
  LAYER M1 ;
        RECT 20.864 34.404 20.896 36.912 ;
  LAYER M1 ;
        RECT 20.928 34.404 20.96 36.912 ;
  LAYER M1 ;
        RECT 20.992 34.404 21.024 36.912 ;
  LAYER M1 ;
        RECT 21.056 34.404 21.088 36.912 ;
  LAYER M1 ;
        RECT 21.12 34.404 21.152 36.912 ;
  LAYER M1 ;
        RECT 21.184 34.404 21.216 36.912 ;
  LAYER M1 ;
        RECT 21.248 34.404 21.28 36.912 ;
  LAYER M2 ;
        RECT 18.924 36.796 21.396 36.828 ;
  LAYER M2 ;
        RECT 18.924 36.732 21.396 36.764 ;
  LAYER M2 ;
        RECT 18.924 36.668 21.396 36.7 ;
  LAYER M2 ;
        RECT 18.924 36.604 21.396 36.636 ;
  LAYER M2 ;
        RECT 18.924 36.54 21.396 36.572 ;
  LAYER M2 ;
        RECT 18.924 36.476 21.396 36.508 ;
  LAYER M2 ;
        RECT 18.924 36.412 21.396 36.444 ;
  LAYER M2 ;
        RECT 18.924 36.348 21.396 36.38 ;
  LAYER M2 ;
        RECT 18.924 36.284 21.396 36.316 ;
  LAYER M2 ;
        RECT 18.924 36.22 21.396 36.252 ;
  LAYER M2 ;
        RECT 18.924 36.156 21.396 36.188 ;
  LAYER M2 ;
        RECT 18.924 36.092 21.396 36.124 ;
  LAYER M2 ;
        RECT 18.924 36.028 21.396 36.06 ;
  LAYER M2 ;
        RECT 18.924 35.964 21.396 35.996 ;
  LAYER M2 ;
        RECT 18.924 35.9 21.396 35.932 ;
  LAYER M2 ;
        RECT 18.924 35.836 21.396 35.868 ;
  LAYER M2 ;
        RECT 18.924 35.772 21.396 35.804 ;
  LAYER M2 ;
        RECT 18.924 35.708 21.396 35.74 ;
  LAYER M2 ;
        RECT 18.924 35.644 21.396 35.676 ;
  LAYER M2 ;
        RECT 18.924 35.58 21.396 35.612 ;
  LAYER M2 ;
        RECT 18.924 35.516 21.396 35.548 ;
  LAYER M2 ;
        RECT 18.924 35.452 21.396 35.484 ;
  LAYER M2 ;
        RECT 18.924 35.388 21.396 35.42 ;
  LAYER M2 ;
        RECT 18.924 35.324 21.396 35.356 ;
  LAYER M2 ;
        RECT 18.924 35.26 21.396 35.292 ;
  LAYER M2 ;
        RECT 18.924 35.196 21.396 35.228 ;
  LAYER M2 ;
        RECT 18.924 35.132 21.396 35.164 ;
  LAYER M2 ;
        RECT 18.924 35.068 21.396 35.1 ;
  LAYER M2 ;
        RECT 18.924 35.004 21.396 35.036 ;
  LAYER M2 ;
        RECT 18.924 34.94 21.396 34.972 ;
  LAYER M2 ;
        RECT 18.924 34.876 21.396 34.908 ;
  LAYER M2 ;
        RECT 18.924 34.812 21.396 34.844 ;
  LAYER M2 ;
        RECT 18.924 34.748 21.396 34.78 ;
  LAYER M2 ;
        RECT 18.924 34.684 21.396 34.716 ;
  LAYER M2 ;
        RECT 18.924 34.62 21.396 34.652 ;
  LAYER M2 ;
        RECT 18.924 34.556 21.396 34.588 ;
  LAYER M3 ;
        RECT 18.944 34.404 18.976 36.912 ;
  LAYER M3 ;
        RECT 19.008 34.404 19.04 36.912 ;
  LAYER M3 ;
        RECT 19.072 34.404 19.104 36.912 ;
  LAYER M3 ;
        RECT 19.136 34.404 19.168 36.912 ;
  LAYER M3 ;
        RECT 19.2 34.404 19.232 36.912 ;
  LAYER M3 ;
        RECT 19.264 34.404 19.296 36.912 ;
  LAYER M3 ;
        RECT 19.328 34.404 19.36 36.912 ;
  LAYER M3 ;
        RECT 19.392 34.404 19.424 36.912 ;
  LAYER M3 ;
        RECT 19.456 34.404 19.488 36.912 ;
  LAYER M3 ;
        RECT 19.52 34.404 19.552 36.912 ;
  LAYER M3 ;
        RECT 19.584 34.404 19.616 36.912 ;
  LAYER M3 ;
        RECT 19.648 34.404 19.68 36.912 ;
  LAYER M3 ;
        RECT 19.712 34.404 19.744 36.912 ;
  LAYER M3 ;
        RECT 19.776 34.404 19.808 36.912 ;
  LAYER M3 ;
        RECT 19.84 34.404 19.872 36.912 ;
  LAYER M3 ;
        RECT 19.904 34.404 19.936 36.912 ;
  LAYER M3 ;
        RECT 19.968 34.404 20 36.912 ;
  LAYER M3 ;
        RECT 20.032 34.404 20.064 36.912 ;
  LAYER M3 ;
        RECT 20.096 34.404 20.128 36.912 ;
  LAYER M3 ;
        RECT 20.16 34.404 20.192 36.912 ;
  LAYER M3 ;
        RECT 20.224 34.404 20.256 36.912 ;
  LAYER M3 ;
        RECT 20.288 34.404 20.32 36.912 ;
  LAYER M3 ;
        RECT 20.352 34.404 20.384 36.912 ;
  LAYER M3 ;
        RECT 20.416 34.404 20.448 36.912 ;
  LAYER M3 ;
        RECT 20.48 34.404 20.512 36.912 ;
  LAYER M3 ;
        RECT 20.544 34.404 20.576 36.912 ;
  LAYER M3 ;
        RECT 20.608 34.404 20.64 36.912 ;
  LAYER M3 ;
        RECT 20.672 34.404 20.704 36.912 ;
  LAYER M3 ;
        RECT 20.736 34.404 20.768 36.912 ;
  LAYER M3 ;
        RECT 20.8 34.404 20.832 36.912 ;
  LAYER M3 ;
        RECT 20.864 34.404 20.896 36.912 ;
  LAYER M3 ;
        RECT 20.928 34.404 20.96 36.912 ;
  LAYER M3 ;
        RECT 20.992 34.404 21.024 36.912 ;
  LAYER M3 ;
        RECT 21.056 34.404 21.088 36.912 ;
  LAYER M3 ;
        RECT 21.12 34.404 21.152 36.912 ;
  LAYER M3 ;
        RECT 21.184 34.404 21.216 36.912 ;
  LAYER M3 ;
        RECT 21.248 34.404 21.28 36.912 ;
  LAYER M3 ;
        RECT 21.344 34.404 21.376 36.912 ;
  LAYER M1 ;
        RECT 18.959 34.44 18.961 36.876 ;
  LAYER M1 ;
        RECT 19.039 34.44 19.041 36.876 ;
  LAYER M1 ;
        RECT 19.119 34.44 19.121 36.876 ;
  LAYER M1 ;
        RECT 19.199 34.44 19.201 36.876 ;
  LAYER M1 ;
        RECT 19.279 34.44 19.281 36.876 ;
  LAYER M1 ;
        RECT 19.359 34.44 19.361 36.876 ;
  LAYER M1 ;
        RECT 19.439 34.44 19.441 36.876 ;
  LAYER M1 ;
        RECT 19.519 34.44 19.521 36.876 ;
  LAYER M1 ;
        RECT 19.599 34.44 19.601 36.876 ;
  LAYER M1 ;
        RECT 19.679 34.44 19.681 36.876 ;
  LAYER M1 ;
        RECT 19.759 34.44 19.761 36.876 ;
  LAYER M1 ;
        RECT 19.839 34.44 19.841 36.876 ;
  LAYER M1 ;
        RECT 19.919 34.44 19.921 36.876 ;
  LAYER M1 ;
        RECT 19.999 34.44 20.001 36.876 ;
  LAYER M1 ;
        RECT 20.079 34.44 20.081 36.876 ;
  LAYER M1 ;
        RECT 20.159 34.44 20.161 36.876 ;
  LAYER M1 ;
        RECT 20.239 34.44 20.241 36.876 ;
  LAYER M1 ;
        RECT 20.319 34.44 20.321 36.876 ;
  LAYER M1 ;
        RECT 20.399 34.44 20.401 36.876 ;
  LAYER M1 ;
        RECT 20.479 34.44 20.481 36.876 ;
  LAYER M1 ;
        RECT 20.559 34.44 20.561 36.876 ;
  LAYER M1 ;
        RECT 20.639 34.44 20.641 36.876 ;
  LAYER M1 ;
        RECT 20.719 34.44 20.721 36.876 ;
  LAYER M1 ;
        RECT 20.799 34.44 20.801 36.876 ;
  LAYER M1 ;
        RECT 20.879 34.44 20.881 36.876 ;
  LAYER M1 ;
        RECT 20.959 34.44 20.961 36.876 ;
  LAYER M1 ;
        RECT 21.039 34.44 21.041 36.876 ;
  LAYER M1 ;
        RECT 21.119 34.44 21.121 36.876 ;
  LAYER M1 ;
        RECT 21.199 34.44 21.201 36.876 ;
  LAYER M1 ;
        RECT 21.279 34.44 21.281 36.876 ;
  LAYER M2 ;
        RECT 18.96 36.875 21.36 36.877 ;
  LAYER M2 ;
        RECT 18.96 36.791 21.36 36.793 ;
  LAYER M2 ;
        RECT 18.96 36.707 21.36 36.709 ;
  LAYER M2 ;
        RECT 18.96 36.623 21.36 36.625 ;
  LAYER M2 ;
        RECT 18.96 36.539 21.36 36.541 ;
  LAYER M2 ;
        RECT 18.96 36.455 21.36 36.457 ;
  LAYER M2 ;
        RECT 18.96 36.371 21.36 36.373 ;
  LAYER M2 ;
        RECT 18.96 36.287 21.36 36.289 ;
  LAYER M2 ;
        RECT 18.96 36.203 21.36 36.205 ;
  LAYER M2 ;
        RECT 18.96 36.119 21.36 36.121 ;
  LAYER M2 ;
        RECT 18.96 36.035 21.36 36.037 ;
  LAYER M2 ;
        RECT 18.96 35.951 21.36 35.953 ;
  LAYER M2 ;
        RECT 18.96 35.8675 21.36 35.8695 ;
  LAYER M2 ;
        RECT 18.96 35.783 21.36 35.785 ;
  LAYER M2 ;
        RECT 18.96 35.699 21.36 35.701 ;
  LAYER M2 ;
        RECT 18.96 35.615 21.36 35.617 ;
  LAYER M2 ;
        RECT 18.96 35.531 21.36 35.533 ;
  LAYER M2 ;
        RECT 18.96 35.447 21.36 35.449 ;
  LAYER M2 ;
        RECT 18.96 35.363 21.36 35.365 ;
  LAYER M2 ;
        RECT 18.96 35.279 21.36 35.281 ;
  LAYER M2 ;
        RECT 18.96 35.195 21.36 35.197 ;
  LAYER M2 ;
        RECT 18.96 35.111 21.36 35.113 ;
  LAYER M2 ;
        RECT 18.96 35.027 21.36 35.029 ;
  LAYER M2 ;
        RECT 18.96 34.943 21.36 34.945 ;
  LAYER M2 ;
        RECT 18.96 34.859 21.36 34.861 ;
  LAYER M2 ;
        RECT 18.96 34.775 21.36 34.777 ;
  LAYER M2 ;
        RECT 18.96 34.691 21.36 34.693 ;
  LAYER M2 ;
        RECT 18.96 34.607 21.36 34.609 ;
  LAYER M2 ;
        RECT 18.96 34.523 21.36 34.525 ;
  LAYER M1 ;
        RECT 18.944 31.464 18.976 33.972 ;
  LAYER M1 ;
        RECT 19.008 31.464 19.04 33.972 ;
  LAYER M1 ;
        RECT 19.072 31.464 19.104 33.972 ;
  LAYER M1 ;
        RECT 19.136 31.464 19.168 33.972 ;
  LAYER M1 ;
        RECT 19.2 31.464 19.232 33.972 ;
  LAYER M1 ;
        RECT 19.264 31.464 19.296 33.972 ;
  LAYER M1 ;
        RECT 19.328 31.464 19.36 33.972 ;
  LAYER M1 ;
        RECT 19.392 31.464 19.424 33.972 ;
  LAYER M1 ;
        RECT 19.456 31.464 19.488 33.972 ;
  LAYER M1 ;
        RECT 19.52 31.464 19.552 33.972 ;
  LAYER M1 ;
        RECT 19.584 31.464 19.616 33.972 ;
  LAYER M1 ;
        RECT 19.648 31.464 19.68 33.972 ;
  LAYER M1 ;
        RECT 19.712 31.464 19.744 33.972 ;
  LAYER M1 ;
        RECT 19.776 31.464 19.808 33.972 ;
  LAYER M1 ;
        RECT 19.84 31.464 19.872 33.972 ;
  LAYER M1 ;
        RECT 19.904 31.464 19.936 33.972 ;
  LAYER M1 ;
        RECT 19.968 31.464 20 33.972 ;
  LAYER M1 ;
        RECT 20.032 31.464 20.064 33.972 ;
  LAYER M1 ;
        RECT 20.096 31.464 20.128 33.972 ;
  LAYER M1 ;
        RECT 20.16 31.464 20.192 33.972 ;
  LAYER M1 ;
        RECT 20.224 31.464 20.256 33.972 ;
  LAYER M1 ;
        RECT 20.288 31.464 20.32 33.972 ;
  LAYER M1 ;
        RECT 20.352 31.464 20.384 33.972 ;
  LAYER M1 ;
        RECT 20.416 31.464 20.448 33.972 ;
  LAYER M1 ;
        RECT 20.48 31.464 20.512 33.972 ;
  LAYER M1 ;
        RECT 20.544 31.464 20.576 33.972 ;
  LAYER M1 ;
        RECT 20.608 31.464 20.64 33.972 ;
  LAYER M1 ;
        RECT 20.672 31.464 20.704 33.972 ;
  LAYER M1 ;
        RECT 20.736 31.464 20.768 33.972 ;
  LAYER M1 ;
        RECT 20.8 31.464 20.832 33.972 ;
  LAYER M1 ;
        RECT 20.864 31.464 20.896 33.972 ;
  LAYER M1 ;
        RECT 20.928 31.464 20.96 33.972 ;
  LAYER M1 ;
        RECT 20.992 31.464 21.024 33.972 ;
  LAYER M1 ;
        RECT 21.056 31.464 21.088 33.972 ;
  LAYER M1 ;
        RECT 21.12 31.464 21.152 33.972 ;
  LAYER M1 ;
        RECT 21.184 31.464 21.216 33.972 ;
  LAYER M1 ;
        RECT 21.248 31.464 21.28 33.972 ;
  LAYER M2 ;
        RECT 18.924 33.856 21.396 33.888 ;
  LAYER M2 ;
        RECT 18.924 33.792 21.396 33.824 ;
  LAYER M2 ;
        RECT 18.924 33.728 21.396 33.76 ;
  LAYER M2 ;
        RECT 18.924 33.664 21.396 33.696 ;
  LAYER M2 ;
        RECT 18.924 33.6 21.396 33.632 ;
  LAYER M2 ;
        RECT 18.924 33.536 21.396 33.568 ;
  LAYER M2 ;
        RECT 18.924 33.472 21.396 33.504 ;
  LAYER M2 ;
        RECT 18.924 33.408 21.396 33.44 ;
  LAYER M2 ;
        RECT 18.924 33.344 21.396 33.376 ;
  LAYER M2 ;
        RECT 18.924 33.28 21.396 33.312 ;
  LAYER M2 ;
        RECT 18.924 33.216 21.396 33.248 ;
  LAYER M2 ;
        RECT 18.924 33.152 21.396 33.184 ;
  LAYER M2 ;
        RECT 18.924 33.088 21.396 33.12 ;
  LAYER M2 ;
        RECT 18.924 33.024 21.396 33.056 ;
  LAYER M2 ;
        RECT 18.924 32.96 21.396 32.992 ;
  LAYER M2 ;
        RECT 18.924 32.896 21.396 32.928 ;
  LAYER M2 ;
        RECT 18.924 32.832 21.396 32.864 ;
  LAYER M2 ;
        RECT 18.924 32.768 21.396 32.8 ;
  LAYER M2 ;
        RECT 18.924 32.704 21.396 32.736 ;
  LAYER M2 ;
        RECT 18.924 32.64 21.396 32.672 ;
  LAYER M2 ;
        RECT 18.924 32.576 21.396 32.608 ;
  LAYER M2 ;
        RECT 18.924 32.512 21.396 32.544 ;
  LAYER M2 ;
        RECT 18.924 32.448 21.396 32.48 ;
  LAYER M2 ;
        RECT 18.924 32.384 21.396 32.416 ;
  LAYER M2 ;
        RECT 18.924 32.32 21.396 32.352 ;
  LAYER M2 ;
        RECT 18.924 32.256 21.396 32.288 ;
  LAYER M2 ;
        RECT 18.924 32.192 21.396 32.224 ;
  LAYER M2 ;
        RECT 18.924 32.128 21.396 32.16 ;
  LAYER M2 ;
        RECT 18.924 32.064 21.396 32.096 ;
  LAYER M2 ;
        RECT 18.924 32 21.396 32.032 ;
  LAYER M2 ;
        RECT 18.924 31.936 21.396 31.968 ;
  LAYER M2 ;
        RECT 18.924 31.872 21.396 31.904 ;
  LAYER M2 ;
        RECT 18.924 31.808 21.396 31.84 ;
  LAYER M2 ;
        RECT 18.924 31.744 21.396 31.776 ;
  LAYER M2 ;
        RECT 18.924 31.68 21.396 31.712 ;
  LAYER M2 ;
        RECT 18.924 31.616 21.396 31.648 ;
  LAYER M3 ;
        RECT 18.944 31.464 18.976 33.972 ;
  LAYER M3 ;
        RECT 19.008 31.464 19.04 33.972 ;
  LAYER M3 ;
        RECT 19.072 31.464 19.104 33.972 ;
  LAYER M3 ;
        RECT 19.136 31.464 19.168 33.972 ;
  LAYER M3 ;
        RECT 19.2 31.464 19.232 33.972 ;
  LAYER M3 ;
        RECT 19.264 31.464 19.296 33.972 ;
  LAYER M3 ;
        RECT 19.328 31.464 19.36 33.972 ;
  LAYER M3 ;
        RECT 19.392 31.464 19.424 33.972 ;
  LAYER M3 ;
        RECT 19.456 31.464 19.488 33.972 ;
  LAYER M3 ;
        RECT 19.52 31.464 19.552 33.972 ;
  LAYER M3 ;
        RECT 19.584 31.464 19.616 33.972 ;
  LAYER M3 ;
        RECT 19.648 31.464 19.68 33.972 ;
  LAYER M3 ;
        RECT 19.712 31.464 19.744 33.972 ;
  LAYER M3 ;
        RECT 19.776 31.464 19.808 33.972 ;
  LAYER M3 ;
        RECT 19.84 31.464 19.872 33.972 ;
  LAYER M3 ;
        RECT 19.904 31.464 19.936 33.972 ;
  LAYER M3 ;
        RECT 19.968 31.464 20 33.972 ;
  LAYER M3 ;
        RECT 20.032 31.464 20.064 33.972 ;
  LAYER M3 ;
        RECT 20.096 31.464 20.128 33.972 ;
  LAYER M3 ;
        RECT 20.16 31.464 20.192 33.972 ;
  LAYER M3 ;
        RECT 20.224 31.464 20.256 33.972 ;
  LAYER M3 ;
        RECT 20.288 31.464 20.32 33.972 ;
  LAYER M3 ;
        RECT 20.352 31.464 20.384 33.972 ;
  LAYER M3 ;
        RECT 20.416 31.464 20.448 33.972 ;
  LAYER M3 ;
        RECT 20.48 31.464 20.512 33.972 ;
  LAYER M3 ;
        RECT 20.544 31.464 20.576 33.972 ;
  LAYER M3 ;
        RECT 20.608 31.464 20.64 33.972 ;
  LAYER M3 ;
        RECT 20.672 31.464 20.704 33.972 ;
  LAYER M3 ;
        RECT 20.736 31.464 20.768 33.972 ;
  LAYER M3 ;
        RECT 20.8 31.464 20.832 33.972 ;
  LAYER M3 ;
        RECT 20.864 31.464 20.896 33.972 ;
  LAYER M3 ;
        RECT 20.928 31.464 20.96 33.972 ;
  LAYER M3 ;
        RECT 20.992 31.464 21.024 33.972 ;
  LAYER M3 ;
        RECT 21.056 31.464 21.088 33.972 ;
  LAYER M3 ;
        RECT 21.12 31.464 21.152 33.972 ;
  LAYER M3 ;
        RECT 21.184 31.464 21.216 33.972 ;
  LAYER M3 ;
        RECT 21.248 31.464 21.28 33.972 ;
  LAYER M3 ;
        RECT 21.344 31.464 21.376 33.972 ;
  LAYER M1 ;
        RECT 18.959 31.5 18.961 33.936 ;
  LAYER M1 ;
        RECT 19.039 31.5 19.041 33.936 ;
  LAYER M1 ;
        RECT 19.119 31.5 19.121 33.936 ;
  LAYER M1 ;
        RECT 19.199 31.5 19.201 33.936 ;
  LAYER M1 ;
        RECT 19.279 31.5 19.281 33.936 ;
  LAYER M1 ;
        RECT 19.359 31.5 19.361 33.936 ;
  LAYER M1 ;
        RECT 19.439 31.5 19.441 33.936 ;
  LAYER M1 ;
        RECT 19.519 31.5 19.521 33.936 ;
  LAYER M1 ;
        RECT 19.599 31.5 19.601 33.936 ;
  LAYER M1 ;
        RECT 19.679 31.5 19.681 33.936 ;
  LAYER M1 ;
        RECT 19.759 31.5 19.761 33.936 ;
  LAYER M1 ;
        RECT 19.839 31.5 19.841 33.936 ;
  LAYER M1 ;
        RECT 19.919 31.5 19.921 33.936 ;
  LAYER M1 ;
        RECT 19.999 31.5 20.001 33.936 ;
  LAYER M1 ;
        RECT 20.079 31.5 20.081 33.936 ;
  LAYER M1 ;
        RECT 20.159 31.5 20.161 33.936 ;
  LAYER M1 ;
        RECT 20.239 31.5 20.241 33.936 ;
  LAYER M1 ;
        RECT 20.319 31.5 20.321 33.936 ;
  LAYER M1 ;
        RECT 20.399 31.5 20.401 33.936 ;
  LAYER M1 ;
        RECT 20.479 31.5 20.481 33.936 ;
  LAYER M1 ;
        RECT 20.559 31.5 20.561 33.936 ;
  LAYER M1 ;
        RECT 20.639 31.5 20.641 33.936 ;
  LAYER M1 ;
        RECT 20.719 31.5 20.721 33.936 ;
  LAYER M1 ;
        RECT 20.799 31.5 20.801 33.936 ;
  LAYER M1 ;
        RECT 20.879 31.5 20.881 33.936 ;
  LAYER M1 ;
        RECT 20.959 31.5 20.961 33.936 ;
  LAYER M1 ;
        RECT 21.039 31.5 21.041 33.936 ;
  LAYER M1 ;
        RECT 21.119 31.5 21.121 33.936 ;
  LAYER M1 ;
        RECT 21.199 31.5 21.201 33.936 ;
  LAYER M1 ;
        RECT 21.279 31.5 21.281 33.936 ;
  LAYER M2 ;
        RECT 18.96 33.935 21.36 33.937 ;
  LAYER M2 ;
        RECT 18.96 33.851 21.36 33.853 ;
  LAYER M2 ;
        RECT 18.96 33.767 21.36 33.769 ;
  LAYER M2 ;
        RECT 18.96 33.683 21.36 33.685 ;
  LAYER M2 ;
        RECT 18.96 33.599 21.36 33.601 ;
  LAYER M2 ;
        RECT 18.96 33.515 21.36 33.517 ;
  LAYER M2 ;
        RECT 18.96 33.431 21.36 33.433 ;
  LAYER M2 ;
        RECT 18.96 33.347 21.36 33.349 ;
  LAYER M2 ;
        RECT 18.96 33.263 21.36 33.265 ;
  LAYER M2 ;
        RECT 18.96 33.179 21.36 33.181 ;
  LAYER M2 ;
        RECT 18.96 33.095 21.36 33.097 ;
  LAYER M2 ;
        RECT 18.96 33.011 21.36 33.013 ;
  LAYER M2 ;
        RECT 18.96 32.9275 21.36 32.9295 ;
  LAYER M2 ;
        RECT 18.96 32.843 21.36 32.845 ;
  LAYER M2 ;
        RECT 18.96 32.759 21.36 32.761 ;
  LAYER M2 ;
        RECT 18.96 32.675 21.36 32.677 ;
  LAYER M2 ;
        RECT 18.96 32.591 21.36 32.593 ;
  LAYER M2 ;
        RECT 18.96 32.507 21.36 32.509 ;
  LAYER M2 ;
        RECT 18.96 32.423 21.36 32.425 ;
  LAYER M2 ;
        RECT 18.96 32.339 21.36 32.341 ;
  LAYER M2 ;
        RECT 18.96 32.255 21.36 32.257 ;
  LAYER M2 ;
        RECT 18.96 32.171 21.36 32.173 ;
  LAYER M2 ;
        RECT 18.96 32.087 21.36 32.089 ;
  LAYER M2 ;
        RECT 18.96 32.003 21.36 32.005 ;
  LAYER M2 ;
        RECT 18.96 31.919 21.36 31.921 ;
  LAYER M2 ;
        RECT 18.96 31.835 21.36 31.837 ;
  LAYER M2 ;
        RECT 18.96 31.751 21.36 31.753 ;
  LAYER M2 ;
        RECT 18.96 31.667 21.36 31.669 ;
  LAYER M2 ;
        RECT 18.96 31.583 21.36 31.585 ;
  LAYER M1 ;
        RECT 18.944 28.524 18.976 31.032 ;
  LAYER M1 ;
        RECT 19.008 28.524 19.04 31.032 ;
  LAYER M1 ;
        RECT 19.072 28.524 19.104 31.032 ;
  LAYER M1 ;
        RECT 19.136 28.524 19.168 31.032 ;
  LAYER M1 ;
        RECT 19.2 28.524 19.232 31.032 ;
  LAYER M1 ;
        RECT 19.264 28.524 19.296 31.032 ;
  LAYER M1 ;
        RECT 19.328 28.524 19.36 31.032 ;
  LAYER M1 ;
        RECT 19.392 28.524 19.424 31.032 ;
  LAYER M1 ;
        RECT 19.456 28.524 19.488 31.032 ;
  LAYER M1 ;
        RECT 19.52 28.524 19.552 31.032 ;
  LAYER M1 ;
        RECT 19.584 28.524 19.616 31.032 ;
  LAYER M1 ;
        RECT 19.648 28.524 19.68 31.032 ;
  LAYER M1 ;
        RECT 19.712 28.524 19.744 31.032 ;
  LAYER M1 ;
        RECT 19.776 28.524 19.808 31.032 ;
  LAYER M1 ;
        RECT 19.84 28.524 19.872 31.032 ;
  LAYER M1 ;
        RECT 19.904 28.524 19.936 31.032 ;
  LAYER M1 ;
        RECT 19.968 28.524 20 31.032 ;
  LAYER M1 ;
        RECT 20.032 28.524 20.064 31.032 ;
  LAYER M1 ;
        RECT 20.096 28.524 20.128 31.032 ;
  LAYER M1 ;
        RECT 20.16 28.524 20.192 31.032 ;
  LAYER M1 ;
        RECT 20.224 28.524 20.256 31.032 ;
  LAYER M1 ;
        RECT 20.288 28.524 20.32 31.032 ;
  LAYER M1 ;
        RECT 20.352 28.524 20.384 31.032 ;
  LAYER M1 ;
        RECT 20.416 28.524 20.448 31.032 ;
  LAYER M1 ;
        RECT 20.48 28.524 20.512 31.032 ;
  LAYER M1 ;
        RECT 20.544 28.524 20.576 31.032 ;
  LAYER M1 ;
        RECT 20.608 28.524 20.64 31.032 ;
  LAYER M1 ;
        RECT 20.672 28.524 20.704 31.032 ;
  LAYER M1 ;
        RECT 20.736 28.524 20.768 31.032 ;
  LAYER M1 ;
        RECT 20.8 28.524 20.832 31.032 ;
  LAYER M1 ;
        RECT 20.864 28.524 20.896 31.032 ;
  LAYER M1 ;
        RECT 20.928 28.524 20.96 31.032 ;
  LAYER M1 ;
        RECT 20.992 28.524 21.024 31.032 ;
  LAYER M1 ;
        RECT 21.056 28.524 21.088 31.032 ;
  LAYER M1 ;
        RECT 21.12 28.524 21.152 31.032 ;
  LAYER M1 ;
        RECT 21.184 28.524 21.216 31.032 ;
  LAYER M1 ;
        RECT 21.248 28.524 21.28 31.032 ;
  LAYER M2 ;
        RECT 18.924 30.916 21.396 30.948 ;
  LAYER M2 ;
        RECT 18.924 30.852 21.396 30.884 ;
  LAYER M2 ;
        RECT 18.924 30.788 21.396 30.82 ;
  LAYER M2 ;
        RECT 18.924 30.724 21.396 30.756 ;
  LAYER M2 ;
        RECT 18.924 30.66 21.396 30.692 ;
  LAYER M2 ;
        RECT 18.924 30.596 21.396 30.628 ;
  LAYER M2 ;
        RECT 18.924 30.532 21.396 30.564 ;
  LAYER M2 ;
        RECT 18.924 30.468 21.396 30.5 ;
  LAYER M2 ;
        RECT 18.924 30.404 21.396 30.436 ;
  LAYER M2 ;
        RECT 18.924 30.34 21.396 30.372 ;
  LAYER M2 ;
        RECT 18.924 30.276 21.396 30.308 ;
  LAYER M2 ;
        RECT 18.924 30.212 21.396 30.244 ;
  LAYER M2 ;
        RECT 18.924 30.148 21.396 30.18 ;
  LAYER M2 ;
        RECT 18.924 30.084 21.396 30.116 ;
  LAYER M2 ;
        RECT 18.924 30.02 21.396 30.052 ;
  LAYER M2 ;
        RECT 18.924 29.956 21.396 29.988 ;
  LAYER M2 ;
        RECT 18.924 29.892 21.396 29.924 ;
  LAYER M2 ;
        RECT 18.924 29.828 21.396 29.86 ;
  LAYER M2 ;
        RECT 18.924 29.764 21.396 29.796 ;
  LAYER M2 ;
        RECT 18.924 29.7 21.396 29.732 ;
  LAYER M2 ;
        RECT 18.924 29.636 21.396 29.668 ;
  LAYER M2 ;
        RECT 18.924 29.572 21.396 29.604 ;
  LAYER M2 ;
        RECT 18.924 29.508 21.396 29.54 ;
  LAYER M2 ;
        RECT 18.924 29.444 21.396 29.476 ;
  LAYER M2 ;
        RECT 18.924 29.38 21.396 29.412 ;
  LAYER M2 ;
        RECT 18.924 29.316 21.396 29.348 ;
  LAYER M2 ;
        RECT 18.924 29.252 21.396 29.284 ;
  LAYER M2 ;
        RECT 18.924 29.188 21.396 29.22 ;
  LAYER M2 ;
        RECT 18.924 29.124 21.396 29.156 ;
  LAYER M2 ;
        RECT 18.924 29.06 21.396 29.092 ;
  LAYER M2 ;
        RECT 18.924 28.996 21.396 29.028 ;
  LAYER M2 ;
        RECT 18.924 28.932 21.396 28.964 ;
  LAYER M2 ;
        RECT 18.924 28.868 21.396 28.9 ;
  LAYER M2 ;
        RECT 18.924 28.804 21.396 28.836 ;
  LAYER M2 ;
        RECT 18.924 28.74 21.396 28.772 ;
  LAYER M2 ;
        RECT 18.924 28.676 21.396 28.708 ;
  LAYER M3 ;
        RECT 18.944 28.524 18.976 31.032 ;
  LAYER M3 ;
        RECT 19.008 28.524 19.04 31.032 ;
  LAYER M3 ;
        RECT 19.072 28.524 19.104 31.032 ;
  LAYER M3 ;
        RECT 19.136 28.524 19.168 31.032 ;
  LAYER M3 ;
        RECT 19.2 28.524 19.232 31.032 ;
  LAYER M3 ;
        RECT 19.264 28.524 19.296 31.032 ;
  LAYER M3 ;
        RECT 19.328 28.524 19.36 31.032 ;
  LAYER M3 ;
        RECT 19.392 28.524 19.424 31.032 ;
  LAYER M3 ;
        RECT 19.456 28.524 19.488 31.032 ;
  LAYER M3 ;
        RECT 19.52 28.524 19.552 31.032 ;
  LAYER M3 ;
        RECT 19.584 28.524 19.616 31.032 ;
  LAYER M3 ;
        RECT 19.648 28.524 19.68 31.032 ;
  LAYER M3 ;
        RECT 19.712 28.524 19.744 31.032 ;
  LAYER M3 ;
        RECT 19.776 28.524 19.808 31.032 ;
  LAYER M3 ;
        RECT 19.84 28.524 19.872 31.032 ;
  LAYER M3 ;
        RECT 19.904 28.524 19.936 31.032 ;
  LAYER M3 ;
        RECT 19.968 28.524 20 31.032 ;
  LAYER M3 ;
        RECT 20.032 28.524 20.064 31.032 ;
  LAYER M3 ;
        RECT 20.096 28.524 20.128 31.032 ;
  LAYER M3 ;
        RECT 20.16 28.524 20.192 31.032 ;
  LAYER M3 ;
        RECT 20.224 28.524 20.256 31.032 ;
  LAYER M3 ;
        RECT 20.288 28.524 20.32 31.032 ;
  LAYER M3 ;
        RECT 20.352 28.524 20.384 31.032 ;
  LAYER M3 ;
        RECT 20.416 28.524 20.448 31.032 ;
  LAYER M3 ;
        RECT 20.48 28.524 20.512 31.032 ;
  LAYER M3 ;
        RECT 20.544 28.524 20.576 31.032 ;
  LAYER M3 ;
        RECT 20.608 28.524 20.64 31.032 ;
  LAYER M3 ;
        RECT 20.672 28.524 20.704 31.032 ;
  LAYER M3 ;
        RECT 20.736 28.524 20.768 31.032 ;
  LAYER M3 ;
        RECT 20.8 28.524 20.832 31.032 ;
  LAYER M3 ;
        RECT 20.864 28.524 20.896 31.032 ;
  LAYER M3 ;
        RECT 20.928 28.524 20.96 31.032 ;
  LAYER M3 ;
        RECT 20.992 28.524 21.024 31.032 ;
  LAYER M3 ;
        RECT 21.056 28.524 21.088 31.032 ;
  LAYER M3 ;
        RECT 21.12 28.524 21.152 31.032 ;
  LAYER M3 ;
        RECT 21.184 28.524 21.216 31.032 ;
  LAYER M3 ;
        RECT 21.248 28.524 21.28 31.032 ;
  LAYER M3 ;
        RECT 21.344 28.524 21.376 31.032 ;
  LAYER M1 ;
        RECT 18.959 28.56 18.961 30.996 ;
  LAYER M1 ;
        RECT 19.039 28.56 19.041 30.996 ;
  LAYER M1 ;
        RECT 19.119 28.56 19.121 30.996 ;
  LAYER M1 ;
        RECT 19.199 28.56 19.201 30.996 ;
  LAYER M1 ;
        RECT 19.279 28.56 19.281 30.996 ;
  LAYER M1 ;
        RECT 19.359 28.56 19.361 30.996 ;
  LAYER M1 ;
        RECT 19.439 28.56 19.441 30.996 ;
  LAYER M1 ;
        RECT 19.519 28.56 19.521 30.996 ;
  LAYER M1 ;
        RECT 19.599 28.56 19.601 30.996 ;
  LAYER M1 ;
        RECT 19.679 28.56 19.681 30.996 ;
  LAYER M1 ;
        RECT 19.759 28.56 19.761 30.996 ;
  LAYER M1 ;
        RECT 19.839 28.56 19.841 30.996 ;
  LAYER M1 ;
        RECT 19.919 28.56 19.921 30.996 ;
  LAYER M1 ;
        RECT 19.999 28.56 20.001 30.996 ;
  LAYER M1 ;
        RECT 20.079 28.56 20.081 30.996 ;
  LAYER M1 ;
        RECT 20.159 28.56 20.161 30.996 ;
  LAYER M1 ;
        RECT 20.239 28.56 20.241 30.996 ;
  LAYER M1 ;
        RECT 20.319 28.56 20.321 30.996 ;
  LAYER M1 ;
        RECT 20.399 28.56 20.401 30.996 ;
  LAYER M1 ;
        RECT 20.479 28.56 20.481 30.996 ;
  LAYER M1 ;
        RECT 20.559 28.56 20.561 30.996 ;
  LAYER M1 ;
        RECT 20.639 28.56 20.641 30.996 ;
  LAYER M1 ;
        RECT 20.719 28.56 20.721 30.996 ;
  LAYER M1 ;
        RECT 20.799 28.56 20.801 30.996 ;
  LAYER M1 ;
        RECT 20.879 28.56 20.881 30.996 ;
  LAYER M1 ;
        RECT 20.959 28.56 20.961 30.996 ;
  LAYER M1 ;
        RECT 21.039 28.56 21.041 30.996 ;
  LAYER M1 ;
        RECT 21.119 28.56 21.121 30.996 ;
  LAYER M1 ;
        RECT 21.199 28.56 21.201 30.996 ;
  LAYER M1 ;
        RECT 21.279 28.56 21.281 30.996 ;
  LAYER M2 ;
        RECT 18.96 30.995 21.36 30.997 ;
  LAYER M2 ;
        RECT 18.96 30.911 21.36 30.913 ;
  LAYER M2 ;
        RECT 18.96 30.827 21.36 30.829 ;
  LAYER M2 ;
        RECT 18.96 30.743 21.36 30.745 ;
  LAYER M2 ;
        RECT 18.96 30.659 21.36 30.661 ;
  LAYER M2 ;
        RECT 18.96 30.575 21.36 30.577 ;
  LAYER M2 ;
        RECT 18.96 30.491 21.36 30.493 ;
  LAYER M2 ;
        RECT 18.96 30.407 21.36 30.409 ;
  LAYER M2 ;
        RECT 18.96 30.323 21.36 30.325 ;
  LAYER M2 ;
        RECT 18.96 30.239 21.36 30.241 ;
  LAYER M2 ;
        RECT 18.96 30.155 21.36 30.157 ;
  LAYER M2 ;
        RECT 18.96 30.071 21.36 30.073 ;
  LAYER M2 ;
        RECT 18.96 29.9875 21.36 29.9895 ;
  LAYER M2 ;
        RECT 18.96 29.903 21.36 29.905 ;
  LAYER M2 ;
        RECT 18.96 29.819 21.36 29.821 ;
  LAYER M2 ;
        RECT 18.96 29.735 21.36 29.737 ;
  LAYER M2 ;
        RECT 18.96 29.651 21.36 29.653 ;
  LAYER M2 ;
        RECT 18.96 29.567 21.36 29.569 ;
  LAYER M2 ;
        RECT 18.96 29.483 21.36 29.485 ;
  LAYER M2 ;
        RECT 18.96 29.399 21.36 29.401 ;
  LAYER M2 ;
        RECT 18.96 29.315 21.36 29.317 ;
  LAYER M2 ;
        RECT 18.96 29.231 21.36 29.233 ;
  LAYER M2 ;
        RECT 18.96 29.147 21.36 29.149 ;
  LAYER M2 ;
        RECT 18.96 29.063 21.36 29.065 ;
  LAYER M2 ;
        RECT 18.96 28.979 21.36 28.981 ;
  LAYER M2 ;
        RECT 18.96 28.895 21.36 28.897 ;
  LAYER M2 ;
        RECT 18.96 28.811 21.36 28.813 ;
  LAYER M2 ;
        RECT 18.96 28.727 21.36 28.729 ;
  LAYER M2 ;
        RECT 18.96 28.643 21.36 28.645 ;
  LAYER M1 ;
        RECT 18.944 25.584 18.976 28.092 ;
  LAYER M1 ;
        RECT 19.008 25.584 19.04 28.092 ;
  LAYER M1 ;
        RECT 19.072 25.584 19.104 28.092 ;
  LAYER M1 ;
        RECT 19.136 25.584 19.168 28.092 ;
  LAYER M1 ;
        RECT 19.2 25.584 19.232 28.092 ;
  LAYER M1 ;
        RECT 19.264 25.584 19.296 28.092 ;
  LAYER M1 ;
        RECT 19.328 25.584 19.36 28.092 ;
  LAYER M1 ;
        RECT 19.392 25.584 19.424 28.092 ;
  LAYER M1 ;
        RECT 19.456 25.584 19.488 28.092 ;
  LAYER M1 ;
        RECT 19.52 25.584 19.552 28.092 ;
  LAYER M1 ;
        RECT 19.584 25.584 19.616 28.092 ;
  LAYER M1 ;
        RECT 19.648 25.584 19.68 28.092 ;
  LAYER M1 ;
        RECT 19.712 25.584 19.744 28.092 ;
  LAYER M1 ;
        RECT 19.776 25.584 19.808 28.092 ;
  LAYER M1 ;
        RECT 19.84 25.584 19.872 28.092 ;
  LAYER M1 ;
        RECT 19.904 25.584 19.936 28.092 ;
  LAYER M1 ;
        RECT 19.968 25.584 20 28.092 ;
  LAYER M1 ;
        RECT 20.032 25.584 20.064 28.092 ;
  LAYER M1 ;
        RECT 20.096 25.584 20.128 28.092 ;
  LAYER M1 ;
        RECT 20.16 25.584 20.192 28.092 ;
  LAYER M1 ;
        RECT 20.224 25.584 20.256 28.092 ;
  LAYER M1 ;
        RECT 20.288 25.584 20.32 28.092 ;
  LAYER M1 ;
        RECT 20.352 25.584 20.384 28.092 ;
  LAYER M1 ;
        RECT 20.416 25.584 20.448 28.092 ;
  LAYER M1 ;
        RECT 20.48 25.584 20.512 28.092 ;
  LAYER M1 ;
        RECT 20.544 25.584 20.576 28.092 ;
  LAYER M1 ;
        RECT 20.608 25.584 20.64 28.092 ;
  LAYER M1 ;
        RECT 20.672 25.584 20.704 28.092 ;
  LAYER M1 ;
        RECT 20.736 25.584 20.768 28.092 ;
  LAYER M1 ;
        RECT 20.8 25.584 20.832 28.092 ;
  LAYER M1 ;
        RECT 20.864 25.584 20.896 28.092 ;
  LAYER M1 ;
        RECT 20.928 25.584 20.96 28.092 ;
  LAYER M1 ;
        RECT 20.992 25.584 21.024 28.092 ;
  LAYER M1 ;
        RECT 21.056 25.584 21.088 28.092 ;
  LAYER M1 ;
        RECT 21.12 25.584 21.152 28.092 ;
  LAYER M1 ;
        RECT 21.184 25.584 21.216 28.092 ;
  LAYER M1 ;
        RECT 21.248 25.584 21.28 28.092 ;
  LAYER M2 ;
        RECT 18.924 27.976 21.396 28.008 ;
  LAYER M2 ;
        RECT 18.924 27.912 21.396 27.944 ;
  LAYER M2 ;
        RECT 18.924 27.848 21.396 27.88 ;
  LAYER M2 ;
        RECT 18.924 27.784 21.396 27.816 ;
  LAYER M2 ;
        RECT 18.924 27.72 21.396 27.752 ;
  LAYER M2 ;
        RECT 18.924 27.656 21.396 27.688 ;
  LAYER M2 ;
        RECT 18.924 27.592 21.396 27.624 ;
  LAYER M2 ;
        RECT 18.924 27.528 21.396 27.56 ;
  LAYER M2 ;
        RECT 18.924 27.464 21.396 27.496 ;
  LAYER M2 ;
        RECT 18.924 27.4 21.396 27.432 ;
  LAYER M2 ;
        RECT 18.924 27.336 21.396 27.368 ;
  LAYER M2 ;
        RECT 18.924 27.272 21.396 27.304 ;
  LAYER M2 ;
        RECT 18.924 27.208 21.396 27.24 ;
  LAYER M2 ;
        RECT 18.924 27.144 21.396 27.176 ;
  LAYER M2 ;
        RECT 18.924 27.08 21.396 27.112 ;
  LAYER M2 ;
        RECT 18.924 27.016 21.396 27.048 ;
  LAYER M2 ;
        RECT 18.924 26.952 21.396 26.984 ;
  LAYER M2 ;
        RECT 18.924 26.888 21.396 26.92 ;
  LAYER M2 ;
        RECT 18.924 26.824 21.396 26.856 ;
  LAYER M2 ;
        RECT 18.924 26.76 21.396 26.792 ;
  LAYER M2 ;
        RECT 18.924 26.696 21.396 26.728 ;
  LAYER M2 ;
        RECT 18.924 26.632 21.396 26.664 ;
  LAYER M2 ;
        RECT 18.924 26.568 21.396 26.6 ;
  LAYER M2 ;
        RECT 18.924 26.504 21.396 26.536 ;
  LAYER M2 ;
        RECT 18.924 26.44 21.396 26.472 ;
  LAYER M2 ;
        RECT 18.924 26.376 21.396 26.408 ;
  LAYER M2 ;
        RECT 18.924 26.312 21.396 26.344 ;
  LAYER M2 ;
        RECT 18.924 26.248 21.396 26.28 ;
  LAYER M2 ;
        RECT 18.924 26.184 21.396 26.216 ;
  LAYER M2 ;
        RECT 18.924 26.12 21.396 26.152 ;
  LAYER M2 ;
        RECT 18.924 26.056 21.396 26.088 ;
  LAYER M2 ;
        RECT 18.924 25.992 21.396 26.024 ;
  LAYER M2 ;
        RECT 18.924 25.928 21.396 25.96 ;
  LAYER M2 ;
        RECT 18.924 25.864 21.396 25.896 ;
  LAYER M2 ;
        RECT 18.924 25.8 21.396 25.832 ;
  LAYER M2 ;
        RECT 18.924 25.736 21.396 25.768 ;
  LAYER M3 ;
        RECT 18.944 25.584 18.976 28.092 ;
  LAYER M3 ;
        RECT 19.008 25.584 19.04 28.092 ;
  LAYER M3 ;
        RECT 19.072 25.584 19.104 28.092 ;
  LAYER M3 ;
        RECT 19.136 25.584 19.168 28.092 ;
  LAYER M3 ;
        RECT 19.2 25.584 19.232 28.092 ;
  LAYER M3 ;
        RECT 19.264 25.584 19.296 28.092 ;
  LAYER M3 ;
        RECT 19.328 25.584 19.36 28.092 ;
  LAYER M3 ;
        RECT 19.392 25.584 19.424 28.092 ;
  LAYER M3 ;
        RECT 19.456 25.584 19.488 28.092 ;
  LAYER M3 ;
        RECT 19.52 25.584 19.552 28.092 ;
  LAYER M3 ;
        RECT 19.584 25.584 19.616 28.092 ;
  LAYER M3 ;
        RECT 19.648 25.584 19.68 28.092 ;
  LAYER M3 ;
        RECT 19.712 25.584 19.744 28.092 ;
  LAYER M3 ;
        RECT 19.776 25.584 19.808 28.092 ;
  LAYER M3 ;
        RECT 19.84 25.584 19.872 28.092 ;
  LAYER M3 ;
        RECT 19.904 25.584 19.936 28.092 ;
  LAYER M3 ;
        RECT 19.968 25.584 20 28.092 ;
  LAYER M3 ;
        RECT 20.032 25.584 20.064 28.092 ;
  LAYER M3 ;
        RECT 20.096 25.584 20.128 28.092 ;
  LAYER M3 ;
        RECT 20.16 25.584 20.192 28.092 ;
  LAYER M3 ;
        RECT 20.224 25.584 20.256 28.092 ;
  LAYER M3 ;
        RECT 20.288 25.584 20.32 28.092 ;
  LAYER M3 ;
        RECT 20.352 25.584 20.384 28.092 ;
  LAYER M3 ;
        RECT 20.416 25.584 20.448 28.092 ;
  LAYER M3 ;
        RECT 20.48 25.584 20.512 28.092 ;
  LAYER M3 ;
        RECT 20.544 25.584 20.576 28.092 ;
  LAYER M3 ;
        RECT 20.608 25.584 20.64 28.092 ;
  LAYER M3 ;
        RECT 20.672 25.584 20.704 28.092 ;
  LAYER M3 ;
        RECT 20.736 25.584 20.768 28.092 ;
  LAYER M3 ;
        RECT 20.8 25.584 20.832 28.092 ;
  LAYER M3 ;
        RECT 20.864 25.584 20.896 28.092 ;
  LAYER M3 ;
        RECT 20.928 25.584 20.96 28.092 ;
  LAYER M3 ;
        RECT 20.992 25.584 21.024 28.092 ;
  LAYER M3 ;
        RECT 21.056 25.584 21.088 28.092 ;
  LAYER M3 ;
        RECT 21.12 25.584 21.152 28.092 ;
  LAYER M3 ;
        RECT 21.184 25.584 21.216 28.092 ;
  LAYER M3 ;
        RECT 21.248 25.584 21.28 28.092 ;
  LAYER M3 ;
        RECT 21.344 25.584 21.376 28.092 ;
  LAYER M1 ;
        RECT 18.959 25.62 18.961 28.056 ;
  LAYER M1 ;
        RECT 19.039 25.62 19.041 28.056 ;
  LAYER M1 ;
        RECT 19.119 25.62 19.121 28.056 ;
  LAYER M1 ;
        RECT 19.199 25.62 19.201 28.056 ;
  LAYER M1 ;
        RECT 19.279 25.62 19.281 28.056 ;
  LAYER M1 ;
        RECT 19.359 25.62 19.361 28.056 ;
  LAYER M1 ;
        RECT 19.439 25.62 19.441 28.056 ;
  LAYER M1 ;
        RECT 19.519 25.62 19.521 28.056 ;
  LAYER M1 ;
        RECT 19.599 25.62 19.601 28.056 ;
  LAYER M1 ;
        RECT 19.679 25.62 19.681 28.056 ;
  LAYER M1 ;
        RECT 19.759 25.62 19.761 28.056 ;
  LAYER M1 ;
        RECT 19.839 25.62 19.841 28.056 ;
  LAYER M1 ;
        RECT 19.919 25.62 19.921 28.056 ;
  LAYER M1 ;
        RECT 19.999 25.62 20.001 28.056 ;
  LAYER M1 ;
        RECT 20.079 25.62 20.081 28.056 ;
  LAYER M1 ;
        RECT 20.159 25.62 20.161 28.056 ;
  LAYER M1 ;
        RECT 20.239 25.62 20.241 28.056 ;
  LAYER M1 ;
        RECT 20.319 25.62 20.321 28.056 ;
  LAYER M1 ;
        RECT 20.399 25.62 20.401 28.056 ;
  LAYER M1 ;
        RECT 20.479 25.62 20.481 28.056 ;
  LAYER M1 ;
        RECT 20.559 25.62 20.561 28.056 ;
  LAYER M1 ;
        RECT 20.639 25.62 20.641 28.056 ;
  LAYER M1 ;
        RECT 20.719 25.62 20.721 28.056 ;
  LAYER M1 ;
        RECT 20.799 25.62 20.801 28.056 ;
  LAYER M1 ;
        RECT 20.879 25.62 20.881 28.056 ;
  LAYER M1 ;
        RECT 20.959 25.62 20.961 28.056 ;
  LAYER M1 ;
        RECT 21.039 25.62 21.041 28.056 ;
  LAYER M1 ;
        RECT 21.119 25.62 21.121 28.056 ;
  LAYER M1 ;
        RECT 21.199 25.62 21.201 28.056 ;
  LAYER M1 ;
        RECT 21.279 25.62 21.281 28.056 ;
  LAYER M2 ;
        RECT 18.96 28.055 21.36 28.057 ;
  LAYER M2 ;
        RECT 18.96 27.971 21.36 27.973 ;
  LAYER M2 ;
        RECT 18.96 27.887 21.36 27.889 ;
  LAYER M2 ;
        RECT 18.96 27.803 21.36 27.805 ;
  LAYER M2 ;
        RECT 18.96 27.719 21.36 27.721 ;
  LAYER M2 ;
        RECT 18.96 27.635 21.36 27.637 ;
  LAYER M2 ;
        RECT 18.96 27.551 21.36 27.553 ;
  LAYER M2 ;
        RECT 18.96 27.467 21.36 27.469 ;
  LAYER M2 ;
        RECT 18.96 27.383 21.36 27.385 ;
  LAYER M2 ;
        RECT 18.96 27.299 21.36 27.301 ;
  LAYER M2 ;
        RECT 18.96 27.215 21.36 27.217 ;
  LAYER M2 ;
        RECT 18.96 27.131 21.36 27.133 ;
  LAYER M2 ;
        RECT 18.96 27.0475 21.36 27.0495 ;
  LAYER M2 ;
        RECT 18.96 26.963 21.36 26.965 ;
  LAYER M2 ;
        RECT 18.96 26.879 21.36 26.881 ;
  LAYER M2 ;
        RECT 18.96 26.795 21.36 26.797 ;
  LAYER M2 ;
        RECT 18.96 26.711 21.36 26.713 ;
  LAYER M2 ;
        RECT 18.96 26.627 21.36 26.629 ;
  LAYER M2 ;
        RECT 18.96 26.543 21.36 26.545 ;
  LAYER M2 ;
        RECT 18.96 26.459 21.36 26.461 ;
  LAYER M2 ;
        RECT 18.96 26.375 21.36 26.377 ;
  LAYER M2 ;
        RECT 18.96 26.291 21.36 26.293 ;
  LAYER M2 ;
        RECT 18.96 26.207 21.36 26.209 ;
  LAYER M2 ;
        RECT 18.96 26.123 21.36 26.125 ;
  LAYER M2 ;
        RECT 18.96 26.039 21.36 26.041 ;
  LAYER M2 ;
        RECT 18.96 25.955 21.36 25.957 ;
  LAYER M2 ;
        RECT 18.96 25.871 21.36 25.873 ;
  LAYER M2 ;
        RECT 18.96 25.787 21.36 25.789 ;
  LAYER M2 ;
        RECT 18.96 25.703 21.36 25.705 ;
  LAYER M1 ;
        RECT 18.944 22.644 18.976 25.152 ;
  LAYER M1 ;
        RECT 19.008 22.644 19.04 25.152 ;
  LAYER M1 ;
        RECT 19.072 22.644 19.104 25.152 ;
  LAYER M1 ;
        RECT 19.136 22.644 19.168 25.152 ;
  LAYER M1 ;
        RECT 19.2 22.644 19.232 25.152 ;
  LAYER M1 ;
        RECT 19.264 22.644 19.296 25.152 ;
  LAYER M1 ;
        RECT 19.328 22.644 19.36 25.152 ;
  LAYER M1 ;
        RECT 19.392 22.644 19.424 25.152 ;
  LAYER M1 ;
        RECT 19.456 22.644 19.488 25.152 ;
  LAYER M1 ;
        RECT 19.52 22.644 19.552 25.152 ;
  LAYER M1 ;
        RECT 19.584 22.644 19.616 25.152 ;
  LAYER M1 ;
        RECT 19.648 22.644 19.68 25.152 ;
  LAYER M1 ;
        RECT 19.712 22.644 19.744 25.152 ;
  LAYER M1 ;
        RECT 19.776 22.644 19.808 25.152 ;
  LAYER M1 ;
        RECT 19.84 22.644 19.872 25.152 ;
  LAYER M1 ;
        RECT 19.904 22.644 19.936 25.152 ;
  LAYER M1 ;
        RECT 19.968 22.644 20 25.152 ;
  LAYER M1 ;
        RECT 20.032 22.644 20.064 25.152 ;
  LAYER M1 ;
        RECT 20.096 22.644 20.128 25.152 ;
  LAYER M1 ;
        RECT 20.16 22.644 20.192 25.152 ;
  LAYER M1 ;
        RECT 20.224 22.644 20.256 25.152 ;
  LAYER M1 ;
        RECT 20.288 22.644 20.32 25.152 ;
  LAYER M1 ;
        RECT 20.352 22.644 20.384 25.152 ;
  LAYER M1 ;
        RECT 20.416 22.644 20.448 25.152 ;
  LAYER M1 ;
        RECT 20.48 22.644 20.512 25.152 ;
  LAYER M1 ;
        RECT 20.544 22.644 20.576 25.152 ;
  LAYER M1 ;
        RECT 20.608 22.644 20.64 25.152 ;
  LAYER M1 ;
        RECT 20.672 22.644 20.704 25.152 ;
  LAYER M1 ;
        RECT 20.736 22.644 20.768 25.152 ;
  LAYER M1 ;
        RECT 20.8 22.644 20.832 25.152 ;
  LAYER M1 ;
        RECT 20.864 22.644 20.896 25.152 ;
  LAYER M1 ;
        RECT 20.928 22.644 20.96 25.152 ;
  LAYER M1 ;
        RECT 20.992 22.644 21.024 25.152 ;
  LAYER M1 ;
        RECT 21.056 22.644 21.088 25.152 ;
  LAYER M1 ;
        RECT 21.12 22.644 21.152 25.152 ;
  LAYER M1 ;
        RECT 21.184 22.644 21.216 25.152 ;
  LAYER M1 ;
        RECT 21.248 22.644 21.28 25.152 ;
  LAYER M2 ;
        RECT 18.924 25.036 21.396 25.068 ;
  LAYER M2 ;
        RECT 18.924 24.972 21.396 25.004 ;
  LAYER M2 ;
        RECT 18.924 24.908 21.396 24.94 ;
  LAYER M2 ;
        RECT 18.924 24.844 21.396 24.876 ;
  LAYER M2 ;
        RECT 18.924 24.78 21.396 24.812 ;
  LAYER M2 ;
        RECT 18.924 24.716 21.396 24.748 ;
  LAYER M2 ;
        RECT 18.924 24.652 21.396 24.684 ;
  LAYER M2 ;
        RECT 18.924 24.588 21.396 24.62 ;
  LAYER M2 ;
        RECT 18.924 24.524 21.396 24.556 ;
  LAYER M2 ;
        RECT 18.924 24.46 21.396 24.492 ;
  LAYER M2 ;
        RECT 18.924 24.396 21.396 24.428 ;
  LAYER M2 ;
        RECT 18.924 24.332 21.396 24.364 ;
  LAYER M2 ;
        RECT 18.924 24.268 21.396 24.3 ;
  LAYER M2 ;
        RECT 18.924 24.204 21.396 24.236 ;
  LAYER M2 ;
        RECT 18.924 24.14 21.396 24.172 ;
  LAYER M2 ;
        RECT 18.924 24.076 21.396 24.108 ;
  LAYER M2 ;
        RECT 18.924 24.012 21.396 24.044 ;
  LAYER M2 ;
        RECT 18.924 23.948 21.396 23.98 ;
  LAYER M2 ;
        RECT 18.924 23.884 21.396 23.916 ;
  LAYER M2 ;
        RECT 18.924 23.82 21.396 23.852 ;
  LAYER M2 ;
        RECT 18.924 23.756 21.396 23.788 ;
  LAYER M2 ;
        RECT 18.924 23.692 21.396 23.724 ;
  LAYER M2 ;
        RECT 18.924 23.628 21.396 23.66 ;
  LAYER M2 ;
        RECT 18.924 23.564 21.396 23.596 ;
  LAYER M2 ;
        RECT 18.924 23.5 21.396 23.532 ;
  LAYER M2 ;
        RECT 18.924 23.436 21.396 23.468 ;
  LAYER M2 ;
        RECT 18.924 23.372 21.396 23.404 ;
  LAYER M2 ;
        RECT 18.924 23.308 21.396 23.34 ;
  LAYER M2 ;
        RECT 18.924 23.244 21.396 23.276 ;
  LAYER M2 ;
        RECT 18.924 23.18 21.396 23.212 ;
  LAYER M2 ;
        RECT 18.924 23.116 21.396 23.148 ;
  LAYER M2 ;
        RECT 18.924 23.052 21.396 23.084 ;
  LAYER M2 ;
        RECT 18.924 22.988 21.396 23.02 ;
  LAYER M2 ;
        RECT 18.924 22.924 21.396 22.956 ;
  LAYER M2 ;
        RECT 18.924 22.86 21.396 22.892 ;
  LAYER M2 ;
        RECT 18.924 22.796 21.396 22.828 ;
  LAYER M3 ;
        RECT 18.944 22.644 18.976 25.152 ;
  LAYER M3 ;
        RECT 19.008 22.644 19.04 25.152 ;
  LAYER M3 ;
        RECT 19.072 22.644 19.104 25.152 ;
  LAYER M3 ;
        RECT 19.136 22.644 19.168 25.152 ;
  LAYER M3 ;
        RECT 19.2 22.644 19.232 25.152 ;
  LAYER M3 ;
        RECT 19.264 22.644 19.296 25.152 ;
  LAYER M3 ;
        RECT 19.328 22.644 19.36 25.152 ;
  LAYER M3 ;
        RECT 19.392 22.644 19.424 25.152 ;
  LAYER M3 ;
        RECT 19.456 22.644 19.488 25.152 ;
  LAYER M3 ;
        RECT 19.52 22.644 19.552 25.152 ;
  LAYER M3 ;
        RECT 19.584 22.644 19.616 25.152 ;
  LAYER M3 ;
        RECT 19.648 22.644 19.68 25.152 ;
  LAYER M3 ;
        RECT 19.712 22.644 19.744 25.152 ;
  LAYER M3 ;
        RECT 19.776 22.644 19.808 25.152 ;
  LAYER M3 ;
        RECT 19.84 22.644 19.872 25.152 ;
  LAYER M3 ;
        RECT 19.904 22.644 19.936 25.152 ;
  LAYER M3 ;
        RECT 19.968 22.644 20 25.152 ;
  LAYER M3 ;
        RECT 20.032 22.644 20.064 25.152 ;
  LAYER M3 ;
        RECT 20.096 22.644 20.128 25.152 ;
  LAYER M3 ;
        RECT 20.16 22.644 20.192 25.152 ;
  LAYER M3 ;
        RECT 20.224 22.644 20.256 25.152 ;
  LAYER M3 ;
        RECT 20.288 22.644 20.32 25.152 ;
  LAYER M3 ;
        RECT 20.352 22.644 20.384 25.152 ;
  LAYER M3 ;
        RECT 20.416 22.644 20.448 25.152 ;
  LAYER M3 ;
        RECT 20.48 22.644 20.512 25.152 ;
  LAYER M3 ;
        RECT 20.544 22.644 20.576 25.152 ;
  LAYER M3 ;
        RECT 20.608 22.644 20.64 25.152 ;
  LAYER M3 ;
        RECT 20.672 22.644 20.704 25.152 ;
  LAYER M3 ;
        RECT 20.736 22.644 20.768 25.152 ;
  LAYER M3 ;
        RECT 20.8 22.644 20.832 25.152 ;
  LAYER M3 ;
        RECT 20.864 22.644 20.896 25.152 ;
  LAYER M3 ;
        RECT 20.928 22.644 20.96 25.152 ;
  LAYER M3 ;
        RECT 20.992 22.644 21.024 25.152 ;
  LAYER M3 ;
        RECT 21.056 22.644 21.088 25.152 ;
  LAYER M3 ;
        RECT 21.12 22.644 21.152 25.152 ;
  LAYER M3 ;
        RECT 21.184 22.644 21.216 25.152 ;
  LAYER M3 ;
        RECT 21.248 22.644 21.28 25.152 ;
  LAYER M3 ;
        RECT 21.344 22.644 21.376 25.152 ;
  LAYER M1 ;
        RECT 18.959 22.68 18.961 25.116 ;
  LAYER M1 ;
        RECT 19.039 22.68 19.041 25.116 ;
  LAYER M1 ;
        RECT 19.119 22.68 19.121 25.116 ;
  LAYER M1 ;
        RECT 19.199 22.68 19.201 25.116 ;
  LAYER M1 ;
        RECT 19.279 22.68 19.281 25.116 ;
  LAYER M1 ;
        RECT 19.359 22.68 19.361 25.116 ;
  LAYER M1 ;
        RECT 19.439 22.68 19.441 25.116 ;
  LAYER M1 ;
        RECT 19.519 22.68 19.521 25.116 ;
  LAYER M1 ;
        RECT 19.599 22.68 19.601 25.116 ;
  LAYER M1 ;
        RECT 19.679 22.68 19.681 25.116 ;
  LAYER M1 ;
        RECT 19.759 22.68 19.761 25.116 ;
  LAYER M1 ;
        RECT 19.839 22.68 19.841 25.116 ;
  LAYER M1 ;
        RECT 19.919 22.68 19.921 25.116 ;
  LAYER M1 ;
        RECT 19.999 22.68 20.001 25.116 ;
  LAYER M1 ;
        RECT 20.079 22.68 20.081 25.116 ;
  LAYER M1 ;
        RECT 20.159 22.68 20.161 25.116 ;
  LAYER M1 ;
        RECT 20.239 22.68 20.241 25.116 ;
  LAYER M1 ;
        RECT 20.319 22.68 20.321 25.116 ;
  LAYER M1 ;
        RECT 20.399 22.68 20.401 25.116 ;
  LAYER M1 ;
        RECT 20.479 22.68 20.481 25.116 ;
  LAYER M1 ;
        RECT 20.559 22.68 20.561 25.116 ;
  LAYER M1 ;
        RECT 20.639 22.68 20.641 25.116 ;
  LAYER M1 ;
        RECT 20.719 22.68 20.721 25.116 ;
  LAYER M1 ;
        RECT 20.799 22.68 20.801 25.116 ;
  LAYER M1 ;
        RECT 20.879 22.68 20.881 25.116 ;
  LAYER M1 ;
        RECT 20.959 22.68 20.961 25.116 ;
  LAYER M1 ;
        RECT 21.039 22.68 21.041 25.116 ;
  LAYER M1 ;
        RECT 21.119 22.68 21.121 25.116 ;
  LAYER M1 ;
        RECT 21.199 22.68 21.201 25.116 ;
  LAYER M1 ;
        RECT 21.279 22.68 21.281 25.116 ;
  LAYER M2 ;
        RECT 18.96 25.115 21.36 25.117 ;
  LAYER M2 ;
        RECT 18.96 25.031 21.36 25.033 ;
  LAYER M2 ;
        RECT 18.96 24.947 21.36 24.949 ;
  LAYER M2 ;
        RECT 18.96 24.863 21.36 24.865 ;
  LAYER M2 ;
        RECT 18.96 24.779 21.36 24.781 ;
  LAYER M2 ;
        RECT 18.96 24.695 21.36 24.697 ;
  LAYER M2 ;
        RECT 18.96 24.611 21.36 24.613 ;
  LAYER M2 ;
        RECT 18.96 24.527 21.36 24.529 ;
  LAYER M2 ;
        RECT 18.96 24.443 21.36 24.445 ;
  LAYER M2 ;
        RECT 18.96 24.359 21.36 24.361 ;
  LAYER M2 ;
        RECT 18.96 24.275 21.36 24.277 ;
  LAYER M2 ;
        RECT 18.96 24.191 21.36 24.193 ;
  LAYER M2 ;
        RECT 18.96 24.1075 21.36 24.1095 ;
  LAYER M2 ;
        RECT 18.96 24.023 21.36 24.025 ;
  LAYER M2 ;
        RECT 18.96 23.939 21.36 23.941 ;
  LAYER M2 ;
        RECT 18.96 23.855 21.36 23.857 ;
  LAYER M2 ;
        RECT 18.96 23.771 21.36 23.773 ;
  LAYER M2 ;
        RECT 18.96 23.687 21.36 23.689 ;
  LAYER M2 ;
        RECT 18.96 23.603 21.36 23.605 ;
  LAYER M2 ;
        RECT 18.96 23.519 21.36 23.521 ;
  LAYER M2 ;
        RECT 18.96 23.435 21.36 23.437 ;
  LAYER M2 ;
        RECT 18.96 23.351 21.36 23.353 ;
  LAYER M2 ;
        RECT 18.96 23.267 21.36 23.269 ;
  LAYER M2 ;
        RECT 18.96 23.183 21.36 23.185 ;
  LAYER M2 ;
        RECT 18.96 23.099 21.36 23.101 ;
  LAYER M2 ;
        RECT 18.96 23.015 21.36 23.017 ;
  LAYER M2 ;
        RECT 18.96 22.931 21.36 22.933 ;
  LAYER M2 ;
        RECT 18.96 22.847 21.36 22.849 ;
  LAYER M2 ;
        RECT 18.96 22.763 21.36 22.765 ;
  LAYER M1 ;
        RECT 18.944 19.704 18.976 22.212 ;
  LAYER M1 ;
        RECT 19.008 19.704 19.04 22.212 ;
  LAYER M1 ;
        RECT 19.072 19.704 19.104 22.212 ;
  LAYER M1 ;
        RECT 19.136 19.704 19.168 22.212 ;
  LAYER M1 ;
        RECT 19.2 19.704 19.232 22.212 ;
  LAYER M1 ;
        RECT 19.264 19.704 19.296 22.212 ;
  LAYER M1 ;
        RECT 19.328 19.704 19.36 22.212 ;
  LAYER M1 ;
        RECT 19.392 19.704 19.424 22.212 ;
  LAYER M1 ;
        RECT 19.456 19.704 19.488 22.212 ;
  LAYER M1 ;
        RECT 19.52 19.704 19.552 22.212 ;
  LAYER M1 ;
        RECT 19.584 19.704 19.616 22.212 ;
  LAYER M1 ;
        RECT 19.648 19.704 19.68 22.212 ;
  LAYER M1 ;
        RECT 19.712 19.704 19.744 22.212 ;
  LAYER M1 ;
        RECT 19.776 19.704 19.808 22.212 ;
  LAYER M1 ;
        RECT 19.84 19.704 19.872 22.212 ;
  LAYER M1 ;
        RECT 19.904 19.704 19.936 22.212 ;
  LAYER M1 ;
        RECT 19.968 19.704 20 22.212 ;
  LAYER M1 ;
        RECT 20.032 19.704 20.064 22.212 ;
  LAYER M1 ;
        RECT 20.096 19.704 20.128 22.212 ;
  LAYER M1 ;
        RECT 20.16 19.704 20.192 22.212 ;
  LAYER M1 ;
        RECT 20.224 19.704 20.256 22.212 ;
  LAYER M1 ;
        RECT 20.288 19.704 20.32 22.212 ;
  LAYER M1 ;
        RECT 20.352 19.704 20.384 22.212 ;
  LAYER M1 ;
        RECT 20.416 19.704 20.448 22.212 ;
  LAYER M1 ;
        RECT 20.48 19.704 20.512 22.212 ;
  LAYER M1 ;
        RECT 20.544 19.704 20.576 22.212 ;
  LAYER M1 ;
        RECT 20.608 19.704 20.64 22.212 ;
  LAYER M1 ;
        RECT 20.672 19.704 20.704 22.212 ;
  LAYER M1 ;
        RECT 20.736 19.704 20.768 22.212 ;
  LAYER M1 ;
        RECT 20.8 19.704 20.832 22.212 ;
  LAYER M1 ;
        RECT 20.864 19.704 20.896 22.212 ;
  LAYER M1 ;
        RECT 20.928 19.704 20.96 22.212 ;
  LAYER M1 ;
        RECT 20.992 19.704 21.024 22.212 ;
  LAYER M1 ;
        RECT 21.056 19.704 21.088 22.212 ;
  LAYER M1 ;
        RECT 21.12 19.704 21.152 22.212 ;
  LAYER M1 ;
        RECT 21.184 19.704 21.216 22.212 ;
  LAYER M1 ;
        RECT 21.248 19.704 21.28 22.212 ;
  LAYER M2 ;
        RECT 18.924 22.096 21.396 22.128 ;
  LAYER M2 ;
        RECT 18.924 22.032 21.396 22.064 ;
  LAYER M2 ;
        RECT 18.924 21.968 21.396 22 ;
  LAYER M2 ;
        RECT 18.924 21.904 21.396 21.936 ;
  LAYER M2 ;
        RECT 18.924 21.84 21.396 21.872 ;
  LAYER M2 ;
        RECT 18.924 21.776 21.396 21.808 ;
  LAYER M2 ;
        RECT 18.924 21.712 21.396 21.744 ;
  LAYER M2 ;
        RECT 18.924 21.648 21.396 21.68 ;
  LAYER M2 ;
        RECT 18.924 21.584 21.396 21.616 ;
  LAYER M2 ;
        RECT 18.924 21.52 21.396 21.552 ;
  LAYER M2 ;
        RECT 18.924 21.456 21.396 21.488 ;
  LAYER M2 ;
        RECT 18.924 21.392 21.396 21.424 ;
  LAYER M2 ;
        RECT 18.924 21.328 21.396 21.36 ;
  LAYER M2 ;
        RECT 18.924 21.264 21.396 21.296 ;
  LAYER M2 ;
        RECT 18.924 21.2 21.396 21.232 ;
  LAYER M2 ;
        RECT 18.924 21.136 21.396 21.168 ;
  LAYER M2 ;
        RECT 18.924 21.072 21.396 21.104 ;
  LAYER M2 ;
        RECT 18.924 21.008 21.396 21.04 ;
  LAYER M2 ;
        RECT 18.924 20.944 21.396 20.976 ;
  LAYER M2 ;
        RECT 18.924 20.88 21.396 20.912 ;
  LAYER M2 ;
        RECT 18.924 20.816 21.396 20.848 ;
  LAYER M2 ;
        RECT 18.924 20.752 21.396 20.784 ;
  LAYER M2 ;
        RECT 18.924 20.688 21.396 20.72 ;
  LAYER M2 ;
        RECT 18.924 20.624 21.396 20.656 ;
  LAYER M2 ;
        RECT 18.924 20.56 21.396 20.592 ;
  LAYER M2 ;
        RECT 18.924 20.496 21.396 20.528 ;
  LAYER M2 ;
        RECT 18.924 20.432 21.396 20.464 ;
  LAYER M2 ;
        RECT 18.924 20.368 21.396 20.4 ;
  LAYER M2 ;
        RECT 18.924 20.304 21.396 20.336 ;
  LAYER M2 ;
        RECT 18.924 20.24 21.396 20.272 ;
  LAYER M2 ;
        RECT 18.924 20.176 21.396 20.208 ;
  LAYER M2 ;
        RECT 18.924 20.112 21.396 20.144 ;
  LAYER M2 ;
        RECT 18.924 20.048 21.396 20.08 ;
  LAYER M2 ;
        RECT 18.924 19.984 21.396 20.016 ;
  LAYER M2 ;
        RECT 18.924 19.92 21.396 19.952 ;
  LAYER M2 ;
        RECT 18.924 19.856 21.396 19.888 ;
  LAYER M3 ;
        RECT 18.944 19.704 18.976 22.212 ;
  LAYER M3 ;
        RECT 19.008 19.704 19.04 22.212 ;
  LAYER M3 ;
        RECT 19.072 19.704 19.104 22.212 ;
  LAYER M3 ;
        RECT 19.136 19.704 19.168 22.212 ;
  LAYER M3 ;
        RECT 19.2 19.704 19.232 22.212 ;
  LAYER M3 ;
        RECT 19.264 19.704 19.296 22.212 ;
  LAYER M3 ;
        RECT 19.328 19.704 19.36 22.212 ;
  LAYER M3 ;
        RECT 19.392 19.704 19.424 22.212 ;
  LAYER M3 ;
        RECT 19.456 19.704 19.488 22.212 ;
  LAYER M3 ;
        RECT 19.52 19.704 19.552 22.212 ;
  LAYER M3 ;
        RECT 19.584 19.704 19.616 22.212 ;
  LAYER M3 ;
        RECT 19.648 19.704 19.68 22.212 ;
  LAYER M3 ;
        RECT 19.712 19.704 19.744 22.212 ;
  LAYER M3 ;
        RECT 19.776 19.704 19.808 22.212 ;
  LAYER M3 ;
        RECT 19.84 19.704 19.872 22.212 ;
  LAYER M3 ;
        RECT 19.904 19.704 19.936 22.212 ;
  LAYER M3 ;
        RECT 19.968 19.704 20 22.212 ;
  LAYER M3 ;
        RECT 20.032 19.704 20.064 22.212 ;
  LAYER M3 ;
        RECT 20.096 19.704 20.128 22.212 ;
  LAYER M3 ;
        RECT 20.16 19.704 20.192 22.212 ;
  LAYER M3 ;
        RECT 20.224 19.704 20.256 22.212 ;
  LAYER M3 ;
        RECT 20.288 19.704 20.32 22.212 ;
  LAYER M3 ;
        RECT 20.352 19.704 20.384 22.212 ;
  LAYER M3 ;
        RECT 20.416 19.704 20.448 22.212 ;
  LAYER M3 ;
        RECT 20.48 19.704 20.512 22.212 ;
  LAYER M3 ;
        RECT 20.544 19.704 20.576 22.212 ;
  LAYER M3 ;
        RECT 20.608 19.704 20.64 22.212 ;
  LAYER M3 ;
        RECT 20.672 19.704 20.704 22.212 ;
  LAYER M3 ;
        RECT 20.736 19.704 20.768 22.212 ;
  LAYER M3 ;
        RECT 20.8 19.704 20.832 22.212 ;
  LAYER M3 ;
        RECT 20.864 19.704 20.896 22.212 ;
  LAYER M3 ;
        RECT 20.928 19.704 20.96 22.212 ;
  LAYER M3 ;
        RECT 20.992 19.704 21.024 22.212 ;
  LAYER M3 ;
        RECT 21.056 19.704 21.088 22.212 ;
  LAYER M3 ;
        RECT 21.12 19.704 21.152 22.212 ;
  LAYER M3 ;
        RECT 21.184 19.704 21.216 22.212 ;
  LAYER M3 ;
        RECT 21.248 19.704 21.28 22.212 ;
  LAYER M3 ;
        RECT 21.344 19.704 21.376 22.212 ;
  LAYER M1 ;
        RECT 18.959 19.74 18.961 22.176 ;
  LAYER M1 ;
        RECT 19.039 19.74 19.041 22.176 ;
  LAYER M1 ;
        RECT 19.119 19.74 19.121 22.176 ;
  LAYER M1 ;
        RECT 19.199 19.74 19.201 22.176 ;
  LAYER M1 ;
        RECT 19.279 19.74 19.281 22.176 ;
  LAYER M1 ;
        RECT 19.359 19.74 19.361 22.176 ;
  LAYER M1 ;
        RECT 19.439 19.74 19.441 22.176 ;
  LAYER M1 ;
        RECT 19.519 19.74 19.521 22.176 ;
  LAYER M1 ;
        RECT 19.599 19.74 19.601 22.176 ;
  LAYER M1 ;
        RECT 19.679 19.74 19.681 22.176 ;
  LAYER M1 ;
        RECT 19.759 19.74 19.761 22.176 ;
  LAYER M1 ;
        RECT 19.839 19.74 19.841 22.176 ;
  LAYER M1 ;
        RECT 19.919 19.74 19.921 22.176 ;
  LAYER M1 ;
        RECT 19.999 19.74 20.001 22.176 ;
  LAYER M1 ;
        RECT 20.079 19.74 20.081 22.176 ;
  LAYER M1 ;
        RECT 20.159 19.74 20.161 22.176 ;
  LAYER M1 ;
        RECT 20.239 19.74 20.241 22.176 ;
  LAYER M1 ;
        RECT 20.319 19.74 20.321 22.176 ;
  LAYER M1 ;
        RECT 20.399 19.74 20.401 22.176 ;
  LAYER M1 ;
        RECT 20.479 19.74 20.481 22.176 ;
  LAYER M1 ;
        RECT 20.559 19.74 20.561 22.176 ;
  LAYER M1 ;
        RECT 20.639 19.74 20.641 22.176 ;
  LAYER M1 ;
        RECT 20.719 19.74 20.721 22.176 ;
  LAYER M1 ;
        RECT 20.799 19.74 20.801 22.176 ;
  LAYER M1 ;
        RECT 20.879 19.74 20.881 22.176 ;
  LAYER M1 ;
        RECT 20.959 19.74 20.961 22.176 ;
  LAYER M1 ;
        RECT 21.039 19.74 21.041 22.176 ;
  LAYER M1 ;
        RECT 21.119 19.74 21.121 22.176 ;
  LAYER M1 ;
        RECT 21.199 19.74 21.201 22.176 ;
  LAYER M1 ;
        RECT 21.279 19.74 21.281 22.176 ;
  LAYER M2 ;
        RECT 18.96 22.175 21.36 22.177 ;
  LAYER M2 ;
        RECT 18.96 22.091 21.36 22.093 ;
  LAYER M2 ;
        RECT 18.96 22.007 21.36 22.009 ;
  LAYER M2 ;
        RECT 18.96 21.923 21.36 21.925 ;
  LAYER M2 ;
        RECT 18.96 21.839 21.36 21.841 ;
  LAYER M2 ;
        RECT 18.96 21.755 21.36 21.757 ;
  LAYER M2 ;
        RECT 18.96 21.671 21.36 21.673 ;
  LAYER M2 ;
        RECT 18.96 21.587 21.36 21.589 ;
  LAYER M2 ;
        RECT 18.96 21.503 21.36 21.505 ;
  LAYER M2 ;
        RECT 18.96 21.419 21.36 21.421 ;
  LAYER M2 ;
        RECT 18.96 21.335 21.36 21.337 ;
  LAYER M2 ;
        RECT 18.96 21.251 21.36 21.253 ;
  LAYER M2 ;
        RECT 18.96 21.1675 21.36 21.1695 ;
  LAYER M2 ;
        RECT 18.96 21.083 21.36 21.085 ;
  LAYER M2 ;
        RECT 18.96 20.999 21.36 21.001 ;
  LAYER M2 ;
        RECT 18.96 20.915 21.36 20.917 ;
  LAYER M2 ;
        RECT 18.96 20.831 21.36 20.833 ;
  LAYER M2 ;
        RECT 18.96 20.747 21.36 20.749 ;
  LAYER M2 ;
        RECT 18.96 20.663 21.36 20.665 ;
  LAYER M2 ;
        RECT 18.96 20.579 21.36 20.581 ;
  LAYER M2 ;
        RECT 18.96 20.495 21.36 20.497 ;
  LAYER M2 ;
        RECT 18.96 20.411 21.36 20.413 ;
  LAYER M2 ;
        RECT 18.96 20.327 21.36 20.329 ;
  LAYER M2 ;
        RECT 18.96 20.243 21.36 20.245 ;
  LAYER M2 ;
        RECT 18.96 20.159 21.36 20.161 ;
  LAYER M2 ;
        RECT 18.96 20.075 21.36 20.077 ;
  LAYER M2 ;
        RECT 18.96 19.991 21.36 19.993 ;
  LAYER M2 ;
        RECT 18.96 19.907 21.36 19.909 ;
  LAYER M2 ;
        RECT 18.96 19.823 21.36 19.825 ;
  LAYER M1 ;
        RECT 21.824 34.404 21.856 36.912 ;
  LAYER M1 ;
        RECT 21.888 34.404 21.92 36.912 ;
  LAYER M1 ;
        RECT 21.952 34.404 21.984 36.912 ;
  LAYER M1 ;
        RECT 22.016 34.404 22.048 36.912 ;
  LAYER M1 ;
        RECT 22.08 34.404 22.112 36.912 ;
  LAYER M1 ;
        RECT 22.144 34.404 22.176 36.912 ;
  LAYER M1 ;
        RECT 22.208 34.404 22.24 36.912 ;
  LAYER M1 ;
        RECT 22.272 34.404 22.304 36.912 ;
  LAYER M1 ;
        RECT 22.336 34.404 22.368 36.912 ;
  LAYER M1 ;
        RECT 22.4 34.404 22.432 36.912 ;
  LAYER M1 ;
        RECT 22.464 34.404 22.496 36.912 ;
  LAYER M1 ;
        RECT 22.528 34.404 22.56 36.912 ;
  LAYER M1 ;
        RECT 22.592 34.404 22.624 36.912 ;
  LAYER M1 ;
        RECT 22.656 34.404 22.688 36.912 ;
  LAYER M1 ;
        RECT 22.72 34.404 22.752 36.912 ;
  LAYER M1 ;
        RECT 22.784 34.404 22.816 36.912 ;
  LAYER M1 ;
        RECT 22.848 34.404 22.88 36.912 ;
  LAYER M1 ;
        RECT 22.912 34.404 22.944 36.912 ;
  LAYER M1 ;
        RECT 22.976 34.404 23.008 36.912 ;
  LAYER M1 ;
        RECT 23.04 34.404 23.072 36.912 ;
  LAYER M1 ;
        RECT 23.104 34.404 23.136 36.912 ;
  LAYER M1 ;
        RECT 23.168 34.404 23.2 36.912 ;
  LAYER M1 ;
        RECT 23.232 34.404 23.264 36.912 ;
  LAYER M1 ;
        RECT 23.296 34.404 23.328 36.912 ;
  LAYER M1 ;
        RECT 23.36 34.404 23.392 36.912 ;
  LAYER M1 ;
        RECT 23.424 34.404 23.456 36.912 ;
  LAYER M1 ;
        RECT 23.488 34.404 23.52 36.912 ;
  LAYER M1 ;
        RECT 23.552 34.404 23.584 36.912 ;
  LAYER M1 ;
        RECT 23.616 34.404 23.648 36.912 ;
  LAYER M1 ;
        RECT 23.68 34.404 23.712 36.912 ;
  LAYER M1 ;
        RECT 23.744 34.404 23.776 36.912 ;
  LAYER M1 ;
        RECT 23.808 34.404 23.84 36.912 ;
  LAYER M1 ;
        RECT 23.872 34.404 23.904 36.912 ;
  LAYER M1 ;
        RECT 23.936 34.404 23.968 36.912 ;
  LAYER M1 ;
        RECT 24 34.404 24.032 36.912 ;
  LAYER M1 ;
        RECT 24.064 34.404 24.096 36.912 ;
  LAYER M1 ;
        RECT 24.128 34.404 24.16 36.912 ;
  LAYER M2 ;
        RECT 21.804 36.796 24.276 36.828 ;
  LAYER M2 ;
        RECT 21.804 36.732 24.276 36.764 ;
  LAYER M2 ;
        RECT 21.804 36.668 24.276 36.7 ;
  LAYER M2 ;
        RECT 21.804 36.604 24.276 36.636 ;
  LAYER M2 ;
        RECT 21.804 36.54 24.276 36.572 ;
  LAYER M2 ;
        RECT 21.804 36.476 24.276 36.508 ;
  LAYER M2 ;
        RECT 21.804 36.412 24.276 36.444 ;
  LAYER M2 ;
        RECT 21.804 36.348 24.276 36.38 ;
  LAYER M2 ;
        RECT 21.804 36.284 24.276 36.316 ;
  LAYER M2 ;
        RECT 21.804 36.22 24.276 36.252 ;
  LAYER M2 ;
        RECT 21.804 36.156 24.276 36.188 ;
  LAYER M2 ;
        RECT 21.804 36.092 24.276 36.124 ;
  LAYER M2 ;
        RECT 21.804 36.028 24.276 36.06 ;
  LAYER M2 ;
        RECT 21.804 35.964 24.276 35.996 ;
  LAYER M2 ;
        RECT 21.804 35.9 24.276 35.932 ;
  LAYER M2 ;
        RECT 21.804 35.836 24.276 35.868 ;
  LAYER M2 ;
        RECT 21.804 35.772 24.276 35.804 ;
  LAYER M2 ;
        RECT 21.804 35.708 24.276 35.74 ;
  LAYER M2 ;
        RECT 21.804 35.644 24.276 35.676 ;
  LAYER M2 ;
        RECT 21.804 35.58 24.276 35.612 ;
  LAYER M2 ;
        RECT 21.804 35.516 24.276 35.548 ;
  LAYER M2 ;
        RECT 21.804 35.452 24.276 35.484 ;
  LAYER M2 ;
        RECT 21.804 35.388 24.276 35.42 ;
  LAYER M2 ;
        RECT 21.804 35.324 24.276 35.356 ;
  LAYER M2 ;
        RECT 21.804 35.26 24.276 35.292 ;
  LAYER M2 ;
        RECT 21.804 35.196 24.276 35.228 ;
  LAYER M2 ;
        RECT 21.804 35.132 24.276 35.164 ;
  LAYER M2 ;
        RECT 21.804 35.068 24.276 35.1 ;
  LAYER M2 ;
        RECT 21.804 35.004 24.276 35.036 ;
  LAYER M2 ;
        RECT 21.804 34.94 24.276 34.972 ;
  LAYER M2 ;
        RECT 21.804 34.876 24.276 34.908 ;
  LAYER M2 ;
        RECT 21.804 34.812 24.276 34.844 ;
  LAYER M2 ;
        RECT 21.804 34.748 24.276 34.78 ;
  LAYER M2 ;
        RECT 21.804 34.684 24.276 34.716 ;
  LAYER M2 ;
        RECT 21.804 34.62 24.276 34.652 ;
  LAYER M2 ;
        RECT 21.804 34.556 24.276 34.588 ;
  LAYER M3 ;
        RECT 21.824 34.404 21.856 36.912 ;
  LAYER M3 ;
        RECT 21.888 34.404 21.92 36.912 ;
  LAYER M3 ;
        RECT 21.952 34.404 21.984 36.912 ;
  LAYER M3 ;
        RECT 22.016 34.404 22.048 36.912 ;
  LAYER M3 ;
        RECT 22.08 34.404 22.112 36.912 ;
  LAYER M3 ;
        RECT 22.144 34.404 22.176 36.912 ;
  LAYER M3 ;
        RECT 22.208 34.404 22.24 36.912 ;
  LAYER M3 ;
        RECT 22.272 34.404 22.304 36.912 ;
  LAYER M3 ;
        RECT 22.336 34.404 22.368 36.912 ;
  LAYER M3 ;
        RECT 22.4 34.404 22.432 36.912 ;
  LAYER M3 ;
        RECT 22.464 34.404 22.496 36.912 ;
  LAYER M3 ;
        RECT 22.528 34.404 22.56 36.912 ;
  LAYER M3 ;
        RECT 22.592 34.404 22.624 36.912 ;
  LAYER M3 ;
        RECT 22.656 34.404 22.688 36.912 ;
  LAYER M3 ;
        RECT 22.72 34.404 22.752 36.912 ;
  LAYER M3 ;
        RECT 22.784 34.404 22.816 36.912 ;
  LAYER M3 ;
        RECT 22.848 34.404 22.88 36.912 ;
  LAYER M3 ;
        RECT 22.912 34.404 22.944 36.912 ;
  LAYER M3 ;
        RECT 22.976 34.404 23.008 36.912 ;
  LAYER M3 ;
        RECT 23.04 34.404 23.072 36.912 ;
  LAYER M3 ;
        RECT 23.104 34.404 23.136 36.912 ;
  LAYER M3 ;
        RECT 23.168 34.404 23.2 36.912 ;
  LAYER M3 ;
        RECT 23.232 34.404 23.264 36.912 ;
  LAYER M3 ;
        RECT 23.296 34.404 23.328 36.912 ;
  LAYER M3 ;
        RECT 23.36 34.404 23.392 36.912 ;
  LAYER M3 ;
        RECT 23.424 34.404 23.456 36.912 ;
  LAYER M3 ;
        RECT 23.488 34.404 23.52 36.912 ;
  LAYER M3 ;
        RECT 23.552 34.404 23.584 36.912 ;
  LAYER M3 ;
        RECT 23.616 34.404 23.648 36.912 ;
  LAYER M3 ;
        RECT 23.68 34.404 23.712 36.912 ;
  LAYER M3 ;
        RECT 23.744 34.404 23.776 36.912 ;
  LAYER M3 ;
        RECT 23.808 34.404 23.84 36.912 ;
  LAYER M3 ;
        RECT 23.872 34.404 23.904 36.912 ;
  LAYER M3 ;
        RECT 23.936 34.404 23.968 36.912 ;
  LAYER M3 ;
        RECT 24 34.404 24.032 36.912 ;
  LAYER M3 ;
        RECT 24.064 34.404 24.096 36.912 ;
  LAYER M3 ;
        RECT 24.128 34.404 24.16 36.912 ;
  LAYER M3 ;
        RECT 24.224 34.404 24.256 36.912 ;
  LAYER M1 ;
        RECT 21.839 34.44 21.841 36.876 ;
  LAYER M1 ;
        RECT 21.919 34.44 21.921 36.876 ;
  LAYER M1 ;
        RECT 21.999 34.44 22.001 36.876 ;
  LAYER M1 ;
        RECT 22.079 34.44 22.081 36.876 ;
  LAYER M1 ;
        RECT 22.159 34.44 22.161 36.876 ;
  LAYER M1 ;
        RECT 22.239 34.44 22.241 36.876 ;
  LAYER M1 ;
        RECT 22.319 34.44 22.321 36.876 ;
  LAYER M1 ;
        RECT 22.399 34.44 22.401 36.876 ;
  LAYER M1 ;
        RECT 22.479 34.44 22.481 36.876 ;
  LAYER M1 ;
        RECT 22.559 34.44 22.561 36.876 ;
  LAYER M1 ;
        RECT 22.639 34.44 22.641 36.876 ;
  LAYER M1 ;
        RECT 22.719 34.44 22.721 36.876 ;
  LAYER M1 ;
        RECT 22.799 34.44 22.801 36.876 ;
  LAYER M1 ;
        RECT 22.879 34.44 22.881 36.876 ;
  LAYER M1 ;
        RECT 22.959 34.44 22.961 36.876 ;
  LAYER M1 ;
        RECT 23.039 34.44 23.041 36.876 ;
  LAYER M1 ;
        RECT 23.119 34.44 23.121 36.876 ;
  LAYER M1 ;
        RECT 23.199 34.44 23.201 36.876 ;
  LAYER M1 ;
        RECT 23.279 34.44 23.281 36.876 ;
  LAYER M1 ;
        RECT 23.359 34.44 23.361 36.876 ;
  LAYER M1 ;
        RECT 23.439 34.44 23.441 36.876 ;
  LAYER M1 ;
        RECT 23.519 34.44 23.521 36.876 ;
  LAYER M1 ;
        RECT 23.599 34.44 23.601 36.876 ;
  LAYER M1 ;
        RECT 23.679 34.44 23.681 36.876 ;
  LAYER M1 ;
        RECT 23.759 34.44 23.761 36.876 ;
  LAYER M1 ;
        RECT 23.839 34.44 23.841 36.876 ;
  LAYER M1 ;
        RECT 23.919 34.44 23.921 36.876 ;
  LAYER M1 ;
        RECT 23.999 34.44 24.001 36.876 ;
  LAYER M1 ;
        RECT 24.079 34.44 24.081 36.876 ;
  LAYER M1 ;
        RECT 24.159 34.44 24.161 36.876 ;
  LAYER M2 ;
        RECT 21.84 36.875 24.24 36.877 ;
  LAYER M2 ;
        RECT 21.84 36.791 24.24 36.793 ;
  LAYER M2 ;
        RECT 21.84 36.707 24.24 36.709 ;
  LAYER M2 ;
        RECT 21.84 36.623 24.24 36.625 ;
  LAYER M2 ;
        RECT 21.84 36.539 24.24 36.541 ;
  LAYER M2 ;
        RECT 21.84 36.455 24.24 36.457 ;
  LAYER M2 ;
        RECT 21.84 36.371 24.24 36.373 ;
  LAYER M2 ;
        RECT 21.84 36.287 24.24 36.289 ;
  LAYER M2 ;
        RECT 21.84 36.203 24.24 36.205 ;
  LAYER M2 ;
        RECT 21.84 36.119 24.24 36.121 ;
  LAYER M2 ;
        RECT 21.84 36.035 24.24 36.037 ;
  LAYER M2 ;
        RECT 21.84 35.951 24.24 35.953 ;
  LAYER M2 ;
        RECT 21.84 35.8675 24.24 35.8695 ;
  LAYER M2 ;
        RECT 21.84 35.783 24.24 35.785 ;
  LAYER M2 ;
        RECT 21.84 35.699 24.24 35.701 ;
  LAYER M2 ;
        RECT 21.84 35.615 24.24 35.617 ;
  LAYER M2 ;
        RECT 21.84 35.531 24.24 35.533 ;
  LAYER M2 ;
        RECT 21.84 35.447 24.24 35.449 ;
  LAYER M2 ;
        RECT 21.84 35.363 24.24 35.365 ;
  LAYER M2 ;
        RECT 21.84 35.279 24.24 35.281 ;
  LAYER M2 ;
        RECT 21.84 35.195 24.24 35.197 ;
  LAYER M2 ;
        RECT 21.84 35.111 24.24 35.113 ;
  LAYER M2 ;
        RECT 21.84 35.027 24.24 35.029 ;
  LAYER M2 ;
        RECT 21.84 34.943 24.24 34.945 ;
  LAYER M2 ;
        RECT 21.84 34.859 24.24 34.861 ;
  LAYER M2 ;
        RECT 21.84 34.775 24.24 34.777 ;
  LAYER M2 ;
        RECT 21.84 34.691 24.24 34.693 ;
  LAYER M2 ;
        RECT 21.84 34.607 24.24 34.609 ;
  LAYER M2 ;
        RECT 21.84 34.523 24.24 34.525 ;
  LAYER M1 ;
        RECT 21.824 31.464 21.856 33.972 ;
  LAYER M1 ;
        RECT 21.888 31.464 21.92 33.972 ;
  LAYER M1 ;
        RECT 21.952 31.464 21.984 33.972 ;
  LAYER M1 ;
        RECT 22.016 31.464 22.048 33.972 ;
  LAYER M1 ;
        RECT 22.08 31.464 22.112 33.972 ;
  LAYER M1 ;
        RECT 22.144 31.464 22.176 33.972 ;
  LAYER M1 ;
        RECT 22.208 31.464 22.24 33.972 ;
  LAYER M1 ;
        RECT 22.272 31.464 22.304 33.972 ;
  LAYER M1 ;
        RECT 22.336 31.464 22.368 33.972 ;
  LAYER M1 ;
        RECT 22.4 31.464 22.432 33.972 ;
  LAYER M1 ;
        RECT 22.464 31.464 22.496 33.972 ;
  LAYER M1 ;
        RECT 22.528 31.464 22.56 33.972 ;
  LAYER M1 ;
        RECT 22.592 31.464 22.624 33.972 ;
  LAYER M1 ;
        RECT 22.656 31.464 22.688 33.972 ;
  LAYER M1 ;
        RECT 22.72 31.464 22.752 33.972 ;
  LAYER M1 ;
        RECT 22.784 31.464 22.816 33.972 ;
  LAYER M1 ;
        RECT 22.848 31.464 22.88 33.972 ;
  LAYER M1 ;
        RECT 22.912 31.464 22.944 33.972 ;
  LAYER M1 ;
        RECT 22.976 31.464 23.008 33.972 ;
  LAYER M1 ;
        RECT 23.04 31.464 23.072 33.972 ;
  LAYER M1 ;
        RECT 23.104 31.464 23.136 33.972 ;
  LAYER M1 ;
        RECT 23.168 31.464 23.2 33.972 ;
  LAYER M1 ;
        RECT 23.232 31.464 23.264 33.972 ;
  LAYER M1 ;
        RECT 23.296 31.464 23.328 33.972 ;
  LAYER M1 ;
        RECT 23.36 31.464 23.392 33.972 ;
  LAYER M1 ;
        RECT 23.424 31.464 23.456 33.972 ;
  LAYER M1 ;
        RECT 23.488 31.464 23.52 33.972 ;
  LAYER M1 ;
        RECT 23.552 31.464 23.584 33.972 ;
  LAYER M1 ;
        RECT 23.616 31.464 23.648 33.972 ;
  LAYER M1 ;
        RECT 23.68 31.464 23.712 33.972 ;
  LAYER M1 ;
        RECT 23.744 31.464 23.776 33.972 ;
  LAYER M1 ;
        RECT 23.808 31.464 23.84 33.972 ;
  LAYER M1 ;
        RECT 23.872 31.464 23.904 33.972 ;
  LAYER M1 ;
        RECT 23.936 31.464 23.968 33.972 ;
  LAYER M1 ;
        RECT 24 31.464 24.032 33.972 ;
  LAYER M1 ;
        RECT 24.064 31.464 24.096 33.972 ;
  LAYER M1 ;
        RECT 24.128 31.464 24.16 33.972 ;
  LAYER M2 ;
        RECT 21.804 33.856 24.276 33.888 ;
  LAYER M2 ;
        RECT 21.804 33.792 24.276 33.824 ;
  LAYER M2 ;
        RECT 21.804 33.728 24.276 33.76 ;
  LAYER M2 ;
        RECT 21.804 33.664 24.276 33.696 ;
  LAYER M2 ;
        RECT 21.804 33.6 24.276 33.632 ;
  LAYER M2 ;
        RECT 21.804 33.536 24.276 33.568 ;
  LAYER M2 ;
        RECT 21.804 33.472 24.276 33.504 ;
  LAYER M2 ;
        RECT 21.804 33.408 24.276 33.44 ;
  LAYER M2 ;
        RECT 21.804 33.344 24.276 33.376 ;
  LAYER M2 ;
        RECT 21.804 33.28 24.276 33.312 ;
  LAYER M2 ;
        RECT 21.804 33.216 24.276 33.248 ;
  LAYER M2 ;
        RECT 21.804 33.152 24.276 33.184 ;
  LAYER M2 ;
        RECT 21.804 33.088 24.276 33.12 ;
  LAYER M2 ;
        RECT 21.804 33.024 24.276 33.056 ;
  LAYER M2 ;
        RECT 21.804 32.96 24.276 32.992 ;
  LAYER M2 ;
        RECT 21.804 32.896 24.276 32.928 ;
  LAYER M2 ;
        RECT 21.804 32.832 24.276 32.864 ;
  LAYER M2 ;
        RECT 21.804 32.768 24.276 32.8 ;
  LAYER M2 ;
        RECT 21.804 32.704 24.276 32.736 ;
  LAYER M2 ;
        RECT 21.804 32.64 24.276 32.672 ;
  LAYER M2 ;
        RECT 21.804 32.576 24.276 32.608 ;
  LAYER M2 ;
        RECT 21.804 32.512 24.276 32.544 ;
  LAYER M2 ;
        RECT 21.804 32.448 24.276 32.48 ;
  LAYER M2 ;
        RECT 21.804 32.384 24.276 32.416 ;
  LAYER M2 ;
        RECT 21.804 32.32 24.276 32.352 ;
  LAYER M2 ;
        RECT 21.804 32.256 24.276 32.288 ;
  LAYER M2 ;
        RECT 21.804 32.192 24.276 32.224 ;
  LAYER M2 ;
        RECT 21.804 32.128 24.276 32.16 ;
  LAYER M2 ;
        RECT 21.804 32.064 24.276 32.096 ;
  LAYER M2 ;
        RECT 21.804 32 24.276 32.032 ;
  LAYER M2 ;
        RECT 21.804 31.936 24.276 31.968 ;
  LAYER M2 ;
        RECT 21.804 31.872 24.276 31.904 ;
  LAYER M2 ;
        RECT 21.804 31.808 24.276 31.84 ;
  LAYER M2 ;
        RECT 21.804 31.744 24.276 31.776 ;
  LAYER M2 ;
        RECT 21.804 31.68 24.276 31.712 ;
  LAYER M2 ;
        RECT 21.804 31.616 24.276 31.648 ;
  LAYER M3 ;
        RECT 21.824 31.464 21.856 33.972 ;
  LAYER M3 ;
        RECT 21.888 31.464 21.92 33.972 ;
  LAYER M3 ;
        RECT 21.952 31.464 21.984 33.972 ;
  LAYER M3 ;
        RECT 22.016 31.464 22.048 33.972 ;
  LAYER M3 ;
        RECT 22.08 31.464 22.112 33.972 ;
  LAYER M3 ;
        RECT 22.144 31.464 22.176 33.972 ;
  LAYER M3 ;
        RECT 22.208 31.464 22.24 33.972 ;
  LAYER M3 ;
        RECT 22.272 31.464 22.304 33.972 ;
  LAYER M3 ;
        RECT 22.336 31.464 22.368 33.972 ;
  LAYER M3 ;
        RECT 22.4 31.464 22.432 33.972 ;
  LAYER M3 ;
        RECT 22.464 31.464 22.496 33.972 ;
  LAYER M3 ;
        RECT 22.528 31.464 22.56 33.972 ;
  LAYER M3 ;
        RECT 22.592 31.464 22.624 33.972 ;
  LAYER M3 ;
        RECT 22.656 31.464 22.688 33.972 ;
  LAYER M3 ;
        RECT 22.72 31.464 22.752 33.972 ;
  LAYER M3 ;
        RECT 22.784 31.464 22.816 33.972 ;
  LAYER M3 ;
        RECT 22.848 31.464 22.88 33.972 ;
  LAYER M3 ;
        RECT 22.912 31.464 22.944 33.972 ;
  LAYER M3 ;
        RECT 22.976 31.464 23.008 33.972 ;
  LAYER M3 ;
        RECT 23.04 31.464 23.072 33.972 ;
  LAYER M3 ;
        RECT 23.104 31.464 23.136 33.972 ;
  LAYER M3 ;
        RECT 23.168 31.464 23.2 33.972 ;
  LAYER M3 ;
        RECT 23.232 31.464 23.264 33.972 ;
  LAYER M3 ;
        RECT 23.296 31.464 23.328 33.972 ;
  LAYER M3 ;
        RECT 23.36 31.464 23.392 33.972 ;
  LAYER M3 ;
        RECT 23.424 31.464 23.456 33.972 ;
  LAYER M3 ;
        RECT 23.488 31.464 23.52 33.972 ;
  LAYER M3 ;
        RECT 23.552 31.464 23.584 33.972 ;
  LAYER M3 ;
        RECT 23.616 31.464 23.648 33.972 ;
  LAYER M3 ;
        RECT 23.68 31.464 23.712 33.972 ;
  LAYER M3 ;
        RECT 23.744 31.464 23.776 33.972 ;
  LAYER M3 ;
        RECT 23.808 31.464 23.84 33.972 ;
  LAYER M3 ;
        RECT 23.872 31.464 23.904 33.972 ;
  LAYER M3 ;
        RECT 23.936 31.464 23.968 33.972 ;
  LAYER M3 ;
        RECT 24 31.464 24.032 33.972 ;
  LAYER M3 ;
        RECT 24.064 31.464 24.096 33.972 ;
  LAYER M3 ;
        RECT 24.128 31.464 24.16 33.972 ;
  LAYER M3 ;
        RECT 24.224 31.464 24.256 33.972 ;
  LAYER M1 ;
        RECT 21.839 31.5 21.841 33.936 ;
  LAYER M1 ;
        RECT 21.919 31.5 21.921 33.936 ;
  LAYER M1 ;
        RECT 21.999 31.5 22.001 33.936 ;
  LAYER M1 ;
        RECT 22.079 31.5 22.081 33.936 ;
  LAYER M1 ;
        RECT 22.159 31.5 22.161 33.936 ;
  LAYER M1 ;
        RECT 22.239 31.5 22.241 33.936 ;
  LAYER M1 ;
        RECT 22.319 31.5 22.321 33.936 ;
  LAYER M1 ;
        RECT 22.399 31.5 22.401 33.936 ;
  LAYER M1 ;
        RECT 22.479 31.5 22.481 33.936 ;
  LAYER M1 ;
        RECT 22.559 31.5 22.561 33.936 ;
  LAYER M1 ;
        RECT 22.639 31.5 22.641 33.936 ;
  LAYER M1 ;
        RECT 22.719 31.5 22.721 33.936 ;
  LAYER M1 ;
        RECT 22.799 31.5 22.801 33.936 ;
  LAYER M1 ;
        RECT 22.879 31.5 22.881 33.936 ;
  LAYER M1 ;
        RECT 22.959 31.5 22.961 33.936 ;
  LAYER M1 ;
        RECT 23.039 31.5 23.041 33.936 ;
  LAYER M1 ;
        RECT 23.119 31.5 23.121 33.936 ;
  LAYER M1 ;
        RECT 23.199 31.5 23.201 33.936 ;
  LAYER M1 ;
        RECT 23.279 31.5 23.281 33.936 ;
  LAYER M1 ;
        RECT 23.359 31.5 23.361 33.936 ;
  LAYER M1 ;
        RECT 23.439 31.5 23.441 33.936 ;
  LAYER M1 ;
        RECT 23.519 31.5 23.521 33.936 ;
  LAYER M1 ;
        RECT 23.599 31.5 23.601 33.936 ;
  LAYER M1 ;
        RECT 23.679 31.5 23.681 33.936 ;
  LAYER M1 ;
        RECT 23.759 31.5 23.761 33.936 ;
  LAYER M1 ;
        RECT 23.839 31.5 23.841 33.936 ;
  LAYER M1 ;
        RECT 23.919 31.5 23.921 33.936 ;
  LAYER M1 ;
        RECT 23.999 31.5 24.001 33.936 ;
  LAYER M1 ;
        RECT 24.079 31.5 24.081 33.936 ;
  LAYER M1 ;
        RECT 24.159 31.5 24.161 33.936 ;
  LAYER M2 ;
        RECT 21.84 33.935 24.24 33.937 ;
  LAYER M2 ;
        RECT 21.84 33.851 24.24 33.853 ;
  LAYER M2 ;
        RECT 21.84 33.767 24.24 33.769 ;
  LAYER M2 ;
        RECT 21.84 33.683 24.24 33.685 ;
  LAYER M2 ;
        RECT 21.84 33.599 24.24 33.601 ;
  LAYER M2 ;
        RECT 21.84 33.515 24.24 33.517 ;
  LAYER M2 ;
        RECT 21.84 33.431 24.24 33.433 ;
  LAYER M2 ;
        RECT 21.84 33.347 24.24 33.349 ;
  LAYER M2 ;
        RECT 21.84 33.263 24.24 33.265 ;
  LAYER M2 ;
        RECT 21.84 33.179 24.24 33.181 ;
  LAYER M2 ;
        RECT 21.84 33.095 24.24 33.097 ;
  LAYER M2 ;
        RECT 21.84 33.011 24.24 33.013 ;
  LAYER M2 ;
        RECT 21.84 32.9275 24.24 32.9295 ;
  LAYER M2 ;
        RECT 21.84 32.843 24.24 32.845 ;
  LAYER M2 ;
        RECT 21.84 32.759 24.24 32.761 ;
  LAYER M2 ;
        RECT 21.84 32.675 24.24 32.677 ;
  LAYER M2 ;
        RECT 21.84 32.591 24.24 32.593 ;
  LAYER M2 ;
        RECT 21.84 32.507 24.24 32.509 ;
  LAYER M2 ;
        RECT 21.84 32.423 24.24 32.425 ;
  LAYER M2 ;
        RECT 21.84 32.339 24.24 32.341 ;
  LAYER M2 ;
        RECT 21.84 32.255 24.24 32.257 ;
  LAYER M2 ;
        RECT 21.84 32.171 24.24 32.173 ;
  LAYER M2 ;
        RECT 21.84 32.087 24.24 32.089 ;
  LAYER M2 ;
        RECT 21.84 32.003 24.24 32.005 ;
  LAYER M2 ;
        RECT 21.84 31.919 24.24 31.921 ;
  LAYER M2 ;
        RECT 21.84 31.835 24.24 31.837 ;
  LAYER M2 ;
        RECT 21.84 31.751 24.24 31.753 ;
  LAYER M2 ;
        RECT 21.84 31.667 24.24 31.669 ;
  LAYER M2 ;
        RECT 21.84 31.583 24.24 31.585 ;
  LAYER M1 ;
        RECT 21.824 28.524 21.856 31.032 ;
  LAYER M1 ;
        RECT 21.888 28.524 21.92 31.032 ;
  LAYER M1 ;
        RECT 21.952 28.524 21.984 31.032 ;
  LAYER M1 ;
        RECT 22.016 28.524 22.048 31.032 ;
  LAYER M1 ;
        RECT 22.08 28.524 22.112 31.032 ;
  LAYER M1 ;
        RECT 22.144 28.524 22.176 31.032 ;
  LAYER M1 ;
        RECT 22.208 28.524 22.24 31.032 ;
  LAYER M1 ;
        RECT 22.272 28.524 22.304 31.032 ;
  LAYER M1 ;
        RECT 22.336 28.524 22.368 31.032 ;
  LAYER M1 ;
        RECT 22.4 28.524 22.432 31.032 ;
  LAYER M1 ;
        RECT 22.464 28.524 22.496 31.032 ;
  LAYER M1 ;
        RECT 22.528 28.524 22.56 31.032 ;
  LAYER M1 ;
        RECT 22.592 28.524 22.624 31.032 ;
  LAYER M1 ;
        RECT 22.656 28.524 22.688 31.032 ;
  LAYER M1 ;
        RECT 22.72 28.524 22.752 31.032 ;
  LAYER M1 ;
        RECT 22.784 28.524 22.816 31.032 ;
  LAYER M1 ;
        RECT 22.848 28.524 22.88 31.032 ;
  LAYER M1 ;
        RECT 22.912 28.524 22.944 31.032 ;
  LAYER M1 ;
        RECT 22.976 28.524 23.008 31.032 ;
  LAYER M1 ;
        RECT 23.04 28.524 23.072 31.032 ;
  LAYER M1 ;
        RECT 23.104 28.524 23.136 31.032 ;
  LAYER M1 ;
        RECT 23.168 28.524 23.2 31.032 ;
  LAYER M1 ;
        RECT 23.232 28.524 23.264 31.032 ;
  LAYER M1 ;
        RECT 23.296 28.524 23.328 31.032 ;
  LAYER M1 ;
        RECT 23.36 28.524 23.392 31.032 ;
  LAYER M1 ;
        RECT 23.424 28.524 23.456 31.032 ;
  LAYER M1 ;
        RECT 23.488 28.524 23.52 31.032 ;
  LAYER M1 ;
        RECT 23.552 28.524 23.584 31.032 ;
  LAYER M1 ;
        RECT 23.616 28.524 23.648 31.032 ;
  LAYER M1 ;
        RECT 23.68 28.524 23.712 31.032 ;
  LAYER M1 ;
        RECT 23.744 28.524 23.776 31.032 ;
  LAYER M1 ;
        RECT 23.808 28.524 23.84 31.032 ;
  LAYER M1 ;
        RECT 23.872 28.524 23.904 31.032 ;
  LAYER M1 ;
        RECT 23.936 28.524 23.968 31.032 ;
  LAYER M1 ;
        RECT 24 28.524 24.032 31.032 ;
  LAYER M1 ;
        RECT 24.064 28.524 24.096 31.032 ;
  LAYER M1 ;
        RECT 24.128 28.524 24.16 31.032 ;
  LAYER M2 ;
        RECT 21.804 30.916 24.276 30.948 ;
  LAYER M2 ;
        RECT 21.804 30.852 24.276 30.884 ;
  LAYER M2 ;
        RECT 21.804 30.788 24.276 30.82 ;
  LAYER M2 ;
        RECT 21.804 30.724 24.276 30.756 ;
  LAYER M2 ;
        RECT 21.804 30.66 24.276 30.692 ;
  LAYER M2 ;
        RECT 21.804 30.596 24.276 30.628 ;
  LAYER M2 ;
        RECT 21.804 30.532 24.276 30.564 ;
  LAYER M2 ;
        RECT 21.804 30.468 24.276 30.5 ;
  LAYER M2 ;
        RECT 21.804 30.404 24.276 30.436 ;
  LAYER M2 ;
        RECT 21.804 30.34 24.276 30.372 ;
  LAYER M2 ;
        RECT 21.804 30.276 24.276 30.308 ;
  LAYER M2 ;
        RECT 21.804 30.212 24.276 30.244 ;
  LAYER M2 ;
        RECT 21.804 30.148 24.276 30.18 ;
  LAYER M2 ;
        RECT 21.804 30.084 24.276 30.116 ;
  LAYER M2 ;
        RECT 21.804 30.02 24.276 30.052 ;
  LAYER M2 ;
        RECT 21.804 29.956 24.276 29.988 ;
  LAYER M2 ;
        RECT 21.804 29.892 24.276 29.924 ;
  LAYER M2 ;
        RECT 21.804 29.828 24.276 29.86 ;
  LAYER M2 ;
        RECT 21.804 29.764 24.276 29.796 ;
  LAYER M2 ;
        RECT 21.804 29.7 24.276 29.732 ;
  LAYER M2 ;
        RECT 21.804 29.636 24.276 29.668 ;
  LAYER M2 ;
        RECT 21.804 29.572 24.276 29.604 ;
  LAYER M2 ;
        RECT 21.804 29.508 24.276 29.54 ;
  LAYER M2 ;
        RECT 21.804 29.444 24.276 29.476 ;
  LAYER M2 ;
        RECT 21.804 29.38 24.276 29.412 ;
  LAYER M2 ;
        RECT 21.804 29.316 24.276 29.348 ;
  LAYER M2 ;
        RECT 21.804 29.252 24.276 29.284 ;
  LAYER M2 ;
        RECT 21.804 29.188 24.276 29.22 ;
  LAYER M2 ;
        RECT 21.804 29.124 24.276 29.156 ;
  LAYER M2 ;
        RECT 21.804 29.06 24.276 29.092 ;
  LAYER M2 ;
        RECT 21.804 28.996 24.276 29.028 ;
  LAYER M2 ;
        RECT 21.804 28.932 24.276 28.964 ;
  LAYER M2 ;
        RECT 21.804 28.868 24.276 28.9 ;
  LAYER M2 ;
        RECT 21.804 28.804 24.276 28.836 ;
  LAYER M2 ;
        RECT 21.804 28.74 24.276 28.772 ;
  LAYER M2 ;
        RECT 21.804 28.676 24.276 28.708 ;
  LAYER M3 ;
        RECT 21.824 28.524 21.856 31.032 ;
  LAYER M3 ;
        RECT 21.888 28.524 21.92 31.032 ;
  LAYER M3 ;
        RECT 21.952 28.524 21.984 31.032 ;
  LAYER M3 ;
        RECT 22.016 28.524 22.048 31.032 ;
  LAYER M3 ;
        RECT 22.08 28.524 22.112 31.032 ;
  LAYER M3 ;
        RECT 22.144 28.524 22.176 31.032 ;
  LAYER M3 ;
        RECT 22.208 28.524 22.24 31.032 ;
  LAYER M3 ;
        RECT 22.272 28.524 22.304 31.032 ;
  LAYER M3 ;
        RECT 22.336 28.524 22.368 31.032 ;
  LAYER M3 ;
        RECT 22.4 28.524 22.432 31.032 ;
  LAYER M3 ;
        RECT 22.464 28.524 22.496 31.032 ;
  LAYER M3 ;
        RECT 22.528 28.524 22.56 31.032 ;
  LAYER M3 ;
        RECT 22.592 28.524 22.624 31.032 ;
  LAYER M3 ;
        RECT 22.656 28.524 22.688 31.032 ;
  LAYER M3 ;
        RECT 22.72 28.524 22.752 31.032 ;
  LAYER M3 ;
        RECT 22.784 28.524 22.816 31.032 ;
  LAYER M3 ;
        RECT 22.848 28.524 22.88 31.032 ;
  LAYER M3 ;
        RECT 22.912 28.524 22.944 31.032 ;
  LAYER M3 ;
        RECT 22.976 28.524 23.008 31.032 ;
  LAYER M3 ;
        RECT 23.04 28.524 23.072 31.032 ;
  LAYER M3 ;
        RECT 23.104 28.524 23.136 31.032 ;
  LAYER M3 ;
        RECT 23.168 28.524 23.2 31.032 ;
  LAYER M3 ;
        RECT 23.232 28.524 23.264 31.032 ;
  LAYER M3 ;
        RECT 23.296 28.524 23.328 31.032 ;
  LAYER M3 ;
        RECT 23.36 28.524 23.392 31.032 ;
  LAYER M3 ;
        RECT 23.424 28.524 23.456 31.032 ;
  LAYER M3 ;
        RECT 23.488 28.524 23.52 31.032 ;
  LAYER M3 ;
        RECT 23.552 28.524 23.584 31.032 ;
  LAYER M3 ;
        RECT 23.616 28.524 23.648 31.032 ;
  LAYER M3 ;
        RECT 23.68 28.524 23.712 31.032 ;
  LAYER M3 ;
        RECT 23.744 28.524 23.776 31.032 ;
  LAYER M3 ;
        RECT 23.808 28.524 23.84 31.032 ;
  LAYER M3 ;
        RECT 23.872 28.524 23.904 31.032 ;
  LAYER M3 ;
        RECT 23.936 28.524 23.968 31.032 ;
  LAYER M3 ;
        RECT 24 28.524 24.032 31.032 ;
  LAYER M3 ;
        RECT 24.064 28.524 24.096 31.032 ;
  LAYER M3 ;
        RECT 24.128 28.524 24.16 31.032 ;
  LAYER M3 ;
        RECT 24.224 28.524 24.256 31.032 ;
  LAYER M1 ;
        RECT 21.839 28.56 21.841 30.996 ;
  LAYER M1 ;
        RECT 21.919 28.56 21.921 30.996 ;
  LAYER M1 ;
        RECT 21.999 28.56 22.001 30.996 ;
  LAYER M1 ;
        RECT 22.079 28.56 22.081 30.996 ;
  LAYER M1 ;
        RECT 22.159 28.56 22.161 30.996 ;
  LAYER M1 ;
        RECT 22.239 28.56 22.241 30.996 ;
  LAYER M1 ;
        RECT 22.319 28.56 22.321 30.996 ;
  LAYER M1 ;
        RECT 22.399 28.56 22.401 30.996 ;
  LAYER M1 ;
        RECT 22.479 28.56 22.481 30.996 ;
  LAYER M1 ;
        RECT 22.559 28.56 22.561 30.996 ;
  LAYER M1 ;
        RECT 22.639 28.56 22.641 30.996 ;
  LAYER M1 ;
        RECT 22.719 28.56 22.721 30.996 ;
  LAYER M1 ;
        RECT 22.799 28.56 22.801 30.996 ;
  LAYER M1 ;
        RECT 22.879 28.56 22.881 30.996 ;
  LAYER M1 ;
        RECT 22.959 28.56 22.961 30.996 ;
  LAYER M1 ;
        RECT 23.039 28.56 23.041 30.996 ;
  LAYER M1 ;
        RECT 23.119 28.56 23.121 30.996 ;
  LAYER M1 ;
        RECT 23.199 28.56 23.201 30.996 ;
  LAYER M1 ;
        RECT 23.279 28.56 23.281 30.996 ;
  LAYER M1 ;
        RECT 23.359 28.56 23.361 30.996 ;
  LAYER M1 ;
        RECT 23.439 28.56 23.441 30.996 ;
  LAYER M1 ;
        RECT 23.519 28.56 23.521 30.996 ;
  LAYER M1 ;
        RECT 23.599 28.56 23.601 30.996 ;
  LAYER M1 ;
        RECT 23.679 28.56 23.681 30.996 ;
  LAYER M1 ;
        RECT 23.759 28.56 23.761 30.996 ;
  LAYER M1 ;
        RECT 23.839 28.56 23.841 30.996 ;
  LAYER M1 ;
        RECT 23.919 28.56 23.921 30.996 ;
  LAYER M1 ;
        RECT 23.999 28.56 24.001 30.996 ;
  LAYER M1 ;
        RECT 24.079 28.56 24.081 30.996 ;
  LAYER M1 ;
        RECT 24.159 28.56 24.161 30.996 ;
  LAYER M2 ;
        RECT 21.84 30.995 24.24 30.997 ;
  LAYER M2 ;
        RECT 21.84 30.911 24.24 30.913 ;
  LAYER M2 ;
        RECT 21.84 30.827 24.24 30.829 ;
  LAYER M2 ;
        RECT 21.84 30.743 24.24 30.745 ;
  LAYER M2 ;
        RECT 21.84 30.659 24.24 30.661 ;
  LAYER M2 ;
        RECT 21.84 30.575 24.24 30.577 ;
  LAYER M2 ;
        RECT 21.84 30.491 24.24 30.493 ;
  LAYER M2 ;
        RECT 21.84 30.407 24.24 30.409 ;
  LAYER M2 ;
        RECT 21.84 30.323 24.24 30.325 ;
  LAYER M2 ;
        RECT 21.84 30.239 24.24 30.241 ;
  LAYER M2 ;
        RECT 21.84 30.155 24.24 30.157 ;
  LAYER M2 ;
        RECT 21.84 30.071 24.24 30.073 ;
  LAYER M2 ;
        RECT 21.84 29.9875 24.24 29.9895 ;
  LAYER M2 ;
        RECT 21.84 29.903 24.24 29.905 ;
  LAYER M2 ;
        RECT 21.84 29.819 24.24 29.821 ;
  LAYER M2 ;
        RECT 21.84 29.735 24.24 29.737 ;
  LAYER M2 ;
        RECT 21.84 29.651 24.24 29.653 ;
  LAYER M2 ;
        RECT 21.84 29.567 24.24 29.569 ;
  LAYER M2 ;
        RECT 21.84 29.483 24.24 29.485 ;
  LAYER M2 ;
        RECT 21.84 29.399 24.24 29.401 ;
  LAYER M2 ;
        RECT 21.84 29.315 24.24 29.317 ;
  LAYER M2 ;
        RECT 21.84 29.231 24.24 29.233 ;
  LAYER M2 ;
        RECT 21.84 29.147 24.24 29.149 ;
  LAYER M2 ;
        RECT 21.84 29.063 24.24 29.065 ;
  LAYER M2 ;
        RECT 21.84 28.979 24.24 28.981 ;
  LAYER M2 ;
        RECT 21.84 28.895 24.24 28.897 ;
  LAYER M2 ;
        RECT 21.84 28.811 24.24 28.813 ;
  LAYER M2 ;
        RECT 21.84 28.727 24.24 28.729 ;
  LAYER M2 ;
        RECT 21.84 28.643 24.24 28.645 ;
  LAYER M1 ;
        RECT 21.824 25.584 21.856 28.092 ;
  LAYER M1 ;
        RECT 21.888 25.584 21.92 28.092 ;
  LAYER M1 ;
        RECT 21.952 25.584 21.984 28.092 ;
  LAYER M1 ;
        RECT 22.016 25.584 22.048 28.092 ;
  LAYER M1 ;
        RECT 22.08 25.584 22.112 28.092 ;
  LAYER M1 ;
        RECT 22.144 25.584 22.176 28.092 ;
  LAYER M1 ;
        RECT 22.208 25.584 22.24 28.092 ;
  LAYER M1 ;
        RECT 22.272 25.584 22.304 28.092 ;
  LAYER M1 ;
        RECT 22.336 25.584 22.368 28.092 ;
  LAYER M1 ;
        RECT 22.4 25.584 22.432 28.092 ;
  LAYER M1 ;
        RECT 22.464 25.584 22.496 28.092 ;
  LAYER M1 ;
        RECT 22.528 25.584 22.56 28.092 ;
  LAYER M1 ;
        RECT 22.592 25.584 22.624 28.092 ;
  LAYER M1 ;
        RECT 22.656 25.584 22.688 28.092 ;
  LAYER M1 ;
        RECT 22.72 25.584 22.752 28.092 ;
  LAYER M1 ;
        RECT 22.784 25.584 22.816 28.092 ;
  LAYER M1 ;
        RECT 22.848 25.584 22.88 28.092 ;
  LAYER M1 ;
        RECT 22.912 25.584 22.944 28.092 ;
  LAYER M1 ;
        RECT 22.976 25.584 23.008 28.092 ;
  LAYER M1 ;
        RECT 23.04 25.584 23.072 28.092 ;
  LAYER M1 ;
        RECT 23.104 25.584 23.136 28.092 ;
  LAYER M1 ;
        RECT 23.168 25.584 23.2 28.092 ;
  LAYER M1 ;
        RECT 23.232 25.584 23.264 28.092 ;
  LAYER M1 ;
        RECT 23.296 25.584 23.328 28.092 ;
  LAYER M1 ;
        RECT 23.36 25.584 23.392 28.092 ;
  LAYER M1 ;
        RECT 23.424 25.584 23.456 28.092 ;
  LAYER M1 ;
        RECT 23.488 25.584 23.52 28.092 ;
  LAYER M1 ;
        RECT 23.552 25.584 23.584 28.092 ;
  LAYER M1 ;
        RECT 23.616 25.584 23.648 28.092 ;
  LAYER M1 ;
        RECT 23.68 25.584 23.712 28.092 ;
  LAYER M1 ;
        RECT 23.744 25.584 23.776 28.092 ;
  LAYER M1 ;
        RECT 23.808 25.584 23.84 28.092 ;
  LAYER M1 ;
        RECT 23.872 25.584 23.904 28.092 ;
  LAYER M1 ;
        RECT 23.936 25.584 23.968 28.092 ;
  LAYER M1 ;
        RECT 24 25.584 24.032 28.092 ;
  LAYER M1 ;
        RECT 24.064 25.584 24.096 28.092 ;
  LAYER M1 ;
        RECT 24.128 25.584 24.16 28.092 ;
  LAYER M2 ;
        RECT 21.804 27.976 24.276 28.008 ;
  LAYER M2 ;
        RECT 21.804 27.912 24.276 27.944 ;
  LAYER M2 ;
        RECT 21.804 27.848 24.276 27.88 ;
  LAYER M2 ;
        RECT 21.804 27.784 24.276 27.816 ;
  LAYER M2 ;
        RECT 21.804 27.72 24.276 27.752 ;
  LAYER M2 ;
        RECT 21.804 27.656 24.276 27.688 ;
  LAYER M2 ;
        RECT 21.804 27.592 24.276 27.624 ;
  LAYER M2 ;
        RECT 21.804 27.528 24.276 27.56 ;
  LAYER M2 ;
        RECT 21.804 27.464 24.276 27.496 ;
  LAYER M2 ;
        RECT 21.804 27.4 24.276 27.432 ;
  LAYER M2 ;
        RECT 21.804 27.336 24.276 27.368 ;
  LAYER M2 ;
        RECT 21.804 27.272 24.276 27.304 ;
  LAYER M2 ;
        RECT 21.804 27.208 24.276 27.24 ;
  LAYER M2 ;
        RECT 21.804 27.144 24.276 27.176 ;
  LAYER M2 ;
        RECT 21.804 27.08 24.276 27.112 ;
  LAYER M2 ;
        RECT 21.804 27.016 24.276 27.048 ;
  LAYER M2 ;
        RECT 21.804 26.952 24.276 26.984 ;
  LAYER M2 ;
        RECT 21.804 26.888 24.276 26.92 ;
  LAYER M2 ;
        RECT 21.804 26.824 24.276 26.856 ;
  LAYER M2 ;
        RECT 21.804 26.76 24.276 26.792 ;
  LAYER M2 ;
        RECT 21.804 26.696 24.276 26.728 ;
  LAYER M2 ;
        RECT 21.804 26.632 24.276 26.664 ;
  LAYER M2 ;
        RECT 21.804 26.568 24.276 26.6 ;
  LAYER M2 ;
        RECT 21.804 26.504 24.276 26.536 ;
  LAYER M2 ;
        RECT 21.804 26.44 24.276 26.472 ;
  LAYER M2 ;
        RECT 21.804 26.376 24.276 26.408 ;
  LAYER M2 ;
        RECT 21.804 26.312 24.276 26.344 ;
  LAYER M2 ;
        RECT 21.804 26.248 24.276 26.28 ;
  LAYER M2 ;
        RECT 21.804 26.184 24.276 26.216 ;
  LAYER M2 ;
        RECT 21.804 26.12 24.276 26.152 ;
  LAYER M2 ;
        RECT 21.804 26.056 24.276 26.088 ;
  LAYER M2 ;
        RECT 21.804 25.992 24.276 26.024 ;
  LAYER M2 ;
        RECT 21.804 25.928 24.276 25.96 ;
  LAYER M2 ;
        RECT 21.804 25.864 24.276 25.896 ;
  LAYER M2 ;
        RECT 21.804 25.8 24.276 25.832 ;
  LAYER M2 ;
        RECT 21.804 25.736 24.276 25.768 ;
  LAYER M3 ;
        RECT 21.824 25.584 21.856 28.092 ;
  LAYER M3 ;
        RECT 21.888 25.584 21.92 28.092 ;
  LAYER M3 ;
        RECT 21.952 25.584 21.984 28.092 ;
  LAYER M3 ;
        RECT 22.016 25.584 22.048 28.092 ;
  LAYER M3 ;
        RECT 22.08 25.584 22.112 28.092 ;
  LAYER M3 ;
        RECT 22.144 25.584 22.176 28.092 ;
  LAYER M3 ;
        RECT 22.208 25.584 22.24 28.092 ;
  LAYER M3 ;
        RECT 22.272 25.584 22.304 28.092 ;
  LAYER M3 ;
        RECT 22.336 25.584 22.368 28.092 ;
  LAYER M3 ;
        RECT 22.4 25.584 22.432 28.092 ;
  LAYER M3 ;
        RECT 22.464 25.584 22.496 28.092 ;
  LAYER M3 ;
        RECT 22.528 25.584 22.56 28.092 ;
  LAYER M3 ;
        RECT 22.592 25.584 22.624 28.092 ;
  LAYER M3 ;
        RECT 22.656 25.584 22.688 28.092 ;
  LAYER M3 ;
        RECT 22.72 25.584 22.752 28.092 ;
  LAYER M3 ;
        RECT 22.784 25.584 22.816 28.092 ;
  LAYER M3 ;
        RECT 22.848 25.584 22.88 28.092 ;
  LAYER M3 ;
        RECT 22.912 25.584 22.944 28.092 ;
  LAYER M3 ;
        RECT 22.976 25.584 23.008 28.092 ;
  LAYER M3 ;
        RECT 23.04 25.584 23.072 28.092 ;
  LAYER M3 ;
        RECT 23.104 25.584 23.136 28.092 ;
  LAYER M3 ;
        RECT 23.168 25.584 23.2 28.092 ;
  LAYER M3 ;
        RECT 23.232 25.584 23.264 28.092 ;
  LAYER M3 ;
        RECT 23.296 25.584 23.328 28.092 ;
  LAYER M3 ;
        RECT 23.36 25.584 23.392 28.092 ;
  LAYER M3 ;
        RECT 23.424 25.584 23.456 28.092 ;
  LAYER M3 ;
        RECT 23.488 25.584 23.52 28.092 ;
  LAYER M3 ;
        RECT 23.552 25.584 23.584 28.092 ;
  LAYER M3 ;
        RECT 23.616 25.584 23.648 28.092 ;
  LAYER M3 ;
        RECT 23.68 25.584 23.712 28.092 ;
  LAYER M3 ;
        RECT 23.744 25.584 23.776 28.092 ;
  LAYER M3 ;
        RECT 23.808 25.584 23.84 28.092 ;
  LAYER M3 ;
        RECT 23.872 25.584 23.904 28.092 ;
  LAYER M3 ;
        RECT 23.936 25.584 23.968 28.092 ;
  LAYER M3 ;
        RECT 24 25.584 24.032 28.092 ;
  LAYER M3 ;
        RECT 24.064 25.584 24.096 28.092 ;
  LAYER M3 ;
        RECT 24.128 25.584 24.16 28.092 ;
  LAYER M3 ;
        RECT 24.224 25.584 24.256 28.092 ;
  LAYER M1 ;
        RECT 21.839 25.62 21.841 28.056 ;
  LAYER M1 ;
        RECT 21.919 25.62 21.921 28.056 ;
  LAYER M1 ;
        RECT 21.999 25.62 22.001 28.056 ;
  LAYER M1 ;
        RECT 22.079 25.62 22.081 28.056 ;
  LAYER M1 ;
        RECT 22.159 25.62 22.161 28.056 ;
  LAYER M1 ;
        RECT 22.239 25.62 22.241 28.056 ;
  LAYER M1 ;
        RECT 22.319 25.62 22.321 28.056 ;
  LAYER M1 ;
        RECT 22.399 25.62 22.401 28.056 ;
  LAYER M1 ;
        RECT 22.479 25.62 22.481 28.056 ;
  LAYER M1 ;
        RECT 22.559 25.62 22.561 28.056 ;
  LAYER M1 ;
        RECT 22.639 25.62 22.641 28.056 ;
  LAYER M1 ;
        RECT 22.719 25.62 22.721 28.056 ;
  LAYER M1 ;
        RECT 22.799 25.62 22.801 28.056 ;
  LAYER M1 ;
        RECT 22.879 25.62 22.881 28.056 ;
  LAYER M1 ;
        RECT 22.959 25.62 22.961 28.056 ;
  LAYER M1 ;
        RECT 23.039 25.62 23.041 28.056 ;
  LAYER M1 ;
        RECT 23.119 25.62 23.121 28.056 ;
  LAYER M1 ;
        RECT 23.199 25.62 23.201 28.056 ;
  LAYER M1 ;
        RECT 23.279 25.62 23.281 28.056 ;
  LAYER M1 ;
        RECT 23.359 25.62 23.361 28.056 ;
  LAYER M1 ;
        RECT 23.439 25.62 23.441 28.056 ;
  LAYER M1 ;
        RECT 23.519 25.62 23.521 28.056 ;
  LAYER M1 ;
        RECT 23.599 25.62 23.601 28.056 ;
  LAYER M1 ;
        RECT 23.679 25.62 23.681 28.056 ;
  LAYER M1 ;
        RECT 23.759 25.62 23.761 28.056 ;
  LAYER M1 ;
        RECT 23.839 25.62 23.841 28.056 ;
  LAYER M1 ;
        RECT 23.919 25.62 23.921 28.056 ;
  LAYER M1 ;
        RECT 23.999 25.62 24.001 28.056 ;
  LAYER M1 ;
        RECT 24.079 25.62 24.081 28.056 ;
  LAYER M1 ;
        RECT 24.159 25.62 24.161 28.056 ;
  LAYER M2 ;
        RECT 21.84 28.055 24.24 28.057 ;
  LAYER M2 ;
        RECT 21.84 27.971 24.24 27.973 ;
  LAYER M2 ;
        RECT 21.84 27.887 24.24 27.889 ;
  LAYER M2 ;
        RECT 21.84 27.803 24.24 27.805 ;
  LAYER M2 ;
        RECT 21.84 27.719 24.24 27.721 ;
  LAYER M2 ;
        RECT 21.84 27.635 24.24 27.637 ;
  LAYER M2 ;
        RECT 21.84 27.551 24.24 27.553 ;
  LAYER M2 ;
        RECT 21.84 27.467 24.24 27.469 ;
  LAYER M2 ;
        RECT 21.84 27.383 24.24 27.385 ;
  LAYER M2 ;
        RECT 21.84 27.299 24.24 27.301 ;
  LAYER M2 ;
        RECT 21.84 27.215 24.24 27.217 ;
  LAYER M2 ;
        RECT 21.84 27.131 24.24 27.133 ;
  LAYER M2 ;
        RECT 21.84 27.0475 24.24 27.0495 ;
  LAYER M2 ;
        RECT 21.84 26.963 24.24 26.965 ;
  LAYER M2 ;
        RECT 21.84 26.879 24.24 26.881 ;
  LAYER M2 ;
        RECT 21.84 26.795 24.24 26.797 ;
  LAYER M2 ;
        RECT 21.84 26.711 24.24 26.713 ;
  LAYER M2 ;
        RECT 21.84 26.627 24.24 26.629 ;
  LAYER M2 ;
        RECT 21.84 26.543 24.24 26.545 ;
  LAYER M2 ;
        RECT 21.84 26.459 24.24 26.461 ;
  LAYER M2 ;
        RECT 21.84 26.375 24.24 26.377 ;
  LAYER M2 ;
        RECT 21.84 26.291 24.24 26.293 ;
  LAYER M2 ;
        RECT 21.84 26.207 24.24 26.209 ;
  LAYER M2 ;
        RECT 21.84 26.123 24.24 26.125 ;
  LAYER M2 ;
        RECT 21.84 26.039 24.24 26.041 ;
  LAYER M2 ;
        RECT 21.84 25.955 24.24 25.957 ;
  LAYER M2 ;
        RECT 21.84 25.871 24.24 25.873 ;
  LAYER M2 ;
        RECT 21.84 25.787 24.24 25.789 ;
  LAYER M2 ;
        RECT 21.84 25.703 24.24 25.705 ;
  LAYER M1 ;
        RECT 21.824 22.644 21.856 25.152 ;
  LAYER M1 ;
        RECT 21.888 22.644 21.92 25.152 ;
  LAYER M1 ;
        RECT 21.952 22.644 21.984 25.152 ;
  LAYER M1 ;
        RECT 22.016 22.644 22.048 25.152 ;
  LAYER M1 ;
        RECT 22.08 22.644 22.112 25.152 ;
  LAYER M1 ;
        RECT 22.144 22.644 22.176 25.152 ;
  LAYER M1 ;
        RECT 22.208 22.644 22.24 25.152 ;
  LAYER M1 ;
        RECT 22.272 22.644 22.304 25.152 ;
  LAYER M1 ;
        RECT 22.336 22.644 22.368 25.152 ;
  LAYER M1 ;
        RECT 22.4 22.644 22.432 25.152 ;
  LAYER M1 ;
        RECT 22.464 22.644 22.496 25.152 ;
  LAYER M1 ;
        RECT 22.528 22.644 22.56 25.152 ;
  LAYER M1 ;
        RECT 22.592 22.644 22.624 25.152 ;
  LAYER M1 ;
        RECT 22.656 22.644 22.688 25.152 ;
  LAYER M1 ;
        RECT 22.72 22.644 22.752 25.152 ;
  LAYER M1 ;
        RECT 22.784 22.644 22.816 25.152 ;
  LAYER M1 ;
        RECT 22.848 22.644 22.88 25.152 ;
  LAYER M1 ;
        RECT 22.912 22.644 22.944 25.152 ;
  LAYER M1 ;
        RECT 22.976 22.644 23.008 25.152 ;
  LAYER M1 ;
        RECT 23.04 22.644 23.072 25.152 ;
  LAYER M1 ;
        RECT 23.104 22.644 23.136 25.152 ;
  LAYER M1 ;
        RECT 23.168 22.644 23.2 25.152 ;
  LAYER M1 ;
        RECT 23.232 22.644 23.264 25.152 ;
  LAYER M1 ;
        RECT 23.296 22.644 23.328 25.152 ;
  LAYER M1 ;
        RECT 23.36 22.644 23.392 25.152 ;
  LAYER M1 ;
        RECT 23.424 22.644 23.456 25.152 ;
  LAYER M1 ;
        RECT 23.488 22.644 23.52 25.152 ;
  LAYER M1 ;
        RECT 23.552 22.644 23.584 25.152 ;
  LAYER M1 ;
        RECT 23.616 22.644 23.648 25.152 ;
  LAYER M1 ;
        RECT 23.68 22.644 23.712 25.152 ;
  LAYER M1 ;
        RECT 23.744 22.644 23.776 25.152 ;
  LAYER M1 ;
        RECT 23.808 22.644 23.84 25.152 ;
  LAYER M1 ;
        RECT 23.872 22.644 23.904 25.152 ;
  LAYER M1 ;
        RECT 23.936 22.644 23.968 25.152 ;
  LAYER M1 ;
        RECT 24 22.644 24.032 25.152 ;
  LAYER M1 ;
        RECT 24.064 22.644 24.096 25.152 ;
  LAYER M1 ;
        RECT 24.128 22.644 24.16 25.152 ;
  LAYER M2 ;
        RECT 21.804 25.036 24.276 25.068 ;
  LAYER M2 ;
        RECT 21.804 24.972 24.276 25.004 ;
  LAYER M2 ;
        RECT 21.804 24.908 24.276 24.94 ;
  LAYER M2 ;
        RECT 21.804 24.844 24.276 24.876 ;
  LAYER M2 ;
        RECT 21.804 24.78 24.276 24.812 ;
  LAYER M2 ;
        RECT 21.804 24.716 24.276 24.748 ;
  LAYER M2 ;
        RECT 21.804 24.652 24.276 24.684 ;
  LAYER M2 ;
        RECT 21.804 24.588 24.276 24.62 ;
  LAYER M2 ;
        RECT 21.804 24.524 24.276 24.556 ;
  LAYER M2 ;
        RECT 21.804 24.46 24.276 24.492 ;
  LAYER M2 ;
        RECT 21.804 24.396 24.276 24.428 ;
  LAYER M2 ;
        RECT 21.804 24.332 24.276 24.364 ;
  LAYER M2 ;
        RECT 21.804 24.268 24.276 24.3 ;
  LAYER M2 ;
        RECT 21.804 24.204 24.276 24.236 ;
  LAYER M2 ;
        RECT 21.804 24.14 24.276 24.172 ;
  LAYER M2 ;
        RECT 21.804 24.076 24.276 24.108 ;
  LAYER M2 ;
        RECT 21.804 24.012 24.276 24.044 ;
  LAYER M2 ;
        RECT 21.804 23.948 24.276 23.98 ;
  LAYER M2 ;
        RECT 21.804 23.884 24.276 23.916 ;
  LAYER M2 ;
        RECT 21.804 23.82 24.276 23.852 ;
  LAYER M2 ;
        RECT 21.804 23.756 24.276 23.788 ;
  LAYER M2 ;
        RECT 21.804 23.692 24.276 23.724 ;
  LAYER M2 ;
        RECT 21.804 23.628 24.276 23.66 ;
  LAYER M2 ;
        RECT 21.804 23.564 24.276 23.596 ;
  LAYER M2 ;
        RECT 21.804 23.5 24.276 23.532 ;
  LAYER M2 ;
        RECT 21.804 23.436 24.276 23.468 ;
  LAYER M2 ;
        RECT 21.804 23.372 24.276 23.404 ;
  LAYER M2 ;
        RECT 21.804 23.308 24.276 23.34 ;
  LAYER M2 ;
        RECT 21.804 23.244 24.276 23.276 ;
  LAYER M2 ;
        RECT 21.804 23.18 24.276 23.212 ;
  LAYER M2 ;
        RECT 21.804 23.116 24.276 23.148 ;
  LAYER M2 ;
        RECT 21.804 23.052 24.276 23.084 ;
  LAYER M2 ;
        RECT 21.804 22.988 24.276 23.02 ;
  LAYER M2 ;
        RECT 21.804 22.924 24.276 22.956 ;
  LAYER M2 ;
        RECT 21.804 22.86 24.276 22.892 ;
  LAYER M2 ;
        RECT 21.804 22.796 24.276 22.828 ;
  LAYER M3 ;
        RECT 21.824 22.644 21.856 25.152 ;
  LAYER M3 ;
        RECT 21.888 22.644 21.92 25.152 ;
  LAYER M3 ;
        RECT 21.952 22.644 21.984 25.152 ;
  LAYER M3 ;
        RECT 22.016 22.644 22.048 25.152 ;
  LAYER M3 ;
        RECT 22.08 22.644 22.112 25.152 ;
  LAYER M3 ;
        RECT 22.144 22.644 22.176 25.152 ;
  LAYER M3 ;
        RECT 22.208 22.644 22.24 25.152 ;
  LAYER M3 ;
        RECT 22.272 22.644 22.304 25.152 ;
  LAYER M3 ;
        RECT 22.336 22.644 22.368 25.152 ;
  LAYER M3 ;
        RECT 22.4 22.644 22.432 25.152 ;
  LAYER M3 ;
        RECT 22.464 22.644 22.496 25.152 ;
  LAYER M3 ;
        RECT 22.528 22.644 22.56 25.152 ;
  LAYER M3 ;
        RECT 22.592 22.644 22.624 25.152 ;
  LAYER M3 ;
        RECT 22.656 22.644 22.688 25.152 ;
  LAYER M3 ;
        RECT 22.72 22.644 22.752 25.152 ;
  LAYER M3 ;
        RECT 22.784 22.644 22.816 25.152 ;
  LAYER M3 ;
        RECT 22.848 22.644 22.88 25.152 ;
  LAYER M3 ;
        RECT 22.912 22.644 22.944 25.152 ;
  LAYER M3 ;
        RECT 22.976 22.644 23.008 25.152 ;
  LAYER M3 ;
        RECT 23.04 22.644 23.072 25.152 ;
  LAYER M3 ;
        RECT 23.104 22.644 23.136 25.152 ;
  LAYER M3 ;
        RECT 23.168 22.644 23.2 25.152 ;
  LAYER M3 ;
        RECT 23.232 22.644 23.264 25.152 ;
  LAYER M3 ;
        RECT 23.296 22.644 23.328 25.152 ;
  LAYER M3 ;
        RECT 23.36 22.644 23.392 25.152 ;
  LAYER M3 ;
        RECT 23.424 22.644 23.456 25.152 ;
  LAYER M3 ;
        RECT 23.488 22.644 23.52 25.152 ;
  LAYER M3 ;
        RECT 23.552 22.644 23.584 25.152 ;
  LAYER M3 ;
        RECT 23.616 22.644 23.648 25.152 ;
  LAYER M3 ;
        RECT 23.68 22.644 23.712 25.152 ;
  LAYER M3 ;
        RECT 23.744 22.644 23.776 25.152 ;
  LAYER M3 ;
        RECT 23.808 22.644 23.84 25.152 ;
  LAYER M3 ;
        RECT 23.872 22.644 23.904 25.152 ;
  LAYER M3 ;
        RECT 23.936 22.644 23.968 25.152 ;
  LAYER M3 ;
        RECT 24 22.644 24.032 25.152 ;
  LAYER M3 ;
        RECT 24.064 22.644 24.096 25.152 ;
  LAYER M3 ;
        RECT 24.128 22.644 24.16 25.152 ;
  LAYER M3 ;
        RECT 24.224 22.644 24.256 25.152 ;
  LAYER M1 ;
        RECT 21.839 22.68 21.841 25.116 ;
  LAYER M1 ;
        RECT 21.919 22.68 21.921 25.116 ;
  LAYER M1 ;
        RECT 21.999 22.68 22.001 25.116 ;
  LAYER M1 ;
        RECT 22.079 22.68 22.081 25.116 ;
  LAYER M1 ;
        RECT 22.159 22.68 22.161 25.116 ;
  LAYER M1 ;
        RECT 22.239 22.68 22.241 25.116 ;
  LAYER M1 ;
        RECT 22.319 22.68 22.321 25.116 ;
  LAYER M1 ;
        RECT 22.399 22.68 22.401 25.116 ;
  LAYER M1 ;
        RECT 22.479 22.68 22.481 25.116 ;
  LAYER M1 ;
        RECT 22.559 22.68 22.561 25.116 ;
  LAYER M1 ;
        RECT 22.639 22.68 22.641 25.116 ;
  LAYER M1 ;
        RECT 22.719 22.68 22.721 25.116 ;
  LAYER M1 ;
        RECT 22.799 22.68 22.801 25.116 ;
  LAYER M1 ;
        RECT 22.879 22.68 22.881 25.116 ;
  LAYER M1 ;
        RECT 22.959 22.68 22.961 25.116 ;
  LAYER M1 ;
        RECT 23.039 22.68 23.041 25.116 ;
  LAYER M1 ;
        RECT 23.119 22.68 23.121 25.116 ;
  LAYER M1 ;
        RECT 23.199 22.68 23.201 25.116 ;
  LAYER M1 ;
        RECT 23.279 22.68 23.281 25.116 ;
  LAYER M1 ;
        RECT 23.359 22.68 23.361 25.116 ;
  LAYER M1 ;
        RECT 23.439 22.68 23.441 25.116 ;
  LAYER M1 ;
        RECT 23.519 22.68 23.521 25.116 ;
  LAYER M1 ;
        RECT 23.599 22.68 23.601 25.116 ;
  LAYER M1 ;
        RECT 23.679 22.68 23.681 25.116 ;
  LAYER M1 ;
        RECT 23.759 22.68 23.761 25.116 ;
  LAYER M1 ;
        RECT 23.839 22.68 23.841 25.116 ;
  LAYER M1 ;
        RECT 23.919 22.68 23.921 25.116 ;
  LAYER M1 ;
        RECT 23.999 22.68 24.001 25.116 ;
  LAYER M1 ;
        RECT 24.079 22.68 24.081 25.116 ;
  LAYER M1 ;
        RECT 24.159 22.68 24.161 25.116 ;
  LAYER M2 ;
        RECT 21.84 25.115 24.24 25.117 ;
  LAYER M2 ;
        RECT 21.84 25.031 24.24 25.033 ;
  LAYER M2 ;
        RECT 21.84 24.947 24.24 24.949 ;
  LAYER M2 ;
        RECT 21.84 24.863 24.24 24.865 ;
  LAYER M2 ;
        RECT 21.84 24.779 24.24 24.781 ;
  LAYER M2 ;
        RECT 21.84 24.695 24.24 24.697 ;
  LAYER M2 ;
        RECT 21.84 24.611 24.24 24.613 ;
  LAYER M2 ;
        RECT 21.84 24.527 24.24 24.529 ;
  LAYER M2 ;
        RECT 21.84 24.443 24.24 24.445 ;
  LAYER M2 ;
        RECT 21.84 24.359 24.24 24.361 ;
  LAYER M2 ;
        RECT 21.84 24.275 24.24 24.277 ;
  LAYER M2 ;
        RECT 21.84 24.191 24.24 24.193 ;
  LAYER M2 ;
        RECT 21.84 24.1075 24.24 24.1095 ;
  LAYER M2 ;
        RECT 21.84 24.023 24.24 24.025 ;
  LAYER M2 ;
        RECT 21.84 23.939 24.24 23.941 ;
  LAYER M2 ;
        RECT 21.84 23.855 24.24 23.857 ;
  LAYER M2 ;
        RECT 21.84 23.771 24.24 23.773 ;
  LAYER M2 ;
        RECT 21.84 23.687 24.24 23.689 ;
  LAYER M2 ;
        RECT 21.84 23.603 24.24 23.605 ;
  LAYER M2 ;
        RECT 21.84 23.519 24.24 23.521 ;
  LAYER M2 ;
        RECT 21.84 23.435 24.24 23.437 ;
  LAYER M2 ;
        RECT 21.84 23.351 24.24 23.353 ;
  LAYER M2 ;
        RECT 21.84 23.267 24.24 23.269 ;
  LAYER M2 ;
        RECT 21.84 23.183 24.24 23.185 ;
  LAYER M2 ;
        RECT 21.84 23.099 24.24 23.101 ;
  LAYER M2 ;
        RECT 21.84 23.015 24.24 23.017 ;
  LAYER M2 ;
        RECT 21.84 22.931 24.24 22.933 ;
  LAYER M2 ;
        RECT 21.84 22.847 24.24 22.849 ;
  LAYER M2 ;
        RECT 21.84 22.763 24.24 22.765 ;
  LAYER M1 ;
        RECT 21.824 19.704 21.856 22.212 ;
  LAYER M1 ;
        RECT 21.888 19.704 21.92 22.212 ;
  LAYER M1 ;
        RECT 21.952 19.704 21.984 22.212 ;
  LAYER M1 ;
        RECT 22.016 19.704 22.048 22.212 ;
  LAYER M1 ;
        RECT 22.08 19.704 22.112 22.212 ;
  LAYER M1 ;
        RECT 22.144 19.704 22.176 22.212 ;
  LAYER M1 ;
        RECT 22.208 19.704 22.24 22.212 ;
  LAYER M1 ;
        RECT 22.272 19.704 22.304 22.212 ;
  LAYER M1 ;
        RECT 22.336 19.704 22.368 22.212 ;
  LAYER M1 ;
        RECT 22.4 19.704 22.432 22.212 ;
  LAYER M1 ;
        RECT 22.464 19.704 22.496 22.212 ;
  LAYER M1 ;
        RECT 22.528 19.704 22.56 22.212 ;
  LAYER M1 ;
        RECT 22.592 19.704 22.624 22.212 ;
  LAYER M1 ;
        RECT 22.656 19.704 22.688 22.212 ;
  LAYER M1 ;
        RECT 22.72 19.704 22.752 22.212 ;
  LAYER M1 ;
        RECT 22.784 19.704 22.816 22.212 ;
  LAYER M1 ;
        RECT 22.848 19.704 22.88 22.212 ;
  LAYER M1 ;
        RECT 22.912 19.704 22.944 22.212 ;
  LAYER M1 ;
        RECT 22.976 19.704 23.008 22.212 ;
  LAYER M1 ;
        RECT 23.04 19.704 23.072 22.212 ;
  LAYER M1 ;
        RECT 23.104 19.704 23.136 22.212 ;
  LAYER M1 ;
        RECT 23.168 19.704 23.2 22.212 ;
  LAYER M1 ;
        RECT 23.232 19.704 23.264 22.212 ;
  LAYER M1 ;
        RECT 23.296 19.704 23.328 22.212 ;
  LAYER M1 ;
        RECT 23.36 19.704 23.392 22.212 ;
  LAYER M1 ;
        RECT 23.424 19.704 23.456 22.212 ;
  LAYER M1 ;
        RECT 23.488 19.704 23.52 22.212 ;
  LAYER M1 ;
        RECT 23.552 19.704 23.584 22.212 ;
  LAYER M1 ;
        RECT 23.616 19.704 23.648 22.212 ;
  LAYER M1 ;
        RECT 23.68 19.704 23.712 22.212 ;
  LAYER M1 ;
        RECT 23.744 19.704 23.776 22.212 ;
  LAYER M1 ;
        RECT 23.808 19.704 23.84 22.212 ;
  LAYER M1 ;
        RECT 23.872 19.704 23.904 22.212 ;
  LAYER M1 ;
        RECT 23.936 19.704 23.968 22.212 ;
  LAYER M1 ;
        RECT 24 19.704 24.032 22.212 ;
  LAYER M1 ;
        RECT 24.064 19.704 24.096 22.212 ;
  LAYER M1 ;
        RECT 24.128 19.704 24.16 22.212 ;
  LAYER M2 ;
        RECT 21.804 22.096 24.276 22.128 ;
  LAYER M2 ;
        RECT 21.804 22.032 24.276 22.064 ;
  LAYER M2 ;
        RECT 21.804 21.968 24.276 22 ;
  LAYER M2 ;
        RECT 21.804 21.904 24.276 21.936 ;
  LAYER M2 ;
        RECT 21.804 21.84 24.276 21.872 ;
  LAYER M2 ;
        RECT 21.804 21.776 24.276 21.808 ;
  LAYER M2 ;
        RECT 21.804 21.712 24.276 21.744 ;
  LAYER M2 ;
        RECT 21.804 21.648 24.276 21.68 ;
  LAYER M2 ;
        RECT 21.804 21.584 24.276 21.616 ;
  LAYER M2 ;
        RECT 21.804 21.52 24.276 21.552 ;
  LAYER M2 ;
        RECT 21.804 21.456 24.276 21.488 ;
  LAYER M2 ;
        RECT 21.804 21.392 24.276 21.424 ;
  LAYER M2 ;
        RECT 21.804 21.328 24.276 21.36 ;
  LAYER M2 ;
        RECT 21.804 21.264 24.276 21.296 ;
  LAYER M2 ;
        RECT 21.804 21.2 24.276 21.232 ;
  LAYER M2 ;
        RECT 21.804 21.136 24.276 21.168 ;
  LAYER M2 ;
        RECT 21.804 21.072 24.276 21.104 ;
  LAYER M2 ;
        RECT 21.804 21.008 24.276 21.04 ;
  LAYER M2 ;
        RECT 21.804 20.944 24.276 20.976 ;
  LAYER M2 ;
        RECT 21.804 20.88 24.276 20.912 ;
  LAYER M2 ;
        RECT 21.804 20.816 24.276 20.848 ;
  LAYER M2 ;
        RECT 21.804 20.752 24.276 20.784 ;
  LAYER M2 ;
        RECT 21.804 20.688 24.276 20.72 ;
  LAYER M2 ;
        RECT 21.804 20.624 24.276 20.656 ;
  LAYER M2 ;
        RECT 21.804 20.56 24.276 20.592 ;
  LAYER M2 ;
        RECT 21.804 20.496 24.276 20.528 ;
  LAYER M2 ;
        RECT 21.804 20.432 24.276 20.464 ;
  LAYER M2 ;
        RECT 21.804 20.368 24.276 20.4 ;
  LAYER M2 ;
        RECT 21.804 20.304 24.276 20.336 ;
  LAYER M2 ;
        RECT 21.804 20.24 24.276 20.272 ;
  LAYER M2 ;
        RECT 21.804 20.176 24.276 20.208 ;
  LAYER M2 ;
        RECT 21.804 20.112 24.276 20.144 ;
  LAYER M2 ;
        RECT 21.804 20.048 24.276 20.08 ;
  LAYER M2 ;
        RECT 21.804 19.984 24.276 20.016 ;
  LAYER M2 ;
        RECT 21.804 19.92 24.276 19.952 ;
  LAYER M2 ;
        RECT 21.804 19.856 24.276 19.888 ;
  LAYER M3 ;
        RECT 21.824 19.704 21.856 22.212 ;
  LAYER M3 ;
        RECT 21.888 19.704 21.92 22.212 ;
  LAYER M3 ;
        RECT 21.952 19.704 21.984 22.212 ;
  LAYER M3 ;
        RECT 22.016 19.704 22.048 22.212 ;
  LAYER M3 ;
        RECT 22.08 19.704 22.112 22.212 ;
  LAYER M3 ;
        RECT 22.144 19.704 22.176 22.212 ;
  LAYER M3 ;
        RECT 22.208 19.704 22.24 22.212 ;
  LAYER M3 ;
        RECT 22.272 19.704 22.304 22.212 ;
  LAYER M3 ;
        RECT 22.336 19.704 22.368 22.212 ;
  LAYER M3 ;
        RECT 22.4 19.704 22.432 22.212 ;
  LAYER M3 ;
        RECT 22.464 19.704 22.496 22.212 ;
  LAYER M3 ;
        RECT 22.528 19.704 22.56 22.212 ;
  LAYER M3 ;
        RECT 22.592 19.704 22.624 22.212 ;
  LAYER M3 ;
        RECT 22.656 19.704 22.688 22.212 ;
  LAYER M3 ;
        RECT 22.72 19.704 22.752 22.212 ;
  LAYER M3 ;
        RECT 22.784 19.704 22.816 22.212 ;
  LAYER M3 ;
        RECT 22.848 19.704 22.88 22.212 ;
  LAYER M3 ;
        RECT 22.912 19.704 22.944 22.212 ;
  LAYER M3 ;
        RECT 22.976 19.704 23.008 22.212 ;
  LAYER M3 ;
        RECT 23.04 19.704 23.072 22.212 ;
  LAYER M3 ;
        RECT 23.104 19.704 23.136 22.212 ;
  LAYER M3 ;
        RECT 23.168 19.704 23.2 22.212 ;
  LAYER M3 ;
        RECT 23.232 19.704 23.264 22.212 ;
  LAYER M3 ;
        RECT 23.296 19.704 23.328 22.212 ;
  LAYER M3 ;
        RECT 23.36 19.704 23.392 22.212 ;
  LAYER M3 ;
        RECT 23.424 19.704 23.456 22.212 ;
  LAYER M3 ;
        RECT 23.488 19.704 23.52 22.212 ;
  LAYER M3 ;
        RECT 23.552 19.704 23.584 22.212 ;
  LAYER M3 ;
        RECT 23.616 19.704 23.648 22.212 ;
  LAYER M3 ;
        RECT 23.68 19.704 23.712 22.212 ;
  LAYER M3 ;
        RECT 23.744 19.704 23.776 22.212 ;
  LAYER M3 ;
        RECT 23.808 19.704 23.84 22.212 ;
  LAYER M3 ;
        RECT 23.872 19.704 23.904 22.212 ;
  LAYER M3 ;
        RECT 23.936 19.704 23.968 22.212 ;
  LAYER M3 ;
        RECT 24 19.704 24.032 22.212 ;
  LAYER M3 ;
        RECT 24.064 19.704 24.096 22.212 ;
  LAYER M3 ;
        RECT 24.128 19.704 24.16 22.212 ;
  LAYER M3 ;
        RECT 24.224 19.704 24.256 22.212 ;
  LAYER M1 ;
        RECT 21.839 19.74 21.841 22.176 ;
  LAYER M1 ;
        RECT 21.919 19.74 21.921 22.176 ;
  LAYER M1 ;
        RECT 21.999 19.74 22.001 22.176 ;
  LAYER M1 ;
        RECT 22.079 19.74 22.081 22.176 ;
  LAYER M1 ;
        RECT 22.159 19.74 22.161 22.176 ;
  LAYER M1 ;
        RECT 22.239 19.74 22.241 22.176 ;
  LAYER M1 ;
        RECT 22.319 19.74 22.321 22.176 ;
  LAYER M1 ;
        RECT 22.399 19.74 22.401 22.176 ;
  LAYER M1 ;
        RECT 22.479 19.74 22.481 22.176 ;
  LAYER M1 ;
        RECT 22.559 19.74 22.561 22.176 ;
  LAYER M1 ;
        RECT 22.639 19.74 22.641 22.176 ;
  LAYER M1 ;
        RECT 22.719 19.74 22.721 22.176 ;
  LAYER M1 ;
        RECT 22.799 19.74 22.801 22.176 ;
  LAYER M1 ;
        RECT 22.879 19.74 22.881 22.176 ;
  LAYER M1 ;
        RECT 22.959 19.74 22.961 22.176 ;
  LAYER M1 ;
        RECT 23.039 19.74 23.041 22.176 ;
  LAYER M1 ;
        RECT 23.119 19.74 23.121 22.176 ;
  LAYER M1 ;
        RECT 23.199 19.74 23.201 22.176 ;
  LAYER M1 ;
        RECT 23.279 19.74 23.281 22.176 ;
  LAYER M1 ;
        RECT 23.359 19.74 23.361 22.176 ;
  LAYER M1 ;
        RECT 23.439 19.74 23.441 22.176 ;
  LAYER M1 ;
        RECT 23.519 19.74 23.521 22.176 ;
  LAYER M1 ;
        RECT 23.599 19.74 23.601 22.176 ;
  LAYER M1 ;
        RECT 23.679 19.74 23.681 22.176 ;
  LAYER M1 ;
        RECT 23.759 19.74 23.761 22.176 ;
  LAYER M1 ;
        RECT 23.839 19.74 23.841 22.176 ;
  LAYER M1 ;
        RECT 23.919 19.74 23.921 22.176 ;
  LAYER M1 ;
        RECT 23.999 19.74 24.001 22.176 ;
  LAYER M1 ;
        RECT 24.079 19.74 24.081 22.176 ;
  LAYER M1 ;
        RECT 24.159 19.74 24.161 22.176 ;
  LAYER M2 ;
        RECT 21.84 22.175 24.24 22.177 ;
  LAYER M2 ;
        RECT 21.84 22.091 24.24 22.093 ;
  LAYER M2 ;
        RECT 21.84 22.007 24.24 22.009 ;
  LAYER M2 ;
        RECT 21.84 21.923 24.24 21.925 ;
  LAYER M2 ;
        RECT 21.84 21.839 24.24 21.841 ;
  LAYER M2 ;
        RECT 21.84 21.755 24.24 21.757 ;
  LAYER M2 ;
        RECT 21.84 21.671 24.24 21.673 ;
  LAYER M2 ;
        RECT 21.84 21.587 24.24 21.589 ;
  LAYER M2 ;
        RECT 21.84 21.503 24.24 21.505 ;
  LAYER M2 ;
        RECT 21.84 21.419 24.24 21.421 ;
  LAYER M2 ;
        RECT 21.84 21.335 24.24 21.337 ;
  LAYER M2 ;
        RECT 21.84 21.251 24.24 21.253 ;
  LAYER M2 ;
        RECT 21.84 21.1675 24.24 21.1695 ;
  LAYER M2 ;
        RECT 21.84 21.083 24.24 21.085 ;
  LAYER M2 ;
        RECT 21.84 20.999 24.24 21.001 ;
  LAYER M2 ;
        RECT 21.84 20.915 24.24 20.917 ;
  LAYER M2 ;
        RECT 21.84 20.831 24.24 20.833 ;
  LAYER M2 ;
        RECT 21.84 20.747 24.24 20.749 ;
  LAYER M2 ;
        RECT 21.84 20.663 24.24 20.665 ;
  LAYER M2 ;
        RECT 21.84 20.579 24.24 20.581 ;
  LAYER M2 ;
        RECT 21.84 20.495 24.24 20.497 ;
  LAYER M2 ;
        RECT 21.84 20.411 24.24 20.413 ;
  LAYER M2 ;
        RECT 21.84 20.327 24.24 20.329 ;
  LAYER M2 ;
        RECT 21.84 20.243 24.24 20.245 ;
  LAYER M2 ;
        RECT 21.84 20.159 24.24 20.161 ;
  LAYER M2 ;
        RECT 21.84 20.075 24.24 20.077 ;
  LAYER M2 ;
        RECT 21.84 19.991 24.24 19.993 ;
  LAYER M2 ;
        RECT 21.84 19.907 24.24 19.909 ;
  LAYER M2 ;
        RECT 21.84 19.823 24.24 19.825 ;
  LAYER M1 ;
        RECT 24.704 34.404 24.736 36.912 ;
  LAYER M1 ;
        RECT 24.768 34.404 24.8 36.912 ;
  LAYER M1 ;
        RECT 24.832 34.404 24.864 36.912 ;
  LAYER M1 ;
        RECT 24.896 34.404 24.928 36.912 ;
  LAYER M1 ;
        RECT 24.96 34.404 24.992 36.912 ;
  LAYER M1 ;
        RECT 25.024 34.404 25.056 36.912 ;
  LAYER M1 ;
        RECT 25.088 34.404 25.12 36.912 ;
  LAYER M1 ;
        RECT 25.152 34.404 25.184 36.912 ;
  LAYER M1 ;
        RECT 25.216 34.404 25.248 36.912 ;
  LAYER M1 ;
        RECT 25.28 34.404 25.312 36.912 ;
  LAYER M1 ;
        RECT 25.344 34.404 25.376 36.912 ;
  LAYER M1 ;
        RECT 25.408 34.404 25.44 36.912 ;
  LAYER M1 ;
        RECT 25.472 34.404 25.504 36.912 ;
  LAYER M1 ;
        RECT 25.536 34.404 25.568 36.912 ;
  LAYER M1 ;
        RECT 25.6 34.404 25.632 36.912 ;
  LAYER M1 ;
        RECT 25.664 34.404 25.696 36.912 ;
  LAYER M1 ;
        RECT 25.728 34.404 25.76 36.912 ;
  LAYER M1 ;
        RECT 25.792 34.404 25.824 36.912 ;
  LAYER M1 ;
        RECT 25.856 34.404 25.888 36.912 ;
  LAYER M1 ;
        RECT 25.92 34.404 25.952 36.912 ;
  LAYER M1 ;
        RECT 25.984 34.404 26.016 36.912 ;
  LAYER M1 ;
        RECT 26.048 34.404 26.08 36.912 ;
  LAYER M1 ;
        RECT 26.112 34.404 26.144 36.912 ;
  LAYER M1 ;
        RECT 26.176 34.404 26.208 36.912 ;
  LAYER M1 ;
        RECT 26.24 34.404 26.272 36.912 ;
  LAYER M1 ;
        RECT 26.304 34.404 26.336 36.912 ;
  LAYER M1 ;
        RECT 26.368 34.404 26.4 36.912 ;
  LAYER M1 ;
        RECT 26.432 34.404 26.464 36.912 ;
  LAYER M1 ;
        RECT 26.496 34.404 26.528 36.912 ;
  LAYER M1 ;
        RECT 26.56 34.404 26.592 36.912 ;
  LAYER M1 ;
        RECT 26.624 34.404 26.656 36.912 ;
  LAYER M1 ;
        RECT 26.688 34.404 26.72 36.912 ;
  LAYER M1 ;
        RECT 26.752 34.404 26.784 36.912 ;
  LAYER M1 ;
        RECT 26.816 34.404 26.848 36.912 ;
  LAYER M1 ;
        RECT 26.88 34.404 26.912 36.912 ;
  LAYER M1 ;
        RECT 26.944 34.404 26.976 36.912 ;
  LAYER M1 ;
        RECT 27.008 34.404 27.04 36.912 ;
  LAYER M2 ;
        RECT 24.684 36.796 27.156 36.828 ;
  LAYER M2 ;
        RECT 24.684 36.732 27.156 36.764 ;
  LAYER M2 ;
        RECT 24.684 36.668 27.156 36.7 ;
  LAYER M2 ;
        RECT 24.684 36.604 27.156 36.636 ;
  LAYER M2 ;
        RECT 24.684 36.54 27.156 36.572 ;
  LAYER M2 ;
        RECT 24.684 36.476 27.156 36.508 ;
  LAYER M2 ;
        RECT 24.684 36.412 27.156 36.444 ;
  LAYER M2 ;
        RECT 24.684 36.348 27.156 36.38 ;
  LAYER M2 ;
        RECT 24.684 36.284 27.156 36.316 ;
  LAYER M2 ;
        RECT 24.684 36.22 27.156 36.252 ;
  LAYER M2 ;
        RECT 24.684 36.156 27.156 36.188 ;
  LAYER M2 ;
        RECT 24.684 36.092 27.156 36.124 ;
  LAYER M2 ;
        RECT 24.684 36.028 27.156 36.06 ;
  LAYER M2 ;
        RECT 24.684 35.964 27.156 35.996 ;
  LAYER M2 ;
        RECT 24.684 35.9 27.156 35.932 ;
  LAYER M2 ;
        RECT 24.684 35.836 27.156 35.868 ;
  LAYER M2 ;
        RECT 24.684 35.772 27.156 35.804 ;
  LAYER M2 ;
        RECT 24.684 35.708 27.156 35.74 ;
  LAYER M2 ;
        RECT 24.684 35.644 27.156 35.676 ;
  LAYER M2 ;
        RECT 24.684 35.58 27.156 35.612 ;
  LAYER M2 ;
        RECT 24.684 35.516 27.156 35.548 ;
  LAYER M2 ;
        RECT 24.684 35.452 27.156 35.484 ;
  LAYER M2 ;
        RECT 24.684 35.388 27.156 35.42 ;
  LAYER M2 ;
        RECT 24.684 35.324 27.156 35.356 ;
  LAYER M2 ;
        RECT 24.684 35.26 27.156 35.292 ;
  LAYER M2 ;
        RECT 24.684 35.196 27.156 35.228 ;
  LAYER M2 ;
        RECT 24.684 35.132 27.156 35.164 ;
  LAYER M2 ;
        RECT 24.684 35.068 27.156 35.1 ;
  LAYER M2 ;
        RECT 24.684 35.004 27.156 35.036 ;
  LAYER M2 ;
        RECT 24.684 34.94 27.156 34.972 ;
  LAYER M2 ;
        RECT 24.684 34.876 27.156 34.908 ;
  LAYER M2 ;
        RECT 24.684 34.812 27.156 34.844 ;
  LAYER M2 ;
        RECT 24.684 34.748 27.156 34.78 ;
  LAYER M2 ;
        RECT 24.684 34.684 27.156 34.716 ;
  LAYER M2 ;
        RECT 24.684 34.62 27.156 34.652 ;
  LAYER M2 ;
        RECT 24.684 34.556 27.156 34.588 ;
  LAYER M3 ;
        RECT 24.704 34.404 24.736 36.912 ;
  LAYER M3 ;
        RECT 24.768 34.404 24.8 36.912 ;
  LAYER M3 ;
        RECT 24.832 34.404 24.864 36.912 ;
  LAYER M3 ;
        RECT 24.896 34.404 24.928 36.912 ;
  LAYER M3 ;
        RECT 24.96 34.404 24.992 36.912 ;
  LAYER M3 ;
        RECT 25.024 34.404 25.056 36.912 ;
  LAYER M3 ;
        RECT 25.088 34.404 25.12 36.912 ;
  LAYER M3 ;
        RECT 25.152 34.404 25.184 36.912 ;
  LAYER M3 ;
        RECT 25.216 34.404 25.248 36.912 ;
  LAYER M3 ;
        RECT 25.28 34.404 25.312 36.912 ;
  LAYER M3 ;
        RECT 25.344 34.404 25.376 36.912 ;
  LAYER M3 ;
        RECT 25.408 34.404 25.44 36.912 ;
  LAYER M3 ;
        RECT 25.472 34.404 25.504 36.912 ;
  LAYER M3 ;
        RECT 25.536 34.404 25.568 36.912 ;
  LAYER M3 ;
        RECT 25.6 34.404 25.632 36.912 ;
  LAYER M3 ;
        RECT 25.664 34.404 25.696 36.912 ;
  LAYER M3 ;
        RECT 25.728 34.404 25.76 36.912 ;
  LAYER M3 ;
        RECT 25.792 34.404 25.824 36.912 ;
  LAYER M3 ;
        RECT 25.856 34.404 25.888 36.912 ;
  LAYER M3 ;
        RECT 25.92 34.404 25.952 36.912 ;
  LAYER M3 ;
        RECT 25.984 34.404 26.016 36.912 ;
  LAYER M3 ;
        RECT 26.048 34.404 26.08 36.912 ;
  LAYER M3 ;
        RECT 26.112 34.404 26.144 36.912 ;
  LAYER M3 ;
        RECT 26.176 34.404 26.208 36.912 ;
  LAYER M3 ;
        RECT 26.24 34.404 26.272 36.912 ;
  LAYER M3 ;
        RECT 26.304 34.404 26.336 36.912 ;
  LAYER M3 ;
        RECT 26.368 34.404 26.4 36.912 ;
  LAYER M3 ;
        RECT 26.432 34.404 26.464 36.912 ;
  LAYER M3 ;
        RECT 26.496 34.404 26.528 36.912 ;
  LAYER M3 ;
        RECT 26.56 34.404 26.592 36.912 ;
  LAYER M3 ;
        RECT 26.624 34.404 26.656 36.912 ;
  LAYER M3 ;
        RECT 26.688 34.404 26.72 36.912 ;
  LAYER M3 ;
        RECT 26.752 34.404 26.784 36.912 ;
  LAYER M3 ;
        RECT 26.816 34.404 26.848 36.912 ;
  LAYER M3 ;
        RECT 26.88 34.404 26.912 36.912 ;
  LAYER M3 ;
        RECT 26.944 34.404 26.976 36.912 ;
  LAYER M3 ;
        RECT 27.008 34.404 27.04 36.912 ;
  LAYER M3 ;
        RECT 27.104 34.404 27.136 36.912 ;
  LAYER M1 ;
        RECT 24.719 34.44 24.721 36.876 ;
  LAYER M1 ;
        RECT 24.799 34.44 24.801 36.876 ;
  LAYER M1 ;
        RECT 24.879 34.44 24.881 36.876 ;
  LAYER M1 ;
        RECT 24.959 34.44 24.961 36.876 ;
  LAYER M1 ;
        RECT 25.039 34.44 25.041 36.876 ;
  LAYER M1 ;
        RECT 25.119 34.44 25.121 36.876 ;
  LAYER M1 ;
        RECT 25.199 34.44 25.201 36.876 ;
  LAYER M1 ;
        RECT 25.279 34.44 25.281 36.876 ;
  LAYER M1 ;
        RECT 25.359 34.44 25.361 36.876 ;
  LAYER M1 ;
        RECT 25.439 34.44 25.441 36.876 ;
  LAYER M1 ;
        RECT 25.519 34.44 25.521 36.876 ;
  LAYER M1 ;
        RECT 25.599 34.44 25.601 36.876 ;
  LAYER M1 ;
        RECT 25.679 34.44 25.681 36.876 ;
  LAYER M1 ;
        RECT 25.759 34.44 25.761 36.876 ;
  LAYER M1 ;
        RECT 25.839 34.44 25.841 36.876 ;
  LAYER M1 ;
        RECT 25.919 34.44 25.921 36.876 ;
  LAYER M1 ;
        RECT 25.999 34.44 26.001 36.876 ;
  LAYER M1 ;
        RECT 26.079 34.44 26.081 36.876 ;
  LAYER M1 ;
        RECT 26.159 34.44 26.161 36.876 ;
  LAYER M1 ;
        RECT 26.239 34.44 26.241 36.876 ;
  LAYER M1 ;
        RECT 26.319 34.44 26.321 36.876 ;
  LAYER M1 ;
        RECT 26.399 34.44 26.401 36.876 ;
  LAYER M1 ;
        RECT 26.479 34.44 26.481 36.876 ;
  LAYER M1 ;
        RECT 26.559 34.44 26.561 36.876 ;
  LAYER M1 ;
        RECT 26.639 34.44 26.641 36.876 ;
  LAYER M1 ;
        RECT 26.719 34.44 26.721 36.876 ;
  LAYER M1 ;
        RECT 26.799 34.44 26.801 36.876 ;
  LAYER M1 ;
        RECT 26.879 34.44 26.881 36.876 ;
  LAYER M1 ;
        RECT 26.959 34.44 26.961 36.876 ;
  LAYER M1 ;
        RECT 27.039 34.44 27.041 36.876 ;
  LAYER M2 ;
        RECT 24.72 36.875 27.12 36.877 ;
  LAYER M2 ;
        RECT 24.72 36.791 27.12 36.793 ;
  LAYER M2 ;
        RECT 24.72 36.707 27.12 36.709 ;
  LAYER M2 ;
        RECT 24.72 36.623 27.12 36.625 ;
  LAYER M2 ;
        RECT 24.72 36.539 27.12 36.541 ;
  LAYER M2 ;
        RECT 24.72 36.455 27.12 36.457 ;
  LAYER M2 ;
        RECT 24.72 36.371 27.12 36.373 ;
  LAYER M2 ;
        RECT 24.72 36.287 27.12 36.289 ;
  LAYER M2 ;
        RECT 24.72 36.203 27.12 36.205 ;
  LAYER M2 ;
        RECT 24.72 36.119 27.12 36.121 ;
  LAYER M2 ;
        RECT 24.72 36.035 27.12 36.037 ;
  LAYER M2 ;
        RECT 24.72 35.951 27.12 35.953 ;
  LAYER M2 ;
        RECT 24.72 35.8675 27.12 35.8695 ;
  LAYER M2 ;
        RECT 24.72 35.783 27.12 35.785 ;
  LAYER M2 ;
        RECT 24.72 35.699 27.12 35.701 ;
  LAYER M2 ;
        RECT 24.72 35.615 27.12 35.617 ;
  LAYER M2 ;
        RECT 24.72 35.531 27.12 35.533 ;
  LAYER M2 ;
        RECT 24.72 35.447 27.12 35.449 ;
  LAYER M2 ;
        RECT 24.72 35.363 27.12 35.365 ;
  LAYER M2 ;
        RECT 24.72 35.279 27.12 35.281 ;
  LAYER M2 ;
        RECT 24.72 35.195 27.12 35.197 ;
  LAYER M2 ;
        RECT 24.72 35.111 27.12 35.113 ;
  LAYER M2 ;
        RECT 24.72 35.027 27.12 35.029 ;
  LAYER M2 ;
        RECT 24.72 34.943 27.12 34.945 ;
  LAYER M2 ;
        RECT 24.72 34.859 27.12 34.861 ;
  LAYER M2 ;
        RECT 24.72 34.775 27.12 34.777 ;
  LAYER M2 ;
        RECT 24.72 34.691 27.12 34.693 ;
  LAYER M2 ;
        RECT 24.72 34.607 27.12 34.609 ;
  LAYER M2 ;
        RECT 24.72 34.523 27.12 34.525 ;
  LAYER M1 ;
        RECT 24.704 31.464 24.736 33.972 ;
  LAYER M1 ;
        RECT 24.768 31.464 24.8 33.972 ;
  LAYER M1 ;
        RECT 24.832 31.464 24.864 33.972 ;
  LAYER M1 ;
        RECT 24.896 31.464 24.928 33.972 ;
  LAYER M1 ;
        RECT 24.96 31.464 24.992 33.972 ;
  LAYER M1 ;
        RECT 25.024 31.464 25.056 33.972 ;
  LAYER M1 ;
        RECT 25.088 31.464 25.12 33.972 ;
  LAYER M1 ;
        RECT 25.152 31.464 25.184 33.972 ;
  LAYER M1 ;
        RECT 25.216 31.464 25.248 33.972 ;
  LAYER M1 ;
        RECT 25.28 31.464 25.312 33.972 ;
  LAYER M1 ;
        RECT 25.344 31.464 25.376 33.972 ;
  LAYER M1 ;
        RECT 25.408 31.464 25.44 33.972 ;
  LAYER M1 ;
        RECT 25.472 31.464 25.504 33.972 ;
  LAYER M1 ;
        RECT 25.536 31.464 25.568 33.972 ;
  LAYER M1 ;
        RECT 25.6 31.464 25.632 33.972 ;
  LAYER M1 ;
        RECT 25.664 31.464 25.696 33.972 ;
  LAYER M1 ;
        RECT 25.728 31.464 25.76 33.972 ;
  LAYER M1 ;
        RECT 25.792 31.464 25.824 33.972 ;
  LAYER M1 ;
        RECT 25.856 31.464 25.888 33.972 ;
  LAYER M1 ;
        RECT 25.92 31.464 25.952 33.972 ;
  LAYER M1 ;
        RECT 25.984 31.464 26.016 33.972 ;
  LAYER M1 ;
        RECT 26.048 31.464 26.08 33.972 ;
  LAYER M1 ;
        RECT 26.112 31.464 26.144 33.972 ;
  LAYER M1 ;
        RECT 26.176 31.464 26.208 33.972 ;
  LAYER M1 ;
        RECT 26.24 31.464 26.272 33.972 ;
  LAYER M1 ;
        RECT 26.304 31.464 26.336 33.972 ;
  LAYER M1 ;
        RECT 26.368 31.464 26.4 33.972 ;
  LAYER M1 ;
        RECT 26.432 31.464 26.464 33.972 ;
  LAYER M1 ;
        RECT 26.496 31.464 26.528 33.972 ;
  LAYER M1 ;
        RECT 26.56 31.464 26.592 33.972 ;
  LAYER M1 ;
        RECT 26.624 31.464 26.656 33.972 ;
  LAYER M1 ;
        RECT 26.688 31.464 26.72 33.972 ;
  LAYER M1 ;
        RECT 26.752 31.464 26.784 33.972 ;
  LAYER M1 ;
        RECT 26.816 31.464 26.848 33.972 ;
  LAYER M1 ;
        RECT 26.88 31.464 26.912 33.972 ;
  LAYER M1 ;
        RECT 26.944 31.464 26.976 33.972 ;
  LAYER M1 ;
        RECT 27.008 31.464 27.04 33.972 ;
  LAYER M2 ;
        RECT 24.684 33.856 27.156 33.888 ;
  LAYER M2 ;
        RECT 24.684 33.792 27.156 33.824 ;
  LAYER M2 ;
        RECT 24.684 33.728 27.156 33.76 ;
  LAYER M2 ;
        RECT 24.684 33.664 27.156 33.696 ;
  LAYER M2 ;
        RECT 24.684 33.6 27.156 33.632 ;
  LAYER M2 ;
        RECT 24.684 33.536 27.156 33.568 ;
  LAYER M2 ;
        RECT 24.684 33.472 27.156 33.504 ;
  LAYER M2 ;
        RECT 24.684 33.408 27.156 33.44 ;
  LAYER M2 ;
        RECT 24.684 33.344 27.156 33.376 ;
  LAYER M2 ;
        RECT 24.684 33.28 27.156 33.312 ;
  LAYER M2 ;
        RECT 24.684 33.216 27.156 33.248 ;
  LAYER M2 ;
        RECT 24.684 33.152 27.156 33.184 ;
  LAYER M2 ;
        RECT 24.684 33.088 27.156 33.12 ;
  LAYER M2 ;
        RECT 24.684 33.024 27.156 33.056 ;
  LAYER M2 ;
        RECT 24.684 32.96 27.156 32.992 ;
  LAYER M2 ;
        RECT 24.684 32.896 27.156 32.928 ;
  LAYER M2 ;
        RECT 24.684 32.832 27.156 32.864 ;
  LAYER M2 ;
        RECT 24.684 32.768 27.156 32.8 ;
  LAYER M2 ;
        RECT 24.684 32.704 27.156 32.736 ;
  LAYER M2 ;
        RECT 24.684 32.64 27.156 32.672 ;
  LAYER M2 ;
        RECT 24.684 32.576 27.156 32.608 ;
  LAYER M2 ;
        RECT 24.684 32.512 27.156 32.544 ;
  LAYER M2 ;
        RECT 24.684 32.448 27.156 32.48 ;
  LAYER M2 ;
        RECT 24.684 32.384 27.156 32.416 ;
  LAYER M2 ;
        RECT 24.684 32.32 27.156 32.352 ;
  LAYER M2 ;
        RECT 24.684 32.256 27.156 32.288 ;
  LAYER M2 ;
        RECT 24.684 32.192 27.156 32.224 ;
  LAYER M2 ;
        RECT 24.684 32.128 27.156 32.16 ;
  LAYER M2 ;
        RECT 24.684 32.064 27.156 32.096 ;
  LAYER M2 ;
        RECT 24.684 32 27.156 32.032 ;
  LAYER M2 ;
        RECT 24.684 31.936 27.156 31.968 ;
  LAYER M2 ;
        RECT 24.684 31.872 27.156 31.904 ;
  LAYER M2 ;
        RECT 24.684 31.808 27.156 31.84 ;
  LAYER M2 ;
        RECT 24.684 31.744 27.156 31.776 ;
  LAYER M2 ;
        RECT 24.684 31.68 27.156 31.712 ;
  LAYER M2 ;
        RECT 24.684 31.616 27.156 31.648 ;
  LAYER M3 ;
        RECT 24.704 31.464 24.736 33.972 ;
  LAYER M3 ;
        RECT 24.768 31.464 24.8 33.972 ;
  LAYER M3 ;
        RECT 24.832 31.464 24.864 33.972 ;
  LAYER M3 ;
        RECT 24.896 31.464 24.928 33.972 ;
  LAYER M3 ;
        RECT 24.96 31.464 24.992 33.972 ;
  LAYER M3 ;
        RECT 25.024 31.464 25.056 33.972 ;
  LAYER M3 ;
        RECT 25.088 31.464 25.12 33.972 ;
  LAYER M3 ;
        RECT 25.152 31.464 25.184 33.972 ;
  LAYER M3 ;
        RECT 25.216 31.464 25.248 33.972 ;
  LAYER M3 ;
        RECT 25.28 31.464 25.312 33.972 ;
  LAYER M3 ;
        RECT 25.344 31.464 25.376 33.972 ;
  LAYER M3 ;
        RECT 25.408 31.464 25.44 33.972 ;
  LAYER M3 ;
        RECT 25.472 31.464 25.504 33.972 ;
  LAYER M3 ;
        RECT 25.536 31.464 25.568 33.972 ;
  LAYER M3 ;
        RECT 25.6 31.464 25.632 33.972 ;
  LAYER M3 ;
        RECT 25.664 31.464 25.696 33.972 ;
  LAYER M3 ;
        RECT 25.728 31.464 25.76 33.972 ;
  LAYER M3 ;
        RECT 25.792 31.464 25.824 33.972 ;
  LAYER M3 ;
        RECT 25.856 31.464 25.888 33.972 ;
  LAYER M3 ;
        RECT 25.92 31.464 25.952 33.972 ;
  LAYER M3 ;
        RECT 25.984 31.464 26.016 33.972 ;
  LAYER M3 ;
        RECT 26.048 31.464 26.08 33.972 ;
  LAYER M3 ;
        RECT 26.112 31.464 26.144 33.972 ;
  LAYER M3 ;
        RECT 26.176 31.464 26.208 33.972 ;
  LAYER M3 ;
        RECT 26.24 31.464 26.272 33.972 ;
  LAYER M3 ;
        RECT 26.304 31.464 26.336 33.972 ;
  LAYER M3 ;
        RECT 26.368 31.464 26.4 33.972 ;
  LAYER M3 ;
        RECT 26.432 31.464 26.464 33.972 ;
  LAYER M3 ;
        RECT 26.496 31.464 26.528 33.972 ;
  LAYER M3 ;
        RECT 26.56 31.464 26.592 33.972 ;
  LAYER M3 ;
        RECT 26.624 31.464 26.656 33.972 ;
  LAYER M3 ;
        RECT 26.688 31.464 26.72 33.972 ;
  LAYER M3 ;
        RECT 26.752 31.464 26.784 33.972 ;
  LAYER M3 ;
        RECT 26.816 31.464 26.848 33.972 ;
  LAYER M3 ;
        RECT 26.88 31.464 26.912 33.972 ;
  LAYER M3 ;
        RECT 26.944 31.464 26.976 33.972 ;
  LAYER M3 ;
        RECT 27.008 31.464 27.04 33.972 ;
  LAYER M3 ;
        RECT 27.104 31.464 27.136 33.972 ;
  LAYER M1 ;
        RECT 24.719 31.5 24.721 33.936 ;
  LAYER M1 ;
        RECT 24.799 31.5 24.801 33.936 ;
  LAYER M1 ;
        RECT 24.879 31.5 24.881 33.936 ;
  LAYER M1 ;
        RECT 24.959 31.5 24.961 33.936 ;
  LAYER M1 ;
        RECT 25.039 31.5 25.041 33.936 ;
  LAYER M1 ;
        RECT 25.119 31.5 25.121 33.936 ;
  LAYER M1 ;
        RECT 25.199 31.5 25.201 33.936 ;
  LAYER M1 ;
        RECT 25.279 31.5 25.281 33.936 ;
  LAYER M1 ;
        RECT 25.359 31.5 25.361 33.936 ;
  LAYER M1 ;
        RECT 25.439 31.5 25.441 33.936 ;
  LAYER M1 ;
        RECT 25.519 31.5 25.521 33.936 ;
  LAYER M1 ;
        RECT 25.599 31.5 25.601 33.936 ;
  LAYER M1 ;
        RECT 25.679 31.5 25.681 33.936 ;
  LAYER M1 ;
        RECT 25.759 31.5 25.761 33.936 ;
  LAYER M1 ;
        RECT 25.839 31.5 25.841 33.936 ;
  LAYER M1 ;
        RECT 25.919 31.5 25.921 33.936 ;
  LAYER M1 ;
        RECT 25.999 31.5 26.001 33.936 ;
  LAYER M1 ;
        RECT 26.079 31.5 26.081 33.936 ;
  LAYER M1 ;
        RECT 26.159 31.5 26.161 33.936 ;
  LAYER M1 ;
        RECT 26.239 31.5 26.241 33.936 ;
  LAYER M1 ;
        RECT 26.319 31.5 26.321 33.936 ;
  LAYER M1 ;
        RECT 26.399 31.5 26.401 33.936 ;
  LAYER M1 ;
        RECT 26.479 31.5 26.481 33.936 ;
  LAYER M1 ;
        RECT 26.559 31.5 26.561 33.936 ;
  LAYER M1 ;
        RECT 26.639 31.5 26.641 33.936 ;
  LAYER M1 ;
        RECT 26.719 31.5 26.721 33.936 ;
  LAYER M1 ;
        RECT 26.799 31.5 26.801 33.936 ;
  LAYER M1 ;
        RECT 26.879 31.5 26.881 33.936 ;
  LAYER M1 ;
        RECT 26.959 31.5 26.961 33.936 ;
  LAYER M1 ;
        RECT 27.039 31.5 27.041 33.936 ;
  LAYER M2 ;
        RECT 24.72 33.935 27.12 33.937 ;
  LAYER M2 ;
        RECT 24.72 33.851 27.12 33.853 ;
  LAYER M2 ;
        RECT 24.72 33.767 27.12 33.769 ;
  LAYER M2 ;
        RECT 24.72 33.683 27.12 33.685 ;
  LAYER M2 ;
        RECT 24.72 33.599 27.12 33.601 ;
  LAYER M2 ;
        RECT 24.72 33.515 27.12 33.517 ;
  LAYER M2 ;
        RECT 24.72 33.431 27.12 33.433 ;
  LAYER M2 ;
        RECT 24.72 33.347 27.12 33.349 ;
  LAYER M2 ;
        RECT 24.72 33.263 27.12 33.265 ;
  LAYER M2 ;
        RECT 24.72 33.179 27.12 33.181 ;
  LAYER M2 ;
        RECT 24.72 33.095 27.12 33.097 ;
  LAYER M2 ;
        RECT 24.72 33.011 27.12 33.013 ;
  LAYER M2 ;
        RECT 24.72 32.9275 27.12 32.9295 ;
  LAYER M2 ;
        RECT 24.72 32.843 27.12 32.845 ;
  LAYER M2 ;
        RECT 24.72 32.759 27.12 32.761 ;
  LAYER M2 ;
        RECT 24.72 32.675 27.12 32.677 ;
  LAYER M2 ;
        RECT 24.72 32.591 27.12 32.593 ;
  LAYER M2 ;
        RECT 24.72 32.507 27.12 32.509 ;
  LAYER M2 ;
        RECT 24.72 32.423 27.12 32.425 ;
  LAYER M2 ;
        RECT 24.72 32.339 27.12 32.341 ;
  LAYER M2 ;
        RECT 24.72 32.255 27.12 32.257 ;
  LAYER M2 ;
        RECT 24.72 32.171 27.12 32.173 ;
  LAYER M2 ;
        RECT 24.72 32.087 27.12 32.089 ;
  LAYER M2 ;
        RECT 24.72 32.003 27.12 32.005 ;
  LAYER M2 ;
        RECT 24.72 31.919 27.12 31.921 ;
  LAYER M2 ;
        RECT 24.72 31.835 27.12 31.837 ;
  LAYER M2 ;
        RECT 24.72 31.751 27.12 31.753 ;
  LAYER M2 ;
        RECT 24.72 31.667 27.12 31.669 ;
  LAYER M2 ;
        RECT 24.72 31.583 27.12 31.585 ;
  LAYER M1 ;
        RECT 24.704 28.524 24.736 31.032 ;
  LAYER M1 ;
        RECT 24.768 28.524 24.8 31.032 ;
  LAYER M1 ;
        RECT 24.832 28.524 24.864 31.032 ;
  LAYER M1 ;
        RECT 24.896 28.524 24.928 31.032 ;
  LAYER M1 ;
        RECT 24.96 28.524 24.992 31.032 ;
  LAYER M1 ;
        RECT 25.024 28.524 25.056 31.032 ;
  LAYER M1 ;
        RECT 25.088 28.524 25.12 31.032 ;
  LAYER M1 ;
        RECT 25.152 28.524 25.184 31.032 ;
  LAYER M1 ;
        RECT 25.216 28.524 25.248 31.032 ;
  LAYER M1 ;
        RECT 25.28 28.524 25.312 31.032 ;
  LAYER M1 ;
        RECT 25.344 28.524 25.376 31.032 ;
  LAYER M1 ;
        RECT 25.408 28.524 25.44 31.032 ;
  LAYER M1 ;
        RECT 25.472 28.524 25.504 31.032 ;
  LAYER M1 ;
        RECT 25.536 28.524 25.568 31.032 ;
  LAYER M1 ;
        RECT 25.6 28.524 25.632 31.032 ;
  LAYER M1 ;
        RECT 25.664 28.524 25.696 31.032 ;
  LAYER M1 ;
        RECT 25.728 28.524 25.76 31.032 ;
  LAYER M1 ;
        RECT 25.792 28.524 25.824 31.032 ;
  LAYER M1 ;
        RECT 25.856 28.524 25.888 31.032 ;
  LAYER M1 ;
        RECT 25.92 28.524 25.952 31.032 ;
  LAYER M1 ;
        RECT 25.984 28.524 26.016 31.032 ;
  LAYER M1 ;
        RECT 26.048 28.524 26.08 31.032 ;
  LAYER M1 ;
        RECT 26.112 28.524 26.144 31.032 ;
  LAYER M1 ;
        RECT 26.176 28.524 26.208 31.032 ;
  LAYER M1 ;
        RECT 26.24 28.524 26.272 31.032 ;
  LAYER M1 ;
        RECT 26.304 28.524 26.336 31.032 ;
  LAYER M1 ;
        RECT 26.368 28.524 26.4 31.032 ;
  LAYER M1 ;
        RECT 26.432 28.524 26.464 31.032 ;
  LAYER M1 ;
        RECT 26.496 28.524 26.528 31.032 ;
  LAYER M1 ;
        RECT 26.56 28.524 26.592 31.032 ;
  LAYER M1 ;
        RECT 26.624 28.524 26.656 31.032 ;
  LAYER M1 ;
        RECT 26.688 28.524 26.72 31.032 ;
  LAYER M1 ;
        RECT 26.752 28.524 26.784 31.032 ;
  LAYER M1 ;
        RECT 26.816 28.524 26.848 31.032 ;
  LAYER M1 ;
        RECT 26.88 28.524 26.912 31.032 ;
  LAYER M1 ;
        RECT 26.944 28.524 26.976 31.032 ;
  LAYER M1 ;
        RECT 27.008 28.524 27.04 31.032 ;
  LAYER M2 ;
        RECT 24.684 30.916 27.156 30.948 ;
  LAYER M2 ;
        RECT 24.684 30.852 27.156 30.884 ;
  LAYER M2 ;
        RECT 24.684 30.788 27.156 30.82 ;
  LAYER M2 ;
        RECT 24.684 30.724 27.156 30.756 ;
  LAYER M2 ;
        RECT 24.684 30.66 27.156 30.692 ;
  LAYER M2 ;
        RECT 24.684 30.596 27.156 30.628 ;
  LAYER M2 ;
        RECT 24.684 30.532 27.156 30.564 ;
  LAYER M2 ;
        RECT 24.684 30.468 27.156 30.5 ;
  LAYER M2 ;
        RECT 24.684 30.404 27.156 30.436 ;
  LAYER M2 ;
        RECT 24.684 30.34 27.156 30.372 ;
  LAYER M2 ;
        RECT 24.684 30.276 27.156 30.308 ;
  LAYER M2 ;
        RECT 24.684 30.212 27.156 30.244 ;
  LAYER M2 ;
        RECT 24.684 30.148 27.156 30.18 ;
  LAYER M2 ;
        RECT 24.684 30.084 27.156 30.116 ;
  LAYER M2 ;
        RECT 24.684 30.02 27.156 30.052 ;
  LAYER M2 ;
        RECT 24.684 29.956 27.156 29.988 ;
  LAYER M2 ;
        RECT 24.684 29.892 27.156 29.924 ;
  LAYER M2 ;
        RECT 24.684 29.828 27.156 29.86 ;
  LAYER M2 ;
        RECT 24.684 29.764 27.156 29.796 ;
  LAYER M2 ;
        RECT 24.684 29.7 27.156 29.732 ;
  LAYER M2 ;
        RECT 24.684 29.636 27.156 29.668 ;
  LAYER M2 ;
        RECT 24.684 29.572 27.156 29.604 ;
  LAYER M2 ;
        RECT 24.684 29.508 27.156 29.54 ;
  LAYER M2 ;
        RECT 24.684 29.444 27.156 29.476 ;
  LAYER M2 ;
        RECT 24.684 29.38 27.156 29.412 ;
  LAYER M2 ;
        RECT 24.684 29.316 27.156 29.348 ;
  LAYER M2 ;
        RECT 24.684 29.252 27.156 29.284 ;
  LAYER M2 ;
        RECT 24.684 29.188 27.156 29.22 ;
  LAYER M2 ;
        RECT 24.684 29.124 27.156 29.156 ;
  LAYER M2 ;
        RECT 24.684 29.06 27.156 29.092 ;
  LAYER M2 ;
        RECT 24.684 28.996 27.156 29.028 ;
  LAYER M2 ;
        RECT 24.684 28.932 27.156 28.964 ;
  LAYER M2 ;
        RECT 24.684 28.868 27.156 28.9 ;
  LAYER M2 ;
        RECT 24.684 28.804 27.156 28.836 ;
  LAYER M2 ;
        RECT 24.684 28.74 27.156 28.772 ;
  LAYER M2 ;
        RECT 24.684 28.676 27.156 28.708 ;
  LAYER M3 ;
        RECT 24.704 28.524 24.736 31.032 ;
  LAYER M3 ;
        RECT 24.768 28.524 24.8 31.032 ;
  LAYER M3 ;
        RECT 24.832 28.524 24.864 31.032 ;
  LAYER M3 ;
        RECT 24.896 28.524 24.928 31.032 ;
  LAYER M3 ;
        RECT 24.96 28.524 24.992 31.032 ;
  LAYER M3 ;
        RECT 25.024 28.524 25.056 31.032 ;
  LAYER M3 ;
        RECT 25.088 28.524 25.12 31.032 ;
  LAYER M3 ;
        RECT 25.152 28.524 25.184 31.032 ;
  LAYER M3 ;
        RECT 25.216 28.524 25.248 31.032 ;
  LAYER M3 ;
        RECT 25.28 28.524 25.312 31.032 ;
  LAYER M3 ;
        RECT 25.344 28.524 25.376 31.032 ;
  LAYER M3 ;
        RECT 25.408 28.524 25.44 31.032 ;
  LAYER M3 ;
        RECT 25.472 28.524 25.504 31.032 ;
  LAYER M3 ;
        RECT 25.536 28.524 25.568 31.032 ;
  LAYER M3 ;
        RECT 25.6 28.524 25.632 31.032 ;
  LAYER M3 ;
        RECT 25.664 28.524 25.696 31.032 ;
  LAYER M3 ;
        RECT 25.728 28.524 25.76 31.032 ;
  LAYER M3 ;
        RECT 25.792 28.524 25.824 31.032 ;
  LAYER M3 ;
        RECT 25.856 28.524 25.888 31.032 ;
  LAYER M3 ;
        RECT 25.92 28.524 25.952 31.032 ;
  LAYER M3 ;
        RECT 25.984 28.524 26.016 31.032 ;
  LAYER M3 ;
        RECT 26.048 28.524 26.08 31.032 ;
  LAYER M3 ;
        RECT 26.112 28.524 26.144 31.032 ;
  LAYER M3 ;
        RECT 26.176 28.524 26.208 31.032 ;
  LAYER M3 ;
        RECT 26.24 28.524 26.272 31.032 ;
  LAYER M3 ;
        RECT 26.304 28.524 26.336 31.032 ;
  LAYER M3 ;
        RECT 26.368 28.524 26.4 31.032 ;
  LAYER M3 ;
        RECT 26.432 28.524 26.464 31.032 ;
  LAYER M3 ;
        RECT 26.496 28.524 26.528 31.032 ;
  LAYER M3 ;
        RECT 26.56 28.524 26.592 31.032 ;
  LAYER M3 ;
        RECT 26.624 28.524 26.656 31.032 ;
  LAYER M3 ;
        RECT 26.688 28.524 26.72 31.032 ;
  LAYER M3 ;
        RECT 26.752 28.524 26.784 31.032 ;
  LAYER M3 ;
        RECT 26.816 28.524 26.848 31.032 ;
  LAYER M3 ;
        RECT 26.88 28.524 26.912 31.032 ;
  LAYER M3 ;
        RECT 26.944 28.524 26.976 31.032 ;
  LAYER M3 ;
        RECT 27.008 28.524 27.04 31.032 ;
  LAYER M3 ;
        RECT 27.104 28.524 27.136 31.032 ;
  LAYER M1 ;
        RECT 24.719 28.56 24.721 30.996 ;
  LAYER M1 ;
        RECT 24.799 28.56 24.801 30.996 ;
  LAYER M1 ;
        RECT 24.879 28.56 24.881 30.996 ;
  LAYER M1 ;
        RECT 24.959 28.56 24.961 30.996 ;
  LAYER M1 ;
        RECT 25.039 28.56 25.041 30.996 ;
  LAYER M1 ;
        RECT 25.119 28.56 25.121 30.996 ;
  LAYER M1 ;
        RECT 25.199 28.56 25.201 30.996 ;
  LAYER M1 ;
        RECT 25.279 28.56 25.281 30.996 ;
  LAYER M1 ;
        RECT 25.359 28.56 25.361 30.996 ;
  LAYER M1 ;
        RECT 25.439 28.56 25.441 30.996 ;
  LAYER M1 ;
        RECT 25.519 28.56 25.521 30.996 ;
  LAYER M1 ;
        RECT 25.599 28.56 25.601 30.996 ;
  LAYER M1 ;
        RECT 25.679 28.56 25.681 30.996 ;
  LAYER M1 ;
        RECT 25.759 28.56 25.761 30.996 ;
  LAYER M1 ;
        RECT 25.839 28.56 25.841 30.996 ;
  LAYER M1 ;
        RECT 25.919 28.56 25.921 30.996 ;
  LAYER M1 ;
        RECT 25.999 28.56 26.001 30.996 ;
  LAYER M1 ;
        RECT 26.079 28.56 26.081 30.996 ;
  LAYER M1 ;
        RECT 26.159 28.56 26.161 30.996 ;
  LAYER M1 ;
        RECT 26.239 28.56 26.241 30.996 ;
  LAYER M1 ;
        RECT 26.319 28.56 26.321 30.996 ;
  LAYER M1 ;
        RECT 26.399 28.56 26.401 30.996 ;
  LAYER M1 ;
        RECT 26.479 28.56 26.481 30.996 ;
  LAYER M1 ;
        RECT 26.559 28.56 26.561 30.996 ;
  LAYER M1 ;
        RECT 26.639 28.56 26.641 30.996 ;
  LAYER M1 ;
        RECT 26.719 28.56 26.721 30.996 ;
  LAYER M1 ;
        RECT 26.799 28.56 26.801 30.996 ;
  LAYER M1 ;
        RECT 26.879 28.56 26.881 30.996 ;
  LAYER M1 ;
        RECT 26.959 28.56 26.961 30.996 ;
  LAYER M1 ;
        RECT 27.039 28.56 27.041 30.996 ;
  LAYER M2 ;
        RECT 24.72 30.995 27.12 30.997 ;
  LAYER M2 ;
        RECT 24.72 30.911 27.12 30.913 ;
  LAYER M2 ;
        RECT 24.72 30.827 27.12 30.829 ;
  LAYER M2 ;
        RECT 24.72 30.743 27.12 30.745 ;
  LAYER M2 ;
        RECT 24.72 30.659 27.12 30.661 ;
  LAYER M2 ;
        RECT 24.72 30.575 27.12 30.577 ;
  LAYER M2 ;
        RECT 24.72 30.491 27.12 30.493 ;
  LAYER M2 ;
        RECT 24.72 30.407 27.12 30.409 ;
  LAYER M2 ;
        RECT 24.72 30.323 27.12 30.325 ;
  LAYER M2 ;
        RECT 24.72 30.239 27.12 30.241 ;
  LAYER M2 ;
        RECT 24.72 30.155 27.12 30.157 ;
  LAYER M2 ;
        RECT 24.72 30.071 27.12 30.073 ;
  LAYER M2 ;
        RECT 24.72 29.9875 27.12 29.9895 ;
  LAYER M2 ;
        RECT 24.72 29.903 27.12 29.905 ;
  LAYER M2 ;
        RECT 24.72 29.819 27.12 29.821 ;
  LAYER M2 ;
        RECT 24.72 29.735 27.12 29.737 ;
  LAYER M2 ;
        RECT 24.72 29.651 27.12 29.653 ;
  LAYER M2 ;
        RECT 24.72 29.567 27.12 29.569 ;
  LAYER M2 ;
        RECT 24.72 29.483 27.12 29.485 ;
  LAYER M2 ;
        RECT 24.72 29.399 27.12 29.401 ;
  LAYER M2 ;
        RECT 24.72 29.315 27.12 29.317 ;
  LAYER M2 ;
        RECT 24.72 29.231 27.12 29.233 ;
  LAYER M2 ;
        RECT 24.72 29.147 27.12 29.149 ;
  LAYER M2 ;
        RECT 24.72 29.063 27.12 29.065 ;
  LAYER M2 ;
        RECT 24.72 28.979 27.12 28.981 ;
  LAYER M2 ;
        RECT 24.72 28.895 27.12 28.897 ;
  LAYER M2 ;
        RECT 24.72 28.811 27.12 28.813 ;
  LAYER M2 ;
        RECT 24.72 28.727 27.12 28.729 ;
  LAYER M2 ;
        RECT 24.72 28.643 27.12 28.645 ;
  LAYER M1 ;
        RECT 24.704 25.584 24.736 28.092 ;
  LAYER M1 ;
        RECT 24.768 25.584 24.8 28.092 ;
  LAYER M1 ;
        RECT 24.832 25.584 24.864 28.092 ;
  LAYER M1 ;
        RECT 24.896 25.584 24.928 28.092 ;
  LAYER M1 ;
        RECT 24.96 25.584 24.992 28.092 ;
  LAYER M1 ;
        RECT 25.024 25.584 25.056 28.092 ;
  LAYER M1 ;
        RECT 25.088 25.584 25.12 28.092 ;
  LAYER M1 ;
        RECT 25.152 25.584 25.184 28.092 ;
  LAYER M1 ;
        RECT 25.216 25.584 25.248 28.092 ;
  LAYER M1 ;
        RECT 25.28 25.584 25.312 28.092 ;
  LAYER M1 ;
        RECT 25.344 25.584 25.376 28.092 ;
  LAYER M1 ;
        RECT 25.408 25.584 25.44 28.092 ;
  LAYER M1 ;
        RECT 25.472 25.584 25.504 28.092 ;
  LAYER M1 ;
        RECT 25.536 25.584 25.568 28.092 ;
  LAYER M1 ;
        RECT 25.6 25.584 25.632 28.092 ;
  LAYER M1 ;
        RECT 25.664 25.584 25.696 28.092 ;
  LAYER M1 ;
        RECT 25.728 25.584 25.76 28.092 ;
  LAYER M1 ;
        RECT 25.792 25.584 25.824 28.092 ;
  LAYER M1 ;
        RECT 25.856 25.584 25.888 28.092 ;
  LAYER M1 ;
        RECT 25.92 25.584 25.952 28.092 ;
  LAYER M1 ;
        RECT 25.984 25.584 26.016 28.092 ;
  LAYER M1 ;
        RECT 26.048 25.584 26.08 28.092 ;
  LAYER M1 ;
        RECT 26.112 25.584 26.144 28.092 ;
  LAYER M1 ;
        RECT 26.176 25.584 26.208 28.092 ;
  LAYER M1 ;
        RECT 26.24 25.584 26.272 28.092 ;
  LAYER M1 ;
        RECT 26.304 25.584 26.336 28.092 ;
  LAYER M1 ;
        RECT 26.368 25.584 26.4 28.092 ;
  LAYER M1 ;
        RECT 26.432 25.584 26.464 28.092 ;
  LAYER M1 ;
        RECT 26.496 25.584 26.528 28.092 ;
  LAYER M1 ;
        RECT 26.56 25.584 26.592 28.092 ;
  LAYER M1 ;
        RECT 26.624 25.584 26.656 28.092 ;
  LAYER M1 ;
        RECT 26.688 25.584 26.72 28.092 ;
  LAYER M1 ;
        RECT 26.752 25.584 26.784 28.092 ;
  LAYER M1 ;
        RECT 26.816 25.584 26.848 28.092 ;
  LAYER M1 ;
        RECT 26.88 25.584 26.912 28.092 ;
  LAYER M1 ;
        RECT 26.944 25.584 26.976 28.092 ;
  LAYER M1 ;
        RECT 27.008 25.584 27.04 28.092 ;
  LAYER M2 ;
        RECT 24.684 27.976 27.156 28.008 ;
  LAYER M2 ;
        RECT 24.684 27.912 27.156 27.944 ;
  LAYER M2 ;
        RECT 24.684 27.848 27.156 27.88 ;
  LAYER M2 ;
        RECT 24.684 27.784 27.156 27.816 ;
  LAYER M2 ;
        RECT 24.684 27.72 27.156 27.752 ;
  LAYER M2 ;
        RECT 24.684 27.656 27.156 27.688 ;
  LAYER M2 ;
        RECT 24.684 27.592 27.156 27.624 ;
  LAYER M2 ;
        RECT 24.684 27.528 27.156 27.56 ;
  LAYER M2 ;
        RECT 24.684 27.464 27.156 27.496 ;
  LAYER M2 ;
        RECT 24.684 27.4 27.156 27.432 ;
  LAYER M2 ;
        RECT 24.684 27.336 27.156 27.368 ;
  LAYER M2 ;
        RECT 24.684 27.272 27.156 27.304 ;
  LAYER M2 ;
        RECT 24.684 27.208 27.156 27.24 ;
  LAYER M2 ;
        RECT 24.684 27.144 27.156 27.176 ;
  LAYER M2 ;
        RECT 24.684 27.08 27.156 27.112 ;
  LAYER M2 ;
        RECT 24.684 27.016 27.156 27.048 ;
  LAYER M2 ;
        RECT 24.684 26.952 27.156 26.984 ;
  LAYER M2 ;
        RECT 24.684 26.888 27.156 26.92 ;
  LAYER M2 ;
        RECT 24.684 26.824 27.156 26.856 ;
  LAYER M2 ;
        RECT 24.684 26.76 27.156 26.792 ;
  LAYER M2 ;
        RECT 24.684 26.696 27.156 26.728 ;
  LAYER M2 ;
        RECT 24.684 26.632 27.156 26.664 ;
  LAYER M2 ;
        RECT 24.684 26.568 27.156 26.6 ;
  LAYER M2 ;
        RECT 24.684 26.504 27.156 26.536 ;
  LAYER M2 ;
        RECT 24.684 26.44 27.156 26.472 ;
  LAYER M2 ;
        RECT 24.684 26.376 27.156 26.408 ;
  LAYER M2 ;
        RECT 24.684 26.312 27.156 26.344 ;
  LAYER M2 ;
        RECT 24.684 26.248 27.156 26.28 ;
  LAYER M2 ;
        RECT 24.684 26.184 27.156 26.216 ;
  LAYER M2 ;
        RECT 24.684 26.12 27.156 26.152 ;
  LAYER M2 ;
        RECT 24.684 26.056 27.156 26.088 ;
  LAYER M2 ;
        RECT 24.684 25.992 27.156 26.024 ;
  LAYER M2 ;
        RECT 24.684 25.928 27.156 25.96 ;
  LAYER M2 ;
        RECT 24.684 25.864 27.156 25.896 ;
  LAYER M2 ;
        RECT 24.684 25.8 27.156 25.832 ;
  LAYER M2 ;
        RECT 24.684 25.736 27.156 25.768 ;
  LAYER M3 ;
        RECT 24.704 25.584 24.736 28.092 ;
  LAYER M3 ;
        RECT 24.768 25.584 24.8 28.092 ;
  LAYER M3 ;
        RECT 24.832 25.584 24.864 28.092 ;
  LAYER M3 ;
        RECT 24.896 25.584 24.928 28.092 ;
  LAYER M3 ;
        RECT 24.96 25.584 24.992 28.092 ;
  LAYER M3 ;
        RECT 25.024 25.584 25.056 28.092 ;
  LAYER M3 ;
        RECT 25.088 25.584 25.12 28.092 ;
  LAYER M3 ;
        RECT 25.152 25.584 25.184 28.092 ;
  LAYER M3 ;
        RECT 25.216 25.584 25.248 28.092 ;
  LAYER M3 ;
        RECT 25.28 25.584 25.312 28.092 ;
  LAYER M3 ;
        RECT 25.344 25.584 25.376 28.092 ;
  LAYER M3 ;
        RECT 25.408 25.584 25.44 28.092 ;
  LAYER M3 ;
        RECT 25.472 25.584 25.504 28.092 ;
  LAYER M3 ;
        RECT 25.536 25.584 25.568 28.092 ;
  LAYER M3 ;
        RECT 25.6 25.584 25.632 28.092 ;
  LAYER M3 ;
        RECT 25.664 25.584 25.696 28.092 ;
  LAYER M3 ;
        RECT 25.728 25.584 25.76 28.092 ;
  LAYER M3 ;
        RECT 25.792 25.584 25.824 28.092 ;
  LAYER M3 ;
        RECT 25.856 25.584 25.888 28.092 ;
  LAYER M3 ;
        RECT 25.92 25.584 25.952 28.092 ;
  LAYER M3 ;
        RECT 25.984 25.584 26.016 28.092 ;
  LAYER M3 ;
        RECT 26.048 25.584 26.08 28.092 ;
  LAYER M3 ;
        RECT 26.112 25.584 26.144 28.092 ;
  LAYER M3 ;
        RECT 26.176 25.584 26.208 28.092 ;
  LAYER M3 ;
        RECT 26.24 25.584 26.272 28.092 ;
  LAYER M3 ;
        RECT 26.304 25.584 26.336 28.092 ;
  LAYER M3 ;
        RECT 26.368 25.584 26.4 28.092 ;
  LAYER M3 ;
        RECT 26.432 25.584 26.464 28.092 ;
  LAYER M3 ;
        RECT 26.496 25.584 26.528 28.092 ;
  LAYER M3 ;
        RECT 26.56 25.584 26.592 28.092 ;
  LAYER M3 ;
        RECT 26.624 25.584 26.656 28.092 ;
  LAYER M3 ;
        RECT 26.688 25.584 26.72 28.092 ;
  LAYER M3 ;
        RECT 26.752 25.584 26.784 28.092 ;
  LAYER M3 ;
        RECT 26.816 25.584 26.848 28.092 ;
  LAYER M3 ;
        RECT 26.88 25.584 26.912 28.092 ;
  LAYER M3 ;
        RECT 26.944 25.584 26.976 28.092 ;
  LAYER M3 ;
        RECT 27.008 25.584 27.04 28.092 ;
  LAYER M3 ;
        RECT 27.104 25.584 27.136 28.092 ;
  LAYER M1 ;
        RECT 24.719 25.62 24.721 28.056 ;
  LAYER M1 ;
        RECT 24.799 25.62 24.801 28.056 ;
  LAYER M1 ;
        RECT 24.879 25.62 24.881 28.056 ;
  LAYER M1 ;
        RECT 24.959 25.62 24.961 28.056 ;
  LAYER M1 ;
        RECT 25.039 25.62 25.041 28.056 ;
  LAYER M1 ;
        RECT 25.119 25.62 25.121 28.056 ;
  LAYER M1 ;
        RECT 25.199 25.62 25.201 28.056 ;
  LAYER M1 ;
        RECT 25.279 25.62 25.281 28.056 ;
  LAYER M1 ;
        RECT 25.359 25.62 25.361 28.056 ;
  LAYER M1 ;
        RECT 25.439 25.62 25.441 28.056 ;
  LAYER M1 ;
        RECT 25.519 25.62 25.521 28.056 ;
  LAYER M1 ;
        RECT 25.599 25.62 25.601 28.056 ;
  LAYER M1 ;
        RECT 25.679 25.62 25.681 28.056 ;
  LAYER M1 ;
        RECT 25.759 25.62 25.761 28.056 ;
  LAYER M1 ;
        RECT 25.839 25.62 25.841 28.056 ;
  LAYER M1 ;
        RECT 25.919 25.62 25.921 28.056 ;
  LAYER M1 ;
        RECT 25.999 25.62 26.001 28.056 ;
  LAYER M1 ;
        RECT 26.079 25.62 26.081 28.056 ;
  LAYER M1 ;
        RECT 26.159 25.62 26.161 28.056 ;
  LAYER M1 ;
        RECT 26.239 25.62 26.241 28.056 ;
  LAYER M1 ;
        RECT 26.319 25.62 26.321 28.056 ;
  LAYER M1 ;
        RECT 26.399 25.62 26.401 28.056 ;
  LAYER M1 ;
        RECT 26.479 25.62 26.481 28.056 ;
  LAYER M1 ;
        RECT 26.559 25.62 26.561 28.056 ;
  LAYER M1 ;
        RECT 26.639 25.62 26.641 28.056 ;
  LAYER M1 ;
        RECT 26.719 25.62 26.721 28.056 ;
  LAYER M1 ;
        RECT 26.799 25.62 26.801 28.056 ;
  LAYER M1 ;
        RECT 26.879 25.62 26.881 28.056 ;
  LAYER M1 ;
        RECT 26.959 25.62 26.961 28.056 ;
  LAYER M1 ;
        RECT 27.039 25.62 27.041 28.056 ;
  LAYER M2 ;
        RECT 24.72 28.055 27.12 28.057 ;
  LAYER M2 ;
        RECT 24.72 27.971 27.12 27.973 ;
  LAYER M2 ;
        RECT 24.72 27.887 27.12 27.889 ;
  LAYER M2 ;
        RECT 24.72 27.803 27.12 27.805 ;
  LAYER M2 ;
        RECT 24.72 27.719 27.12 27.721 ;
  LAYER M2 ;
        RECT 24.72 27.635 27.12 27.637 ;
  LAYER M2 ;
        RECT 24.72 27.551 27.12 27.553 ;
  LAYER M2 ;
        RECT 24.72 27.467 27.12 27.469 ;
  LAYER M2 ;
        RECT 24.72 27.383 27.12 27.385 ;
  LAYER M2 ;
        RECT 24.72 27.299 27.12 27.301 ;
  LAYER M2 ;
        RECT 24.72 27.215 27.12 27.217 ;
  LAYER M2 ;
        RECT 24.72 27.131 27.12 27.133 ;
  LAYER M2 ;
        RECT 24.72 27.0475 27.12 27.0495 ;
  LAYER M2 ;
        RECT 24.72 26.963 27.12 26.965 ;
  LAYER M2 ;
        RECT 24.72 26.879 27.12 26.881 ;
  LAYER M2 ;
        RECT 24.72 26.795 27.12 26.797 ;
  LAYER M2 ;
        RECT 24.72 26.711 27.12 26.713 ;
  LAYER M2 ;
        RECT 24.72 26.627 27.12 26.629 ;
  LAYER M2 ;
        RECT 24.72 26.543 27.12 26.545 ;
  LAYER M2 ;
        RECT 24.72 26.459 27.12 26.461 ;
  LAYER M2 ;
        RECT 24.72 26.375 27.12 26.377 ;
  LAYER M2 ;
        RECT 24.72 26.291 27.12 26.293 ;
  LAYER M2 ;
        RECT 24.72 26.207 27.12 26.209 ;
  LAYER M2 ;
        RECT 24.72 26.123 27.12 26.125 ;
  LAYER M2 ;
        RECT 24.72 26.039 27.12 26.041 ;
  LAYER M2 ;
        RECT 24.72 25.955 27.12 25.957 ;
  LAYER M2 ;
        RECT 24.72 25.871 27.12 25.873 ;
  LAYER M2 ;
        RECT 24.72 25.787 27.12 25.789 ;
  LAYER M2 ;
        RECT 24.72 25.703 27.12 25.705 ;
  LAYER M1 ;
        RECT 24.704 22.644 24.736 25.152 ;
  LAYER M1 ;
        RECT 24.768 22.644 24.8 25.152 ;
  LAYER M1 ;
        RECT 24.832 22.644 24.864 25.152 ;
  LAYER M1 ;
        RECT 24.896 22.644 24.928 25.152 ;
  LAYER M1 ;
        RECT 24.96 22.644 24.992 25.152 ;
  LAYER M1 ;
        RECT 25.024 22.644 25.056 25.152 ;
  LAYER M1 ;
        RECT 25.088 22.644 25.12 25.152 ;
  LAYER M1 ;
        RECT 25.152 22.644 25.184 25.152 ;
  LAYER M1 ;
        RECT 25.216 22.644 25.248 25.152 ;
  LAYER M1 ;
        RECT 25.28 22.644 25.312 25.152 ;
  LAYER M1 ;
        RECT 25.344 22.644 25.376 25.152 ;
  LAYER M1 ;
        RECT 25.408 22.644 25.44 25.152 ;
  LAYER M1 ;
        RECT 25.472 22.644 25.504 25.152 ;
  LAYER M1 ;
        RECT 25.536 22.644 25.568 25.152 ;
  LAYER M1 ;
        RECT 25.6 22.644 25.632 25.152 ;
  LAYER M1 ;
        RECT 25.664 22.644 25.696 25.152 ;
  LAYER M1 ;
        RECT 25.728 22.644 25.76 25.152 ;
  LAYER M1 ;
        RECT 25.792 22.644 25.824 25.152 ;
  LAYER M1 ;
        RECT 25.856 22.644 25.888 25.152 ;
  LAYER M1 ;
        RECT 25.92 22.644 25.952 25.152 ;
  LAYER M1 ;
        RECT 25.984 22.644 26.016 25.152 ;
  LAYER M1 ;
        RECT 26.048 22.644 26.08 25.152 ;
  LAYER M1 ;
        RECT 26.112 22.644 26.144 25.152 ;
  LAYER M1 ;
        RECT 26.176 22.644 26.208 25.152 ;
  LAYER M1 ;
        RECT 26.24 22.644 26.272 25.152 ;
  LAYER M1 ;
        RECT 26.304 22.644 26.336 25.152 ;
  LAYER M1 ;
        RECT 26.368 22.644 26.4 25.152 ;
  LAYER M1 ;
        RECT 26.432 22.644 26.464 25.152 ;
  LAYER M1 ;
        RECT 26.496 22.644 26.528 25.152 ;
  LAYER M1 ;
        RECT 26.56 22.644 26.592 25.152 ;
  LAYER M1 ;
        RECT 26.624 22.644 26.656 25.152 ;
  LAYER M1 ;
        RECT 26.688 22.644 26.72 25.152 ;
  LAYER M1 ;
        RECT 26.752 22.644 26.784 25.152 ;
  LAYER M1 ;
        RECT 26.816 22.644 26.848 25.152 ;
  LAYER M1 ;
        RECT 26.88 22.644 26.912 25.152 ;
  LAYER M1 ;
        RECT 26.944 22.644 26.976 25.152 ;
  LAYER M1 ;
        RECT 27.008 22.644 27.04 25.152 ;
  LAYER M2 ;
        RECT 24.684 25.036 27.156 25.068 ;
  LAYER M2 ;
        RECT 24.684 24.972 27.156 25.004 ;
  LAYER M2 ;
        RECT 24.684 24.908 27.156 24.94 ;
  LAYER M2 ;
        RECT 24.684 24.844 27.156 24.876 ;
  LAYER M2 ;
        RECT 24.684 24.78 27.156 24.812 ;
  LAYER M2 ;
        RECT 24.684 24.716 27.156 24.748 ;
  LAYER M2 ;
        RECT 24.684 24.652 27.156 24.684 ;
  LAYER M2 ;
        RECT 24.684 24.588 27.156 24.62 ;
  LAYER M2 ;
        RECT 24.684 24.524 27.156 24.556 ;
  LAYER M2 ;
        RECT 24.684 24.46 27.156 24.492 ;
  LAYER M2 ;
        RECT 24.684 24.396 27.156 24.428 ;
  LAYER M2 ;
        RECT 24.684 24.332 27.156 24.364 ;
  LAYER M2 ;
        RECT 24.684 24.268 27.156 24.3 ;
  LAYER M2 ;
        RECT 24.684 24.204 27.156 24.236 ;
  LAYER M2 ;
        RECT 24.684 24.14 27.156 24.172 ;
  LAYER M2 ;
        RECT 24.684 24.076 27.156 24.108 ;
  LAYER M2 ;
        RECT 24.684 24.012 27.156 24.044 ;
  LAYER M2 ;
        RECT 24.684 23.948 27.156 23.98 ;
  LAYER M2 ;
        RECT 24.684 23.884 27.156 23.916 ;
  LAYER M2 ;
        RECT 24.684 23.82 27.156 23.852 ;
  LAYER M2 ;
        RECT 24.684 23.756 27.156 23.788 ;
  LAYER M2 ;
        RECT 24.684 23.692 27.156 23.724 ;
  LAYER M2 ;
        RECT 24.684 23.628 27.156 23.66 ;
  LAYER M2 ;
        RECT 24.684 23.564 27.156 23.596 ;
  LAYER M2 ;
        RECT 24.684 23.5 27.156 23.532 ;
  LAYER M2 ;
        RECT 24.684 23.436 27.156 23.468 ;
  LAYER M2 ;
        RECT 24.684 23.372 27.156 23.404 ;
  LAYER M2 ;
        RECT 24.684 23.308 27.156 23.34 ;
  LAYER M2 ;
        RECT 24.684 23.244 27.156 23.276 ;
  LAYER M2 ;
        RECT 24.684 23.18 27.156 23.212 ;
  LAYER M2 ;
        RECT 24.684 23.116 27.156 23.148 ;
  LAYER M2 ;
        RECT 24.684 23.052 27.156 23.084 ;
  LAYER M2 ;
        RECT 24.684 22.988 27.156 23.02 ;
  LAYER M2 ;
        RECT 24.684 22.924 27.156 22.956 ;
  LAYER M2 ;
        RECT 24.684 22.86 27.156 22.892 ;
  LAYER M2 ;
        RECT 24.684 22.796 27.156 22.828 ;
  LAYER M3 ;
        RECT 24.704 22.644 24.736 25.152 ;
  LAYER M3 ;
        RECT 24.768 22.644 24.8 25.152 ;
  LAYER M3 ;
        RECT 24.832 22.644 24.864 25.152 ;
  LAYER M3 ;
        RECT 24.896 22.644 24.928 25.152 ;
  LAYER M3 ;
        RECT 24.96 22.644 24.992 25.152 ;
  LAYER M3 ;
        RECT 25.024 22.644 25.056 25.152 ;
  LAYER M3 ;
        RECT 25.088 22.644 25.12 25.152 ;
  LAYER M3 ;
        RECT 25.152 22.644 25.184 25.152 ;
  LAYER M3 ;
        RECT 25.216 22.644 25.248 25.152 ;
  LAYER M3 ;
        RECT 25.28 22.644 25.312 25.152 ;
  LAYER M3 ;
        RECT 25.344 22.644 25.376 25.152 ;
  LAYER M3 ;
        RECT 25.408 22.644 25.44 25.152 ;
  LAYER M3 ;
        RECT 25.472 22.644 25.504 25.152 ;
  LAYER M3 ;
        RECT 25.536 22.644 25.568 25.152 ;
  LAYER M3 ;
        RECT 25.6 22.644 25.632 25.152 ;
  LAYER M3 ;
        RECT 25.664 22.644 25.696 25.152 ;
  LAYER M3 ;
        RECT 25.728 22.644 25.76 25.152 ;
  LAYER M3 ;
        RECT 25.792 22.644 25.824 25.152 ;
  LAYER M3 ;
        RECT 25.856 22.644 25.888 25.152 ;
  LAYER M3 ;
        RECT 25.92 22.644 25.952 25.152 ;
  LAYER M3 ;
        RECT 25.984 22.644 26.016 25.152 ;
  LAYER M3 ;
        RECT 26.048 22.644 26.08 25.152 ;
  LAYER M3 ;
        RECT 26.112 22.644 26.144 25.152 ;
  LAYER M3 ;
        RECT 26.176 22.644 26.208 25.152 ;
  LAYER M3 ;
        RECT 26.24 22.644 26.272 25.152 ;
  LAYER M3 ;
        RECT 26.304 22.644 26.336 25.152 ;
  LAYER M3 ;
        RECT 26.368 22.644 26.4 25.152 ;
  LAYER M3 ;
        RECT 26.432 22.644 26.464 25.152 ;
  LAYER M3 ;
        RECT 26.496 22.644 26.528 25.152 ;
  LAYER M3 ;
        RECT 26.56 22.644 26.592 25.152 ;
  LAYER M3 ;
        RECT 26.624 22.644 26.656 25.152 ;
  LAYER M3 ;
        RECT 26.688 22.644 26.72 25.152 ;
  LAYER M3 ;
        RECT 26.752 22.644 26.784 25.152 ;
  LAYER M3 ;
        RECT 26.816 22.644 26.848 25.152 ;
  LAYER M3 ;
        RECT 26.88 22.644 26.912 25.152 ;
  LAYER M3 ;
        RECT 26.944 22.644 26.976 25.152 ;
  LAYER M3 ;
        RECT 27.008 22.644 27.04 25.152 ;
  LAYER M3 ;
        RECT 27.104 22.644 27.136 25.152 ;
  LAYER M1 ;
        RECT 24.719 22.68 24.721 25.116 ;
  LAYER M1 ;
        RECT 24.799 22.68 24.801 25.116 ;
  LAYER M1 ;
        RECT 24.879 22.68 24.881 25.116 ;
  LAYER M1 ;
        RECT 24.959 22.68 24.961 25.116 ;
  LAYER M1 ;
        RECT 25.039 22.68 25.041 25.116 ;
  LAYER M1 ;
        RECT 25.119 22.68 25.121 25.116 ;
  LAYER M1 ;
        RECT 25.199 22.68 25.201 25.116 ;
  LAYER M1 ;
        RECT 25.279 22.68 25.281 25.116 ;
  LAYER M1 ;
        RECT 25.359 22.68 25.361 25.116 ;
  LAYER M1 ;
        RECT 25.439 22.68 25.441 25.116 ;
  LAYER M1 ;
        RECT 25.519 22.68 25.521 25.116 ;
  LAYER M1 ;
        RECT 25.599 22.68 25.601 25.116 ;
  LAYER M1 ;
        RECT 25.679 22.68 25.681 25.116 ;
  LAYER M1 ;
        RECT 25.759 22.68 25.761 25.116 ;
  LAYER M1 ;
        RECT 25.839 22.68 25.841 25.116 ;
  LAYER M1 ;
        RECT 25.919 22.68 25.921 25.116 ;
  LAYER M1 ;
        RECT 25.999 22.68 26.001 25.116 ;
  LAYER M1 ;
        RECT 26.079 22.68 26.081 25.116 ;
  LAYER M1 ;
        RECT 26.159 22.68 26.161 25.116 ;
  LAYER M1 ;
        RECT 26.239 22.68 26.241 25.116 ;
  LAYER M1 ;
        RECT 26.319 22.68 26.321 25.116 ;
  LAYER M1 ;
        RECT 26.399 22.68 26.401 25.116 ;
  LAYER M1 ;
        RECT 26.479 22.68 26.481 25.116 ;
  LAYER M1 ;
        RECT 26.559 22.68 26.561 25.116 ;
  LAYER M1 ;
        RECT 26.639 22.68 26.641 25.116 ;
  LAYER M1 ;
        RECT 26.719 22.68 26.721 25.116 ;
  LAYER M1 ;
        RECT 26.799 22.68 26.801 25.116 ;
  LAYER M1 ;
        RECT 26.879 22.68 26.881 25.116 ;
  LAYER M1 ;
        RECT 26.959 22.68 26.961 25.116 ;
  LAYER M1 ;
        RECT 27.039 22.68 27.041 25.116 ;
  LAYER M2 ;
        RECT 24.72 25.115 27.12 25.117 ;
  LAYER M2 ;
        RECT 24.72 25.031 27.12 25.033 ;
  LAYER M2 ;
        RECT 24.72 24.947 27.12 24.949 ;
  LAYER M2 ;
        RECT 24.72 24.863 27.12 24.865 ;
  LAYER M2 ;
        RECT 24.72 24.779 27.12 24.781 ;
  LAYER M2 ;
        RECT 24.72 24.695 27.12 24.697 ;
  LAYER M2 ;
        RECT 24.72 24.611 27.12 24.613 ;
  LAYER M2 ;
        RECT 24.72 24.527 27.12 24.529 ;
  LAYER M2 ;
        RECT 24.72 24.443 27.12 24.445 ;
  LAYER M2 ;
        RECT 24.72 24.359 27.12 24.361 ;
  LAYER M2 ;
        RECT 24.72 24.275 27.12 24.277 ;
  LAYER M2 ;
        RECT 24.72 24.191 27.12 24.193 ;
  LAYER M2 ;
        RECT 24.72 24.1075 27.12 24.1095 ;
  LAYER M2 ;
        RECT 24.72 24.023 27.12 24.025 ;
  LAYER M2 ;
        RECT 24.72 23.939 27.12 23.941 ;
  LAYER M2 ;
        RECT 24.72 23.855 27.12 23.857 ;
  LAYER M2 ;
        RECT 24.72 23.771 27.12 23.773 ;
  LAYER M2 ;
        RECT 24.72 23.687 27.12 23.689 ;
  LAYER M2 ;
        RECT 24.72 23.603 27.12 23.605 ;
  LAYER M2 ;
        RECT 24.72 23.519 27.12 23.521 ;
  LAYER M2 ;
        RECT 24.72 23.435 27.12 23.437 ;
  LAYER M2 ;
        RECT 24.72 23.351 27.12 23.353 ;
  LAYER M2 ;
        RECT 24.72 23.267 27.12 23.269 ;
  LAYER M2 ;
        RECT 24.72 23.183 27.12 23.185 ;
  LAYER M2 ;
        RECT 24.72 23.099 27.12 23.101 ;
  LAYER M2 ;
        RECT 24.72 23.015 27.12 23.017 ;
  LAYER M2 ;
        RECT 24.72 22.931 27.12 22.933 ;
  LAYER M2 ;
        RECT 24.72 22.847 27.12 22.849 ;
  LAYER M2 ;
        RECT 24.72 22.763 27.12 22.765 ;
  LAYER M1 ;
        RECT 24.704 19.704 24.736 22.212 ;
  LAYER M1 ;
        RECT 24.768 19.704 24.8 22.212 ;
  LAYER M1 ;
        RECT 24.832 19.704 24.864 22.212 ;
  LAYER M1 ;
        RECT 24.896 19.704 24.928 22.212 ;
  LAYER M1 ;
        RECT 24.96 19.704 24.992 22.212 ;
  LAYER M1 ;
        RECT 25.024 19.704 25.056 22.212 ;
  LAYER M1 ;
        RECT 25.088 19.704 25.12 22.212 ;
  LAYER M1 ;
        RECT 25.152 19.704 25.184 22.212 ;
  LAYER M1 ;
        RECT 25.216 19.704 25.248 22.212 ;
  LAYER M1 ;
        RECT 25.28 19.704 25.312 22.212 ;
  LAYER M1 ;
        RECT 25.344 19.704 25.376 22.212 ;
  LAYER M1 ;
        RECT 25.408 19.704 25.44 22.212 ;
  LAYER M1 ;
        RECT 25.472 19.704 25.504 22.212 ;
  LAYER M1 ;
        RECT 25.536 19.704 25.568 22.212 ;
  LAYER M1 ;
        RECT 25.6 19.704 25.632 22.212 ;
  LAYER M1 ;
        RECT 25.664 19.704 25.696 22.212 ;
  LAYER M1 ;
        RECT 25.728 19.704 25.76 22.212 ;
  LAYER M1 ;
        RECT 25.792 19.704 25.824 22.212 ;
  LAYER M1 ;
        RECT 25.856 19.704 25.888 22.212 ;
  LAYER M1 ;
        RECT 25.92 19.704 25.952 22.212 ;
  LAYER M1 ;
        RECT 25.984 19.704 26.016 22.212 ;
  LAYER M1 ;
        RECT 26.048 19.704 26.08 22.212 ;
  LAYER M1 ;
        RECT 26.112 19.704 26.144 22.212 ;
  LAYER M1 ;
        RECT 26.176 19.704 26.208 22.212 ;
  LAYER M1 ;
        RECT 26.24 19.704 26.272 22.212 ;
  LAYER M1 ;
        RECT 26.304 19.704 26.336 22.212 ;
  LAYER M1 ;
        RECT 26.368 19.704 26.4 22.212 ;
  LAYER M1 ;
        RECT 26.432 19.704 26.464 22.212 ;
  LAYER M1 ;
        RECT 26.496 19.704 26.528 22.212 ;
  LAYER M1 ;
        RECT 26.56 19.704 26.592 22.212 ;
  LAYER M1 ;
        RECT 26.624 19.704 26.656 22.212 ;
  LAYER M1 ;
        RECT 26.688 19.704 26.72 22.212 ;
  LAYER M1 ;
        RECT 26.752 19.704 26.784 22.212 ;
  LAYER M1 ;
        RECT 26.816 19.704 26.848 22.212 ;
  LAYER M1 ;
        RECT 26.88 19.704 26.912 22.212 ;
  LAYER M1 ;
        RECT 26.944 19.704 26.976 22.212 ;
  LAYER M1 ;
        RECT 27.008 19.704 27.04 22.212 ;
  LAYER M2 ;
        RECT 24.684 22.096 27.156 22.128 ;
  LAYER M2 ;
        RECT 24.684 22.032 27.156 22.064 ;
  LAYER M2 ;
        RECT 24.684 21.968 27.156 22 ;
  LAYER M2 ;
        RECT 24.684 21.904 27.156 21.936 ;
  LAYER M2 ;
        RECT 24.684 21.84 27.156 21.872 ;
  LAYER M2 ;
        RECT 24.684 21.776 27.156 21.808 ;
  LAYER M2 ;
        RECT 24.684 21.712 27.156 21.744 ;
  LAYER M2 ;
        RECT 24.684 21.648 27.156 21.68 ;
  LAYER M2 ;
        RECT 24.684 21.584 27.156 21.616 ;
  LAYER M2 ;
        RECT 24.684 21.52 27.156 21.552 ;
  LAYER M2 ;
        RECT 24.684 21.456 27.156 21.488 ;
  LAYER M2 ;
        RECT 24.684 21.392 27.156 21.424 ;
  LAYER M2 ;
        RECT 24.684 21.328 27.156 21.36 ;
  LAYER M2 ;
        RECT 24.684 21.264 27.156 21.296 ;
  LAYER M2 ;
        RECT 24.684 21.2 27.156 21.232 ;
  LAYER M2 ;
        RECT 24.684 21.136 27.156 21.168 ;
  LAYER M2 ;
        RECT 24.684 21.072 27.156 21.104 ;
  LAYER M2 ;
        RECT 24.684 21.008 27.156 21.04 ;
  LAYER M2 ;
        RECT 24.684 20.944 27.156 20.976 ;
  LAYER M2 ;
        RECT 24.684 20.88 27.156 20.912 ;
  LAYER M2 ;
        RECT 24.684 20.816 27.156 20.848 ;
  LAYER M2 ;
        RECT 24.684 20.752 27.156 20.784 ;
  LAYER M2 ;
        RECT 24.684 20.688 27.156 20.72 ;
  LAYER M2 ;
        RECT 24.684 20.624 27.156 20.656 ;
  LAYER M2 ;
        RECT 24.684 20.56 27.156 20.592 ;
  LAYER M2 ;
        RECT 24.684 20.496 27.156 20.528 ;
  LAYER M2 ;
        RECT 24.684 20.432 27.156 20.464 ;
  LAYER M2 ;
        RECT 24.684 20.368 27.156 20.4 ;
  LAYER M2 ;
        RECT 24.684 20.304 27.156 20.336 ;
  LAYER M2 ;
        RECT 24.684 20.24 27.156 20.272 ;
  LAYER M2 ;
        RECT 24.684 20.176 27.156 20.208 ;
  LAYER M2 ;
        RECT 24.684 20.112 27.156 20.144 ;
  LAYER M2 ;
        RECT 24.684 20.048 27.156 20.08 ;
  LAYER M2 ;
        RECT 24.684 19.984 27.156 20.016 ;
  LAYER M2 ;
        RECT 24.684 19.92 27.156 19.952 ;
  LAYER M2 ;
        RECT 24.684 19.856 27.156 19.888 ;
  LAYER M3 ;
        RECT 24.704 19.704 24.736 22.212 ;
  LAYER M3 ;
        RECT 24.768 19.704 24.8 22.212 ;
  LAYER M3 ;
        RECT 24.832 19.704 24.864 22.212 ;
  LAYER M3 ;
        RECT 24.896 19.704 24.928 22.212 ;
  LAYER M3 ;
        RECT 24.96 19.704 24.992 22.212 ;
  LAYER M3 ;
        RECT 25.024 19.704 25.056 22.212 ;
  LAYER M3 ;
        RECT 25.088 19.704 25.12 22.212 ;
  LAYER M3 ;
        RECT 25.152 19.704 25.184 22.212 ;
  LAYER M3 ;
        RECT 25.216 19.704 25.248 22.212 ;
  LAYER M3 ;
        RECT 25.28 19.704 25.312 22.212 ;
  LAYER M3 ;
        RECT 25.344 19.704 25.376 22.212 ;
  LAYER M3 ;
        RECT 25.408 19.704 25.44 22.212 ;
  LAYER M3 ;
        RECT 25.472 19.704 25.504 22.212 ;
  LAYER M3 ;
        RECT 25.536 19.704 25.568 22.212 ;
  LAYER M3 ;
        RECT 25.6 19.704 25.632 22.212 ;
  LAYER M3 ;
        RECT 25.664 19.704 25.696 22.212 ;
  LAYER M3 ;
        RECT 25.728 19.704 25.76 22.212 ;
  LAYER M3 ;
        RECT 25.792 19.704 25.824 22.212 ;
  LAYER M3 ;
        RECT 25.856 19.704 25.888 22.212 ;
  LAYER M3 ;
        RECT 25.92 19.704 25.952 22.212 ;
  LAYER M3 ;
        RECT 25.984 19.704 26.016 22.212 ;
  LAYER M3 ;
        RECT 26.048 19.704 26.08 22.212 ;
  LAYER M3 ;
        RECT 26.112 19.704 26.144 22.212 ;
  LAYER M3 ;
        RECT 26.176 19.704 26.208 22.212 ;
  LAYER M3 ;
        RECT 26.24 19.704 26.272 22.212 ;
  LAYER M3 ;
        RECT 26.304 19.704 26.336 22.212 ;
  LAYER M3 ;
        RECT 26.368 19.704 26.4 22.212 ;
  LAYER M3 ;
        RECT 26.432 19.704 26.464 22.212 ;
  LAYER M3 ;
        RECT 26.496 19.704 26.528 22.212 ;
  LAYER M3 ;
        RECT 26.56 19.704 26.592 22.212 ;
  LAYER M3 ;
        RECT 26.624 19.704 26.656 22.212 ;
  LAYER M3 ;
        RECT 26.688 19.704 26.72 22.212 ;
  LAYER M3 ;
        RECT 26.752 19.704 26.784 22.212 ;
  LAYER M3 ;
        RECT 26.816 19.704 26.848 22.212 ;
  LAYER M3 ;
        RECT 26.88 19.704 26.912 22.212 ;
  LAYER M3 ;
        RECT 26.944 19.704 26.976 22.212 ;
  LAYER M3 ;
        RECT 27.008 19.704 27.04 22.212 ;
  LAYER M3 ;
        RECT 27.104 19.704 27.136 22.212 ;
  LAYER M1 ;
        RECT 24.719 19.74 24.721 22.176 ;
  LAYER M1 ;
        RECT 24.799 19.74 24.801 22.176 ;
  LAYER M1 ;
        RECT 24.879 19.74 24.881 22.176 ;
  LAYER M1 ;
        RECT 24.959 19.74 24.961 22.176 ;
  LAYER M1 ;
        RECT 25.039 19.74 25.041 22.176 ;
  LAYER M1 ;
        RECT 25.119 19.74 25.121 22.176 ;
  LAYER M1 ;
        RECT 25.199 19.74 25.201 22.176 ;
  LAYER M1 ;
        RECT 25.279 19.74 25.281 22.176 ;
  LAYER M1 ;
        RECT 25.359 19.74 25.361 22.176 ;
  LAYER M1 ;
        RECT 25.439 19.74 25.441 22.176 ;
  LAYER M1 ;
        RECT 25.519 19.74 25.521 22.176 ;
  LAYER M1 ;
        RECT 25.599 19.74 25.601 22.176 ;
  LAYER M1 ;
        RECT 25.679 19.74 25.681 22.176 ;
  LAYER M1 ;
        RECT 25.759 19.74 25.761 22.176 ;
  LAYER M1 ;
        RECT 25.839 19.74 25.841 22.176 ;
  LAYER M1 ;
        RECT 25.919 19.74 25.921 22.176 ;
  LAYER M1 ;
        RECT 25.999 19.74 26.001 22.176 ;
  LAYER M1 ;
        RECT 26.079 19.74 26.081 22.176 ;
  LAYER M1 ;
        RECT 26.159 19.74 26.161 22.176 ;
  LAYER M1 ;
        RECT 26.239 19.74 26.241 22.176 ;
  LAYER M1 ;
        RECT 26.319 19.74 26.321 22.176 ;
  LAYER M1 ;
        RECT 26.399 19.74 26.401 22.176 ;
  LAYER M1 ;
        RECT 26.479 19.74 26.481 22.176 ;
  LAYER M1 ;
        RECT 26.559 19.74 26.561 22.176 ;
  LAYER M1 ;
        RECT 26.639 19.74 26.641 22.176 ;
  LAYER M1 ;
        RECT 26.719 19.74 26.721 22.176 ;
  LAYER M1 ;
        RECT 26.799 19.74 26.801 22.176 ;
  LAYER M1 ;
        RECT 26.879 19.74 26.881 22.176 ;
  LAYER M1 ;
        RECT 26.959 19.74 26.961 22.176 ;
  LAYER M1 ;
        RECT 27.039 19.74 27.041 22.176 ;
  LAYER M2 ;
        RECT 24.72 22.175 27.12 22.177 ;
  LAYER M2 ;
        RECT 24.72 22.091 27.12 22.093 ;
  LAYER M2 ;
        RECT 24.72 22.007 27.12 22.009 ;
  LAYER M2 ;
        RECT 24.72 21.923 27.12 21.925 ;
  LAYER M2 ;
        RECT 24.72 21.839 27.12 21.841 ;
  LAYER M2 ;
        RECT 24.72 21.755 27.12 21.757 ;
  LAYER M2 ;
        RECT 24.72 21.671 27.12 21.673 ;
  LAYER M2 ;
        RECT 24.72 21.587 27.12 21.589 ;
  LAYER M2 ;
        RECT 24.72 21.503 27.12 21.505 ;
  LAYER M2 ;
        RECT 24.72 21.419 27.12 21.421 ;
  LAYER M2 ;
        RECT 24.72 21.335 27.12 21.337 ;
  LAYER M2 ;
        RECT 24.72 21.251 27.12 21.253 ;
  LAYER M2 ;
        RECT 24.72 21.1675 27.12 21.1695 ;
  LAYER M2 ;
        RECT 24.72 21.083 27.12 21.085 ;
  LAYER M2 ;
        RECT 24.72 20.999 27.12 21.001 ;
  LAYER M2 ;
        RECT 24.72 20.915 27.12 20.917 ;
  LAYER M2 ;
        RECT 24.72 20.831 27.12 20.833 ;
  LAYER M2 ;
        RECT 24.72 20.747 27.12 20.749 ;
  LAYER M2 ;
        RECT 24.72 20.663 27.12 20.665 ;
  LAYER M2 ;
        RECT 24.72 20.579 27.12 20.581 ;
  LAYER M2 ;
        RECT 24.72 20.495 27.12 20.497 ;
  LAYER M2 ;
        RECT 24.72 20.411 27.12 20.413 ;
  LAYER M2 ;
        RECT 24.72 20.327 27.12 20.329 ;
  LAYER M2 ;
        RECT 24.72 20.243 27.12 20.245 ;
  LAYER M2 ;
        RECT 24.72 20.159 27.12 20.161 ;
  LAYER M2 ;
        RECT 24.72 20.075 27.12 20.077 ;
  LAYER M2 ;
        RECT 24.72 19.991 27.12 19.993 ;
  LAYER M2 ;
        RECT 24.72 19.907 27.12 19.909 ;
  LAYER M2 ;
        RECT 24.72 19.823 27.12 19.825 ;
  LAYER M1 ;
        RECT 27.584 34.404 27.616 36.912 ;
  LAYER M1 ;
        RECT 27.648 34.404 27.68 36.912 ;
  LAYER M1 ;
        RECT 27.712 34.404 27.744 36.912 ;
  LAYER M1 ;
        RECT 27.776 34.404 27.808 36.912 ;
  LAYER M1 ;
        RECT 27.84 34.404 27.872 36.912 ;
  LAYER M1 ;
        RECT 27.904 34.404 27.936 36.912 ;
  LAYER M1 ;
        RECT 27.968 34.404 28 36.912 ;
  LAYER M1 ;
        RECT 28.032 34.404 28.064 36.912 ;
  LAYER M1 ;
        RECT 28.096 34.404 28.128 36.912 ;
  LAYER M1 ;
        RECT 28.16 34.404 28.192 36.912 ;
  LAYER M1 ;
        RECT 28.224 34.404 28.256 36.912 ;
  LAYER M1 ;
        RECT 28.288 34.404 28.32 36.912 ;
  LAYER M1 ;
        RECT 28.352 34.404 28.384 36.912 ;
  LAYER M1 ;
        RECT 28.416 34.404 28.448 36.912 ;
  LAYER M1 ;
        RECT 28.48 34.404 28.512 36.912 ;
  LAYER M1 ;
        RECT 28.544 34.404 28.576 36.912 ;
  LAYER M1 ;
        RECT 28.608 34.404 28.64 36.912 ;
  LAYER M1 ;
        RECT 28.672 34.404 28.704 36.912 ;
  LAYER M1 ;
        RECT 28.736 34.404 28.768 36.912 ;
  LAYER M1 ;
        RECT 28.8 34.404 28.832 36.912 ;
  LAYER M1 ;
        RECT 28.864 34.404 28.896 36.912 ;
  LAYER M1 ;
        RECT 28.928 34.404 28.96 36.912 ;
  LAYER M1 ;
        RECT 28.992 34.404 29.024 36.912 ;
  LAYER M1 ;
        RECT 29.056 34.404 29.088 36.912 ;
  LAYER M1 ;
        RECT 29.12 34.404 29.152 36.912 ;
  LAYER M1 ;
        RECT 29.184 34.404 29.216 36.912 ;
  LAYER M1 ;
        RECT 29.248 34.404 29.28 36.912 ;
  LAYER M1 ;
        RECT 29.312 34.404 29.344 36.912 ;
  LAYER M1 ;
        RECT 29.376 34.404 29.408 36.912 ;
  LAYER M1 ;
        RECT 29.44 34.404 29.472 36.912 ;
  LAYER M1 ;
        RECT 29.504 34.404 29.536 36.912 ;
  LAYER M1 ;
        RECT 29.568 34.404 29.6 36.912 ;
  LAYER M1 ;
        RECT 29.632 34.404 29.664 36.912 ;
  LAYER M1 ;
        RECT 29.696 34.404 29.728 36.912 ;
  LAYER M1 ;
        RECT 29.76 34.404 29.792 36.912 ;
  LAYER M1 ;
        RECT 29.824 34.404 29.856 36.912 ;
  LAYER M1 ;
        RECT 29.888 34.404 29.92 36.912 ;
  LAYER M2 ;
        RECT 27.564 36.796 30.036 36.828 ;
  LAYER M2 ;
        RECT 27.564 36.732 30.036 36.764 ;
  LAYER M2 ;
        RECT 27.564 36.668 30.036 36.7 ;
  LAYER M2 ;
        RECT 27.564 36.604 30.036 36.636 ;
  LAYER M2 ;
        RECT 27.564 36.54 30.036 36.572 ;
  LAYER M2 ;
        RECT 27.564 36.476 30.036 36.508 ;
  LAYER M2 ;
        RECT 27.564 36.412 30.036 36.444 ;
  LAYER M2 ;
        RECT 27.564 36.348 30.036 36.38 ;
  LAYER M2 ;
        RECT 27.564 36.284 30.036 36.316 ;
  LAYER M2 ;
        RECT 27.564 36.22 30.036 36.252 ;
  LAYER M2 ;
        RECT 27.564 36.156 30.036 36.188 ;
  LAYER M2 ;
        RECT 27.564 36.092 30.036 36.124 ;
  LAYER M2 ;
        RECT 27.564 36.028 30.036 36.06 ;
  LAYER M2 ;
        RECT 27.564 35.964 30.036 35.996 ;
  LAYER M2 ;
        RECT 27.564 35.9 30.036 35.932 ;
  LAYER M2 ;
        RECT 27.564 35.836 30.036 35.868 ;
  LAYER M2 ;
        RECT 27.564 35.772 30.036 35.804 ;
  LAYER M2 ;
        RECT 27.564 35.708 30.036 35.74 ;
  LAYER M2 ;
        RECT 27.564 35.644 30.036 35.676 ;
  LAYER M2 ;
        RECT 27.564 35.58 30.036 35.612 ;
  LAYER M2 ;
        RECT 27.564 35.516 30.036 35.548 ;
  LAYER M2 ;
        RECT 27.564 35.452 30.036 35.484 ;
  LAYER M2 ;
        RECT 27.564 35.388 30.036 35.42 ;
  LAYER M2 ;
        RECT 27.564 35.324 30.036 35.356 ;
  LAYER M2 ;
        RECT 27.564 35.26 30.036 35.292 ;
  LAYER M2 ;
        RECT 27.564 35.196 30.036 35.228 ;
  LAYER M2 ;
        RECT 27.564 35.132 30.036 35.164 ;
  LAYER M2 ;
        RECT 27.564 35.068 30.036 35.1 ;
  LAYER M2 ;
        RECT 27.564 35.004 30.036 35.036 ;
  LAYER M2 ;
        RECT 27.564 34.94 30.036 34.972 ;
  LAYER M2 ;
        RECT 27.564 34.876 30.036 34.908 ;
  LAYER M2 ;
        RECT 27.564 34.812 30.036 34.844 ;
  LAYER M2 ;
        RECT 27.564 34.748 30.036 34.78 ;
  LAYER M2 ;
        RECT 27.564 34.684 30.036 34.716 ;
  LAYER M2 ;
        RECT 27.564 34.62 30.036 34.652 ;
  LAYER M2 ;
        RECT 27.564 34.556 30.036 34.588 ;
  LAYER M3 ;
        RECT 27.584 34.404 27.616 36.912 ;
  LAYER M3 ;
        RECT 27.648 34.404 27.68 36.912 ;
  LAYER M3 ;
        RECT 27.712 34.404 27.744 36.912 ;
  LAYER M3 ;
        RECT 27.776 34.404 27.808 36.912 ;
  LAYER M3 ;
        RECT 27.84 34.404 27.872 36.912 ;
  LAYER M3 ;
        RECT 27.904 34.404 27.936 36.912 ;
  LAYER M3 ;
        RECT 27.968 34.404 28 36.912 ;
  LAYER M3 ;
        RECT 28.032 34.404 28.064 36.912 ;
  LAYER M3 ;
        RECT 28.096 34.404 28.128 36.912 ;
  LAYER M3 ;
        RECT 28.16 34.404 28.192 36.912 ;
  LAYER M3 ;
        RECT 28.224 34.404 28.256 36.912 ;
  LAYER M3 ;
        RECT 28.288 34.404 28.32 36.912 ;
  LAYER M3 ;
        RECT 28.352 34.404 28.384 36.912 ;
  LAYER M3 ;
        RECT 28.416 34.404 28.448 36.912 ;
  LAYER M3 ;
        RECT 28.48 34.404 28.512 36.912 ;
  LAYER M3 ;
        RECT 28.544 34.404 28.576 36.912 ;
  LAYER M3 ;
        RECT 28.608 34.404 28.64 36.912 ;
  LAYER M3 ;
        RECT 28.672 34.404 28.704 36.912 ;
  LAYER M3 ;
        RECT 28.736 34.404 28.768 36.912 ;
  LAYER M3 ;
        RECT 28.8 34.404 28.832 36.912 ;
  LAYER M3 ;
        RECT 28.864 34.404 28.896 36.912 ;
  LAYER M3 ;
        RECT 28.928 34.404 28.96 36.912 ;
  LAYER M3 ;
        RECT 28.992 34.404 29.024 36.912 ;
  LAYER M3 ;
        RECT 29.056 34.404 29.088 36.912 ;
  LAYER M3 ;
        RECT 29.12 34.404 29.152 36.912 ;
  LAYER M3 ;
        RECT 29.184 34.404 29.216 36.912 ;
  LAYER M3 ;
        RECT 29.248 34.404 29.28 36.912 ;
  LAYER M3 ;
        RECT 29.312 34.404 29.344 36.912 ;
  LAYER M3 ;
        RECT 29.376 34.404 29.408 36.912 ;
  LAYER M3 ;
        RECT 29.44 34.404 29.472 36.912 ;
  LAYER M3 ;
        RECT 29.504 34.404 29.536 36.912 ;
  LAYER M3 ;
        RECT 29.568 34.404 29.6 36.912 ;
  LAYER M3 ;
        RECT 29.632 34.404 29.664 36.912 ;
  LAYER M3 ;
        RECT 29.696 34.404 29.728 36.912 ;
  LAYER M3 ;
        RECT 29.76 34.404 29.792 36.912 ;
  LAYER M3 ;
        RECT 29.824 34.404 29.856 36.912 ;
  LAYER M3 ;
        RECT 29.888 34.404 29.92 36.912 ;
  LAYER M3 ;
        RECT 29.984 34.404 30.016 36.912 ;
  LAYER M1 ;
        RECT 27.599 34.44 27.601 36.876 ;
  LAYER M1 ;
        RECT 27.679 34.44 27.681 36.876 ;
  LAYER M1 ;
        RECT 27.759 34.44 27.761 36.876 ;
  LAYER M1 ;
        RECT 27.839 34.44 27.841 36.876 ;
  LAYER M1 ;
        RECT 27.919 34.44 27.921 36.876 ;
  LAYER M1 ;
        RECT 27.999 34.44 28.001 36.876 ;
  LAYER M1 ;
        RECT 28.079 34.44 28.081 36.876 ;
  LAYER M1 ;
        RECT 28.159 34.44 28.161 36.876 ;
  LAYER M1 ;
        RECT 28.239 34.44 28.241 36.876 ;
  LAYER M1 ;
        RECT 28.319 34.44 28.321 36.876 ;
  LAYER M1 ;
        RECT 28.399 34.44 28.401 36.876 ;
  LAYER M1 ;
        RECT 28.479 34.44 28.481 36.876 ;
  LAYER M1 ;
        RECT 28.559 34.44 28.561 36.876 ;
  LAYER M1 ;
        RECT 28.639 34.44 28.641 36.876 ;
  LAYER M1 ;
        RECT 28.719 34.44 28.721 36.876 ;
  LAYER M1 ;
        RECT 28.799 34.44 28.801 36.876 ;
  LAYER M1 ;
        RECT 28.879 34.44 28.881 36.876 ;
  LAYER M1 ;
        RECT 28.959 34.44 28.961 36.876 ;
  LAYER M1 ;
        RECT 29.039 34.44 29.041 36.876 ;
  LAYER M1 ;
        RECT 29.119 34.44 29.121 36.876 ;
  LAYER M1 ;
        RECT 29.199 34.44 29.201 36.876 ;
  LAYER M1 ;
        RECT 29.279 34.44 29.281 36.876 ;
  LAYER M1 ;
        RECT 29.359 34.44 29.361 36.876 ;
  LAYER M1 ;
        RECT 29.439 34.44 29.441 36.876 ;
  LAYER M1 ;
        RECT 29.519 34.44 29.521 36.876 ;
  LAYER M1 ;
        RECT 29.599 34.44 29.601 36.876 ;
  LAYER M1 ;
        RECT 29.679 34.44 29.681 36.876 ;
  LAYER M1 ;
        RECT 29.759 34.44 29.761 36.876 ;
  LAYER M1 ;
        RECT 29.839 34.44 29.841 36.876 ;
  LAYER M1 ;
        RECT 29.919 34.44 29.921 36.876 ;
  LAYER M2 ;
        RECT 27.6 36.875 30 36.877 ;
  LAYER M2 ;
        RECT 27.6 36.791 30 36.793 ;
  LAYER M2 ;
        RECT 27.6 36.707 30 36.709 ;
  LAYER M2 ;
        RECT 27.6 36.623 30 36.625 ;
  LAYER M2 ;
        RECT 27.6 36.539 30 36.541 ;
  LAYER M2 ;
        RECT 27.6 36.455 30 36.457 ;
  LAYER M2 ;
        RECT 27.6 36.371 30 36.373 ;
  LAYER M2 ;
        RECT 27.6 36.287 30 36.289 ;
  LAYER M2 ;
        RECT 27.6 36.203 30 36.205 ;
  LAYER M2 ;
        RECT 27.6 36.119 30 36.121 ;
  LAYER M2 ;
        RECT 27.6 36.035 30 36.037 ;
  LAYER M2 ;
        RECT 27.6 35.951 30 35.953 ;
  LAYER M2 ;
        RECT 27.6 35.8675 30 35.8695 ;
  LAYER M2 ;
        RECT 27.6 35.783 30 35.785 ;
  LAYER M2 ;
        RECT 27.6 35.699 30 35.701 ;
  LAYER M2 ;
        RECT 27.6 35.615 30 35.617 ;
  LAYER M2 ;
        RECT 27.6 35.531 30 35.533 ;
  LAYER M2 ;
        RECT 27.6 35.447 30 35.449 ;
  LAYER M2 ;
        RECT 27.6 35.363 30 35.365 ;
  LAYER M2 ;
        RECT 27.6 35.279 30 35.281 ;
  LAYER M2 ;
        RECT 27.6 35.195 30 35.197 ;
  LAYER M2 ;
        RECT 27.6 35.111 30 35.113 ;
  LAYER M2 ;
        RECT 27.6 35.027 30 35.029 ;
  LAYER M2 ;
        RECT 27.6 34.943 30 34.945 ;
  LAYER M2 ;
        RECT 27.6 34.859 30 34.861 ;
  LAYER M2 ;
        RECT 27.6 34.775 30 34.777 ;
  LAYER M2 ;
        RECT 27.6 34.691 30 34.693 ;
  LAYER M2 ;
        RECT 27.6 34.607 30 34.609 ;
  LAYER M2 ;
        RECT 27.6 34.523 30 34.525 ;
  LAYER M1 ;
        RECT 27.584 31.464 27.616 33.972 ;
  LAYER M1 ;
        RECT 27.648 31.464 27.68 33.972 ;
  LAYER M1 ;
        RECT 27.712 31.464 27.744 33.972 ;
  LAYER M1 ;
        RECT 27.776 31.464 27.808 33.972 ;
  LAYER M1 ;
        RECT 27.84 31.464 27.872 33.972 ;
  LAYER M1 ;
        RECT 27.904 31.464 27.936 33.972 ;
  LAYER M1 ;
        RECT 27.968 31.464 28 33.972 ;
  LAYER M1 ;
        RECT 28.032 31.464 28.064 33.972 ;
  LAYER M1 ;
        RECT 28.096 31.464 28.128 33.972 ;
  LAYER M1 ;
        RECT 28.16 31.464 28.192 33.972 ;
  LAYER M1 ;
        RECT 28.224 31.464 28.256 33.972 ;
  LAYER M1 ;
        RECT 28.288 31.464 28.32 33.972 ;
  LAYER M1 ;
        RECT 28.352 31.464 28.384 33.972 ;
  LAYER M1 ;
        RECT 28.416 31.464 28.448 33.972 ;
  LAYER M1 ;
        RECT 28.48 31.464 28.512 33.972 ;
  LAYER M1 ;
        RECT 28.544 31.464 28.576 33.972 ;
  LAYER M1 ;
        RECT 28.608 31.464 28.64 33.972 ;
  LAYER M1 ;
        RECT 28.672 31.464 28.704 33.972 ;
  LAYER M1 ;
        RECT 28.736 31.464 28.768 33.972 ;
  LAYER M1 ;
        RECT 28.8 31.464 28.832 33.972 ;
  LAYER M1 ;
        RECT 28.864 31.464 28.896 33.972 ;
  LAYER M1 ;
        RECT 28.928 31.464 28.96 33.972 ;
  LAYER M1 ;
        RECT 28.992 31.464 29.024 33.972 ;
  LAYER M1 ;
        RECT 29.056 31.464 29.088 33.972 ;
  LAYER M1 ;
        RECT 29.12 31.464 29.152 33.972 ;
  LAYER M1 ;
        RECT 29.184 31.464 29.216 33.972 ;
  LAYER M1 ;
        RECT 29.248 31.464 29.28 33.972 ;
  LAYER M1 ;
        RECT 29.312 31.464 29.344 33.972 ;
  LAYER M1 ;
        RECT 29.376 31.464 29.408 33.972 ;
  LAYER M1 ;
        RECT 29.44 31.464 29.472 33.972 ;
  LAYER M1 ;
        RECT 29.504 31.464 29.536 33.972 ;
  LAYER M1 ;
        RECT 29.568 31.464 29.6 33.972 ;
  LAYER M1 ;
        RECT 29.632 31.464 29.664 33.972 ;
  LAYER M1 ;
        RECT 29.696 31.464 29.728 33.972 ;
  LAYER M1 ;
        RECT 29.76 31.464 29.792 33.972 ;
  LAYER M1 ;
        RECT 29.824 31.464 29.856 33.972 ;
  LAYER M1 ;
        RECT 29.888 31.464 29.92 33.972 ;
  LAYER M2 ;
        RECT 27.564 33.856 30.036 33.888 ;
  LAYER M2 ;
        RECT 27.564 33.792 30.036 33.824 ;
  LAYER M2 ;
        RECT 27.564 33.728 30.036 33.76 ;
  LAYER M2 ;
        RECT 27.564 33.664 30.036 33.696 ;
  LAYER M2 ;
        RECT 27.564 33.6 30.036 33.632 ;
  LAYER M2 ;
        RECT 27.564 33.536 30.036 33.568 ;
  LAYER M2 ;
        RECT 27.564 33.472 30.036 33.504 ;
  LAYER M2 ;
        RECT 27.564 33.408 30.036 33.44 ;
  LAYER M2 ;
        RECT 27.564 33.344 30.036 33.376 ;
  LAYER M2 ;
        RECT 27.564 33.28 30.036 33.312 ;
  LAYER M2 ;
        RECT 27.564 33.216 30.036 33.248 ;
  LAYER M2 ;
        RECT 27.564 33.152 30.036 33.184 ;
  LAYER M2 ;
        RECT 27.564 33.088 30.036 33.12 ;
  LAYER M2 ;
        RECT 27.564 33.024 30.036 33.056 ;
  LAYER M2 ;
        RECT 27.564 32.96 30.036 32.992 ;
  LAYER M2 ;
        RECT 27.564 32.896 30.036 32.928 ;
  LAYER M2 ;
        RECT 27.564 32.832 30.036 32.864 ;
  LAYER M2 ;
        RECT 27.564 32.768 30.036 32.8 ;
  LAYER M2 ;
        RECT 27.564 32.704 30.036 32.736 ;
  LAYER M2 ;
        RECT 27.564 32.64 30.036 32.672 ;
  LAYER M2 ;
        RECT 27.564 32.576 30.036 32.608 ;
  LAYER M2 ;
        RECT 27.564 32.512 30.036 32.544 ;
  LAYER M2 ;
        RECT 27.564 32.448 30.036 32.48 ;
  LAYER M2 ;
        RECT 27.564 32.384 30.036 32.416 ;
  LAYER M2 ;
        RECT 27.564 32.32 30.036 32.352 ;
  LAYER M2 ;
        RECT 27.564 32.256 30.036 32.288 ;
  LAYER M2 ;
        RECT 27.564 32.192 30.036 32.224 ;
  LAYER M2 ;
        RECT 27.564 32.128 30.036 32.16 ;
  LAYER M2 ;
        RECT 27.564 32.064 30.036 32.096 ;
  LAYER M2 ;
        RECT 27.564 32 30.036 32.032 ;
  LAYER M2 ;
        RECT 27.564 31.936 30.036 31.968 ;
  LAYER M2 ;
        RECT 27.564 31.872 30.036 31.904 ;
  LAYER M2 ;
        RECT 27.564 31.808 30.036 31.84 ;
  LAYER M2 ;
        RECT 27.564 31.744 30.036 31.776 ;
  LAYER M2 ;
        RECT 27.564 31.68 30.036 31.712 ;
  LAYER M2 ;
        RECT 27.564 31.616 30.036 31.648 ;
  LAYER M3 ;
        RECT 27.584 31.464 27.616 33.972 ;
  LAYER M3 ;
        RECT 27.648 31.464 27.68 33.972 ;
  LAYER M3 ;
        RECT 27.712 31.464 27.744 33.972 ;
  LAYER M3 ;
        RECT 27.776 31.464 27.808 33.972 ;
  LAYER M3 ;
        RECT 27.84 31.464 27.872 33.972 ;
  LAYER M3 ;
        RECT 27.904 31.464 27.936 33.972 ;
  LAYER M3 ;
        RECT 27.968 31.464 28 33.972 ;
  LAYER M3 ;
        RECT 28.032 31.464 28.064 33.972 ;
  LAYER M3 ;
        RECT 28.096 31.464 28.128 33.972 ;
  LAYER M3 ;
        RECT 28.16 31.464 28.192 33.972 ;
  LAYER M3 ;
        RECT 28.224 31.464 28.256 33.972 ;
  LAYER M3 ;
        RECT 28.288 31.464 28.32 33.972 ;
  LAYER M3 ;
        RECT 28.352 31.464 28.384 33.972 ;
  LAYER M3 ;
        RECT 28.416 31.464 28.448 33.972 ;
  LAYER M3 ;
        RECT 28.48 31.464 28.512 33.972 ;
  LAYER M3 ;
        RECT 28.544 31.464 28.576 33.972 ;
  LAYER M3 ;
        RECT 28.608 31.464 28.64 33.972 ;
  LAYER M3 ;
        RECT 28.672 31.464 28.704 33.972 ;
  LAYER M3 ;
        RECT 28.736 31.464 28.768 33.972 ;
  LAYER M3 ;
        RECT 28.8 31.464 28.832 33.972 ;
  LAYER M3 ;
        RECT 28.864 31.464 28.896 33.972 ;
  LAYER M3 ;
        RECT 28.928 31.464 28.96 33.972 ;
  LAYER M3 ;
        RECT 28.992 31.464 29.024 33.972 ;
  LAYER M3 ;
        RECT 29.056 31.464 29.088 33.972 ;
  LAYER M3 ;
        RECT 29.12 31.464 29.152 33.972 ;
  LAYER M3 ;
        RECT 29.184 31.464 29.216 33.972 ;
  LAYER M3 ;
        RECT 29.248 31.464 29.28 33.972 ;
  LAYER M3 ;
        RECT 29.312 31.464 29.344 33.972 ;
  LAYER M3 ;
        RECT 29.376 31.464 29.408 33.972 ;
  LAYER M3 ;
        RECT 29.44 31.464 29.472 33.972 ;
  LAYER M3 ;
        RECT 29.504 31.464 29.536 33.972 ;
  LAYER M3 ;
        RECT 29.568 31.464 29.6 33.972 ;
  LAYER M3 ;
        RECT 29.632 31.464 29.664 33.972 ;
  LAYER M3 ;
        RECT 29.696 31.464 29.728 33.972 ;
  LAYER M3 ;
        RECT 29.76 31.464 29.792 33.972 ;
  LAYER M3 ;
        RECT 29.824 31.464 29.856 33.972 ;
  LAYER M3 ;
        RECT 29.888 31.464 29.92 33.972 ;
  LAYER M3 ;
        RECT 29.984 31.464 30.016 33.972 ;
  LAYER M1 ;
        RECT 27.599 31.5 27.601 33.936 ;
  LAYER M1 ;
        RECT 27.679 31.5 27.681 33.936 ;
  LAYER M1 ;
        RECT 27.759 31.5 27.761 33.936 ;
  LAYER M1 ;
        RECT 27.839 31.5 27.841 33.936 ;
  LAYER M1 ;
        RECT 27.919 31.5 27.921 33.936 ;
  LAYER M1 ;
        RECT 27.999 31.5 28.001 33.936 ;
  LAYER M1 ;
        RECT 28.079 31.5 28.081 33.936 ;
  LAYER M1 ;
        RECT 28.159 31.5 28.161 33.936 ;
  LAYER M1 ;
        RECT 28.239 31.5 28.241 33.936 ;
  LAYER M1 ;
        RECT 28.319 31.5 28.321 33.936 ;
  LAYER M1 ;
        RECT 28.399 31.5 28.401 33.936 ;
  LAYER M1 ;
        RECT 28.479 31.5 28.481 33.936 ;
  LAYER M1 ;
        RECT 28.559 31.5 28.561 33.936 ;
  LAYER M1 ;
        RECT 28.639 31.5 28.641 33.936 ;
  LAYER M1 ;
        RECT 28.719 31.5 28.721 33.936 ;
  LAYER M1 ;
        RECT 28.799 31.5 28.801 33.936 ;
  LAYER M1 ;
        RECT 28.879 31.5 28.881 33.936 ;
  LAYER M1 ;
        RECT 28.959 31.5 28.961 33.936 ;
  LAYER M1 ;
        RECT 29.039 31.5 29.041 33.936 ;
  LAYER M1 ;
        RECT 29.119 31.5 29.121 33.936 ;
  LAYER M1 ;
        RECT 29.199 31.5 29.201 33.936 ;
  LAYER M1 ;
        RECT 29.279 31.5 29.281 33.936 ;
  LAYER M1 ;
        RECT 29.359 31.5 29.361 33.936 ;
  LAYER M1 ;
        RECT 29.439 31.5 29.441 33.936 ;
  LAYER M1 ;
        RECT 29.519 31.5 29.521 33.936 ;
  LAYER M1 ;
        RECT 29.599 31.5 29.601 33.936 ;
  LAYER M1 ;
        RECT 29.679 31.5 29.681 33.936 ;
  LAYER M1 ;
        RECT 29.759 31.5 29.761 33.936 ;
  LAYER M1 ;
        RECT 29.839 31.5 29.841 33.936 ;
  LAYER M1 ;
        RECT 29.919 31.5 29.921 33.936 ;
  LAYER M2 ;
        RECT 27.6 33.935 30 33.937 ;
  LAYER M2 ;
        RECT 27.6 33.851 30 33.853 ;
  LAYER M2 ;
        RECT 27.6 33.767 30 33.769 ;
  LAYER M2 ;
        RECT 27.6 33.683 30 33.685 ;
  LAYER M2 ;
        RECT 27.6 33.599 30 33.601 ;
  LAYER M2 ;
        RECT 27.6 33.515 30 33.517 ;
  LAYER M2 ;
        RECT 27.6 33.431 30 33.433 ;
  LAYER M2 ;
        RECT 27.6 33.347 30 33.349 ;
  LAYER M2 ;
        RECT 27.6 33.263 30 33.265 ;
  LAYER M2 ;
        RECT 27.6 33.179 30 33.181 ;
  LAYER M2 ;
        RECT 27.6 33.095 30 33.097 ;
  LAYER M2 ;
        RECT 27.6 33.011 30 33.013 ;
  LAYER M2 ;
        RECT 27.6 32.9275 30 32.9295 ;
  LAYER M2 ;
        RECT 27.6 32.843 30 32.845 ;
  LAYER M2 ;
        RECT 27.6 32.759 30 32.761 ;
  LAYER M2 ;
        RECT 27.6 32.675 30 32.677 ;
  LAYER M2 ;
        RECT 27.6 32.591 30 32.593 ;
  LAYER M2 ;
        RECT 27.6 32.507 30 32.509 ;
  LAYER M2 ;
        RECT 27.6 32.423 30 32.425 ;
  LAYER M2 ;
        RECT 27.6 32.339 30 32.341 ;
  LAYER M2 ;
        RECT 27.6 32.255 30 32.257 ;
  LAYER M2 ;
        RECT 27.6 32.171 30 32.173 ;
  LAYER M2 ;
        RECT 27.6 32.087 30 32.089 ;
  LAYER M2 ;
        RECT 27.6 32.003 30 32.005 ;
  LAYER M2 ;
        RECT 27.6 31.919 30 31.921 ;
  LAYER M2 ;
        RECT 27.6 31.835 30 31.837 ;
  LAYER M2 ;
        RECT 27.6 31.751 30 31.753 ;
  LAYER M2 ;
        RECT 27.6 31.667 30 31.669 ;
  LAYER M2 ;
        RECT 27.6 31.583 30 31.585 ;
  LAYER M1 ;
        RECT 27.584 28.524 27.616 31.032 ;
  LAYER M1 ;
        RECT 27.648 28.524 27.68 31.032 ;
  LAYER M1 ;
        RECT 27.712 28.524 27.744 31.032 ;
  LAYER M1 ;
        RECT 27.776 28.524 27.808 31.032 ;
  LAYER M1 ;
        RECT 27.84 28.524 27.872 31.032 ;
  LAYER M1 ;
        RECT 27.904 28.524 27.936 31.032 ;
  LAYER M1 ;
        RECT 27.968 28.524 28 31.032 ;
  LAYER M1 ;
        RECT 28.032 28.524 28.064 31.032 ;
  LAYER M1 ;
        RECT 28.096 28.524 28.128 31.032 ;
  LAYER M1 ;
        RECT 28.16 28.524 28.192 31.032 ;
  LAYER M1 ;
        RECT 28.224 28.524 28.256 31.032 ;
  LAYER M1 ;
        RECT 28.288 28.524 28.32 31.032 ;
  LAYER M1 ;
        RECT 28.352 28.524 28.384 31.032 ;
  LAYER M1 ;
        RECT 28.416 28.524 28.448 31.032 ;
  LAYER M1 ;
        RECT 28.48 28.524 28.512 31.032 ;
  LAYER M1 ;
        RECT 28.544 28.524 28.576 31.032 ;
  LAYER M1 ;
        RECT 28.608 28.524 28.64 31.032 ;
  LAYER M1 ;
        RECT 28.672 28.524 28.704 31.032 ;
  LAYER M1 ;
        RECT 28.736 28.524 28.768 31.032 ;
  LAYER M1 ;
        RECT 28.8 28.524 28.832 31.032 ;
  LAYER M1 ;
        RECT 28.864 28.524 28.896 31.032 ;
  LAYER M1 ;
        RECT 28.928 28.524 28.96 31.032 ;
  LAYER M1 ;
        RECT 28.992 28.524 29.024 31.032 ;
  LAYER M1 ;
        RECT 29.056 28.524 29.088 31.032 ;
  LAYER M1 ;
        RECT 29.12 28.524 29.152 31.032 ;
  LAYER M1 ;
        RECT 29.184 28.524 29.216 31.032 ;
  LAYER M1 ;
        RECT 29.248 28.524 29.28 31.032 ;
  LAYER M1 ;
        RECT 29.312 28.524 29.344 31.032 ;
  LAYER M1 ;
        RECT 29.376 28.524 29.408 31.032 ;
  LAYER M1 ;
        RECT 29.44 28.524 29.472 31.032 ;
  LAYER M1 ;
        RECT 29.504 28.524 29.536 31.032 ;
  LAYER M1 ;
        RECT 29.568 28.524 29.6 31.032 ;
  LAYER M1 ;
        RECT 29.632 28.524 29.664 31.032 ;
  LAYER M1 ;
        RECT 29.696 28.524 29.728 31.032 ;
  LAYER M1 ;
        RECT 29.76 28.524 29.792 31.032 ;
  LAYER M1 ;
        RECT 29.824 28.524 29.856 31.032 ;
  LAYER M1 ;
        RECT 29.888 28.524 29.92 31.032 ;
  LAYER M2 ;
        RECT 27.564 30.916 30.036 30.948 ;
  LAYER M2 ;
        RECT 27.564 30.852 30.036 30.884 ;
  LAYER M2 ;
        RECT 27.564 30.788 30.036 30.82 ;
  LAYER M2 ;
        RECT 27.564 30.724 30.036 30.756 ;
  LAYER M2 ;
        RECT 27.564 30.66 30.036 30.692 ;
  LAYER M2 ;
        RECT 27.564 30.596 30.036 30.628 ;
  LAYER M2 ;
        RECT 27.564 30.532 30.036 30.564 ;
  LAYER M2 ;
        RECT 27.564 30.468 30.036 30.5 ;
  LAYER M2 ;
        RECT 27.564 30.404 30.036 30.436 ;
  LAYER M2 ;
        RECT 27.564 30.34 30.036 30.372 ;
  LAYER M2 ;
        RECT 27.564 30.276 30.036 30.308 ;
  LAYER M2 ;
        RECT 27.564 30.212 30.036 30.244 ;
  LAYER M2 ;
        RECT 27.564 30.148 30.036 30.18 ;
  LAYER M2 ;
        RECT 27.564 30.084 30.036 30.116 ;
  LAYER M2 ;
        RECT 27.564 30.02 30.036 30.052 ;
  LAYER M2 ;
        RECT 27.564 29.956 30.036 29.988 ;
  LAYER M2 ;
        RECT 27.564 29.892 30.036 29.924 ;
  LAYER M2 ;
        RECT 27.564 29.828 30.036 29.86 ;
  LAYER M2 ;
        RECT 27.564 29.764 30.036 29.796 ;
  LAYER M2 ;
        RECT 27.564 29.7 30.036 29.732 ;
  LAYER M2 ;
        RECT 27.564 29.636 30.036 29.668 ;
  LAYER M2 ;
        RECT 27.564 29.572 30.036 29.604 ;
  LAYER M2 ;
        RECT 27.564 29.508 30.036 29.54 ;
  LAYER M2 ;
        RECT 27.564 29.444 30.036 29.476 ;
  LAYER M2 ;
        RECT 27.564 29.38 30.036 29.412 ;
  LAYER M2 ;
        RECT 27.564 29.316 30.036 29.348 ;
  LAYER M2 ;
        RECT 27.564 29.252 30.036 29.284 ;
  LAYER M2 ;
        RECT 27.564 29.188 30.036 29.22 ;
  LAYER M2 ;
        RECT 27.564 29.124 30.036 29.156 ;
  LAYER M2 ;
        RECT 27.564 29.06 30.036 29.092 ;
  LAYER M2 ;
        RECT 27.564 28.996 30.036 29.028 ;
  LAYER M2 ;
        RECT 27.564 28.932 30.036 28.964 ;
  LAYER M2 ;
        RECT 27.564 28.868 30.036 28.9 ;
  LAYER M2 ;
        RECT 27.564 28.804 30.036 28.836 ;
  LAYER M2 ;
        RECT 27.564 28.74 30.036 28.772 ;
  LAYER M2 ;
        RECT 27.564 28.676 30.036 28.708 ;
  LAYER M3 ;
        RECT 27.584 28.524 27.616 31.032 ;
  LAYER M3 ;
        RECT 27.648 28.524 27.68 31.032 ;
  LAYER M3 ;
        RECT 27.712 28.524 27.744 31.032 ;
  LAYER M3 ;
        RECT 27.776 28.524 27.808 31.032 ;
  LAYER M3 ;
        RECT 27.84 28.524 27.872 31.032 ;
  LAYER M3 ;
        RECT 27.904 28.524 27.936 31.032 ;
  LAYER M3 ;
        RECT 27.968 28.524 28 31.032 ;
  LAYER M3 ;
        RECT 28.032 28.524 28.064 31.032 ;
  LAYER M3 ;
        RECT 28.096 28.524 28.128 31.032 ;
  LAYER M3 ;
        RECT 28.16 28.524 28.192 31.032 ;
  LAYER M3 ;
        RECT 28.224 28.524 28.256 31.032 ;
  LAYER M3 ;
        RECT 28.288 28.524 28.32 31.032 ;
  LAYER M3 ;
        RECT 28.352 28.524 28.384 31.032 ;
  LAYER M3 ;
        RECT 28.416 28.524 28.448 31.032 ;
  LAYER M3 ;
        RECT 28.48 28.524 28.512 31.032 ;
  LAYER M3 ;
        RECT 28.544 28.524 28.576 31.032 ;
  LAYER M3 ;
        RECT 28.608 28.524 28.64 31.032 ;
  LAYER M3 ;
        RECT 28.672 28.524 28.704 31.032 ;
  LAYER M3 ;
        RECT 28.736 28.524 28.768 31.032 ;
  LAYER M3 ;
        RECT 28.8 28.524 28.832 31.032 ;
  LAYER M3 ;
        RECT 28.864 28.524 28.896 31.032 ;
  LAYER M3 ;
        RECT 28.928 28.524 28.96 31.032 ;
  LAYER M3 ;
        RECT 28.992 28.524 29.024 31.032 ;
  LAYER M3 ;
        RECT 29.056 28.524 29.088 31.032 ;
  LAYER M3 ;
        RECT 29.12 28.524 29.152 31.032 ;
  LAYER M3 ;
        RECT 29.184 28.524 29.216 31.032 ;
  LAYER M3 ;
        RECT 29.248 28.524 29.28 31.032 ;
  LAYER M3 ;
        RECT 29.312 28.524 29.344 31.032 ;
  LAYER M3 ;
        RECT 29.376 28.524 29.408 31.032 ;
  LAYER M3 ;
        RECT 29.44 28.524 29.472 31.032 ;
  LAYER M3 ;
        RECT 29.504 28.524 29.536 31.032 ;
  LAYER M3 ;
        RECT 29.568 28.524 29.6 31.032 ;
  LAYER M3 ;
        RECT 29.632 28.524 29.664 31.032 ;
  LAYER M3 ;
        RECT 29.696 28.524 29.728 31.032 ;
  LAYER M3 ;
        RECT 29.76 28.524 29.792 31.032 ;
  LAYER M3 ;
        RECT 29.824 28.524 29.856 31.032 ;
  LAYER M3 ;
        RECT 29.888 28.524 29.92 31.032 ;
  LAYER M3 ;
        RECT 29.984 28.524 30.016 31.032 ;
  LAYER M1 ;
        RECT 27.599 28.56 27.601 30.996 ;
  LAYER M1 ;
        RECT 27.679 28.56 27.681 30.996 ;
  LAYER M1 ;
        RECT 27.759 28.56 27.761 30.996 ;
  LAYER M1 ;
        RECT 27.839 28.56 27.841 30.996 ;
  LAYER M1 ;
        RECT 27.919 28.56 27.921 30.996 ;
  LAYER M1 ;
        RECT 27.999 28.56 28.001 30.996 ;
  LAYER M1 ;
        RECT 28.079 28.56 28.081 30.996 ;
  LAYER M1 ;
        RECT 28.159 28.56 28.161 30.996 ;
  LAYER M1 ;
        RECT 28.239 28.56 28.241 30.996 ;
  LAYER M1 ;
        RECT 28.319 28.56 28.321 30.996 ;
  LAYER M1 ;
        RECT 28.399 28.56 28.401 30.996 ;
  LAYER M1 ;
        RECT 28.479 28.56 28.481 30.996 ;
  LAYER M1 ;
        RECT 28.559 28.56 28.561 30.996 ;
  LAYER M1 ;
        RECT 28.639 28.56 28.641 30.996 ;
  LAYER M1 ;
        RECT 28.719 28.56 28.721 30.996 ;
  LAYER M1 ;
        RECT 28.799 28.56 28.801 30.996 ;
  LAYER M1 ;
        RECT 28.879 28.56 28.881 30.996 ;
  LAYER M1 ;
        RECT 28.959 28.56 28.961 30.996 ;
  LAYER M1 ;
        RECT 29.039 28.56 29.041 30.996 ;
  LAYER M1 ;
        RECT 29.119 28.56 29.121 30.996 ;
  LAYER M1 ;
        RECT 29.199 28.56 29.201 30.996 ;
  LAYER M1 ;
        RECT 29.279 28.56 29.281 30.996 ;
  LAYER M1 ;
        RECT 29.359 28.56 29.361 30.996 ;
  LAYER M1 ;
        RECT 29.439 28.56 29.441 30.996 ;
  LAYER M1 ;
        RECT 29.519 28.56 29.521 30.996 ;
  LAYER M1 ;
        RECT 29.599 28.56 29.601 30.996 ;
  LAYER M1 ;
        RECT 29.679 28.56 29.681 30.996 ;
  LAYER M1 ;
        RECT 29.759 28.56 29.761 30.996 ;
  LAYER M1 ;
        RECT 29.839 28.56 29.841 30.996 ;
  LAYER M1 ;
        RECT 29.919 28.56 29.921 30.996 ;
  LAYER M2 ;
        RECT 27.6 30.995 30 30.997 ;
  LAYER M2 ;
        RECT 27.6 30.911 30 30.913 ;
  LAYER M2 ;
        RECT 27.6 30.827 30 30.829 ;
  LAYER M2 ;
        RECT 27.6 30.743 30 30.745 ;
  LAYER M2 ;
        RECT 27.6 30.659 30 30.661 ;
  LAYER M2 ;
        RECT 27.6 30.575 30 30.577 ;
  LAYER M2 ;
        RECT 27.6 30.491 30 30.493 ;
  LAYER M2 ;
        RECT 27.6 30.407 30 30.409 ;
  LAYER M2 ;
        RECT 27.6 30.323 30 30.325 ;
  LAYER M2 ;
        RECT 27.6 30.239 30 30.241 ;
  LAYER M2 ;
        RECT 27.6 30.155 30 30.157 ;
  LAYER M2 ;
        RECT 27.6 30.071 30 30.073 ;
  LAYER M2 ;
        RECT 27.6 29.9875 30 29.9895 ;
  LAYER M2 ;
        RECT 27.6 29.903 30 29.905 ;
  LAYER M2 ;
        RECT 27.6 29.819 30 29.821 ;
  LAYER M2 ;
        RECT 27.6 29.735 30 29.737 ;
  LAYER M2 ;
        RECT 27.6 29.651 30 29.653 ;
  LAYER M2 ;
        RECT 27.6 29.567 30 29.569 ;
  LAYER M2 ;
        RECT 27.6 29.483 30 29.485 ;
  LAYER M2 ;
        RECT 27.6 29.399 30 29.401 ;
  LAYER M2 ;
        RECT 27.6 29.315 30 29.317 ;
  LAYER M2 ;
        RECT 27.6 29.231 30 29.233 ;
  LAYER M2 ;
        RECT 27.6 29.147 30 29.149 ;
  LAYER M2 ;
        RECT 27.6 29.063 30 29.065 ;
  LAYER M2 ;
        RECT 27.6 28.979 30 28.981 ;
  LAYER M2 ;
        RECT 27.6 28.895 30 28.897 ;
  LAYER M2 ;
        RECT 27.6 28.811 30 28.813 ;
  LAYER M2 ;
        RECT 27.6 28.727 30 28.729 ;
  LAYER M2 ;
        RECT 27.6 28.643 30 28.645 ;
  LAYER M1 ;
        RECT 27.584 25.584 27.616 28.092 ;
  LAYER M1 ;
        RECT 27.648 25.584 27.68 28.092 ;
  LAYER M1 ;
        RECT 27.712 25.584 27.744 28.092 ;
  LAYER M1 ;
        RECT 27.776 25.584 27.808 28.092 ;
  LAYER M1 ;
        RECT 27.84 25.584 27.872 28.092 ;
  LAYER M1 ;
        RECT 27.904 25.584 27.936 28.092 ;
  LAYER M1 ;
        RECT 27.968 25.584 28 28.092 ;
  LAYER M1 ;
        RECT 28.032 25.584 28.064 28.092 ;
  LAYER M1 ;
        RECT 28.096 25.584 28.128 28.092 ;
  LAYER M1 ;
        RECT 28.16 25.584 28.192 28.092 ;
  LAYER M1 ;
        RECT 28.224 25.584 28.256 28.092 ;
  LAYER M1 ;
        RECT 28.288 25.584 28.32 28.092 ;
  LAYER M1 ;
        RECT 28.352 25.584 28.384 28.092 ;
  LAYER M1 ;
        RECT 28.416 25.584 28.448 28.092 ;
  LAYER M1 ;
        RECT 28.48 25.584 28.512 28.092 ;
  LAYER M1 ;
        RECT 28.544 25.584 28.576 28.092 ;
  LAYER M1 ;
        RECT 28.608 25.584 28.64 28.092 ;
  LAYER M1 ;
        RECT 28.672 25.584 28.704 28.092 ;
  LAYER M1 ;
        RECT 28.736 25.584 28.768 28.092 ;
  LAYER M1 ;
        RECT 28.8 25.584 28.832 28.092 ;
  LAYER M1 ;
        RECT 28.864 25.584 28.896 28.092 ;
  LAYER M1 ;
        RECT 28.928 25.584 28.96 28.092 ;
  LAYER M1 ;
        RECT 28.992 25.584 29.024 28.092 ;
  LAYER M1 ;
        RECT 29.056 25.584 29.088 28.092 ;
  LAYER M1 ;
        RECT 29.12 25.584 29.152 28.092 ;
  LAYER M1 ;
        RECT 29.184 25.584 29.216 28.092 ;
  LAYER M1 ;
        RECT 29.248 25.584 29.28 28.092 ;
  LAYER M1 ;
        RECT 29.312 25.584 29.344 28.092 ;
  LAYER M1 ;
        RECT 29.376 25.584 29.408 28.092 ;
  LAYER M1 ;
        RECT 29.44 25.584 29.472 28.092 ;
  LAYER M1 ;
        RECT 29.504 25.584 29.536 28.092 ;
  LAYER M1 ;
        RECT 29.568 25.584 29.6 28.092 ;
  LAYER M1 ;
        RECT 29.632 25.584 29.664 28.092 ;
  LAYER M1 ;
        RECT 29.696 25.584 29.728 28.092 ;
  LAYER M1 ;
        RECT 29.76 25.584 29.792 28.092 ;
  LAYER M1 ;
        RECT 29.824 25.584 29.856 28.092 ;
  LAYER M1 ;
        RECT 29.888 25.584 29.92 28.092 ;
  LAYER M2 ;
        RECT 27.564 27.976 30.036 28.008 ;
  LAYER M2 ;
        RECT 27.564 27.912 30.036 27.944 ;
  LAYER M2 ;
        RECT 27.564 27.848 30.036 27.88 ;
  LAYER M2 ;
        RECT 27.564 27.784 30.036 27.816 ;
  LAYER M2 ;
        RECT 27.564 27.72 30.036 27.752 ;
  LAYER M2 ;
        RECT 27.564 27.656 30.036 27.688 ;
  LAYER M2 ;
        RECT 27.564 27.592 30.036 27.624 ;
  LAYER M2 ;
        RECT 27.564 27.528 30.036 27.56 ;
  LAYER M2 ;
        RECT 27.564 27.464 30.036 27.496 ;
  LAYER M2 ;
        RECT 27.564 27.4 30.036 27.432 ;
  LAYER M2 ;
        RECT 27.564 27.336 30.036 27.368 ;
  LAYER M2 ;
        RECT 27.564 27.272 30.036 27.304 ;
  LAYER M2 ;
        RECT 27.564 27.208 30.036 27.24 ;
  LAYER M2 ;
        RECT 27.564 27.144 30.036 27.176 ;
  LAYER M2 ;
        RECT 27.564 27.08 30.036 27.112 ;
  LAYER M2 ;
        RECT 27.564 27.016 30.036 27.048 ;
  LAYER M2 ;
        RECT 27.564 26.952 30.036 26.984 ;
  LAYER M2 ;
        RECT 27.564 26.888 30.036 26.92 ;
  LAYER M2 ;
        RECT 27.564 26.824 30.036 26.856 ;
  LAYER M2 ;
        RECT 27.564 26.76 30.036 26.792 ;
  LAYER M2 ;
        RECT 27.564 26.696 30.036 26.728 ;
  LAYER M2 ;
        RECT 27.564 26.632 30.036 26.664 ;
  LAYER M2 ;
        RECT 27.564 26.568 30.036 26.6 ;
  LAYER M2 ;
        RECT 27.564 26.504 30.036 26.536 ;
  LAYER M2 ;
        RECT 27.564 26.44 30.036 26.472 ;
  LAYER M2 ;
        RECT 27.564 26.376 30.036 26.408 ;
  LAYER M2 ;
        RECT 27.564 26.312 30.036 26.344 ;
  LAYER M2 ;
        RECT 27.564 26.248 30.036 26.28 ;
  LAYER M2 ;
        RECT 27.564 26.184 30.036 26.216 ;
  LAYER M2 ;
        RECT 27.564 26.12 30.036 26.152 ;
  LAYER M2 ;
        RECT 27.564 26.056 30.036 26.088 ;
  LAYER M2 ;
        RECT 27.564 25.992 30.036 26.024 ;
  LAYER M2 ;
        RECT 27.564 25.928 30.036 25.96 ;
  LAYER M2 ;
        RECT 27.564 25.864 30.036 25.896 ;
  LAYER M2 ;
        RECT 27.564 25.8 30.036 25.832 ;
  LAYER M2 ;
        RECT 27.564 25.736 30.036 25.768 ;
  LAYER M3 ;
        RECT 27.584 25.584 27.616 28.092 ;
  LAYER M3 ;
        RECT 27.648 25.584 27.68 28.092 ;
  LAYER M3 ;
        RECT 27.712 25.584 27.744 28.092 ;
  LAYER M3 ;
        RECT 27.776 25.584 27.808 28.092 ;
  LAYER M3 ;
        RECT 27.84 25.584 27.872 28.092 ;
  LAYER M3 ;
        RECT 27.904 25.584 27.936 28.092 ;
  LAYER M3 ;
        RECT 27.968 25.584 28 28.092 ;
  LAYER M3 ;
        RECT 28.032 25.584 28.064 28.092 ;
  LAYER M3 ;
        RECT 28.096 25.584 28.128 28.092 ;
  LAYER M3 ;
        RECT 28.16 25.584 28.192 28.092 ;
  LAYER M3 ;
        RECT 28.224 25.584 28.256 28.092 ;
  LAYER M3 ;
        RECT 28.288 25.584 28.32 28.092 ;
  LAYER M3 ;
        RECT 28.352 25.584 28.384 28.092 ;
  LAYER M3 ;
        RECT 28.416 25.584 28.448 28.092 ;
  LAYER M3 ;
        RECT 28.48 25.584 28.512 28.092 ;
  LAYER M3 ;
        RECT 28.544 25.584 28.576 28.092 ;
  LAYER M3 ;
        RECT 28.608 25.584 28.64 28.092 ;
  LAYER M3 ;
        RECT 28.672 25.584 28.704 28.092 ;
  LAYER M3 ;
        RECT 28.736 25.584 28.768 28.092 ;
  LAYER M3 ;
        RECT 28.8 25.584 28.832 28.092 ;
  LAYER M3 ;
        RECT 28.864 25.584 28.896 28.092 ;
  LAYER M3 ;
        RECT 28.928 25.584 28.96 28.092 ;
  LAYER M3 ;
        RECT 28.992 25.584 29.024 28.092 ;
  LAYER M3 ;
        RECT 29.056 25.584 29.088 28.092 ;
  LAYER M3 ;
        RECT 29.12 25.584 29.152 28.092 ;
  LAYER M3 ;
        RECT 29.184 25.584 29.216 28.092 ;
  LAYER M3 ;
        RECT 29.248 25.584 29.28 28.092 ;
  LAYER M3 ;
        RECT 29.312 25.584 29.344 28.092 ;
  LAYER M3 ;
        RECT 29.376 25.584 29.408 28.092 ;
  LAYER M3 ;
        RECT 29.44 25.584 29.472 28.092 ;
  LAYER M3 ;
        RECT 29.504 25.584 29.536 28.092 ;
  LAYER M3 ;
        RECT 29.568 25.584 29.6 28.092 ;
  LAYER M3 ;
        RECT 29.632 25.584 29.664 28.092 ;
  LAYER M3 ;
        RECT 29.696 25.584 29.728 28.092 ;
  LAYER M3 ;
        RECT 29.76 25.584 29.792 28.092 ;
  LAYER M3 ;
        RECT 29.824 25.584 29.856 28.092 ;
  LAYER M3 ;
        RECT 29.888 25.584 29.92 28.092 ;
  LAYER M3 ;
        RECT 29.984 25.584 30.016 28.092 ;
  LAYER M1 ;
        RECT 27.599 25.62 27.601 28.056 ;
  LAYER M1 ;
        RECT 27.679 25.62 27.681 28.056 ;
  LAYER M1 ;
        RECT 27.759 25.62 27.761 28.056 ;
  LAYER M1 ;
        RECT 27.839 25.62 27.841 28.056 ;
  LAYER M1 ;
        RECT 27.919 25.62 27.921 28.056 ;
  LAYER M1 ;
        RECT 27.999 25.62 28.001 28.056 ;
  LAYER M1 ;
        RECT 28.079 25.62 28.081 28.056 ;
  LAYER M1 ;
        RECT 28.159 25.62 28.161 28.056 ;
  LAYER M1 ;
        RECT 28.239 25.62 28.241 28.056 ;
  LAYER M1 ;
        RECT 28.319 25.62 28.321 28.056 ;
  LAYER M1 ;
        RECT 28.399 25.62 28.401 28.056 ;
  LAYER M1 ;
        RECT 28.479 25.62 28.481 28.056 ;
  LAYER M1 ;
        RECT 28.559 25.62 28.561 28.056 ;
  LAYER M1 ;
        RECT 28.639 25.62 28.641 28.056 ;
  LAYER M1 ;
        RECT 28.719 25.62 28.721 28.056 ;
  LAYER M1 ;
        RECT 28.799 25.62 28.801 28.056 ;
  LAYER M1 ;
        RECT 28.879 25.62 28.881 28.056 ;
  LAYER M1 ;
        RECT 28.959 25.62 28.961 28.056 ;
  LAYER M1 ;
        RECT 29.039 25.62 29.041 28.056 ;
  LAYER M1 ;
        RECT 29.119 25.62 29.121 28.056 ;
  LAYER M1 ;
        RECT 29.199 25.62 29.201 28.056 ;
  LAYER M1 ;
        RECT 29.279 25.62 29.281 28.056 ;
  LAYER M1 ;
        RECT 29.359 25.62 29.361 28.056 ;
  LAYER M1 ;
        RECT 29.439 25.62 29.441 28.056 ;
  LAYER M1 ;
        RECT 29.519 25.62 29.521 28.056 ;
  LAYER M1 ;
        RECT 29.599 25.62 29.601 28.056 ;
  LAYER M1 ;
        RECT 29.679 25.62 29.681 28.056 ;
  LAYER M1 ;
        RECT 29.759 25.62 29.761 28.056 ;
  LAYER M1 ;
        RECT 29.839 25.62 29.841 28.056 ;
  LAYER M1 ;
        RECT 29.919 25.62 29.921 28.056 ;
  LAYER M2 ;
        RECT 27.6 28.055 30 28.057 ;
  LAYER M2 ;
        RECT 27.6 27.971 30 27.973 ;
  LAYER M2 ;
        RECT 27.6 27.887 30 27.889 ;
  LAYER M2 ;
        RECT 27.6 27.803 30 27.805 ;
  LAYER M2 ;
        RECT 27.6 27.719 30 27.721 ;
  LAYER M2 ;
        RECT 27.6 27.635 30 27.637 ;
  LAYER M2 ;
        RECT 27.6 27.551 30 27.553 ;
  LAYER M2 ;
        RECT 27.6 27.467 30 27.469 ;
  LAYER M2 ;
        RECT 27.6 27.383 30 27.385 ;
  LAYER M2 ;
        RECT 27.6 27.299 30 27.301 ;
  LAYER M2 ;
        RECT 27.6 27.215 30 27.217 ;
  LAYER M2 ;
        RECT 27.6 27.131 30 27.133 ;
  LAYER M2 ;
        RECT 27.6 27.0475 30 27.0495 ;
  LAYER M2 ;
        RECT 27.6 26.963 30 26.965 ;
  LAYER M2 ;
        RECT 27.6 26.879 30 26.881 ;
  LAYER M2 ;
        RECT 27.6 26.795 30 26.797 ;
  LAYER M2 ;
        RECT 27.6 26.711 30 26.713 ;
  LAYER M2 ;
        RECT 27.6 26.627 30 26.629 ;
  LAYER M2 ;
        RECT 27.6 26.543 30 26.545 ;
  LAYER M2 ;
        RECT 27.6 26.459 30 26.461 ;
  LAYER M2 ;
        RECT 27.6 26.375 30 26.377 ;
  LAYER M2 ;
        RECT 27.6 26.291 30 26.293 ;
  LAYER M2 ;
        RECT 27.6 26.207 30 26.209 ;
  LAYER M2 ;
        RECT 27.6 26.123 30 26.125 ;
  LAYER M2 ;
        RECT 27.6 26.039 30 26.041 ;
  LAYER M2 ;
        RECT 27.6 25.955 30 25.957 ;
  LAYER M2 ;
        RECT 27.6 25.871 30 25.873 ;
  LAYER M2 ;
        RECT 27.6 25.787 30 25.789 ;
  LAYER M2 ;
        RECT 27.6 25.703 30 25.705 ;
  LAYER M1 ;
        RECT 27.584 22.644 27.616 25.152 ;
  LAYER M1 ;
        RECT 27.648 22.644 27.68 25.152 ;
  LAYER M1 ;
        RECT 27.712 22.644 27.744 25.152 ;
  LAYER M1 ;
        RECT 27.776 22.644 27.808 25.152 ;
  LAYER M1 ;
        RECT 27.84 22.644 27.872 25.152 ;
  LAYER M1 ;
        RECT 27.904 22.644 27.936 25.152 ;
  LAYER M1 ;
        RECT 27.968 22.644 28 25.152 ;
  LAYER M1 ;
        RECT 28.032 22.644 28.064 25.152 ;
  LAYER M1 ;
        RECT 28.096 22.644 28.128 25.152 ;
  LAYER M1 ;
        RECT 28.16 22.644 28.192 25.152 ;
  LAYER M1 ;
        RECT 28.224 22.644 28.256 25.152 ;
  LAYER M1 ;
        RECT 28.288 22.644 28.32 25.152 ;
  LAYER M1 ;
        RECT 28.352 22.644 28.384 25.152 ;
  LAYER M1 ;
        RECT 28.416 22.644 28.448 25.152 ;
  LAYER M1 ;
        RECT 28.48 22.644 28.512 25.152 ;
  LAYER M1 ;
        RECT 28.544 22.644 28.576 25.152 ;
  LAYER M1 ;
        RECT 28.608 22.644 28.64 25.152 ;
  LAYER M1 ;
        RECT 28.672 22.644 28.704 25.152 ;
  LAYER M1 ;
        RECT 28.736 22.644 28.768 25.152 ;
  LAYER M1 ;
        RECT 28.8 22.644 28.832 25.152 ;
  LAYER M1 ;
        RECT 28.864 22.644 28.896 25.152 ;
  LAYER M1 ;
        RECT 28.928 22.644 28.96 25.152 ;
  LAYER M1 ;
        RECT 28.992 22.644 29.024 25.152 ;
  LAYER M1 ;
        RECT 29.056 22.644 29.088 25.152 ;
  LAYER M1 ;
        RECT 29.12 22.644 29.152 25.152 ;
  LAYER M1 ;
        RECT 29.184 22.644 29.216 25.152 ;
  LAYER M1 ;
        RECT 29.248 22.644 29.28 25.152 ;
  LAYER M1 ;
        RECT 29.312 22.644 29.344 25.152 ;
  LAYER M1 ;
        RECT 29.376 22.644 29.408 25.152 ;
  LAYER M1 ;
        RECT 29.44 22.644 29.472 25.152 ;
  LAYER M1 ;
        RECT 29.504 22.644 29.536 25.152 ;
  LAYER M1 ;
        RECT 29.568 22.644 29.6 25.152 ;
  LAYER M1 ;
        RECT 29.632 22.644 29.664 25.152 ;
  LAYER M1 ;
        RECT 29.696 22.644 29.728 25.152 ;
  LAYER M1 ;
        RECT 29.76 22.644 29.792 25.152 ;
  LAYER M1 ;
        RECT 29.824 22.644 29.856 25.152 ;
  LAYER M1 ;
        RECT 29.888 22.644 29.92 25.152 ;
  LAYER M2 ;
        RECT 27.564 25.036 30.036 25.068 ;
  LAYER M2 ;
        RECT 27.564 24.972 30.036 25.004 ;
  LAYER M2 ;
        RECT 27.564 24.908 30.036 24.94 ;
  LAYER M2 ;
        RECT 27.564 24.844 30.036 24.876 ;
  LAYER M2 ;
        RECT 27.564 24.78 30.036 24.812 ;
  LAYER M2 ;
        RECT 27.564 24.716 30.036 24.748 ;
  LAYER M2 ;
        RECT 27.564 24.652 30.036 24.684 ;
  LAYER M2 ;
        RECT 27.564 24.588 30.036 24.62 ;
  LAYER M2 ;
        RECT 27.564 24.524 30.036 24.556 ;
  LAYER M2 ;
        RECT 27.564 24.46 30.036 24.492 ;
  LAYER M2 ;
        RECT 27.564 24.396 30.036 24.428 ;
  LAYER M2 ;
        RECT 27.564 24.332 30.036 24.364 ;
  LAYER M2 ;
        RECT 27.564 24.268 30.036 24.3 ;
  LAYER M2 ;
        RECT 27.564 24.204 30.036 24.236 ;
  LAYER M2 ;
        RECT 27.564 24.14 30.036 24.172 ;
  LAYER M2 ;
        RECT 27.564 24.076 30.036 24.108 ;
  LAYER M2 ;
        RECT 27.564 24.012 30.036 24.044 ;
  LAYER M2 ;
        RECT 27.564 23.948 30.036 23.98 ;
  LAYER M2 ;
        RECT 27.564 23.884 30.036 23.916 ;
  LAYER M2 ;
        RECT 27.564 23.82 30.036 23.852 ;
  LAYER M2 ;
        RECT 27.564 23.756 30.036 23.788 ;
  LAYER M2 ;
        RECT 27.564 23.692 30.036 23.724 ;
  LAYER M2 ;
        RECT 27.564 23.628 30.036 23.66 ;
  LAYER M2 ;
        RECT 27.564 23.564 30.036 23.596 ;
  LAYER M2 ;
        RECT 27.564 23.5 30.036 23.532 ;
  LAYER M2 ;
        RECT 27.564 23.436 30.036 23.468 ;
  LAYER M2 ;
        RECT 27.564 23.372 30.036 23.404 ;
  LAYER M2 ;
        RECT 27.564 23.308 30.036 23.34 ;
  LAYER M2 ;
        RECT 27.564 23.244 30.036 23.276 ;
  LAYER M2 ;
        RECT 27.564 23.18 30.036 23.212 ;
  LAYER M2 ;
        RECT 27.564 23.116 30.036 23.148 ;
  LAYER M2 ;
        RECT 27.564 23.052 30.036 23.084 ;
  LAYER M2 ;
        RECT 27.564 22.988 30.036 23.02 ;
  LAYER M2 ;
        RECT 27.564 22.924 30.036 22.956 ;
  LAYER M2 ;
        RECT 27.564 22.86 30.036 22.892 ;
  LAYER M2 ;
        RECT 27.564 22.796 30.036 22.828 ;
  LAYER M3 ;
        RECT 27.584 22.644 27.616 25.152 ;
  LAYER M3 ;
        RECT 27.648 22.644 27.68 25.152 ;
  LAYER M3 ;
        RECT 27.712 22.644 27.744 25.152 ;
  LAYER M3 ;
        RECT 27.776 22.644 27.808 25.152 ;
  LAYER M3 ;
        RECT 27.84 22.644 27.872 25.152 ;
  LAYER M3 ;
        RECT 27.904 22.644 27.936 25.152 ;
  LAYER M3 ;
        RECT 27.968 22.644 28 25.152 ;
  LAYER M3 ;
        RECT 28.032 22.644 28.064 25.152 ;
  LAYER M3 ;
        RECT 28.096 22.644 28.128 25.152 ;
  LAYER M3 ;
        RECT 28.16 22.644 28.192 25.152 ;
  LAYER M3 ;
        RECT 28.224 22.644 28.256 25.152 ;
  LAYER M3 ;
        RECT 28.288 22.644 28.32 25.152 ;
  LAYER M3 ;
        RECT 28.352 22.644 28.384 25.152 ;
  LAYER M3 ;
        RECT 28.416 22.644 28.448 25.152 ;
  LAYER M3 ;
        RECT 28.48 22.644 28.512 25.152 ;
  LAYER M3 ;
        RECT 28.544 22.644 28.576 25.152 ;
  LAYER M3 ;
        RECT 28.608 22.644 28.64 25.152 ;
  LAYER M3 ;
        RECT 28.672 22.644 28.704 25.152 ;
  LAYER M3 ;
        RECT 28.736 22.644 28.768 25.152 ;
  LAYER M3 ;
        RECT 28.8 22.644 28.832 25.152 ;
  LAYER M3 ;
        RECT 28.864 22.644 28.896 25.152 ;
  LAYER M3 ;
        RECT 28.928 22.644 28.96 25.152 ;
  LAYER M3 ;
        RECT 28.992 22.644 29.024 25.152 ;
  LAYER M3 ;
        RECT 29.056 22.644 29.088 25.152 ;
  LAYER M3 ;
        RECT 29.12 22.644 29.152 25.152 ;
  LAYER M3 ;
        RECT 29.184 22.644 29.216 25.152 ;
  LAYER M3 ;
        RECT 29.248 22.644 29.28 25.152 ;
  LAYER M3 ;
        RECT 29.312 22.644 29.344 25.152 ;
  LAYER M3 ;
        RECT 29.376 22.644 29.408 25.152 ;
  LAYER M3 ;
        RECT 29.44 22.644 29.472 25.152 ;
  LAYER M3 ;
        RECT 29.504 22.644 29.536 25.152 ;
  LAYER M3 ;
        RECT 29.568 22.644 29.6 25.152 ;
  LAYER M3 ;
        RECT 29.632 22.644 29.664 25.152 ;
  LAYER M3 ;
        RECT 29.696 22.644 29.728 25.152 ;
  LAYER M3 ;
        RECT 29.76 22.644 29.792 25.152 ;
  LAYER M3 ;
        RECT 29.824 22.644 29.856 25.152 ;
  LAYER M3 ;
        RECT 29.888 22.644 29.92 25.152 ;
  LAYER M3 ;
        RECT 29.984 22.644 30.016 25.152 ;
  LAYER M1 ;
        RECT 27.599 22.68 27.601 25.116 ;
  LAYER M1 ;
        RECT 27.679 22.68 27.681 25.116 ;
  LAYER M1 ;
        RECT 27.759 22.68 27.761 25.116 ;
  LAYER M1 ;
        RECT 27.839 22.68 27.841 25.116 ;
  LAYER M1 ;
        RECT 27.919 22.68 27.921 25.116 ;
  LAYER M1 ;
        RECT 27.999 22.68 28.001 25.116 ;
  LAYER M1 ;
        RECT 28.079 22.68 28.081 25.116 ;
  LAYER M1 ;
        RECT 28.159 22.68 28.161 25.116 ;
  LAYER M1 ;
        RECT 28.239 22.68 28.241 25.116 ;
  LAYER M1 ;
        RECT 28.319 22.68 28.321 25.116 ;
  LAYER M1 ;
        RECT 28.399 22.68 28.401 25.116 ;
  LAYER M1 ;
        RECT 28.479 22.68 28.481 25.116 ;
  LAYER M1 ;
        RECT 28.559 22.68 28.561 25.116 ;
  LAYER M1 ;
        RECT 28.639 22.68 28.641 25.116 ;
  LAYER M1 ;
        RECT 28.719 22.68 28.721 25.116 ;
  LAYER M1 ;
        RECT 28.799 22.68 28.801 25.116 ;
  LAYER M1 ;
        RECT 28.879 22.68 28.881 25.116 ;
  LAYER M1 ;
        RECT 28.959 22.68 28.961 25.116 ;
  LAYER M1 ;
        RECT 29.039 22.68 29.041 25.116 ;
  LAYER M1 ;
        RECT 29.119 22.68 29.121 25.116 ;
  LAYER M1 ;
        RECT 29.199 22.68 29.201 25.116 ;
  LAYER M1 ;
        RECT 29.279 22.68 29.281 25.116 ;
  LAYER M1 ;
        RECT 29.359 22.68 29.361 25.116 ;
  LAYER M1 ;
        RECT 29.439 22.68 29.441 25.116 ;
  LAYER M1 ;
        RECT 29.519 22.68 29.521 25.116 ;
  LAYER M1 ;
        RECT 29.599 22.68 29.601 25.116 ;
  LAYER M1 ;
        RECT 29.679 22.68 29.681 25.116 ;
  LAYER M1 ;
        RECT 29.759 22.68 29.761 25.116 ;
  LAYER M1 ;
        RECT 29.839 22.68 29.841 25.116 ;
  LAYER M1 ;
        RECT 29.919 22.68 29.921 25.116 ;
  LAYER M2 ;
        RECT 27.6 25.115 30 25.117 ;
  LAYER M2 ;
        RECT 27.6 25.031 30 25.033 ;
  LAYER M2 ;
        RECT 27.6 24.947 30 24.949 ;
  LAYER M2 ;
        RECT 27.6 24.863 30 24.865 ;
  LAYER M2 ;
        RECT 27.6 24.779 30 24.781 ;
  LAYER M2 ;
        RECT 27.6 24.695 30 24.697 ;
  LAYER M2 ;
        RECT 27.6 24.611 30 24.613 ;
  LAYER M2 ;
        RECT 27.6 24.527 30 24.529 ;
  LAYER M2 ;
        RECT 27.6 24.443 30 24.445 ;
  LAYER M2 ;
        RECT 27.6 24.359 30 24.361 ;
  LAYER M2 ;
        RECT 27.6 24.275 30 24.277 ;
  LAYER M2 ;
        RECT 27.6 24.191 30 24.193 ;
  LAYER M2 ;
        RECT 27.6 24.1075 30 24.1095 ;
  LAYER M2 ;
        RECT 27.6 24.023 30 24.025 ;
  LAYER M2 ;
        RECT 27.6 23.939 30 23.941 ;
  LAYER M2 ;
        RECT 27.6 23.855 30 23.857 ;
  LAYER M2 ;
        RECT 27.6 23.771 30 23.773 ;
  LAYER M2 ;
        RECT 27.6 23.687 30 23.689 ;
  LAYER M2 ;
        RECT 27.6 23.603 30 23.605 ;
  LAYER M2 ;
        RECT 27.6 23.519 30 23.521 ;
  LAYER M2 ;
        RECT 27.6 23.435 30 23.437 ;
  LAYER M2 ;
        RECT 27.6 23.351 30 23.353 ;
  LAYER M2 ;
        RECT 27.6 23.267 30 23.269 ;
  LAYER M2 ;
        RECT 27.6 23.183 30 23.185 ;
  LAYER M2 ;
        RECT 27.6 23.099 30 23.101 ;
  LAYER M2 ;
        RECT 27.6 23.015 30 23.017 ;
  LAYER M2 ;
        RECT 27.6 22.931 30 22.933 ;
  LAYER M2 ;
        RECT 27.6 22.847 30 22.849 ;
  LAYER M2 ;
        RECT 27.6 22.763 30 22.765 ;
  LAYER M1 ;
        RECT 27.584 19.704 27.616 22.212 ;
  LAYER M1 ;
        RECT 27.648 19.704 27.68 22.212 ;
  LAYER M1 ;
        RECT 27.712 19.704 27.744 22.212 ;
  LAYER M1 ;
        RECT 27.776 19.704 27.808 22.212 ;
  LAYER M1 ;
        RECT 27.84 19.704 27.872 22.212 ;
  LAYER M1 ;
        RECT 27.904 19.704 27.936 22.212 ;
  LAYER M1 ;
        RECT 27.968 19.704 28 22.212 ;
  LAYER M1 ;
        RECT 28.032 19.704 28.064 22.212 ;
  LAYER M1 ;
        RECT 28.096 19.704 28.128 22.212 ;
  LAYER M1 ;
        RECT 28.16 19.704 28.192 22.212 ;
  LAYER M1 ;
        RECT 28.224 19.704 28.256 22.212 ;
  LAYER M1 ;
        RECT 28.288 19.704 28.32 22.212 ;
  LAYER M1 ;
        RECT 28.352 19.704 28.384 22.212 ;
  LAYER M1 ;
        RECT 28.416 19.704 28.448 22.212 ;
  LAYER M1 ;
        RECT 28.48 19.704 28.512 22.212 ;
  LAYER M1 ;
        RECT 28.544 19.704 28.576 22.212 ;
  LAYER M1 ;
        RECT 28.608 19.704 28.64 22.212 ;
  LAYER M1 ;
        RECT 28.672 19.704 28.704 22.212 ;
  LAYER M1 ;
        RECT 28.736 19.704 28.768 22.212 ;
  LAYER M1 ;
        RECT 28.8 19.704 28.832 22.212 ;
  LAYER M1 ;
        RECT 28.864 19.704 28.896 22.212 ;
  LAYER M1 ;
        RECT 28.928 19.704 28.96 22.212 ;
  LAYER M1 ;
        RECT 28.992 19.704 29.024 22.212 ;
  LAYER M1 ;
        RECT 29.056 19.704 29.088 22.212 ;
  LAYER M1 ;
        RECT 29.12 19.704 29.152 22.212 ;
  LAYER M1 ;
        RECT 29.184 19.704 29.216 22.212 ;
  LAYER M1 ;
        RECT 29.248 19.704 29.28 22.212 ;
  LAYER M1 ;
        RECT 29.312 19.704 29.344 22.212 ;
  LAYER M1 ;
        RECT 29.376 19.704 29.408 22.212 ;
  LAYER M1 ;
        RECT 29.44 19.704 29.472 22.212 ;
  LAYER M1 ;
        RECT 29.504 19.704 29.536 22.212 ;
  LAYER M1 ;
        RECT 29.568 19.704 29.6 22.212 ;
  LAYER M1 ;
        RECT 29.632 19.704 29.664 22.212 ;
  LAYER M1 ;
        RECT 29.696 19.704 29.728 22.212 ;
  LAYER M1 ;
        RECT 29.76 19.704 29.792 22.212 ;
  LAYER M1 ;
        RECT 29.824 19.704 29.856 22.212 ;
  LAYER M1 ;
        RECT 29.888 19.704 29.92 22.212 ;
  LAYER M2 ;
        RECT 27.564 22.096 30.036 22.128 ;
  LAYER M2 ;
        RECT 27.564 22.032 30.036 22.064 ;
  LAYER M2 ;
        RECT 27.564 21.968 30.036 22 ;
  LAYER M2 ;
        RECT 27.564 21.904 30.036 21.936 ;
  LAYER M2 ;
        RECT 27.564 21.84 30.036 21.872 ;
  LAYER M2 ;
        RECT 27.564 21.776 30.036 21.808 ;
  LAYER M2 ;
        RECT 27.564 21.712 30.036 21.744 ;
  LAYER M2 ;
        RECT 27.564 21.648 30.036 21.68 ;
  LAYER M2 ;
        RECT 27.564 21.584 30.036 21.616 ;
  LAYER M2 ;
        RECT 27.564 21.52 30.036 21.552 ;
  LAYER M2 ;
        RECT 27.564 21.456 30.036 21.488 ;
  LAYER M2 ;
        RECT 27.564 21.392 30.036 21.424 ;
  LAYER M2 ;
        RECT 27.564 21.328 30.036 21.36 ;
  LAYER M2 ;
        RECT 27.564 21.264 30.036 21.296 ;
  LAYER M2 ;
        RECT 27.564 21.2 30.036 21.232 ;
  LAYER M2 ;
        RECT 27.564 21.136 30.036 21.168 ;
  LAYER M2 ;
        RECT 27.564 21.072 30.036 21.104 ;
  LAYER M2 ;
        RECT 27.564 21.008 30.036 21.04 ;
  LAYER M2 ;
        RECT 27.564 20.944 30.036 20.976 ;
  LAYER M2 ;
        RECT 27.564 20.88 30.036 20.912 ;
  LAYER M2 ;
        RECT 27.564 20.816 30.036 20.848 ;
  LAYER M2 ;
        RECT 27.564 20.752 30.036 20.784 ;
  LAYER M2 ;
        RECT 27.564 20.688 30.036 20.72 ;
  LAYER M2 ;
        RECT 27.564 20.624 30.036 20.656 ;
  LAYER M2 ;
        RECT 27.564 20.56 30.036 20.592 ;
  LAYER M2 ;
        RECT 27.564 20.496 30.036 20.528 ;
  LAYER M2 ;
        RECT 27.564 20.432 30.036 20.464 ;
  LAYER M2 ;
        RECT 27.564 20.368 30.036 20.4 ;
  LAYER M2 ;
        RECT 27.564 20.304 30.036 20.336 ;
  LAYER M2 ;
        RECT 27.564 20.24 30.036 20.272 ;
  LAYER M2 ;
        RECT 27.564 20.176 30.036 20.208 ;
  LAYER M2 ;
        RECT 27.564 20.112 30.036 20.144 ;
  LAYER M2 ;
        RECT 27.564 20.048 30.036 20.08 ;
  LAYER M2 ;
        RECT 27.564 19.984 30.036 20.016 ;
  LAYER M2 ;
        RECT 27.564 19.92 30.036 19.952 ;
  LAYER M2 ;
        RECT 27.564 19.856 30.036 19.888 ;
  LAYER M3 ;
        RECT 27.584 19.704 27.616 22.212 ;
  LAYER M3 ;
        RECT 27.648 19.704 27.68 22.212 ;
  LAYER M3 ;
        RECT 27.712 19.704 27.744 22.212 ;
  LAYER M3 ;
        RECT 27.776 19.704 27.808 22.212 ;
  LAYER M3 ;
        RECT 27.84 19.704 27.872 22.212 ;
  LAYER M3 ;
        RECT 27.904 19.704 27.936 22.212 ;
  LAYER M3 ;
        RECT 27.968 19.704 28 22.212 ;
  LAYER M3 ;
        RECT 28.032 19.704 28.064 22.212 ;
  LAYER M3 ;
        RECT 28.096 19.704 28.128 22.212 ;
  LAYER M3 ;
        RECT 28.16 19.704 28.192 22.212 ;
  LAYER M3 ;
        RECT 28.224 19.704 28.256 22.212 ;
  LAYER M3 ;
        RECT 28.288 19.704 28.32 22.212 ;
  LAYER M3 ;
        RECT 28.352 19.704 28.384 22.212 ;
  LAYER M3 ;
        RECT 28.416 19.704 28.448 22.212 ;
  LAYER M3 ;
        RECT 28.48 19.704 28.512 22.212 ;
  LAYER M3 ;
        RECT 28.544 19.704 28.576 22.212 ;
  LAYER M3 ;
        RECT 28.608 19.704 28.64 22.212 ;
  LAYER M3 ;
        RECT 28.672 19.704 28.704 22.212 ;
  LAYER M3 ;
        RECT 28.736 19.704 28.768 22.212 ;
  LAYER M3 ;
        RECT 28.8 19.704 28.832 22.212 ;
  LAYER M3 ;
        RECT 28.864 19.704 28.896 22.212 ;
  LAYER M3 ;
        RECT 28.928 19.704 28.96 22.212 ;
  LAYER M3 ;
        RECT 28.992 19.704 29.024 22.212 ;
  LAYER M3 ;
        RECT 29.056 19.704 29.088 22.212 ;
  LAYER M3 ;
        RECT 29.12 19.704 29.152 22.212 ;
  LAYER M3 ;
        RECT 29.184 19.704 29.216 22.212 ;
  LAYER M3 ;
        RECT 29.248 19.704 29.28 22.212 ;
  LAYER M3 ;
        RECT 29.312 19.704 29.344 22.212 ;
  LAYER M3 ;
        RECT 29.376 19.704 29.408 22.212 ;
  LAYER M3 ;
        RECT 29.44 19.704 29.472 22.212 ;
  LAYER M3 ;
        RECT 29.504 19.704 29.536 22.212 ;
  LAYER M3 ;
        RECT 29.568 19.704 29.6 22.212 ;
  LAYER M3 ;
        RECT 29.632 19.704 29.664 22.212 ;
  LAYER M3 ;
        RECT 29.696 19.704 29.728 22.212 ;
  LAYER M3 ;
        RECT 29.76 19.704 29.792 22.212 ;
  LAYER M3 ;
        RECT 29.824 19.704 29.856 22.212 ;
  LAYER M3 ;
        RECT 29.888 19.704 29.92 22.212 ;
  LAYER M3 ;
        RECT 29.984 19.704 30.016 22.212 ;
  LAYER M1 ;
        RECT 27.599 19.74 27.601 22.176 ;
  LAYER M1 ;
        RECT 27.679 19.74 27.681 22.176 ;
  LAYER M1 ;
        RECT 27.759 19.74 27.761 22.176 ;
  LAYER M1 ;
        RECT 27.839 19.74 27.841 22.176 ;
  LAYER M1 ;
        RECT 27.919 19.74 27.921 22.176 ;
  LAYER M1 ;
        RECT 27.999 19.74 28.001 22.176 ;
  LAYER M1 ;
        RECT 28.079 19.74 28.081 22.176 ;
  LAYER M1 ;
        RECT 28.159 19.74 28.161 22.176 ;
  LAYER M1 ;
        RECT 28.239 19.74 28.241 22.176 ;
  LAYER M1 ;
        RECT 28.319 19.74 28.321 22.176 ;
  LAYER M1 ;
        RECT 28.399 19.74 28.401 22.176 ;
  LAYER M1 ;
        RECT 28.479 19.74 28.481 22.176 ;
  LAYER M1 ;
        RECT 28.559 19.74 28.561 22.176 ;
  LAYER M1 ;
        RECT 28.639 19.74 28.641 22.176 ;
  LAYER M1 ;
        RECT 28.719 19.74 28.721 22.176 ;
  LAYER M1 ;
        RECT 28.799 19.74 28.801 22.176 ;
  LAYER M1 ;
        RECT 28.879 19.74 28.881 22.176 ;
  LAYER M1 ;
        RECT 28.959 19.74 28.961 22.176 ;
  LAYER M1 ;
        RECT 29.039 19.74 29.041 22.176 ;
  LAYER M1 ;
        RECT 29.119 19.74 29.121 22.176 ;
  LAYER M1 ;
        RECT 29.199 19.74 29.201 22.176 ;
  LAYER M1 ;
        RECT 29.279 19.74 29.281 22.176 ;
  LAYER M1 ;
        RECT 29.359 19.74 29.361 22.176 ;
  LAYER M1 ;
        RECT 29.439 19.74 29.441 22.176 ;
  LAYER M1 ;
        RECT 29.519 19.74 29.521 22.176 ;
  LAYER M1 ;
        RECT 29.599 19.74 29.601 22.176 ;
  LAYER M1 ;
        RECT 29.679 19.74 29.681 22.176 ;
  LAYER M1 ;
        RECT 29.759 19.74 29.761 22.176 ;
  LAYER M1 ;
        RECT 29.839 19.74 29.841 22.176 ;
  LAYER M1 ;
        RECT 29.919 19.74 29.921 22.176 ;
  LAYER M2 ;
        RECT 27.6 22.175 30 22.177 ;
  LAYER M2 ;
        RECT 27.6 22.091 30 22.093 ;
  LAYER M2 ;
        RECT 27.6 22.007 30 22.009 ;
  LAYER M2 ;
        RECT 27.6 21.923 30 21.925 ;
  LAYER M2 ;
        RECT 27.6 21.839 30 21.841 ;
  LAYER M2 ;
        RECT 27.6 21.755 30 21.757 ;
  LAYER M2 ;
        RECT 27.6 21.671 30 21.673 ;
  LAYER M2 ;
        RECT 27.6 21.587 30 21.589 ;
  LAYER M2 ;
        RECT 27.6 21.503 30 21.505 ;
  LAYER M2 ;
        RECT 27.6 21.419 30 21.421 ;
  LAYER M2 ;
        RECT 27.6 21.335 30 21.337 ;
  LAYER M2 ;
        RECT 27.6 21.251 30 21.253 ;
  LAYER M2 ;
        RECT 27.6 21.1675 30 21.1695 ;
  LAYER M2 ;
        RECT 27.6 21.083 30 21.085 ;
  LAYER M2 ;
        RECT 27.6 20.999 30 21.001 ;
  LAYER M2 ;
        RECT 27.6 20.915 30 20.917 ;
  LAYER M2 ;
        RECT 27.6 20.831 30 20.833 ;
  LAYER M2 ;
        RECT 27.6 20.747 30 20.749 ;
  LAYER M2 ;
        RECT 27.6 20.663 30 20.665 ;
  LAYER M2 ;
        RECT 27.6 20.579 30 20.581 ;
  LAYER M2 ;
        RECT 27.6 20.495 30 20.497 ;
  LAYER M2 ;
        RECT 27.6 20.411 30 20.413 ;
  LAYER M2 ;
        RECT 27.6 20.327 30 20.329 ;
  LAYER M2 ;
        RECT 27.6 20.243 30 20.245 ;
  LAYER M2 ;
        RECT 27.6 20.159 30 20.161 ;
  LAYER M2 ;
        RECT 27.6 20.075 30 20.077 ;
  LAYER M2 ;
        RECT 27.6 19.991 30 19.993 ;
  LAYER M2 ;
        RECT 27.6 19.907 30 19.909 ;
  LAYER M2 ;
        RECT 27.6 19.823 30 19.825 ;
  END 
END switched_capacitor_filter
