.PARAM wdef=60n
.PARAM minl=20n

.subckt Tristate_buffer vin vout enable VDD VSS

M5 inv_out enable VSS VSS nfet l=minl w=wdef nfin=20
M1 vout vin net26 VSS nfet l=minl w=wdef nfin=20
M0 net26 enable VSS VSS nfet l=minl w=wdef nfin=20
M3 net30 inv_out VDD VDD pfet l=minl w=wdef nfin=20
M4 inv_out enable VDD VDD pfet  l=minl w=wdef nfin=20
M2 vout vin net30 VDD pfet l=minl w=wdef nfin=20
.ends

