
.subckt Sanitized_model3x_MDLL_TOP EN_DLL MD_SAR MD_TRK SCLK0 VDD VSS FRCODE<6> FRCODE<5> FRCODE<4> FRCODE<3> FRCODE<2> FRCODE<1> FRCODE<0> NDIV<5> NDIV<4> NDIV<3> NDIV<2> NDIV<1> NDIV<0> CKOUT
XI0 EN_DLL FR MD_SAR MD_TRK net15 net19 SCLK0 SEL_RST net20 VDD VSS MDLL_CKGEN_V1
XI1 net17 EN_DLL CODE<2> CODE<1> CODE<0> net15 CODE<3> CODE<4> CODE<5> CODE<6> net013 VDD VSS DEL_7b
XI3 CODE<6> CODE<5> CODE<4> CODE<3> CODE<2> CODE<1> CODE<0> COMP EN_DLL FRCODE<6> FRCODE<5> FRCODE<4> FRCODE<3> FRCODE<2> FRCODE<1> FRCODE<0> FR net15 net19 net016<0> net016<1> net016<2> net20 VDD VSS MDLL_LOGIC_VLOG
XI10<131> VDD VSS DCAP8
XI10<130> VDD VSS DCAP8
XI10<129> VDD VSS DCAP8
XI10<128> VDD VSS DCAP8
XI10<127> VDD VSS DCAP8
XI10<126> VDD VSS DCAP8
XI10<125> VDD VSS DCAP8
XI10<124> VDD VSS DCAP8
XI10<123> VDD VSS DCAP8
XI10<122> VDD VSS DCAP8
XI10<121> VDD VSS DCAP8
XI10<120> VDD VSS DCAP8
XI10<119> VDD VSS DCAP8
XI10<118> VDD VSS DCAP8
XI10<117> VDD VSS DCAP8
XI10<116> VDD VSS DCAP8
XI10<115> VDD VSS DCAP8
XI10<114> VDD VSS DCAP8
XI10<113> VDD VSS DCAP8
XI10<112> VDD VSS DCAP8
XI10<111> VDD VSS DCAP8
XI10<110> VDD VSS DCAP8
XI10<109> VDD VSS DCAP8
XI10<108> VDD VSS DCAP8
XI10<107> VDD VSS DCAP8
XI10<106> VDD VSS DCAP8
XI10<105> VDD VSS DCAP8
XI10<104> VDD VSS DCAP8
XI10<103> VDD VSS DCAP8
XI10<102> VDD VSS DCAP8
XI10<101> VDD VSS DCAP8
XI10<100> VDD VSS DCAP8
XI10<99> VDD VSS DCAP8
XI10<98> VDD VSS DCAP8
XI10<97> VDD VSS DCAP8
XI10<96> VDD VSS DCAP8
XI10<95> VDD VSS DCAP8
XI10<94> VDD VSS DCAP8
XI10<93> VDD VSS DCAP8
XI10<92> VDD VSS DCAP8
XI10<91> VDD VSS DCAP8
XI10<90> VDD VSS DCAP8
XI10<89> VDD VSS DCAP8
XI10<88> VDD VSS DCAP8
XI10<87> VDD VSS DCAP8
XI10<86> VDD VSS DCAP8
XI10<85> VDD VSS DCAP8
XI10<84> VDD VSS DCAP8
XI10<83> VDD VSS DCAP8
XI10<82> VDD VSS DCAP8
XI10<81> VDD VSS DCAP8
XI10<80> VDD VSS DCAP8
XI10<79> VDD VSS DCAP8
XI10<78> VDD VSS DCAP8
XI10<77> VDD VSS DCAP8
XI10<76> VDD VSS DCAP8
XI10<75> VDD VSS DCAP8
XI10<74> VDD VSS DCAP8
XI10<73> VDD VSS DCAP8
XI10<72> VDD VSS DCAP8
XI10<71> VDD VSS DCAP8
XI10<70> VDD VSS DCAP8
XI10<69> VDD VSS DCAP8
XI10<68> VDD VSS DCAP8
XI10<67> VDD VSS DCAP8
XI10<66> VDD VSS DCAP8
XI10<65> VDD VSS DCAP8
XI10<64> VDD VSS DCAP8
XI10<63> VDD VSS DCAP8
XI10<62> VDD VSS DCAP8
XI10<61> VDD VSS DCAP8
XI10<60> VDD VSS DCAP8
XI10<59> VDD VSS DCAP8
XI10<58> VDD VSS DCAP8
XI10<57> VDD VSS DCAP8
XI10<56> VDD VSS DCAP8
XI10<55> VDD VSS DCAP8
XI10<54> VDD VSS DCAP8
XI10<53> VDD VSS DCAP8
XI10<52> VDD VSS DCAP8
XI10<51> VDD VSS DCAP8
XI10<50> VDD VSS DCAP8
XI10<49> VDD VSS DCAP8
XI10<48> VDD VSS DCAP8
XI10<47> VDD VSS DCAP8
XI10<46> VDD VSS DCAP8
XI10<45> VDD VSS DCAP8
XI10<44> VDD VSS DCAP8
XI10<43> VDD VSS DCAP8
XI10<42> VDD VSS DCAP8
XI10<41> VDD VSS DCAP8
XI10<40> VDD VSS DCAP8
XI10<39> VDD VSS DCAP8
XI10<38> VDD VSS DCAP8
XI10<37> VDD VSS DCAP8
XI10<36> VDD VSS DCAP8
XI10<35> VDD VSS DCAP8
XI10<34> VDD VSS DCAP8
XI10<33> VDD VSS DCAP8
XI10<32> VDD VSS DCAP8
XI10<31> VDD VSS DCAP8
XI10<30> VDD VSS DCAP8
XI10<29> VDD VSS DCAP8
XI10<28> VDD VSS DCAP8
XI10<27> VDD VSS DCAP8
XI10<26> VDD VSS DCAP8
XI10<25> VDD VSS DCAP8
XI10<24> VDD VSS DCAP8
XI10<23> VDD VSS DCAP8
XI10<22> VDD VSS DCAP8
XI10<21> VDD VSS DCAP8
XI10<20> VDD VSS DCAP8
XI10<19> VDD VSS DCAP8
XI10<18> VDD VSS DCAP8
XI10<17> VDD VSS DCAP8
XI10<16> VDD VSS DCAP8
XI10<15> VDD VSS DCAP8
XI10<14> VDD VSS DCAP8
XI10<13> VDD VSS DCAP8
XI10<12> VDD VSS DCAP8
XI10<11> VDD VSS DCAP8
XI10<10> VDD VSS DCAP8
XI10<9> VDD VSS DCAP8
XI10<8> VDD VSS DCAP8
XI10<7> VDD VSS DCAP8
XI10<6> VDD VSS DCAP8
XI10<5> VDD VSS DCAP8
XI10<4> VDD VSS DCAP8
XI10<3> VDD VSS DCAP8
XI10<2> VDD VSS DCAP8
XI10<1> VDD VSS DCAP8
XI10<0> VDD VSS DCAP8
XI2 net17 NDIV<5> NDIV<4> NDIV<3> NDIV<2> NDIV<1> NDIV<0> net16 SEL_RST VDD VSS SEL_LOGIC_V2
XI8 net16 VDD VSS COMP INVD0
XI7 net17 VDD VSS CKOUT CKBD2
XI16 net16 FR VDD VSS net013 OR2D1
.ends Sanitized_model3x_MDLL_TOP

.subckt MDLL_CKGEN_V1 EN_DLL FREE_RUN MD_SAR MD_TRK REF_CLK SAR_EN SCLK0 SEL_RST TRK_EN
XI9 net31 VDD VSS net17 INVD0
XI40 net042 EN_DLL MD_SAR VDD VSS SAR_EN AN3D2
XI45 SCLK net010 net25 VDD VSS net048 AN3D2
XI25 net010 VDD VSS FREE_RUN INVD1
XI5 net37 VDD VSS net25 INVD1
XI0 MD_SAR MD_TRK VDD VSS net36 NR2D0
XI43 SCLK0 EN_DLL net032 net045 VDD VSS DFND1
XI44 net048 VDD VSS SEL_RST INVD8
XI15 VDD VSS net32 TIEL
XI22 SCLK net30 net27 net14 VDD VSS DFSNQD1
XI21 SCLK net29 net30 net14 VDD VSS DFSNQD1
XI20 SCLK net27 net021 net14 VDD VSS DFSNQD1
XI19 SCLK net34 net33 net14 VDD VSS DFSNQD1
XI18 SCLK net33 net29 net14 VDD VSS DFSNQD1
XI17 SCLK net35 net34 net14 VDD VSS DFSNQD1
XI16 SCLK net32 net35 net14 VDD VSS DFSNQD1
XI24 net36 EN_DLL VDD VSS net010 ND2D0
XI8 EN_DLL VDD VSS net31 DEL015
XI4 SCLK VDD VSS net37 DEL015
XI27 SCLK net021 net042 net026 net14 VDD VSS DFSND1
XI28 net026 EN_DLL VDD VSS TRK_RST AN2D0
XI30 TRK_RST net020 net039 net027 net039 VDD VSS DFCND1
XI29 TRK_RST SCLK net015 net020 net015 VDD VSS DFCND1
XI36 net032 SCLK0 VDD VSS SCLK AN2D2
XI35 SCLK VDD VSS REF_CLK CKBD4
XI38 EN_DLL net17 MD_SAR VDD VSS net14 ND3D3
XI42 net027 net015 MD_TRK VDD VSS TRK_EN AN3D1
.ends MDLL_CKGEN_V1

.subckt INVD0 I ZN
xMMU1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD0

.subckt Switch_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_NMOS_n12_X1_Y1

.subckt Switch_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_PMOS_n12_X1_Y1

.subckt AN3D2 A1 A2 A3 Z
xMM_u3_1_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u6 net13 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u5 net9 A2 net13 VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u4 net5 A1 net9 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_0_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u3 net5 A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_1_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_0_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AN3D2

.subckt INVD1 I ZN
xMMU1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD1

.subckt NR2D0 A1 A2 ZN
xMMI1_M_u3 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 net13 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A1 net13 VDD Switch_PMOS_n12_X1_Y1
.ends NR2D0

.subckt DFND1 CPN D Q QN
xMMI53_M_u2 net63 net100 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI29_M_u2 QN net97 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI4 net24 net67 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55 net97 net67 net100 VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net11 net1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI50 net11 net95 net100 VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u2 net67 net95 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net1 D net24 VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u2 net95 CPN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI56_M_u2 net97 net63 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net9 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 Q net63 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net1 net95 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI53_M_u3 net63 net100 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI54 net97 net95 net100 VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u3 net67 net95 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI43 net60 net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net1 D net53 VDD Switch_PMOS_n12_X1_Y1
xMMI29_M_u3 QN net97 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u3 net95 CPN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 Q net63 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net11 net1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI52 net11 net67 net100 VDD Switch_PMOS_n12_X1_Y1
xMMI56_M_u3 net97 net63 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI45 net1 net67 net60 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net53 net95 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DFND1

.subckt INVD8 I ZN
xMMU1_5_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_0_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_3_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_7_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_4_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_6_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_2_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_0_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_4_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_5_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_3_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_7_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_6_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_2_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD8

.subckt TIEL ZN
xMM_u2 ZN net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u1 net5 VDD VDD VDD DCL_PMOS_n12_X1_Y1
.ends TIEL

.subckt DCL_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends DCL_PMOS_n12_X1_Y1

.subckt DFSNQD1 CP D Q SDN
xMMI32_M_u4 net44 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u2 net11 CP VSS VSS Switch_NMOS_n12_X1_Y1
xMMI60_M_u2 Q net13 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u3 net7 SDN net44 VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u4 net37 net13 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u3 net33 SDN net37 VSS Switch_NMOS_n12_X1_Y1
xMMI20 net7 net83 net63 VSS Switch_NMOS_n12_X1_Y1
xMMI23 net25 net83 net5 VSS Switch_NMOS_n12_X1_Y1
xMMI22 net33 net11 net63 VSS Switch_NMOS_n12_X1_Y1
xMMI21 net25 D net20 VSS Switch_NMOS_n12_X1_Y1
xMMI25_M_u2 net13 net63 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI19 net20 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI24 net5 net7 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI40_M_u2 net83 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u3 net11 CP VDD VDD Switch_PMOS_n12_X1_Y1
xMMI33 net33 net83 net63 VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u1 net7 SDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI60_M_u3 Q net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI34 net25 net11 net96 VDD Switch_PMOS_n12_X1_Y1
xMMI30 net7 net11 net63 VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u2 net7 net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI28 net81 net83 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI40_M_u3 net83 net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u2 net33 net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI35 net96 net7 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u1 net33 SDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI25_M_u3 net13 net63 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI26 net25 D net81 VDD Switch_PMOS_n12_X1_Y1
.ends DFSNQD1

.subckt ND2D0 A1 A2 ZN
xMMI0_M_u3 ZN A1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u4 net1 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends ND2D0

.subckt DEL015 I Z
xMMI2_M_u2 Z net13 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI29 net25 net9 net28 VSS Switch_NMOS_n12_X1_Y1
xMMI30 net28 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI37 net17 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI28 net13 net9 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI35 net9 net5 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u2 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMI36 net44 net5 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u3 Z net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI20 net57 net9 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI23 net13 net9 net25 VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21 net25 net9 net57 VDD Switch_PMOS_n12_X1_Y1
xMMI32 net9 net5 net44 VDD Switch_PMOS_n12_X1_Y1
xMMI31 net44 net5 net33 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net33 net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DEL015

.subckt DFSND1 CP D Q QN SDN
xMMI32_M_u4 net57 net61 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u2 net11 CP VSS VSS Switch_NMOS_n12_X1_Y1
xMMI60_M_u2 Q net79 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u3 net97 SDN net57 VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u4 net40 net79 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u3 net25 SDN net40 VSS Switch_NMOS_n12_X1_Y1
xMMI20 net97 net81 net67 VSS Switch_NMOS_n12_X1_Y1
xMMI23 net61 net81 net5 VSS Switch_NMOS_n12_X1_Y1
xMMI22 net25 net11 net67 VSS Switch_NMOS_n12_X1_Y1
xMMI21 net61 D net9 VSS Switch_NMOS_n12_X1_Y1
xMMI25_M_u2 net79 net67 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI57_M_u2 QN net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI19 net9 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI24 net5 net97 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI40_M_u2 net81 net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u3 net11 CP VDD VDD Switch_PMOS_n12_X1_Y1
xMMI33 net25 net81 net67 VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u1 net97 SDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI60_M_u3 Q net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI34 net61 net11 net104 VDD Switch_PMOS_n12_X1_Y1
xMMI30 net97 net11 net67 VDD Switch_PMOS_n12_X1_Y1
xMMI57_M_u3 QN net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u2 net97 net61 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI28 net85 net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI40_M_u3 net81 net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u2 net25 net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI35 net104 net97 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u1 net25 SDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI25_M_u3 net79 net67 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI26 net61 D net85 VDD Switch_PMOS_n12_X1_Y1
.ends DFSND1

.subckt AN2D0 A1 A2 Z
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u4 net17 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net17 VSS Switch_NMOS_n12_X1_Y1
.ends AN2D0

.subckt DFCND1 CDN CP D Q QN
xMMI29_M_u2 QN net33 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI4 net53 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI18 net33 net5 net79 VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u3 net95 net79 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net81 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI15 net81 net67 net79 VSS Switch_NMOS_n12_X1_Y1
xMMI14_M_u2 net33 net95 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u2 net67 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net25 D net53 VSS Switch_NMOS_n12_X1_Y1
xMMI49 net20 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net17 net81 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 Q net95 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u4 net9 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI22_M_u2 net5 CP VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net25 net67 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI14_M_u3 net33 net95 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI22_M_u3 net5 CP VDD VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u3 net67 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI43 net72 net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net25 D net104 VDD Switch_PMOS_n12_X1_Y1
xMMI29_M_u3 QN net33 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 Q net95 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI44 net72 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI17 net33 net67 net79 VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net81 net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u1 net95 net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16 net81 net5 net79 VDD Switch_PMOS_n12_X1_Y1
xMMI45 net25 net5 net72 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net104 net67 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u2 net95 CDN VDD VDD Switch_PMOS_n12_X1_Y1
.ends DFCND1

.subckt AN2D2 A1 A2 Z
xMM_u3_1_M_u3 Z net9 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u2 net9 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_0_M_u3 Z net9 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net9 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u4 net29 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net9 A1 net29 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_1_M_u2 Z net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_0_M_u2 Z net9 VSS VSS Switch_NMOS_n12_X1_Y1
.ends AN2D2

.subckt CKBD4 I Z
xMM_u15_1 net11 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU23_1 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU23_3 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU23_0 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU23_2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u15_0 net11 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU21_0 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU21_1 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_0 net11 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU21_3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_1 net11 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU21_2 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKBD4

.subckt ND3D3 A1 A2 A3 ZN
xMMI0_0_M_u3 ZN A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_0_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_2_M_u3 ZN A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_2_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u3 ZN A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_0_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_2_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u5 net69 A2 net72 VSS Switch_NMOS_n12_X1_Y1
xMMI0_2_M_u6 net56 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_1_M_u4 ZN A1 net69 VSS Switch_NMOS_n12_X1_Y1
xMMI0_2_M_u4 ZN A1 net53 VSS Switch_NMOS_n12_X1_Y1
xMMI0_2_M_u5 net53 A2 net56 VSS Switch_NMOS_n12_X1_Y1
xMMI0_1_M_u6 net72 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_0_M_u6 net44 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_0_M_u5 net40 A2 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI0_0_M_u4 ZN A1 net40 VSS Switch_NMOS_n12_X1_Y1
.ends ND3D3

.subckt AN3D1 A1 A2 A3 Z
xMM_u4_M_u6 net13 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u5 net5 A2 net13 VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u4 net11 A1 net5 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 net11 A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u1 net11 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u2 net11 A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AN3D1

.subckt DEL_7b CKOUT EN LSB<3> LSB<2> LSB<1> REF_CLK SEL0 SEL1 SEL2 SEL3 SEL_DL
XI29 net87 net82 LSB<3> LSB<2> LSB<1> VDD VSS DEL_3x1_BIN
XI14 SEL3 SEL2 VDD VSS S2T<1> OR2D0
XI23 SEL1 S2T<1> VDD VSS net90 OR2D0
XI27 SEL1 S2T<3> VDD VSS net88 OR2D0
XI25 SEL1 S2T<2> VDD VSS net89 OR2D0
XI24 SEL0 S2T<1> VDD VSS net83 OR2D0
XI28 SEL0 S2T<3> VDD VSS net85 OR2D0
XI26 SEL0 S2T<2> VDD VSS net84 OR2D0
XI0 REF_CLK net82 SEL_DL VDD VSS net91 MUX2D0
XI19 net91 net76 S2T<0> net83 net90 VDD VSS DEL_3x1
XI22 net80 net86 S2T<3> SEL0 SEL1 VDD VSS DEL_4x1
XI21 net78 net80 S2T<2> net85 net88 VDD VSS DEL_4x1
XI20 net76 net78 S2T<1> net84 net89 VDD VSS DEL_4x1
XI18 SEL3 SEL2 VDD VSS S2T<3> AN2D0
XI16 EN VDD VSS S2T<0> BUFFD0
XI17 SEL3 VDD VSS S2T<2> BUFFD0
XI2 net82 VDD VSS CKOUT CKBD2
XI3 net76 net78 net80 net86 SEL2 SEL3 VDD VSS net87 MUX4ND0
.ends DEL_7b

.subckt DEL_3x1_BIN DEL_IN DEL_OUT LSB<3> LSB<2> LSB<1>
XI9 net020 net027 net033 VDD VSS DEL_OUT MUX2D1
XI1 net010 VDD VSS net032 DEL0
XI19 LSB<3> VDD VSS net013 DEL0
XI20 LSB<2> VDD VSS net035 DEL015
XI5 net030 VDD VSS net029 DEL015
XI21 LSB<1> VDD VSS net033 DEL015
XI3 DEL_IN net032 net013 VDD VSS net019 MUX2D0
XI6 net019 net029 net035 VDD VSS net020 MUX2D0
XI8 net028 VDD VSS net027 DEL005
XI14 DEL_IN VDD VSS net05 INVD0
XI16 net019 VDD VSS net018 INVD0
XI17 net020 VDD VSS net023 INVD0
XI15 net018 LSB<2> VDD VSS net030 ND2D0
XI13 net05 LSB<3> VDD VSS net010 ND2D0
XI18 net023 LSB<1> VDD VSS net028 ND2D0
.ends DEL_3x1_BIN

.subckt MUX2D1 I0 I1 S Z
xMMI14_M_u3 net5 I1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16_M_u3 net37 I0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU29_M_u3 Z net27 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI15_M_u3 net9 S VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u2 net5 net9 net27 VDD Switch_PMOS_n12_X1_Y1
xMMU18_M_u2 net37 S net27 VDD Switch_PMOS_n12_X1_Y1
xMMU18_M_u3 net37 net9 net27 VSS Switch_NMOS_n12_X1_Y1
xMMI15_M_u2 net9 S VSS VSS Switch_NMOS_n12_X1_Y1
xMMI16_M_u2 net37 I0 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u3 net5 S net27 VSS Switch_NMOS_n12_X1_Y1
xMMI14_M_u2 net5 I1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU29_M_u2 Z net27 VSS VSS Switch_NMOS_n12_X1_Y1
.ends MUX2D1

.subckt DEL0 I Z
xMMU7_M_u2 net11 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u2 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU5_M_u2 net25 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU5_M_u3 net25 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU7_M_u3 net11 net25 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DEL0

.subckt MUX2D0 I0 I1 S Z
xMMU29_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI15_M_u3 net17 S VDD VDD Switch_PMOS_n12_X1_Y1
xMMI111 net13 I0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI24 net9 I1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 net5 S net13 VDD Switch_PMOS_n12_X1_Y1
xMMI25 net5 net17 net9 VDD Switch_PMOS_n12_X1_Y1
xMMI15_M_u2 net17 S VSS VSS Switch_NMOS_n12_X1_Y1
xMMI20 net36 I1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 net5 net17 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI21 net5 S net36 VSS Switch_NMOS_n12_X1_Y1
xMMU29_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI19 net25 I0 VSS VSS Switch_NMOS_n12_X1_Y1
.ends MUX2D0

.subckt DEL005 I Z
xMMI2_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMI10 net11 I net5 VDD Switch_PMOS_n12_X1_Y1
xMMI13 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 net11 I net5 VSS Switch_NMOS_n12_X1_Y1
.ends DEL005

.subckt OR2D0 A1 A2 Z
xMMU1_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u4 net5 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u3 net5 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u1 net17 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u2 net5 A1 net17 VDD Switch_PMOS_n12_X1_Y1
.ends OR2D0

.subckt DEL_3x1 DEL_IN DEL_OUT EN SEL0 SEL1
XI18 SEL1 SEL0 VDD VSS S2T<3> AN2D0
XI8 net12 S2T<3> VDD VSS net18 AN2D0
XI6 net11 S2T<2> VDD VSS net19 AN2D0
XI4 net21 S2T<1> VDD VSS net20 AN2D0
XI2 DEL_IN S2T<0> VDD VSS net21 AN2D0
XI9 net18 VDD VSS net17 DEL1
XI7 net19 VDD VSS net12 DEL1
XI5 net20 VDD VSS net11 DEL1
XI11 net21 net11 net12 net17 SEL0 SEL1 VDD VSS DEL_OUT MUX4D0
XI17 SEL1 VDD VSS S2T<2> BUFFD0
XI16 EN VDD VSS S2T<0> BUFFD0
XI14 SEL1 SEL0 VDD VSS S2T<1> OR2D0
.ends DEL_3x1

.subckt DEL1 I Z
xMMU7_M_u2 net11 net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u2 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU5_M_u2 net25 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU5_M_u3 net25 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU7_M_u3 net11 net25 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DEL1

.subckt MUX4D0 I0 I1 I2 I3 S0 S1 Z
xMMU18_M_u3 Z net20 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI53_M_u2 net97 S1 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI51_M_u3 net37 I3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI55_M_u2 net37 net61 net104 VDD Switch_PMOS_n12_X1_Y1
xMMI50_M_u3 net33 S1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI48_M_u3 net61 S0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI49_M_u3 net81 I2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI47_M_u3 net5 I1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI56_M_u2 net104 net33 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI54_M_u2 net81 S0 net104 VDD Switch_PMOS_n12_X1_Y1
xMMI40_M_u2 net9 S0 net97 VDD Switch_PMOS_n12_X1_Y1
xMMI52_M_u2 net5 net61 net97 VDD Switch_PMOS_n12_X1_Y1
xMMI46_M_u3 net9 I0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI55_M_u3 net37 S0 net104 VSS Switch_NMOS_n12_X1_Y1
xMMI53_M_u3 net97 net33 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI47_M_u2 net5 I1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI51_M_u2 net37 I3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI52_M_u3 net5 S0 net97 VSS Switch_NMOS_n12_X1_Y1
xMMI54_M_u3 net81 net61 net104 VSS Switch_NMOS_n12_X1_Y1
xMMI56_M_u3 net104 S1 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI40_M_u3 net9 net61 net97 VSS Switch_NMOS_n12_X1_Y1
xMMI49_M_u2 net81 I2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU18_M_u2 Z net20 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48_M_u2 net61 S0 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI46_M_u2 net9 I0 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI50_M_u2 net33 S1 VSS VSS Switch_NMOS_n12_X1_Y1
.ends MUX4D0

.subckt BUFFD0 I Z
xMMI2_M_u2 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends BUFFD0

.subckt DEL_4x1 DEL_IN DEL_OUT EN SEL0 SEL1
XI18 SEL1 SEL0 VDD VSS S2T<3> AN2D0
XI8 net12 S2T<3> VDD VSS net18 AN2D0
XI6 net11 S2T<2> VDD VSS net19 AN2D0
XI4 net10 S2T<1> VDD VSS net20 AN2D0
XI2 DEL_IN S2T<0> VDD VSS net21 AN2D0
XI9 net18 VDD VSS net17 DEL1
XI7 net19 VDD VSS net12 DEL1
XI5 net20 VDD VSS net11 DEL1
XI3 net21 VDD VSS net10 DEL1
XI11 net10 net11 net12 net17 SEL0 SEL1 VDD VSS DEL_OUT MUX4D0
XI17 SEL1 VDD VSS S2T<2> BUFFD0
XI16 EN VDD VSS S2T<0> BUFFD0
XI14 SEL1 SEL0 VDD VSS S2T<1> OR2D0
.ends DEL_4x1

.subckt CKBD2 I Z
xMMU23_1 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u15 net5 I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU23_0 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3 net5 I VDD VDD Switch_PMOS_n12_X1_Y1
xMMU21_0 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU21_1 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKBD2

.subckt MUX4ND0 I0 I1 I2 I3 S0 S1 ZN
xMMI47_M_u2 net17 I2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI51_M_u3 net20 S1 ZN VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u2 net61 I0 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI50_M_u3 net33 net83 ZN VSS Switch_NMOS_n12_X1_Y1
xMMI48_M_u3 net61 net67 net33 VSS Switch_NMOS_n12_X1_Y1
xMMI58_M_u2 net67 S0 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI49_M_u3 net5 S0 net33 VSS Switch_NMOS_n12_X1_Y1
xMMI52_M_u3 net17 net67 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI54_M_u3 net9 S0 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI57_M_u2 net9 I3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI56_M_u2 net5 I1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU18_M_u2 net83 S1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI55_M_u3 net61 I0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU18_M_u3 net83 S1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI58_M_u3 net67 S0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI51_M_u2 net20 net83 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI57_M_u3 net9 I3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI56_M_u3 net5 I1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI47_M_u3 net17 I2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI49_M_u2 net5 net67 net33 VDD Switch_PMOS_n12_X1_Y1
xMMI48_M_u2 net61 S0 net33 VDD Switch_PMOS_n12_X1_Y1
xMMI54_M_u2 net9 net67 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI52_M_u2 net17 S0 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI50_M_u2 net33 S1 ZN VDD Switch_PMOS_n12_X1_Y1
.ends MUX4ND0

.subckt MDLL_LOGIC_VLOG CODE<6> CODE<5> CODE<4> CODE<3> CODE<2> CODE<1> CODE<0> COMP EN0DLL FRCODE<6> FRCODE<5> FRCODE<4> FRCODE<3> FRCODE<2> FRCODE<1> FRCODE<0> FREE0RUN REFCLK SAR0EN STATUS<2> STATUS<1> STATUS<0> TRK0EN
XU85 N130 VDD VSS N131 CKND0
XU2 SAR0CODE<5> VDD VSS N2 CKND0
XU3 SAR0CODE<2> VDD VSS N3 CKND0
XU4 SAR0CODE<4> VDD VSS N4 CKND0
XU5 SAR0CODE<0> VDD VSS N5 CKND0
XU6 STATUS<0> VDD VSS N6 CKND0
XU1 FREE0RUN VDD VSS N1 CKND0
XU56 N41 N75 N27 N53 VDD VSS N89 AO22D0
XU100 N39 N75 N25 N53 VDD VSS N125 AO22D0
XU106 N1 SAR0CODE<3> FRCODE<3> FREE0RUN VDD VSS CODE<3> AO22D0
XU105 N1 SAR0CODE<2> FRCODE<2> FREE0RUN VDD VSS CODE<2> AO22D0
XU104 N1 SAR0CODE<1> FRCODE<1> FREE0RUN VDD VSS CODE<1> AO22D0
XU103 N1 SAR0CODE<0> FRCODE<0> FREE0RUN VDD VSS CODE<0> AO22D0
XU156 N136 FREE0RUN FRCODE<6> FREE0RUN VDD VSS CODE<6> MOAI22D1
XU155 FREE0RUN N2 FRCODE<5> FREE0RUN VDD VSS CODE<5> MOAI22D1
XU154 FREE0RUN N4 FRCODE<4> FREE0RUN VDD VSS CODE<4> MOAI22D1
XU75 N111 N6 VDD VSS N620 CKAN2D0
XU69 N110 N56 VDD VSS N71 CKAN2D0
XU90 N69 N110 VDD VSS N70 CKAN2D0
XU107 N64 N73 VDD VSS N76 AN2XD1
XU68 N113 N6 VDD VSS N56 AN2XD1
XU63 N640 N108 VDD VSS N55 AN2XD1
XU92 N113 STATUS<0> VDD VSS N69 AN2XD1
XU65 N55 N69 VDD VSS N68 AN2XD1
XU81 N82 N130 N81 VDD VSS N73 AN3D0
XU89 N111 N6 N110 VDD VSS N74 AN3D0
XU57 COMP N88 N118 VDD VSS N53 AN3XD1
XU91 N55 STATUS<0> N111 VDD VSS N67 AN3XD1
XU73 N29 N53 VDD VSS N610 ND2D1
XU72 SAR0CODE<4> N101 VDD VSS N600 ND2D1
XU96 N45 N75 VDD VSS N119 ND2D1
XU95 N31 N53 VDD VSS N120 ND2D1
XU101 N6 N85 VDD VSS N107 ND2D1
XU67 STATUS<1> STATUS<0> VDD VSS N590 ND2D1
XU79 N630 N590 VDD VSS N640 ND2D1
XU66 N640 N108 VDD VSS N110 ND2D1
XU80 STATUS<2> VDD VSS N630 INVD1
XU58 N590 VDD VSS N109 INVD1
XU77 N111 VDD VSS N113 INVD1
XU55 N107 N590 VDD VSS N111 CKND2D2
XU133 N97 N96 VDD VSS N46 CKND2D1
XU153 N133 N132 VDD VSS N48 CKND2D1
XU121 N129 N91 VDD VSS N84 CKND2D1
XU60 STATUS<2> N109 VDD VSS N108 CKND2D1
XU150 SAR0CODE<1> VDD VSS N127 CKND1
XU141 N115 VDD VSS N103 CKND1
XU123 N94 VDD VSS N83 CKND1
XU138 N104 VDD VSS N114 CKND1
XU125 SAR0EN VDD VSS N87 CKND1
XU139 N101 VDD VSS N102 CKND1
XU126 STATUS<1> VDD VSS N85 CKND1
XU129 SAR0CODE<3> VDD VSS N92 CKND1
XU134 N98 VDD VSS N99 CKND1
XU120 N137 VDD VSS N91 CKND1
XU119 N124 VDD VSS N129 CKND1
XU117 COMP VDD VSS N86 CKND1
XU115 N80 VDD VSS N88 CKND1
XU87 N114 N2 VDD VSS N117 CKND2D0
XU71 STATUS<2> N109 VDD VSS N58 CKND2D0
XU157 SAR0CODE<1> N5 VDD VSS N137 IND2D0
XU82 N107 N630 VDD VSS N118 IND2D0
XSUB049 SAR0CODE<6> N2 SAR0CODE<4> SAR0CODE<3> N3 SAR0CODE<1> N5 N74 N70 N71 N67 N72 N68 N66 N45 N44 N43 N42 N41 N40 N39 SAR0CODE<0> SAR0CODE<2> SAR0CODE<5> VDD VSS MDLL_LOGIC_VLOG_DW01_sub_J17_0
XADD049 SAR0CODE<6> SAR0CODE<5> N4 SAR0CODE<3> N3 SAR0CODE<1> SAR0CODE<0> N74 N70 N71 N67 N72 N68 N66 SAR0CODE<4> SAR0CODE<2> N31 N30 N29 N28 N27 N26 N25 VDD VSS MDLL_LOGIC_VLOG_DW01_add_J16_0
XU114 N58 VDD VSS N82 INVD0
XU99 N123 N122 VDD VSS N430 IND2D1
XU118 COMP0REG N86 VDD VSS N81 IND2D1
XU116 TRK0EN N82 VDD VSS N130 IND2D1
XU93 N81 N82 N130 VDD VSS N124 IND3D1
XADD051 SAR0CODE<6> SAR0CODE<5> SAR0CODE<4> SAR0CODE<3> SAR0CODE<2> SAR0CODE<1> SAR0CODE<0> N64 N63 N62 N61 N60 N59 VDD VSS MDLL_LOGIC_VLOG_DW01_inc_0
XU131 N3 N92 N98 VDD VSS N95 OAI21D1
XU151 N5 N127 N137 VDD VSS N128 OAI21D1
XU140 N4 N124 N102 VDD VSS N115 OAI21D1
XU135 N99 N124 N130 VDD VSS N101 OAI21D1
XU122 N91 N124 N130 VDD VSS N94 OAI21D1
XU74 N600 N610 N104 VDD VSS N100 ND3D1
XU94 N120 N119 N118 VDD VSS N121 ND3D1
XU130 N91 N92 N3 VDD VSS N98 ND3D1
XU137 N99 N129 N4 VDD VSS N104 ND3D1
XU70 N113 N6 VDD VSS N65 CKAN2D1
XU64 N55 N65 VDD VSS N66 AN2D2
XU76 N55 N620 VDD VSS N72 AN2D1
XSAR0CODE0REG030 EN0DLL REFCLK N46 SAR0CODE<3> VDD VSS DFCNQD1
XSAR0CODE0REG040 EN0DLL REFCLK N450 SAR0CODE<4> VDD VSS DFCNQD1
XSAR0CODE0REG010 EN0DLL REFCLK N48 SAR0CODE<1> VDD VSS DFCNQD1
XSAR0CODE0REG050 EN0DLL REFCLK N440 SAR0CODE<5> VDD VSS DFCNQD1
XSAR0CODE0REG020 EN0DLL REFCLK N47 SAR0CODE<2> VDD VSS DFCNQD1
XCOMP0REG0REG EN0DLL REFCLK N54 COMP0REG VDD VSS DFCNQD1
XSTATUS0REG010 EN0DLL REFCLK N51 STATUS<1> VDD VSS DFCNQD1
XSTATUS0REG000 EN0DLL REFCLK N52 STATUS<0> VDD VSS DFCNQD1
XSTATUS0REG020 EN0DLL REFCLK N50 STATUS<2> VDD VSS DFCNQD1
XU109 N590 N80 N630 VDD VSS N50 OAI21D0
XU78 STATUS<1> N79 VDD VSS N51 CKXOR2D0
XU112 STATUS<0> N88 VDD VSS N52 CKXOR2D0
XU110 N6 N80 VDD VSS N79 NR2D0
XU113 SAR0EN N58 VDD VSS N80 ND2D0
XU83 N87 N86 N118 N58 VDD VSS N75 OA211D0
XU59 COMP VDD VSS N54 DEL005
XU144 N63 N73 N106 N105 VDD VSS N440 AO211D1
XU127 N60 N73 N90 N89 VDD VSS N47 AO211D1
XU148 N5 N73 N126 N125 VDD VSS N49 AO211D1
XU142 N104 N103 SAR0CODE<5> VDD VSS N106 MUX2ND0
XU124 N84 N83 SAR0CODE<2> VDD VSS N90 MUX2ND0
XU146 N117 N116 SAR0CODE<6> VDD VSS N123 MUX2ND0
XU147 N124 N130 SAR0CODE<0> VDD VSS N126 MUX2ND0
XSAR0CODE0REG000 EN0DLL REFCLK N49 SAR0CODE<0> VDD VSS DFCNQD4
XU88 N121 N76 VDD VSS N122 NR2XD0
XSAR0CODE0REG060 REFCLK N430 SAR0CODE<6> N136 EN0DLL VDD VSS DFSND1
XU84 N129 SAR0CODE<5> N115 VDD VSS N116 AOI21D0
XU143 N44 N75 N30 N53 VDD VSS N105 AO22D1
XU132 N42 N75 N61 N73 VDD VSS N96 AOI22D1
XU152 N59 N73 N131 SAR0CODE<1> VDD VSS N132 AOI22D1
XU98 N28 N53 N129 N95 SAR0CODE<3> N94 VDD VSS N97 AOI222D0
XU97 N40 N75 N129 N128 N26 N53 VDD VSS N133 AOI222D0
XU86 N43 N75 N62 N73 N100 VDD VSS N450 AO221D1
.ends MDLL_LOGIC_VLOG

.subckt CKND0 I ZN
xMM_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u1 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKND0

.subckt AO22D0 A1 A2 B1 B2 Z
xMMI23 net17 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI8_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI16 net5 B1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI24 net5 A1 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI22 net1 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI20 net5 A1 net33 VDD Switch_PMOS_n12_X1_Y1
xMM_u2 net33 B2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI19 net5 A2 net33 VDD Switch_PMOS_n12_X1_Y1
xMMI8_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21 net33 B1 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AO22D0

.subckt MOAI22D1 A1 A2 B1 B2 ZN
xMMU1 net37 B1 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI6 net9 net37 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU9 net9 A1 ZN VSS Switch_NMOS_n12_X1_Y1
xMMI5 net20 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU10 net9 A2 ZN VSS Switch_NMOS_n12_X1_Y1
xMMI1 net37 B1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI3 net33 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI4 ZN A1 net33 VDD Switch_PMOS_n12_X1_Y1
xMMI2 ZN net37 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU3 net37 B2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends MOAI22D1

.subckt CKAN2D0 A1 A2 Z
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u4 net21 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net21 VSS Switch_NMOS_n12_X1_Y1
.ends CKAN2D0

.subckt AN2XD1 A1 A2 Z
xMM_u2_M_u4 net9 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net9 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AN2XD1

.subckt AN3D0 A1 A2 A3 Z
xMM_u4_M_u6 net13 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u5 net5 A2 net13 VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u4 net11 A1 net5 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 net11 A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u1 net11 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u2 net11 A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AN3D0

.subckt AN3XD1 A1 A2 A3 Z
xMM_u4_M_u6 net13 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u5 net5 A2 net13 VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u4 net11 A1 net5 VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u3 Z net11 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 net11 A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u1 net11 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u2 net11 A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AN3XD1

.subckt ND2D1 A1 A2 ZN
xMMI1_M_u3 ZN A1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 net1 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends ND2D1

.subckt CKND2D2 A1 A2 ZN
xMMI0_0_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_0_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_1_M_u4 net24 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_0_M_u3 ZN A1 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI0_1_M_u3 ZN A1 net24 VSS Switch_NMOS_n12_X1_Y1
xMMI0_0_M_u4 net17 A2 VSS VSS Switch_NMOS_n12_X1_Y1
.ends CKND2D2

.subckt CKND2D1 A1 A2 ZN
xMMI0_M_u3 ZN A1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u4 net1 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKND2D1

.subckt CKND1 I ZN
xMM_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u1 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKND1

.subckt CKND2D0 A1 A2 ZN
xMMU1_M_u3 ZN A1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u4 net1 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
.ends CKND2D0

.subckt IND2D0 A1 B1 ZN
xMMI2_M_u3 net9 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI11 VDD B1 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u16 VDD net9 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI13 net21 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 net9 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 ZN B1 net21 VSS Switch_NMOS_n12_X1_Y1
.ends IND2D0

.subckt MDLL_LOGIC_VLOG_DW01_sub_J17_0 A<6> A<5> A<4> A<3> A<2> A<1> A<0> B<6> B<5> B<4> B<3> B<2> B<1> B<0> DIFF<6> DIFF<5> DIFF<4> DIFF<3> DIFF<2> DIFF<1> DIFF<0> IN0 IN1 IN2
XU35 N1 N16 VDD VSS N15 ND2D1
XU45 N10 N12 VDD VSS N22 ND2D1
XU34 N1 N18 VDD VSS N24 ND2D1
XU38 A<3> N41 VDD VSS N36 ND2D1
XU15 IN1 N44 VDD VSS N35 ND2D1
XU6 B<3> N42 VDD VSS N37 ND2D1
XU37 A<1> N54 VDD VSS N27 ND2D1
XU7 B<1> N55 VDD VSS N29 ND2D1
XU10 N23 N18 VDD VSS N10 ND2D1
XU32 N48 N29 VDD VSS N26 ND2D1
XU9 B<0> IN0 VDD VSS N51 IND2D2
XU55 N18 VDD VSS N17 CKND1
XU62 N35 VDD VSS N43 CKND1
XU13 N25 VDD VSS N14 CKND1
XU60 N37 VDD VSS N34 CKND1
XU54 N9 VDD VSS N11 CKND1
XU64 N51 VDD VSS N48 CKND1
XU26 B<0> A<0> N48 VDD VSS DIFF<0> AO21D0
XU8 N37 N36 VDD VSS N40 CKND2D0
XU25 N51 N52 VDD VSS N50 CKND2D0
XU24 N29 N27 VDD VSS N49 CKND2D0
XU20 B<2> A<2> VDD VSS N38 CKND2D0
XU30 N38 N35 VDD VSS N2 AN2XD1
XU28 N38 N37 VDD VSS N1 AN2XD1
XU46 IN2 B<5> VDD VSS N9 IND2D1
XU42 B<4> A<4> VDD VSS N12 IND2D1
XU40 A<4> B<4> VDD VSS N18 IND2D1
XU49 B<2> VDD VSS N44 INVD1
XU43 A<3> VDD VSS N42 INVD1
XU39 A<1> VDD VSS N55 INVD1
XU48 B<0> VDD VSS N53 CKND0
XU21 B<3> VDD VSS N41 CKND0
XU19 B<1> VDD VSS N54 CKND0
XU52 N4 N5 VDD VSS DIFF<6> CKXOR2D1
XU53 B<6> A<6> VDD VSS N5 CKXOR2D1
XU56 N19 N20 VDD VSS DIFF<5> CKXOR2D1
XU57 B<5> IN2 VDD VSS N20 CKXOR2D1
XU59 B<4> A<4> VDD VSS N32 CKXOR2D1
XU58 N31 N32 VDD VSS DIFF<4> CKXOR2D1
XU61 N39 N40 VDD VSS DIFF<3> CKXOR2D1
XU29 N33 N2 VDD VSS DIFF<2> CKXOR2D1
XU27 N34 N35 N36 VDD VSS N23 OAI21D1
XU51 IN0 B<0> VDD VSS N30 IND2D0
XU50 IN0 B<0> VDD VSS N47 IND2D0
XU12 N29 N30 VDD VSS N28 ND2D0
XU11 N29 N47 VDD VSS N46 ND2D0
XU47 N26 N27 N28 VDD VSS N25 ND3D1
XU5 N26 N27 N46 VDD VSS N33 ND3D1
XU63 N49 N50 VDD VSS DIFF<1> XNR2D1
XU17 N14 N15 VDD VSS N6 NR2D0
XU23 IN0 N53 VDD VSS N52 NR2D0
XU16 N1 N33 N23 VDD VSS N31 AOI21D0
XU18 N33 N38 N43 VDD VSS N39 AOI21D0
XU22 N21 N22 VDD VSS N19 NR2XD0
XU36 N17 N11 VDD VSS N16 NR2D1
XU33 N14 N24 VDD VSS N21 NR2D1
XU3 N6 N7 N8 VDD VSS N4 NR3D0
XU31 N9 N10 VDD VSS N8 INR2D1
XU14 N11 N12 B<5> A<5> VDD VSS N7 OAI22D0
.ends MDLL_LOGIC_VLOG_DW01_sub_J17_0

.subckt IND2D2 A1 B1 ZN
xMMI3 VDD net11 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u16 VDD B1 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI9_M_u3 net11 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI9_M_u2 net11 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI4 net20 B1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI11 net21 B1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 ZN net11 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI10 ZN net11 net21 VSS Switch_NMOS_n12_X1_Y1
.ends IND2D2

.subckt AO21D0 A1 A2 B Z
xMMI9 net5 A2 net9 VDD Switch_PMOS_n12_X1_Y1
xMM_u2 net9 B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI10 net5 A1 net9 VDD Switch_PMOS_n12_X1_Y1
xMMI8_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI11 net5 A1 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI12 net25 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI8_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI6 net5 B VSS VSS Switch_NMOS_n12_X1_Y1
.ends AO21D0

.subckt IND2D1 A1 B1 ZN
xMMI2_M_u3 net9 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI11 VDD B1 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u16 VDD net9 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI13 net21 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 net9 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 ZN B1 net21 VSS Switch_NMOS_n12_X1_Y1
.ends IND2D1

.subckt CKXOR2D1 A1 A2 Z
xMM_u6_M_u2 net27 A1 net44 VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 Z net44 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u5_M_u3 net5 net27 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u8_M_u3 net9 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_M_u2 net5 net9 net44 VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u3 net27 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u6_M_u3 net27 net9 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u3 net5 A1 net44 VSS Switch_NMOS_n12_X1_Y1
xMM_u8_M_u2 net9 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u2 Z net44 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u2 net27 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u5_M_u2 net5 net27 VSS VSS Switch_NMOS_n12_X1_Y1
.ends CKXOR2D1

.subckt OAI21D1 A1 A2 B ZN
xMMI16_MI13 net9 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u9 ZN B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16_MI12 ZN A1 net9 VDD Switch_PMOS_n12_X1_Y1
xMM_u3 ZN A2 net24 VSS Switch_NMOS_n12_X1_Y1
xMM_u4 net24 B VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2 ZN A1 net24 VSS Switch_NMOS_n12_X1_Y1
.ends OAI21D1

.subckt ND3D1 A1 A2 A3 ZN
xMMI1_M_u5 net9 A2 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 ZN A1 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u6 net1 A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 ZN A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends ND3D1

.subckt XNR2D1 A1 A2 ZN
xMM_u6_M_u2 net27 net9 net44 VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 ZN net44 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u5_M_u3 net5 net27 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u8_M_u3 net9 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0_M_u2 net5 A1 net44 VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u3 net27 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u6_M_u3 net27 A1 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI0_M_u3 net5 net9 net44 VSS Switch_NMOS_n12_X1_Y1
xMM_u8_M_u2 net9 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u2 ZN net44 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u2 net27 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u5_M_u2 net5 net27 VSS VSS Switch_NMOS_n12_X1_Y1
.ends XNR2D1

.subckt AOI21D0 A1 A2 B ZN
xMMI9 ZN A1 net5 VDD Switch_PMOS_n12_X1_Y1
xMM_u2 net5 B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI8 ZN A2 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI2 ZN A1 net13 VSS Switch_NMOS_n12_X1_Y1
xMMI11 ZN B VSS VSS Switch_NMOS_n12_X1_Y1
xMMI10 net13 A2 VSS VSS Switch_NMOS_n12_X1_Y1
.ends AOI21D0

.subckt NR2XD0 A1 A2 ZN
xMMI1_M_u3 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 net13 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A1 net13 VDD Switch_PMOS_n12_X1_Y1
.ends NR2XD0

.subckt NR2D1 A1 A2 ZN
xMMI1_M_u3 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 net13 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A1 net13 VDD Switch_PMOS_n12_X1_Y1
.ends NR2D1

.subckt NR3D0 A1 A2 A3 ZN
xMMI3 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4 ZN A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1 ZN A1 net13 VDD Switch_PMOS_n12_X1_Y1
xMM_u1 net17 A3 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI0 net13 A2 net17 VDD Switch_PMOS_n12_X1_Y1
.ends NR3D0

.subckt INR2D1 A1 B1 ZN
xMMU1_M_u3 ZN net11 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u4 ZN B1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU6_M_u2 net11 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU6_M_u3 net11 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU1_M_u2 ZN B1 net20 VDD Switch_PMOS_n12_X1_Y1
xMMU1_M_u1 net20 net11 VDD VDD Switch_PMOS_n12_X1_Y1
.ends INR2D1

.subckt OAI22D0 A1 A2 B1 B2 ZN
xMM_u4 net13 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI8 ZN A2 net13 VSS Switch_NMOS_n12_X1_Y1
xMMI9 ZN A1 net13 VSS Switch_NMOS_n12_X1_Y1
xMMI7 net13 B1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI4 ZN B1 net32 VDD Switch_PMOS_n12_X1_Y1
xMMI6 ZN A1 net17 VDD Switch_PMOS_n12_X1_Y1
xMMU24 net32 B2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 net17 A2 VDD VDD Switch_PMOS_n12_X1_Y1
.ends OAI22D0

.subckt MDLL_LOGIC_VLOG_DW01_add_J16_0 A<6> A<5> A<4> A<3> A<2> A<1> A<0> B<6> B<5> B<4> B<3> B<2> B<1> B<0> IN0 IN1 SUM<6> SUM<5> SUM<4> SUM<3> SUM<2> SUM<1> SUM<0>
XU41 A<0> B<0> VDD VSS N19 CKND2D0
XU17 N30 N28 VDD VSS N32 CKND2D0
XU18 B<2> IN1 VDD VSS N34 CKND2D0
XU39 N21 N20 VDD VSS N37 CKND2D0
XU19 B<3> A<3> VDD VSS N28 CKND2D0
XU35 B<0> A<0> VDD VSS N38 CKND2D0
XU14 N11 N12 VDD VSS N10 ND2D1
XU11 N36 N20 VDD VSS N26 ND2D1
XU30 B<1> A<1> VDD VSS N20 ND2D1
XU32 B<3> A<3> VDD VSS N30 OR2D1
XU10 B<1> A<1> VDD VSS N21 OR2D1
XU3 B<2> A<2> VDD VSS N29 IND2D1
XU31 B<4> A<4> VDD VSS N15 IND2D1
XU47 N34 VDD VSS N33 CKND1
XU16 N30 VDD VSS N16 CKND1
XU45 N29 VDD VSS N17 CKND1
XU36 N24 N7 VDD VSS SUM<4> XNR2D1
XU43 B<6> A<6> VDD VSS N9 XNR2D1
XU20 N10 N5 VDD VSS SUM<5> XNR2D1
XU21 B<5> A<5> VDD VSS N5 XNR2D1
XU34 A<0> B<0> VDD VSS N39 NR2D0
XU33 N38 N39 VDD VSS SUM<0> INR2D1
XU27 B<4> IN0 VDD VSS N7 CKXOR2D1
XU42 N8 N9 VDD VSS SUM<6> CKXOR2D1
XU46 N31 N32 VDD VSS SUM<3> CKXOR2D1
XU24 N26 N6 VDD VSS SUM<2> CKXOR2D1
XU23 N37 N38 VDD VSS SUM<1> CKXOR2D1
XU6 B<4> IN0 VDD VSS N2 AN2XD1
XU5 B<5> A<5> VDD VSS N1 AN2XD1
XU8 B<0> A<0> VDD VSS N4 AN2XD1
XU25 N29 N34 VDD VSS N6 AN2XD1
XU13 N21 N4 VDD VSS N36 ND2D0
XU38 IN1 B<2> VDD VSS N27 CKND2D1
XU44 N18 N19 N20 VDD VSS N13 OAI21D1
XU26 N16 N27 N28 VDD VSS N22 OAI21D1
XU15 N26 N29 N33 VDD VSS N31 AOI21D0
XU28 N25 N26 N22 VDD VSS N24 AOI21D1
XU9 N22 N15 N2 VDD VSS N11 AOI21D1
XU29 N3 N10 N1 VDD VSS N8 AOI21D1
XU7 A<5> B<5> VDD VSS N3 OR2XD1
XU37 N21 VDD VSS N18 INVD1
XU12 N16 N17 VDD VSS N14 NR2XD0
XU22 N14 N15 N13 VDD VSS N12 ND3D1
XU40 N16 N17 VDD VSS N25 NR2D1
.ends MDLL_LOGIC_VLOG_DW01_add_J16_0

.subckt OR2D1 A1 A2 Z
xMMU1_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u4 net5 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u3 net5 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u1 net17 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u2 net5 A1 net17 VDD Switch_PMOS_n12_X1_Y1
.ends OR2D1

.subckt AOI21D1 A1 A2 B ZN
xMM_u3 net5 A1 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u2 net5 B VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4 net5 A2 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI2 ZN A1 net13 VSS Switch_NMOS_n12_X1_Y1
xMM_u7 ZN B VSS VSS Switch_NMOS_n12_X1_Y1
xMMI3 net13 A2 VSS VSS Switch_NMOS_n12_X1_Y1
.ends AOI21D1

.subckt OR2XD1 A1 A2 Z
xMMU1_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u4 net5 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u7_M_u3 net5 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u1 net17 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u7_M_u2 net5 A1 net17 VDD Switch_PMOS_n12_X1_Y1
.ends OR2XD1

.subckt IND3D1 A1 B1 B2 ZN
xMMI4 VDD net19 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI11 VDD B2 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u16 VDD B1 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI5_M_u3 net19 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5_M_u2 net19 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI6 net25 B1 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI12 ZN B2 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI7 net17 net19 VSS VSS Switch_NMOS_n12_X1_Y1
.ends IND3D1

.subckt MDLL_LOGIC_VLOG_DW01_inc_0 A<6> A<5> A<4> A<3> A<2> A<1> A<0> SUM<6> SUM<5> SUM<4> SUM<3> SUM<2> SUM<1>
XU10103 A<3> CARRY<3> CARRY<4> SUM<3> VDD VSS HA1D0
XU10101 A<1> A<0> CARRY<2> SUM<1> VDD VSS HA1D0
XU10102 A<2> CARRY<2> CARRY<3> SUM<2> VDD VSS HA1D0
XU10104 A<4> CARRY<4> CARRY<5> SUM<4> VDD VSS HA1D0
XU10105 A<5> CARRY<5> CARRY<6> SUM<5> VDD VSS HA1D0
XU2 CARRY<6> A<6> VDD VSS SUM<6> CKXOR2D0
.ends MDLL_LOGIC_VLOG_DW01_inc_0

.subckt INV_LVT zn i SN SP
xxm0 zn i SN SN Switch_NMOS_n12_X1_Y1
xxm1 zn i SP SP Switch_PMOS_n12_X1_Y1
.ends INV_LVT

.subckt stage2_inv G1 SN G2 SP
MM0_MM2 D SN SP G1 INV_LVT
MM1_MM3 G2 SN SP D INV_LVT
.ends stage2_inv

.subckt tgate D GA S GB
xM0 D GA S BN Switch_NMOS_n12_X1_Y1
xM1 D GB S BP Switch_PMOS_n12_X1_Y1
.ends tgate

.subckt HA1D0 A B CO S
xMMU9_M_u1 net25 A VDD VDD Switch_PMOS_n12_X1_Y1
xMMU9_M_u2 net25 B VDD VDD Switch_PMOS_n12_X1_Y1
xMMU9_M_u4 net56 B VSS VSS Switch_NMOS_n12_X1_Y1
xMMU9_M_u3 net25 A net56 VSS Switch_NMOS_n12_X1_Y1
MMU2_M_u2_MMU1_M_u2_MMU2_M_u3_MMU1_M_u3 VSS A VDD net13 stage2_inv
MMU3_M_u2_MMU3_M_u3 B VSS VDD net5 INV_LVT
MMU5_M_u2_MMU5_M_u3 net25 VSS VDD CO INV_LVT
MMU4_M_u2_MMU4_M_u3 net72 VSS VDD S INV_LVT
MMU7_M_u3_MMU7_M_u2 B net72 net5 net13 tgate
MMU8_M_u3_MMU8_M_u2 net5 net72 B net9 tgate
.ends HA1D0

.subckt CKXOR2D0 A1 A2 Z
xMM_u6_M_u3 net37 net17 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u2 net17 A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4_M_u2 Z net44 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI3_M_u3 net5 A1 net44 VSS Switch_NMOS_n12_X1_Y1
xMM_u5_M_u2 net5 net37 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u2 net37 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2_M_u3 net17 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u6_M_u2 net37 A1 net44 VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u3 net37 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u4_M_u3 Z net44 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u5_M_u3 net5 net37 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI3_M_u2 net5 net17 net44 VDD Switch_PMOS_n12_X1_Y1
.ends CKXOR2D0

.subckt CKAN2D1 A1 A2 Z
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u4 net21 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net21 VSS Switch_NMOS_n12_X1_Y1
.ends CKAN2D1

.subckt AN2D1 A1 A2 Z
xMM_u3_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u1 net5 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u2_M_u2 net5 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u3_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u4 net17 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2_M_u3 net5 A1 net17 VSS Switch_NMOS_n12_X1_Y1
.ends AN2D1

.subckt DFCNQD1 CDN CP D Q
xMMI4 net53 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u3 net81 net51 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net37 net97 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI29 net51 net5 net44 VSS Switch_NMOS_n12_X1_Y1
xMMI15 net37 net63 net51 VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u2 net63 net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net97 D net53 VSS Switch_NMOS_n12_X1_Y1
xMMI49 net20 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI26 net44 net81 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net17 net37 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 Q net81 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u4 net9 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI22_M_u2 net5 CP VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net97 net63 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI22_M_u3 net5 CP VDD VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u3 net63 net5 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI43 net101 net37 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net97 D net100 VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 Q net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI44 net101 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net37 net97 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u1 net81 net51 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16 net37 net5 net51 VDD Switch_PMOS_n12_X1_Y1
xMMI24 net72 net81 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI28 net51 net63 net72 VDD Switch_PMOS_n12_X1_Y1
xMMI45 net97 net5 net101 VDD Switch_PMOS_n12_X1_Y1
xMMI7 net100 net63 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI21_M_u2 net81 CDN VDD VDD Switch_PMOS_n12_X1_Y1
.ends DFCNQD1

.subckt OAI21D0 A1 A2 B ZN
xMMI16_MI13 net9 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u9 ZN B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16_MI12 ZN A1 net9 VDD Switch_PMOS_n12_X1_Y1
xMM_u3 ZN A2 net24 VSS Switch_NMOS_n12_X1_Y1
xMM_u4 net24 B VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2 ZN A1 net24 VSS Switch_NMOS_n12_X1_Y1
.ends OAI21D0

.subckt OA211D0 A1 A2 B C Z
xMMI8 net17 B net20 VSS Switch_NMOS_n12_X1_Y1
xMMI11_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI9 net20 C VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u2 net5 A1 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI7 net5 A2 net17 VSS Switch_NMOS_n12_X1_Y1
xMMI4 net5 C VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net5 A2 net25 VDD Switch_PMOS_n12_X1_Y1
xMM_u12 net5 B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 net25 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI11_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends OA211D0

.subckt AO211D1 A1 A2 B C Z
xMM_u12 net5 C VSS VSS Switch_NMOS_n12_X1_Y1
xMMI8_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12_M_u10 net5 A1 net1 VSS Switch_NMOS_n12_X1_Y1
xMM_u13 net5 B VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12_M_u11 net1 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI16_MI12 net33 B net25 VDD Switch_PMOS_n12_X1_Y1
xMM_u3 net33 A1 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI0 net33 A2 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI16_MI13 net25 C VDD VDD Switch_PMOS_n12_X1_Y1
xMMI8_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AO211D1

.subckt MUX2ND0 I0 I1 S ZN
xMMI15_M_u3 net37 S VDD VDD Switch_PMOS_n12_X1_Y1
xMMI111 net13 I0 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI24 net9 I1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 ZN S net13 VDD Switch_PMOS_n12_X1_Y1
xMMI25 ZN net37 net9 VDD Switch_PMOS_n12_X1_Y1
xMMI15_M_u2 net37 S VSS VSS Switch_NMOS_n12_X1_Y1
xMMI20 net33 I1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI12 ZN net37 net32 VSS Switch_NMOS_n12_X1_Y1
xMMI21 ZN S net33 VSS Switch_NMOS_n12_X1_Y1
xMMI19 net32 I0 VSS VSS Switch_NMOS_n12_X1_Y1
.ends MUX2ND0

.subckt DFCNQD4 CDN CP D Q
xMMI22_M_u3 Q net123 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI38 net16 net123 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI32_M_u3 net79 net67 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI43 net61 net125 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI6 net9 D net1 VDD Switch_PMOS_n12_X1_Y1
xMMI31_M_u3 net67 CP VDD VDD Switch_PMOS_n12_X1_Y1
xMMI27_M_u3 Q net123 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI36_M_u2 net123 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI44 net61 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI36_M_u1 net123 net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI13_M_u3 net125 net9 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI24_M_u3 Q net123 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI16 net125 net67 net13 VDD Switch_PMOS_n12_X1_Y1
xMMI30_M_u1 net123 net13 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI30_M_u2 net123 CDN VDD VDD Switch_PMOS_n12_X1_Y1
xMMI28 net13 net79 net16 VDD Switch_PMOS_n12_X1_Y1
xMMI45 net9 net67 net61 VDD Switch_PMOS_n12_X1_Y1
xMMI25_M_u3 Q net123 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI7 net1 net79 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI24_M_u2 Q net123 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI30_M_u4 net145 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI4 net112 net67 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI13_M_u2 net125 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI30_M_u3 net123 net13 net145 VSS Switch_NMOS_n12_X1_Y1
xMMI29 net13 net67 net93 VSS Switch_NMOS_n12_X1_Y1
xMMI15 net125 net79 net13 VSS Switch_NMOS_n12_X1_Y1
xMMI25_M_u2 Q net123 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI36_M_u3 net123 net13 net97 VSS Switch_NMOS_n12_X1_Y1
xMMI32_M_u2 net79 net67 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net9 D net112 VSS Switch_NMOS_n12_X1_Y1
xMMI31_M_u2 net67 CP VSS VSS Switch_NMOS_n12_X1_Y1
xMMI49 net92 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI36_M_u4 net97 CDN VSS VSS Switch_NMOS_n12_X1_Y1
xMMI26 net93 net123 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI48 net80 net125 net92 VSS Switch_NMOS_n12_X1_Y1
xMMI27_M_u2 Q net123 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI22_M_u2 Q net123 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI47 net9 net79 net80 VSS Switch_NMOS_n12_X1_Y1
.ends DFCNQD4

.subckt AO22D1 A1 A2 B1 B2 Z
xMMI20_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI29 net13 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI22 net9 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI28 net5 A1 net13 VSS Switch_NMOS_n12_X1_Y1
xMMI21 net5 B1 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI17 net25 B1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI19 net5 A1 net25 VDD Switch_PMOS_n12_X1_Y1
xMMI18 net5 A2 net25 VDD Switch_PMOS_n12_X1_Y1
xMMI15 net25 B2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI20_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AO22D1

.subckt AOI22D1 A1 A2 B1 B2 ZN
xMMI3 ZN B1 net1 VSS Switch_NMOS_n12_X1_Y1
xMMI9 ZN A1 net5 VSS Switch_NMOS_n12_X1_Y1
xMMI10 net5 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI8 net1 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u3 net20 A2 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u5 VDD B2 net20 VDD Switch_PMOS_n12_X1_Y1
xMM_u2 net20 A1 ZN VDD Switch_PMOS_n12_X1_Y1
xMM_u4 VDD B1 net20 VDD Switch_PMOS_n12_X1_Y1
.ends AOI22D1

.subckt AOI222D0 A1 A2 B1 B2 C1 C2 ZN
xMMI17 net17 B1 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI16 net17 B2 net20 VDD Switch_PMOS_n12_X1_Y1
xMMI19 net20 A1 ZN VDD Switch_PMOS_n12_X1_Y1
xMMU27 VDD C2 net17 VDD Switch_PMOS_n12_X1_Y1
xMMI18 net20 A2 ZN VDD Switch_PMOS_n12_X1_Y1
xMMI15 VDD C1 net17 VDD Switch_PMOS_n12_X1_Y1
xMMI20_M_u10 ZN B1 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI6_M_u11 net40 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI6_M_u10 ZN A1 net40 VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u10 ZN C1 net36 VSS Switch_NMOS_n12_X1_Y1
xMMI21_M_u11 net36 C2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI20_M_u11 net25 B2 VSS VSS Switch_NMOS_n12_X1_Y1
.ends AOI222D0

.subckt AO221D1 A1 A2 B1 B2 C Z
xMMI1_M_u10 net5 A1 net9 VSS Switch_NMOS_n12_X1_Y1
xMMI17_M_u10 net5 B1 net20 VSS Switch_NMOS_n12_X1_Y1
xMMI8_M_u2 Z net5 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u11 net9 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU20 net5 C VSS VSS Switch_NMOS_n12_X1_Y1
xMMI17_M_u11 net20 B2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI5 net44 A1 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI2 net33 B2 net44 VDD Switch_PMOS_n12_X1_Y1
xMMU22 VDD C net33 VDD Switch_PMOS_n12_X1_Y1
xMMI3 net33 B1 net44 VDD Switch_PMOS_n12_X1_Y1
xMMI4 net44 A2 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI8_M_u3 Z net5 VDD VDD Switch_PMOS_n12_X1_Y1
.ends AO221D1

.subckt DCAP8 
xMMI4 VSS net9 VSS Dcap_NMOS_n12_X1_Y1
xMM_u2 net11 net9 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI3 VDD net11 VDD Dcap_PMOS_n12_X1_Y1
xMM_u1 net9 net11 VDD VDD Switch_PMOS_n12_X1_Y1
.ends DCAP8

.subckt Dcap_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_NMOS_n12_X1_Y1

.subckt Dcap_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Dcap_PMOS_n12_X1_Y1

.subckt SEL_LOGIC_V2 MDLCLK NDIV<5> NDIV<4> NDIV<3> NDIV<2> NDIV<1> NDIV<0> SEL SRST
XCYLCNT0REG010 SRST MDLCLK N1 CYLCNT<1> VDD VSS DFCNQD1
XCYLCNT0REG020 SRST MDLCLK N2 CYLCNT<2> VDD VSS DFCNQD1
XCYLCNT0REG030 SRST MDLCLK N3 CYLCNT<3> VDD VSS DFCNQD1
XCYLCNT0REG040 SRST MDLCLK N4 CYLCNT<4> VDD VSS DFCNQD1
XCYLCNT0REG050 SRST MDLCLK N5 CYLCNT<5> VDD VSS DFCNQD1
XCYLCNT0REG000 SRST MDLCLK N14 CYLCNT<0> VDD VSS DFCNQD1
XU22 CYLCNT<0> VDD VSS N14 INVD1
XU5 N15 N16 N17 SEL VDD VSS N10 OA31D1
XU11 NDIV<4> CYLCNT<4> VDD VSS N20 XNR2D1
XU12 NDIV<2> CYLCNT<2> VDD VSS N19 XNR2D1
XU13 NDIV<5> CYLCNT<5> VDD VSS N18 XNR2D1
XU16 NDIV<3> CYLCNT<3> VDD VSS N21 XNR2D1
XU15 NDIV<1> CYLCNT<1> VDD VSS N22 XNR2D1
XU17 NDIV<0> N14 VDD VSS N15 XNR2D1
XSEL0REG MDLCLK N10 SEL SRST VDD VSS DFSNQD1
XU20 N21 N22 VDD VSS N16 ND2D1
XU6 CYLCNT<1> CYLCNT<0> ADD0190CARRY020 N1 VDD VSS HA1D0
XU7 CYLCNT<3> ADD0190CARRY030 ADD0190CARRY040 N3 VDD VSS HA1D0
XU8 CYLCNT<2> ADD0190CARRY020 ADD0190CARRY030 N2 VDD VSS HA1D0
XU9 CYLCNT<4> ADD0190CARRY040 ADD0190CARRY050 N4 VDD VSS HA1D0
XU18 ADD0190CARRY050 CYLCNT<5> VDD VSS N5 CKXOR2D1
XU21 N18 N19 N20 VDD VSS N17 ND3D1
.ends SEL_LOGIC_V2

.subckt OA31D1 A1 A2 A3 B Z
xMMU1_M_u2 Z net25 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI6 net5 A1 net25 VSS Switch_NMOS_n12_X1_Y1
xMM_u5 VSS B net5 VSS Switch_NMOS_n12_X1_Y1
xMMI8 net5 A3 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI7 net5 A2 net25 VSS Switch_NMOS_n12_X1_Y1
xMMI3 net37 A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI4 net33 A2 net37 VDD Switch_PMOS_n12_X1_Y1
xMMU1_M_u3 Z net25 VDD VDD Switch_PMOS_n12_X1_Y1
xMM_u11 net25 B VDD VDD Switch_PMOS_n12_X1_Y1
xMMI5 net25 A3 net33 VDD Switch_PMOS_n12_X1_Y1
.ends OA31D1
