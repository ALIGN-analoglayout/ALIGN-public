VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

 
MACRO CAP_MIM_wt32_lt32
  ORIGIN 0 0 ;
  FOREIGN CAP_MIM_wt32_lt32 0 0 ;
  SIZE 52.8 BY 56.8 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
        RECT 8.4 12.8 9.52 44.16 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
        RECT 43.12 11.52 44.24 45.44 ;
    END
  END MINUS
  OBS
    LAYER M7 ;
      RECT 7 6.96 46 49 ;
    LAYER M8 ;
      RECT 10 10 42.8 46.8 ;
  END
END CAP_MIM_wt32_lt32

END LIBRARY
