MACRO switched_capacitor_combination
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_combination 0 0 ;
  SIZE 15.52 BY 29.904 ;
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.46 0.384 10.5 0.708 ;
      LAYER M3 ;
        RECT 10.22 0.384 10.26 0.708 ;
      LAYER M2 ;
        RECT 9.564 0.488 9.796 0.52 ;
      LAYER M2 ;
        RECT 7.724 0.488 7.956 0.52 ;
      LAYER M3 ;
        RECT 10.46 0.484 10.5 0.524 ;
      LAYER M4 ;
        RECT 10 0.484 10.48 0.524 ;
      LAYER M3 ;
        RECT 9.98 0.484 10.02 0.524 ;
      LAYER M2 ;
        RECT 9.76 0.488 10 0.52 ;
      LAYER M2 ;
        RECT 7.92 0.488 9.6 0.52 ;
    END
  END phi2
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.62 0.552 10.66 0.876 ;
      LAYER M3 ;
        RECT 10.38 0.552 10.42 0.876 ;
      LAYER M2 ;
        RECT 9.644 0.656 9.876 0.688 ;
      LAYER M2 ;
        RECT 7.644 0.656 7.876 0.688 ;
      LAYER M3 ;
        RECT 10.38 0.652 10.42 0.692 ;
      LAYER M4 ;
        RECT 10.08 0.652 10.4 0.692 ;
      LAYER M3 ;
        RECT 10.06 0.652 10.1 0.692 ;
      LAYER M2 ;
        RECT 9.84 0.656 10.08 0.688 ;
      LAYER M2 ;
        RECT 7.76 0.656 9.68 0.688 ;
    END
  END agnd
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.38 17.436 0.42 17.76 ;
      LAYER M3 ;
        RECT 0.14 17.436 0.18 17.76 ;
      LAYER M2 ;
        RECT 9.084 0.572 9.316 0.604 ;
      LAYER M2 ;
        RECT 8.204 0.572 8.436 0.604 ;
      LAYER M3 ;
        RECT 0.38 10.416 0.42 17.472 ;
      LAYER M2 ;
        RECT 0.4 10.4 8.32 10.432 ;
      LAYER M3 ;
        RECT 8.3 0.588 8.34 10.416 ;
      LAYER M2 ;
        RECT 8.304 0.572 8.336 0.604 ;
      LAYER M2 ;
        RECT 8.4 0.572 9.12 0.604 ;
    END
  END phi1
  PIN Vin
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.54 17.604 0.58 17.928 ;
      LAYER M3 ;
        RECT 0.3 17.604 0.34 17.928 ;
    END
  END Vin
  PIN Vin_ota
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.164 0.74 9.396 0.772 ;
      LAYER M1 ;
        RECT 3.664 16.764 3.696 16.836 ;
      LAYER M2 ;
        RECT 3.644 16.784 3.716 16.816 ;
      LAYER M1 ;
        RECT 12.304 16.764 12.336 16.836 ;
      LAYER M2 ;
        RECT 12.284 16.784 12.356 16.816 ;
      LAYER M2 ;
        RECT 3.68 16.784 12.32 16.816 ;
      LAYER M2 ;
        RECT 8.96 0.74 9.2 0.772 ;
      LAYER M3 ;
        RECT 8.94 0.756 8.98 16.128 ;
      LAYER M4 ;
        RECT 8.64 16.108 8.96 16.148 ;
      LAYER M5 ;
        RECT 8.608 16.128 8.672 16.548 ;
      LAYER M4 ;
        RECT 8.62 16.528 8.66 16.568 ;
      LAYER M3 ;
        RECT 8.62 16.548 8.66 16.8 ;
      LAYER M2 ;
        RECT 8.624 16.784 8.656 16.816 ;
    END
  END Vin_ota
  PIN Voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.124 0.74 8.356 0.772 ;
      LAYER M1 ;
        RECT 3.824 1.224 3.856 1.296 ;
      LAYER M2 ;
        RECT 3.804 1.244 3.876 1.276 ;
      LAYER M1 ;
        RECT 12.464 1.224 12.496 1.296 ;
      LAYER M2 ;
        RECT 12.444 1.244 12.516 1.276 ;
      LAYER M2 ;
        RECT 3.84 1.244 12.48 1.276 ;
      LAYER M2 ;
        RECT 8.144 0.74 8.176 0.772 ;
      LAYER M3 ;
        RECT 8.14 0.756 8.18 1.26 ;
      LAYER M2 ;
        RECT 8.144 1.244 8.176 1.276 ;
    END
  END Voutn
  OBS 
  LAYER M1 ;
        RECT 9.344 29.616 9.376 29.688 ;
  LAYER M2 ;
        RECT 9.324 29.636 9.396 29.668 ;
  LAYER M1 ;
        RECT 6.464 29.616 6.496 29.688 ;
  LAYER M2 ;
        RECT 6.444 29.636 6.516 29.668 ;
  LAYER M2 ;
        RECT 6.48 29.636 9.36 29.668 ;
  LAYER M2 ;
        RECT 9.004 0.824 9.716 0.856 ;
  LAYER M1 ;
        RECT 6.544 16.596 6.576 16.668 ;
  LAYER M2 ;
        RECT 6.524 16.616 6.596 16.648 ;
  LAYER M1 ;
        RECT 9.424 16.596 9.456 16.668 ;
  LAYER M2 ;
        RECT 9.404 16.616 9.476 16.648 ;
  LAYER M2 ;
        RECT 6.56 16.616 9.44 16.648 ;
  LAYER M2 ;
        RECT 7.184 29.636 7.216 29.668 ;
  LAYER M3 ;
        RECT 7.18 29.4 7.22 29.652 ;
  LAYER M4 ;
        RECT 7.18 29.38 7.22 29.42 ;
  LAYER M5 ;
        RECT 7.168 16.884 7.232 29.4 ;
  LAYER M4 ;
        RECT 7.18 16.864 7.22 16.904 ;
  LAYER M3 ;
        RECT 7.18 16.632 7.22 16.884 ;
  LAYER M2 ;
        RECT 7.184 16.616 7.216 16.648 ;
  LAYER M2 ;
        RECT 9.344 16.616 9.376 16.648 ;
  LAYER M3 ;
        RECT 9.34 1.512 9.38 16.632 ;
  LAYER M4 ;
        RECT 9.34 1.492 9.38 1.532 ;
  LAYER M5 ;
        RECT 9.328 1.344 9.392 1.512 ;
  LAYER M4 ;
        RECT 9.34 1.324 9.38 1.364 ;
  LAYER M3 ;
        RECT 9.34 0.84 9.38 1.344 ;
  LAYER M2 ;
        RECT 9.344 0.824 9.376 0.856 ;
  LAYER M1 ;
        RECT 9.504 17.352 9.536 17.424 ;
  LAYER M2 ;
        RECT 9.484 17.372 9.556 17.404 ;
  LAYER M1 ;
        RECT 6.624 17.352 6.656 17.424 ;
  LAYER M2 ;
        RECT 6.604 17.372 6.676 17.404 ;
  LAYER M2 ;
        RECT 6.64 17.372 9.52 17.404 ;
  LAYER M3 ;
        RECT 10.54 0.468 10.58 0.792 ;
  LAYER M3 ;
        RECT 10.3 0.468 10.34 0.792 ;
  LAYER M3 ;
        RECT 0.46 17.52 0.5 17.844 ;
  LAYER M3 ;
        RECT 0.22 17.52 0.26 17.844 ;
  LAYER M2 ;
        RECT 0.48 17.372 6.72 17.404 ;
  LAYER M3 ;
        RECT 0.46 17.388 0.5 17.64 ;
  LAYER M2 ;
        RECT 9.504 17.372 9.536 17.404 ;
  LAYER M3 ;
        RECT 9.5 0.756 9.54 17.388 ;
  LAYER M4 ;
        RECT 9.52 0.736 10.32 0.776 ;
  LAYER M3 ;
        RECT 10.3 0.736 10.34 0.776 ;
  LAYER M2 ;
        RECT 7.804 0.824 8.516 0.856 ;
  LAYER M1 ;
        RECT 6.704 1.392 6.736 1.464 ;
  LAYER M2 ;
        RECT 6.684 1.412 6.756 1.444 ;
  LAYER M1 ;
        RECT 9.584 1.392 9.616 1.464 ;
  LAYER M2 ;
        RECT 9.564 1.412 9.636 1.444 ;
  LAYER M2 ;
        RECT 6.72 1.412 9.6 1.444 ;
  LAYER M2 ;
        RECT 7.904 0.824 7.936 0.856 ;
  LAYER M3 ;
        RECT 7.9 0.84 7.94 1.344 ;
  LAYER M4 ;
        RECT 7.9 1.324 7.94 1.364 ;
  LAYER M5 ;
        RECT 7.888 1.344 7.952 1.428 ;
  LAYER M4 ;
        RECT 7.9 1.408 7.94 1.448 ;
  LAYER M3 ;
        RECT 7.9 1.408 7.94 1.448 ;
  LAYER M2 ;
        RECT 7.904 1.412 7.936 1.444 ;
  LAYER M1 ;
        RECT 9.184 20.796 9.216 20.868 ;
  LAYER M2 ;
        RECT 9.164 20.816 9.236 20.848 ;
  LAYER M2 ;
        RECT 9.2 20.816 9.52 20.848 ;
  LAYER M1 ;
        RECT 9.504 20.796 9.536 20.868 ;
  LAYER M2 ;
        RECT 9.484 20.816 9.556 20.848 ;
  LAYER M1 ;
        RECT 9.184 23.736 9.216 23.808 ;
  LAYER M2 ;
        RECT 9.164 23.756 9.236 23.788 ;
  LAYER M2 ;
        RECT 9.2 23.756 9.52 23.788 ;
  LAYER M1 ;
        RECT 9.504 23.736 9.536 23.808 ;
  LAYER M2 ;
        RECT 9.484 23.756 9.556 23.788 ;
  LAYER M1 ;
        RECT 12.064 20.796 12.096 20.868 ;
  LAYER M2 ;
        RECT 12.044 20.816 12.116 20.848 ;
  LAYER M1 ;
        RECT 12.064 20.664 12.096 20.832 ;
  LAYER M1 ;
        RECT 12.064 20.628 12.096 20.7 ;
  LAYER M2 ;
        RECT 12.044 20.648 12.116 20.68 ;
  LAYER M2 ;
        RECT 9.52 20.648 12.08 20.68 ;
  LAYER M1 ;
        RECT 9.504 20.628 9.536 20.7 ;
  LAYER M2 ;
        RECT 9.484 20.648 9.556 20.68 ;
  LAYER M1 ;
        RECT 12.064 23.736 12.096 23.808 ;
  LAYER M2 ;
        RECT 12.044 23.756 12.116 23.788 ;
  LAYER M1 ;
        RECT 12.064 23.604 12.096 23.772 ;
  LAYER M1 ;
        RECT 12.064 23.568 12.096 23.64 ;
  LAYER M2 ;
        RECT 12.044 23.588 12.116 23.62 ;
  LAYER M2 ;
        RECT 9.52 23.588 12.08 23.62 ;
  LAYER M1 ;
        RECT 9.504 23.568 9.536 23.64 ;
  LAYER M2 ;
        RECT 9.484 23.588 9.556 23.62 ;
  LAYER M1 ;
        RECT 9.504 17.352 9.536 17.424 ;
  LAYER M2 ;
        RECT 9.484 17.372 9.556 17.404 ;
  LAYER M1 ;
        RECT 9.504 17.388 9.536 17.556 ;
  LAYER M1 ;
        RECT 9.504 17.556 9.536 23.772 ;
  LAYER M1 ;
        RECT 6.304 23.736 6.336 23.808 ;
  LAYER M2 ;
        RECT 6.284 23.756 6.356 23.788 ;
  LAYER M2 ;
        RECT 6.32 23.756 6.64 23.788 ;
  LAYER M1 ;
        RECT 6.624 23.736 6.656 23.808 ;
  LAYER M2 ;
        RECT 6.604 23.756 6.676 23.788 ;
  LAYER M1 ;
        RECT 6.304 20.796 6.336 20.868 ;
  LAYER M2 ;
        RECT 6.284 20.816 6.356 20.848 ;
  LAYER M2 ;
        RECT 6.32 20.816 6.64 20.848 ;
  LAYER M1 ;
        RECT 6.624 20.796 6.656 20.868 ;
  LAYER M2 ;
        RECT 6.604 20.816 6.676 20.848 ;
  LAYER M1 ;
        RECT 6.624 17.352 6.656 17.424 ;
  LAYER M2 ;
        RECT 6.604 17.372 6.676 17.404 ;
  LAYER M1 ;
        RECT 6.624 17.388 6.656 17.556 ;
  LAYER M1 ;
        RECT 6.624 17.556 6.656 23.772 ;
  LAYER M2 ;
        RECT 6.64 17.372 9.52 17.404 ;
  LAYER M1 ;
        RECT 14.944 17.856 14.976 17.928 ;
  LAYER M2 ;
        RECT 14.924 17.876 14.996 17.908 ;
  LAYER M1 ;
        RECT 14.944 17.724 14.976 17.892 ;
  LAYER M1 ;
        RECT 14.944 17.688 14.976 17.76 ;
  LAYER M2 ;
        RECT 14.924 17.708 14.996 17.74 ;
  LAYER M2 ;
        RECT 12.4 17.708 14.96 17.74 ;
  LAYER M1 ;
        RECT 12.384 17.688 12.416 17.76 ;
  LAYER M2 ;
        RECT 12.364 17.708 12.436 17.74 ;
  LAYER M1 ;
        RECT 14.944 20.796 14.976 20.868 ;
  LAYER M2 ;
        RECT 14.924 20.816 14.996 20.848 ;
  LAYER M1 ;
        RECT 14.944 20.664 14.976 20.832 ;
  LAYER M1 ;
        RECT 14.944 20.628 14.976 20.7 ;
  LAYER M2 ;
        RECT 14.924 20.648 14.996 20.68 ;
  LAYER M2 ;
        RECT 12.4 20.648 14.96 20.68 ;
  LAYER M1 ;
        RECT 12.384 20.628 12.416 20.7 ;
  LAYER M2 ;
        RECT 12.364 20.648 12.436 20.68 ;
  LAYER M1 ;
        RECT 14.944 23.736 14.976 23.808 ;
  LAYER M2 ;
        RECT 14.924 23.756 14.996 23.788 ;
  LAYER M1 ;
        RECT 14.944 23.604 14.976 23.772 ;
  LAYER M1 ;
        RECT 14.944 23.568 14.976 23.64 ;
  LAYER M2 ;
        RECT 14.924 23.588 14.996 23.62 ;
  LAYER M2 ;
        RECT 12.4 23.588 14.96 23.62 ;
  LAYER M1 ;
        RECT 12.384 23.568 12.416 23.64 ;
  LAYER M2 ;
        RECT 12.364 23.588 12.436 23.62 ;
  LAYER M1 ;
        RECT 14.944 26.676 14.976 26.748 ;
  LAYER M2 ;
        RECT 14.924 26.696 14.996 26.728 ;
  LAYER M1 ;
        RECT 14.944 26.544 14.976 26.712 ;
  LAYER M1 ;
        RECT 14.944 26.508 14.976 26.58 ;
  LAYER M2 ;
        RECT 14.924 26.528 14.996 26.56 ;
  LAYER M2 ;
        RECT 12.4 26.528 14.96 26.56 ;
  LAYER M1 ;
        RECT 12.384 26.508 12.416 26.58 ;
  LAYER M2 ;
        RECT 12.364 26.528 12.436 26.56 ;
  LAYER M1 ;
        RECT 12.064 17.856 12.096 17.928 ;
  LAYER M2 ;
        RECT 12.044 17.876 12.116 17.908 ;
  LAYER M2 ;
        RECT 12.08 17.876 12.4 17.908 ;
  LAYER M1 ;
        RECT 12.384 17.856 12.416 17.928 ;
  LAYER M2 ;
        RECT 12.364 17.876 12.436 17.908 ;
  LAYER M1 ;
        RECT 12.064 26.676 12.096 26.748 ;
  LAYER M2 ;
        RECT 12.044 26.696 12.116 26.728 ;
  LAYER M2 ;
        RECT 12.08 26.696 12.4 26.728 ;
  LAYER M1 ;
        RECT 12.384 26.676 12.416 26.748 ;
  LAYER M2 ;
        RECT 12.364 26.696 12.436 26.728 ;
  LAYER M1 ;
        RECT 12.384 17.184 12.416 17.256 ;
  LAYER M2 ;
        RECT 12.364 17.204 12.436 17.236 ;
  LAYER M1 ;
        RECT 12.384 17.22 12.416 17.556 ;
  LAYER M1 ;
        RECT 12.384 17.556 12.416 26.712 ;
  LAYER M1 ;
        RECT 6.304 17.856 6.336 17.928 ;
  LAYER M2 ;
        RECT 6.284 17.876 6.356 17.908 ;
  LAYER M1 ;
        RECT 6.304 17.724 6.336 17.892 ;
  LAYER M1 ;
        RECT 6.304 17.688 6.336 17.76 ;
  LAYER M2 ;
        RECT 6.284 17.708 6.356 17.74 ;
  LAYER M2 ;
        RECT 3.76 17.708 6.32 17.74 ;
  LAYER M1 ;
        RECT 3.744 17.688 3.776 17.76 ;
  LAYER M2 ;
        RECT 3.724 17.708 3.796 17.74 ;
  LAYER M1 ;
        RECT 6.304 26.676 6.336 26.748 ;
  LAYER M2 ;
        RECT 6.284 26.696 6.356 26.728 ;
  LAYER M1 ;
        RECT 6.304 26.544 6.336 26.712 ;
  LAYER M1 ;
        RECT 6.304 26.508 6.336 26.58 ;
  LAYER M2 ;
        RECT 6.284 26.528 6.356 26.56 ;
  LAYER M2 ;
        RECT 3.76 26.528 6.32 26.56 ;
  LAYER M1 ;
        RECT 3.744 26.508 3.776 26.58 ;
  LAYER M2 ;
        RECT 3.724 26.528 3.796 26.56 ;
  LAYER M1 ;
        RECT 3.424 17.856 3.456 17.928 ;
  LAYER M2 ;
        RECT 3.404 17.876 3.476 17.908 ;
  LAYER M2 ;
        RECT 3.44 17.876 3.76 17.908 ;
  LAYER M1 ;
        RECT 3.744 17.856 3.776 17.928 ;
  LAYER M2 ;
        RECT 3.724 17.876 3.796 17.908 ;
  LAYER M1 ;
        RECT 3.424 20.796 3.456 20.868 ;
  LAYER M2 ;
        RECT 3.404 20.816 3.476 20.848 ;
  LAYER M2 ;
        RECT 3.44 20.816 3.76 20.848 ;
  LAYER M1 ;
        RECT 3.744 20.796 3.776 20.868 ;
  LAYER M2 ;
        RECT 3.724 20.816 3.796 20.848 ;
  LAYER M1 ;
        RECT 3.424 23.736 3.456 23.808 ;
  LAYER M2 ;
        RECT 3.404 23.756 3.476 23.788 ;
  LAYER M2 ;
        RECT 3.44 23.756 3.76 23.788 ;
  LAYER M1 ;
        RECT 3.744 23.736 3.776 23.808 ;
  LAYER M2 ;
        RECT 3.724 23.756 3.796 23.788 ;
  LAYER M1 ;
        RECT 3.424 26.676 3.456 26.748 ;
  LAYER M2 ;
        RECT 3.404 26.696 3.476 26.728 ;
  LAYER M2 ;
        RECT 3.44 26.696 3.76 26.728 ;
  LAYER M1 ;
        RECT 3.744 26.676 3.776 26.748 ;
  LAYER M2 ;
        RECT 3.724 26.696 3.796 26.728 ;
  LAYER M1 ;
        RECT 3.744 17.184 3.776 17.256 ;
  LAYER M2 ;
        RECT 3.724 17.204 3.796 17.236 ;
  LAYER M1 ;
        RECT 3.744 17.22 3.776 17.556 ;
  LAYER M1 ;
        RECT 3.744 17.556 3.776 26.712 ;
  LAYER M2 ;
        RECT 3.76 17.204 12.4 17.236 ;
  LAYER M1 ;
        RECT 9.184 26.676 9.216 26.748 ;
  LAYER M2 ;
        RECT 9.164 26.696 9.236 26.728 ;
  LAYER M2 ;
        RECT 9.2 26.696 12.08 26.728 ;
  LAYER M1 ;
        RECT 12.064 26.676 12.096 26.748 ;
  LAYER M2 ;
        RECT 12.044 26.696 12.116 26.728 ;
  LAYER M1 ;
        RECT 9.184 17.856 9.216 17.928 ;
  LAYER M2 ;
        RECT 9.164 17.876 9.236 17.908 ;
  LAYER M2 ;
        RECT 6.32 17.876 9.2 17.908 ;
  LAYER M1 ;
        RECT 6.304 17.856 6.336 17.928 ;
  LAYER M2 ;
        RECT 6.284 17.876 6.356 17.908 ;
  LAYER M1 ;
        RECT 6.784 23.232 6.816 23.304 ;
  LAYER M2 ;
        RECT 6.764 23.252 6.836 23.284 ;
  LAYER M2 ;
        RECT 6.8 23.252 9.36 23.284 ;
  LAYER M1 ;
        RECT 9.344 23.232 9.376 23.304 ;
  LAYER M2 ;
        RECT 9.324 23.252 9.396 23.284 ;
  LAYER M1 ;
        RECT 6.784 26.172 6.816 26.244 ;
  LAYER M2 ;
        RECT 6.764 26.192 6.836 26.224 ;
  LAYER M2 ;
        RECT 6.8 26.192 9.36 26.224 ;
  LAYER M1 ;
        RECT 9.344 26.172 9.376 26.244 ;
  LAYER M2 ;
        RECT 9.324 26.192 9.396 26.224 ;
  LAYER M1 ;
        RECT 9.664 23.232 9.696 23.304 ;
  LAYER M2 ;
        RECT 9.644 23.252 9.716 23.284 ;
  LAYER M1 ;
        RECT 9.664 23.268 9.696 23.436 ;
  LAYER M1 ;
        RECT 9.664 23.4 9.696 23.472 ;
  LAYER M2 ;
        RECT 9.644 23.42 9.716 23.452 ;
  LAYER M2 ;
        RECT 9.36 23.42 9.68 23.452 ;
  LAYER M1 ;
        RECT 9.344 23.4 9.376 23.472 ;
  LAYER M2 ;
        RECT 9.324 23.42 9.396 23.452 ;
  LAYER M1 ;
        RECT 9.664 26.172 9.696 26.244 ;
  LAYER M2 ;
        RECT 9.644 26.192 9.716 26.224 ;
  LAYER M1 ;
        RECT 9.664 26.208 9.696 26.376 ;
  LAYER M1 ;
        RECT 9.664 26.34 9.696 26.412 ;
  LAYER M2 ;
        RECT 9.644 26.36 9.716 26.392 ;
  LAYER M2 ;
        RECT 9.36 26.36 9.68 26.392 ;
  LAYER M1 ;
        RECT 9.344 26.34 9.376 26.412 ;
  LAYER M2 ;
        RECT 9.324 26.36 9.396 26.392 ;
  LAYER M1 ;
        RECT 9.344 29.616 9.376 29.688 ;
  LAYER M2 ;
        RECT 9.324 29.636 9.396 29.668 ;
  LAYER M1 ;
        RECT 9.344 29.484 9.376 29.652 ;
  LAYER M1 ;
        RECT 9.344 23.268 9.376 29.484 ;
  LAYER M1 ;
        RECT 3.904 26.172 3.936 26.244 ;
  LAYER M2 ;
        RECT 3.884 26.192 3.956 26.224 ;
  LAYER M2 ;
        RECT 3.92 26.192 6.48 26.224 ;
  LAYER M1 ;
        RECT 6.464 26.172 6.496 26.244 ;
  LAYER M2 ;
        RECT 6.444 26.192 6.516 26.224 ;
  LAYER M1 ;
        RECT 3.904 23.232 3.936 23.304 ;
  LAYER M2 ;
        RECT 3.884 23.252 3.956 23.284 ;
  LAYER M2 ;
        RECT 3.92 23.252 6.48 23.284 ;
  LAYER M1 ;
        RECT 6.464 23.232 6.496 23.304 ;
  LAYER M2 ;
        RECT 6.444 23.252 6.516 23.284 ;
  LAYER M1 ;
        RECT 6.464 29.616 6.496 29.688 ;
  LAYER M2 ;
        RECT 6.444 29.636 6.516 29.668 ;
  LAYER M1 ;
        RECT 6.464 29.484 6.496 29.652 ;
  LAYER M1 ;
        RECT 6.464 23.268 6.496 29.484 ;
  LAYER M2 ;
        RECT 6.48 29.636 9.36 29.668 ;
  LAYER M1 ;
        RECT 12.544 20.292 12.576 20.364 ;
  LAYER M2 ;
        RECT 12.524 20.312 12.596 20.344 ;
  LAYER M2 ;
        RECT 12.56 20.312 15.28 20.344 ;
  LAYER M1 ;
        RECT 15.264 20.292 15.296 20.364 ;
  LAYER M2 ;
        RECT 15.244 20.312 15.316 20.344 ;
  LAYER M1 ;
        RECT 12.544 23.232 12.576 23.304 ;
  LAYER M2 ;
        RECT 12.524 23.252 12.596 23.284 ;
  LAYER M2 ;
        RECT 12.56 23.252 15.28 23.284 ;
  LAYER M1 ;
        RECT 15.264 23.232 15.296 23.304 ;
  LAYER M2 ;
        RECT 15.244 23.252 15.316 23.284 ;
  LAYER M1 ;
        RECT 12.544 26.172 12.576 26.244 ;
  LAYER M2 ;
        RECT 12.524 26.192 12.596 26.224 ;
  LAYER M2 ;
        RECT 12.56 26.192 15.28 26.224 ;
  LAYER M1 ;
        RECT 15.264 26.172 15.296 26.244 ;
  LAYER M2 ;
        RECT 15.244 26.192 15.316 26.224 ;
  LAYER M1 ;
        RECT 12.544 29.112 12.576 29.184 ;
  LAYER M2 ;
        RECT 12.524 29.132 12.596 29.164 ;
  LAYER M2 ;
        RECT 12.56 29.132 15.28 29.164 ;
  LAYER M1 ;
        RECT 15.264 29.112 15.296 29.184 ;
  LAYER M2 ;
        RECT 15.244 29.132 15.316 29.164 ;
  LAYER M1 ;
        RECT 15.264 29.784 15.296 29.856 ;
  LAYER M2 ;
        RECT 15.244 29.804 15.316 29.836 ;
  LAYER M1 ;
        RECT 15.264 29.484 15.296 29.82 ;
  LAYER M1 ;
        RECT 15.264 20.328 15.296 29.484 ;
  LAYER M1 ;
        RECT 1.024 20.292 1.056 20.364 ;
  LAYER M2 ;
        RECT 1.004 20.312 1.076 20.344 ;
  LAYER M1 ;
        RECT 1.024 20.328 1.056 20.496 ;
  LAYER M1 ;
        RECT 1.024 20.46 1.056 20.532 ;
  LAYER M2 ;
        RECT 1.004 20.48 1.076 20.512 ;
  LAYER M2 ;
        RECT 0.88 20.48 1.04 20.512 ;
  LAYER M1 ;
        RECT 0.864 20.46 0.896 20.532 ;
  LAYER M2 ;
        RECT 0.844 20.48 0.916 20.512 ;
  LAYER M1 ;
        RECT 1.024 23.232 1.056 23.304 ;
  LAYER M2 ;
        RECT 1.004 23.252 1.076 23.284 ;
  LAYER M1 ;
        RECT 1.024 23.268 1.056 23.436 ;
  LAYER M1 ;
        RECT 1.024 23.4 1.056 23.472 ;
  LAYER M2 ;
        RECT 1.004 23.42 1.076 23.452 ;
  LAYER M2 ;
        RECT 0.88 23.42 1.04 23.452 ;
  LAYER M1 ;
        RECT 0.864 23.4 0.896 23.472 ;
  LAYER M2 ;
        RECT 0.844 23.42 0.916 23.452 ;
  LAYER M1 ;
        RECT 1.024 26.172 1.056 26.244 ;
  LAYER M2 ;
        RECT 1.004 26.192 1.076 26.224 ;
  LAYER M1 ;
        RECT 1.024 26.208 1.056 26.376 ;
  LAYER M1 ;
        RECT 1.024 26.34 1.056 26.412 ;
  LAYER M2 ;
        RECT 1.004 26.36 1.076 26.392 ;
  LAYER M2 ;
        RECT 0.88 26.36 1.04 26.392 ;
  LAYER M1 ;
        RECT 0.864 26.34 0.896 26.412 ;
  LAYER M2 ;
        RECT 0.844 26.36 0.916 26.392 ;
  LAYER M1 ;
        RECT 1.024 29.112 1.056 29.184 ;
  LAYER M2 ;
        RECT 1.004 29.132 1.076 29.164 ;
  LAYER M1 ;
        RECT 1.024 29.148 1.056 29.316 ;
  LAYER M1 ;
        RECT 1.024 29.28 1.056 29.352 ;
  LAYER M2 ;
        RECT 1.004 29.3 1.076 29.332 ;
  LAYER M2 ;
        RECT 0.88 29.3 1.04 29.332 ;
  LAYER M1 ;
        RECT 0.864 29.28 0.896 29.352 ;
  LAYER M2 ;
        RECT 0.844 29.3 0.916 29.332 ;
  LAYER M1 ;
        RECT 0.864 29.784 0.896 29.856 ;
  LAYER M2 ;
        RECT 0.844 29.804 0.916 29.836 ;
  LAYER M1 ;
        RECT 0.864 29.484 0.896 29.82 ;
  LAYER M1 ;
        RECT 0.864 20.496 0.896 29.484 ;
  LAYER M2 ;
        RECT 0.88 29.804 15.28 29.836 ;
  LAYER M1 ;
        RECT 9.664 20.292 9.696 20.364 ;
  LAYER M2 ;
        RECT 9.644 20.312 9.716 20.344 ;
  LAYER M2 ;
        RECT 9.68 20.312 12.56 20.344 ;
  LAYER M1 ;
        RECT 12.544 20.292 12.576 20.364 ;
  LAYER M2 ;
        RECT 12.524 20.312 12.596 20.344 ;
  LAYER M1 ;
        RECT 9.664 29.112 9.696 29.184 ;
  LAYER M2 ;
        RECT 9.644 29.132 9.716 29.164 ;
  LAYER M2 ;
        RECT 9.68 29.132 12.56 29.164 ;
  LAYER M1 ;
        RECT 12.544 29.112 12.576 29.184 ;
  LAYER M2 ;
        RECT 12.524 29.132 12.596 29.164 ;
  LAYER M1 ;
        RECT 6.784 29.112 6.816 29.184 ;
  LAYER M2 ;
        RECT 6.764 29.132 6.836 29.164 ;
  LAYER M2 ;
        RECT 6.8 29.132 9.68 29.164 ;
  LAYER M1 ;
        RECT 9.664 29.112 9.696 29.184 ;
  LAYER M2 ;
        RECT 9.644 29.132 9.716 29.164 ;
  LAYER M1 ;
        RECT 3.904 29.112 3.936 29.184 ;
  LAYER M2 ;
        RECT 3.884 29.132 3.956 29.164 ;
  LAYER M2 ;
        RECT 3.92 29.132 6.8 29.164 ;
  LAYER M1 ;
        RECT 6.784 29.112 6.816 29.184 ;
  LAYER M2 ;
        RECT 6.764 29.132 6.836 29.164 ;
  LAYER M1 ;
        RECT 3.904 20.292 3.936 20.364 ;
  LAYER M2 ;
        RECT 3.884 20.312 3.956 20.344 ;
  LAYER M2 ;
        RECT 1.04 20.312 3.92 20.344 ;
  LAYER M1 ;
        RECT 1.024 20.292 1.056 20.364 ;
  LAYER M2 ;
        RECT 1.004 20.312 1.076 20.344 ;
  LAYER M1 ;
        RECT 6.784 20.292 6.816 20.364 ;
  LAYER M2 ;
        RECT 6.764 20.312 6.836 20.344 ;
  LAYER M2 ;
        RECT 3.92 20.312 6.8 20.344 ;
  LAYER M1 ;
        RECT 3.904 20.292 3.936 20.364 ;
  LAYER M2 ;
        RECT 3.884 20.312 3.956 20.344 ;
  LAYER M1 ;
        RECT 14.944 17.856 14.976 20.364 ;
  LAYER M1 ;
        RECT 14.88 17.856 14.912 20.364 ;
  LAYER M1 ;
        RECT 14.816 17.856 14.848 20.364 ;
  LAYER M1 ;
        RECT 14.752 17.856 14.784 20.364 ;
  LAYER M1 ;
        RECT 14.688 17.856 14.72 20.364 ;
  LAYER M1 ;
        RECT 14.624 17.856 14.656 20.364 ;
  LAYER M1 ;
        RECT 14.56 17.856 14.592 20.364 ;
  LAYER M1 ;
        RECT 14.496 17.856 14.528 20.364 ;
  LAYER M1 ;
        RECT 14.432 17.856 14.464 20.364 ;
  LAYER M1 ;
        RECT 14.368 17.856 14.4 20.364 ;
  LAYER M1 ;
        RECT 14.304 17.856 14.336 20.364 ;
  LAYER M1 ;
        RECT 14.24 17.856 14.272 20.364 ;
  LAYER M1 ;
        RECT 14.176 17.856 14.208 20.364 ;
  LAYER M1 ;
        RECT 14.112 17.856 14.144 20.364 ;
  LAYER M1 ;
        RECT 14.048 17.856 14.08 20.364 ;
  LAYER M1 ;
        RECT 13.984 17.856 14.016 20.364 ;
  LAYER M1 ;
        RECT 13.92 17.856 13.952 20.364 ;
  LAYER M1 ;
        RECT 13.856 17.856 13.888 20.364 ;
  LAYER M1 ;
        RECT 13.792 17.856 13.824 20.364 ;
  LAYER M1 ;
        RECT 13.728 17.856 13.76 20.364 ;
  LAYER M1 ;
        RECT 13.664 17.856 13.696 20.364 ;
  LAYER M1 ;
        RECT 13.6 17.856 13.632 20.364 ;
  LAYER M1 ;
        RECT 13.536 17.856 13.568 20.364 ;
  LAYER M1 ;
        RECT 13.472 17.856 13.504 20.364 ;
  LAYER M1 ;
        RECT 13.408 17.856 13.44 20.364 ;
  LAYER M1 ;
        RECT 13.344 17.856 13.376 20.364 ;
  LAYER M1 ;
        RECT 13.28 17.856 13.312 20.364 ;
  LAYER M1 ;
        RECT 13.216 17.856 13.248 20.364 ;
  LAYER M1 ;
        RECT 13.152 17.856 13.184 20.364 ;
  LAYER M1 ;
        RECT 13.088 17.856 13.12 20.364 ;
  LAYER M1 ;
        RECT 13.024 17.856 13.056 20.364 ;
  LAYER M1 ;
        RECT 12.96 17.856 12.992 20.364 ;
  LAYER M1 ;
        RECT 12.896 17.856 12.928 20.364 ;
  LAYER M1 ;
        RECT 12.832 17.856 12.864 20.364 ;
  LAYER M1 ;
        RECT 12.768 17.856 12.8 20.364 ;
  LAYER M1 ;
        RECT 12.704 17.856 12.736 20.364 ;
  LAYER M1 ;
        RECT 12.64 17.856 12.672 20.364 ;
  LAYER M2 ;
        RECT 12.524 17.94 14.996 17.972 ;
  LAYER M2 ;
        RECT 12.524 18.004 14.996 18.036 ;
  LAYER M2 ;
        RECT 12.524 18.068 14.996 18.1 ;
  LAYER M2 ;
        RECT 12.524 18.132 14.996 18.164 ;
  LAYER M2 ;
        RECT 12.524 18.196 14.996 18.228 ;
  LAYER M2 ;
        RECT 12.524 18.26 14.996 18.292 ;
  LAYER M2 ;
        RECT 12.524 18.324 14.996 18.356 ;
  LAYER M2 ;
        RECT 12.524 18.388 14.996 18.42 ;
  LAYER M2 ;
        RECT 12.524 18.452 14.996 18.484 ;
  LAYER M2 ;
        RECT 12.524 18.516 14.996 18.548 ;
  LAYER M2 ;
        RECT 12.524 18.58 14.996 18.612 ;
  LAYER M2 ;
        RECT 12.524 18.644 14.996 18.676 ;
  LAYER M2 ;
        RECT 12.524 18.708 14.996 18.74 ;
  LAYER M2 ;
        RECT 12.524 18.772 14.996 18.804 ;
  LAYER M2 ;
        RECT 12.524 18.836 14.996 18.868 ;
  LAYER M2 ;
        RECT 12.524 18.9 14.996 18.932 ;
  LAYER M2 ;
        RECT 12.524 18.964 14.996 18.996 ;
  LAYER M2 ;
        RECT 12.524 19.028 14.996 19.06 ;
  LAYER M2 ;
        RECT 12.524 19.092 14.996 19.124 ;
  LAYER M2 ;
        RECT 12.524 19.156 14.996 19.188 ;
  LAYER M2 ;
        RECT 12.524 19.22 14.996 19.252 ;
  LAYER M2 ;
        RECT 12.524 19.284 14.996 19.316 ;
  LAYER M2 ;
        RECT 12.524 19.348 14.996 19.38 ;
  LAYER M2 ;
        RECT 12.524 19.412 14.996 19.444 ;
  LAYER M2 ;
        RECT 12.524 19.476 14.996 19.508 ;
  LAYER M2 ;
        RECT 12.524 19.54 14.996 19.572 ;
  LAYER M2 ;
        RECT 12.524 19.604 14.996 19.636 ;
  LAYER M2 ;
        RECT 12.524 19.668 14.996 19.7 ;
  LAYER M2 ;
        RECT 12.524 19.732 14.996 19.764 ;
  LAYER M2 ;
        RECT 12.524 19.796 14.996 19.828 ;
  LAYER M2 ;
        RECT 12.524 19.86 14.996 19.892 ;
  LAYER M2 ;
        RECT 12.524 19.924 14.996 19.956 ;
  LAYER M2 ;
        RECT 12.524 19.988 14.996 20.02 ;
  LAYER M2 ;
        RECT 12.524 20.052 14.996 20.084 ;
  LAYER M2 ;
        RECT 12.524 20.116 14.996 20.148 ;
  LAYER M2 ;
        RECT 12.524 20.18 14.996 20.212 ;
  LAYER M3 ;
        RECT 14.944 17.856 14.976 20.364 ;
  LAYER M3 ;
        RECT 14.88 17.856 14.912 20.364 ;
  LAYER M3 ;
        RECT 14.816 17.856 14.848 20.364 ;
  LAYER M3 ;
        RECT 14.752 17.856 14.784 20.364 ;
  LAYER M3 ;
        RECT 14.688 17.856 14.72 20.364 ;
  LAYER M3 ;
        RECT 14.624 17.856 14.656 20.364 ;
  LAYER M3 ;
        RECT 14.56 17.856 14.592 20.364 ;
  LAYER M3 ;
        RECT 14.496 17.856 14.528 20.364 ;
  LAYER M3 ;
        RECT 14.432 17.856 14.464 20.364 ;
  LAYER M3 ;
        RECT 14.368 17.856 14.4 20.364 ;
  LAYER M3 ;
        RECT 14.304 17.856 14.336 20.364 ;
  LAYER M3 ;
        RECT 14.24 17.856 14.272 20.364 ;
  LAYER M3 ;
        RECT 14.176 17.856 14.208 20.364 ;
  LAYER M3 ;
        RECT 14.112 17.856 14.144 20.364 ;
  LAYER M3 ;
        RECT 14.048 17.856 14.08 20.364 ;
  LAYER M3 ;
        RECT 13.984 17.856 14.016 20.364 ;
  LAYER M3 ;
        RECT 13.92 17.856 13.952 20.364 ;
  LAYER M3 ;
        RECT 13.856 17.856 13.888 20.364 ;
  LAYER M3 ;
        RECT 13.792 17.856 13.824 20.364 ;
  LAYER M3 ;
        RECT 13.728 17.856 13.76 20.364 ;
  LAYER M3 ;
        RECT 13.664 17.856 13.696 20.364 ;
  LAYER M3 ;
        RECT 13.6 17.856 13.632 20.364 ;
  LAYER M3 ;
        RECT 13.536 17.856 13.568 20.364 ;
  LAYER M3 ;
        RECT 13.472 17.856 13.504 20.364 ;
  LAYER M3 ;
        RECT 13.408 17.856 13.44 20.364 ;
  LAYER M3 ;
        RECT 13.344 17.856 13.376 20.364 ;
  LAYER M3 ;
        RECT 13.28 17.856 13.312 20.364 ;
  LAYER M3 ;
        RECT 13.216 17.856 13.248 20.364 ;
  LAYER M3 ;
        RECT 13.152 17.856 13.184 20.364 ;
  LAYER M3 ;
        RECT 13.088 17.856 13.12 20.364 ;
  LAYER M3 ;
        RECT 13.024 17.856 13.056 20.364 ;
  LAYER M3 ;
        RECT 12.96 17.856 12.992 20.364 ;
  LAYER M3 ;
        RECT 12.896 17.856 12.928 20.364 ;
  LAYER M3 ;
        RECT 12.832 17.856 12.864 20.364 ;
  LAYER M3 ;
        RECT 12.768 17.856 12.8 20.364 ;
  LAYER M3 ;
        RECT 12.704 17.856 12.736 20.364 ;
  LAYER M3 ;
        RECT 12.64 17.856 12.672 20.364 ;
  LAYER M3 ;
        RECT 12.544 17.856 12.576 20.364 ;
  LAYER M1 ;
        RECT 14.959 17.892 14.961 20.328 ;
  LAYER M1 ;
        RECT 14.879 17.892 14.881 20.328 ;
  LAYER M1 ;
        RECT 14.799 17.892 14.801 20.328 ;
  LAYER M1 ;
        RECT 14.719 17.892 14.721 20.328 ;
  LAYER M1 ;
        RECT 14.639 17.892 14.641 20.328 ;
  LAYER M1 ;
        RECT 14.559 17.892 14.561 20.328 ;
  LAYER M1 ;
        RECT 14.479 17.892 14.481 20.328 ;
  LAYER M1 ;
        RECT 14.399 17.892 14.401 20.328 ;
  LAYER M1 ;
        RECT 14.319 17.892 14.321 20.328 ;
  LAYER M1 ;
        RECT 14.239 17.892 14.241 20.328 ;
  LAYER M1 ;
        RECT 14.159 17.892 14.161 20.328 ;
  LAYER M1 ;
        RECT 14.079 17.892 14.081 20.328 ;
  LAYER M1 ;
        RECT 13.999 17.892 14.001 20.328 ;
  LAYER M1 ;
        RECT 13.919 17.892 13.921 20.328 ;
  LAYER M1 ;
        RECT 13.839 17.892 13.841 20.328 ;
  LAYER M1 ;
        RECT 13.759 17.892 13.761 20.328 ;
  LAYER M1 ;
        RECT 13.679 17.892 13.681 20.328 ;
  LAYER M1 ;
        RECT 13.599 17.892 13.601 20.328 ;
  LAYER M1 ;
        RECT 13.519 17.892 13.521 20.328 ;
  LAYER M1 ;
        RECT 13.439 17.892 13.441 20.328 ;
  LAYER M1 ;
        RECT 13.359 17.892 13.361 20.328 ;
  LAYER M1 ;
        RECT 13.279 17.892 13.281 20.328 ;
  LAYER M1 ;
        RECT 13.199 17.892 13.201 20.328 ;
  LAYER M1 ;
        RECT 13.119 17.892 13.121 20.328 ;
  LAYER M1 ;
        RECT 13.039 17.892 13.041 20.328 ;
  LAYER M1 ;
        RECT 12.959 17.892 12.961 20.328 ;
  LAYER M1 ;
        RECT 12.879 17.892 12.881 20.328 ;
  LAYER M1 ;
        RECT 12.799 17.892 12.801 20.328 ;
  LAYER M1 ;
        RECT 12.719 17.892 12.721 20.328 ;
  LAYER M1 ;
        RECT 12.639 17.892 12.641 20.328 ;
  LAYER M2 ;
        RECT 12.56 17.891 14.96 17.893 ;
  LAYER M2 ;
        RECT 12.56 17.975 14.96 17.977 ;
  LAYER M2 ;
        RECT 12.56 18.059 14.96 18.061 ;
  LAYER M2 ;
        RECT 12.56 18.143 14.96 18.145 ;
  LAYER M2 ;
        RECT 12.56 18.227 14.96 18.229 ;
  LAYER M2 ;
        RECT 12.56 18.311 14.96 18.313 ;
  LAYER M2 ;
        RECT 12.56 18.395 14.96 18.397 ;
  LAYER M2 ;
        RECT 12.56 18.479 14.96 18.481 ;
  LAYER M2 ;
        RECT 12.56 18.563 14.96 18.565 ;
  LAYER M2 ;
        RECT 12.56 18.647 14.96 18.649 ;
  LAYER M2 ;
        RECT 12.56 18.731 14.96 18.733 ;
  LAYER M2 ;
        RECT 12.56 18.815 14.96 18.817 ;
  LAYER M2 ;
        RECT 12.56 18.8985 14.96 18.9005 ;
  LAYER M2 ;
        RECT 12.56 18.983 14.96 18.985 ;
  LAYER M2 ;
        RECT 12.56 19.067 14.96 19.069 ;
  LAYER M2 ;
        RECT 12.56 19.151 14.96 19.153 ;
  LAYER M2 ;
        RECT 12.56 19.235 14.96 19.237 ;
  LAYER M2 ;
        RECT 12.56 19.319 14.96 19.321 ;
  LAYER M2 ;
        RECT 12.56 19.403 14.96 19.405 ;
  LAYER M2 ;
        RECT 12.56 19.487 14.96 19.489 ;
  LAYER M2 ;
        RECT 12.56 19.571 14.96 19.573 ;
  LAYER M2 ;
        RECT 12.56 19.655 14.96 19.657 ;
  LAYER M2 ;
        RECT 12.56 19.739 14.96 19.741 ;
  LAYER M2 ;
        RECT 12.56 19.823 14.96 19.825 ;
  LAYER M2 ;
        RECT 12.56 19.907 14.96 19.909 ;
  LAYER M2 ;
        RECT 12.56 19.991 14.96 19.993 ;
  LAYER M2 ;
        RECT 12.56 20.075 14.96 20.077 ;
  LAYER M2 ;
        RECT 12.56 20.159 14.96 20.161 ;
  LAYER M2 ;
        RECT 12.56 20.243 14.96 20.245 ;
  LAYER M1 ;
        RECT 14.944 20.796 14.976 23.304 ;
  LAYER M1 ;
        RECT 14.88 20.796 14.912 23.304 ;
  LAYER M1 ;
        RECT 14.816 20.796 14.848 23.304 ;
  LAYER M1 ;
        RECT 14.752 20.796 14.784 23.304 ;
  LAYER M1 ;
        RECT 14.688 20.796 14.72 23.304 ;
  LAYER M1 ;
        RECT 14.624 20.796 14.656 23.304 ;
  LAYER M1 ;
        RECT 14.56 20.796 14.592 23.304 ;
  LAYER M1 ;
        RECT 14.496 20.796 14.528 23.304 ;
  LAYER M1 ;
        RECT 14.432 20.796 14.464 23.304 ;
  LAYER M1 ;
        RECT 14.368 20.796 14.4 23.304 ;
  LAYER M1 ;
        RECT 14.304 20.796 14.336 23.304 ;
  LAYER M1 ;
        RECT 14.24 20.796 14.272 23.304 ;
  LAYER M1 ;
        RECT 14.176 20.796 14.208 23.304 ;
  LAYER M1 ;
        RECT 14.112 20.796 14.144 23.304 ;
  LAYER M1 ;
        RECT 14.048 20.796 14.08 23.304 ;
  LAYER M1 ;
        RECT 13.984 20.796 14.016 23.304 ;
  LAYER M1 ;
        RECT 13.92 20.796 13.952 23.304 ;
  LAYER M1 ;
        RECT 13.856 20.796 13.888 23.304 ;
  LAYER M1 ;
        RECT 13.792 20.796 13.824 23.304 ;
  LAYER M1 ;
        RECT 13.728 20.796 13.76 23.304 ;
  LAYER M1 ;
        RECT 13.664 20.796 13.696 23.304 ;
  LAYER M1 ;
        RECT 13.6 20.796 13.632 23.304 ;
  LAYER M1 ;
        RECT 13.536 20.796 13.568 23.304 ;
  LAYER M1 ;
        RECT 13.472 20.796 13.504 23.304 ;
  LAYER M1 ;
        RECT 13.408 20.796 13.44 23.304 ;
  LAYER M1 ;
        RECT 13.344 20.796 13.376 23.304 ;
  LAYER M1 ;
        RECT 13.28 20.796 13.312 23.304 ;
  LAYER M1 ;
        RECT 13.216 20.796 13.248 23.304 ;
  LAYER M1 ;
        RECT 13.152 20.796 13.184 23.304 ;
  LAYER M1 ;
        RECT 13.088 20.796 13.12 23.304 ;
  LAYER M1 ;
        RECT 13.024 20.796 13.056 23.304 ;
  LAYER M1 ;
        RECT 12.96 20.796 12.992 23.304 ;
  LAYER M1 ;
        RECT 12.896 20.796 12.928 23.304 ;
  LAYER M1 ;
        RECT 12.832 20.796 12.864 23.304 ;
  LAYER M1 ;
        RECT 12.768 20.796 12.8 23.304 ;
  LAYER M1 ;
        RECT 12.704 20.796 12.736 23.304 ;
  LAYER M1 ;
        RECT 12.64 20.796 12.672 23.304 ;
  LAYER M2 ;
        RECT 12.524 20.88 14.996 20.912 ;
  LAYER M2 ;
        RECT 12.524 20.944 14.996 20.976 ;
  LAYER M2 ;
        RECT 12.524 21.008 14.996 21.04 ;
  LAYER M2 ;
        RECT 12.524 21.072 14.996 21.104 ;
  LAYER M2 ;
        RECT 12.524 21.136 14.996 21.168 ;
  LAYER M2 ;
        RECT 12.524 21.2 14.996 21.232 ;
  LAYER M2 ;
        RECT 12.524 21.264 14.996 21.296 ;
  LAYER M2 ;
        RECT 12.524 21.328 14.996 21.36 ;
  LAYER M2 ;
        RECT 12.524 21.392 14.996 21.424 ;
  LAYER M2 ;
        RECT 12.524 21.456 14.996 21.488 ;
  LAYER M2 ;
        RECT 12.524 21.52 14.996 21.552 ;
  LAYER M2 ;
        RECT 12.524 21.584 14.996 21.616 ;
  LAYER M2 ;
        RECT 12.524 21.648 14.996 21.68 ;
  LAYER M2 ;
        RECT 12.524 21.712 14.996 21.744 ;
  LAYER M2 ;
        RECT 12.524 21.776 14.996 21.808 ;
  LAYER M2 ;
        RECT 12.524 21.84 14.996 21.872 ;
  LAYER M2 ;
        RECT 12.524 21.904 14.996 21.936 ;
  LAYER M2 ;
        RECT 12.524 21.968 14.996 22 ;
  LAYER M2 ;
        RECT 12.524 22.032 14.996 22.064 ;
  LAYER M2 ;
        RECT 12.524 22.096 14.996 22.128 ;
  LAYER M2 ;
        RECT 12.524 22.16 14.996 22.192 ;
  LAYER M2 ;
        RECT 12.524 22.224 14.996 22.256 ;
  LAYER M2 ;
        RECT 12.524 22.288 14.996 22.32 ;
  LAYER M2 ;
        RECT 12.524 22.352 14.996 22.384 ;
  LAYER M2 ;
        RECT 12.524 22.416 14.996 22.448 ;
  LAYER M2 ;
        RECT 12.524 22.48 14.996 22.512 ;
  LAYER M2 ;
        RECT 12.524 22.544 14.996 22.576 ;
  LAYER M2 ;
        RECT 12.524 22.608 14.996 22.64 ;
  LAYER M2 ;
        RECT 12.524 22.672 14.996 22.704 ;
  LAYER M2 ;
        RECT 12.524 22.736 14.996 22.768 ;
  LAYER M2 ;
        RECT 12.524 22.8 14.996 22.832 ;
  LAYER M2 ;
        RECT 12.524 22.864 14.996 22.896 ;
  LAYER M2 ;
        RECT 12.524 22.928 14.996 22.96 ;
  LAYER M2 ;
        RECT 12.524 22.992 14.996 23.024 ;
  LAYER M2 ;
        RECT 12.524 23.056 14.996 23.088 ;
  LAYER M2 ;
        RECT 12.524 23.12 14.996 23.152 ;
  LAYER M3 ;
        RECT 14.944 20.796 14.976 23.304 ;
  LAYER M3 ;
        RECT 14.88 20.796 14.912 23.304 ;
  LAYER M3 ;
        RECT 14.816 20.796 14.848 23.304 ;
  LAYER M3 ;
        RECT 14.752 20.796 14.784 23.304 ;
  LAYER M3 ;
        RECT 14.688 20.796 14.72 23.304 ;
  LAYER M3 ;
        RECT 14.624 20.796 14.656 23.304 ;
  LAYER M3 ;
        RECT 14.56 20.796 14.592 23.304 ;
  LAYER M3 ;
        RECT 14.496 20.796 14.528 23.304 ;
  LAYER M3 ;
        RECT 14.432 20.796 14.464 23.304 ;
  LAYER M3 ;
        RECT 14.368 20.796 14.4 23.304 ;
  LAYER M3 ;
        RECT 14.304 20.796 14.336 23.304 ;
  LAYER M3 ;
        RECT 14.24 20.796 14.272 23.304 ;
  LAYER M3 ;
        RECT 14.176 20.796 14.208 23.304 ;
  LAYER M3 ;
        RECT 14.112 20.796 14.144 23.304 ;
  LAYER M3 ;
        RECT 14.048 20.796 14.08 23.304 ;
  LAYER M3 ;
        RECT 13.984 20.796 14.016 23.304 ;
  LAYER M3 ;
        RECT 13.92 20.796 13.952 23.304 ;
  LAYER M3 ;
        RECT 13.856 20.796 13.888 23.304 ;
  LAYER M3 ;
        RECT 13.792 20.796 13.824 23.304 ;
  LAYER M3 ;
        RECT 13.728 20.796 13.76 23.304 ;
  LAYER M3 ;
        RECT 13.664 20.796 13.696 23.304 ;
  LAYER M3 ;
        RECT 13.6 20.796 13.632 23.304 ;
  LAYER M3 ;
        RECT 13.536 20.796 13.568 23.304 ;
  LAYER M3 ;
        RECT 13.472 20.796 13.504 23.304 ;
  LAYER M3 ;
        RECT 13.408 20.796 13.44 23.304 ;
  LAYER M3 ;
        RECT 13.344 20.796 13.376 23.304 ;
  LAYER M3 ;
        RECT 13.28 20.796 13.312 23.304 ;
  LAYER M3 ;
        RECT 13.216 20.796 13.248 23.304 ;
  LAYER M3 ;
        RECT 13.152 20.796 13.184 23.304 ;
  LAYER M3 ;
        RECT 13.088 20.796 13.12 23.304 ;
  LAYER M3 ;
        RECT 13.024 20.796 13.056 23.304 ;
  LAYER M3 ;
        RECT 12.96 20.796 12.992 23.304 ;
  LAYER M3 ;
        RECT 12.896 20.796 12.928 23.304 ;
  LAYER M3 ;
        RECT 12.832 20.796 12.864 23.304 ;
  LAYER M3 ;
        RECT 12.768 20.796 12.8 23.304 ;
  LAYER M3 ;
        RECT 12.704 20.796 12.736 23.304 ;
  LAYER M3 ;
        RECT 12.64 20.796 12.672 23.304 ;
  LAYER M3 ;
        RECT 12.544 20.796 12.576 23.304 ;
  LAYER M1 ;
        RECT 14.959 20.832 14.961 23.268 ;
  LAYER M1 ;
        RECT 14.879 20.832 14.881 23.268 ;
  LAYER M1 ;
        RECT 14.799 20.832 14.801 23.268 ;
  LAYER M1 ;
        RECT 14.719 20.832 14.721 23.268 ;
  LAYER M1 ;
        RECT 14.639 20.832 14.641 23.268 ;
  LAYER M1 ;
        RECT 14.559 20.832 14.561 23.268 ;
  LAYER M1 ;
        RECT 14.479 20.832 14.481 23.268 ;
  LAYER M1 ;
        RECT 14.399 20.832 14.401 23.268 ;
  LAYER M1 ;
        RECT 14.319 20.832 14.321 23.268 ;
  LAYER M1 ;
        RECT 14.239 20.832 14.241 23.268 ;
  LAYER M1 ;
        RECT 14.159 20.832 14.161 23.268 ;
  LAYER M1 ;
        RECT 14.079 20.832 14.081 23.268 ;
  LAYER M1 ;
        RECT 13.999 20.832 14.001 23.268 ;
  LAYER M1 ;
        RECT 13.919 20.832 13.921 23.268 ;
  LAYER M1 ;
        RECT 13.839 20.832 13.841 23.268 ;
  LAYER M1 ;
        RECT 13.759 20.832 13.761 23.268 ;
  LAYER M1 ;
        RECT 13.679 20.832 13.681 23.268 ;
  LAYER M1 ;
        RECT 13.599 20.832 13.601 23.268 ;
  LAYER M1 ;
        RECT 13.519 20.832 13.521 23.268 ;
  LAYER M1 ;
        RECT 13.439 20.832 13.441 23.268 ;
  LAYER M1 ;
        RECT 13.359 20.832 13.361 23.268 ;
  LAYER M1 ;
        RECT 13.279 20.832 13.281 23.268 ;
  LAYER M1 ;
        RECT 13.199 20.832 13.201 23.268 ;
  LAYER M1 ;
        RECT 13.119 20.832 13.121 23.268 ;
  LAYER M1 ;
        RECT 13.039 20.832 13.041 23.268 ;
  LAYER M1 ;
        RECT 12.959 20.832 12.961 23.268 ;
  LAYER M1 ;
        RECT 12.879 20.832 12.881 23.268 ;
  LAYER M1 ;
        RECT 12.799 20.832 12.801 23.268 ;
  LAYER M1 ;
        RECT 12.719 20.832 12.721 23.268 ;
  LAYER M1 ;
        RECT 12.639 20.832 12.641 23.268 ;
  LAYER M2 ;
        RECT 12.56 20.831 14.96 20.833 ;
  LAYER M2 ;
        RECT 12.56 20.915 14.96 20.917 ;
  LAYER M2 ;
        RECT 12.56 20.999 14.96 21.001 ;
  LAYER M2 ;
        RECT 12.56 21.083 14.96 21.085 ;
  LAYER M2 ;
        RECT 12.56 21.167 14.96 21.169 ;
  LAYER M2 ;
        RECT 12.56 21.251 14.96 21.253 ;
  LAYER M2 ;
        RECT 12.56 21.335 14.96 21.337 ;
  LAYER M2 ;
        RECT 12.56 21.419 14.96 21.421 ;
  LAYER M2 ;
        RECT 12.56 21.503 14.96 21.505 ;
  LAYER M2 ;
        RECT 12.56 21.587 14.96 21.589 ;
  LAYER M2 ;
        RECT 12.56 21.671 14.96 21.673 ;
  LAYER M2 ;
        RECT 12.56 21.755 14.96 21.757 ;
  LAYER M2 ;
        RECT 12.56 21.8385 14.96 21.8405 ;
  LAYER M2 ;
        RECT 12.56 21.923 14.96 21.925 ;
  LAYER M2 ;
        RECT 12.56 22.007 14.96 22.009 ;
  LAYER M2 ;
        RECT 12.56 22.091 14.96 22.093 ;
  LAYER M2 ;
        RECT 12.56 22.175 14.96 22.177 ;
  LAYER M2 ;
        RECT 12.56 22.259 14.96 22.261 ;
  LAYER M2 ;
        RECT 12.56 22.343 14.96 22.345 ;
  LAYER M2 ;
        RECT 12.56 22.427 14.96 22.429 ;
  LAYER M2 ;
        RECT 12.56 22.511 14.96 22.513 ;
  LAYER M2 ;
        RECT 12.56 22.595 14.96 22.597 ;
  LAYER M2 ;
        RECT 12.56 22.679 14.96 22.681 ;
  LAYER M2 ;
        RECT 12.56 22.763 14.96 22.765 ;
  LAYER M2 ;
        RECT 12.56 22.847 14.96 22.849 ;
  LAYER M2 ;
        RECT 12.56 22.931 14.96 22.933 ;
  LAYER M2 ;
        RECT 12.56 23.015 14.96 23.017 ;
  LAYER M2 ;
        RECT 12.56 23.099 14.96 23.101 ;
  LAYER M2 ;
        RECT 12.56 23.183 14.96 23.185 ;
  LAYER M1 ;
        RECT 14.944 23.736 14.976 26.244 ;
  LAYER M1 ;
        RECT 14.88 23.736 14.912 26.244 ;
  LAYER M1 ;
        RECT 14.816 23.736 14.848 26.244 ;
  LAYER M1 ;
        RECT 14.752 23.736 14.784 26.244 ;
  LAYER M1 ;
        RECT 14.688 23.736 14.72 26.244 ;
  LAYER M1 ;
        RECT 14.624 23.736 14.656 26.244 ;
  LAYER M1 ;
        RECT 14.56 23.736 14.592 26.244 ;
  LAYER M1 ;
        RECT 14.496 23.736 14.528 26.244 ;
  LAYER M1 ;
        RECT 14.432 23.736 14.464 26.244 ;
  LAYER M1 ;
        RECT 14.368 23.736 14.4 26.244 ;
  LAYER M1 ;
        RECT 14.304 23.736 14.336 26.244 ;
  LAYER M1 ;
        RECT 14.24 23.736 14.272 26.244 ;
  LAYER M1 ;
        RECT 14.176 23.736 14.208 26.244 ;
  LAYER M1 ;
        RECT 14.112 23.736 14.144 26.244 ;
  LAYER M1 ;
        RECT 14.048 23.736 14.08 26.244 ;
  LAYER M1 ;
        RECT 13.984 23.736 14.016 26.244 ;
  LAYER M1 ;
        RECT 13.92 23.736 13.952 26.244 ;
  LAYER M1 ;
        RECT 13.856 23.736 13.888 26.244 ;
  LAYER M1 ;
        RECT 13.792 23.736 13.824 26.244 ;
  LAYER M1 ;
        RECT 13.728 23.736 13.76 26.244 ;
  LAYER M1 ;
        RECT 13.664 23.736 13.696 26.244 ;
  LAYER M1 ;
        RECT 13.6 23.736 13.632 26.244 ;
  LAYER M1 ;
        RECT 13.536 23.736 13.568 26.244 ;
  LAYER M1 ;
        RECT 13.472 23.736 13.504 26.244 ;
  LAYER M1 ;
        RECT 13.408 23.736 13.44 26.244 ;
  LAYER M1 ;
        RECT 13.344 23.736 13.376 26.244 ;
  LAYER M1 ;
        RECT 13.28 23.736 13.312 26.244 ;
  LAYER M1 ;
        RECT 13.216 23.736 13.248 26.244 ;
  LAYER M1 ;
        RECT 13.152 23.736 13.184 26.244 ;
  LAYER M1 ;
        RECT 13.088 23.736 13.12 26.244 ;
  LAYER M1 ;
        RECT 13.024 23.736 13.056 26.244 ;
  LAYER M1 ;
        RECT 12.96 23.736 12.992 26.244 ;
  LAYER M1 ;
        RECT 12.896 23.736 12.928 26.244 ;
  LAYER M1 ;
        RECT 12.832 23.736 12.864 26.244 ;
  LAYER M1 ;
        RECT 12.768 23.736 12.8 26.244 ;
  LAYER M1 ;
        RECT 12.704 23.736 12.736 26.244 ;
  LAYER M1 ;
        RECT 12.64 23.736 12.672 26.244 ;
  LAYER M2 ;
        RECT 12.524 23.82 14.996 23.852 ;
  LAYER M2 ;
        RECT 12.524 23.884 14.996 23.916 ;
  LAYER M2 ;
        RECT 12.524 23.948 14.996 23.98 ;
  LAYER M2 ;
        RECT 12.524 24.012 14.996 24.044 ;
  LAYER M2 ;
        RECT 12.524 24.076 14.996 24.108 ;
  LAYER M2 ;
        RECT 12.524 24.14 14.996 24.172 ;
  LAYER M2 ;
        RECT 12.524 24.204 14.996 24.236 ;
  LAYER M2 ;
        RECT 12.524 24.268 14.996 24.3 ;
  LAYER M2 ;
        RECT 12.524 24.332 14.996 24.364 ;
  LAYER M2 ;
        RECT 12.524 24.396 14.996 24.428 ;
  LAYER M2 ;
        RECT 12.524 24.46 14.996 24.492 ;
  LAYER M2 ;
        RECT 12.524 24.524 14.996 24.556 ;
  LAYER M2 ;
        RECT 12.524 24.588 14.996 24.62 ;
  LAYER M2 ;
        RECT 12.524 24.652 14.996 24.684 ;
  LAYER M2 ;
        RECT 12.524 24.716 14.996 24.748 ;
  LAYER M2 ;
        RECT 12.524 24.78 14.996 24.812 ;
  LAYER M2 ;
        RECT 12.524 24.844 14.996 24.876 ;
  LAYER M2 ;
        RECT 12.524 24.908 14.996 24.94 ;
  LAYER M2 ;
        RECT 12.524 24.972 14.996 25.004 ;
  LAYER M2 ;
        RECT 12.524 25.036 14.996 25.068 ;
  LAYER M2 ;
        RECT 12.524 25.1 14.996 25.132 ;
  LAYER M2 ;
        RECT 12.524 25.164 14.996 25.196 ;
  LAYER M2 ;
        RECT 12.524 25.228 14.996 25.26 ;
  LAYER M2 ;
        RECT 12.524 25.292 14.996 25.324 ;
  LAYER M2 ;
        RECT 12.524 25.356 14.996 25.388 ;
  LAYER M2 ;
        RECT 12.524 25.42 14.996 25.452 ;
  LAYER M2 ;
        RECT 12.524 25.484 14.996 25.516 ;
  LAYER M2 ;
        RECT 12.524 25.548 14.996 25.58 ;
  LAYER M2 ;
        RECT 12.524 25.612 14.996 25.644 ;
  LAYER M2 ;
        RECT 12.524 25.676 14.996 25.708 ;
  LAYER M2 ;
        RECT 12.524 25.74 14.996 25.772 ;
  LAYER M2 ;
        RECT 12.524 25.804 14.996 25.836 ;
  LAYER M2 ;
        RECT 12.524 25.868 14.996 25.9 ;
  LAYER M2 ;
        RECT 12.524 25.932 14.996 25.964 ;
  LAYER M2 ;
        RECT 12.524 25.996 14.996 26.028 ;
  LAYER M2 ;
        RECT 12.524 26.06 14.996 26.092 ;
  LAYER M3 ;
        RECT 14.944 23.736 14.976 26.244 ;
  LAYER M3 ;
        RECT 14.88 23.736 14.912 26.244 ;
  LAYER M3 ;
        RECT 14.816 23.736 14.848 26.244 ;
  LAYER M3 ;
        RECT 14.752 23.736 14.784 26.244 ;
  LAYER M3 ;
        RECT 14.688 23.736 14.72 26.244 ;
  LAYER M3 ;
        RECT 14.624 23.736 14.656 26.244 ;
  LAYER M3 ;
        RECT 14.56 23.736 14.592 26.244 ;
  LAYER M3 ;
        RECT 14.496 23.736 14.528 26.244 ;
  LAYER M3 ;
        RECT 14.432 23.736 14.464 26.244 ;
  LAYER M3 ;
        RECT 14.368 23.736 14.4 26.244 ;
  LAYER M3 ;
        RECT 14.304 23.736 14.336 26.244 ;
  LAYER M3 ;
        RECT 14.24 23.736 14.272 26.244 ;
  LAYER M3 ;
        RECT 14.176 23.736 14.208 26.244 ;
  LAYER M3 ;
        RECT 14.112 23.736 14.144 26.244 ;
  LAYER M3 ;
        RECT 14.048 23.736 14.08 26.244 ;
  LAYER M3 ;
        RECT 13.984 23.736 14.016 26.244 ;
  LAYER M3 ;
        RECT 13.92 23.736 13.952 26.244 ;
  LAYER M3 ;
        RECT 13.856 23.736 13.888 26.244 ;
  LAYER M3 ;
        RECT 13.792 23.736 13.824 26.244 ;
  LAYER M3 ;
        RECT 13.728 23.736 13.76 26.244 ;
  LAYER M3 ;
        RECT 13.664 23.736 13.696 26.244 ;
  LAYER M3 ;
        RECT 13.6 23.736 13.632 26.244 ;
  LAYER M3 ;
        RECT 13.536 23.736 13.568 26.244 ;
  LAYER M3 ;
        RECT 13.472 23.736 13.504 26.244 ;
  LAYER M3 ;
        RECT 13.408 23.736 13.44 26.244 ;
  LAYER M3 ;
        RECT 13.344 23.736 13.376 26.244 ;
  LAYER M3 ;
        RECT 13.28 23.736 13.312 26.244 ;
  LAYER M3 ;
        RECT 13.216 23.736 13.248 26.244 ;
  LAYER M3 ;
        RECT 13.152 23.736 13.184 26.244 ;
  LAYER M3 ;
        RECT 13.088 23.736 13.12 26.244 ;
  LAYER M3 ;
        RECT 13.024 23.736 13.056 26.244 ;
  LAYER M3 ;
        RECT 12.96 23.736 12.992 26.244 ;
  LAYER M3 ;
        RECT 12.896 23.736 12.928 26.244 ;
  LAYER M3 ;
        RECT 12.832 23.736 12.864 26.244 ;
  LAYER M3 ;
        RECT 12.768 23.736 12.8 26.244 ;
  LAYER M3 ;
        RECT 12.704 23.736 12.736 26.244 ;
  LAYER M3 ;
        RECT 12.64 23.736 12.672 26.244 ;
  LAYER M3 ;
        RECT 12.544 23.736 12.576 26.244 ;
  LAYER M1 ;
        RECT 14.959 23.772 14.961 26.208 ;
  LAYER M1 ;
        RECT 14.879 23.772 14.881 26.208 ;
  LAYER M1 ;
        RECT 14.799 23.772 14.801 26.208 ;
  LAYER M1 ;
        RECT 14.719 23.772 14.721 26.208 ;
  LAYER M1 ;
        RECT 14.639 23.772 14.641 26.208 ;
  LAYER M1 ;
        RECT 14.559 23.772 14.561 26.208 ;
  LAYER M1 ;
        RECT 14.479 23.772 14.481 26.208 ;
  LAYER M1 ;
        RECT 14.399 23.772 14.401 26.208 ;
  LAYER M1 ;
        RECT 14.319 23.772 14.321 26.208 ;
  LAYER M1 ;
        RECT 14.239 23.772 14.241 26.208 ;
  LAYER M1 ;
        RECT 14.159 23.772 14.161 26.208 ;
  LAYER M1 ;
        RECT 14.079 23.772 14.081 26.208 ;
  LAYER M1 ;
        RECT 13.999 23.772 14.001 26.208 ;
  LAYER M1 ;
        RECT 13.919 23.772 13.921 26.208 ;
  LAYER M1 ;
        RECT 13.839 23.772 13.841 26.208 ;
  LAYER M1 ;
        RECT 13.759 23.772 13.761 26.208 ;
  LAYER M1 ;
        RECT 13.679 23.772 13.681 26.208 ;
  LAYER M1 ;
        RECT 13.599 23.772 13.601 26.208 ;
  LAYER M1 ;
        RECT 13.519 23.772 13.521 26.208 ;
  LAYER M1 ;
        RECT 13.439 23.772 13.441 26.208 ;
  LAYER M1 ;
        RECT 13.359 23.772 13.361 26.208 ;
  LAYER M1 ;
        RECT 13.279 23.772 13.281 26.208 ;
  LAYER M1 ;
        RECT 13.199 23.772 13.201 26.208 ;
  LAYER M1 ;
        RECT 13.119 23.772 13.121 26.208 ;
  LAYER M1 ;
        RECT 13.039 23.772 13.041 26.208 ;
  LAYER M1 ;
        RECT 12.959 23.772 12.961 26.208 ;
  LAYER M1 ;
        RECT 12.879 23.772 12.881 26.208 ;
  LAYER M1 ;
        RECT 12.799 23.772 12.801 26.208 ;
  LAYER M1 ;
        RECT 12.719 23.772 12.721 26.208 ;
  LAYER M1 ;
        RECT 12.639 23.772 12.641 26.208 ;
  LAYER M2 ;
        RECT 12.56 23.771 14.96 23.773 ;
  LAYER M2 ;
        RECT 12.56 23.855 14.96 23.857 ;
  LAYER M2 ;
        RECT 12.56 23.939 14.96 23.941 ;
  LAYER M2 ;
        RECT 12.56 24.023 14.96 24.025 ;
  LAYER M2 ;
        RECT 12.56 24.107 14.96 24.109 ;
  LAYER M2 ;
        RECT 12.56 24.191 14.96 24.193 ;
  LAYER M2 ;
        RECT 12.56 24.275 14.96 24.277 ;
  LAYER M2 ;
        RECT 12.56 24.359 14.96 24.361 ;
  LAYER M2 ;
        RECT 12.56 24.443 14.96 24.445 ;
  LAYER M2 ;
        RECT 12.56 24.527 14.96 24.529 ;
  LAYER M2 ;
        RECT 12.56 24.611 14.96 24.613 ;
  LAYER M2 ;
        RECT 12.56 24.695 14.96 24.697 ;
  LAYER M2 ;
        RECT 12.56 24.7785 14.96 24.7805 ;
  LAYER M2 ;
        RECT 12.56 24.863 14.96 24.865 ;
  LAYER M2 ;
        RECT 12.56 24.947 14.96 24.949 ;
  LAYER M2 ;
        RECT 12.56 25.031 14.96 25.033 ;
  LAYER M2 ;
        RECT 12.56 25.115 14.96 25.117 ;
  LAYER M2 ;
        RECT 12.56 25.199 14.96 25.201 ;
  LAYER M2 ;
        RECT 12.56 25.283 14.96 25.285 ;
  LAYER M2 ;
        RECT 12.56 25.367 14.96 25.369 ;
  LAYER M2 ;
        RECT 12.56 25.451 14.96 25.453 ;
  LAYER M2 ;
        RECT 12.56 25.535 14.96 25.537 ;
  LAYER M2 ;
        RECT 12.56 25.619 14.96 25.621 ;
  LAYER M2 ;
        RECT 12.56 25.703 14.96 25.705 ;
  LAYER M2 ;
        RECT 12.56 25.787 14.96 25.789 ;
  LAYER M2 ;
        RECT 12.56 25.871 14.96 25.873 ;
  LAYER M2 ;
        RECT 12.56 25.955 14.96 25.957 ;
  LAYER M2 ;
        RECT 12.56 26.039 14.96 26.041 ;
  LAYER M2 ;
        RECT 12.56 26.123 14.96 26.125 ;
  LAYER M1 ;
        RECT 14.944 26.676 14.976 29.184 ;
  LAYER M1 ;
        RECT 14.88 26.676 14.912 29.184 ;
  LAYER M1 ;
        RECT 14.816 26.676 14.848 29.184 ;
  LAYER M1 ;
        RECT 14.752 26.676 14.784 29.184 ;
  LAYER M1 ;
        RECT 14.688 26.676 14.72 29.184 ;
  LAYER M1 ;
        RECT 14.624 26.676 14.656 29.184 ;
  LAYER M1 ;
        RECT 14.56 26.676 14.592 29.184 ;
  LAYER M1 ;
        RECT 14.496 26.676 14.528 29.184 ;
  LAYER M1 ;
        RECT 14.432 26.676 14.464 29.184 ;
  LAYER M1 ;
        RECT 14.368 26.676 14.4 29.184 ;
  LAYER M1 ;
        RECT 14.304 26.676 14.336 29.184 ;
  LAYER M1 ;
        RECT 14.24 26.676 14.272 29.184 ;
  LAYER M1 ;
        RECT 14.176 26.676 14.208 29.184 ;
  LAYER M1 ;
        RECT 14.112 26.676 14.144 29.184 ;
  LAYER M1 ;
        RECT 14.048 26.676 14.08 29.184 ;
  LAYER M1 ;
        RECT 13.984 26.676 14.016 29.184 ;
  LAYER M1 ;
        RECT 13.92 26.676 13.952 29.184 ;
  LAYER M1 ;
        RECT 13.856 26.676 13.888 29.184 ;
  LAYER M1 ;
        RECT 13.792 26.676 13.824 29.184 ;
  LAYER M1 ;
        RECT 13.728 26.676 13.76 29.184 ;
  LAYER M1 ;
        RECT 13.664 26.676 13.696 29.184 ;
  LAYER M1 ;
        RECT 13.6 26.676 13.632 29.184 ;
  LAYER M1 ;
        RECT 13.536 26.676 13.568 29.184 ;
  LAYER M1 ;
        RECT 13.472 26.676 13.504 29.184 ;
  LAYER M1 ;
        RECT 13.408 26.676 13.44 29.184 ;
  LAYER M1 ;
        RECT 13.344 26.676 13.376 29.184 ;
  LAYER M1 ;
        RECT 13.28 26.676 13.312 29.184 ;
  LAYER M1 ;
        RECT 13.216 26.676 13.248 29.184 ;
  LAYER M1 ;
        RECT 13.152 26.676 13.184 29.184 ;
  LAYER M1 ;
        RECT 13.088 26.676 13.12 29.184 ;
  LAYER M1 ;
        RECT 13.024 26.676 13.056 29.184 ;
  LAYER M1 ;
        RECT 12.96 26.676 12.992 29.184 ;
  LAYER M1 ;
        RECT 12.896 26.676 12.928 29.184 ;
  LAYER M1 ;
        RECT 12.832 26.676 12.864 29.184 ;
  LAYER M1 ;
        RECT 12.768 26.676 12.8 29.184 ;
  LAYER M1 ;
        RECT 12.704 26.676 12.736 29.184 ;
  LAYER M1 ;
        RECT 12.64 26.676 12.672 29.184 ;
  LAYER M2 ;
        RECT 12.524 26.76 14.996 26.792 ;
  LAYER M2 ;
        RECT 12.524 26.824 14.996 26.856 ;
  LAYER M2 ;
        RECT 12.524 26.888 14.996 26.92 ;
  LAYER M2 ;
        RECT 12.524 26.952 14.996 26.984 ;
  LAYER M2 ;
        RECT 12.524 27.016 14.996 27.048 ;
  LAYER M2 ;
        RECT 12.524 27.08 14.996 27.112 ;
  LAYER M2 ;
        RECT 12.524 27.144 14.996 27.176 ;
  LAYER M2 ;
        RECT 12.524 27.208 14.996 27.24 ;
  LAYER M2 ;
        RECT 12.524 27.272 14.996 27.304 ;
  LAYER M2 ;
        RECT 12.524 27.336 14.996 27.368 ;
  LAYER M2 ;
        RECT 12.524 27.4 14.996 27.432 ;
  LAYER M2 ;
        RECT 12.524 27.464 14.996 27.496 ;
  LAYER M2 ;
        RECT 12.524 27.528 14.996 27.56 ;
  LAYER M2 ;
        RECT 12.524 27.592 14.996 27.624 ;
  LAYER M2 ;
        RECT 12.524 27.656 14.996 27.688 ;
  LAYER M2 ;
        RECT 12.524 27.72 14.996 27.752 ;
  LAYER M2 ;
        RECT 12.524 27.784 14.996 27.816 ;
  LAYER M2 ;
        RECT 12.524 27.848 14.996 27.88 ;
  LAYER M2 ;
        RECT 12.524 27.912 14.996 27.944 ;
  LAYER M2 ;
        RECT 12.524 27.976 14.996 28.008 ;
  LAYER M2 ;
        RECT 12.524 28.04 14.996 28.072 ;
  LAYER M2 ;
        RECT 12.524 28.104 14.996 28.136 ;
  LAYER M2 ;
        RECT 12.524 28.168 14.996 28.2 ;
  LAYER M2 ;
        RECT 12.524 28.232 14.996 28.264 ;
  LAYER M2 ;
        RECT 12.524 28.296 14.996 28.328 ;
  LAYER M2 ;
        RECT 12.524 28.36 14.996 28.392 ;
  LAYER M2 ;
        RECT 12.524 28.424 14.996 28.456 ;
  LAYER M2 ;
        RECT 12.524 28.488 14.996 28.52 ;
  LAYER M2 ;
        RECT 12.524 28.552 14.996 28.584 ;
  LAYER M2 ;
        RECT 12.524 28.616 14.996 28.648 ;
  LAYER M2 ;
        RECT 12.524 28.68 14.996 28.712 ;
  LAYER M2 ;
        RECT 12.524 28.744 14.996 28.776 ;
  LAYER M2 ;
        RECT 12.524 28.808 14.996 28.84 ;
  LAYER M2 ;
        RECT 12.524 28.872 14.996 28.904 ;
  LAYER M2 ;
        RECT 12.524 28.936 14.996 28.968 ;
  LAYER M2 ;
        RECT 12.524 29 14.996 29.032 ;
  LAYER M3 ;
        RECT 14.944 26.676 14.976 29.184 ;
  LAYER M3 ;
        RECT 14.88 26.676 14.912 29.184 ;
  LAYER M3 ;
        RECT 14.816 26.676 14.848 29.184 ;
  LAYER M3 ;
        RECT 14.752 26.676 14.784 29.184 ;
  LAYER M3 ;
        RECT 14.688 26.676 14.72 29.184 ;
  LAYER M3 ;
        RECT 14.624 26.676 14.656 29.184 ;
  LAYER M3 ;
        RECT 14.56 26.676 14.592 29.184 ;
  LAYER M3 ;
        RECT 14.496 26.676 14.528 29.184 ;
  LAYER M3 ;
        RECT 14.432 26.676 14.464 29.184 ;
  LAYER M3 ;
        RECT 14.368 26.676 14.4 29.184 ;
  LAYER M3 ;
        RECT 14.304 26.676 14.336 29.184 ;
  LAYER M3 ;
        RECT 14.24 26.676 14.272 29.184 ;
  LAYER M3 ;
        RECT 14.176 26.676 14.208 29.184 ;
  LAYER M3 ;
        RECT 14.112 26.676 14.144 29.184 ;
  LAYER M3 ;
        RECT 14.048 26.676 14.08 29.184 ;
  LAYER M3 ;
        RECT 13.984 26.676 14.016 29.184 ;
  LAYER M3 ;
        RECT 13.92 26.676 13.952 29.184 ;
  LAYER M3 ;
        RECT 13.856 26.676 13.888 29.184 ;
  LAYER M3 ;
        RECT 13.792 26.676 13.824 29.184 ;
  LAYER M3 ;
        RECT 13.728 26.676 13.76 29.184 ;
  LAYER M3 ;
        RECT 13.664 26.676 13.696 29.184 ;
  LAYER M3 ;
        RECT 13.6 26.676 13.632 29.184 ;
  LAYER M3 ;
        RECT 13.536 26.676 13.568 29.184 ;
  LAYER M3 ;
        RECT 13.472 26.676 13.504 29.184 ;
  LAYER M3 ;
        RECT 13.408 26.676 13.44 29.184 ;
  LAYER M3 ;
        RECT 13.344 26.676 13.376 29.184 ;
  LAYER M3 ;
        RECT 13.28 26.676 13.312 29.184 ;
  LAYER M3 ;
        RECT 13.216 26.676 13.248 29.184 ;
  LAYER M3 ;
        RECT 13.152 26.676 13.184 29.184 ;
  LAYER M3 ;
        RECT 13.088 26.676 13.12 29.184 ;
  LAYER M3 ;
        RECT 13.024 26.676 13.056 29.184 ;
  LAYER M3 ;
        RECT 12.96 26.676 12.992 29.184 ;
  LAYER M3 ;
        RECT 12.896 26.676 12.928 29.184 ;
  LAYER M3 ;
        RECT 12.832 26.676 12.864 29.184 ;
  LAYER M3 ;
        RECT 12.768 26.676 12.8 29.184 ;
  LAYER M3 ;
        RECT 12.704 26.676 12.736 29.184 ;
  LAYER M3 ;
        RECT 12.64 26.676 12.672 29.184 ;
  LAYER M3 ;
        RECT 12.544 26.676 12.576 29.184 ;
  LAYER M1 ;
        RECT 14.959 26.712 14.961 29.148 ;
  LAYER M1 ;
        RECT 14.879 26.712 14.881 29.148 ;
  LAYER M1 ;
        RECT 14.799 26.712 14.801 29.148 ;
  LAYER M1 ;
        RECT 14.719 26.712 14.721 29.148 ;
  LAYER M1 ;
        RECT 14.639 26.712 14.641 29.148 ;
  LAYER M1 ;
        RECT 14.559 26.712 14.561 29.148 ;
  LAYER M1 ;
        RECT 14.479 26.712 14.481 29.148 ;
  LAYER M1 ;
        RECT 14.399 26.712 14.401 29.148 ;
  LAYER M1 ;
        RECT 14.319 26.712 14.321 29.148 ;
  LAYER M1 ;
        RECT 14.239 26.712 14.241 29.148 ;
  LAYER M1 ;
        RECT 14.159 26.712 14.161 29.148 ;
  LAYER M1 ;
        RECT 14.079 26.712 14.081 29.148 ;
  LAYER M1 ;
        RECT 13.999 26.712 14.001 29.148 ;
  LAYER M1 ;
        RECT 13.919 26.712 13.921 29.148 ;
  LAYER M1 ;
        RECT 13.839 26.712 13.841 29.148 ;
  LAYER M1 ;
        RECT 13.759 26.712 13.761 29.148 ;
  LAYER M1 ;
        RECT 13.679 26.712 13.681 29.148 ;
  LAYER M1 ;
        RECT 13.599 26.712 13.601 29.148 ;
  LAYER M1 ;
        RECT 13.519 26.712 13.521 29.148 ;
  LAYER M1 ;
        RECT 13.439 26.712 13.441 29.148 ;
  LAYER M1 ;
        RECT 13.359 26.712 13.361 29.148 ;
  LAYER M1 ;
        RECT 13.279 26.712 13.281 29.148 ;
  LAYER M1 ;
        RECT 13.199 26.712 13.201 29.148 ;
  LAYER M1 ;
        RECT 13.119 26.712 13.121 29.148 ;
  LAYER M1 ;
        RECT 13.039 26.712 13.041 29.148 ;
  LAYER M1 ;
        RECT 12.959 26.712 12.961 29.148 ;
  LAYER M1 ;
        RECT 12.879 26.712 12.881 29.148 ;
  LAYER M1 ;
        RECT 12.799 26.712 12.801 29.148 ;
  LAYER M1 ;
        RECT 12.719 26.712 12.721 29.148 ;
  LAYER M1 ;
        RECT 12.639 26.712 12.641 29.148 ;
  LAYER M2 ;
        RECT 12.56 26.711 14.96 26.713 ;
  LAYER M2 ;
        RECT 12.56 26.795 14.96 26.797 ;
  LAYER M2 ;
        RECT 12.56 26.879 14.96 26.881 ;
  LAYER M2 ;
        RECT 12.56 26.963 14.96 26.965 ;
  LAYER M2 ;
        RECT 12.56 27.047 14.96 27.049 ;
  LAYER M2 ;
        RECT 12.56 27.131 14.96 27.133 ;
  LAYER M2 ;
        RECT 12.56 27.215 14.96 27.217 ;
  LAYER M2 ;
        RECT 12.56 27.299 14.96 27.301 ;
  LAYER M2 ;
        RECT 12.56 27.383 14.96 27.385 ;
  LAYER M2 ;
        RECT 12.56 27.467 14.96 27.469 ;
  LAYER M2 ;
        RECT 12.56 27.551 14.96 27.553 ;
  LAYER M2 ;
        RECT 12.56 27.635 14.96 27.637 ;
  LAYER M2 ;
        RECT 12.56 27.7185 14.96 27.7205 ;
  LAYER M2 ;
        RECT 12.56 27.803 14.96 27.805 ;
  LAYER M2 ;
        RECT 12.56 27.887 14.96 27.889 ;
  LAYER M2 ;
        RECT 12.56 27.971 14.96 27.973 ;
  LAYER M2 ;
        RECT 12.56 28.055 14.96 28.057 ;
  LAYER M2 ;
        RECT 12.56 28.139 14.96 28.141 ;
  LAYER M2 ;
        RECT 12.56 28.223 14.96 28.225 ;
  LAYER M2 ;
        RECT 12.56 28.307 14.96 28.309 ;
  LAYER M2 ;
        RECT 12.56 28.391 14.96 28.393 ;
  LAYER M2 ;
        RECT 12.56 28.475 14.96 28.477 ;
  LAYER M2 ;
        RECT 12.56 28.559 14.96 28.561 ;
  LAYER M2 ;
        RECT 12.56 28.643 14.96 28.645 ;
  LAYER M2 ;
        RECT 12.56 28.727 14.96 28.729 ;
  LAYER M2 ;
        RECT 12.56 28.811 14.96 28.813 ;
  LAYER M2 ;
        RECT 12.56 28.895 14.96 28.897 ;
  LAYER M2 ;
        RECT 12.56 28.979 14.96 28.981 ;
  LAYER M2 ;
        RECT 12.56 29.063 14.96 29.065 ;
  LAYER M1 ;
        RECT 12.064 17.856 12.096 20.364 ;
  LAYER M1 ;
        RECT 12 17.856 12.032 20.364 ;
  LAYER M1 ;
        RECT 11.936 17.856 11.968 20.364 ;
  LAYER M1 ;
        RECT 11.872 17.856 11.904 20.364 ;
  LAYER M1 ;
        RECT 11.808 17.856 11.84 20.364 ;
  LAYER M1 ;
        RECT 11.744 17.856 11.776 20.364 ;
  LAYER M1 ;
        RECT 11.68 17.856 11.712 20.364 ;
  LAYER M1 ;
        RECT 11.616 17.856 11.648 20.364 ;
  LAYER M1 ;
        RECT 11.552 17.856 11.584 20.364 ;
  LAYER M1 ;
        RECT 11.488 17.856 11.52 20.364 ;
  LAYER M1 ;
        RECT 11.424 17.856 11.456 20.364 ;
  LAYER M1 ;
        RECT 11.36 17.856 11.392 20.364 ;
  LAYER M1 ;
        RECT 11.296 17.856 11.328 20.364 ;
  LAYER M1 ;
        RECT 11.232 17.856 11.264 20.364 ;
  LAYER M1 ;
        RECT 11.168 17.856 11.2 20.364 ;
  LAYER M1 ;
        RECT 11.104 17.856 11.136 20.364 ;
  LAYER M1 ;
        RECT 11.04 17.856 11.072 20.364 ;
  LAYER M1 ;
        RECT 10.976 17.856 11.008 20.364 ;
  LAYER M1 ;
        RECT 10.912 17.856 10.944 20.364 ;
  LAYER M1 ;
        RECT 10.848 17.856 10.88 20.364 ;
  LAYER M1 ;
        RECT 10.784 17.856 10.816 20.364 ;
  LAYER M1 ;
        RECT 10.72 17.856 10.752 20.364 ;
  LAYER M1 ;
        RECT 10.656 17.856 10.688 20.364 ;
  LAYER M1 ;
        RECT 10.592 17.856 10.624 20.364 ;
  LAYER M1 ;
        RECT 10.528 17.856 10.56 20.364 ;
  LAYER M1 ;
        RECT 10.464 17.856 10.496 20.364 ;
  LAYER M1 ;
        RECT 10.4 17.856 10.432 20.364 ;
  LAYER M1 ;
        RECT 10.336 17.856 10.368 20.364 ;
  LAYER M1 ;
        RECT 10.272 17.856 10.304 20.364 ;
  LAYER M1 ;
        RECT 10.208 17.856 10.24 20.364 ;
  LAYER M1 ;
        RECT 10.144 17.856 10.176 20.364 ;
  LAYER M1 ;
        RECT 10.08 17.856 10.112 20.364 ;
  LAYER M1 ;
        RECT 10.016 17.856 10.048 20.364 ;
  LAYER M1 ;
        RECT 9.952 17.856 9.984 20.364 ;
  LAYER M1 ;
        RECT 9.888 17.856 9.92 20.364 ;
  LAYER M1 ;
        RECT 9.824 17.856 9.856 20.364 ;
  LAYER M1 ;
        RECT 9.76 17.856 9.792 20.364 ;
  LAYER M2 ;
        RECT 9.644 17.94 12.116 17.972 ;
  LAYER M2 ;
        RECT 9.644 18.004 12.116 18.036 ;
  LAYER M2 ;
        RECT 9.644 18.068 12.116 18.1 ;
  LAYER M2 ;
        RECT 9.644 18.132 12.116 18.164 ;
  LAYER M2 ;
        RECT 9.644 18.196 12.116 18.228 ;
  LAYER M2 ;
        RECT 9.644 18.26 12.116 18.292 ;
  LAYER M2 ;
        RECT 9.644 18.324 12.116 18.356 ;
  LAYER M2 ;
        RECT 9.644 18.388 12.116 18.42 ;
  LAYER M2 ;
        RECT 9.644 18.452 12.116 18.484 ;
  LAYER M2 ;
        RECT 9.644 18.516 12.116 18.548 ;
  LAYER M2 ;
        RECT 9.644 18.58 12.116 18.612 ;
  LAYER M2 ;
        RECT 9.644 18.644 12.116 18.676 ;
  LAYER M2 ;
        RECT 9.644 18.708 12.116 18.74 ;
  LAYER M2 ;
        RECT 9.644 18.772 12.116 18.804 ;
  LAYER M2 ;
        RECT 9.644 18.836 12.116 18.868 ;
  LAYER M2 ;
        RECT 9.644 18.9 12.116 18.932 ;
  LAYER M2 ;
        RECT 9.644 18.964 12.116 18.996 ;
  LAYER M2 ;
        RECT 9.644 19.028 12.116 19.06 ;
  LAYER M2 ;
        RECT 9.644 19.092 12.116 19.124 ;
  LAYER M2 ;
        RECT 9.644 19.156 12.116 19.188 ;
  LAYER M2 ;
        RECT 9.644 19.22 12.116 19.252 ;
  LAYER M2 ;
        RECT 9.644 19.284 12.116 19.316 ;
  LAYER M2 ;
        RECT 9.644 19.348 12.116 19.38 ;
  LAYER M2 ;
        RECT 9.644 19.412 12.116 19.444 ;
  LAYER M2 ;
        RECT 9.644 19.476 12.116 19.508 ;
  LAYER M2 ;
        RECT 9.644 19.54 12.116 19.572 ;
  LAYER M2 ;
        RECT 9.644 19.604 12.116 19.636 ;
  LAYER M2 ;
        RECT 9.644 19.668 12.116 19.7 ;
  LAYER M2 ;
        RECT 9.644 19.732 12.116 19.764 ;
  LAYER M2 ;
        RECT 9.644 19.796 12.116 19.828 ;
  LAYER M2 ;
        RECT 9.644 19.86 12.116 19.892 ;
  LAYER M2 ;
        RECT 9.644 19.924 12.116 19.956 ;
  LAYER M2 ;
        RECT 9.644 19.988 12.116 20.02 ;
  LAYER M2 ;
        RECT 9.644 20.052 12.116 20.084 ;
  LAYER M2 ;
        RECT 9.644 20.116 12.116 20.148 ;
  LAYER M2 ;
        RECT 9.644 20.18 12.116 20.212 ;
  LAYER M3 ;
        RECT 12.064 17.856 12.096 20.364 ;
  LAYER M3 ;
        RECT 12 17.856 12.032 20.364 ;
  LAYER M3 ;
        RECT 11.936 17.856 11.968 20.364 ;
  LAYER M3 ;
        RECT 11.872 17.856 11.904 20.364 ;
  LAYER M3 ;
        RECT 11.808 17.856 11.84 20.364 ;
  LAYER M3 ;
        RECT 11.744 17.856 11.776 20.364 ;
  LAYER M3 ;
        RECT 11.68 17.856 11.712 20.364 ;
  LAYER M3 ;
        RECT 11.616 17.856 11.648 20.364 ;
  LAYER M3 ;
        RECT 11.552 17.856 11.584 20.364 ;
  LAYER M3 ;
        RECT 11.488 17.856 11.52 20.364 ;
  LAYER M3 ;
        RECT 11.424 17.856 11.456 20.364 ;
  LAYER M3 ;
        RECT 11.36 17.856 11.392 20.364 ;
  LAYER M3 ;
        RECT 11.296 17.856 11.328 20.364 ;
  LAYER M3 ;
        RECT 11.232 17.856 11.264 20.364 ;
  LAYER M3 ;
        RECT 11.168 17.856 11.2 20.364 ;
  LAYER M3 ;
        RECT 11.104 17.856 11.136 20.364 ;
  LAYER M3 ;
        RECT 11.04 17.856 11.072 20.364 ;
  LAYER M3 ;
        RECT 10.976 17.856 11.008 20.364 ;
  LAYER M3 ;
        RECT 10.912 17.856 10.944 20.364 ;
  LAYER M3 ;
        RECT 10.848 17.856 10.88 20.364 ;
  LAYER M3 ;
        RECT 10.784 17.856 10.816 20.364 ;
  LAYER M3 ;
        RECT 10.72 17.856 10.752 20.364 ;
  LAYER M3 ;
        RECT 10.656 17.856 10.688 20.364 ;
  LAYER M3 ;
        RECT 10.592 17.856 10.624 20.364 ;
  LAYER M3 ;
        RECT 10.528 17.856 10.56 20.364 ;
  LAYER M3 ;
        RECT 10.464 17.856 10.496 20.364 ;
  LAYER M3 ;
        RECT 10.4 17.856 10.432 20.364 ;
  LAYER M3 ;
        RECT 10.336 17.856 10.368 20.364 ;
  LAYER M3 ;
        RECT 10.272 17.856 10.304 20.364 ;
  LAYER M3 ;
        RECT 10.208 17.856 10.24 20.364 ;
  LAYER M3 ;
        RECT 10.144 17.856 10.176 20.364 ;
  LAYER M3 ;
        RECT 10.08 17.856 10.112 20.364 ;
  LAYER M3 ;
        RECT 10.016 17.856 10.048 20.364 ;
  LAYER M3 ;
        RECT 9.952 17.856 9.984 20.364 ;
  LAYER M3 ;
        RECT 9.888 17.856 9.92 20.364 ;
  LAYER M3 ;
        RECT 9.824 17.856 9.856 20.364 ;
  LAYER M3 ;
        RECT 9.76 17.856 9.792 20.364 ;
  LAYER M3 ;
        RECT 9.664 17.856 9.696 20.364 ;
  LAYER M1 ;
        RECT 12.079 17.892 12.081 20.328 ;
  LAYER M1 ;
        RECT 11.999 17.892 12.001 20.328 ;
  LAYER M1 ;
        RECT 11.919 17.892 11.921 20.328 ;
  LAYER M1 ;
        RECT 11.839 17.892 11.841 20.328 ;
  LAYER M1 ;
        RECT 11.759 17.892 11.761 20.328 ;
  LAYER M1 ;
        RECT 11.679 17.892 11.681 20.328 ;
  LAYER M1 ;
        RECT 11.599 17.892 11.601 20.328 ;
  LAYER M1 ;
        RECT 11.519 17.892 11.521 20.328 ;
  LAYER M1 ;
        RECT 11.439 17.892 11.441 20.328 ;
  LAYER M1 ;
        RECT 11.359 17.892 11.361 20.328 ;
  LAYER M1 ;
        RECT 11.279 17.892 11.281 20.328 ;
  LAYER M1 ;
        RECT 11.199 17.892 11.201 20.328 ;
  LAYER M1 ;
        RECT 11.119 17.892 11.121 20.328 ;
  LAYER M1 ;
        RECT 11.039 17.892 11.041 20.328 ;
  LAYER M1 ;
        RECT 10.959 17.892 10.961 20.328 ;
  LAYER M1 ;
        RECT 10.879 17.892 10.881 20.328 ;
  LAYER M1 ;
        RECT 10.799 17.892 10.801 20.328 ;
  LAYER M1 ;
        RECT 10.719 17.892 10.721 20.328 ;
  LAYER M1 ;
        RECT 10.639 17.892 10.641 20.328 ;
  LAYER M1 ;
        RECT 10.559 17.892 10.561 20.328 ;
  LAYER M1 ;
        RECT 10.479 17.892 10.481 20.328 ;
  LAYER M1 ;
        RECT 10.399 17.892 10.401 20.328 ;
  LAYER M1 ;
        RECT 10.319 17.892 10.321 20.328 ;
  LAYER M1 ;
        RECT 10.239 17.892 10.241 20.328 ;
  LAYER M1 ;
        RECT 10.159 17.892 10.161 20.328 ;
  LAYER M1 ;
        RECT 10.079 17.892 10.081 20.328 ;
  LAYER M1 ;
        RECT 9.999 17.892 10.001 20.328 ;
  LAYER M1 ;
        RECT 9.919 17.892 9.921 20.328 ;
  LAYER M1 ;
        RECT 9.839 17.892 9.841 20.328 ;
  LAYER M1 ;
        RECT 9.759 17.892 9.761 20.328 ;
  LAYER M2 ;
        RECT 9.68 17.891 12.08 17.893 ;
  LAYER M2 ;
        RECT 9.68 17.975 12.08 17.977 ;
  LAYER M2 ;
        RECT 9.68 18.059 12.08 18.061 ;
  LAYER M2 ;
        RECT 9.68 18.143 12.08 18.145 ;
  LAYER M2 ;
        RECT 9.68 18.227 12.08 18.229 ;
  LAYER M2 ;
        RECT 9.68 18.311 12.08 18.313 ;
  LAYER M2 ;
        RECT 9.68 18.395 12.08 18.397 ;
  LAYER M2 ;
        RECT 9.68 18.479 12.08 18.481 ;
  LAYER M2 ;
        RECT 9.68 18.563 12.08 18.565 ;
  LAYER M2 ;
        RECT 9.68 18.647 12.08 18.649 ;
  LAYER M2 ;
        RECT 9.68 18.731 12.08 18.733 ;
  LAYER M2 ;
        RECT 9.68 18.815 12.08 18.817 ;
  LAYER M2 ;
        RECT 9.68 18.8985 12.08 18.9005 ;
  LAYER M2 ;
        RECT 9.68 18.983 12.08 18.985 ;
  LAYER M2 ;
        RECT 9.68 19.067 12.08 19.069 ;
  LAYER M2 ;
        RECT 9.68 19.151 12.08 19.153 ;
  LAYER M2 ;
        RECT 9.68 19.235 12.08 19.237 ;
  LAYER M2 ;
        RECT 9.68 19.319 12.08 19.321 ;
  LAYER M2 ;
        RECT 9.68 19.403 12.08 19.405 ;
  LAYER M2 ;
        RECT 9.68 19.487 12.08 19.489 ;
  LAYER M2 ;
        RECT 9.68 19.571 12.08 19.573 ;
  LAYER M2 ;
        RECT 9.68 19.655 12.08 19.657 ;
  LAYER M2 ;
        RECT 9.68 19.739 12.08 19.741 ;
  LAYER M2 ;
        RECT 9.68 19.823 12.08 19.825 ;
  LAYER M2 ;
        RECT 9.68 19.907 12.08 19.909 ;
  LAYER M2 ;
        RECT 9.68 19.991 12.08 19.993 ;
  LAYER M2 ;
        RECT 9.68 20.075 12.08 20.077 ;
  LAYER M2 ;
        RECT 9.68 20.159 12.08 20.161 ;
  LAYER M2 ;
        RECT 9.68 20.243 12.08 20.245 ;
  LAYER M1 ;
        RECT 12.064 20.796 12.096 23.304 ;
  LAYER M1 ;
        RECT 12 20.796 12.032 23.304 ;
  LAYER M1 ;
        RECT 11.936 20.796 11.968 23.304 ;
  LAYER M1 ;
        RECT 11.872 20.796 11.904 23.304 ;
  LAYER M1 ;
        RECT 11.808 20.796 11.84 23.304 ;
  LAYER M1 ;
        RECT 11.744 20.796 11.776 23.304 ;
  LAYER M1 ;
        RECT 11.68 20.796 11.712 23.304 ;
  LAYER M1 ;
        RECT 11.616 20.796 11.648 23.304 ;
  LAYER M1 ;
        RECT 11.552 20.796 11.584 23.304 ;
  LAYER M1 ;
        RECT 11.488 20.796 11.52 23.304 ;
  LAYER M1 ;
        RECT 11.424 20.796 11.456 23.304 ;
  LAYER M1 ;
        RECT 11.36 20.796 11.392 23.304 ;
  LAYER M1 ;
        RECT 11.296 20.796 11.328 23.304 ;
  LAYER M1 ;
        RECT 11.232 20.796 11.264 23.304 ;
  LAYER M1 ;
        RECT 11.168 20.796 11.2 23.304 ;
  LAYER M1 ;
        RECT 11.104 20.796 11.136 23.304 ;
  LAYER M1 ;
        RECT 11.04 20.796 11.072 23.304 ;
  LAYER M1 ;
        RECT 10.976 20.796 11.008 23.304 ;
  LAYER M1 ;
        RECT 10.912 20.796 10.944 23.304 ;
  LAYER M1 ;
        RECT 10.848 20.796 10.88 23.304 ;
  LAYER M1 ;
        RECT 10.784 20.796 10.816 23.304 ;
  LAYER M1 ;
        RECT 10.72 20.796 10.752 23.304 ;
  LAYER M1 ;
        RECT 10.656 20.796 10.688 23.304 ;
  LAYER M1 ;
        RECT 10.592 20.796 10.624 23.304 ;
  LAYER M1 ;
        RECT 10.528 20.796 10.56 23.304 ;
  LAYER M1 ;
        RECT 10.464 20.796 10.496 23.304 ;
  LAYER M1 ;
        RECT 10.4 20.796 10.432 23.304 ;
  LAYER M1 ;
        RECT 10.336 20.796 10.368 23.304 ;
  LAYER M1 ;
        RECT 10.272 20.796 10.304 23.304 ;
  LAYER M1 ;
        RECT 10.208 20.796 10.24 23.304 ;
  LAYER M1 ;
        RECT 10.144 20.796 10.176 23.304 ;
  LAYER M1 ;
        RECT 10.08 20.796 10.112 23.304 ;
  LAYER M1 ;
        RECT 10.016 20.796 10.048 23.304 ;
  LAYER M1 ;
        RECT 9.952 20.796 9.984 23.304 ;
  LAYER M1 ;
        RECT 9.888 20.796 9.92 23.304 ;
  LAYER M1 ;
        RECT 9.824 20.796 9.856 23.304 ;
  LAYER M1 ;
        RECT 9.76 20.796 9.792 23.304 ;
  LAYER M2 ;
        RECT 9.644 20.88 12.116 20.912 ;
  LAYER M2 ;
        RECT 9.644 20.944 12.116 20.976 ;
  LAYER M2 ;
        RECT 9.644 21.008 12.116 21.04 ;
  LAYER M2 ;
        RECT 9.644 21.072 12.116 21.104 ;
  LAYER M2 ;
        RECT 9.644 21.136 12.116 21.168 ;
  LAYER M2 ;
        RECT 9.644 21.2 12.116 21.232 ;
  LAYER M2 ;
        RECT 9.644 21.264 12.116 21.296 ;
  LAYER M2 ;
        RECT 9.644 21.328 12.116 21.36 ;
  LAYER M2 ;
        RECT 9.644 21.392 12.116 21.424 ;
  LAYER M2 ;
        RECT 9.644 21.456 12.116 21.488 ;
  LAYER M2 ;
        RECT 9.644 21.52 12.116 21.552 ;
  LAYER M2 ;
        RECT 9.644 21.584 12.116 21.616 ;
  LAYER M2 ;
        RECT 9.644 21.648 12.116 21.68 ;
  LAYER M2 ;
        RECT 9.644 21.712 12.116 21.744 ;
  LAYER M2 ;
        RECT 9.644 21.776 12.116 21.808 ;
  LAYER M2 ;
        RECT 9.644 21.84 12.116 21.872 ;
  LAYER M2 ;
        RECT 9.644 21.904 12.116 21.936 ;
  LAYER M2 ;
        RECT 9.644 21.968 12.116 22 ;
  LAYER M2 ;
        RECT 9.644 22.032 12.116 22.064 ;
  LAYER M2 ;
        RECT 9.644 22.096 12.116 22.128 ;
  LAYER M2 ;
        RECT 9.644 22.16 12.116 22.192 ;
  LAYER M2 ;
        RECT 9.644 22.224 12.116 22.256 ;
  LAYER M2 ;
        RECT 9.644 22.288 12.116 22.32 ;
  LAYER M2 ;
        RECT 9.644 22.352 12.116 22.384 ;
  LAYER M2 ;
        RECT 9.644 22.416 12.116 22.448 ;
  LAYER M2 ;
        RECT 9.644 22.48 12.116 22.512 ;
  LAYER M2 ;
        RECT 9.644 22.544 12.116 22.576 ;
  LAYER M2 ;
        RECT 9.644 22.608 12.116 22.64 ;
  LAYER M2 ;
        RECT 9.644 22.672 12.116 22.704 ;
  LAYER M2 ;
        RECT 9.644 22.736 12.116 22.768 ;
  LAYER M2 ;
        RECT 9.644 22.8 12.116 22.832 ;
  LAYER M2 ;
        RECT 9.644 22.864 12.116 22.896 ;
  LAYER M2 ;
        RECT 9.644 22.928 12.116 22.96 ;
  LAYER M2 ;
        RECT 9.644 22.992 12.116 23.024 ;
  LAYER M2 ;
        RECT 9.644 23.056 12.116 23.088 ;
  LAYER M2 ;
        RECT 9.644 23.12 12.116 23.152 ;
  LAYER M3 ;
        RECT 12.064 20.796 12.096 23.304 ;
  LAYER M3 ;
        RECT 12 20.796 12.032 23.304 ;
  LAYER M3 ;
        RECT 11.936 20.796 11.968 23.304 ;
  LAYER M3 ;
        RECT 11.872 20.796 11.904 23.304 ;
  LAYER M3 ;
        RECT 11.808 20.796 11.84 23.304 ;
  LAYER M3 ;
        RECT 11.744 20.796 11.776 23.304 ;
  LAYER M3 ;
        RECT 11.68 20.796 11.712 23.304 ;
  LAYER M3 ;
        RECT 11.616 20.796 11.648 23.304 ;
  LAYER M3 ;
        RECT 11.552 20.796 11.584 23.304 ;
  LAYER M3 ;
        RECT 11.488 20.796 11.52 23.304 ;
  LAYER M3 ;
        RECT 11.424 20.796 11.456 23.304 ;
  LAYER M3 ;
        RECT 11.36 20.796 11.392 23.304 ;
  LAYER M3 ;
        RECT 11.296 20.796 11.328 23.304 ;
  LAYER M3 ;
        RECT 11.232 20.796 11.264 23.304 ;
  LAYER M3 ;
        RECT 11.168 20.796 11.2 23.304 ;
  LAYER M3 ;
        RECT 11.104 20.796 11.136 23.304 ;
  LAYER M3 ;
        RECT 11.04 20.796 11.072 23.304 ;
  LAYER M3 ;
        RECT 10.976 20.796 11.008 23.304 ;
  LAYER M3 ;
        RECT 10.912 20.796 10.944 23.304 ;
  LAYER M3 ;
        RECT 10.848 20.796 10.88 23.304 ;
  LAYER M3 ;
        RECT 10.784 20.796 10.816 23.304 ;
  LAYER M3 ;
        RECT 10.72 20.796 10.752 23.304 ;
  LAYER M3 ;
        RECT 10.656 20.796 10.688 23.304 ;
  LAYER M3 ;
        RECT 10.592 20.796 10.624 23.304 ;
  LAYER M3 ;
        RECT 10.528 20.796 10.56 23.304 ;
  LAYER M3 ;
        RECT 10.464 20.796 10.496 23.304 ;
  LAYER M3 ;
        RECT 10.4 20.796 10.432 23.304 ;
  LAYER M3 ;
        RECT 10.336 20.796 10.368 23.304 ;
  LAYER M3 ;
        RECT 10.272 20.796 10.304 23.304 ;
  LAYER M3 ;
        RECT 10.208 20.796 10.24 23.304 ;
  LAYER M3 ;
        RECT 10.144 20.796 10.176 23.304 ;
  LAYER M3 ;
        RECT 10.08 20.796 10.112 23.304 ;
  LAYER M3 ;
        RECT 10.016 20.796 10.048 23.304 ;
  LAYER M3 ;
        RECT 9.952 20.796 9.984 23.304 ;
  LAYER M3 ;
        RECT 9.888 20.796 9.92 23.304 ;
  LAYER M3 ;
        RECT 9.824 20.796 9.856 23.304 ;
  LAYER M3 ;
        RECT 9.76 20.796 9.792 23.304 ;
  LAYER M3 ;
        RECT 9.664 20.796 9.696 23.304 ;
  LAYER M1 ;
        RECT 12.079 20.832 12.081 23.268 ;
  LAYER M1 ;
        RECT 11.999 20.832 12.001 23.268 ;
  LAYER M1 ;
        RECT 11.919 20.832 11.921 23.268 ;
  LAYER M1 ;
        RECT 11.839 20.832 11.841 23.268 ;
  LAYER M1 ;
        RECT 11.759 20.832 11.761 23.268 ;
  LAYER M1 ;
        RECT 11.679 20.832 11.681 23.268 ;
  LAYER M1 ;
        RECT 11.599 20.832 11.601 23.268 ;
  LAYER M1 ;
        RECT 11.519 20.832 11.521 23.268 ;
  LAYER M1 ;
        RECT 11.439 20.832 11.441 23.268 ;
  LAYER M1 ;
        RECT 11.359 20.832 11.361 23.268 ;
  LAYER M1 ;
        RECT 11.279 20.832 11.281 23.268 ;
  LAYER M1 ;
        RECT 11.199 20.832 11.201 23.268 ;
  LAYER M1 ;
        RECT 11.119 20.832 11.121 23.268 ;
  LAYER M1 ;
        RECT 11.039 20.832 11.041 23.268 ;
  LAYER M1 ;
        RECT 10.959 20.832 10.961 23.268 ;
  LAYER M1 ;
        RECT 10.879 20.832 10.881 23.268 ;
  LAYER M1 ;
        RECT 10.799 20.832 10.801 23.268 ;
  LAYER M1 ;
        RECT 10.719 20.832 10.721 23.268 ;
  LAYER M1 ;
        RECT 10.639 20.832 10.641 23.268 ;
  LAYER M1 ;
        RECT 10.559 20.832 10.561 23.268 ;
  LAYER M1 ;
        RECT 10.479 20.832 10.481 23.268 ;
  LAYER M1 ;
        RECT 10.399 20.832 10.401 23.268 ;
  LAYER M1 ;
        RECT 10.319 20.832 10.321 23.268 ;
  LAYER M1 ;
        RECT 10.239 20.832 10.241 23.268 ;
  LAYER M1 ;
        RECT 10.159 20.832 10.161 23.268 ;
  LAYER M1 ;
        RECT 10.079 20.832 10.081 23.268 ;
  LAYER M1 ;
        RECT 9.999 20.832 10.001 23.268 ;
  LAYER M1 ;
        RECT 9.919 20.832 9.921 23.268 ;
  LAYER M1 ;
        RECT 9.839 20.832 9.841 23.268 ;
  LAYER M1 ;
        RECT 9.759 20.832 9.761 23.268 ;
  LAYER M2 ;
        RECT 9.68 20.831 12.08 20.833 ;
  LAYER M2 ;
        RECT 9.68 20.915 12.08 20.917 ;
  LAYER M2 ;
        RECT 9.68 20.999 12.08 21.001 ;
  LAYER M2 ;
        RECT 9.68 21.083 12.08 21.085 ;
  LAYER M2 ;
        RECT 9.68 21.167 12.08 21.169 ;
  LAYER M2 ;
        RECT 9.68 21.251 12.08 21.253 ;
  LAYER M2 ;
        RECT 9.68 21.335 12.08 21.337 ;
  LAYER M2 ;
        RECT 9.68 21.419 12.08 21.421 ;
  LAYER M2 ;
        RECT 9.68 21.503 12.08 21.505 ;
  LAYER M2 ;
        RECT 9.68 21.587 12.08 21.589 ;
  LAYER M2 ;
        RECT 9.68 21.671 12.08 21.673 ;
  LAYER M2 ;
        RECT 9.68 21.755 12.08 21.757 ;
  LAYER M2 ;
        RECT 9.68 21.8385 12.08 21.8405 ;
  LAYER M2 ;
        RECT 9.68 21.923 12.08 21.925 ;
  LAYER M2 ;
        RECT 9.68 22.007 12.08 22.009 ;
  LAYER M2 ;
        RECT 9.68 22.091 12.08 22.093 ;
  LAYER M2 ;
        RECT 9.68 22.175 12.08 22.177 ;
  LAYER M2 ;
        RECT 9.68 22.259 12.08 22.261 ;
  LAYER M2 ;
        RECT 9.68 22.343 12.08 22.345 ;
  LAYER M2 ;
        RECT 9.68 22.427 12.08 22.429 ;
  LAYER M2 ;
        RECT 9.68 22.511 12.08 22.513 ;
  LAYER M2 ;
        RECT 9.68 22.595 12.08 22.597 ;
  LAYER M2 ;
        RECT 9.68 22.679 12.08 22.681 ;
  LAYER M2 ;
        RECT 9.68 22.763 12.08 22.765 ;
  LAYER M2 ;
        RECT 9.68 22.847 12.08 22.849 ;
  LAYER M2 ;
        RECT 9.68 22.931 12.08 22.933 ;
  LAYER M2 ;
        RECT 9.68 23.015 12.08 23.017 ;
  LAYER M2 ;
        RECT 9.68 23.099 12.08 23.101 ;
  LAYER M2 ;
        RECT 9.68 23.183 12.08 23.185 ;
  LAYER M1 ;
        RECT 12.064 23.736 12.096 26.244 ;
  LAYER M1 ;
        RECT 12 23.736 12.032 26.244 ;
  LAYER M1 ;
        RECT 11.936 23.736 11.968 26.244 ;
  LAYER M1 ;
        RECT 11.872 23.736 11.904 26.244 ;
  LAYER M1 ;
        RECT 11.808 23.736 11.84 26.244 ;
  LAYER M1 ;
        RECT 11.744 23.736 11.776 26.244 ;
  LAYER M1 ;
        RECT 11.68 23.736 11.712 26.244 ;
  LAYER M1 ;
        RECT 11.616 23.736 11.648 26.244 ;
  LAYER M1 ;
        RECT 11.552 23.736 11.584 26.244 ;
  LAYER M1 ;
        RECT 11.488 23.736 11.52 26.244 ;
  LAYER M1 ;
        RECT 11.424 23.736 11.456 26.244 ;
  LAYER M1 ;
        RECT 11.36 23.736 11.392 26.244 ;
  LAYER M1 ;
        RECT 11.296 23.736 11.328 26.244 ;
  LAYER M1 ;
        RECT 11.232 23.736 11.264 26.244 ;
  LAYER M1 ;
        RECT 11.168 23.736 11.2 26.244 ;
  LAYER M1 ;
        RECT 11.104 23.736 11.136 26.244 ;
  LAYER M1 ;
        RECT 11.04 23.736 11.072 26.244 ;
  LAYER M1 ;
        RECT 10.976 23.736 11.008 26.244 ;
  LAYER M1 ;
        RECT 10.912 23.736 10.944 26.244 ;
  LAYER M1 ;
        RECT 10.848 23.736 10.88 26.244 ;
  LAYER M1 ;
        RECT 10.784 23.736 10.816 26.244 ;
  LAYER M1 ;
        RECT 10.72 23.736 10.752 26.244 ;
  LAYER M1 ;
        RECT 10.656 23.736 10.688 26.244 ;
  LAYER M1 ;
        RECT 10.592 23.736 10.624 26.244 ;
  LAYER M1 ;
        RECT 10.528 23.736 10.56 26.244 ;
  LAYER M1 ;
        RECT 10.464 23.736 10.496 26.244 ;
  LAYER M1 ;
        RECT 10.4 23.736 10.432 26.244 ;
  LAYER M1 ;
        RECT 10.336 23.736 10.368 26.244 ;
  LAYER M1 ;
        RECT 10.272 23.736 10.304 26.244 ;
  LAYER M1 ;
        RECT 10.208 23.736 10.24 26.244 ;
  LAYER M1 ;
        RECT 10.144 23.736 10.176 26.244 ;
  LAYER M1 ;
        RECT 10.08 23.736 10.112 26.244 ;
  LAYER M1 ;
        RECT 10.016 23.736 10.048 26.244 ;
  LAYER M1 ;
        RECT 9.952 23.736 9.984 26.244 ;
  LAYER M1 ;
        RECT 9.888 23.736 9.92 26.244 ;
  LAYER M1 ;
        RECT 9.824 23.736 9.856 26.244 ;
  LAYER M1 ;
        RECT 9.76 23.736 9.792 26.244 ;
  LAYER M2 ;
        RECT 9.644 23.82 12.116 23.852 ;
  LAYER M2 ;
        RECT 9.644 23.884 12.116 23.916 ;
  LAYER M2 ;
        RECT 9.644 23.948 12.116 23.98 ;
  LAYER M2 ;
        RECT 9.644 24.012 12.116 24.044 ;
  LAYER M2 ;
        RECT 9.644 24.076 12.116 24.108 ;
  LAYER M2 ;
        RECT 9.644 24.14 12.116 24.172 ;
  LAYER M2 ;
        RECT 9.644 24.204 12.116 24.236 ;
  LAYER M2 ;
        RECT 9.644 24.268 12.116 24.3 ;
  LAYER M2 ;
        RECT 9.644 24.332 12.116 24.364 ;
  LAYER M2 ;
        RECT 9.644 24.396 12.116 24.428 ;
  LAYER M2 ;
        RECT 9.644 24.46 12.116 24.492 ;
  LAYER M2 ;
        RECT 9.644 24.524 12.116 24.556 ;
  LAYER M2 ;
        RECT 9.644 24.588 12.116 24.62 ;
  LAYER M2 ;
        RECT 9.644 24.652 12.116 24.684 ;
  LAYER M2 ;
        RECT 9.644 24.716 12.116 24.748 ;
  LAYER M2 ;
        RECT 9.644 24.78 12.116 24.812 ;
  LAYER M2 ;
        RECT 9.644 24.844 12.116 24.876 ;
  LAYER M2 ;
        RECT 9.644 24.908 12.116 24.94 ;
  LAYER M2 ;
        RECT 9.644 24.972 12.116 25.004 ;
  LAYER M2 ;
        RECT 9.644 25.036 12.116 25.068 ;
  LAYER M2 ;
        RECT 9.644 25.1 12.116 25.132 ;
  LAYER M2 ;
        RECT 9.644 25.164 12.116 25.196 ;
  LAYER M2 ;
        RECT 9.644 25.228 12.116 25.26 ;
  LAYER M2 ;
        RECT 9.644 25.292 12.116 25.324 ;
  LAYER M2 ;
        RECT 9.644 25.356 12.116 25.388 ;
  LAYER M2 ;
        RECT 9.644 25.42 12.116 25.452 ;
  LAYER M2 ;
        RECT 9.644 25.484 12.116 25.516 ;
  LAYER M2 ;
        RECT 9.644 25.548 12.116 25.58 ;
  LAYER M2 ;
        RECT 9.644 25.612 12.116 25.644 ;
  LAYER M2 ;
        RECT 9.644 25.676 12.116 25.708 ;
  LAYER M2 ;
        RECT 9.644 25.74 12.116 25.772 ;
  LAYER M2 ;
        RECT 9.644 25.804 12.116 25.836 ;
  LAYER M2 ;
        RECT 9.644 25.868 12.116 25.9 ;
  LAYER M2 ;
        RECT 9.644 25.932 12.116 25.964 ;
  LAYER M2 ;
        RECT 9.644 25.996 12.116 26.028 ;
  LAYER M2 ;
        RECT 9.644 26.06 12.116 26.092 ;
  LAYER M3 ;
        RECT 12.064 23.736 12.096 26.244 ;
  LAYER M3 ;
        RECT 12 23.736 12.032 26.244 ;
  LAYER M3 ;
        RECT 11.936 23.736 11.968 26.244 ;
  LAYER M3 ;
        RECT 11.872 23.736 11.904 26.244 ;
  LAYER M3 ;
        RECT 11.808 23.736 11.84 26.244 ;
  LAYER M3 ;
        RECT 11.744 23.736 11.776 26.244 ;
  LAYER M3 ;
        RECT 11.68 23.736 11.712 26.244 ;
  LAYER M3 ;
        RECT 11.616 23.736 11.648 26.244 ;
  LAYER M3 ;
        RECT 11.552 23.736 11.584 26.244 ;
  LAYER M3 ;
        RECT 11.488 23.736 11.52 26.244 ;
  LAYER M3 ;
        RECT 11.424 23.736 11.456 26.244 ;
  LAYER M3 ;
        RECT 11.36 23.736 11.392 26.244 ;
  LAYER M3 ;
        RECT 11.296 23.736 11.328 26.244 ;
  LAYER M3 ;
        RECT 11.232 23.736 11.264 26.244 ;
  LAYER M3 ;
        RECT 11.168 23.736 11.2 26.244 ;
  LAYER M3 ;
        RECT 11.104 23.736 11.136 26.244 ;
  LAYER M3 ;
        RECT 11.04 23.736 11.072 26.244 ;
  LAYER M3 ;
        RECT 10.976 23.736 11.008 26.244 ;
  LAYER M3 ;
        RECT 10.912 23.736 10.944 26.244 ;
  LAYER M3 ;
        RECT 10.848 23.736 10.88 26.244 ;
  LAYER M3 ;
        RECT 10.784 23.736 10.816 26.244 ;
  LAYER M3 ;
        RECT 10.72 23.736 10.752 26.244 ;
  LAYER M3 ;
        RECT 10.656 23.736 10.688 26.244 ;
  LAYER M3 ;
        RECT 10.592 23.736 10.624 26.244 ;
  LAYER M3 ;
        RECT 10.528 23.736 10.56 26.244 ;
  LAYER M3 ;
        RECT 10.464 23.736 10.496 26.244 ;
  LAYER M3 ;
        RECT 10.4 23.736 10.432 26.244 ;
  LAYER M3 ;
        RECT 10.336 23.736 10.368 26.244 ;
  LAYER M3 ;
        RECT 10.272 23.736 10.304 26.244 ;
  LAYER M3 ;
        RECT 10.208 23.736 10.24 26.244 ;
  LAYER M3 ;
        RECT 10.144 23.736 10.176 26.244 ;
  LAYER M3 ;
        RECT 10.08 23.736 10.112 26.244 ;
  LAYER M3 ;
        RECT 10.016 23.736 10.048 26.244 ;
  LAYER M3 ;
        RECT 9.952 23.736 9.984 26.244 ;
  LAYER M3 ;
        RECT 9.888 23.736 9.92 26.244 ;
  LAYER M3 ;
        RECT 9.824 23.736 9.856 26.244 ;
  LAYER M3 ;
        RECT 9.76 23.736 9.792 26.244 ;
  LAYER M3 ;
        RECT 9.664 23.736 9.696 26.244 ;
  LAYER M1 ;
        RECT 12.079 23.772 12.081 26.208 ;
  LAYER M1 ;
        RECT 11.999 23.772 12.001 26.208 ;
  LAYER M1 ;
        RECT 11.919 23.772 11.921 26.208 ;
  LAYER M1 ;
        RECT 11.839 23.772 11.841 26.208 ;
  LAYER M1 ;
        RECT 11.759 23.772 11.761 26.208 ;
  LAYER M1 ;
        RECT 11.679 23.772 11.681 26.208 ;
  LAYER M1 ;
        RECT 11.599 23.772 11.601 26.208 ;
  LAYER M1 ;
        RECT 11.519 23.772 11.521 26.208 ;
  LAYER M1 ;
        RECT 11.439 23.772 11.441 26.208 ;
  LAYER M1 ;
        RECT 11.359 23.772 11.361 26.208 ;
  LAYER M1 ;
        RECT 11.279 23.772 11.281 26.208 ;
  LAYER M1 ;
        RECT 11.199 23.772 11.201 26.208 ;
  LAYER M1 ;
        RECT 11.119 23.772 11.121 26.208 ;
  LAYER M1 ;
        RECT 11.039 23.772 11.041 26.208 ;
  LAYER M1 ;
        RECT 10.959 23.772 10.961 26.208 ;
  LAYER M1 ;
        RECT 10.879 23.772 10.881 26.208 ;
  LAYER M1 ;
        RECT 10.799 23.772 10.801 26.208 ;
  LAYER M1 ;
        RECT 10.719 23.772 10.721 26.208 ;
  LAYER M1 ;
        RECT 10.639 23.772 10.641 26.208 ;
  LAYER M1 ;
        RECT 10.559 23.772 10.561 26.208 ;
  LAYER M1 ;
        RECT 10.479 23.772 10.481 26.208 ;
  LAYER M1 ;
        RECT 10.399 23.772 10.401 26.208 ;
  LAYER M1 ;
        RECT 10.319 23.772 10.321 26.208 ;
  LAYER M1 ;
        RECT 10.239 23.772 10.241 26.208 ;
  LAYER M1 ;
        RECT 10.159 23.772 10.161 26.208 ;
  LAYER M1 ;
        RECT 10.079 23.772 10.081 26.208 ;
  LAYER M1 ;
        RECT 9.999 23.772 10.001 26.208 ;
  LAYER M1 ;
        RECT 9.919 23.772 9.921 26.208 ;
  LAYER M1 ;
        RECT 9.839 23.772 9.841 26.208 ;
  LAYER M1 ;
        RECT 9.759 23.772 9.761 26.208 ;
  LAYER M2 ;
        RECT 9.68 23.771 12.08 23.773 ;
  LAYER M2 ;
        RECT 9.68 23.855 12.08 23.857 ;
  LAYER M2 ;
        RECT 9.68 23.939 12.08 23.941 ;
  LAYER M2 ;
        RECT 9.68 24.023 12.08 24.025 ;
  LAYER M2 ;
        RECT 9.68 24.107 12.08 24.109 ;
  LAYER M2 ;
        RECT 9.68 24.191 12.08 24.193 ;
  LAYER M2 ;
        RECT 9.68 24.275 12.08 24.277 ;
  LAYER M2 ;
        RECT 9.68 24.359 12.08 24.361 ;
  LAYER M2 ;
        RECT 9.68 24.443 12.08 24.445 ;
  LAYER M2 ;
        RECT 9.68 24.527 12.08 24.529 ;
  LAYER M2 ;
        RECT 9.68 24.611 12.08 24.613 ;
  LAYER M2 ;
        RECT 9.68 24.695 12.08 24.697 ;
  LAYER M2 ;
        RECT 9.68 24.7785 12.08 24.7805 ;
  LAYER M2 ;
        RECT 9.68 24.863 12.08 24.865 ;
  LAYER M2 ;
        RECT 9.68 24.947 12.08 24.949 ;
  LAYER M2 ;
        RECT 9.68 25.031 12.08 25.033 ;
  LAYER M2 ;
        RECT 9.68 25.115 12.08 25.117 ;
  LAYER M2 ;
        RECT 9.68 25.199 12.08 25.201 ;
  LAYER M2 ;
        RECT 9.68 25.283 12.08 25.285 ;
  LAYER M2 ;
        RECT 9.68 25.367 12.08 25.369 ;
  LAYER M2 ;
        RECT 9.68 25.451 12.08 25.453 ;
  LAYER M2 ;
        RECT 9.68 25.535 12.08 25.537 ;
  LAYER M2 ;
        RECT 9.68 25.619 12.08 25.621 ;
  LAYER M2 ;
        RECT 9.68 25.703 12.08 25.705 ;
  LAYER M2 ;
        RECT 9.68 25.787 12.08 25.789 ;
  LAYER M2 ;
        RECT 9.68 25.871 12.08 25.873 ;
  LAYER M2 ;
        RECT 9.68 25.955 12.08 25.957 ;
  LAYER M2 ;
        RECT 9.68 26.039 12.08 26.041 ;
  LAYER M2 ;
        RECT 9.68 26.123 12.08 26.125 ;
  LAYER M1 ;
        RECT 12.064 26.676 12.096 29.184 ;
  LAYER M1 ;
        RECT 12 26.676 12.032 29.184 ;
  LAYER M1 ;
        RECT 11.936 26.676 11.968 29.184 ;
  LAYER M1 ;
        RECT 11.872 26.676 11.904 29.184 ;
  LAYER M1 ;
        RECT 11.808 26.676 11.84 29.184 ;
  LAYER M1 ;
        RECT 11.744 26.676 11.776 29.184 ;
  LAYER M1 ;
        RECT 11.68 26.676 11.712 29.184 ;
  LAYER M1 ;
        RECT 11.616 26.676 11.648 29.184 ;
  LAYER M1 ;
        RECT 11.552 26.676 11.584 29.184 ;
  LAYER M1 ;
        RECT 11.488 26.676 11.52 29.184 ;
  LAYER M1 ;
        RECT 11.424 26.676 11.456 29.184 ;
  LAYER M1 ;
        RECT 11.36 26.676 11.392 29.184 ;
  LAYER M1 ;
        RECT 11.296 26.676 11.328 29.184 ;
  LAYER M1 ;
        RECT 11.232 26.676 11.264 29.184 ;
  LAYER M1 ;
        RECT 11.168 26.676 11.2 29.184 ;
  LAYER M1 ;
        RECT 11.104 26.676 11.136 29.184 ;
  LAYER M1 ;
        RECT 11.04 26.676 11.072 29.184 ;
  LAYER M1 ;
        RECT 10.976 26.676 11.008 29.184 ;
  LAYER M1 ;
        RECT 10.912 26.676 10.944 29.184 ;
  LAYER M1 ;
        RECT 10.848 26.676 10.88 29.184 ;
  LAYER M1 ;
        RECT 10.784 26.676 10.816 29.184 ;
  LAYER M1 ;
        RECT 10.72 26.676 10.752 29.184 ;
  LAYER M1 ;
        RECT 10.656 26.676 10.688 29.184 ;
  LAYER M1 ;
        RECT 10.592 26.676 10.624 29.184 ;
  LAYER M1 ;
        RECT 10.528 26.676 10.56 29.184 ;
  LAYER M1 ;
        RECT 10.464 26.676 10.496 29.184 ;
  LAYER M1 ;
        RECT 10.4 26.676 10.432 29.184 ;
  LAYER M1 ;
        RECT 10.336 26.676 10.368 29.184 ;
  LAYER M1 ;
        RECT 10.272 26.676 10.304 29.184 ;
  LAYER M1 ;
        RECT 10.208 26.676 10.24 29.184 ;
  LAYER M1 ;
        RECT 10.144 26.676 10.176 29.184 ;
  LAYER M1 ;
        RECT 10.08 26.676 10.112 29.184 ;
  LAYER M1 ;
        RECT 10.016 26.676 10.048 29.184 ;
  LAYER M1 ;
        RECT 9.952 26.676 9.984 29.184 ;
  LAYER M1 ;
        RECT 9.888 26.676 9.92 29.184 ;
  LAYER M1 ;
        RECT 9.824 26.676 9.856 29.184 ;
  LAYER M1 ;
        RECT 9.76 26.676 9.792 29.184 ;
  LAYER M2 ;
        RECT 9.644 26.76 12.116 26.792 ;
  LAYER M2 ;
        RECT 9.644 26.824 12.116 26.856 ;
  LAYER M2 ;
        RECT 9.644 26.888 12.116 26.92 ;
  LAYER M2 ;
        RECT 9.644 26.952 12.116 26.984 ;
  LAYER M2 ;
        RECT 9.644 27.016 12.116 27.048 ;
  LAYER M2 ;
        RECT 9.644 27.08 12.116 27.112 ;
  LAYER M2 ;
        RECT 9.644 27.144 12.116 27.176 ;
  LAYER M2 ;
        RECT 9.644 27.208 12.116 27.24 ;
  LAYER M2 ;
        RECT 9.644 27.272 12.116 27.304 ;
  LAYER M2 ;
        RECT 9.644 27.336 12.116 27.368 ;
  LAYER M2 ;
        RECT 9.644 27.4 12.116 27.432 ;
  LAYER M2 ;
        RECT 9.644 27.464 12.116 27.496 ;
  LAYER M2 ;
        RECT 9.644 27.528 12.116 27.56 ;
  LAYER M2 ;
        RECT 9.644 27.592 12.116 27.624 ;
  LAYER M2 ;
        RECT 9.644 27.656 12.116 27.688 ;
  LAYER M2 ;
        RECT 9.644 27.72 12.116 27.752 ;
  LAYER M2 ;
        RECT 9.644 27.784 12.116 27.816 ;
  LAYER M2 ;
        RECT 9.644 27.848 12.116 27.88 ;
  LAYER M2 ;
        RECT 9.644 27.912 12.116 27.944 ;
  LAYER M2 ;
        RECT 9.644 27.976 12.116 28.008 ;
  LAYER M2 ;
        RECT 9.644 28.04 12.116 28.072 ;
  LAYER M2 ;
        RECT 9.644 28.104 12.116 28.136 ;
  LAYER M2 ;
        RECT 9.644 28.168 12.116 28.2 ;
  LAYER M2 ;
        RECT 9.644 28.232 12.116 28.264 ;
  LAYER M2 ;
        RECT 9.644 28.296 12.116 28.328 ;
  LAYER M2 ;
        RECT 9.644 28.36 12.116 28.392 ;
  LAYER M2 ;
        RECT 9.644 28.424 12.116 28.456 ;
  LAYER M2 ;
        RECT 9.644 28.488 12.116 28.52 ;
  LAYER M2 ;
        RECT 9.644 28.552 12.116 28.584 ;
  LAYER M2 ;
        RECT 9.644 28.616 12.116 28.648 ;
  LAYER M2 ;
        RECT 9.644 28.68 12.116 28.712 ;
  LAYER M2 ;
        RECT 9.644 28.744 12.116 28.776 ;
  LAYER M2 ;
        RECT 9.644 28.808 12.116 28.84 ;
  LAYER M2 ;
        RECT 9.644 28.872 12.116 28.904 ;
  LAYER M2 ;
        RECT 9.644 28.936 12.116 28.968 ;
  LAYER M2 ;
        RECT 9.644 29 12.116 29.032 ;
  LAYER M3 ;
        RECT 12.064 26.676 12.096 29.184 ;
  LAYER M3 ;
        RECT 12 26.676 12.032 29.184 ;
  LAYER M3 ;
        RECT 11.936 26.676 11.968 29.184 ;
  LAYER M3 ;
        RECT 11.872 26.676 11.904 29.184 ;
  LAYER M3 ;
        RECT 11.808 26.676 11.84 29.184 ;
  LAYER M3 ;
        RECT 11.744 26.676 11.776 29.184 ;
  LAYER M3 ;
        RECT 11.68 26.676 11.712 29.184 ;
  LAYER M3 ;
        RECT 11.616 26.676 11.648 29.184 ;
  LAYER M3 ;
        RECT 11.552 26.676 11.584 29.184 ;
  LAYER M3 ;
        RECT 11.488 26.676 11.52 29.184 ;
  LAYER M3 ;
        RECT 11.424 26.676 11.456 29.184 ;
  LAYER M3 ;
        RECT 11.36 26.676 11.392 29.184 ;
  LAYER M3 ;
        RECT 11.296 26.676 11.328 29.184 ;
  LAYER M3 ;
        RECT 11.232 26.676 11.264 29.184 ;
  LAYER M3 ;
        RECT 11.168 26.676 11.2 29.184 ;
  LAYER M3 ;
        RECT 11.104 26.676 11.136 29.184 ;
  LAYER M3 ;
        RECT 11.04 26.676 11.072 29.184 ;
  LAYER M3 ;
        RECT 10.976 26.676 11.008 29.184 ;
  LAYER M3 ;
        RECT 10.912 26.676 10.944 29.184 ;
  LAYER M3 ;
        RECT 10.848 26.676 10.88 29.184 ;
  LAYER M3 ;
        RECT 10.784 26.676 10.816 29.184 ;
  LAYER M3 ;
        RECT 10.72 26.676 10.752 29.184 ;
  LAYER M3 ;
        RECT 10.656 26.676 10.688 29.184 ;
  LAYER M3 ;
        RECT 10.592 26.676 10.624 29.184 ;
  LAYER M3 ;
        RECT 10.528 26.676 10.56 29.184 ;
  LAYER M3 ;
        RECT 10.464 26.676 10.496 29.184 ;
  LAYER M3 ;
        RECT 10.4 26.676 10.432 29.184 ;
  LAYER M3 ;
        RECT 10.336 26.676 10.368 29.184 ;
  LAYER M3 ;
        RECT 10.272 26.676 10.304 29.184 ;
  LAYER M3 ;
        RECT 10.208 26.676 10.24 29.184 ;
  LAYER M3 ;
        RECT 10.144 26.676 10.176 29.184 ;
  LAYER M3 ;
        RECT 10.08 26.676 10.112 29.184 ;
  LAYER M3 ;
        RECT 10.016 26.676 10.048 29.184 ;
  LAYER M3 ;
        RECT 9.952 26.676 9.984 29.184 ;
  LAYER M3 ;
        RECT 9.888 26.676 9.92 29.184 ;
  LAYER M3 ;
        RECT 9.824 26.676 9.856 29.184 ;
  LAYER M3 ;
        RECT 9.76 26.676 9.792 29.184 ;
  LAYER M3 ;
        RECT 9.664 26.676 9.696 29.184 ;
  LAYER M1 ;
        RECT 12.079 26.712 12.081 29.148 ;
  LAYER M1 ;
        RECT 11.999 26.712 12.001 29.148 ;
  LAYER M1 ;
        RECT 11.919 26.712 11.921 29.148 ;
  LAYER M1 ;
        RECT 11.839 26.712 11.841 29.148 ;
  LAYER M1 ;
        RECT 11.759 26.712 11.761 29.148 ;
  LAYER M1 ;
        RECT 11.679 26.712 11.681 29.148 ;
  LAYER M1 ;
        RECT 11.599 26.712 11.601 29.148 ;
  LAYER M1 ;
        RECT 11.519 26.712 11.521 29.148 ;
  LAYER M1 ;
        RECT 11.439 26.712 11.441 29.148 ;
  LAYER M1 ;
        RECT 11.359 26.712 11.361 29.148 ;
  LAYER M1 ;
        RECT 11.279 26.712 11.281 29.148 ;
  LAYER M1 ;
        RECT 11.199 26.712 11.201 29.148 ;
  LAYER M1 ;
        RECT 11.119 26.712 11.121 29.148 ;
  LAYER M1 ;
        RECT 11.039 26.712 11.041 29.148 ;
  LAYER M1 ;
        RECT 10.959 26.712 10.961 29.148 ;
  LAYER M1 ;
        RECT 10.879 26.712 10.881 29.148 ;
  LAYER M1 ;
        RECT 10.799 26.712 10.801 29.148 ;
  LAYER M1 ;
        RECT 10.719 26.712 10.721 29.148 ;
  LAYER M1 ;
        RECT 10.639 26.712 10.641 29.148 ;
  LAYER M1 ;
        RECT 10.559 26.712 10.561 29.148 ;
  LAYER M1 ;
        RECT 10.479 26.712 10.481 29.148 ;
  LAYER M1 ;
        RECT 10.399 26.712 10.401 29.148 ;
  LAYER M1 ;
        RECT 10.319 26.712 10.321 29.148 ;
  LAYER M1 ;
        RECT 10.239 26.712 10.241 29.148 ;
  LAYER M1 ;
        RECT 10.159 26.712 10.161 29.148 ;
  LAYER M1 ;
        RECT 10.079 26.712 10.081 29.148 ;
  LAYER M1 ;
        RECT 9.999 26.712 10.001 29.148 ;
  LAYER M1 ;
        RECT 9.919 26.712 9.921 29.148 ;
  LAYER M1 ;
        RECT 9.839 26.712 9.841 29.148 ;
  LAYER M1 ;
        RECT 9.759 26.712 9.761 29.148 ;
  LAYER M2 ;
        RECT 9.68 26.711 12.08 26.713 ;
  LAYER M2 ;
        RECT 9.68 26.795 12.08 26.797 ;
  LAYER M2 ;
        RECT 9.68 26.879 12.08 26.881 ;
  LAYER M2 ;
        RECT 9.68 26.963 12.08 26.965 ;
  LAYER M2 ;
        RECT 9.68 27.047 12.08 27.049 ;
  LAYER M2 ;
        RECT 9.68 27.131 12.08 27.133 ;
  LAYER M2 ;
        RECT 9.68 27.215 12.08 27.217 ;
  LAYER M2 ;
        RECT 9.68 27.299 12.08 27.301 ;
  LAYER M2 ;
        RECT 9.68 27.383 12.08 27.385 ;
  LAYER M2 ;
        RECT 9.68 27.467 12.08 27.469 ;
  LAYER M2 ;
        RECT 9.68 27.551 12.08 27.553 ;
  LAYER M2 ;
        RECT 9.68 27.635 12.08 27.637 ;
  LAYER M2 ;
        RECT 9.68 27.7185 12.08 27.7205 ;
  LAYER M2 ;
        RECT 9.68 27.803 12.08 27.805 ;
  LAYER M2 ;
        RECT 9.68 27.887 12.08 27.889 ;
  LAYER M2 ;
        RECT 9.68 27.971 12.08 27.973 ;
  LAYER M2 ;
        RECT 9.68 28.055 12.08 28.057 ;
  LAYER M2 ;
        RECT 9.68 28.139 12.08 28.141 ;
  LAYER M2 ;
        RECT 9.68 28.223 12.08 28.225 ;
  LAYER M2 ;
        RECT 9.68 28.307 12.08 28.309 ;
  LAYER M2 ;
        RECT 9.68 28.391 12.08 28.393 ;
  LAYER M2 ;
        RECT 9.68 28.475 12.08 28.477 ;
  LAYER M2 ;
        RECT 9.68 28.559 12.08 28.561 ;
  LAYER M2 ;
        RECT 9.68 28.643 12.08 28.645 ;
  LAYER M2 ;
        RECT 9.68 28.727 12.08 28.729 ;
  LAYER M2 ;
        RECT 9.68 28.811 12.08 28.813 ;
  LAYER M2 ;
        RECT 9.68 28.895 12.08 28.897 ;
  LAYER M2 ;
        RECT 9.68 28.979 12.08 28.981 ;
  LAYER M2 ;
        RECT 9.68 29.063 12.08 29.065 ;
  LAYER M1 ;
        RECT 9.184 17.856 9.216 20.364 ;
  LAYER M1 ;
        RECT 9.12 17.856 9.152 20.364 ;
  LAYER M1 ;
        RECT 9.056 17.856 9.088 20.364 ;
  LAYER M1 ;
        RECT 8.992 17.856 9.024 20.364 ;
  LAYER M1 ;
        RECT 8.928 17.856 8.96 20.364 ;
  LAYER M1 ;
        RECT 8.864 17.856 8.896 20.364 ;
  LAYER M1 ;
        RECT 8.8 17.856 8.832 20.364 ;
  LAYER M1 ;
        RECT 8.736 17.856 8.768 20.364 ;
  LAYER M1 ;
        RECT 8.672 17.856 8.704 20.364 ;
  LAYER M1 ;
        RECT 8.608 17.856 8.64 20.364 ;
  LAYER M1 ;
        RECT 8.544 17.856 8.576 20.364 ;
  LAYER M1 ;
        RECT 8.48 17.856 8.512 20.364 ;
  LAYER M1 ;
        RECT 8.416 17.856 8.448 20.364 ;
  LAYER M1 ;
        RECT 8.352 17.856 8.384 20.364 ;
  LAYER M1 ;
        RECT 8.288 17.856 8.32 20.364 ;
  LAYER M1 ;
        RECT 8.224 17.856 8.256 20.364 ;
  LAYER M1 ;
        RECT 8.16 17.856 8.192 20.364 ;
  LAYER M1 ;
        RECT 8.096 17.856 8.128 20.364 ;
  LAYER M1 ;
        RECT 8.032 17.856 8.064 20.364 ;
  LAYER M1 ;
        RECT 7.968 17.856 8 20.364 ;
  LAYER M1 ;
        RECT 7.904 17.856 7.936 20.364 ;
  LAYER M1 ;
        RECT 7.84 17.856 7.872 20.364 ;
  LAYER M1 ;
        RECT 7.776 17.856 7.808 20.364 ;
  LAYER M1 ;
        RECT 7.712 17.856 7.744 20.364 ;
  LAYER M1 ;
        RECT 7.648 17.856 7.68 20.364 ;
  LAYER M1 ;
        RECT 7.584 17.856 7.616 20.364 ;
  LAYER M1 ;
        RECT 7.52 17.856 7.552 20.364 ;
  LAYER M1 ;
        RECT 7.456 17.856 7.488 20.364 ;
  LAYER M1 ;
        RECT 7.392 17.856 7.424 20.364 ;
  LAYER M1 ;
        RECT 7.328 17.856 7.36 20.364 ;
  LAYER M1 ;
        RECT 7.264 17.856 7.296 20.364 ;
  LAYER M1 ;
        RECT 7.2 17.856 7.232 20.364 ;
  LAYER M1 ;
        RECT 7.136 17.856 7.168 20.364 ;
  LAYER M1 ;
        RECT 7.072 17.856 7.104 20.364 ;
  LAYER M1 ;
        RECT 7.008 17.856 7.04 20.364 ;
  LAYER M1 ;
        RECT 6.944 17.856 6.976 20.364 ;
  LAYER M1 ;
        RECT 6.88 17.856 6.912 20.364 ;
  LAYER M2 ;
        RECT 6.764 17.94 9.236 17.972 ;
  LAYER M2 ;
        RECT 6.764 18.004 9.236 18.036 ;
  LAYER M2 ;
        RECT 6.764 18.068 9.236 18.1 ;
  LAYER M2 ;
        RECT 6.764 18.132 9.236 18.164 ;
  LAYER M2 ;
        RECT 6.764 18.196 9.236 18.228 ;
  LAYER M2 ;
        RECT 6.764 18.26 9.236 18.292 ;
  LAYER M2 ;
        RECT 6.764 18.324 9.236 18.356 ;
  LAYER M2 ;
        RECT 6.764 18.388 9.236 18.42 ;
  LAYER M2 ;
        RECT 6.764 18.452 9.236 18.484 ;
  LAYER M2 ;
        RECT 6.764 18.516 9.236 18.548 ;
  LAYER M2 ;
        RECT 6.764 18.58 9.236 18.612 ;
  LAYER M2 ;
        RECT 6.764 18.644 9.236 18.676 ;
  LAYER M2 ;
        RECT 6.764 18.708 9.236 18.74 ;
  LAYER M2 ;
        RECT 6.764 18.772 9.236 18.804 ;
  LAYER M2 ;
        RECT 6.764 18.836 9.236 18.868 ;
  LAYER M2 ;
        RECT 6.764 18.9 9.236 18.932 ;
  LAYER M2 ;
        RECT 6.764 18.964 9.236 18.996 ;
  LAYER M2 ;
        RECT 6.764 19.028 9.236 19.06 ;
  LAYER M2 ;
        RECT 6.764 19.092 9.236 19.124 ;
  LAYER M2 ;
        RECT 6.764 19.156 9.236 19.188 ;
  LAYER M2 ;
        RECT 6.764 19.22 9.236 19.252 ;
  LAYER M2 ;
        RECT 6.764 19.284 9.236 19.316 ;
  LAYER M2 ;
        RECT 6.764 19.348 9.236 19.38 ;
  LAYER M2 ;
        RECT 6.764 19.412 9.236 19.444 ;
  LAYER M2 ;
        RECT 6.764 19.476 9.236 19.508 ;
  LAYER M2 ;
        RECT 6.764 19.54 9.236 19.572 ;
  LAYER M2 ;
        RECT 6.764 19.604 9.236 19.636 ;
  LAYER M2 ;
        RECT 6.764 19.668 9.236 19.7 ;
  LAYER M2 ;
        RECT 6.764 19.732 9.236 19.764 ;
  LAYER M2 ;
        RECT 6.764 19.796 9.236 19.828 ;
  LAYER M2 ;
        RECT 6.764 19.86 9.236 19.892 ;
  LAYER M2 ;
        RECT 6.764 19.924 9.236 19.956 ;
  LAYER M2 ;
        RECT 6.764 19.988 9.236 20.02 ;
  LAYER M2 ;
        RECT 6.764 20.052 9.236 20.084 ;
  LAYER M2 ;
        RECT 6.764 20.116 9.236 20.148 ;
  LAYER M2 ;
        RECT 6.764 20.18 9.236 20.212 ;
  LAYER M3 ;
        RECT 9.184 17.856 9.216 20.364 ;
  LAYER M3 ;
        RECT 9.12 17.856 9.152 20.364 ;
  LAYER M3 ;
        RECT 9.056 17.856 9.088 20.364 ;
  LAYER M3 ;
        RECT 8.992 17.856 9.024 20.364 ;
  LAYER M3 ;
        RECT 8.928 17.856 8.96 20.364 ;
  LAYER M3 ;
        RECT 8.864 17.856 8.896 20.364 ;
  LAYER M3 ;
        RECT 8.8 17.856 8.832 20.364 ;
  LAYER M3 ;
        RECT 8.736 17.856 8.768 20.364 ;
  LAYER M3 ;
        RECT 8.672 17.856 8.704 20.364 ;
  LAYER M3 ;
        RECT 8.608 17.856 8.64 20.364 ;
  LAYER M3 ;
        RECT 8.544 17.856 8.576 20.364 ;
  LAYER M3 ;
        RECT 8.48 17.856 8.512 20.364 ;
  LAYER M3 ;
        RECT 8.416 17.856 8.448 20.364 ;
  LAYER M3 ;
        RECT 8.352 17.856 8.384 20.364 ;
  LAYER M3 ;
        RECT 8.288 17.856 8.32 20.364 ;
  LAYER M3 ;
        RECT 8.224 17.856 8.256 20.364 ;
  LAYER M3 ;
        RECT 8.16 17.856 8.192 20.364 ;
  LAYER M3 ;
        RECT 8.096 17.856 8.128 20.364 ;
  LAYER M3 ;
        RECT 8.032 17.856 8.064 20.364 ;
  LAYER M3 ;
        RECT 7.968 17.856 8 20.364 ;
  LAYER M3 ;
        RECT 7.904 17.856 7.936 20.364 ;
  LAYER M3 ;
        RECT 7.84 17.856 7.872 20.364 ;
  LAYER M3 ;
        RECT 7.776 17.856 7.808 20.364 ;
  LAYER M3 ;
        RECT 7.712 17.856 7.744 20.364 ;
  LAYER M3 ;
        RECT 7.648 17.856 7.68 20.364 ;
  LAYER M3 ;
        RECT 7.584 17.856 7.616 20.364 ;
  LAYER M3 ;
        RECT 7.52 17.856 7.552 20.364 ;
  LAYER M3 ;
        RECT 7.456 17.856 7.488 20.364 ;
  LAYER M3 ;
        RECT 7.392 17.856 7.424 20.364 ;
  LAYER M3 ;
        RECT 7.328 17.856 7.36 20.364 ;
  LAYER M3 ;
        RECT 7.264 17.856 7.296 20.364 ;
  LAYER M3 ;
        RECT 7.2 17.856 7.232 20.364 ;
  LAYER M3 ;
        RECT 7.136 17.856 7.168 20.364 ;
  LAYER M3 ;
        RECT 7.072 17.856 7.104 20.364 ;
  LAYER M3 ;
        RECT 7.008 17.856 7.04 20.364 ;
  LAYER M3 ;
        RECT 6.944 17.856 6.976 20.364 ;
  LAYER M3 ;
        RECT 6.88 17.856 6.912 20.364 ;
  LAYER M3 ;
        RECT 6.784 17.856 6.816 20.364 ;
  LAYER M1 ;
        RECT 9.199 17.892 9.201 20.328 ;
  LAYER M1 ;
        RECT 9.119 17.892 9.121 20.328 ;
  LAYER M1 ;
        RECT 9.039 17.892 9.041 20.328 ;
  LAYER M1 ;
        RECT 8.959 17.892 8.961 20.328 ;
  LAYER M1 ;
        RECT 8.879 17.892 8.881 20.328 ;
  LAYER M1 ;
        RECT 8.799 17.892 8.801 20.328 ;
  LAYER M1 ;
        RECT 8.719 17.892 8.721 20.328 ;
  LAYER M1 ;
        RECT 8.639 17.892 8.641 20.328 ;
  LAYER M1 ;
        RECT 8.559 17.892 8.561 20.328 ;
  LAYER M1 ;
        RECT 8.479 17.892 8.481 20.328 ;
  LAYER M1 ;
        RECT 8.399 17.892 8.401 20.328 ;
  LAYER M1 ;
        RECT 8.319 17.892 8.321 20.328 ;
  LAYER M1 ;
        RECT 8.239 17.892 8.241 20.328 ;
  LAYER M1 ;
        RECT 8.159 17.892 8.161 20.328 ;
  LAYER M1 ;
        RECT 8.079 17.892 8.081 20.328 ;
  LAYER M1 ;
        RECT 7.999 17.892 8.001 20.328 ;
  LAYER M1 ;
        RECT 7.919 17.892 7.921 20.328 ;
  LAYER M1 ;
        RECT 7.839 17.892 7.841 20.328 ;
  LAYER M1 ;
        RECT 7.759 17.892 7.761 20.328 ;
  LAYER M1 ;
        RECT 7.679 17.892 7.681 20.328 ;
  LAYER M1 ;
        RECT 7.599 17.892 7.601 20.328 ;
  LAYER M1 ;
        RECT 7.519 17.892 7.521 20.328 ;
  LAYER M1 ;
        RECT 7.439 17.892 7.441 20.328 ;
  LAYER M1 ;
        RECT 7.359 17.892 7.361 20.328 ;
  LAYER M1 ;
        RECT 7.279 17.892 7.281 20.328 ;
  LAYER M1 ;
        RECT 7.199 17.892 7.201 20.328 ;
  LAYER M1 ;
        RECT 7.119 17.892 7.121 20.328 ;
  LAYER M1 ;
        RECT 7.039 17.892 7.041 20.328 ;
  LAYER M1 ;
        RECT 6.959 17.892 6.961 20.328 ;
  LAYER M1 ;
        RECT 6.879 17.892 6.881 20.328 ;
  LAYER M2 ;
        RECT 6.8 17.891 9.2 17.893 ;
  LAYER M2 ;
        RECT 6.8 17.975 9.2 17.977 ;
  LAYER M2 ;
        RECT 6.8 18.059 9.2 18.061 ;
  LAYER M2 ;
        RECT 6.8 18.143 9.2 18.145 ;
  LAYER M2 ;
        RECT 6.8 18.227 9.2 18.229 ;
  LAYER M2 ;
        RECT 6.8 18.311 9.2 18.313 ;
  LAYER M2 ;
        RECT 6.8 18.395 9.2 18.397 ;
  LAYER M2 ;
        RECT 6.8 18.479 9.2 18.481 ;
  LAYER M2 ;
        RECT 6.8 18.563 9.2 18.565 ;
  LAYER M2 ;
        RECT 6.8 18.647 9.2 18.649 ;
  LAYER M2 ;
        RECT 6.8 18.731 9.2 18.733 ;
  LAYER M2 ;
        RECT 6.8 18.815 9.2 18.817 ;
  LAYER M2 ;
        RECT 6.8 18.8985 9.2 18.9005 ;
  LAYER M2 ;
        RECT 6.8 18.983 9.2 18.985 ;
  LAYER M2 ;
        RECT 6.8 19.067 9.2 19.069 ;
  LAYER M2 ;
        RECT 6.8 19.151 9.2 19.153 ;
  LAYER M2 ;
        RECT 6.8 19.235 9.2 19.237 ;
  LAYER M2 ;
        RECT 6.8 19.319 9.2 19.321 ;
  LAYER M2 ;
        RECT 6.8 19.403 9.2 19.405 ;
  LAYER M2 ;
        RECT 6.8 19.487 9.2 19.489 ;
  LAYER M2 ;
        RECT 6.8 19.571 9.2 19.573 ;
  LAYER M2 ;
        RECT 6.8 19.655 9.2 19.657 ;
  LAYER M2 ;
        RECT 6.8 19.739 9.2 19.741 ;
  LAYER M2 ;
        RECT 6.8 19.823 9.2 19.825 ;
  LAYER M2 ;
        RECT 6.8 19.907 9.2 19.909 ;
  LAYER M2 ;
        RECT 6.8 19.991 9.2 19.993 ;
  LAYER M2 ;
        RECT 6.8 20.075 9.2 20.077 ;
  LAYER M2 ;
        RECT 6.8 20.159 9.2 20.161 ;
  LAYER M2 ;
        RECT 6.8 20.243 9.2 20.245 ;
  LAYER M1 ;
        RECT 9.184 20.796 9.216 23.304 ;
  LAYER M1 ;
        RECT 9.12 20.796 9.152 23.304 ;
  LAYER M1 ;
        RECT 9.056 20.796 9.088 23.304 ;
  LAYER M1 ;
        RECT 8.992 20.796 9.024 23.304 ;
  LAYER M1 ;
        RECT 8.928 20.796 8.96 23.304 ;
  LAYER M1 ;
        RECT 8.864 20.796 8.896 23.304 ;
  LAYER M1 ;
        RECT 8.8 20.796 8.832 23.304 ;
  LAYER M1 ;
        RECT 8.736 20.796 8.768 23.304 ;
  LAYER M1 ;
        RECT 8.672 20.796 8.704 23.304 ;
  LAYER M1 ;
        RECT 8.608 20.796 8.64 23.304 ;
  LAYER M1 ;
        RECT 8.544 20.796 8.576 23.304 ;
  LAYER M1 ;
        RECT 8.48 20.796 8.512 23.304 ;
  LAYER M1 ;
        RECT 8.416 20.796 8.448 23.304 ;
  LAYER M1 ;
        RECT 8.352 20.796 8.384 23.304 ;
  LAYER M1 ;
        RECT 8.288 20.796 8.32 23.304 ;
  LAYER M1 ;
        RECT 8.224 20.796 8.256 23.304 ;
  LAYER M1 ;
        RECT 8.16 20.796 8.192 23.304 ;
  LAYER M1 ;
        RECT 8.096 20.796 8.128 23.304 ;
  LAYER M1 ;
        RECT 8.032 20.796 8.064 23.304 ;
  LAYER M1 ;
        RECT 7.968 20.796 8 23.304 ;
  LAYER M1 ;
        RECT 7.904 20.796 7.936 23.304 ;
  LAYER M1 ;
        RECT 7.84 20.796 7.872 23.304 ;
  LAYER M1 ;
        RECT 7.776 20.796 7.808 23.304 ;
  LAYER M1 ;
        RECT 7.712 20.796 7.744 23.304 ;
  LAYER M1 ;
        RECT 7.648 20.796 7.68 23.304 ;
  LAYER M1 ;
        RECT 7.584 20.796 7.616 23.304 ;
  LAYER M1 ;
        RECT 7.52 20.796 7.552 23.304 ;
  LAYER M1 ;
        RECT 7.456 20.796 7.488 23.304 ;
  LAYER M1 ;
        RECT 7.392 20.796 7.424 23.304 ;
  LAYER M1 ;
        RECT 7.328 20.796 7.36 23.304 ;
  LAYER M1 ;
        RECT 7.264 20.796 7.296 23.304 ;
  LAYER M1 ;
        RECT 7.2 20.796 7.232 23.304 ;
  LAYER M1 ;
        RECT 7.136 20.796 7.168 23.304 ;
  LAYER M1 ;
        RECT 7.072 20.796 7.104 23.304 ;
  LAYER M1 ;
        RECT 7.008 20.796 7.04 23.304 ;
  LAYER M1 ;
        RECT 6.944 20.796 6.976 23.304 ;
  LAYER M1 ;
        RECT 6.88 20.796 6.912 23.304 ;
  LAYER M2 ;
        RECT 6.764 20.88 9.236 20.912 ;
  LAYER M2 ;
        RECT 6.764 20.944 9.236 20.976 ;
  LAYER M2 ;
        RECT 6.764 21.008 9.236 21.04 ;
  LAYER M2 ;
        RECT 6.764 21.072 9.236 21.104 ;
  LAYER M2 ;
        RECT 6.764 21.136 9.236 21.168 ;
  LAYER M2 ;
        RECT 6.764 21.2 9.236 21.232 ;
  LAYER M2 ;
        RECT 6.764 21.264 9.236 21.296 ;
  LAYER M2 ;
        RECT 6.764 21.328 9.236 21.36 ;
  LAYER M2 ;
        RECT 6.764 21.392 9.236 21.424 ;
  LAYER M2 ;
        RECT 6.764 21.456 9.236 21.488 ;
  LAYER M2 ;
        RECT 6.764 21.52 9.236 21.552 ;
  LAYER M2 ;
        RECT 6.764 21.584 9.236 21.616 ;
  LAYER M2 ;
        RECT 6.764 21.648 9.236 21.68 ;
  LAYER M2 ;
        RECT 6.764 21.712 9.236 21.744 ;
  LAYER M2 ;
        RECT 6.764 21.776 9.236 21.808 ;
  LAYER M2 ;
        RECT 6.764 21.84 9.236 21.872 ;
  LAYER M2 ;
        RECT 6.764 21.904 9.236 21.936 ;
  LAYER M2 ;
        RECT 6.764 21.968 9.236 22 ;
  LAYER M2 ;
        RECT 6.764 22.032 9.236 22.064 ;
  LAYER M2 ;
        RECT 6.764 22.096 9.236 22.128 ;
  LAYER M2 ;
        RECT 6.764 22.16 9.236 22.192 ;
  LAYER M2 ;
        RECT 6.764 22.224 9.236 22.256 ;
  LAYER M2 ;
        RECT 6.764 22.288 9.236 22.32 ;
  LAYER M2 ;
        RECT 6.764 22.352 9.236 22.384 ;
  LAYER M2 ;
        RECT 6.764 22.416 9.236 22.448 ;
  LAYER M2 ;
        RECT 6.764 22.48 9.236 22.512 ;
  LAYER M2 ;
        RECT 6.764 22.544 9.236 22.576 ;
  LAYER M2 ;
        RECT 6.764 22.608 9.236 22.64 ;
  LAYER M2 ;
        RECT 6.764 22.672 9.236 22.704 ;
  LAYER M2 ;
        RECT 6.764 22.736 9.236 22.768 ;
  LAYER M2 ;
        RECT 6.764 22.8 9.236 22.832 ;
  LAYER M2 ;
        RECT 6.764 22.864 9.236 22.896 ;
  LAYER M2 ;
        RECT 6.764 22.928 9.236 22.96 ;
  LAYER M2 ;
        RECT 6.764 22.992 9.236 23.024 ;
  LAYER M2 ;
        RECT 6.764 23.056 9.236 23.088 ;
  LAYER M2 ;
        RECT 6.764 23.12 9.236 23.152 ;
  LAYER M3 ;
        RECT 9.184 20.796 9.216 23.304 ;
  LAYER M3 ;
        RECT 9.12 20.796 9.152 23.304 ;
  LAYER M3 ;
        RECT 9.056 20.796 9.088 23.304 ;
  LAYER M3 ;
        RECT 8.992 20.796 9.024 23.304 ;
  LAYER M3 ;
        RECT 8.928 20.796 8.96 23.304 ;
  LAYER M3 ;
        RECT 8.864 20.796 8.896 23.304 ;
  LAYER M3 ;
        RECT 8.8 20.796 8.832 23.304 ;
  LAYER M3 ;
        RECT 8.736 20.796 8.768 23.304 ;
  LAYER M3 ;
        RECT 8.672 20.796 8.704 23.304 ;
  LAYER M3 ;
        RECT 8.608 20.796 8.64 23.304 ;
  LAYER M3 ;
        RECT 8.544 20.796 8.576 23.304 ;
  LAYER M3 ;
        RECT 8.48 20.796 8.512 23.304 ;
  LAYER M3 ;
        RECT 8.416 20.796 8.448 23.304 ;
  LAYER M3 ;
        RECT 8.352 20.796 8.384 23.304 ;
  LAYER M3 ;
        RECT 8.288 20.796 8.32 23.304 ;
  LAYER M3 ;
        RECT 8.224 20.796 8.256 23.304 ;
  LAYER M3 ;
        RECT 8.16 20.796 8.192 23.304 ;
  LAYER M3 ;
        RECT 8.096 20.796 8.128 23.304 ;
  LAYER M3 ;
        RECT 8.032 20.796 8.064 23.304 ;
  LAYER M3 ;
        RECT 7.968 20.796 8 23.304 ;
  LAYER M3 ;
        RECT 7.904 20.796 7.936 23.304 ;
  LAYER M3 ;
        RECT 7.84 20.796 7.872 23.304 ;
  LAYER M3 ;
        RECT 7.776 20.796 7.808 23.304 ;
  LAYER M3 ;
        RECT 7.712 20.796 7.744 23.304 ;
  LAYER M3 ;
        RECT 7.648 20.796 7.68 23.304 ;
  LAYER M3 ;
        RECT 7.584 20.796 7.616 23.304 ;
  LAYER M3 ;
        RECT 7.52 20.796 7.552 23.304 ;
  LAYER M3 ;
        RECT 7.456 20.796 7.488 23.304 ;
  LAYER M3 ;
        RECT 7.392 20.796 7.424 23.304 ;
  LAYER M3 ;
        RECT 7.328 20.796 7.36 23.304 ;
  LAYER M3 ;
        RECT 7.264 20.796 7.296 23.304 ;
  LAYER M3 ;
        RECT 7.2 20.796 7.232 23.304 ;
  LAYER M3 ;
        RECT 7.136 20.796 7.168 23.304 ;
  LAYER M3 ;
        RECT 7.072 20.796 7.104 23.304 ;
  LAYER M3 ;
        RECT 7.008 20.796 7.04 23.304 ;
  LAYER M3 ;
        RECT 6.944 20.796 6.976 23.304 ;
  LAYER M3 ;
        RECT 6.88 20.796 6.912 23.304 ;
  LAYER M3 ;
        RECT 6.784 20.796 6.816 23.304 ;
  LAYER M1 ;
        RECT 9.199 20.832 9.201 23.268 ;
  LAYER M1 ;
        RECT 9.119 20.832 9.121 23.268 ;
  LAYER M1 ;
        RECT 9.039 20.832 9.041 23.268 ;
  LAYER M1 ;
        RECT 8.959 20.832 8.961 23.268 ;
  LAYER M1 ;
        RECT 8.879 20.832 8.881 23.268 ;
  LAYER M1 ;
        RECT 8.799 20.832 8.801 23.268 ;
  LAYER M1 ;
        RECT 8.719 20.832 8.721 23.268 ;
  LAYER M1 ;
        RECT 8.639 20.832 8.641 23.268 ;
  LAYER M1 ;
        RECT 8.559 20.832 8.561 23.268 ;
  LAYER M1 ;
        RECT 8.479 20.832 8.481 23.268 ;
  LAYER M1 ;
        RECT 8.399 20.832 8.401 23.268 ;
  LAYER M1 ;
        RECT 8.319 20.832 8.321 23.268 ;
  LAYER M1 ;
        RECT 8.239 20.832 8.241 23.268 ;
  LAYER M1 ;
        RECT 8.159 20.832 8.161 23.268 ;
  LAYER M1 ;
        RECT 8.079 20.832 8.081 23.268 ;
  LAYER M1 ;
        RECT 7.999 20.832 8.001 23.268 ;
  LAYER M1 ;
        RECT 7.919 20.832 7.921 23.268 ;
  LAYER M1 ;
        RECT 7.839 20.832 7.841 23.268 ;
  LAYER M1 ;
        RECT 7.759 20.832 7.761 23.268 ;
  LAYER M1 ;
        RECT 7.679 20.832 7.681 23.268 ;
  LAYER M1 ;
        RECT 7.599 20.832 7.601 23.268 ;
  LAYER M1 ;
        RECT 7.519 20.832 7.521 23.268 ;
  LAYER M1 ;
        RECT 7.439 20.832 7.441 23.268 ;
  LAYER M1 ;
        RECT 7.359 20.832 7.361 23.268 ;
  LAYER M1 ;
        RECT 7.279 20.832 7.281 23.268 ;
  LAYER M1 ;
        RECT 7.199 20.832 7.201 23.268 ;
  LAYER M1 ;
        RECT 7.119 20.832 7.121 23.268 ;
  LAYER M1 ;
        RECT 7.039 20.832 7.041 23.268 ;
  LAYER M1 ;
        RECT 6.959 20.832 6.961 23.268 ;
  LAYER M1 ;
        RECT 6.879 20.832 6.881 23.268 ;
  LAYER M2 ;
        RECT 6.8 20.831 9.2 20.833 ;
  LAYER M2 ;
        RECT 6.8 20.915 9.2 20.917 ;
  LAYER M2 ;
        RECT 6.8 20.999 9.2 21.001 ;
  LAYER M2 ;
        RECT 6.8 21.083 9.2 21.085 ;
  LAYER M2 ;
        RECT 6.8 21.167 9.2 21.169 ;
  LAYER M2 ;
        RECT 6.8 21.251 9.2 21.253 ;
  LAYER M2 ;
        RECT 6.8 21.335 9.2 21.337 ;
  LAYER M2 ;
        RECT 6.8 21.419 9.2 21.421 ;
  LAYER M2 ;
        RECT 6.8 21.503 9.2 21.505 ;
  LAYER M2 ;
        RECT 6.8 21.587 9.2 21.589 ;
  LAYER M2 ;
        RECT 6.8 21.671 9.2 21.673 ;
  LAYER M2 ;
        RECT 6.8 21.755 9.2 21.757 ;
  LAYER M2 ;
        RECT 6.8 21.8385 9.2 21.8405 ;
  LAYER M2 ;
        RECT 6.8 21.923 9.2 21.925 ;
  LAYER M2 ;
        RECT 6.8 22.007 9.2 22.009 ;
  LAYER M2 ;
        RECT 6.8 22.091 9.2 22.093 ;
  LAYER M2 ;
        RECT 6.8 22.175 9.2 22.177 ;
  LAYER M2 ;
        RECT 6.8 22.259 9.2 22.261 ;
  LAYER M2 ;
        RECT 6.8 22.343 9.2 22.345 ;
  LAYER M2 ;
        RECT 6.8 22.427 9.2 22.429 ;
  LAYER M2 ;
        RECT 6.8 22.511 9.2 22.513 ;
  LAYER M2 ;
        RECT 6.8 22.595 9.2 22.597 ;
  LAYER M2 ;
        RECT 6.8 22.679 9.2 22.681 ;
  LAYER M2 ;
        RECT 6.8 22.763 9.2 22.765 ;
  LAYER M2 ;
        RECT 6.8 22.847 9.2 22.849 ;
  LAYER M2 ;
        RECT 6.8 22.931 9.2 22.933 ;
  LAYER M2 ;
        RECT 6.8 23.015 9.2 23.017 ;
  LAYER M2 ;
        RECT 6.8 23.099 9.2 23.101 ;
  LAYER M2 ;
        RECT 6.8 23.183 9.2 23.185 ;
  LAYER M1 ;
        RECT 9.184 23.736 9.216 26.244 ;
  LAYER M1 ;
        RECT 9.12 23.736 9.152 26.244 ;
  LAYER M1 ;
        RECT 9.056 23.736 9.088 26.244 ;
  LAYER M1 ;
        RECT 8.992 23.736 9.024 26.244 ;
  LAYER M1 ;
        RECT 8.928 23.736 8.96 26.244 ;
  LAYER M1 ;
        RECT 8.864 23.736 8.896 26.244 ;
  LAYER M1 ;
        RECT 8.8 23.736 8.832 26.244 ;
  LAYER M1 ;
        RECT 8.736 23.736 8.768 26.244 ;
  LAYER M1 ;
        RECT 8.672 23.736 8.704 26.244 ;
  LAYER M1 ;
        RECT 8.608 23.736 8.64 26.244 ;
  LAYER M1 ;
        RECT 8.544 23.736 8.576 26.244 ;
  LAYER M1 ;
        RECT 8.48 23.736 8.512 26.244 ;
  LAYER M1 ;
        RECT 8.416 23.736 8.448 26.244 ;
  LAYER M1 ;
        RECT 8.352 23.736 8.384 26.244 ;
  LAYER M1 ;
        RECT 8.288 23.736 8.32 26.244 ;
  LAYER M1 ;
        RECT 8.224 23.736 8.256 26.244 ;
  LAYER M1 ;
        RECT 8.16 23.736 8.192 26.244 ;
  LAYER M1 ;
        RECT 8.096 23.736 8.128 26.244 ;
  LAYER M1 ;
        RECT 8.032 23.736 8.064 26.244 ;
  LAYER M1 ;
        RECT 7.968 23.736 8 26.244 ;
  LAYER M1 ;
        RECT 7.904 23.736 7.936 26.244 ;
  LAYER M1 ;
        RECT 7.84 23.736 7.872 26.244 ;
  LAYER M1 ;
        RECT 7.776 23.736 7.808 26.244 ;
  LAYER M1 ;
        RECT 7.712 23.736 7.744 26.244 ;
  LAYER M1 ;
        RECT 7.648 23.736 7.68 26.244 ;
  LAYER M1 ;
        RECT 7.584 23.736 7.616 26.244 ;
  LAYER M1 ;
        RECT 7.52 23.736 7.552 26.244 ;
  LAYER M1 ;
        RECT 7.456 23.736 7.488 26.244 ;
  LAYER M1 ;
        RECT 7.392 23.736 7.424 26.244 ;
  LAYER M1 ;
        RECT 7.328 23.736 7.36 26.244 ;
  LAYER M1 ;
        RECT 7.264 23.736 7.296 26.244 ;
  LAYER M1 ;
        RECT 7.2 23.736 7.232 26.244 ;
  LAYER M1 ;
        RECT 7.136 23.736 7.168 26.244 ;
  LAYER M1 ;
        RECT 7.072 23.736 7.104 26.244 ;
  LAYER M1 ;
        RECT 7.008 23.736 7.04 26.244 ;
  LAYER M1 ;
        RECT 6.944 23.736 6.976 26.244 ;
  LAYER M1 ;
        RECT 6.88 23.736 6.912 26.244 ;
  LAYER M2 ;
        RECT 6.764 23.82 9.236 23.852 ;
  LAYER M2 ;
        RECT 6.764 23.884 9.236 23.916 ;
  LAYER M2 ;
        RECT 6.764 23.948 9.236 23.98 ;
  LAYER M2 ;
        RECT 6.764 24.012 9.236 24.044 ;
  LAYER M2 ;
        RECT 6.764 24.076 9.236 24.108 ;
  LAYER M2 ;
        RECT 6.764 24.14 9.236 24.172 ;
  LAYER M2 ;
        RECT 6.764 24.204 9.236 24.236 ;
  LAYER M2 ;
        RECT 6.764 24.268 9.236 24.3 ;
  LAYER M2 ;
        RECT 6.764 24.332 9.236 24.364 ;
  LAYER M2 ;
        RECT 6.764 24.396 9.236 24.428 ;
  LAYER M2 ;
        RECT 6.764 24.46 9.236 24.492 ;
  LAYER M2 ;
        RECT 6.764 24.524 9.236 24.556 ;
  LAYER M2 ;
        RECT 6.764 24.588 9.236 24.62 ;
  LAYER M2 ;
        RECT 6.764 24.652 9.236 24.684 ;
  LAYER M2 ;
        RECT 6.764 24.716 9.236 24.748 ;
  LAYER M2 ;
        RECT 6.764 24.78 9.236 24.812 ;
  LAYER M2 ;
        RECT 6.764 24.844 9.236 24.876 ;
  LAYER M2 ;
        RECT 6.764 24.908 9.236 24.94 ;
  LAYER M2 ;
        RECT 6.764 24.972 9.236 25.004 ;
  LAYER M2 ;
        RECT 6.764 25.036 9.236 25.068 ;
  LAYER M2 ;
        RECT 6.764 25.1 9.236 25.132 ;
  LAYER M2 ;
        RECT 6.764 25.164 9.236 25.196 ;
  LAYER M2 ;
        RECT 6.764 25.228 9.236 25.26 ;
  LAYER M2 ;
        RECT 6.764 25.292 9.236 25.324 ;
  LAYER M2 ;
        RECT 6.764 25.356 9.236 25.388 ;
  LAYER M2 ;
        RECT 6.764 25.42 9.236 25.452 ;
  LAYER M2 ;
        RECT 6.764 25.484 9.236 25.516 ;
  LAYER M2 ;
        RECT 6.764 25.548 9.236 25.58 ;
  LAYER M2 ;
        RECT 6.764 25.612 9.236 25.644 ;
  LAYER M2 ;
        RECT 6.764 25.676 9.236 25.708 ;
  LAYER M2 ;
        RECT 6.764 25.74 9.236 25.772 ;
  LAYER M2 ;
        RECT 6.764 25.804 9.236 25.836 ;
  LAYER M2 ;
        RECT 6.764 25.868 9.236 25.9 ;
  LAYER M2 ;
        RECT 6.764 25.932 9.236 25.964 ;
  LAYER M2 ;
        RECT 6.764 25.996 9.236 26.028 ;
  LAYER M2 ;
        RECT 6.764 26.06 9.236 26.092 ;
  LAYER M3 ;
        RECT 9.184 23.736 9.216 26.244 ;
  LAYER M3 ;
        RECT 9.12 23.736 9.152 26.244 ;
  LAYER M3 ;
        RECT 9.056 23.736 9.088 26.244 ;
  LAYER M3 ;
        RECT 8.992 23.736 9.024 26.244 ;
  LAYER M3 ;
        RECT 8.928 23.736 8.96 26.244 ;
  LAYER M3 ;
        RECT 8.864 23.736 8.896 26.244 ;
  LAYER M3 ;
        RECT 8.8 23.736 8.832 26.244 ;
  LAYER M3 ;
        RECT 8.736 23.736 8.768 26.244 ;
  LAYER M3 ;
        RECT 8.672 23.736 8.704 26.244 ;
  LAYER M3 ;
        RECT 8.608 23.736 8.64 26.244 ;
  LAYER M3 ;
        RECT 8.544 23.736 8.576 26.244 ;
  LAYER M3 ;
        RECT 8.48 23.736 8.512 26.244 ;
  LAYER M3 ;
        RECT 8.416 23.736 8.448 26.244 ;
  LAYER M3 ;
        RECT 8.352 23.736 8.384 26.244 ;
  LAYER M3 ;
        RECT 8.288 23.736 8.32 26.244 ;
  LAYER M3 ;
        RECT 8.224 23.736 8.256 26.244 ;
  LAYER M3 ;
        RECT 8.16 23.736 8.192 26.244 ;
  LAYER M3 ;
        RECT 8.096 23.736 8.128 26.244 ;
  LAYER M3 ;
        RECT 8.032 23.736 8.064 26.244 ;
  LAYER M3 ;
        RECT 7.968 23.736 8 26.244 ;
  LAYER M3 ;
        RECT 7.904 23.736 7.936 26.244 ;
  LAYER M3 ;
        RECT 7.84 23.736 7.872 26.244 ;
  LAYER M3 ;
        RECT 7.776 23.736 7.808 26.244 ;
  LAYER M3 ;
        RECT 7.712 23.736 7.744 26.244 ;
  LAYER M3 ;
        RECT 7.648 23.736 7.68 26.244 ;
  LAYER M3 ;
        RECT 7.584 23.736 7.616 26.244 ;
  LAYER M3 ;
        RECT 7.52 23.736 7.552 26.244 ;
  LAYER M3 ;
        RECT 7.456 23.736 7.488 26.244 ;
  LAYER M3 ;
        RECT 7.392 23.736 7.424 26.244 ;
  LAYER M3 ;
        RECT 7.328 23.736 7.36 26.244 ;
  LAYER M3 ;
        RECT 7.264 23.736 7.296 26.244 ;
  LAYER M3 ;
        RECT 7.2 23.736 7.232 26.244 ;
  LAYER M3 ;
        RECT 7.136 23.736 7.168 26.244 ;
  LAYER M3 ;
        RECT 7.072 23.736 7.104 26.244 ;
  LAYER M3 ;
        RECT 7.008 23.736 7.04 26.244 ;
  LAYER M3 ;
        RECT 6.944 23.736 6.976 26.244 ;
  LAYER M3 ;
        RECT 6.88 23.736 6.912 26.244 ;
  LAYER M3 ;
        RECT 6.784 23.736 6.816 26.244 ;
  LAYER M1 ;
        RECT 9.199 23.772 9.201 26.208 ;
  LAYER M1 ;
        RECT 9.119 23.772 9.121 26.208 ;
  LAYER M1 ;
        RECT 9.039 23.772 9.041 26.208 ;
  LAYER M1 ;
        RECT 8.959 23.772 8.961 26.208 ;
  LAYER M1 ;
        RECT 8.879 23.772 8.881 26.208 ;
  LAYER M1 ;
        RECT 8.799 23.772 8.801 26.208 ;
  LAYER M1 ;
        RECT 8.719 23.772 8.721 26.208 ;
  LAYER M1 ;
        RECT 8.639 23.772 8.641 26.208 ;
  LAYER M1 ;
        RECT 8.559 23.772 8.561 26.208 ;
  LAYER M1 ;
        RECT 8.479 23.772 8.481 26.208 ;
  LAYER M1 ;
        RECT 8.399 23.772 8.401 26.208 ;
  LAYER M1 ;
        RECT 8.319 23.772 8.321 26.208 ;
  LAYER M1 ;
        RECT 8.239 23.772 8.241 26.208 ;
  LAYER M1 ;
        RECT 8.159 23.772 8.161 26.208 ;
  LAYER M1 ;
        RECT 8.079 23.772 8.081 26.208 ;
  LAYER M1 ;
        RECT 7.999 23.772 8.001 26.208 ;
  LAYER M1 ;
        RECT 7.919 23.772 7.921 26.208 ;
  LAYER M1 ;
        RECT 7.839 23.772 7.841 26.208 ;
  LAYER M1 ;
        RECT 7.759 23.772 7.761 26.208 ;
  LAYER M1 ;
        RECT 7.679 23.772 7.681 26.208 ;
  LAYER M1 ;
        RECT 7.599 23.772 7.601 26.208 ;
  LAYER M1 ;
        RECT 7.519 23.772 7.521 26.208 ;
  LAYER M1 ;
        RECT 7.439 23.772 7.441 26.208 ;
  LAYER M1 ;
        RECT 7.359 23.772 7.361 26.208 ;
  LAYER M1 ;
        RECT 7.279 23.772 7.281 26.208 ;
  LAYER M1 ;
        RECT 7.199 23.772 7.201 26.208 ;
  LAYER M1 ;
        RECT 7.119 23.772 7.121 26.208 ;
  LAYER M1 ;
        RECT 7.039 23.772 7.041 26.208 ;
  LAYER M1 ;
        RECT 6.959 23.772 6.961 26.208 ;
  LAYER M1 ;
        RECT 6.879 23.772 6.881 26.208 ;
  LAYER M2 ;
        RECT 6.8 23.771 9.2 23.773 ;
  LAYER M2 ;
        RECT 6.8 23.855 9.2 23.857 ;
  LAYER M2 ;
        RECT 6.8 23.939 9.2 23.941 ;
  LAYER M2 ;
        RECT 6.8 24.023 9.2 24.025 ;
  LAYER M2 ;
        RECT 6.8 24.107 9.2 24.109 ;
  LAYER M2 ;
        RECT 6.8 24.191 9.2 24.193 ;
  LAYER M2 ;
        RECT 6.8 24.275 9.2 24.277 ;
  LAYER M2 ;
        RECT 6.8 24.359 9.2 24.361 ;
  LAYER M2 ;
        RECT 6.8 24.443 9.2 24.445 ;
  LAYER M2 ;
        RECT 6.8 24.527 9.2 24.529 ;
  LAYER M2 ;
        RECT 6.8 24.611 9.2 24.613 ;
  LAYER M2 ;
        RECT 6.8 24.695 9.2 24.697 ;
  LAYER M2 ;
        RECT 6.8 24.7785 9.2 24.7805 ;
  LAYER M2 ;
        RECT 6.8 24.863 9.2 24.865 ;
  LAYER M2 ;
        RECT 6.8 24.947 9.2 24.949 ;
  LAYER M2 ;
        RECT 6.8 25.031 9.2 25.033 ;
  LAYER M2 ;
        RECT 6.8 25.115 9.2 25.117 ;
  LAYER M2 ;
        RECT 6.8 25.199 9.2 25.201 ;
  LAYER M2 ;
        RECT 6.8 25.283 9.2 25.285 ;
  LAYER M2 ;
        RECT 6.8 25.367 9.2 25.369 ;
  LAYER M2 ;
        RECT 6.8 25.451 9.2 25.453 ;
  LAYER M2 ;
        RECT 6.8 25.535 9.2 25.537 ;
  LAYER M2 ;
        RECT 6.8 25.619 9.2 25.621 ;
  LAYER M2 ;
        RECT 6.8 25.703 9.2 25.705 ;
  LAYER M2 ;
        RECT 6.8 25.787 9.2 25.789 ;
  LAYER M2 ;
        RECT 6.8 25.871 9.2 25.873 ;
  LAYER M2 ;
        RECT 6.8 25.955 9.2 25.957 ;
  LAYER M2 ;
        RECT 6.8 26.039 9.2 26.041 ;
  LAYER M2 ;
        RECT 6.8 26.123 9.2 26.125 ;
  LAYER M1 ;
        RECT 9.184 26.676 9.216 29.184 ;
  LAYER M1 ;
        RECT 9.12 26.676 9.152 29.184 ;
  LAYER M1 ;
        RECT 9.056 26.676 9.088 29.184 ;
  LAYER M1 ;
        RECT 8.992 26.676 9.024 29.184 ;
  LAYER M1 ;
        RECT 8.928 26.676 8.96 29.184 ;
  LAYER M1 ;
        RECT 8.864 26.676 8.896 29.184 ;
  LAYER M1 ;
        RECT 8.8 26.676 8.832 29.184 ;
  LAYER M1 ;
        RECT 8.736 26.676 8.768 29.184 ;
  LAYER M1 ;
        RECT 8.672 26.676 8.704 29.184 ;
  LAYER M1 ;
        RECT 8.608 26.676 8.64 29.184 ;
  LAYER M1 ;
        RECT 8.544 26.676 8.576 29.184 ;
  LAYER M1 ;
        RECT 8.48 26.676 8.512 29.184 ;
  LAYER M1 ;
        RECT 8.416 26.676 8.448 29.184 ;
  LAYER M1 ;
        RECT 8.352 26.676 8.384 29.184 ;
  LAYER M1 ;
        RECT 8.288 26.676 8.32 29.184 ;
  LAYER M1 ;
        RECT 8.224 26.676 8.256 29.184 ;
  LAYER M1 ;
        RECT 8.16 26.676 8.192 29.184 ;
  LAYER M1 ;
        RECT 8.096 26.676 8.128 29.184 ;
  LAYER M1 ;
        RECT 8.032 26.676 8.064 29.184 ;
  LAYER M1 ;
        RECT 7.968 26.676 8 29.184 ;
  LAYER M1 ;
        RECT 7.904 26.676 7.936 29.184 ;
  LAYER M1 ;
        RECT 7.84 26.676 7.872 29.184 ;
  LAYER M1 ;
        RECT 7.776 26.676 7.808 29.184 ;
  LAYER M1 ;
        RECT 7.712 26.676 7.744 29.184 ;
  LAYER M1 ;
        RECT 7.648 26.676 7.68 29.184 ;
  LAYER M1 ;
        RECT 7.584 26.676 7.616 29.184 ;
  LAYER M1 ;
        RECT 7.52 26.676 7.552 29.184 ;
  LAYER M1 ;
        RECT 7.456 26.676 7.488 29.184 ;
  LAYER M1 ;
        RECT 7.392 26.676 7.424 29.184 ;
  LAYER M1 ;
        RECT 7.328 26.676 7.36 29.184 ;
  LAYER M1 ;
        RECT 7.264 26.676 7.296 29.184 ;
  LAYER M1 ;
        RECT 7.2 26.676 7.232 29.184 ;
  LAYER M1 ;
        RECT 7.136 26.676 7.168 29.184 ;
  LAYER M1 ;
        RECT 7.072 26.676 7.104 29.184 ;
  LAYER M1 ;
        RECT 7.008 26.676 7.04 29.184 ;
  LAYER M1 ;
        RECT 6.944 26.676 6.976 29.184 ;
  LAYER M1 ;
        RECT 6.88 26.676 6.912 29.184 ;
  LAYER M2 ;
        RECT 6.764 26.76 9.236 26.792 ;
  LAYER M2 ;
        RECT 6.764 26.824 9.236 26.856 ;
  LAYER M2 ;
        RECT 6.764 26.888 9.236 26.92 ;
  LAYER M2 ;
        RECT 6.764 26.952 9.236 26.984 ;
  LAYER M2 ;
        RECT 6.764 27.016 9.236 27.048 ;
  LAYER M2 ;
        RECT 6.764 27.08 9.236 27.112 ;
  LAYER M2 ;
        RECT 6.764 27.144 9.236 27.176 ;
  LAYER M2 ;
        RECT 6.764 27.208 9.236 27.24 ;
  LAYER M2 ;
        RECT 6.764 27.272 9.236 27.304 ;
  LAYER M2 ;
        RECT 6.764 27.336 9.236 27.368 ;
  LAYER M2 ;
        RECT 6.764 27.4 9.236 27.432 ;
  LAYER M2 ;
        RECT 6.764 27.464 9.236 27.496 ;
  LAYER M2 ;
        RECT 6.764 27.528 9.236 27.56 ;
  LAYER M2 ;
        RECT 6.764 27.592 9.236 27.624 ;
  LAYER M2 ;
        RECT 6.764 27.656 9.236 27.688 ;
  LAYER M2 ;
        RECT 6.764 27.72 9.236 27.752 ;
  LAYER M2 ;
        RECT 6.764 27.784 9.236 27.816 ;
  LAYER M2 ;
        RECT 6.764 27.848 9.236 27.88 ;
  LAYER M2 ;
        RECT 6.764 27.912 9.236 27.944 ;
  LAYER M2 ;
        RECT 6.764 27.976 9.236 28.008 ;
  LAYER M2 ;
        RECT 6.764 28.04 9.236 28.072 ;
  LAYER M2 ;
        RECT 6.764 28.104 9.236 28.136 ;
  LAYER M2 ;
        RECT 6.764 28.168 9.236 28.2 ;
  LAYER M2 ;
        RECT 6.764 28.232 9.236 28.264 ;
  LAYER M2 ;
        RECT 6.764 28.296 9.236 28.328 ;
  LAYER M2 ;
        RECT 6.764 28.36 9.236 28.392 ;
  LAYER M2 ;
        RECT 6.764 28.424 9.236 28.456 ;
  LAYER M2 ;
        RECT 6.764 28.488 9.236 28.52 ;
  LAYER M2 ;
        RECT 6.764 28.552 9.236 28.584 ;
  LAYER M2 ;
        RECT 6.764 28.616 9.236 28.648 ;
  LAYER M2 ;
        RECT 6.764 28.68 9.236 28.712 ;
  LAYER M2 ;
        RECT 6.764 28.744 9.236 28.776 ;
  LAYER M2 ;
        RECT 6.764 28.808 9.236 28.84 ;
  LAYER M2 ;
        RECT 6.764 28.872 9.236 28.904 ;
  LAYER M2 ;
        RECT 6.764 28.936 9.236 28.968 ;
  LAYER M2 ;
        RECT 6.764 29 9.236 29.032 ;
  LAYER M3 ;
        RECT 9.184 26.676 9.216 29.184 ;
  LAYER M3 ;
        RECT 9.12 26.676 9.152 29.184 ;
  LAYER M3 ;
        RECT 9.056 26.676 9.088 29.184 ;
  LAYER M3 ;
        RECT 8.992 26.676 9.024 29.184 ;
  LAYER M3 ;
        RECT 8.928 26.676 8.96 29.184 ;
  LAYER M3 ;
        RECT 8.864 26.676 8.896 29.184 ;
  LAYER M3 ;
        RECT 8.8 26.676 8.832 29.184 ;
  LAYER M3 ;
        RECT 8.736 26.676 8.768 29.184 ;
  LAYER M3 ;
        RECT 8.672 26.676 8.704 29.184 ;
  LAYER M3 ;
        RECT 8.608 26.676 8.64 29.184 ;
  LAYER M3 ;
        RECT 8.544 26.676 8.576 29.184 ;
  LAYER M3 ;
        RECT 8.48 26.676 8.512 29.184 ;
  LAYER M3 ;
        RECT 8.416 26.676 8.448 29.184 ;
  LAYER M3 ;
        RECT 8.352 26.676 8.384 29.184 ;
  LAYER M3 ;
        RECT 8.288 26.676 8.32 29.184 ;
  LAYER M3 ;
        RECT 8.224 26.676 8.256 29.184 ;
  LAYER M3 ;
        RECT 8.16 26.676 8.192 29.184 ;
  LAYER M3 ;
        RECT 8.096 26.676 8.128 29.184 ;
  LAYER M3 ;
        RECT 8.032 26.676 8.064 29.184 ;
  LAYER M3 ;
        RECT 7.968 26.676 8 29.184 ;
  LAYER M3 ;
        RECT 7.904 26.676 7.936 29.184 ;
  LAYER M3 ;
        RECT 7.84 26.676 7.872 29.184 ;
  LAYER M3 ;
        RECT 7.776 26.676 7.808 29.184 ;
  LAYER M3 ;
        RECT 7.712 26.676 7.744 29.184 ;
  LAYER M3 ;
        RECT 7.648 26.676 7.68 29.184 ;
  LAYER M3 ;
        RECT 7.584 26.676 7.616 29.184 ;
  LAYER M3 ;
        RECT 7.52 26.676 7.552 29.184 ;
  LAYER M3 ;
        RECT 7.456 26.676 7.488 29.184 ;
  LAYER M3 ;
        RECT 7.392 26.676 7.424 29.184 ;
  LAYER M3 ;
        RECT 7.328 26.676 7.36 29.184 ;
  LAYER M3 ;
        RECT 7.264 26.676 7.296 29.184 ;
  LAYER M3 ;
        RECT 7.2 26.676 7.232 29.184 ;
  LAYER M3 ;
        RECT 7.136 26.676 7.168 29.184 ;
  LAYER M3 ;
        RECT 7.072 26.676 7.104 29.184 ;
  LAYER M3 ;
        RECT 7.008 26.676 7.04 29.184 ;
  LAYER M3 ;
        RECT 6.944 26.676 6.976 29.184 ;
  LAYER M3 ;
        RECT 6.88 26.676 6.912 29.184 ;
  LAYER M3 ;
        RECT 6.784 26.676 6.816 29.184 ;
  LAYER M1 ;
        RECT 9.199 26.712 9.201 29.148 ;
  LAYER M1 ;
        RECT 9.119 26.712 9.121 29.148 ;
  LAYER M1 ;
        RECT 9.039 26.712 9.041 29.148 ;
  LAYER M1 ;
        RECT 8.959 26.712 8.961 29.148 ;
  LAYER M1 ;
        RECT 8.879 26.712 8.881 29.148 ;
  LAYER M1 ;
        RECT 8.799 26.712 8.801 29.148 ;
  LAYER M1 ;
        RECT 8.719 26.712 8.721 29.148 ;
  LAYER M1 ;
        RECT 8.639 26.712 8.641 29.148 ;
  LAYER M1 ;
        RECT 8.559 26.712 8.561 29.148 ;
  LAYER M1 ;
        RECT 8.479 26.712 8.481 29.148 ;
  LAYER M1 ;
        RECT 8.399 26.712 8.401 29.148 ;
  LAYER M1 ;
        RECT 8.319 26.712 8.321 29.148 ;
  LAYER M1 ;
        RECT 8.239 26.712 8.241 29.148 ;
  LAYER M1 ;
        RECT 8.159 26.712 8.161 29.148 ;
  LAYER M1 ;
        RECT 8.079 26.712 8.081 29.148 ;
  LAYER M1 ;
        RECT 7.999 26.712 8.001 29.148 ;
  LAYER M1 ;
        RECT 7.919 26.712 7.921 29.148 ;
  LAYER M1 ;
        RECT 7.839 26.712 7.841 29.148 ;
  LAYER M1 ;
        RECT 7.759 26.712 7.761 29.148 ;
  LAYER M1 ;
        RECT 7.679 26.712 7.681 29.148 ;
  LAYER M1 ;
        RECT 7.599 26.712 7.601 29.148 ;
  LAYER M1 ;
        RECT 7.519 26.712 7.521 29.148 ;
  LAYER M1 ;
        RECT 7.439 26.712 7.441 29.148 ;
  LAYER M1 ;
        RECT 7.359 26.712 7.361 29.148 ;
  LAYER M1 ;
        RECT 7.279 26.712 7.281 29.148 ;
  LAYER M1 ;
        RECT 7.199 26.712 7.201 29.148 ;
  LAYER M1 ;
        RECT 7.119 26.712 7.121 29.148 ;
  LAYER M1 ;
        RECT 7.039 26.712 7.041 29.148 ;
  LAYER M1 ;
        RECT 6.959 26.712 6.961 29.148 ;
  LAYER M1 ;
        RECT 6.879 26.712 6.881 29.148 ;
  LAYER M2 ;
        RECT 6.8 26.711 9.2 26.713 ;
  LAYER M2 ;
        RECT 6.8 26.795 9.2 26.797 ;
  LAYER M2 ;
        RECT 6.8 26.879 9.2 26.881 ;
  LAYER M2 ;
        RECT 6.8 26.963 9.2 26.965 ;
  LAYER M2 ;
        RECT 6.8 27.047 9.2 27.049 ;
  LAYER M2 ;
        RECT 6.8 27.131 9.2 27.133 ;
  LAYER M2 ;
        RECT 6.8 27.215 9.2 27.217 ;
  LAYER M2 ;
        RECT 6.8 27.299 9.2 27.301 ;
  LAYER M2 ;
        RECT 6.8 27.383 9.2 27.385 ;
  LAYER M2 ;
        RECT 6.8 27.467 9.2 27.469 ;
  LAYER M2 ;
        RECT 6.8 27.551 9.2 27.553 ;
  LAYER M2 ;
        RECT 6.8 27.635 9.2 27.637 ;
  LAYER M2 ;
        RECT 6.8 27.7185 9.2 27.7205 ;
  LAYER M2 ;
        RECT 6.8 27.803 9.2 27.805 ;
  LAYER M2 ;
        RECT 6.8 27.887 9.2 27.889 ;
  LAYER M2 ;
        RECT 6.8 27.971 9.2 27.973 ;
  LAYER M2 ;
        RECT 6.8 28.055 9.2 28.057 ;
  LAYER M2 ;
        RECT 6.8 28.139 9.2 28.141 ;
  LAYER M2 ;
        RECT 6.8 28.223 9.2 28.225 ;
  LAYER M2 ;
        RECT 6.8 28.307 9.2 28.309 ;
  LAYER M2 ;
        RECT 6.8 28.391 9.2 28.393 ;
  LAYER M2 ;
        RECT 6.8 28.475 9.2 28.477 ;
  LAYER M2 ;
        RECT 6.8 28.559 9.2 28.561 ;
  LAYER M2 ;
        RECT 6.8 28.643 9.2 28.645 ;
  LAYER M2 ;
        RECT 6.8 28.727 9.2 28.729 ;
  LAYER M2 ;
        RECT 6.8 28.811 9.2 28.813 ;
  LAYER M2 ;
        RECT 6.8 28.895 9.2 28.897 ;
  LAYER M2 ;
        RECT 6.8 28.979 9.2 28.981 ;
  LAYER M2 ;
        RECT 6.8 29.063 9.2 29.065 ;
  LAYER M1 ;
        RECT 6.304 17.856 6.336 20.364 ;
  LAYER M1 ;
        RECT 6.24 17.856 6.272 20.364 ;
  LAYER M1 ;
        RECT 6.176 17.856 6.208 20.364 ;
  LAYER M1 ;
        RECT 6.112 17.856 6.144 20.364 ;
  LAYER M1 ;
        RECT 6.048 17.856 6.08 20.364 ;
  LAYER M1 ;
        RECT 5.984 17.856 6.016 20.364 ;
  LAYER M1 ;
        RECT 5.92 17.856 5.952 20.364 ;
  LAYER M1 ;
        RECT 5.856 17.856 5.888 20.364 ;
  LAYER M1 ;
        RECT 5.792 17.856 5.824 20.364 ;
  LAYER M1 ;
        RECT 5.728 17.856 5.76 20.364 ;
  LAYER M1 ;
        RECT 5.664 17.856 5.696 20.364 ;
  LAYER M1 ;
        RECT 5.6 17.856 5.632 20.364 ;
  LAYER M1 ;
        RECT 5.536 17.856 5.568 20.364 ;
  LAYER M1 ;
        RECT 5.472 17.856 5.504 20.364 ;
  LAYER M1 ;
        RECT 5.408 17.856 5.44 20.364 ;
  LAYER M1 ;
        RECT 5.344 17.856 5.376 20.364 ;
  LAYER M1 ;
        RECT 5.28 17.856 5.312 20.364 ;
  LAYER M1 ;
        RECT 5.216 17.856 5.248 20.364 ;
  LAYER M1 ;
        RECT 5.152 17.856 5.184 20.364 ;
  LAYER M1 ;
        RECT 5.088 17.856 5.12 20.364 ;
  LAYER M1 ;
        RECT 5.024 17.856 5.056 20.364 ;
  LAYER M1 ;
        RECT 4.96 17.856 4.992 20.364 ;
  LAYER M1 ;
        RECT 4.896 17.856 4.928 20.364 ;
  LAYER M1 ;
        RECT 4.832 17.856 4.864 20.364 ;
  LAYER M1 ;
        RECT 4.768 17.856 4.8 20.364 ;
  LAYER M1 ;
        RECT 4.704 17.856 4.736 20.364 ;
  LAYER M1 ;
        RECT 4.64 17.856 4.672 20.364 ;
  LAYER M1 ;
        RECT 4.576 17.856 4.608 20.364 ;
  LAYER M1 ;
        RECT 4.512 17.856 4.544 20.364 ;
  LAYER M1 ;
        RECT 4.448 17.856 4.48 20.364 ;
  LAYER M1 ;
        RECT 4.384 17.856 4.416 20.364 ;
  LAYER M1 ;
        RECT 4.32 17.856 4.352 20.364 ;
  LAYER M1 ;
        RECT 4.256 17.856 4.288 20.364 ;
  LAYER M1 ;
        RECT 4.192 17.856 4.224 20.364 ;
  LAYER M1 ;
        RECT 4.128 17.856 4.16 20.364 ;
  LAYER M1 ;
        RECT 4.064 17.856 4.096 20.364 ;
  LAYER M1 ;
        RECT 4 17.856 4.032 20.364 ;
  LAYER M2 ;
        RECT 3.884 17.94 6.356 17.972 ;
  LAYER M2 ;
        RECT 3.884 18.004 6.356 18.036 ;
  LAYER M2 ;
        RECT 3.884 18.068 6.356 18.1 ;
  LAYER M2 ;
        RECT 3.884 18.132 6.356 18.164 ;
  LAYER M2 ;
        RECT 3.884 18.196 6.356 18.228 ;
  LAYER M2 ;
        RECT 3.884 18.26 6.356 18.292 ;
  LAYER M2 ;
        RECT 3.884 18.324 6.356 18.356 ;
  LAYER M2 ;
        RECT 3.884 18.388 6.356 18.42 ;
  LAYER M2 ;
        RECT 3.884 18.452 6.356 18.484 ;
  LAYER M2 ;
        RECT 3.884 18.516 6.356 18.548 ;
  LAYER M2 ;
        RECT 3.884 18.58 6.356 18.612 ;
  LAYER M2 ;
        RECT 3.884 18.644 6.356 18.676 ;
  LAYER M2 ;
        RECT 3.884 18.708 6.356 18.74 ;
  LAYER M2 ;
        RECT 3.884 18.772 6.356 18.804 ;
  LAYER M2 ;
        RECT 3.884 18.836 6.356 18.868 ;
  LAYER M2 ;
        RECT 3.884 18.9 6.356 18.932 ;
  LAYER M2 ;
        RECT 3.884 18.964 6.356 18.996 ;
  LAYER M2 ;
        RECT 3.884 19.028 6.356 19.06 ;
  LAYER M2 ;
        RECT 3.884 19.092 6.356 19.124 ;
  LAYER M2 ;
        RECT 3.884 19.156 6.356 19.188 ;
  LAYER M2 ;
        RECT 3.884 19.22 6.356 19.252 ;
  LAYER M2 ;
        RECT 3.884 19.284 6.356 19.316 ;
  LAYER M2 ;
        RECT 3.884 19.348 6.356 19.38 ;
  LAYER M2 ;
        RECT 3.884 19.412 6.356 19.444 ;
  LAYER M2 ;
        RECT 3.884 19.476 6.356 19.508 ;
  LAYER M2 ;
        RECT 3.884 19.54 6.356 19.572 ;
  LAYER M2 ;
        RECT 3.884 19.604 6.356 19.636 ;
  LAYER M2 ;
        RECT 3.884 19.668 6.356 19.7 ;
  LAYER M2 ;
        RECT 3.884 19.732 6.356 19.764 ;
  LAYER M2 ;
        RECT 3.884 19.796 6.356 19.828 ;
  LAYER M2 ;
        RECT 3.884 19.86 6.356 19.892 ;
  LAYER M2 ;
        RECT 3.884 19.924 6.356 19.956 ;
  LAYER M2 ;
        RECT 3.884 19.988 6.356 20.02 ;
  LAYER M2 ;
        RECT 3.884 20.052 6.356 20.084 ;
  LAYER M2 ;
        RECT 3.884 20.116 6.356 20.148 ;
  LAYER M2 ;
        RECT 3.884 20.18 6.356 20.212 ;
  LAYER M3 ;
        RECT 6.304 17.856 6.336 20.364 ;
  LAYER M3 ;
        RECT 6.24 17.856 6.272 20.364 ;
  LAYER M3 ;
        RECT 6.176 17.856 6.208 20.364 ;
  LAYER M3 ;
        RECT 6.112 17.856 6.144 20.364 ;
  LAYER M3 ;
        RECT 6.048 17.856 6.08 20.364 ;
  LAYER M3 ;
        RECT 5.984 17.856 6.016 20.364 ;
  LAYER M3 ;
        RECT 5.92 17.856 5.952 20.364 ;
  LAYER M3 ;
        RECT 5.856 17.856 5.888 20.364 ;
  LAYER M3 ;
        RECT 5.792 17.856 5.824 20.364 ;
  LAYER M3 ;
        RECT 5.728 17.856 5.76 20.364 ;
  LAYER M3 ;
        RECT 5.664 17.856 5.696 20.364 ;
  LAYER M3 ;
        RECT 5.6 17.856 5.632 20.364 ;
  LAYER M3 ;
        RECT 5.536 17.856 5.568 20.364 ;
  LAYER M3 ;
        RECT 5.472 17.856 5.504 20.364 ;
  LAYER M3 ;
        RECT 5.408 17.856 5.44 20.364 ;
  LAYER M3 ;
        RECT 5.344 17.856 5.376 20.364 ;
  LAYER M3 ;
        RECT 5.28 17.856 5.312 20.364 ;
  LAYER M3 ;
        RECT 5.216 17.856 5.248 20.364 ;
  LAYER M3 ;
        RECT 5.152 17.856 5.184 20.364 ;
  LAYER M3 ;
        RECT 5.088 17.856 5.12 20.364 ;
  LAYER M3 ;
        RECT 5.024 17.856 5.056 20.364 ;
  LAYER M3 ;
        RECT 4.96 17.856 4.992 20.364 ;
  LAYER M3 ;
        RECT 4.896 17.856 4.928 20.364 ;
  LAYER M3 ;
        RECT 4.832 17.856 4.864 20.364 ;
  LAYER M3 ;
        RECT 4.768 17.856 4.8 20.364 ;
  LAYER M3 ;
        RECT 4.704 17.856 4.736 20.364 ;
  LAYER M3 ;
        RECT 4.64 17.856 4.672 20.364 ;
  LAYER M3 ;
        RECT 4.576 17.856 4.608 20.364 ;
  LAYER M3 ;
        RECT 4.512 17.856 4.544 20.364 ;
  LAYER M3 ;
        RECT 4.448 17.856 4.48 20.364 ;
  LAYER M3 ;
        RECT 4.384 17.856 4.416 20.364 ;
  LAYER M3 ;
        RECT 4.32 17.856 4.352 20.364 ;
  LAYER M3 ;
        RECT 4.256 17.856 4.288 20.364 ;
  LAYER M3 ;
        RECT 4.192 17.856 4.224 20.364 ;
  LAYER M3 ;
        RECT 4.128 17.856 4.16 20.364 ;
  LAYER M3 ;
        RECT 4.064 17.856 4.096 20.364 ;
  LAYER M3 ;
        RECT 4 17.856 4.032 20.364 ;
  LAYER M3 ;
        RECT 3.904 17.856 3.936 20.364 ;
  LAYER M1 ;
        RECT 6.319 17.892 6.321 20.328 ;
  LAYER M1 ;
        RECT 6.239 17.892 6.241 20.328 ;
  LAYER M1 ;
        RECT 6.159 17.892 6.161 20.328 ;
  LAYER M1 ;
        RECT 6.079 17.892 6.081 20.328 ;
  LAYER M1 ;
        RECT 5.999 17.892 6.001 20.328 ;
  LAYER M1 ;
        RECT 5.919 17.892 5.921 20.328 ;
  LAYER M1 ;
        RECT 5.839 17.892 5.841 20.328 ;
  LAYER M1 ;
        RECT 5.759 17.892 5.761 20.328 ;
  LAYER M1 ;
        RECT 5.679 17.892 5.681 20.328 ;
  LAYER M1 ;
        RECT 5.599 17.892 5.601 20.328 ;
  LAYER M1 ;
        RECT 5.519 17.892 5.521 20.328 ;
  LAYER M1 ;
        RECT 5.439 17.892 5.441 20.328 ;
  LAYER M1 ;
        RECT 5.359 17.892 5.361 20.328 ;
  LAYER M1 ;
        RECT 5.279 17.892 5.281 20.328 ;
  LAYER M1 ;
        RECT 5.199 17.892 5.201 20.328 ;
  LAYER M1 ;
        RECT 5.119 17.892 5.121 20.328 ;
  LAYER M1 ;
        RECT 5.039 17.892 5.041 20.328 ;
  LAYER M1 ;
        RECT 4.959 17.892 4.961 20.328 ;
  LAYER M1 ;
        RECT 4.879 17.892 4.881 20.328 ;
  LAYER M1 ;
        RECT 4.799 17.892 4.801 20.328 ;
  LAYER M1 ;
        RECT 4.719 17.892 4.721 20.328 ;
  LAYER M1 ;
        RECT 4.639 17.892 4.641 20.328 ;
  LAYER M1 ;
        RECT 4.559 17.892 4.561 20.328 ;
  LAYER M1 ;
        RECT 4.479 17.892 4.481 20.328 ;
  LAYER M1 ;
        RECT 4.399 17.892 4.401 20.328 ;
  LAYER M1 ;
        RECT 4.319 17.892 4.321 20.328 ;
  LAYER M1 ;
        RECT 4.239 17.892 4.241 20.328 ;
  LAYER M1 ;
        RECT 4.159 17.892 4.161 20.328 ;
  LAYER M1 ;
        RECT 4.079 17.892 4.081 20.328 ;
  LAYER M1 ;
        RECT 3.999 17.892 4.001 20.328 ;
  LAYER M2 ;
        RECT 3.92 17.891 6.32 17.893 ;
  LAYER M2 ;
        RECT 3.92 17.975 6.32 17.977 ;
  LAYER M2 ;
        RECT 3.92 18.059 6.32 18.061 ;
  LAYER M2 ;
        RECT 3.92 18.143 6.32 18.145 ;
  LAYER M2 ;
        RECT 3.92 18.227 6.32 18.229 ;
  LAYER M2 ;
        RECT 3.92 18.311 6.32 18.313 ;
  LAYER M2 ;
        RECT 3.92 18.395 6.32 18.397 ;
  LAYER M2 ;
        RECT 3.92 18.479 6.32 18.481 ;
  LAYER M2 ;
        RECT 3.92 18.563 6.32 18.565 ;
  LAYER M2 ;
        RECT 3.92 18.647 6.32 18.649 ;
  LAYER M2 ;
        RECT 3.92 18.731 6.32 18.733 ;
  LAYER M2 ;
        RECT 3.92 18.815 6.32 18.817 ;
  LAYER M2 ;
        RECT 3.92 18.8985 6.32 18.9005 ;
  LAYER M2 ;
        RECT 3.92 18.983 6.32 18.985 ;
  LAYER M2 ;
        RECT 3.92 19.067 6.32 19.069 ;
  LAYER M2 ;
        RECT 3.92 19.151 6.32 19.153 ;
  LAYER M2 ;
        RECT 3.92 19.235 6.32 19.237 ;
  LAYER M2 ;
        RECT 3.92 19.319 6.32 19.321 ;
  LAYER M2 ;
        RECT 3.92 19.403 6.32 19.405 ;
  LAYER M2 ;
        RECT 3.92 19.487 6.32 19.489 ;
  LAYER M2 ;
        RECT 3.92 19.571 6.32 19.573 ;
  LAYER M2 ;
        RECT 3.92 19.655 6.32 19.657 ;
  LAYER M2 ;
        RECT 3.92 19.739 6.32 19.741 ;
  LAYER M2 ;
        RECT 3.92 19.823 6.32 19.825 ;
  LAYER M2 ;
        RECT 3.92 19.907 6.32 19.909 ;
  LAYER M2 ;
        RECT 3.92 19.991 6.32 19.993 ;
  LAYER M2 ;
        RECT 3.92 20.075 6.32 20.077 ;
  LAYER M2 ;
        RECT 3.92 20.159 6.32 20.161 ;
  LAYER M2 ;
        RECT 3.92 20.243 6.32 20.245 ;
  LAYER M1 ;
        RECT 6.304 20.796 6.336 23.304 ;
  LAYER M1 ;
        RECT 6.24 20.796 6.272 23.304 ;
  LAYER M1 ;
        RECT 6.176 20.796 6.208 23.304 ;
  LAYER M1 ;
        RECT 6.112 20.796 6.144 23.304 ;
  LAYER M1 ;
        RECT 6.048 20.796 6.08 23.304 ;
  LAYER M1 ;
        RECT 5.984 20.796 6.016 23.304 ;
  LAYER M1 ;
        RECT 5.92 20.796 5.952 23.304 ;
  LAYER M1 ;
        RECT 5.856 20.796 5.888 23.304 ;
  LAYER M1 ;
        RECT 5.792 20.796 5.824 23.304 ;
  LAYER M1 ;
        RECT 5.728 20.796 5.76 23.304 ;
  LAYER M1 ;
        RECT 5.664 20.796 5.696 23.304 ;
  LAYER M1 ;
        RECT 5.6 20.796 5.632 23.304 ;
  LAYER M1 ;
        RECT 5.536 20.796 5.568 23.304 ;
  LAYER M1 ;
        RECT 5.472 20.796 5.504 23.304 ;
  LAYER M1 ;
        RECT 5.408 20.796 5.44 23.304 ;
  LAYER M1 ;
        RECT 5.344 20.796 5.376 23.304 ;
  LAYER M1 ;
        RECT 5.28 20.796 5.312 23.304 ;
  LAYER M1 ;
        RECT 5.216 20.796 5.248 23.304 ;
  LAYER M1 ;
        RECT 5.152 20.796 5.184 23.304 ;
  LAYER M1 ;
        RECT 5.088 20.796 5.12 23.304 ;
  LAYER M1 ;
        RECT 5.024 20.796 5.056 23.304 ;
  LAYER M1 ;
        RECT 4.96 20.796 4.992 23.304 ;
  LAYER M1 ;
        RECT 4.896 20.796 4.928 23.304 ;
  LAYER M1 ;
        RECT 4.832 20.796 4.864 23.304 ;
  LAYER M1 ;
        RECT 4.768 20.796 4.8 23.304 ;
  LAYER M1 ;
        RECT 4.704 20.796 4.736 23.304 ;
  LAYER M1 ;
        RECT 4.64 20.796 4.672 23.304 ;
  LAYER M1 ;
        RECT 4.576 20.796 4.608 23.304 ;
  LAYER M1 ;
        RECT 4.512 20.796 4.544 23.304 ;
  LAYER M1 ;
        RECT 4.448 20.796 4.48 23.304 ;
  LAYER M1 ;
        RECT 4.384 20.796 4.416 23.304 ;
  LAYER M1 ;
        RECT 4.32 20.796 4.352 23.304 ;
  LAYER M1 ;
        RECT 4.256 20.796 4.288 23.304 ;
  LAYER M1 ;
        RECT 4.192 20.796 4.224 23.304 ;
  LAYER M1 ;
        RECT 4.128 20.796 4.16 23.304 ;
  LAYER M1 ;
        RECT 4.064 20.796 4.096 23.304 ;
  LAYER M1 ;
        RECT 4 20.796 4.032 23.304 ;
  LAYER M2 ;
        RECT 3.884 20.88 6.356 20.912 ;
  LAYER M2 ;
        RECT 3.884 20.944 6.356 20.976 ;
  LAYER M2 ;
        RECT 3.884 21.008 6.356 21.04 ;
  LAYER M2 ;
        RECT 3.884 21.072 6.356 21.104 ;
  LAYER M2 ;
        RECT 3.884 21.136 6.356 21.168 ;
  LAYER M2 ;
        RECT 3.884 21.2 6.356 21.232 ;
  LAYER M2 ;
        RECT 3.884 21.264 6.356 21.296 ;
  LAYER M2 ;
        RECT 3.884 21.328 6.356 21.36 ;
  LAYER M2 ;
        RECT 3.884 21.392 6.356 21.424 ;
  LAYER M2 ;
        RECT 3.884 21.456 6.356 21.488 ;
  LAYER M2 ;
        RECT 3.884 21.52 6.356 21.552 ;
  LAYER M2 ;
        RECT 3.884 21.584 6.356 21.616 ;
  LAYER M2 ;
        RECT 3.884 21.648 6.356 21.68 ;
  LAYER M2 ;
        RECT 3.884 21.712 6.356 21.744 ;
  LAYER M2 ;
        RECT 3.884 21.776 6.356 21.808 ;
  LAYER M2 ;
        RECT 3.884 21.84 6.356 21.872 ;
  LAYER M2 ;
        RECT 3.884 21.904 6.356 21.936 ;
  LAYER M2 ;
        RECT 3.884 21.968 6.356 22 ;
  LAYER M2 ;
        RECT 3.884 22.032 6.356 22.064 ;
  LAYER M2 ;
        RECT 3.884 22.096 6.356 22.128 ;
  LAYER M2 ;
        RECT 3.884 22.16 6.356 22.192 ;
  LAYER M2 ;
        RECT 3.884 22.224 6.356 22.256 ;
  LAYER M2 ;
        RECT 3.884 22.288 6.356 22.32 ;
  LAYER M2 ;
        RECT 3.884 22.352 6.356 22.384 ;
  LAYER M2 ;
        RECT 3.884 22.416 6.356 22.448 ;
  LAYER M2 ;
        RECT 3.884 22.48 6.356 22.512 ;
  LAYER M2 ;
        RECT 3.884 22.544 6.356 22.576 ;
  LAYER M2 ;
        RECT 3.884 22.608 6.356 22.64 ;
  LAYER M2 ;
        RECT 3.884 22.672 6.356 22.704 ;
  LAYER M2 ;
        RECT 3.884 22.736 6.356 22.768 ;
  LAYER M2 ;
        RECT 3.884 22.8 6.356 22.832 ;
  LAYER M2 ;
        RECT 3.884 22.864 6.356 22.896 ;
  LAYER M2 ;
        RECT 3.884 22.928 6.356 22.96 ;
  LAYER M2 ;
        RECT 3.884 22.992 6.356 23.024 ;
  LAYER M2 ;
        RECT 3.884 23.056 6.356 23.088 ;
  LAYER M2 ;
        RECT 3.884 23.12 6.356 23.152 ;
  LAYER M3 ;
        RECT 6.304 20.796 6.336 23.304 ;
  LAYER M3 ;
        RECT 6.24 20.796 6.272 23.304 ;
  LAYER M3 ;
        RECT 6.176 20.796 6.208 23.304 ;
  LAYER M3 ;
        RECT 6.112 20.796 6.144 23.304 ;
  LAYER M3 ;
        RECT 6.048 20.796 6.08 23.304 ;
  LAYER M3 ;
        RECT 5.984 20.796 6.016 23.304 ;
  LAYER M3 ;
        RECT 5.92 20.796 5.952 23.304 ;
  LAYER M3 ;
        RECT 5.856 20.796 5.888 23.304 ;
  LAYER M3 ;
        RECT 5.792 20.796 5.824 23.304 ;
  LAYER M3 ;
        RECT 5.728 20.796 5.76 23.304 ;
  LAYER M3 ;
        RECT 5.664 20.796 5.696 23.304 ;
  LAYER M3 ;
        RECT 5.6 20.796 5.632 23.304 ;
  LAYER M3 ;
        RECT 5.536 20.796 5.568 23.304 ;
  LAYER M3 ;
        RECT 5.472 20.796 5.504 23.304 ;
  LAYER M3 ;
        RECT 5.408 20.796 5.44 23.304 ;
  LAYER M3 ;
        RECT 5.344 20.796 5.376 23.304 ;
  LAYER M3 ;
        RECT 5.28 20.796 5.312 23.304 ;
  LAYER M3 ;
        RECT 5.216 20.796 5.248 23.304 ;
  LAYER M3 ;
        RECT 5.152 20.796 5.184 23.304 ;
  LAYER M3 ;
        RECT 5.088 20.796 5.12 23.304 ;
  LAYER M3 ;
        RECT 5.024 20.796 5.056 23.304 ;
  LAYER M3 ;
        RECT 4.96 20.796 4.992 23.304 ;
  LAYER M3 ;
        RECT 4.896 20.796 4.928 23.304 ;
  LAYER M3 ;
        RECT 4.832 20.796 4.864 23.304 ;
  LAYER M3 ;
        RECT 4.768 20.796 4.8 23.304 ;
  LAYER M3 ;
        RECT 4.704 20.796 4.736 23.304 ;
  LAYER M3 ;
        RECT 4.64 20.796 4.672 23.304 ;
  LAYER M3 ;
        RECT 4.576 20.796 4.608 23.304 ;
  LAYER M3 ;
        RECT 4.512 20.796 4.544 23.304 ;
  LAYER M3 ;
        RECT 4.448 20.796 4.48 23.304 ;
  LAYER M3 ;
        RECT 4.384 20.796 4.416 23.304 ;
  LAYER M3 ;
        RECT 4.32 20.796 4.352 23.304 ;
  LAYER M3 ;
        RECT 4.256 20.796 4.288 23.304 ;
  LAYER M3 ;
        RECT 4.192 20.796 4.224 23.304 ;
  LAYER M3 ;
        RECT 4.128 20.796 4.16 23.304 ;
  LAYER M3 ;
        RECT 4.064 20.796 4.096 23.304 ;
  LAYER M3 ;
        RECT 4 20.796 4.032 23.304 ;
  LAYER M3 ;
        RECT 3.904 20.796 3.936 23.304 ;
  LAYER M1 ;
        RECT 6.319 20.832 6.321 23.268 ;
  LAYER M1 ;
        RECT 6.239 20.832 6.241 23.268 ;
  LAYER M1 ;
        RECT 6.159 20.832 6.161 23.268 ;
  LAYER M1 ;
        RECT 6.079 20.832 6.081 23.268 ;
  LAYER M1 ;
        RECT 5.999 20.832 6.001 23.268 ;
  LAYER M1 ;
        RECT 5.919 20.832 5.921 23.268 ;
  LAYER M1 ;
        RECT 5.839 20.832 5.841 23.268 ;
  LAYER M1 ;
        RECT 5.759 20.832 5.761 23.268 ;
  LAYER M1 ;
        RECT 5.679 20.832 5.681 23.268 ;
  LAYER M1 ;
        RECT 5.599 20.832 5.601 23.268 ;
  LAYER M1 ;
        RECT 5.519 20.832 5.521 23.268 ;
  LAYER M1 ;
        RECT 5.439 20.832 5.441 23.268 ;
  LAYER M1 ;
        RECT 5.359 20.832 5.361 23.268 ;
  LAYER M1 ;
        RECT 5.279 20.832 5.281 23.268 ;
  LAYER M1 ;
        RECT 5.199 20.832 5.201 23.268 ;
  LAYER M1 ;
        RECT 5.119 20.832 5.121 23.268 ;
  LAYER M1 ;
        RECT 5.039 20.832 5.041 23.268 ;
  LAYER M1 ;
        RECT 4.959 20.832 4.961 23.268 ;
  LAYER M1 ;
        RECT 4.879 20.832 4.881 23.268 ;
  LAYER M1 ;
        RECT 4.799 20.832 4.801 23.268 ;
  LAYER M1 ;
        RECT 4.719 20.832 4.721 23.268 ;
  LAYER M1 ;
        RECT 4.639 20.832 4.641 23.268 ;
  LAYER M1 ;
        RECT 4.559 20.832 4.561 23.268 ;
  LAYER M1 ;
        RECT 4.479 20.832 4.481 23.268 ;
  LAYER M1 ;
        RECT 4.399 20.832 4.401 23.268 ;
  LAYER M1 ;
        RECT 4.319 20.832 4.321 23.268 ;
  LAYER M1 ;
        RECT 4.239 20.832 4.241 23.268 ;
  LAYER M1 ;
        RECT 4.159 20.832 4.161 23.268 ;
  LAYER M1 ;
        RECT 4.079 20.832 4.081 23.268 ;
  LAYER M1 ;
        RECT 3.999 20.832 4.001 23.268 ;
  LAYER M2 ;
        RECT 3.92 20.831 6.32 20.833 ;
  LAYER M2 ;
        RECT 3.92 20.915 6.32 20.917 ;
  LAYER M2 ;
        RECT 3.92 20.999 6.32 21.001 ;
  LAYER M2 ;
        RECT 3.92 21.083 6.32 21.085 ;
  LAYER M2 ;
        RECT 3.92 21.167 6.32 21.169 ;
  LAYER M2 ;
        RECT 3.92 21.251 6.32 21.253 ;
  LAYER M2 ;
        RECT 3.92 21.335 6.32 21.337 ;
  LAYER M2 ;
        RECT 3.92 21.419 6.32 21.421 ;
  LAYER M2 ;
        RECT 3.92 21.503 6.32 21.505 ;
  LAYER M2 ;
        RECT 3.92 21.587 6.32 21.589 ;
  LAYER M2 ;
        RECT 3.92 21.671 6.32 21.673 ;
  LAYER M2 ;
        RECT 3.92 21.755 6.32 21.757 ;
  LAYER M2 ;
        RECT 3.92 21.8385 6.32 21.8405 ;
  LAYER M2 ;
        RECT 3.92 21.923 6.32 21.925 ;
  LAYER M2 ;
        RECT 3.92 22.007 6.32 22.009 ;
  LAYER M2 ;
        RECT 3.92 22.091 6.32 22.093 ;
  LAYER M2 ;
        RECT 3.92 22.175 6.32 22.177 ;
  LAYER M2 ;
        RECT 3.92 22.259 6.32 22.261 ;
  LAYER M2 ;
        RECT 3.92 22.343 6.32 22.345 ;
  LAYER M2 ;
        RECT 3.92 22.427 6.32 22.429 ;
  LAYER M2 ;
        RECT 3.92 22.511 6.32 22.513 ;
  LAYER M2 ;
        RECT 3.92 22.595 6.32 22.597 ;
  LAYER M2 ;
        RECT 3.92 22.679 6.32 22.681 ;
  LAYER M2 ;
        RECT 3.92 22.763 6.32 22.765 ;
  LAYER M2 ;
        RECT 3.92 22.847 6.32 22.849 ;
  LAYER M2 ;
        RECT 3.92 22.931 6.32 22.933 ;
  LAYER M2 ;
        RECT 3.92 23.015 6.32 23.017 ;
  LAYER M2 ;
        RECT 3.92 23.099 6.32 23.101 ;
  LAYER M2 ;
        RECT 3.92 23.183 6.32 23.185 ;
  LAYER M1 ;
        RECT 6.304 23.736 6.336 26.244 ;
  LAYER M1 ;
        RECT 6.24 23.736 6.272 26.244 ;
  LAYER M1 ;
        RECT 6.176 23.736 6.208 26.244 ;
  LAYER M1 ;
        RECT 6.112 23.736 6.144 26.244 ;
  LAYER M1 ;
        RECT 6.048 23.736 6.08 26.244 ;
  LAYER M1 ;
        RECT 5.984 23.736 6.016 26.244 ;
  LAYER M1 ;
        RECT 5.92 23.736 5.952 26.244 ;
  LAYER M1 ;
        RECT 5.856 23.736 5.888 26.244 ;
  LAYER M1 ;
        RECT 5.792 23.736 5.824 26.244 ;
  LAYER M1 ;
        RECT 5.728 23.736 5.76 26.244 ;
  LAYER M1 ;
        RECT 5.664 23.736 5.696 26.244 ;
  LAYER M1 ;
        RECT 5.6 23.736 5.632 26.244 ;
  LAYER M1 ;
        RECT 5.536 23.736 5.568 26.244 ;
  LAYER M1 ;
        RECT 5.472 23.736 5.504 26.244 ;
  LAYER M1 ;
        RECT 5.408 23.736 5.44 26.244 ;
  LAYER M1 ;
        RECT 5.344 23.736 5.376 26.244 ;
  LAYER M1 ;
        RECT 5.28 23.736 5.312 26.244 ;
  LAYER M1 ;
        RECT 5.216 23.736 5.248 26.244 ;
  LAYER M1 ;
        RECT 5.152 23.736 5.184 26.244 ;
  LAYER M1 ;
        RECT 5.088 23.736 5.12 26.244 ;
  LAYER M1 ;
        RECT 5.024 23.736 5.056 26.244 ;
  LAYER M1 ;
        RECT 4.96 23.736 4.992 26.244 ;
  LAYER M1 ;
        RECT 4.896 23.736 4.928 26.244 ;
  LAYER M1 ;
        RECT 4.832 23.736 4.864 26.244 ;
  LAYER M1 ;
        RECT 4.768 23.736 4.8 26.244 ;
  LAYER M1 ;
        RECT 4.704 23.736 4.736 26.244 ;
  LAYER M1 ;
        RECT 4.64 23.736 4.672 26.244 ;
  LAYER M1 ;
        RECT 4.576 23.736 4.608 26.244 ;
  LAYER M1 ;
        RECT 4.512 23.736 4.544 26.244 ;
  LAYER M1 ;
        RECT 4.448 23.736 4.48 26.244 ;
  LAYER M1 ;
        RECT 4.384 23.736 4.416 26.244 ;
  LAYER M1 ;
        RECT 4.32 23.736 4.352 26.244 ;
  LAYER M1 ;
        RECT 4.256 23.736 4.288 26.244 ;
  LAYER M1 ;
        RECT 4.192 23.736 4.224 26.244 ;
  LAYER M1 ;
        RECT 4.128 23.736 4.16 26.244 ;
  LAYER M1 ;
        RECT 4.064 23.736 4.096 26.244 ;
  LAYER M1 ;
        RECT 4 23.736 4.032 26.244 ;
  LAYER M2 ;
        RECT 3.884 23.82 6.356 23.852 ;
  LAYER M2 ;
        RECT 3.884 23.884 6.356 23.916 ;
  LAYER M2 ;
        RECT 3.884 23.948 6.356 23.98 ;
  LAYER M2 ;
        RECT 3.884 24.012 6.356 24.044 ;
  LAYER M2 ;
        RECT 3.884 24.076 6.356 24.108 ;
  LAYER M2 ;
        RECT 3.884 24.14 6.356 24.172 ;
  LAYER M2 ;
        RECT 3.884 24.204 6.356 24.236 ;
  LAYER M2 ;
        RECT 3.884 24.268 6.356 24.3 ;
  LAYER M2 ;
        RECT 3.884 24.332 6.356 24.364 ;
  LAYER M2 ;
        RECT 3.884 24.396 6.356 24.428 ;
  LAYER M2 ;
        RECT 3.884 24.46 6.356 24.492 ;
  LAYER M2 ;
        RECT 3.884 24.524 6.356 24.556 ;
  LAYER M2 ;
        RECT 3.884 24.588 6.356 24.62 ;
  LAYER M2 ;
        RECT 3.884 24.652 6.356 24.684 ;
  LAYER M2 ;
        RECT 3.884 24.716 6.356 24.748 ;
  LAYER M2 ;
        RECT 3.884 24.78 6.356 24.812 ;
  LAYER M2 ;
        RECT 3.884 24.844 6.356 24.876 ;
  LAYER M2 ;
        RECT 3.884 24.908 6.356 24.94 ;
  LAYER M2 ;
        RECT 3.884 24.972 6.356 25.004 ;
  LAYER M2 ;
        RECT 3.884 25.036 6.356 25.068 ;
  LAYER M2 ;
        RECT 3.884 25.1 6.356 25.132 ;
  LAYER M2 ;
        RECT 3.884 25.164 6.356 25.196 ;
  LAYER M2 ;
        RECT 3.884 25.228 6.356 25.26 ;
  LAYER M2 ;
        RECT 3.884 25.292 6.356 25.324 ;
  LAYER M2 ;
        RECT 3.884 25.356 6.356 25.388 ;
  LAYER M2 ;
        RECT 3.884 25.42 6.356 25.452 ;
  LAYER M2 ;
        RECT 3.884 25.484 6.356 25.516 ;
  LAYER M2 ;
        RECT 3.884 25.548 6.356 25.58 ;
  LAYER M2 ;
        RECT 3.884 25.612 6.356 25.644 ;
  LAYER M2 ;
        RECT 3.884 25.676 6.356 25.708 ;
  LAYER M2 ;
        RECT 3.884 25.74 6.356 25.772 ;
  LAYER M2 ;
        RECT 3.884 25.804 6.356 25.836 ;
  LAYER M2 ;
        RECT 3.884 25.868 6.356 25.9 ;
  LAYER M2 ;
        RECT 3.884 25.932 6.356 25.964 ;
  LAYER M2 ;
        RECT 3.884 25.996 6.356 26.028 ;
  LAYER M2 ;
        RECT 3.884 26.06 6.356 26.092 ;
  LAYER M3 ;
        RECT 6.304 23.736 6.336 26.244 ;
  LAYER M3 ;
        RECT 6.24 23.736 6.272 26.244 ;
  LAYER M3 ;
        RECT 6.176 23.736 6.208 26.244 ;
  LAYER M3 ;
        RECT 6.112 23.736 6.144 26.244 ;
  LAYER M3 ;
        RECT 6.048 23.736 6.08 26.244 ;
  LAYER M3 ;
        RECT 5.984 23.736 6.016 26.244 ;
  LAYER M3 ;
        RECT 5.92 23.736 5.952 26.244 ;
  LAYER M3 ;
        RECT 5.856 23.736 5.888 26.244 ;
  LAYER M3 ;
        RECT 5.792 23.736 5.824 26.244 ;
  LAYER M3 ;
        RECT 5.728 23.736 5.76 26.244 ;
  LAYER M3 ;
        RECT 5.664 23.736 5.696 26.244 ;
  LAYER M3 ;
        RECT 5.6 23.736 5.632 26.244 ;
  LAYER M3 ;
        RECT 5.536 23.736 5.568 26.244 ;
  LAYER M3 ;
        RECT 5.472 23.736 5.504 26.244 ;
  LAYER M3 ;
        RECT 5.408 23.736 5.44 26.244 ;
  LAYER M3 ;
        RECT 5.344 23.736 5.376 26.244 ;
  LAYER M3 ;
        RECT 5.28 23.736 5.312 26.244 ;
  LAYER M3 ;
        RECT 5.216 23.736 5.248 26.244 ;
  LAYER M3 ;
        RECT 5.152 23.736 5.184 26.244 ;
  LAYER M3 ;
        RECT 5.088 23.736 5.12 26.244 ;
  LAYER M3 ;
        RECT 5.024 23.736 5.056 26.244 ;
  LAYER M3 ;
        RECT 4.96 23.736 4.992 26.244 ;
  LAYER M3 ;
        RECT 4.896 23.736 4.928 26.244 ;
  LAYER M3 ;
        RECT 4.832 23.736 4.864 26.244 ;
  LAYER M3 ;
        RECT 4.768 23.736 4.8 26.244 ;
  LAYER M3 ;
        RECT 4.704 23.736 4.736 26.244 ;
  LAYER M3 ;
        RECT 4.64 23.736 4.672 26.244 ;
  LAYER M3 ;
        RECT 4.576 23.736 4.608 26.244 ;
  LAYER M3 ;
        RECT 4.512 23.736 4.544 26.244 ;
  LAYER M3 ;
        RECT 4.448 23.736 4.48 26.244 ;
  LAYER M3 ;
        RECT 4.384 23.736 4.416 26.244 ;
  LAYER M3 ;
        RECT 4.32 23.736 4.352 26.244 ;
  LAYER M3 ;
        RECT 4.256 23.736 4.288 26.244 ;
  LAYER M3 ;
        RECT 4.192 23.736 4.224 26.244 ;
  LAYER M3 ;
        RECT 4.128 23.736 4.16 26.244 ;
  LAYER M3 ;
        RECT 4.064 23.736 4.096 26.244 ;
  LAYER M3 ;
        RECT 4 23.736 4.032 26.244 ;
  LAYER M3 ;
        RECT 3.904 23.736 3.936 26.244 ;
  LAYER M1 ;
        RECT 6.319 23.772 6.321 26.208 ;
  LAYER M1 ;
        RECT 6.239 23.772 6.241 26.208 ;
  LAYER M1 ;
        RECT 6.159 23.772 6.161 26.208 ;
  LAYER M1 ;
        RECT 6.079 23.772 6.081 26.208 ;
  LAYER M1 ;
        RECT 5.999 23.772 6.001 26.208 ;
  LAYER M1 ;
        RECT 5.919 23.772 5.921 26.208 ;
  LAYER M1 ;
        RECT 5.839 23.772 5.841 26.208 ;
  LAYER M1 ;
        RECT 5.759 23.772 5.761 26.208 ;
  LAYER M1 ;
        RECT 5.679 23.772 5.681 26.208 ;
  LAYER M1 ;
        RECT 5.599 23.772 5.601 26.208 ;
  LAYER M1 ;
        RECT 5.519 23.772 5.521 26.208 ;
  LAYER M1 ;
        RECT 5.439 23.772 5.441 26.208 ;
  LAYER M1 ;
        RECT 5.359 23.772 5.361 26.208 ;
  LAYER M1 ;
        RECT 5.279 23.772 5.281 26.208 ;
  LAYER M1 ;
        RECT 5.199 23.772 5.201 26.208 ;
  LAYER M1 ;
        RECT 5.119 23.772 5.121 26.208 ;
  LAYER M1 ;
        RECT 5.039 23.772 5.041 26.208 ;
  LAYER M1 ;
        RECT 4.959 23.772 4.961 26.208 ;
  LAYER M1 ;
        RECT 4.879 23.772 4.881 26.208 ;
  LAYER M1 ;
        RECT 4.799 23.772 4.801 26.208 ;
  LAYER M1 ;
        RECT 4.719 23.772 4.721 26.208 ;
  LAYER M1 ;
        RECT 4.639 23.772 4.641 26.208 ;
  LAYER M1 ;
        RECT 4.559 23.772 4.561 26.208 ;
  LAYER M1 ;
        RECT 4.479 23.772 4.481 26.208 ;
  LAYER M1 ;
        RECT 4.399 23.772 4.401 26.208 ;
  LAYER M1 ;
        RECT 4.319 23.772 4.321 26.208 ;
  LAYER M1 ;
        RECT 4.239 23.772 4.241 26.208 ;
  LAYER M1 ;
        RECT 4.159 23.772 4.161 26.208 ;
  LAYER M1 ;
        RECT 4.079 23.772 4.081 26.208 ;
  LAYER M1 ;
        RECT 3.999 23.772 4.001 26.208 ;
  LAYER M2 ;
        RECT 3.92 23.771 6.32 23.773 ;
  LAYER M2 ;
        RECT 3.92 23.855 6.32 23.857 ;
  LAYER M2 ;
        RECT 3.92 23.939 6.32 23.941 ;
  LAYER M2 ;
        RECT 3.92 24.023 6.32 24.025 ;
  LAYER M2 ;
        RECT 3.92 24.107 6.32 24.109 ;
  LAYER M2 ;
        RECT 3.92 24.191 6.32 24.193 ;
  LAYER M2 ;
        RECT 3.92 24.275 6.32 24.277 ;
  LAYER M2 ;
        RECT 3.92 24.359 6.32 24.361 ;
  LAYER M2 ;
        RECT 3.92 24.443 6.32 24.445 ;
  LAYER M2 ;
        RECT 3.92 24.527 6.32 24.529 ;
  LAYER M2 ;
        RECT 3.92 24.611 6.32 24.613 ;
  LAYER M2 ;
        RECT 3.92 24.695 6.32 24.697 ;
  LAYER M2 ;
        RECT 3.92 24.7785 6.32 24.7805 ;
  LAYER M2 ;
        RECT 3.92 24.863 6.32 24.865 ;
  LAYER M2 ;
        RECT 3.92 24.947 6.32 24.949 ;
  LAYER M2 ;
        RECT 3.92 25.031 6.32 25.033 ;
  LAYER M2 ;
        RECT 3.92 25.115 6.32 25.117 ;
  LAYER M2 ;
        RECT 3.92 25.199 6.32 25.201 ;
  LAYER M2 ;
        RECT 3.92 25.283 6.32 25.285 ;
  LAYER M2 ;
        RECT 3.92 25.367 6.32 25.369 ;
  LAYER M2 ;
        RECT 3.92 25.451 6.32 25.453 ;
  LAYER M2 ;
        RECT 3.92 25.535 6.32 25.537 ;
  LAYER M2 ;
        RECT 3.92 25.619 6.32 25.621 ;
  LAYER M2 ;
        RECT 3.92 25.703 6.32 25.705 ;
  LAYER M2 ;
        RECT 3.92 25.787 6.32 25.789 ;
  LAYER M2 ;
        RECT 3.92 25.871 6.32 25.873 ;
  LAYER M2 ;
        RECT 3.92 25.955 6.32 25.957 ;
  LAYER M2 ;
        RECT 3.92 26.039 6.32 26.041 ;
  LAYER M2 ;
        RECT 3.92 26.123 6.32 26.125 ;
  LAYER M1 ;
        RECT 6.304 26.676 6.336 29.184 ;
  LAYER M1 ;
        RECT 6.24 26.676 6.272 29.184 ;
  LAYER M1 ;
        RECT 6.176 26.676 6.208 29.184 ;
  LAYER M1 ;
        RECT 6.112 26.676 6.144 29.184 ;
  LAYER M1 ;
        RECT 6.048 26.676 6.08 29.184 ;
  LAYER M1 ;
        RECT 5.984 26.676 6.016 29.184 ;
  LAYER M1 ;
        RECT 5.92 26.676 5.952 29.184 ;
  LAYER M1 ;
        RECT 5.856 26.676 5.888 29.184 ;
  LAYER M1 ;
        RECT 5.792 26.676 5.824 29.184 ;
  LAYER M1 ;
        RECT 5.728 26.676 5.76 29.184 ;
  LAYER M1 ;
        RECT 5.664 26.676 5.696 29.184 ;
  LAYER M1 ;
        RECT 5.6 26.676 5.632 29.184 ;
  LAYER M1 ;
        RECT 5.536 26.676 5.568 29.184 ;
  LAYER M1 ;
        RECT 5.472 26.676 5.504 29.184 ;
  LAYER M1 ;
        RECT 5.408 26.676 5.44 29.184 ;
  LAYER M1 ;
        RECT 5.344 26.676 5.376 29.184 ;
  LAYER M1 ;
        RECT 5.28 26.676 5.312 29.184 ;
  LAYER M1 ;
        RECT 5.216 26.676 5.248 29.184 ;
  LAYER M1 ;
        RECT 5.152 26.676 5.184 29.184 ;
  LAYER M1 ;
        RECT 5.088 26.676 5.12 29.184 ;
  LAYER M1 ;
        RECT 5.024 26.676 5.056 29.184 ;
  LAYER M1 ;
        RECT 4.96 26.676 4.992 29.184 ;
  LAYER M1 ;
        RECT 4.896 26.676 4.928 29.184 ;
  LAYER M1 ;
        RECT 4.832 26.676 4.864 29.184 ;
  LAYER M1 ;
        RECT 4.768 26.676 4.8 29.184 ;
  LAYER M1 ;
        RECT 4.704 26.676 4.736 29.184 ;
  LAYER M1 ;
        RECT 4.64 26.676 4.672 29.184 ;
  LAYER M1 ;
        RECT 4.576 26.676 4.608 29.184 ;
  LAYER M1 ;
        RECT 4.512 26.676 4.544 29.184 ;
  LAYER M1 ;
        RECT 4.448 26.676 4.48 29.184 ;
  LAYER M1 ;
        RECT 4.384 26.676 4.416 29.184 ;
  LAYER M1 ;
        RECT 4.32 26.676 4.352 29.184 ;
  LAYER M1 ;
        RECT 4.256 26.676 4.288 29.184 ;
  LAYER M1 ;
        RECT 4.192 26.676 4.224 29.184 ;
  LAYER M1 ;
        RECT 4.128 26.676 4.16 29.184 ;
  LAYER M1 ;
        RECT 4.064 26.676 4.096 29.184 ;
  LAYER M1 ;
        RECT 4 26.676 4.032 29.184 ;
  LAYER M2 ;
        RECT 3.884 26.76 6.356 26.792 ;
  LAYER M2 ;
        RECT 3.884 26.824 6.356 26.856 ;
  LAYER M2 ;
        RECT 3.884 26.888 6.356 26.92 ;
  LAYER M2 ;
        RECT 3.884 26.952 6.356 26.984 ;
  LAYER M2 ;
        RECT 3.884 27.016 6.356 27.048 ;
  LAYER M2 ;
        RECT 3.884 27.08 6.356 27.112 ;
  LAYER M2 ;
        RECT 3.884 27.144 6.356 27.176 ;
  LAYER M2 ;
        RECT 3.884 27.208 6.356 27.24 ;
  LAYER M2 ;
        RECT 3.884 27.272 6.356 27.304 ;
  LAYER M2 ;
        RECT 3.884 27.336 6.356 27.368 ;
  LAYER M2 ;
        RECT 3.884 27.4 6.356 27.432 ;
  LAYER M2 ;
        RECT 3.884 27.464 6.356 27.496 ;
  LAYER M2 ;
        RECT 3.884 27.528 6.356 27.56 ;
  LAYER M2 ;
        RECT 3.884 27.592 6.356 27.624 ;
  LAYER M2 ;
        RECT 3.884 27.656 6.356 27.688 ;
  LAYER M2 ;
        RECT 3.884 27.72 6.356 27.752 ;
  LAYER M2 ;
        RECT 3.884 27.784 6.356 27.816 ;
  LAYER M2 ;
        RECT 3.884 27.848 6.356 27.88 ;
  LAYER M2 ;
        RECT 3.884 27.912 6.356 27.944 ;
  LAYER M2 ;
        RECT 3.884 27.976 6.356 28.008 ;
  LAYER M2 ;
        RECT 3.884 28.04 6.356 28.072 ;
  LAYER M2 ;
        RECT 3.884 28.104 6.356 28.136 ;
  LAYER M2 ;
        RECT 3.884 28.168 6.356 28.2 ;
  LAYER M2 ;
        RECT 3.884 28.232 6.356 28.264 ;
  LAYER M2 ;
        RECT 3.884 28.296 6.356 28.328 ;
  LAYER M2 ;
        RECT 3.884 28.36 6.356 28.392 ;
  LAYER M2 ;
        RECT 3.884 28.424 6.356 28.456 ;
  LAYER M2 ;
        RECT 3.884 28.488 6.356 28.52 ;
  LAYER M2 ;
        RECT 3.884 28.552 6.356 28.584 ;
  LAYER M2 ;
        RECT 3.884 28.616 6.356 28.648 ;
  LAYER M2 ;
        RECT 3.884 28.68 6.356 28.712 ;
  LAYER M2 ;
        RECT 3.884 28.744 6.356 28.776 ;
  LAYER M2 ;
        RECT 3.884 28.808 6.356 28.84 ;
  LAYER M2 ;
        RECT 3.884 28.872 6.356 28.904 ;
  LAYER M2 ;
        RECT 3.884 28.936 6.356 28.968 ;
  LAYER M2 ;
        RECT 3.884 29 6.356 29.032 ;
  LAYER M3 ;
        RECT 6.304 26.676 6.336 29.184 ;
  LAYER M3 ;
        RECT 6.24 26.676 6.272 29.184 ;
  LAYER M3 ;
        RECT 6.176 26.676 6.208 29.184 ;
  LAYER M3 ;
        RECT 6.112 26.676 6.144 29.184 ;
  LAYER M3 ;
        RECT 6.048 26.676 6.08 29.184 ;
  LAYER M3 ;
        RECT 5.984 26.676 6.016 29.184 ;
  LAYER M3 ;
        RECT 5.92 26.676 5.952 29.184 ;
  LAYER M3 ;
        RECT 5.856 26.676 5.888 29.184 ;
  LAYER M3 ;
        RECT 5.792 26.676 5.824 29.184 ;
  LAYER M3 ;
        RECT 5.728 26.676 5.76 29.184 ;
  LAYER M3 ;
        RECT 5.664 26.676 5.696 29.184 ;
  LAYER M3 ;
        RECT 5.6 26.676 5.632 29.184 ;
  LAYER M3 ;
        RECT 5.536 26.676 5.568 29.184 ;
  LAYER M3 ;
        RECT 5.472 26.676 5.504 29.184 ;
  LAYER M3 ;
        RECT 5.408 26.676 5.44 29.184 ;
  LAYER M3 ;
        RECT 5.344 26.676 5.376 29.184 ;
  LAYER M3 ;
        RECT 5.28 26.676 5.312 29.184 ;
  LAYER M3 ;
        RECT 5.216 26.676 5.248 29.184 ;
  LAYER M3 ;
        RECT 5.152 26.676 5.184 29.184 ;
  LAYER M3 ;
        RECT 5.088 26.676 5.12 29.184 ;
  LAYER M3 ;
        RECT 5.024 26.676 5.056 29.184 ;
  LAYER M3 ;
        RECT 4.96 26.676 4.992 29.184 ;
  LAYER M3 ;
        RECT 4.896 26.676 4.928 29.184 ;
  LAYER M3 ;
        RECT 4.832 26.676 4.864 29.184 ;
  LAYER M3 ;
        RECT 4.768 26.676 4.8 29.184 ;
  LAYER M3 ;
        RECT 4.704 26.676 4.736 29.184 ;
  LAYER M3 ;
        RECT 4.64 26.676 4.672 29.184 ;
  LAYER M3 ;
        RECT 4.576 26.676 4.608 29.184 ;
  LAYER M3 ;
        RECT 4.512 26.676 4.544 29.184 ;
  LAYER M3 ;
        RECT 4.448 26.676 4.48 29.184 ;
  LAYER M3 ;
        RECT 4.384 26.676 4.416 29.184 ;
  LAYER M3 ;
        RECT 4.32 26.676 4.352 29.184 ;
  LAYER M3 ;
        RECT 4.256 26.676 4.288 29.184 ;
  LAYER M3 ;
        RECT 4.192 26.676 4.224 29.184 ;
  LAYER M3 ;
        RECT 4.128 26.676 4.16 29.184 ;
  LAYER M3 ;
        RECT 4.064 26.676 4.096 29.184 ;
  LAYER M3 ;
        RECT 4 26.676 4.032 29.184 ;
  LAYER M3 ;
        RECT 3.904 26.676 3.936 29.184 ;
  LAYER M1 ;
        RECT 6.319 26.712 6.321 29.148 ;
  LAYER M1 ;
        RECT 6.239 26.712 6.241 29.148 ;
  LAYER M1 ;
        RECT 6.159 26.712 6.161 29.148 ;
  LAYER M1 ;
        RECT 6.079 26.712 6.081 29.148 ;
  LAYER M1 ;
        RECT 5.999 26.712 6.001 29.148 ;
  LAYER M1 ;
        RECT 5.919 26.712 5.921 29.148 ;
  LAYER M1 ;
        RECT 5.839 26.712 5.841 29.148 ;
  LAYER M1 ;
        RECT 5.759 26.712 5.761 29.148 ;
  LAYER M1 ;
        RECT 5.679 26.712 5.681 29.148 ;
  LAYER M1 ;
        RECT 5.599 26.712 5.601 29.148 ;
  LAYER M1 ;
        RECT 5.519 26.712 5.521 29.148 ;
  LAYER M1 ;
        RECT 5.439 26.712 5.441 29.148 ;
  LAYER M1 ;
        RECT 5.359 26.712 5.361 29.148 ;
  LAYER M1 ;
        RECT 5.279 26.712 5.281 29.148 ;
  LAYER M1 ;
        RECT 5.199 26.712 5.201 29.148 ;
  LAYER M1 ;
        RECT 5.119 26.712 5.121 29.148 ;
  LAYER M1 ;
        RECT 5.039 26.712 5.041 29.148 ;
  LAYER M1 ;
        RECT 4.959 26.712 4.961 29.148 ;
  LAYER M1 ;
        RECT 4.879 26.712 4.881 29.148 ;
  LAYER M1 ;
        RECT 4.799 26.712 4.801 29.148 ;
  LAYER M1 ;
        RECT 4.719 26.712 4.721 29.148 ;
  LAYER M1 ;
        RECT 4.639 26.712 4.641 29.148 ;
  LAYER M1 ;
        RECT 4.559 26.712 4.561 29.148 ;
  LAYER M1 ;
        RECT 4.479 26.712 4.481 29.148 ;
  LAYER M1 ;
        RECT 4.399 26.712 4.401 29.148 ;
  LAYER M1 ;
        RECT 4.319 26.712 4.321 29.148 ;
  LAYER M1 ;
        RECT 4.239 26.712 4.241 29.148 ;
  LAYER M1 ;
        RECT 4.159 26.712 4.161 29.148 ;
  LAYER M1 ;
        RECT 4.079 26.712 4.081 29.148 ;
  LAYER M1 ;
        RECT 3.999 26.712 4.001 29.148 ;
  LAYER M2 ;
        RECT 3.92 26.711 6.32 26.713 ;
  LAYER M2 ;
        RECT 3.92 26.795 6.32 26.797 ;
  LAYER M2 ;
        RECT 3.92 26.879 6.32 26.881 ;
  LAYER M2 ;
        RECT 3.92 26.963 6.32 26.965 ;
  LAYER M2 ;
        RECT 3.92 27.047 6.32 27.049 ;
  LAYER M2 ;
        RECT 3.92 27.131 6.32 27.133 ;
  LAYER M2 ;
        RECT 3.92 27.215 6.32 27.217 ;
  LAYER M2 ;
        RECT 3.92 27.299 6.32 27.301 ;
  LAYER M2 ;
        RECT 3.92 27.383 6.32 27.385 ;
  LAYER M2 ;
        RECT 3.92 27.467 6.32 27.469 ;
  LAYER M2 ;
        RECT 3.92 27.551 6.32 27.553 ;
  LAYER M2 ;
        RECT 3.92 27.635 6.32 27.637 ;
  LAYER M2 ;
        RECT 3.92 27.7185 6.32 27.7205 ;
  LAYER M2 ;
        RECT 3.92 27.803 6.32 27.805 ;
  LAYER M2 ;
        RECT 3.92 27.887 6.32 27.889 ;
  LAYER M2 ;
        RECT 3.92 27.971 6.32 27.973 ;
  LAYER M2 ;
        RECT 3.92 28.055 6.32 28.057 ;
  LAYER M2 ;
        RECT 3.92 28.139 6.32 28.141 ;
  LAYER M2 ;
        RECT 3.92 28.223 6.32 28.225 ;
  LAYER M2 ;
        RECT 3.92 28.307 6.32 28.309 ;
  LAYER M2 ;
        RECT 3.92 28.391 6.32 28.393 ;
  LAYER M2 ;
        RECT 3.92 28.475 6.32 28.477 ;
  LAYER M2 ;
        RECT 3.92 28.559 6.32 28.561 ;
  LAYER M2 ;
        RECT 3.92 28.643 6.32 28.645 ;
  LAYER M2 ;
        RECT 3.92 28.727 6.32 28.729 ;
  LAYER M2 ;
        RECT 3.92 28.811 6.32 28.813 ;
  LAYER M2 ;
        RECT 3.92 28.895 6.32 28.897 ;
  LAYER M2 ;
        RECT 3.92 28.979 6.32 28.981 ;
  LAYER M2 ;
        RECT 3.92 29.063 6.32 29.065 ;
  LAYER M1 ;
        RECT 3.424 17.856 3.456 20.364 ;
  LAYER M1 ;
        RECT 3.36 17.856 3.392 20.364 ;
  LAYER M1 ;
        RECT 3.296 17.856 3.328 20.364 ;
  LAYER M1 ;
        RECT 3.232 17.856 3.264 20.364 ;
  LAYER M1 ;
        RECT 3.168 17.856 3.2 20.364 ;
  LAYER M1 ;
        RECT 3.104 17.856 3.136 20.364 ;
  LAYER M1 ;
        RECT 3.04 17.856 3.072 20.364 ;
  LAYER M1 ;
        RECT 2.976 17.856 3.008 20.364 ;
  LAYER M1 ;
        RECT 2.912 17.856 2.944 20.364 ;
  LAYER M1 ;
        RECT 2.848 17.856 2.88 20.364 ;
  LAYER M1 ;
        RECT 2.784 17.856 2.816 20.364 ;
  LAYER M1 ;
        RECT 2.72 17.856 2.752 20.364 ;
  LAYER M1 ;
        RECT 2.656 17.856 2.688 20.364 ;
  LAYER M1 ;
        RECT 2.592 17.856 2.624 20.364 ;
  LAYER M1 ;
        RECT 2.528 17.856 2.56 20.364 ;
  LAYER M1 ;
        RECT 2.464 17.856 2.496 20.364 ;
  LAYER M1 ;
        RECT 2.4 17.856 2.432 20.364 ;
  LAYER M1 ;
        RECT 2.336 17.856 2.368 20.364 ;
  LAYER M1 ;
        RECT 2.272 17.856 2.304 20.364 ;
  LAYER M1 ;
        RECT 2.208 17.856 2.24 20.364 ;
  LAYER M1 ;
        RECT 2.144 17.856 2.176 20.364 ;
  LAYER M1 ;
        RECT 2.08 17.856 2.112 20.364 ;
  LAYER M1 ;
        RECT 2.016 17.856 2.048 20.364 ;
  LAYER M1 ;
        RECT 1.952 17.856 1.984 20.364 ;
  LAYER M1 ;
        RECT 1.888 17.856 1.92 20.364 ;
  LAYER M1 ;
        RECT 1.824 17.856 1.856 20.364 ;
  LAYER M1 ;
        RECT 1.76 17.856 1.792 20.364 ;
  LAYER M1 ;
        RECT 1.696 17.856 1.728 20.364 ;
  LAYER M1 ;
        RECT 1.632 17.856 1.664 20.364 ;
  LAYER M1 ;
        RECT 1.568 17.856 1.6 20.364 ;
  LAYER M1 ;
        RECT 1.504 17.856 1.536 20.364 ;
  LAYER M1 ;
        RECT 1.44 17.856 1.472 20.364 ;
  LAYER M1 ;
        RECT 1.376 17.856 1.408 20.364 ;
  LAYER M1 ;
        RECT 1.312 17.856 1.344 20.364 ;
  LAYER M1 ;
        RECT 1.248 17.856 1.28 20.364 ;
  LAYER M1 ;
        RECT 1.184 17.856 1.216 20.364 ;
  LAYER M1 ;
        RECT 1.12 17.856 1.152 20.364 ;
  LAYER M2 ;
        RECT 1.004 17.94 3.476 17.972 ;
  LAYER M2 ;
        RECT 1.004 18.004 3.476 18.036 ;
  LAYER M2 ;
        RECT 1.004 18.068 3.476 18.1 ;
  LAYER M2 ;
        RECT 1.004 18.132 3.476 18.164 ;
  LAYER M2 ;
        RECT 1.004 18.196 3.476 18.228 ;
  LAYER M2 ;
        RECT 1.004 18.26 3.476 18.292 ;
  LAYER M2 ;
        RECT 1.004 18.324 3.476 18.356 ;
  LAYER M2 ;
        RECT 1.004 18.388 3.476 18.42 ;
  LAYER M2 ;
        RECT 1.004 18.452 3.476 18.484 ;
  LAYER M2 ;
        RECT 1.004 18.516 3.476 18.548 ;
  LAYER M2 ;
        RECT 1.004 18.58 3.476 18.612 ;
  LAYER M2 ;
        RECT 1.004 18.644 3.476 18.676 ;
  LAYER M2 ;
        RECT 1.004 18.708 3.476 18.74 ;
  LAYER M2 ;
        RECT 1.004 18.772 3.476 18.804 ;
  LAYER M2 ;
        RECT 1.004 18.836 3.476 18.868 ;
  LAYER M2 ;
        RECT 1.004 18.9 3.476 18.932 ;
  LAYER M2 ;
        RECT 1.004 18.964 3.476 18.996 ;
  LAYER M2 ;
        RECT 1.004 19.028 3.476 19.06 ;
  LAYER M2 ;
        RECT 1.004 19.092 3.476 19.124 ;
  LAYER M2 ;
        RECT 1.004 19.156 3.476 19.188 ;
  LAYER M2 ;
        RECT 1.004 19.22 3.476 19.252 ;
  LAYER M2 ;
        RECT 1.004 19.284 3.476 19.316 ;
  LAYER M2 ;
        RECT 1.004 19.348 3.476 19.38 ;
  LAYER M2 ;
        RECT 1.004 19.412 3.476 19.444 ;
  LAYER M2 ;
        RECT 1.004 19.476 3.476 19.508 ;
  LAYER M2 ;
        RECT 1.004 19.54 3.476 19.572 ;
  LAYER M2 ;
        RECT 1.004 19.604 3.476 19.636 ;
  LAYER M2 ;
        RECT 1.004 19.668 3.476 19.7 ;
  LAYER M2 ;
        RECT 1.004 19.732 3.476 19.764 ;
  LAYER M2 ;
        RECT 1.004 19.796 3.476 19.828 ;
  LAYER M2 ;
        RECT 1.004 19.86 3.476 19.892 ;
  LAYER M2 ;
        RECT 1.004 19.924 3.476 19.956 ;
  LAYER M2 ;
        RECT 1.004 19.988 3.476 20.02 ;
  LAYER M2 ;
        RECT 1.004 20.052 3.476 20.084 ;
  LAYER M2 ;
        RECT 1.004 20.116 3.476 20.148 ;
  LAYER M2 ;
        RECT 1.004 20.18 3.476 20.212 ;
  LAYER M3 ;
        RECT 3.424 17.856 3.456 20.364 ;
  LAYER M3 ;
        RECT 3.36 17.856 3.392 20.364 ;
  LAYER M3 ;
        RECT 3.296 17.856 3.328 20.364 ;
  LAYER M3 ;
        RECT 3.232 17.856 3.264 20.364 ;
  LAYER M3 ;
        RECT 3.168 17.856 3.2 20.364 ;
  LAYER M3 ;
        RECT 3.104 17.856 3.136 20.364 ;
  LAYER M3 ;
        RECT 3.04 17.856 3.072 20.364 ;
  LAYER M3 ;
        RECT 2.976 17.856 3.008 20.364 ;
  LAYER M3 ;
        RECT 2.912 17.856 2.944 20.364 ;
  LAYER M3 ;
        RECT 2.848 17.856 2.88 20.364 ;
  LAYER M3 ;
        RECT 2.784 17.856 2.816 20.364 ;
  LAYER M3 ;
        RECT 2.72 17.856 2.752 20.364 ;
  LAYER M3 ;
        RECT 2.656 17.856 2.688 20.364 ;
  LAYER M3 ;
        RECT 2.592 17.856 2.624 20.364 ;
  LAYER M3 ;
        RECT 2.528 17.856 2.56 20.364 ;
  LAYER M3 ;
        RECT 2.464 17.856 2.496 20.364 ;
  LAYER M3 ;
        RECT 2.4 17.856 2.432 20.364 ;
  LAYER M3 ;
        RECT 2.336 17.856 2.368 20.364 ;
  LAYER M3 ;
        RECT 2.272 17.856 2.304 20.364 ;
  LAYER M3 ;
        RECT 2.208 17.856 2.24 20.364 ;
  LAYER M3 ;
        RECT 2.144 17.856 2.176 20.364 ;
  LAYER M3 ;
        RECT 2.08 17.856 2.112 20.364 ;
  LAYER M3 ;
        RECT 2.016 17.856 2.048 20.364 ;
  LAYER M3 ;
        RECT 1.952 17.856 1.984 20.364 ;
  LAYER M3 ;
        RECT 1.888 17.856 1.92 20.364 ;
  LAYER M3 ;
        RECT 1.824 17.856 1.856 20.364 ;
  LAYER M3 ;
        RECT 1.76 17.856 1.792 20.364 ;
  LAYER M3 ;
        RECT 1.696 17.856 1.728 20.364 ;
  LAYER M3 ;
        RECT 1.632 17.856 1.664 20.364 ;
  LAYER M3 ;
        RECT 1.568 17.856 1.6 20.364 ;
  LAYER M3 ;
        RECT 1.504 17.856 1.536 20.364 ;
  LAYER M3 ;
        RECT 1.44 17.856 1.472 20.364 ;
  LAYER M3 ;
        RECT 1.376 17.856 1.408 20.364 ;
  LAYER M3 ;
        RECT 1.312 17.856 1.344 20.364 ;
  LAYER M3 ;
        RECT 1.248 17.856 1.28 20.364 ;
  LAYER M3 ;
        RECT 1.184 17.856 1.216 20.364 ;
  LAYER M3 ;
        RECT 1.12 17.856 1.152 20.364 ;
  LAYER M3 ;
        RECT 1.024 17.856 1.056 20.364 ;
  LAYER M1 ;
        RECT 3.439 17.892 3.441 20.328 ;
  LAYER M1 ;
        RECT 3.359 17.892 3.361 20.328 ;
  LAYER M1 ;
        RECT 3.279 17.892 3.281 20.328 ;
  LAYER M1 ;
        RECT 3.199 17.892 3.201 20.328 ;
  LAYER M1 ;
        RECT 3.119 17.892 3.121 20.328 ;
  LAYER M1 ;
        RECT 3.039 17.892 3.041 20.328 ;
  LAYER M1 ;
        RECT 2.959 17.892 2.961 20.328 ;
  LAYER M1 ;
        RECT 2.879 17.892 2.881 20.328 ;
  LAYER M1 ;
        RECT 2.799 17.892 2.801 20.328 ;
  LAYER M1 ;
        RECT 2.719 17.892 2.721 20.328 ;
  LAYER M1 ;
        RECT 2.639 17.892 2.641 20.328 ;
  LAYER M1 ;
        RECT 2.559 17.892 2.561 20.328 ;
  LAYER M1 ;
        RECT 2.479 17.892 2.481 20.328 ;
  LAYER M1 ;
        RECT 2.399 17.892 2.401 20.328 ;
  LAYER M1 ;
        RECT 2.319 17.892 2.321 20.328 ;
  LAYER M1 ;
        RECT 2.239 17.892 2.241 20.328 ;
  LAYER M1 ;
        RECT 2.159 17.892 2.161 20.328 ;
  LAYER M1 ;
        RECT 2.079 17.892 2.081 20.328 ;
  LAYER M1 ;
        RECT 1.999 17.892 2.001 20.328 ;
  LAYER M1 ;
        RECT 1.919 17.892 1.921 20.328 ;
  LAYER M1 ;
        RECT 1.839 17.892 1.841 20.328 ;
  LAYER M1 ;
        RECT 1.759 17.892 1.761 20.328 ;
  LAYER M1 ;
        RECT 1.679 17.892 1.681 20.328 ;
  LAYER M1 ;
        RECT 1.599 17.892 1.601 20.328 ;
  LAYER M1 ;
        RECT 1.519 17.892 1.521 20.328 ;
  LAYER M1 ;
        RECT 1.439 17.892 1.441 20.328 ;
  LAYER M1 ;
        RECT 1.359 17.892 1.361 20.328 ;
  LAYER M1 ;
        RECT 1.279 17.892 1.281 20.328 ;
  LAYER M1 ;
        RECT 1.199 17.892 1.201 20.328 ;
  LAYER M1 ;
        RECT 1.119 17.892 1.121 20.328 ;
  LAYER M2 ;
        RECT 1.04 17.891 3.44 17.893 ;
  LAYER M2 ;
        RECT 1.04 17.975 3.44 17.977 ;
  LAYER M2 ;
        RECT 1.04 18.059 3.44 18.061 ;
  LAYER M2 ;
        RECT 1.04 18.143 3.44 18.145 ;
  LAYER M2 ;
        RECT 1.04 18.227 3.44 18.229 ;
  LAYER M2 ;
        RECT 1.04 18.311 3.44 18.313 ;
  LAYER M2 ;
        RECT 1.04 18.395 3.44 18.397 ;
  LAYER M2 ;
        RECT 1.04 18.479 3.44 18.481 ;
  LAYER M2 ;
        RECT 1.04 18.563 3.44 18.565 ;
  LAYER M2 ;
        RECT 1.04 18.647 3.44 18.649 ;
  LAYER M2 ;
        RECT 1.04 18.731 3.44 18.733 ;
  LAYER M2 ;
        RECT 1.04 18.815 3.44 18.817 ;
  LAYER M2 ;
        RECT 1.04 18.8985 3.44 18.9005 ;
  LAYER M2 ;
        RECT 1.04 18.983 3.44 18.985 ;
  LAYER M2 ;
        RECT 1.04 19.067 3.44 19.069 ;
  LAYER M2 ;
        RECT 1.04 19.151 3.44 19.153 ;
  LAYER M2 ;
        RECT 1.04 19.235 3.44 19.237 ;
  LAYER M2 ;
        RECT 1.04 19.319 3.44 19.321 ;
  LAYER M2 ;
        RECT 1.04 19.403 3.44 19.405 ;
  LAYER M2 ;
        RECT 1.04 19.487 3.44 19.489 ;
  LAYER M2 ;
        RECT 1.04 19.571 3.44 19.573 ;
  LAYER M2 ;
        RECT 1.04 19.655 3.44 19.657 ;
  LAYER M2 ;
        RECT 1.04 19.739 3.44 19.741 ;
  LAYER M2 ;
        RECT 1.04 19.823 3.44 19.825 ;
  LAYER M2 ;
        RECT 1.04 19.907 3.44 19.909 ;
  LAYER M2 ;
        RECT 1.04 19.991 3.44 19.993 ;
  LAYER M2 ;
        RECT 1.04 20.075 3.44 20.077 ;
  LAYER M2 ;
        RECT 1.04 20.159 3.44 20.161 ;
  LAYER M2 ;
        RECT 1.04 20.243 3.44 20.245 ;
  LAYER M1 ;
        RECT 3.424 20.796 3.456 23.304 ;
  LAYER M1 ;
        RECT 3.36 20.796 3.392 23.304 ;
  LAYER M1 ;
        RECT 3.296 20.796 3.328 23.304 ;
  LAYER M1 ;
        RECT 3.232 20.796 3.264 23.304 ;
  LAYER M1 ;
        RECT 3.168 20.796 3.2 23.304 ;
  LAYER M1 ;
        RECT 3.104 20.796 3.136 23.304 ;
  LAYER M1 ;
        RECT 3.04 20.796 3.072 23.304 ;
  LAYER M1 ;
        RECT 2.976 20.796 3.008 23.304 ;
  LAYER M1 ;
        RECT 2.912 20.796 2.944 23.304 ;
  LAYER M1 ;
        RECT 2.848 20.796 2.88 23.304 ;
  LAYER M1 ;
        RECT 2.784 20.796 2.816 23.304 ;
  LAYER M1 ;
        RECT 2.72 20.796 2.752 23.304 ;
  LAYER M1 ;
        RECT 2.656 20.796 2.688 23.304 ;
  LAYER M1 ;
        RECT 2.592 20.796 2.624 23.304 ;
  LAYER M1 ;
        RECT 2.528 20.796 2.56 23.304 ;
  LAYER M1 ;
        RECT 2.464 20.796 2.496 23.304 ;
  LAYER M1 ;
        RECT 2.4 20.796 2.432 23.304 ;
  LAYER M1 ;
        RECT 2.336 20.796 2.368 23.304 ;
  LAYER M1 ;
        RECT 2.272 20.796 2.304 23.304 ;
  LAYER M1 ;
        RECT 2.208 20.796 2.24 23.304 ;
  LAYER M1 ;
        RECT 2.144 20.796 2.176 23.304 ;
  LAYER M1 ;
        RECT 2.08 20.796 2.112 23.304 ;
  LAYER M1 ;
        RECT 2.016 20.796 2.048 23.304 ;
  LAYER M1 ;
        RECT 1.952 20.796 1.984 23.304 ;
  LAYER M1 ;
        RECT 1.888 20.796 1.92 23.304 ;
  LAYER M1 ;
        RECT 1.824 20.796 1.856 23.304 ;
  LAYER M1 ;
        RECT 1.76 20.796 1.792 23.304 ;
  LAYER M1 ;
        RECT 1.696 20.796 1.728 23.304 ;
  LAYER M1 ;
        RECT 1.632 20.796 1.664 23.304 ;
  LAYER M1 ;
        RECT 1.568 20.796 1.6 23.304 ;
  LAYER M1 ;
        RECT 1.504 20.796 1.536 23.304 ;
  LAYER M1 ;
        RECT 1.44 20.796 1.472 23.304 ;
  LAYER M1 ;
        RECT 1.376 20.796 1.408 23.304 ;
  LAYER M1 ;
        RECT 1.312 20.796 1.344 23.304 ;
  LAYER M1 ;
        RECT 1.248 20.796 1.28 23.304 ;
  LAYER M1 ;
        RECT 1.184 20.796 1.216 23.304 ;
  LAYER M1 ;
        RECT 1.12 20.796 1.152 23.304 ;
  LAYER M2 ;
        RECT 1.004 20.88 3.476 20.912 ;
  LAYER M2 ;
        RECT 1.004 20.944 3.476 20.976 ;
  LAYER M2 ;
        RECT 1.004 21.008 3.476 21.04 ;
  LAYER M2 ;
        RECT 1.004 21.072 3.476 21.104 ;
  LAYER M2 ;
        RECT 1.004 21.136 3.476 21.168 ;
  LAYER M2 ;
        RECT 1.004 21.2 3.476 21.232 ;
  LAYER M2 ;
        RECT 1.004 21.264 3.476 21.296 ;
  LAYER M2 ;
        RECT 1.004 21.328 3.476 21.36 ;
  LAYER M2 ;
        RECT 1.004 21.392 3.476 21.424 ;
  LAYER M2 ;
        RECT 1.004 21.456 3.476 21.488 ;
  LAYER M2 ;
        RECT 1.004 21.52 3.476 21.552 ;
  LAYER M2 ;
        RECT 1.004 21.584 3.476 21.616 ;
  LAYER M2 ;
        RECT 1.004 21.648 3.476 21.68 ;
  LAYER M2 ;
        RECT 1.004 21.712 3.476 21.744 ;
  LAYER M2 ;
        RECT 1.004 21.776 3.476 21.808 ;
  LAYER M2 ;
        RECT 1.004 21.84 3.476 21.872 ;
  LAYER M2 ;
        RECT 1.004 21.904 3.476 21.936 ;
  LAYER M2 ;
        RECT 1.004 21.968 3.476 22 ;
  LAYER M2 ;
        RECT 1.004 22.032 3.476 22.064 ;
  LAYER M2 ;
        RECT 1.004 22.096 3.476 22.128 ;
  LAYER M2 ;
        RECT 1.004 22.16 3.476 22.192 ;
  LAYER M2 ;
        RECT 1.004 22.224 3.476 22.256 ;
  LAYER M2 ;
        RECT 1.004 22.288 3.476 22.32 ;
  LAYER M2 ;
        RECT 1.004 22.352 3.476 22.384 ;
  LAYER M2 ;
        RECT 1.004 22.416 3.476 22.448 ;
  LAYER M2 ;
        RECT 1.004 22.48 3.476 22.512 ;
  LAYER M2 ;
        RECT 1.004 22.544 3.476 22.576 ;
  LAYER M2 ;
        RECT 1.004 22.608 3.476 22.64 ;
  LAYER M2 ;
        RECT 1.004 22.672 3.476 22.704 ;
  LAYER M2 ;
        RECT 1.004 22.736 3.476 22.768 ;
  LAYER M2 ;
        RECT 1.004 22.8 3.476 22.832 ;
  LAYER M2 ;
        RECT 1.004 22.864 3.476 22.896 ;
  LAYER M2 ;
        RECT 1.004 22.928 3.476 22.96 ;
  LAYER M2 ;
        RECT 1.004 22.992 3.476 23.024 ;
  LAYER M2 ;
        RECT 1.004 23.056 3.476 23.088 ;
  LAYER M2 ;
        RECT 1.004 23.12 3.476 23.152 ;
  LAYER M3 ;
        RECT 3.424 20.796 3.456 23.304 ;
  LAYER M3 ;
        RECT 3.36 20.796 3.392 23.304 ;
  LAYER M3 ;
        RECT 3.296 20.796 3.328 23.304 ;
  LAYER M3 ;
        RECT 3.232 20.796 3.264 23.304 ;
  LAYER M3 ;
        RECT 3.168 20.796 3.2 23.304 ;
  LAYER M3 ;
        RECT 3.104 20.796 3.136 23.304 ;
  LAYER M3 ;
        RECT 3.04 20.796 3.072 23.304 ;
  LAYER M3 ;
        RECT 2.976 20.796 3.008 23.304 ;
  LAYER M3 ;
        RECT 2.912 20.796 2.944 23.304 ;
  LAYER M3 ;
        RECT 2.848 20.796 2.88 23.304 ;
  LAYER M3 ;
        RECT 2.784 20.796 2.816 23.304 ;
  LAYER M3 ;
        RECT 2.72 20.796 2.752 23.304 ;
  LAYER M3 ;
        RECT 2.656 20.796 2.688 23.304 ;
  LAYER M3 ;
        RECT 2.592 20.796 2.624 23.304 ;
  LAYER M3 ;
        RECT 2.528 20.796 2.56 23.304 ;
  LAYER M3 ;
        RECT 2.464 20.796 2.496 23.304 ;
  LAYER M3 ;
        RECT 2.4 20.796 2.432 23.304 ;
  LAYER M3 ;
        RECT 2.336 20.796 2.368 23.304 ;
  LAYER M3 ;
        RECT 2.272 20.796 2.304 23.304 ;
  LAYER M3 ;
        RECT 2.208 20.796 2.24 23.304 ;
  LAYER M3 ;
        RECT 2.144 20.796 2.176 23.304 ;
  LAYER M3 ;
        RECT 2.08 20.796 2.112 23.304 ;
  LAYER M3 ;
        RECT 2.016 20.796 2.048 23.304 ;
  LAYER M3 ;
        RECT 1.952 20.796 1.984 23.304 ;
  LAYER M3 ;
        RECT 1.888 20.796 1.92 23.304 ;
  LAYER M3 ;
        RECT 1.824 20.796 1.856 23.304 ;
  LAYER M3 ;
        RECT 1.76 20.796 1.792 23.304 ;
  LAYER M3 ;
        RECT 1.696 20.796 1.728 23.304 ;
  LAYER M3 ;
        RECT 1.632 20.796 1.664 23.304 ;
  LAYER M3 ;
        RECT 1.568 20.796 1.6 23.304 ;
  LAYER M3 ;
        RECT 1.504 20.796 1.536 23.304 ;
  LAYER M3 ;
        RECT 1.44 20.796 1.472 23.304 ;
  LAYER M3 ;
        RECT 1.376 20.796 1.408 23.304 ;
  LAYER M3 ;
        RECT 1.312 20.796 1.344 23.304 ;
  LAYER M3 ;
        RECT 1.248 20.796 1.28 23.304 ;
  LAYER M3 ;
        RECT 1.184 20.796 1.216 23.304 ;
  LAYER M3 ;
        RECT 1.12 20.796 1.152 23.304 ;
  LAYER M3 ;
        RECT 1.024 20.796 1.056 23.304 ;
  LAYER M1 ;
        RECT 3.439 20.832 3.441 23.268 ;
  LAYER M1 ;
        RECT 3.359 20.832 3.361 23.268 ;
  LAYER M1 ;
        RECT 3.279 20.832 3.281 23.268 ;
  LAYER M1 ;
        RECT 3.199 20.832 3.201 23.268 ;
  LAYER M1 ;
        RECT 3.119 20.832 3.121 23.268 ;
  LAYER M1 ;
        RECT 3.039 20.832 3.041 23.268 ;
  LAYER M1 ;
        RECT 2.959 20.832 2.961 23.268 ;
  LAYER M1 ;
        RECT 2.879 20.832 2.881 23.268 ;
  LAYER M1 ;
        RECT 2.799 20.832 2.801 23.268 ;
  LAYER M1 ;
        RECT 2.719 20.832 2.721 23.268 ;
  LAYER M1 ;
        RECT 2.639 20.832 2.641 23.268 ;
  LAYER M1 ;
        RECT 2.559 20.832 2.561 23.268 ;
  LAYER M1 ;
        RECT 2.479 20.832 2.481 23.268 ;
  LAYER M1 ;
        RECT 2.399 20.832 2.401 23.268 ;
  LAYER M1 ;
        RECT 2.319 20.832 2.321 23.268 ;
  LAYER M1 ;
        RECT 2.239 20.832 2.241 23.268 ;
  LAYER M1 ;
        RECT 2.159 20.832 2.161 23.268 ;
  LAYER M1 ;
        RECT 2.079 20.832 2.081 23.268 ;
  LAYER M1 ;
        RECT 1.999 20.832 2.001 23.268 ;
  LAYER M1 ;
        RECT 1.919 20.832 1.921 23.268 ;
  LAYER M1 ;
        RECT 1.839 20.832 1.841 23.268 ;
  LAYER M1 ;
        RECT 1.759 20.832 1.761 23.268 ;
  LAYER M1 ;
        RECT 1.679 20.832 1.681 23.268 ;
  LAYER M1 ;
        RECT 1.599 20.832 1.601 23.268 ;
  LAYER M1 ;
        RECT 1.519 20.832 1.521 23.268 ;
  LAYER M1 ;
        RECT 1.439 20.832 1.441 23.268 ;
  LAYER M1 ;
        RECT 1.359 20.832 1.361 23.268 ;
  LAYER M1 ;
        RECT 1.279 20.832 1.281 23.268 ;
  LAYER M1 ;
        RECT 1.199 20.832 1.201 23.268 ;
  LAYER M1 ;
        RECT 1.119 20.832 1.121 23.268 ;
  LAYER M2 ;
        RECT 1.04 20.831 3.44 20.833 ;
  LAYER M2 ;
        RECT 1.04 20.915 3.44 20.917 ;
  LAYER M2 ;
        RECT 1.04 20.999 3.44 21.001 ;
  LAYER M2 ;
        RECT 1.04 21.083 3.44 21.085 ;
  LAYER M2 ;
        RECT 1.04 21.167 3.44 21.169 ;
  LAYER M2 ;
        RECT 1.04 21.251 3.44 21.253 ;
  LAYER M2 ;
        RECT 1.04 21.335 3.44 21.337 ;
  LAYER M2 ;
        RECT 1.04 21.419 3.44 21.421 ;
  LAYER M2 ;
        RECT 1.04 21.503 3.44 21.505 ;
  LAYER M2 ;
        RECT 1.04 21.587 3.44 21.589 ;
  LAYER M2 ;
        RECT 1.04 21.671 3.44 21.673 ;
  LAYER M2 ;
        RECT 1.04 21.755 3.44 21.757 ;
  LAYER M2 ;
        RECT 1.04 21.8385 3.44 21.8405 ;
  LAYER M2 ;
        RECT 1.04 21.923 3.44 21.925 ;
  LAYER M2 ;
        RECT 1.04 22.007 3.44 22.009 ;
  LAYER M2 ;
        RECT 1.04 22.091 3.44 22.093 ;
  LAYER M2 ;
        RECT 1.04 22.175 3.44 22.177 ;
  LAYER M2 ;
        RECT 1.04 22.259 3.44 22.261 ;
  LAYER M2 ;
        RECT 1.04 22.343 3.44 22.345 ;
  LAYER M2 ;
        RECT 1.04 22.427 3.44 22.429 ;
  LAYER M2 ;
        RECT 1.04 22.511 3.44 22.513 ;
  LAYER M2 ;
        RECT 1.04 22.595 3.44 22.597 ;
  LAYER M2 ;
        RECT 1.04 22.679 3.44 22.681 ;
  LAYER M2 ;
        RECT 1.04 22.763 3.44 22.765 ;
  LAYER M2 ;
        RECT 1.04 22.847 3.44 22.849 ;
  LAYER M2 ;
        RECT 1.04 22.931 3.44 22.933 ;
  LAYER M2 ;
        RECT 1.04 23.015 3.44 23.017 ;
  LAYER M2 ;
        RECT 1.04 23.099 3.44 23.101 ;
  LAYER M2 ;
        RECT 1.04 23.183 3.44 23.185 ;
  LAYER M1 ;
        RECT 3.424 23.736 3.456 26.244 ;
  LAYER M1 ;
        RECT 3.36 23.736 3.392 26.244 ;
  LAYER M1 ;
        RECT 3.296 23.736 3.328 26.244 ;
  LAYER M1 ;
        RECT 3.232 23.736 3.264 26.244 ;
  LAYER M1 ;
        RECT 3.168 23.736 3.2 26.244 ;
  LAYER M1 ;
        RECT 3.104 23.736 3.136 26.244 ;
  LAYER M1 ;
        RECT 3.04 23.736 3.072 26.244 ;
  LAYER M1 ;
        RECT 2.976 23.736 3.008 26.244 ;
  LAYER M1 ;
        RECT 2.912 23.736 2.944 26.244 ;
  LAYER M1 ;
        RECT 2.848 23.736 2.88 26.244 ;
  LAYER M1 ;
        RECT 2.784 23.736 2.816 26.244 ;
  LAYER M1 ;
        RECT 2.72 23.736 2.752 26.244 ;
  LAYER M1 ;
        RECT 2.656 23.736 2.688 26.244 ;
  LAYER M1 ;
        RECT 2.592 23.736 2.624 26.244 ;
  LAYER M1 ;
        RECT 2.528 23.736 2.56 26.244 ;
  LAYER M1 ;
        RECT 2.464 23.736 2.496 26.244 ;
  LAYER M1 ;
        RECT 2.4 23.736 2.432 26.244 ;
  LAYER M1 ;
        RECT 2.336 23.736 2.368 26.244 ;
  LAYER M1 ;
        RECT 2.272 23.736 2.304 26.244 ;
  LAYER M1 ;
        RECT 2.208 23.736 2.24 26.244 ;
  LAYER M1 ;
        RECT 2.144 23.736 2.176 26.244 ;
  LAYER M1 ;
        RECT 2.08 23.736 2.112 26.244 ;
  LAYER M1 ;
        RECT 2.016 23.736 2.048 26.244 ;
  LAYER M1 ;
        RECT 1.952 23.736 1.984 26.244 ;
  LAYER M1 ;
        RECT 1.888 23.736 1.92 26.244 ;
  LAYER M1 ;
        RECT 1.824 23.736 1.856 26.244 ;
  LAYER M1 ;
        RECT 1.76 23.736 1.792 26.244 ;
  LAYER M1 ;
        RECT 1.696 23.736 1.728 26.244 ;
  LAYER M1 ;
        RECT 1.632 23.736 1.664 26.244 ;
  LAYER M1 ;
        RECT 1.568 23.736 1.6 26.244 ;
  LAYER M1 ;
        RECT 1.504 23.736 1.536 26.244 ;
  LAYER M1 ;
        RECT 1.44 23.736 1.472 26.244 ;
  LAYER M1 ;
        RECT 1.376 23.736 1.408 26.244 ;
  LAYER M1 ;
        RECT 1.312 23.736 1.344 26.244 ;
  LAYER M1 ;
        RECT 1.248 23.736 1.28 26.244 ;
  LAYER M1 ;
        RECT 1.184 23.736 1.216 26.244 ;
  LAYER M1 ;
        RECT 1.12 23.736 1.152 26.244 ;
  LAYER M2 ;
        RECT 1.004 23.82 3.476 23.852 ;
  LAYER M2 ;
        RECT 1.004 23.884 3.476 23.916 ;
  LAYER M2 ;
        RECT 1.004 23.948 3.476 23.98 ;
  LAYER M2 ;
        RECT 1.004 24.012 3.476 24.044 ;
  LAYER M2 ;
        RECT 1.004 24.076 3.476 24.108 ;
  LAYER M2 ;
        RECT 1.004 24.14 3.476 24.172 ;
  LAYER M2 ;
        RECT 1.004 24.204 3.476 24.236 ;
  LAYER M2 ;
        RECT 1.004 24.268 3.476 24.3 ;
  LAYER M2 ;
        RECT 1.004 24.332 3.476 24.364 ;
  LAYER M2 ;
        RECT 1.004 24.396 3.476 24.428 ;
  LAYER M2 ;
        RECT 1.004 24.46 3.476 24.492 ;
  LAYER M2 ;
        RECT 1.004 24.524 3.476 24.556 ;
  LAYER M2 ;
        RECT 1.004 24.588 3.476 24.62 ;
  LAYER M2 ;
        RECT 1.004 24.652 3.476 24.684 ;
  LAYER M2 ;
        RECT 1.004 24.716 3.476 24.748 ;
  LAYER M2 ;
        RECT 1.004 24.78 3.476 24.812 ;
  LAYER M2 ;
        RECT 1.004 24.844 3.476 24.876 ;
  LAYER M2 ;
        RECT 1.004 24.908 3.476 24.94 ;
  LAYER M2 ;
        RECT 1.004 24.972 3.476 25.004 ;
  LAYER M2 ;
        RECT 1.004 25.036 3.476 25.068 ;
  LAYER M2 ;
        RECT 1.004 25.1 3.476 25.132 ;
  LAYER M2 ;
        RECT 1.004 25.164 3.476 25.196 ;
  LAYER M2 ;
        RECT 1.004 25.228 3.476 25.26 ;
  LAYER M2 ;
        RECT 1.004 25.292 3.476 25.324 ;
  LAYER M2 ;
        RECT 1.004 25.356 3.476 25.388 ;
  LAYER M2 ;
        RECT 1.004 25.42 3.476 25.452 ;
  LAYER M2 ;
        RECT 1.004 25.484 3.476 25.516 ;
  LAYER M2 ;
        RECT 1.004 25.548 3.476 25.58 ;
  LAYER M2 ;
        RECT 1.004 25.612 3.476 25.644 ;
  LAYER M2 ;
        RECT 1.004 25.676 3.476 25.708 ;
  LAYER M2 ;
        RECT 1.004 25.74 3.476 25.772 ;
  LAYER M2 ;
        RECT 1.004 25.804 3.476 25.836 ;
  LAYER M2 ;
        RECT 1.004 25.868 3.476 25.9 ;
  LAYER M2 ;
        RECT 1.004 25.932 3.476 25.964 ;
  LAYER M2 ;
        RECT 1.004 25.996 3.476 26.028 ;
  LAYER M2 ;
        RECT 1.004 26.06 3.476 26.092 ;
  LAYER M3 ;
        RECT 3.424 23.736 3.456 26.244 ;
  LAYER M3 ;
        RECT 3.36 23.736 3.392 26.244 ;
  LAYER M3 ;
        RECT 3.296 23.736 3.328 26.244 ;
  LAYER M3 ;
        RECT 3.232 23.736 3.264 26.244 ;
  LAYER M3 ;
        RECT 3.168 23.736 3.2 26.244 ;
  LAYER M3 ;
        RECT 3.104 23.736 3.136 26.244 ;
  LAYER M3 ;
        RECT 3.04 23.736 3.072 26.244 ;
  LAYER M3 ;
        RECT 2.976 23.736 3.008 26.244 ;
  LAYER M3 ;
        RECT 2.912 23.736 2.944 26.244 ;
  LAYER M3 ;
        RECT 2.848 23.736 2.88 26.244 ;
  LAYER M3 ;
        RECT 2.784 23.736 2.816 26.244 ;
  LAYER M3 ;
        RECT 2.72 23.736 2.752 26.244 ;
  LAYER M3 ;
        RECT 2.656 23.736 2.688 26.244 ;
  LAYER M3 ;
        RECT 2.592 23.736 2.624 26.244 ;
  LAYER M3 ;
        RECT 2.528 23.736 2.56 26.244 ;
  LAYER M3 ;
        RECT 2.464 23.736 2.496 26.244 ;
  LAYER M3 ;
        RECT 2.4 23.736 2.432 26.244 ;
  LAYER M3 ;
        RECT 2.336 23.736 2.368 26.244 ;
  LAYER M3 ;
        RECT 2.272 23.736 2.304 26.244 ;
  LAYER M3 ;
        RECT 2.208 23.736 2.24 26.244 ;
  LAYER M3 ;
        RECT 2.144 23.736 2.176 26.244 ;
  LAYER M3 ;
        RECT 2.08 23.736 2.112 26.244 ;
  LAYER M3 ;
        RECT 2.016 23.736 2.048 26.244 ;
  LAYER M3 ;
        RECT 1.952 23.736 1.984 26.244 ;
  LAYER M3 ;
        RECT 1.888 23.736 1.92 26.244 ;
  LAYER M3 ;
        RECT 1.824 23.736 1.856 26.244 ;
  LAYER M3 ;
        RECT 1.76 23.736 1.792 26.244 ;
  LAYER M3 ;
        RECT 1.696 23.736 1.728 26.244 ;
  LAYER M3 ;
        RECT 1.632 23.736 1.664 26.244 ;
  LAYER M3 ;
        RECT 1.568 23.736 1.6 26.244 ;
  LAYER M3 ;
        RECT 1.504 23.736 1.536 26.244 ;
  LAYER M3 ;
        RECT 1.44 23.736 1.472 26.244 ;
  LAYER M3 ;
        RECT 1.376 23.736 1.408 26.244 ;
  LAYER M3 ;
        RECT 1.312 23.736 1.344 26.244 ;
  LAYER M3 ;
        RECT 1.248 23.736 1.28 26.244 ;
  LAYER M3 ;
        RECT 1.184 23.736 1.216 26.244 ;
  LAYER M3 ;
        RECT 1.12 23.736 1.152 26.244 ;
  LAYER M3 ;
        RECT 1.024 23.736 1.056 26.244 ;
  LAYER M1 ;
        RECT 3.439 23.772 3.441 26.208 ;
  LAYER M1 ;
        RECT 3.359 23.772 3.361 26.208 ;
  LAYER M1 ;
        RECT 3.279 23.772 3.281 26.208 ;
  LAYER M1 ;
        RECT 3.199 23.772 3.201 26.208 ;
  LAYER M1 ;
        RECT 3.119 23.772 3.121 26.208 ;
  LAYER M1 ;
        RECT 3.039 23.772 3.041 26.208 ;
  LAYER M1 ;
        RECT 2.959 23.772 2.961 26.208 ;
  LAYER M1 ;
        RECT 2.879 23.772 2.881 26.208 ;
  LAYER M1 ;
        RECT 2.799 23.772 2.801 26.208 ;
  LAYER M1 ;
        RECT 2.719 23.772 2.721 26.208 ;
  LAYER M1 ;
        RECT 2.639 23.772 2.641 26.208 ;
  LAYER M1 ;
        RECT 2.559 23.772 2.561 26.208 ;
  LAYER M1 ;
        RECT 2.479 23.772 2.481 26.208 ;
  LAYER M1 ;
        RECT 2.399 23.772 2.401 26.208 ;
  LAYER M1 ;
        RECT 2.319 23.772 2.321 26.208 ;
  LAYER M1 ;
        RECT 2.239 23.772 2.241 26.208 ;
  LAYER M1 ;
        RECT 2.159 23.772 2.161 26.208 ;
  LAYER M1 ;
        RECT 2.079 23.772 2.081 26.208 ;
  LAYER M1 ;
        RECT 1.999 23.772 2.001 26.208 ;
  LAYER M1 ;
        RECT 1.919 23.772 1.921 26.208 ;
  LAYER M1 ;
        RECT 1.839 23.772 1.841 26.208 ;
  LAYER M1 ;
        RECT 1.759 23.772 1.761 26.208 ;
  LAYER M1 ;
        RECT 1.679 23.772 1.681 26.208 ;
  LAYER M1 ;
        RECT 1.599 23.772 1.601 26.208 ;
  LAYER M1 ;
        RECT 1.519 23.772 1.521 26.208 ;
  LAYER M1 ;
        RECT 1.439 23.772 1.441 26.208 ;
  LAYER M1 ;
        RECT 1.359 23.772 1.361 26.208 ;
  LAYER M1 ;
        RECT 1.279 23.772 1.281 26.208 ;
  LAYER M1 ;
        RECT 1.199 23.772 1.201 26.208 ;
  LAYER M1 ;
        RECT 1.119 23.772 1.121 26.208 ;
  LAYER M2 ;
        RECT 1.04 23.771 3.44 23.773 ;
  LAYER M2 ;
        RECT 1.04 23.855 3.44 23.857 ;
  LAYER M2 ;
        RECT 1.04 23.939 3.44 23.941 ;
  LAYER M2 ;
        RECT 1.04 24.023 3.44 24.025 ;
  LAYER M2 ;
        RECT 1.04 24.107 3.44 24.109 ;
  LAYER M2 ;
        RECT 1.04 24.191 3.44 24.193 ;
  LAYER M2 ;
        RECT 1.04 24.275 3.44 24.277 ;
  LAYER M2 ;
        RECT 1.04 24.359 3.44 24.361 ;
  LAYER M2 ;
        RECT 1.04 24.443 3.44 24.445 ;
  LAYER M2 ;
        RECT 1.04 24.527 3.44 24.529 ;
  LAYER M2 ;
        RECT 1.04 24.611 3.44 24.613 ;
  LAYER M2 ;
        RECT 1.04 24.695 3.44 24.697 ;
  LAYER M2 ;
        RECT 1.04 24.7785 3.44 24.7805 ;
  LAYER M2 ;
        RECT 1.04 24.863 3.44 24.865 ;
  LAYER M2 ;
        RECT 1.04 24.947 3.44 24.949 ;
  LAYER M2 ;
        RECT 1.04 25.031 3.44 25.033 ;
  LAYER M2 ;
        RECT 1.04 25.115 3.44 25.117 ;
  LAYER M2 ;
        RECT 1.04 25.199 3.44 25.201 ;
  LAYER M2 ;
        RECT 1.04 25.283 3.44 25.285 ;
  LAYER M2 ;
        RECT 1.04 25.367 3.44 25.369 ;
  LAYER M2 ;
        RECT 1.04 25.451 3.44 25.453 ;
  LAYER M2 ;
        RECT 1.04 25.535 3.44 25.537 ;
  LAYER M2 ;
        RECT 1.04 25.619 3.44 25.621 ;
  LAYER M2 ;
        RECT 1.04 25.703 3.44 25.705 ;
  LAYER M2 ;
        RECT 1.04 25.787 3.44 25.789 ;
  LAYER M2 ;
        RECT 1.04 25.871 3.44 25.873 ;
  LAYER M2 ;
        RECT 1.04 25.955 3.44 25.957 ;
  LAYER M2 ;
        RECT 1.04 26.039 3.44 26.041 ;
  LAYER M2 ;
        RECT 1.04 26.123 3.44 26.125 ;
  LAYER M1 ;
        RECT 3.424 26.676 3.456 29.184 ;
  LAYER M1 ;
        RECT 3.36 26.676 3.392 29.184 ;
  LAYER M1 ;
        RECT 3.296 26.676 3.328 29.184 ;
  LAYER M1 ;
        RECT 3.232 26.676 3.264 29.184 ;
  LAYER M1 ;
        RECT 3.168 26.676 3.2 29.184 ;
  LAYER M1 ;
        RECT 3.104 26.676 3.136 29.184 ;
  LAYER M1 ;
        RECT 3.04 26.676 3.072 29.184 ;
  LAYER M1 ;
        RECT 2.976 26.676 3.008 29.184 ;
  LAYER M1 ;
        RECT 2.912 26.676 2.944 29.184 ;
  LAYER M1 ;
        RECT 2.848 26.676 2.88 29.184 ;
  LAYER M1 ;
        RECT 2.784 26.676 2.816 29.184 ;
  LAYER M1 ;
        RECT 2.72 26.676 2.752 29.184 ;
  LAYER M1 ;
        RECT 2.656 26.676 2.688 29.184 ;
  LAYER M1 ;
        RECT 2.592 26.676 2.624 29.184 ;
  LAYER M1 ;
        RECT 2.528 26.676 2.56 29.184 ;
  LAYER M1 ;
        RECT 2.464 26.676 2.496 29.184 ;
  LAYER M1 ;
        RECT 2.4 26.676 2.432 29.184 ;
  LAYER M1 ;
        RECT 2.336 26.676 2.368 29.184 ;
  LAYER M1 ;
        RECT 2.272 26.676 2.304 29.184 ;
  LAYER M1 ;
        RECT 2.208 26.676 2.24 29.184 ;
  LAYER M1 ;
        RECT 2.144 26.676 2.176 29.184 ;
  LAYER M1 ;
        RECT 2.08 26.676 2.112 29.184 ;
  LAYER M1 ;
        RECT 2.016 26.676 2.048 29.184 ;
  LAYER M1 ;
        RECT 1.952 26.676 1.984 29.184 ;
  LAYER M1 ;
        RECT 1.888 26.676 1.92 29.184 ;
  LAYER M1 ;
        RECT 1.824 26.676 1.856 29.184 ;
  LAYER M1 ;
        RECT 1.76 26.676 1.792 29.184 ;
  LAYER M1 ;
        RECT 1.696 26.676 1.728 29.184 ;
  LAYER M1 ;
        RECT 1.632 26.676 1.664 29.184 ;
  LAYER M1 ;
        RECT 1.568 26.676 1.6 29.184 ;
  LAYER M1 ;
        RECT 1.504 26.676 1.536 29.184 ;
  LAYER M1 ;
        RECT 1.44 26.676 1.472 29.184 ;
  LAYER M1 ;
        RECT 1.376 26.676 1.408 29.184 ;
  LAYER M1 ;
        RECT 1.312 26.676 1.344 29.184 ;
  LAYER M1 ;
        RECT 1.248 26.676 1.28 29.184 ;
  LAYER M1 ;
        RECT 1.184 26.676 1.216 29.184 ;
  LAYER M1 ;
        RECT 1.12 26.676 1.152 29.184 ;
  LAYER M2 ;
        RECT 1.004 26.76 3.476 26.792 ;
  LAYER M2 ;
        RECT 1.004 26.824 3.476 26.856 ;
  LAYER M2 ;
        RECT 1.004 26.888 3.476 26.92 ;
  LAYER M2 ;
        RECT 1.004 26.952 3.476 26.984 ;
  LAYER M2 ;
        RECT 1.004 27.016 3.476 27.048 ;
  LAYER M2 ;
        RECT 1.004 27.08 3.476 27.112 ;
  LAYER M2 ;
        RECT 1.004 27.144 3.476 27.176 ;
  LAYER M2 ;
        RECT 1.004 27.208 3.476 27.24 ;
  LAYER M2 ;
        RECT 1.004 27.272 3.476 27.304 ;
  LAYER M2 ;
        RECT 1.004 27.336 3.476 27.368 ;
  LAYER M2 ;
        RECT 1.004 27.4 3.476 27.432 ;
  LAYER M2 ;
        RECT 1.004 27.464 3.476 27.496 ;
  LAYER M2 ;
        RECT 1.004 27.528 3.476 27.56 ;
  LAYER M2 ;
        RECT 1.004 27.592 3.476 27.624 ;
  LAYER M2 ;
        RECT 1.004 27.656 3.476 27.688 ;
  LAYER M2 ;
        RECT 1.004 27.72 3.476 27.752 ;
  LAYER M2 ;
        RECT 1.004 27.784 3.476 27.816 ;
  LAYER M2 ;
        RECT 1.004 27.848 3.476 27.88 ;
  LAYER M2 ;
        RECT 1.004 27.912 3.476 27.944 ;
  LAYER M2 ;
        RECT 1.004 27.976 3.476 28.008 ;
  LAYER M2 ;
        RECT 1.004 28.04 3.476 28.072 ;
  LAYER M2 ;
        RECT 1.004 28.104 3.476 28.136 ;
  LAYER M2 ;
        RECT 1.004 28.168 3.476 28.2 ;
  LAYER M2 ;
        RECT 1.004 28.232 3.476 28.264 ;
  LAYER M2 ;
        RECT 1.004 28.296 3.476 28.328 ;
  LAYER M2 ;
        RECT 1.004 28.36 3.476 28.392 ;
  LAYER M2 ;
        RECT 1.004 28.424 3.476 28.456 ;
  LAYER M2 ;
        RECT 1.004 28.488 3.476 28.52 ;
  LAYER M2 ;
        RECT 1.004 28.552 3.476 28.584 ;
  LAYER M2 ;
        RECT 1.004 28.616 3.476 28.648 ;
  LAYER M2 ;
        RECT 1.004 28.68 3.476 28.712 ;
  LAYER M2 ;
        RECT 1.004 28.744 3.476 28.776 ;
  LAYER M2 ;
        RECT 1.004 28.808 3.476 28.84 ;
  LAYER M2 ;
        RECT 1.004 28.872 3.476 28.904 ;
  LAYER M2 ;
        RECT 1.004 28.936 3.476 28.968 ;
  LAYER M2 ;
        RECT 1.004 29 3.476 29.032 ;
  LAYER M3 ;
        RECT 3.424 26.676 3.456 29.184 ;
  LAYER M3 ;
        RECT 3.36 26.676 3.392 29.184 ;
  LAYER M3 ;
        RECT 3.296 26.676 3.328 29.184 ;
  LAYER M3 ;
        RECT 3.232 26.676 3.264 29.184 ;
  LAYER M3 ;
        RECT 3.168 26.676 3.2 29.184 ;
  LAYER M3 ;
        RECT 3.104 26.676 3.136 29.184 ;
  LAYER M3 ;
        RECT 3.04 26.676 3.072 29.184 ;
  LAYER M3 ;
        RECT 2.976 26.676 3.008 29.184 ;
  LAYER M3 ;
        RECT 2.912 26.676 2.944 29.184 ;
  LAYER M3 ;
        RECT 2.848 26.676 2.88 29.184 ;
  LAYER M3 ;
        RECT 2.784 26.676 2.816 29.184 ;
  LAYER M3 ;
        RECT 2.72 26.676 2.752 29.184 ;
  LAYER M3 ;
        RECT 2.656 26.676 2.688 29.184 ;
  LAYER M3 ;
        RECT 2.592 26.676 2.624 29.184 ;
  LAYER M3 ;
        RECT 2.528 26.676 2.56 29.184 ;
  LAYER M3 ;
        RECT 2.464 26.676 2.496 29.184 ;
  LAYER M3 ;
        RECT 2.4 26.676 2.432 29.184 ;
  LAYER M3 ;
        RECT 2.336 26.676 2.368 29.184 ;
  LAYER M3 ;
        RECT 2.272 26.676 2.304 29.184 ;
  LAYER M3 ;
        RECT 2.208 26.676 2.24 29.184 ;
  LAYER M3 ;
        RECT 2.144 26.676 2.176 29.184 ;
  LAYER M3 ;
        RECT 2.08 26.676 2.112 29.184 ;
  LAYER M3 ;
        RECT 2.016 26.676 2.048 29.184 ;
  LAYER M3 ;
        RECT 1.952 26.676 1.984 29.184 ;
  LAYER M3 ;
        RECT 1.888 26.676 1.92 29.184 ;
  LAYER M3 ;
        RECT 1.824 26.676 1.856 29.184 ;
  LAYER M3 ;
        RECT 1.76 26.676 1.792 29.184 ;
  LAYER M3 ;
        RECT 1.696 26.676 1.728 29.184 ;
  LAYER M3 ;
        RECT 1.632 26.676 1.664 29.184 ;
  LAYER M3 ;
        RECT 1.568 26.676 1.6 29.184 ;
  LAYER M3 ;
        RECT 1.504 26.676 1.536 29.184 ;
  LAYER M3 ;
        RECT 1.44 26.676 1.472 29.184 ;
  LAYER M3 ;
        RECT 1.376 26.676 1.408 29.184 ;
  LAYER M3 ;
        RECT 1.312 26.676 1.344 29.184 ;
  LAYER M3 ;
        RECT 1.248 26.676 1.28 29.184 ;
  LAYER M3 ;
        RECT 1.184 26.676 1.216 29.184 ;
  LAYER M3 ;
        RECT 1.12 26.676 1.152 29.184 ;
  LAYER M3 ;
        RECT 1.024 26.676 1.056 29.184 ;
  LAYER M1 ;
        RECT 3.439 26.712 3.441 29.148 ;
  LAYER M1 ;
        RECT 3.359 26.712 3.361 29.148 ;
  LAYER M1 ;
        RECT 3.279 26.712 3.281 29.148 ;
  LAYER M1 ;
        RECT 3.199 26.712 3.201 29.148 ;
  LAYER M1 ;
        RECT 3.119 26.712 3.121 29.148 ;
  LAYER M1 ;
        RECT 3.039 26.712 3.041 29.148 ;
  LAYER M1 ;
        RECT 2.959 26.712 2.961 29.148 ;
  LAYER M1 ;
        RECT 2.879 26.712 2.881 29.148 ;
  LAYER M1 ;
        RECT 2.799 26.712 2.801 29.148 ;
  LAYER M1 ;
        RECT 2.719 26.712 2.721 29.148 ;
  LAYER M1 ;
        RECT 2.639 26.712 2.641 29.148 ;
  LAYER M1 ;
        RECT 2.559 26.712 2.561 29.148 ;
  LAYER M1 ;
        RECT 2.479 26.712 2.481 29.148 ;
  LAYER M1 ;
        RECT 2.399 26.712 2.401 29.148 ;
  LAYER M1 ;
        RECT 2.319 26.712 2.321 29.148 ;
  LAYER M1 ;
        RECT 2.239 26.712 2.241 29.148 ;
  LAYER M1 ;
        RECT 2.159 26.712 2.161 29.148 ;
  LAYER M1 ;
        RECT 2.079 26.712 2.081 29.148 ;
  LAYER M1 ;
        RECT 1.999 26.712 2.001 29.148 ;
  LAYER M1 ;
        RECT 1.919 26.712 1.921 29.148 ;
  LAYER M1 ;
        RECT 1.839 26.712 1.841 29.148 ;
  LAYER M1 ;
        RECT 1.759 26.712 1.761 29.148 ;
  LAYER M1 ;
        RECT 1.679 26.712 1.681 29.148 ;
  LAYER M1 ;
        RECT 1.599 26.712 1.601 29.148 ;
  LAYER M1 ;
        RECT 1.519 26.712 1.521 29.148 ;
  LAYER M1 ;
        RECT 1.439 26.712 1.441 29.148 ;
  LAYER M1 ;
        RECT 1.359 26.712 1.361 29.148 ;
  LAYER M1 ;
        RECT 1.279 26.712 1.281 29.148 ;
  LAYER M1 ;
        RECT 1.199 26.712 1.201 29.148 ;
  LAYER M1 ;
        RECT 1.119 26.712 1.121 29.148 ;
  LAYER M2 ;
        RECT 1.04 26.711 3.44 26.713 ;
  LAYER M2 ;
        RECT 1.04 26.795 3.44 26.797 ;
  LAYER M2 ;
        RECT 1.04 26.879 3.44 26.881 ;
  LAYER M2 ;
        RECT 1.04 26.963 3.44 26.965 ;
  LAYER M2 ;
        RECT 1.04 27.047 3.44 27.049 ;
  LAYER M2 ;
        RECT 1.04 27.131 3.44 27.133 ;
  LAYER M2 ;
        RECT 1.04 27.215 3.44 27.217 ;
  LAYER M2 ;
        RECT 1.04 27.299 3.44 27.301 ;
  LAYER M2 ;
        RECT 1.04 27.383 3.44 27.385 ;
  LAYER M2 ;
        RECT 1.04 27.467 3.44 27.469 ;
  LAYER M2 ;
        RECT 1.04 27.551 3.44 27.553 ;
  LAYER M2 ;
        RECT 1.04 27.635 3.44 27.637 ;
  LAYER M2 ;
        RECT 1.04 27.7185 3.44 27.7205 ;
  LAYER M2 ;
        RECT 1.04 27.803 3.44 27.805 ;
  LAYER M2 ;
        RECT 1.04 27.887 3.44 27.889 ;
  LAYER M2 ;
        RECT 1.04 27.971 3.44 27.973 ;
  LAYER M2 ;
        RECT 1.04 28.055 3.44 28.057 ;
  LAYER M2 ;
        RECT 1.04 28.139 3.44 28.141 ;
  LAYER M2 ;
        RECT 1.04 28.223 3.44 28.225 ;
  LAYER M2 ;
        RECT 1.04 28.307 3.44 28.309 ;
  LAYER M2 ;
        RECT 1.04 28.391 3.44 28.393 ;
  LAYER M2 ;
        RECT 1.04 28.475 3.44 28.477 ;
  LAYER M2 ;
        RECT 1.04 28.559 3.44 28.561 ;
  LAYER M2 ;
        RECT 1.04 28.643 3.44 28.645 ;
  LAYER M2 ;
        RECT 1.04 28.727 3.44 28.729 ;
  LAYER M2 ;
        RECT 1.04 28.811 3.44 28.813 ;
  LAYER M2 ;
        RECT 1.04 28.895 3.44 28.897 ;
  LAYER M2 ;
        RECT 1.04 28.979 3.44 28.981 ;
  LAYER M2 ;
        RECT 1.04 29.063 3.44 29.065 ;
  LAYER M1 ;
        RECT 10.464 0.216 10.496 0.876 ;
  LAYER M1 ;
        RECT 10.544 0.216 10.576 0.876 ;
  LAYER M1 ;
        RECT 10.384 0.216 10.416 0.876 ;
  LAYER M2 ;
        RECT 10.364 0.824 10.676 0.856 ;
  LAYER M2 ;
        RECT 10.364 0.572 10.676 0.604 ;
  LAYER M2 ;
        RECT 10.284 0.74 10.596 0.772 ;
  LAYER M2 ;
        RECT 10.284 0.488 10.596 0.52 ;
  LAYER M2 ;
        RECT 10.204 0.656 10.596 0.688 ;
  LAYER M2 ;
        RECT 10.431 0.824 10.529 0.856 ;
  LAYER M1 ;
        RECT 0.384 17.268 0.416 17.928 ;
  LAYER M1 ;
        RECT 0.464 17.268 0.496 17.928 ;
  LAYER M1 ;
        RECT 0.304 17.268 0.336 17.928 ;
  LAYER M2 ;
        RECT 0.284 17.876 0.596 17.908 ;
  LAYER M2 ;
        RECT 0.284 17.624 0.596 17.656 ;
  LAYER M2 ;
        RECT 0.204 17.792 0.516 17.824 ;
  LAYER M2 ;
        RECT 0.204 17.54 0.516 17.572 ;
  LAYER M2 ;
        RECT 0.124 17.708 0.516 17.74 ;
  LAYER M2 ;
        RECT 0.351 17.876 0.449 17.908 ;
  LAYER M1 ;
        RECT 9.104 0.216 9.136 0.876 ;
  LAYER M1 ;
        RECT 9.024 0.216 9.056 0.876 ;
  LAYER M1 ;
        RECT 9.184 0.216 9.216 0.876 ;
  LAYER M1 ;
        RECT 9.744 0.216 9.776 0.876 ;
  LAYER M1 ;
        RECT 9.664 0.216 9.696 0.876 ;
  LAYER M1 ;
        RECT 9.711 0.824 9.8085 0.856 ;
  LAYER M1 ;
        RECT 8.384 0.216 8.416 0.876 ;
  LAYER M1 ;
        RECT 8.464 0.216 8.496 0.876 ;
  LAYER M1 ;
        RECT 8.304 0.216 8.336 0.876 ;
  LAYER M1 ;
        RECT 7.744 0.216 7.776 0.876 ;
  LAYER M1 ;
        RECT 7.824 0.216 7.856 0.876 ;
  LAYER M1 ;
        RECT 7.7115 0.824 7.809 0.856 ;
  LAYER M1 ;
        RECT 6.864 10.212 6.896 10.284 ;
  LAYER M2 ;
        RECT 6.844 10.232 6.916 10.264 ;
  LAYER M2 ;
        RECT 6.56 10.232 6.88 10.264 ;
  LAYER M1 ;
        RECT 6.544 10.212 6.576 10.284 ;
  LAYER M2 ;
        RECT 6.524 10.232 6.596 10.264 ;
  LAYER M1 ;
        RECT 3.984 7.272 4.016 7.344 ;
  LAYER M2 ;
        RECT 3.964 7.292 4.036 7.324 ;
  LAYER M1 ;
        RECT 3.984 7.308 4.016 7.476 ;
  LAYER M1 ;
        RECT 3.984 7.44 4.016 7.512 ;
  LAYER M2 ;
        RECT 3.964 7.46 4.036 7.492 ;
  LAYER M2 ;
        RECT 4 7.46 6.56 7.492 ;
  LAYER M1 ;
        RECT 6.544 7.44 6.576 7.512 ;
  LAYER M2 ;
        RECT 6.524 7.46 6.596 7.492 ;
  LAYER M1 ;
        RECT 6.544 16.596 6.576 16.668 ;
  LAYER M2 ;
        RECT 6.524 16.616 6.596 16.648 ;
  LAYER M1 ;
        RECT 6.544 16.464 6.576 16.632 ;
  LAYER M1 ;
        RECT 6.544 7.476 6.576 16.464 ;
  LAYER M1 ;
        RECT 9.744 13.152 9.776 13.224 ;
  LAYER M2 ;
        RECT 9.724 13.172 9.796 13.204 ;
  LAYER M2 ;
        RECT 9.44 13.172 9.76 13.204 ;
  LAYER M1 ;
        RECT 9.424 13.152 9.456 13.224 ;
  LAYER M2 ;
        RECT 9.404 13.172 9.476 13.204 ;
  LAYER M1 ;
        RECT 9.424 16.596 9.456 16.668 ;
  LAYER M2 ;
        RECT 9.404 16.616 9.476 16.648 ;
  LAYER M1 ;
        RECT 9.424 16.464 9.456 16.632 ;
  LAYER M1 ;
        RECT 9.424 13.188 9.456 16.464 ;
  LAYER M2 ;
        RECT 6.56 16.616 9.44 16.648 ;
  LAYER M1 ;
        RECT 3.984 10.212 4.016 10.284 ;
  LAYER M2 ;
        RECT 3.964 10.232 4.036 10.264 ;
  LAYER M2 ;
        RECT 3.68 10.232 4 10.264 ;
  LAYER M1 ;
        RECT 3.664 10.212 3.696 10.284 ;
  LAYER M2 ;
        RECT 3.644 10.232 3.716 10.264 ;
  LAYER M1 ;
        RECT 3.984 13.152 4.016 13.224 ;
  LAYER M2 ;
        RECT 3.964 13.172 4.036 13.204 ;
  LAYER M2 ;
        RECT 3.68 13.172 4 13.204 ;
  LAYER M1 ;
        RECT 3.664 13.152 3.696 13.224 ;
  LAYER M2 ;
        RECT 3.644 13.172 3.716 13.204 ;
  LAYER M1 ;
        RECT 3.664 16.764 3.696 16.836 ;
  LAYER M2 ;
        RECT 3.644 16.784 3.716 16.816 ;
  LAYER M1 ;
        RECT 3.664 16.464 3.696 16.8 ;
  LAYER M1 ;
        RECT 3.664 10.248 3.696 16.464 ;
  LAYER M1 ;
        RECT 9.744 10.212 9.776 10.284 ;
  LAYER M2 ;
        RECT 9.724 10.232 9.796 10.264 ;
  LAYER M1 ;
        RECT 9.744 10.248 9.776 10.416 ;
  LAYER M1 ;
        RECT 9.744 10.38 9.776 10.452 ;
  LAYER M2 ;
        RECT 9.724 10.4 9.796 10.432 ;
  LAYER M2 ;
        RECT 9.76 10.4 12.32 10.432 ;
  LAYER M1 ;
        RECT 12.304 10.38 12.336 10.452 ;
  LAYER M2 ;
        RECT 12.284 10.4 12.356 10.432 ;
  LAYER M1 ;
        RECT 9.744 7.272 9.776 7.344 ;
  LAYER M2 ;
        RECT 9.724 7.292 9.796 7.324 ;
  LAYER M1 ;
        RECT 9.744 7.308 9.776 7.476 ;
  LAYER M1 ;
        RECT 9.744 7.44 9.776 7.512 ;
  LAYER M2 ;
        RECT 9.724 7.46 9.796 7.492 ;
  LAYER M2 ;
        RECT 9.76 7.46 12.32 7.492 ;
  LAYER M1 ;
        RECT 12.304 7.44 12.336 7.512 ;
  LAYER M2 ;
        RECT 12.284 7.46 12.356 7.492 ;
  LAYER M1 ;
        RECT 12.304 16.764 12.336 16.836 ;
  LAYER M2 ;
        RECT 12.284 16.784 12.356 16.816 ;
  LAYER M1 ;
        RECT 12.304 16.464 12.336 16.8 ;
  LAYER M1 ;
        RECT 12.304 7.476 12.336 16.464 ;
  LAYER M2 ;
        RECT 3.68 16.784 12.32 16.816 ;
  LAYER M1 ;
        RECT 6.864 13.152 6.896 13.224 ;
  LAYER M2 ;
        RECT 6.844 13.172 6.916 13.204 ;
  LAYER M2 ;
        RECT 4 13.172 6.88 13.204 ;
  LAYER M1 ;
        RECT 3.984 13.152 4.016 13.224 ;
  LAYER M2 ;
        RECT 3.964 13.172 4.036 13.204 ;
  LAYER M1 ;
        RECT 6.864 7.272 6.896 7.344 ;
  LAYER M2 ;
        RECT 6.844 7.292 6.916 7.324 ;
  LAYER M2 ;
        RECT 6.88 7.292 9.76 7.324 ;
  LAYER M1 ;
        RECT 9.744 7.272 9.776 7.344 ;
  LAYER M2 ;
        RECT 9.724 7.292 9.796 7.324 ;
  LAYER M1 ;
        RECT 1.104 16.092 1.136 16.164 ;
  LAYER M2 ;
        RECT 1.084 16.112 1.156 16.144 ;
  LAYER M2 ;
        RECT 0.8 16.112 1.12 16.144 ;
  LAYER M1 ;
        RECT 0.784 16.092 0.816 16.164 ;
  LAYER M2 ;
        RECT 0.764 16.112 0.836 16.144 ;
  LAYER M1 ;
        RECT 1.104 13.152 1.136 13.224 ;
  LAYER M2 ;
        RECT 1.084 13.172 1.156 13.204 ;
  LAYER M2 ;
        RECT 0.8 13.172 1.12 13.204 ;
  LAYER M1 ;
        RECT 0.784 13.152 0.816 13.224 ;
  LAYER M2 ;
        RECT 0.764 13.172 0.836 13.204 ;
  LAYER M1 ;
        RECT 1.104 10.212 1.136 10.284 ;
  LAYER M2 ;
        RECT 1.084 10.232 1.156 10.264 ;
  LAYER M2 ;
        RECT 0.8 10.232 1.12 10.264 ;
  LAYER M1 ;
        RECT 0.784 10.212 0.816 10.284 ;
  LAYER M2 ;
        RECT 0.764 10.232 0.836 10.264 ;
  LAYER M1 ;
        RECT 1.104 7.272 1.136 7.344 ;
  LAYER M2 ;
        RECT 1.084 7.292 1.156 7.324 ;
  LAYER M2 ;
        RECT 0.8 7.292 1.12 7.324 ;
  LAYER M1 ;
        RECT 0.784 7.272 0.816 7.344 ;
  LAYER M2 ;
        RECT 0.764 7.292 0.836 7.324 ;
  LAYER M1 ;
        RECT 1.104 4.332 1.136 4.404 ;
  LAYER M2 ;
        RECT 1.084 4.352 1.156 4.384 ;
  LAYER M2 ;
        RECT 0.8 4.352 1.12 4.384 ;
  LAYER M1 ;
        RECT 0.784 4.332 0.816 4.404 ;
  LAYER M2 ;
        RECT 0.764 4.352 0.836 4.384 ;
  LAYER M1 ;
        RECT 0.784 16.932 0.816 17.004 ;
  LAYER M2 ;
        RECT 0.764 16.952 0.836 16.984 ;
  LAYER M1 ;
        RECT 0.784 16.464 0.816 16.968 ;
  LAYER M1 ;
        RECT 0.784 4.368 0.816 16.464 ;
  LAYER M1 ;
        RECT 12.624 16.092 12.656 16.164 ;
  LAYER M2 ;
        RECT 12.604 16.112 12.676 16.144 ;
  LAYER M1 ;
        RECT 12.624 16.128 12.656 16.296 ;
  LAYER M1 ;
        RECT 12.624 16.26 12.656 16.332 ;
  LAYER M2 ;
        RECT 12.604 16.28 12.676 16.312 ;
  LAYER M2 ;
        RECT 12.64 16.28 15.2 16.312 ;
  LAYER M1 ;
        RECT 15.184 16.26 15.216 16.332 ;
  LAYER M2 ;
        RECT 15.164 16.28 15.236 16.312 ;
  LAYER M1 ;
        RECT 12.624 13.152 12.656 13.224 ;
  LAYER M2 ;
        RECT 12.604 13.172 12.676 13.204 ;
  LAYER M1 ;
        RECT 12.624 13.188 12.656 13.356 ;
  LAYER M1 ;
        RECT 12.624 13.32 12.656 13.392 ;
  LAYER M2 ;
        RECT 12.604 13.34 12.676 13.372 ;
  LAYER M2 ;
        RECT 12.64 13.34 15.2 13.372 ;
  LAYER M1 ;
        RECT 15.184 13.32 15.216 13.392 ;
  LAYER M2 ;
        RECT 15.164 13.34 15.236 13.372 ;
  LAYER M1 ;
        RECT 12.624 10.212 12.656 10.284 ;
  LAYER M2 ;
        RECT 12.604 10.232 12.676 10.264 ;
  LAYER M1 ;
        RECT 12.624 10.248 12.656 10.416 ;
  LAYER M1 ;
        RECT 12.624 10.38 12.656 10.452 ;
  LAYER M2 ;
        RECT 12.604 10.4 12.676 10.432 ;
  LAYER M2 ;
        RECT 12.64 10.4 15.2 10.432 ;
  LAYER M1 ;
        RECT 15.184 10.38 15.216 10.452 ;
  LAYER M2 ;
        RECT 15.164 10.4 15.236 10.432 ;
  LAYER M1 ;
        RECT 12.624 7.272 12.656 7.344 ;
  LAYER M2 ;
        RECT 12.604 7.292 12.676 7.324 ;
  LAYER M1 ;
        RECT 12.624 7.308 12.656 7.476 ;
  LAYER M1 ;
        RECT 12.624 7.44 12.656 7.512 ;
  LAYER M2 ;
        RECT 12.604 7.46 12.676 7.492 ;
  LAYER M2 ;
        RECT 12.64 7.46 15.2 7.492 ;
  LAYER M1 ;
        RECT 15.184 7.44 15.216 7.512 ;
  LAYER M2 ;
        RECT 15.164 7.46 15.236 7.492 ;
  LAYER M1 ;
        RECT 12.624 4.332 12.656 4.404 ;
  LAYER M2 ;
        RECT 12.604 4.352 12.676 4.384 ;
  LAYER M1 ;
        RECT 12.624 4.368 12.656 4.536 ;
  LAYER M1 ;
        RECT 12.624 4.5 12.656 4.572 ;
  LAYER M2 ;
        RECT 12.604 4.52 12.676 4.552 ;
  LAYER M2 ;
        RECT 12.64 4.52 15.2 4.552 ;
  LAYER M1 ;
        RECT 15.184 4.5 15.216 4.572 ;
  LAYER M2 ;
        RECT 15.164 4.52 15.236 4.552 ;
  LAYER M1 ;
        RECT 15.184 16.932 15.216 17.004 ;
  LAYER M2 ;
        RECT 15.164 16.952 15.236 16.984 ;
  LAYER M1 ;
        RECT 15.184 16.464 15.216 16.968 ;
  LAYER M1 ;
        RECT 15.184 4.536 15.216 16.464 ;
  LAYER M2 ;
        RECT 0.8 16.952 15.2 16.984 ;
  LAYER M1 ;
        RECT 3.984 16.092 4.016 16.164 ;
  LAYER M2 ;
        RECT 3.964 16.112 4.036 16.144 ;
  LAYER M2 ;
        RECT 1.12 16.112 4 16.144 ;
  LAYER M1 ;
        RECT 1.104 16.092 1.136 16.164 ;
  LAYER M2 ;
        RECT 1.084 16.112 1.156 16.144 ;
  LAYER M1 ;
        RECT 3.984 4.332 4.016 4.404 ;
  LAYER M2 ;
        RECT 3.964 4.352 4.036 4.384 ;
  LAYER M2 ;
        RECT 1.12 4.352 4 4.384 ;
  LAYER M1 ;
        RECT 1.104 4.332 1.136 4.404 ;
  LAYER M2 ;
        RECT 1.084 4.352 1.156 4.384 ;
  LAYER M1 ;
        RECT 6.864 4.332 6.896 4.404 ;
  LAYER M2 ;
        RECT 6.844 4.352 6.916 4.384 ;
  LAYER M2 ;
        RECT 4 4.352 6.88 4.384 ;
  LAYER M1 ;
        RECT 3.984 4.332 4.016 4.404 ;
  LAYER M2 ;
        RECT 3.964 4.352 4.036 4.384 ;
  LAYER M1 ;
        RECT 9.744 4.332 9.776 4.404 ;
  LAYER M2 ;
        RECT 9.724 4.352 9.796 4.384 ;
  LAYER M2 ;
        RECT 6.88 4.352 9.76 4.384 ;
  LAYER M1 ;
        RECT 6.864 4.332 6.896 4.404 ;
  LAYER M2 ;
        RECT 6.844 4.352 6.916 4.384 ;
  LAYER M1 ;
        RECT 9.744 16.092 9.776 16.164 ;
  LAYER M2 ;
        RECT 9.724 16.112 9.796 16.144 ;
  LAYER M2 ;
        RECT 9.76 16.112 12.64 16.144 ;
  LAYER M1 ;
        RECT 12.624 16.092 12.656 16.164 ;
  LAYER M2 ;
        RECT 12.604 16.112 12.676 16.144 ;
  LAYER M1 ;
        RECT 6.864 16.092 6.896 16.164 ;
  LAYER M2 ;
        RECT 6.844 16.112 6.916 16.144 ;
  LAYER M2 ;
        RECT 6.88 16.112 9.76 16.144 ;
  LAYER M1 ;
        RECT 9.744 16.092 9.776 16.164 ;
  LAYER M2 ;
        RECT 9.724 16.112 9.796 16.144 ;
  LAYER M1 ;
        RECT 9.264 7.776 9.296 7.848 ;
  LAYER M2 ;
        RECT 9.244 7.796 9.316 7.828 ;
  LAYER M2 ;
        RECT 6.72 7.796 9.28 7.828 ;
  LAYER M1 ;
        RECT 6.704 7.776 6.736 7.848 ;
  LAYER M2 ;
        RECT 6.684 7.796 6.756 7.828 ;
  LAYER M1 ;
        RECT 6.384 4.836 6.416 4.908 ;
  LAYER M2 ;
        RECT 6.364 4.856 6.436 4.888 ;
  LAYER M1 ;
        RECT 6.384 4.704 6.416 4.872 ;
  LAYER M1 ;
        RECT 6.384 4.668 6.416 4.74 ;
  LAYER M2 ;
        RECT 6.364 4.688 6.436 4.72 ;
  LAYER M2 ;
        RECT 6.4 4.688 6.72 4.72 ;
  LAYER M1 ;
        RECT 6.704 4.668 6.736 4.74 ;
  LAYER M2 ;
        RECT 6.684 4.688 6.756 4.72 ;
  LAYER M1 ;
        RECT 6.704 1.392 6.736 1.464 ;
  LAYER M2 ;
        RECT 6.684 1.412 6.756 1.444 ;
  LAYER M1 ;
        RECT 6.704 1.428 6.736 1.596 ;
  LAYER M1 ;
        RECT 6.704 1.596 6.736 7.812 ;
  LAYER M1 ;
        RECT 12.144 10.716 12.176 10.788 ;
  LAYER M2 ;
        RECT 12.124 10.736 12.196 10.768 ;
  LAYER M2 ;
        RECT 9.6 10.736 12.16 10.768 ;
  LAYER M1 ;
        RECT 9.584 10.716 9.616 10.788 ;
  LAYER M2 ;
        RECT 9.564 10.736 9.636 10.768 ;
  LAYER M1 ;
        RECT 9.584 1.392 9.616 1.464 ;
  LAYER M2 ;
        RECT 9.564 1.412 9.636 1.444 ;
  LAYER M1 ;
        RECT 9.584 1.428 9.616 1.596 ;
  LAYER M1 ;
        RECT 9.584 1.596 9.616 10.752 ;
  LAYER M2 ;
        RECT 6.72 1.412 9.6 1.444 ;
  LAYER M1 ;
        RECT 6.384 7.776 6.416 7.848 ;
  LAYER M2 ;
        RECT 6.364 7.796 6.436 7.828 ;
  LAYER M2 ;
        RECT 3.84 7.796 6.4 7.828 ;
  LAYER M1 ;
        RECT 3.824 7.776 3.856 7.848 ;
  LAYER M2 ;
        RECT 3.804 7.796 3.876 7.828 ;
  LAYER M1 ;
        RECT 6.384 10.716 6.416 10.788 ;
  LAYER M2 ;
        RECT 6.364 10.736 6.436 10.768 ;
  LAYER M2 ;
        RECT 3.84 10.736 6.4 10.768 ;
  LAYER M1 ;
        RECT 3.824 10.716 3.856 10.788 ;
  LAYER M2 ;
        RECT 3.804 10.736 3.876 10.768 ;
  LAYER M1 ;
        RECT 3.824 1.224 3.856 1.296 ;
  LAYER M2 ;
        RECT 3.804 1.244 3.876 1.276 ;
  LAYER M1 ;
        RECT 3.824 1.26 3.856 1.596 ;
  LAYER M1 ;
        RECT 3.824 1.596 3.856 10.752 ;
  LAYER M1 ;
        RECT 12.144 7.776 12.176 7.848 ;
  LAYER M2 ;
        RECT 12.124 7.796 12.196 7.828 ;
  LAYER M1 ;
        RECT 12.144 7.644 12.176 7.812 ;
  LAYER M1 ;
        RECT 12.144 7.608 12.176 7.68 ;
  LAYER M2 ;
        RECT 12.124 7.628 12.196 7.66 ;
  LAYER M2 ;
        RECT 12.16 7.628 12.48 7.66 ;
  LAYER M1 ;
        RECT 12.464 7.608 12.496 7.68 ;
  LAYER M2 ;
        RECT 12.444 7.628 12.516 7.66 ;
  LAYER M1 ;
        RECT 12.144 4.836 12.176 4.908 ;
  LAYER M2 ;
        RECT 12.124 4.856 12.196 4.888 ;
  LAYER M1 ;
        RECT 12.144 4.704 12.176 4.872 ;
  LAYER M1 ;
        RECT 12.144 4.668 12.176 4.74 ;
  LAYER M2 ;
        RECT 12.124 4.688 12.196 4.72 ;
  LAYER M2 ;
        RECT 12.16 4.688 12.48 4.72 ;
  LAYER M1 ;
        RECT 12.464 4.668 12.496 4.74 ;
  LAYER M2 ;
        RECT 12.444 4.688 12.516 4.72 ;
  LAYER M1 ;
        RECT 12.464 1.224 12.496 1.296 ;
  LAYER M2 ;
        RECT 12.444 1.244 12.516 1.276 ;
  LAYER M1 ;
        RECT 12.464 1.26 12.496 1.596 ;
  LAYER M1 ;
        RECT 12.464 1.596 12.496 7.644 ;
  LAYER M2 ;
        RECT 3.84 1.244 12.48 1.276 ;
  LAYER M1 ;
        RECT 9.264 10.716 9.296 10.788 ;
  LAYER M2 ;
        RECT 9.244 10.736 9.316 10.768 ;
  LAYER M2 ;
        RECT 6.4 10.736 9.28 10.768 ;
  LAYER M1 ;
        RECT 6.384 10.716 6.416 10.788 ;
  LAYER M2 ;
        RECT 6.364 10.736 6.436 10.768 ;
  LAYER M1 ;
        RECT 9.264 4.836 9.296 4.908 ;
  LAYER M2 ;
        RECT 9.244 4.856 9.316 4.888 ;
  LAYER M2 ;
        RECT 9.28 4.856 12.16 4.888 ;
  LAYER M1 ;
        RECT 12.144 4.836 12.176 4.908 ;
  LAYER M2 ;
        RECT 12.124 4.856 12.196 4.888 ;
  LAYER M1 ;
        RECT 3.504 13.656 3.536 13.728 ;
  LAYER M2 ;
        RECT 3.484 13.676 3.556 13.708 ;
  LAYER M2 ;
        RECT 0.96 13.676 3.52 13.708 ;
  LAYER M1 ;
        RECT 0.944 13.656 0.976 13.728 ;
  LAYER M2 ;
        RECT 0.924 13.676 0.996 13.708 ;
  LAYER M1 ;
        RECT 3.504 10.716 3.536 10.788 ;
  LAYER M2 ;
        RECT 3.484 10.736 3.556 10.768 ;
  LAYER M2 ;
        RECT 0.96 10.736 3.52 10.768 ;
  LAYER M1 ;
        RECT 0.944 10.716 0.976 10.788 ;
  LAYER M2 ;
        RECT 0.924 10.736 0.996 10.768 ;
  LAYER M1 ;
        RECT 3.504 7.776 3.536 7.848 ;
  LAYER M2 ;
        RECT 3.484 7.796 3.556 7.828 ;
  LAYER M2 ;
        RECT 0.96 7.796 3.52 7.828 ;
  LAYER M1 ;
        RECT 0.944 7.776 0.976 7.848 ;
  LAYER M2 ;
        RECT 0.924 7.796 0.996 7.828 ;
  LAYER M1 ;
        RECT 3.504 4.836 3.536 4.908 ;
  LAYER M2 ;
        RECT 3.484 4.856 3.556 4.888 ;
  LAYER M2 ;
        RECT 0.96 4.856 3.52 4.888 ;
  LAYER M1 ;
        RECT 0.944 4.836 0.976 4.908 ;
  LAYER M2 ;
        RECT 0.924 4.856 0.996 4.888 ;
  LAYER M1 ;
        RECT 3.504 1.896 3.536 1.968 ;
  LAYER M2 ;
        RECT 3.484 1.916 3.556 1.948 ;
  LAYER M2 ;
        RECT 0.96 1.916 3.52 1.948 ;
  LAYER M1 ;
        RECT 0.944 1.896 0.976 1.968 ;
  LAYER M2 ;
        RECT 0.924 1.916 0.996 1.948 ;
  LAYER M1 ;
        RECT 0.944 1.056 0.976 1.128 ;
  LAYER M2 ;
        RECT 0.924 1.076 0.996 1.108 ;
  LAYER M1 ;
        RECT 0.944 1.092 0.976 1.596 ;
  LAYER M1 ;
        RECT 0.944 1.596 0.976 13.692 ;
  LAYER M1 ;
        RECT 15.024 13.656 15.056 13.728 ;
  LAYER M2 ;
        RECT 15.004 13.676 15.076 13.708 ;
  LAYER M1 ;
        RECT 15.024 13.524 15.056 13.692 ;
  LAYER M1 ;
        RECT 15.024 13.488 15.056 13.56 ;
  LAYER M2 ;
        RECT 15.004 13.508 15.076 13.54 ;
  LAYER M2 ;
        RECT 15.04 13.508 15.36 13.54 ;
  LAYER M1 ;
        RECT 15.344 13.488 15.376 13.56 ;
  LAYER M2 ;
        RECT 15.324 13.508 15.396 13.54 ;
  LAYER M1 ;
        RECT 15.024 10.716 15.056 10.788 ;
  LAYER M2 ;
        RECT 15.004 10.736 15.076 10.768 ;
  LAYER M1 ;
        RECT 15.024 10.584 15.056 10.752 ;
  LAYER M1 ;
        RECT 15.024 10.548 15.056 10.62 ;
  LAYER M2 ;
        RECT 15.004 10.568 15.076 10.6 ;
  LAYER M2 ;
        RECT 15.04 10.568 15.36 10.6 ;
  LAYER M1 ;
        RECT 15.344 10.548 15.376 10.62 ;
  LAYER M2 ;
        RECT 15.324 10.568 15.396 10.6 ;
  LAYER M1 ;
        RECT 15.024 7.776 15.056 7.848 ;
  LAYER M2 ;
        RECT 15.004 7.796 15.076 7.828 ;
  LAYER M1 ;
        RECT 15.024 7.644 15.056 7.812 ;
  LAYER M1 ;
        RECT 15.024 7.608 15.056 7.68 ;
  LAYER M2 ;
        RECT 15.004 7.628 15.076 7.66 ;
  LAYER M2 ;
        RECT 15.04 7.628 15.36 7.66 ;
  LAYER M1 ;
        RECT 15.344 7.608 15.376 7.68 ;
  LAYER M2 ;
        RECT 15.324 7.628 15.396 7.66 ;
  LAYER M1 ;
        RECT 15.024 4.836 15.056 4.908 ;
  LAYER M2 ;
        RECT 15.004 4.856 15.076 4.888 ;
  LAYER M1 ;
        RECT 15.024 4.704 15.056 4.872 ;
  LAYER M1 ;
        RECT 15.024 4.668 15.056 4.74 ;
  LAYER M2 ;
        RECT 15.004 4.688 15.076 4.72 ;
  LAYER M2 ;
        RECT 15.04 4.688 15.36 4.72 ;
  LAYER M1 ;
        RECT 15.344 4.668 15.376 4.74 ;
  LAYER M2 ;
        RECT 15.324 4.688 15.396 4.72 ;
  LAYER M1 ;
        RECT 15.024 1.896 15.056 1.968 ;
  LAYER M2 ;
        RECT 15.004 1.916 15.076 1.948 ;
  LAYER M1 ;
        RECT 15.024 1.764 15.056 1.932 ;
  LAYER M1 ;
        RECT 15.024 1.728 15.056 1.8 ;
  LAYER M2 ;
        RECT 15.004 1.748 15.076 1.78 ;
  LAYER M2 ;
        RECT 15.04 1.748 15.36 1.78 ;
  LAYER M1 ;
        RECT 15.344 1.728 15.376 1.8 ;
  LAYER M2 ;
        RECT 15.324 1.748 15.396 1.78 ;
  LAYER M1 ;
        RECT 15.344 1.056 15.376 1.128 ;
  LAYER M2 ;
        RECT 15.324 1.076 15.396 1.108 ;
  LAYER M1 ;
        RECT 15.344 1.092 15.376 1.596 ;
  LAYER M1 ;
        RECT 15.344 1.596 15.376 13.524 ;
  LAYER M2 ;
        RECT 0.96 1.076 15.36 1.108 ;
  LAYER M1 ;
        RECT 6.384 13.656 6.416 13.728 ;
  LAYER M2 ;
        RECT 6.364 13.676 6.436 13.708 ;
  LAYER M2 ;
        RECT 3.52 13.676 6.4 13.708 ;
  LAYER M1 ;
        RECT 3.504 13.656 3.536 13.728 ;
  LAYER M2 ;
        RECT 3.484 13.676 3.556 13.708 ;
  LAYER M1 ;
        RECT 6.384 1.896 6.416 1.968 ;
  LAYER M2 ;
        RECT 6.364 1.916 6.436 1.948 ;
  LAYER M2 ;
        RECT 3.52 1.916 6.4 1.948 ;
  LAYER M1 ;
        RECT 3.504 1.896 3.536 1.968 ;
  LAYER M2 ;
        RECT 3.484 1.916 3.556 1.948 ;
  LAYER M1 ;
        RECT 9.264 1.896 9.296 1.968 ;
  LAYER M2 ;
        RECT 9.244 1.916 9.316 1.948 ;
  LAYER M2 ;
        RECT 6.4 1.916 9.28 1.948 ;
  LAYER M1 ;
        RECT 6.384 1.896 6.416 1.968 ;
  LAYER M2 ;
        RECT 6.364 1.916 6.436 1.948 ;
  LAYER M1 ;
        RECT 12.144 1.896 12.176 1.968 ;
  LAYER M2 ;
        RECT 12.124 1.916 12.196 1.948 ;
  LAYER M2 ;
        RECT 9.28 1.916 12.16 1.948 ;
  LAYER M1 ;
        RECT 9.264 1.896 9.296 1.968 ;
  LAYER M2 ;
        RECT 9.244 1.916 9.316 1.948 ;
  LAYER M1 ;
        RECT 12.144 13.656 12.176 13.728 ;
  LAYER M2 ;
        RECT 12.124 13.676 12.196 13.708 ;
  LAYER M2 ;
        RECT 12.16 13.676 15.04 13.708 ;
  LAYER M1 ;
        RECT 15.024 13.656 15.056 13.728 ;
  LAYER M2 ;
        RECT 15.004 13.676 15.076 13.708 ;
  LAYER M1 ;
        RECT 9.264 13.656 9.296 13.728 ;
  LAYER M2 ;
        RECT 9.244 13.676 9.316 13.708 ;
  LAYER M2 ;
        RECT 9.28 13.676 12.16 13.708 ;
  LAYER M1 ;
        RECT 12.144 13.656 12.176 13.728 ;
  LAYER M2 ;
        RECT 12.124 13.676 12.196 13.708 ;
  LAYER M1 ;
        RECT 1.104 13.656 1.136 16.164 ;
  LAYER M1 ;
        RECT 1.168 13.656 1.2 16.164 ;
  LAYER M1 ;
        RECT 1.232 13.656 1.264 16.164 ;
  LAYER M1 ;
        RECT 1.296 13.656 1.328 16.164 ;
  LAYER M1 ;
        RECT 1.36 13.656 1.392 16.164 ;
  LAYER M1 ;
        RECT 1.424 13.656 1.456 16.164 ;
  LAYER M1 ;
        RECT 1.488 13.656 1.52 16.164 ;
  LAYER M1 ;
        RECT 1.552 13.656 1.584 16.164 ;
  LAYER M1 ;
        RECT 1.616 13.656 1.648 16.164 ;
  LAYER M1 ;
        RECT 1.68 13.656 1.712 16.164 ;
  LAYER M1 ;
        RECT 1.744 13.656 1.776 16.164 ;
  LAYER M1 ;
        RECT 1.808 13.656 1.84 16.164 ;
  LAYER M1 ;
        RECT 1.872 13.656 1.904 16.164 ;
  LAYER M1 ;
        RECT 1.936 13.656 1.968 16.164 ;
  LAYER M1 ;
        RECT 2 13.656 2.032 16.164 ;
  LAYER M1 ;
        RECT 2.064 13.656 2.096 16.164 ;
  LAYER M1 ;
        RECT 2.128 13.656 2.16 16.164 ;
  LAYER M1 ;
        RECT 2.192 13.656 2.224 16.164 ;
  LAYER M1 ;
        RECT 2.256 13.656 2.288 16.164 ;
  LAYER M1 ;
        RECT 2.32 13.656 2.352 16.164 ;
  LAYER M1 ;
        RECT 2.384 13.656 2.416 16.164 ;
  LAYER M1 ;
        RECT 2.448 13.656 2.48 16.164 ;
  LAYER M1 ;
        RECT 2.512 13.656 2.544 16.164 ;
  LAYER M1 ;
        RECT 2.576 13.656 2.608 16.164 ;
  LAYER M1 ;
        RECT 2.64 13.656 2.672 16.164 ;
  LAYER M1 ;
        RECT 2.704 13.656 2.736 16.164 ;
  LAYER M1 ;
        RECT 2.768 13.656 2.8 16.164 ;
  LAYER M1 ;
        RECT 2.832 13.656 2.864 16.164 ;
  LAYER M1 ;
        RECT 2.896 13.656 2.928 16.164 ;
  LAYER M1 ;
        RECT 2.96 13.656 2.992 16.164 ;
  LAYER M1 ;
        RECT 3.024 13.656 3.056 16.164 ;
  LAYER M1 ;
        RECT 3.088 13.656 3.12 16.164 ;
  LAYER M1 ;
        RECT 3.152 13.656 3.184 16.164 ;
  LAYER M1 ;
        RECT 3.216 13.656 3.248 16.164 ;
  LAYER M1 ;
        RECT 3.28 13.656 3.312 16.164 ;
  LAYER M1 ;
        RECT 3.344 13.656 3.376 16.164 ;
  LAYER M1 ;
        RECT 3.408 13.656 3.44 16.164 ;
  LAYER M2 ;
        RECT 1.084 16.048 3.556 16.08 ;
  LAYER M2 ;
        RECT 1.084 15.984 3.556 16.016 ;
  LAYER M2 ;
        RECT 1.084 15.92 3.556 15.952 ;
  LAYER M2 ;
        RECT 1.084 15.856 3.556 15.888 ;
  LAYER M2 ;
        RECT 1.084 15.792 3.556 15.824 ;
  LAYER M2 ;
        RECT 1.084 15.728 3.556 15.76 ;
  LAYER M2 ;
        RECT 1.084 15.664 3.556 15.696 ;
  LAYER M2 ;
        RECT 1.084 15.6 3.556 15.632 ;
  LAYER M2 ;
        RECT 1.084 15.536 3.556 15.568 ;
  LAYER M2 ;
        RECT 1.084 15.472 3.556 15.504 ;
  LAYER M2 ;
        RECT 1.084 15.408 3.556 15.44 ;
  LAYER M2 ;
        RECT 1.084 15.344 3.556 15.376 ;
  LAYER M2 ;
        RECT 1.084 15.28 3.556 15.312 ;
  LAYER M2 ;
        RECT 1.084 15.216 3.556 15.248 ;
  LAYER M2 ;
        RECT 1.084 15.152 3.556 15.184 ;
  LAYER M2 ;
        RECT 1.084 15.088 3.556 15.12 ;
  LAYER M2 ;
        RECT 1.084 15.024 3.556 15.056 ;
  LAYER M2 ;
        RECT 1.084 14.96 3.556 14.992 ;
  LAYER M2 ;
        RECT 1.084 14.896 3.556 14.928 ;
  LAYER M2 ;
        RECT 1.084 14.832 3.556 14.864 ;
  LAYER M2 ;
        RECT 1.084 14.768 3.556 14.8 ;
  LAYER M2 ;
        RECT 1.084 14.704 3.556 14.736 ;
  LAYER M2 ;
        RECT 1.084 14.64 3.556 14.672 ;
  LAYER M2 ;
        RECT 1.084 14.576 3.556 14.608 ;
  LAYER M2 ;
        RECT 1.084 14.512 3.556 14.544 ;
  LAYER M2 ;
        RECT 1.084 14.448 3.556 14.48 ;
  LAYER M2 ;
        RECT 1.084 14.384 3.556 14.416 ;
  LAYER M2 ;
        RECT 1.084 14.32 3.556 14.352 ;
  LAYER M2 ;
        RECT 1.084 14.256 3.556 14.288 ;
  LAYER M2 ;
        RECT 1.084 14.192 3.556 14.224 ;
  LAYER M2 ;
        RECT 1.084 14.128 3.556 14.16 ;
  LAYER M2 ;
        RECT 1.084 14.064 3.556 14.096 ;
  LAYER M2 ;
        RECT 1.084 14 3.556 14.032 ;
  LAYER M2 ;
        RECT 1.084 13.936 3.556 13.968 ;
  LAYER M2 ;
        RECT 1.084 13.872 3.556 13.904 ;
  LAYER M2 ;
        RECT 1.084 13.808 3.556 13.84 ;
  LAYER M3 ;
        RECT 1.104 13.656 1.136 16.164 ;
  LAYER M3 ;
        RECT 1.168 13.656 1.2 16.164 ;
  LAYER M3 ;
        RECT 1.232 13.656 1.264 16.164 ;
  LAYER M3 ;
        RECT 1.296 13.656 1.328 16.164 ;
  LAYER M3 ;
        RECT 1.36 13.656 1.392 16.164 ;
  LAYER M3 ;
        RECT 1.424 13.656 1.456 16.164 ;
  LAYER M3 ;
        RECT 1.488 13.656 1.52 16.164 ;
  LAYER M3 ;
        RECT 1.552 13.656 1.584 16.164 ;
  LAYER M3 ;
        RECT 1.616 13.656 1.648 16.164 ;
  LAYER M3 ;
        RECT 1.68 13.656 1.712 16.164 ;
  LAYER M3 ;
        RECT 1.744 13.656 1.776 16.164 ;
  LAYER M3 ;
        RECT 1.808 13.656 1.84 16.164 ;
  LAYER M3 ;
        RECT 1.872 13.656 1.904 16.164 ;
  LAYER M3 ;
        RECT 1.936 13.656 1.968 16.164 ;
  LAYER M3 ;
        RECT 2 13.656 2.032 16.164 ;
  LAYER M3 ;
        RECT 2.064 13.656 2.096 16.164 ;
  LAYER M3 ;
        RECT 2.128 13.656 2.16 16.164 ;
  LAYER M3 ;
        RECT 2.192 13.656 2.224 16.164 ;
  LAYER M3 ;
        RECT 2.256 13.656 2.288 16.164 ;
  LAYER M3 ;
        RECT 2.32 13.656 2.352 16.164 ;
  LAYER M3 ;
        RECT 2.384 13.656 2.416 16.164 ;
  LAYER M3 ;
        RECT 2.448 13.656 2.48 16.164 ;
  LAYER M3 ;
        RECT 2.512 13.656 2.544 16.164 ;
  LAYER M3 ;
        RECT 2.576 13.656 2.608 16.164 ;
  LAYER M3 ;
        RECT 2.64 13.656 2.672 16.164 ;
  LAYER M3 ;
        RECT 2.704 13.656 2.736 16.164 ;
  LAYER M3 ;
        RECT 2.768 13.656 2.8 16.164 ;
  LAYER M3 ;
        RECT 2.832 13.656 2.864 16.164 ;
  LAYER M3 ;
        RECT 2.896 13.656 2.928 16.164 ;
  LAYER M3 ;
        RECT 2.96 13.656 2.992 16.164 ;
  LAYER M3 ;
        RECT 3.024 13.656 3.056 16.164 ;
  LAYER M3 ;
        RECT 3.088 13.656 3.12 16.164 ;
  LAYER M3 ;
        RECT 3.152 13.656 3.184 16.164 ;
  LAYER M3 ;
        RECT 3.216 13.656 3.248 16.164 ;
  LAYER M3 ;
        RECT 3.28 13.656 3.312 16.164 ;
  LAYER M3 ;
        RECT 3.344 13.656 3.376 16.164 ;
  LAYER M3 ;
        RECT 3.408 13.656 3.44 16.164 ;
  LAYER M3 ;
        RECT 3.504 13.656 3.536 16.164 ;
  LAYER M1 ;
        RECT 1.119 13.692 1.121 16.128 ;
  LAYER M1 ;
        RECT 1.199 13.692 1.201 16.128 ;
  LAYER M1 ;
        RECT 1.279 13.692 1.281 16.128 ;
  LAYER M1 ;
        RECT 1.359 13.692 1.361 16.128 ;
  LAYER M1 ;
        RECT 1.439 13.692 1.441 16.128 ;
  LAYER M1 ;
        RECT 1.519 13.692 1.521 16.128 ;
  LAYER M1 ;
        RECT 1.599 13.692 1.601 16.128 ;
  LAYER M1 ;
        RECT 1.679 13.692 1.681 16.128 ;
  LAYER M1 ;
        RECT 1.759 13.692 1.761 16.128 ;
  LAYER M1 ;
        RECT 1.839 13.692 1.841 16.128 ;
  LAYER M1 ;
        RECT 1.919 13.692 1.921 16.128 ;
  LAYER M1 ;
        RECT 1.999 13.692 2.001 16.128 ;
  LAYER M1 ;
        RECT 2.079 13.692 2.081 16.128 ;
  LAYER M1 ;
        RECT 2.159 13.692 2.161 16.128 ;
  LAYER M1 ;
        RECT 2.239 13.692 2.241 16.128 ;
  LAYER M1 ;
        RECT 2.319 13.692 2.321 16.128 ;
  LAYER M1 ;
        RECT 2.399 13.692 2.401 16.128 ;
  LAYER M1 ;
        RECT 2.479 13.692 2.481 16.128 ;
  LAYER M1 ;
        RECT 2.559 13.692 2.561 16.128 ;
  LAYER M1 ;
        RECT 2.639 13.692 2.641 16.128 ;
  LAYER M1 ;
        RECT 2.719 13.692 2.721 16.128 ;
  LAYER M1 ;
        RECT 2.799 13.692 2.801 16.128 ;
  LAYER M1 ;
        RECT 2.879 13.692 2.881 16.128 ;
  LAYER M1 ;
        RECT 2.959 13.692 2.961 16.128 ;
  LAYER M1 ;
        RECT 3.039 13.692 3.041 16.128 ;
  LAYER M1 ;
        RECT 3.119 13.692 3.121 16.128 ;
  LAYER M1 ;
        RECT 3.199 13.692 3.201 16.128 ;
  LAYER M1 ;
        RECT 3.279 13.692 3.281 16.128 ;
  LAYER M1 ;
        RECT 3.359 13.692 3.361 16.128 ;
  LAYER M1 ;
        RECT 3.439 13.692 3.441 16.128 ;
  LAYER M2 ;
        RECT 1.12 16.127 3.52 16.129 ;
  LAYER M2 ;
        RECT 1.12 16.043 3.52 16.045 ;
  LAYER M2 ;
        RECT 1.12 15.959 3.52 15.961 ;
  LAYER M2 ;
        RECT 1.12 15.875 3.52 15.877 ;
  LAYER M2 ;
        RECT 1.12 15.791 3.52 15.793 ;
  LAYER M2 ;
        RECT 1.12 15.707 3.52 15.709 ;
  LAYER M2 ;
        RECT 1.12 15.623 3.52 15.625 ;
  LAYER M2 ;
        RECT 1.12 15.539 3.52 15.541 ;
  LAYER M2 ;
        RECT 1.12 15.455 3.52 15.457 ;
  LAYER M2 ;
        RECT 1.12 15.371 3.52 15.373 ;
  LAYER M2 ;
        RECT 1.12 15.287 3.52 15.289 ;
  LAYER M2 ;
        RECT 1.12 15.203 3.52 15.205 ;
  LAYER M2 ;
        RECT 1.12 15.1195 3.52 15.1215 ;
  LAYER M2 ;
        RECT 1.12 15.035 3.52 15.037 ;
  LAYER M2 ;
        RECT 1.12 14.951 3.52 14.953 ;
  LAYER M2 ;
        RECT 1.12 14.867 3.52 14.869 ;
  LAYER M2 ;
        RECT 1.12 14.783 3.52 14.785 ;
  LAYER M2 ;
        RECT 1.12 14.699 3.52 14.701 ;
  LAYER M2 ;
        RECT 1.12 14.615 3.52 14.617 ;
  LAYER M2 ;
        RECT 1.12 14.531 3.52 14.533 ;
  LAYER M2 ;
        RECT 1.12 14.447 3.52 14.449 ;
  LAYER M2 ;
        RECT 1.12 14.363 3.52 14.365 ;
  LAYER M2 ;
        RECT 1.12 14.279 3.52 14.281 ;
  LAYER M2 ;
        RECT 1.12 14.195 3.52 14.197 ;
  LAYER M2 ;
        RECT 1.12 14.111 3.52 14.113 ;
  LAYER M2 ;
        RECT 1.12 14.027 3.52 14.029 ;
  LAYER M2 ;
        RECT 1.12 13.943 3.52 13.945 ;
  LAYER M2 ;
        RECT 1.12 13.859 3.52 13.861 ;
  LAYER M2 ;
        RECT 1.12 13.775 3.52 13.777 ;
  LAYER M1 ;
        RECT 1.104 10.716 1.136 13.224 ;
  LAYER M1 ;
        RECT 1.168 10.716 1.2 13.224 ;
  LAYER M1 ;
        RECT 1.232 10.716 1.264 13.224 ;
  LAYER M1 ;
        RECT 1.296 10.716 1.328 13.224 ;
  LAYER M1 ;
        RECT 1.36 10.716 1.392 13.224 ;
  LAYER M1 ;
        RECT 1.424 10.716 1.456 13.224 ;
  LAYER M1 ;
        RECT 1.488 10.716 1.52 13.224 ;
  LAYER M1 ;
        RECT 1.552 10.716 1.584 13.224 ;
  LAYER M1 ;
        RECT 1.616 10.716 1.648 13.224 ;
  LAYER M1 ;
        RECT 1.68 10.716 1.712 13.224 ;
  LAYER M1 ;
        RECT 1.744 10.716 1.776 13.224 ;
  LAYER M1 ;
        RECT 1.808 10.716 1.84 13.224 ;
  LAYER M1 ;
        RECT 1.872 10.716 1.904 13.224 ;
  LAYER M1 ;
        RECT 1.936 10.716 1.968 13.224 ;
  LAYER M1 ;
        RECT 2 10.716 2.032 13.224 ;
  LAYER M1 ;
        RECT 2.064 10.716 2.096 13.224 ;
  LAYER M1 ;
        RECT 2.128 10.716 2.16 13.224 ;
  LAYER M1 ;
        RECT 2.192 10.716 2.224 13.224 ;
  LAYER M1 ;
        RECT 2.256 10.716 2.288 13.224 ;
  LAYER M1 ;
        RECT 2.32 10.716 2.352 13.224 ;
  LAYER M1 ;
        RECT 2.384 10.716 2.416 13.224 ;
  LAYER M1 ;
        RECT 2.448 10.716 2.48 13.224 ;
  LAYER M1 ;
        RECT 2.512 10.716 2.544 13.224 ;
  LAYER M1 ;
        RECT 2.576 10.716 2.608 13.224 ;
  LAYER M1 ;
        RECT 2.64 10.716 2.672 13.224 ;
  LAYER M1 ;
        RECT 2.704 10.716 2.736 13.224 ;
  LAYER M1 ;
        RECT 2.768 10.716 2.8 13.224 ;
  LAYER M1 ;
        RECT 2.832 10.716 2.864 13.224 ;
  LAYER M1 ;
        RECT 2.896 10.716 2.928 13.224 ;
  LAYER M1 ;
        RECT 2.96 10.716 2.992 13.224 ;
  LAYER M1 ;
        RECT 3.024 10.716 3.056 13.224 ;
  LAYER M1 ;
        RECT 3.088 10.716 3.12 13.224 ;
  LAYER M1 ;
        RECT 3.152 10.716 3.184 13.224 ;
  LAYER M1 ;
        RECT 3.216 10.716 3.248 13.224 ;
  LAYER M1 ;
        RECT 3.28 10.716 3.312 13.224 ;
  LAYER M1 ;
        RECT 3.344 10.716 3.376 13.224 ;
  LAYER M1 ;
        RECT 3.408 10.716 3.44 13.224 ;
  LAYER M2 ;
        RECT 1.084 13.108 3.556 13.14 ;
  LAYER M2 ;
        RECT 1.084 13.044 3.556 13.076 ;
  LAYER M2 ;
        RECT 1.084 12.98 3.556 13.012 ;
  LAYER M2 ;
        RECT 1.084 12.916 3.556 12.948 ;
  LAYER M2 ;
        RECT 1.084 12.852 3.556 12.884 ;
  LAYER M2 ;
        RECT 1.084 12.788 3.556 12.82 ;
  LAYER M2 ;
        RECT 1.084 12.724 3.556 12.756 ;
  LAYER M2 ;
        RECT 1.084 12.66 3.556 12.692 ;
  LAYER M2 ;
        RECT 1.084 12.596 3.556 12.628 ;
  LAYER M2 ;
        RECT 1.084 12.532 3.556 12.564 ;
  LAYER M2 ;
        RECT 1.084 12.468 3.556 12.5 ;
  LAYER M2 ;
        RECT 1.084 12.404 3.556 12.436 ;
  LAYER M2 ;
        RECT 1.084 12.34 3.556 12.372 ;
  LAYER M2 ;
        RECT 1.084 12.276 3.556 12.308 ;
  LAYER M2 ;
        RECT 1.084 12.212 3.556 12.244 ;
  LAYER M2 ;
        RECT 1.084 12.148 3.556 12.18 ;
  LAYER M2 ;
        RECT 1.084 12.084 3.556 12.116 ;
  LAYER M2 ;
        RECT 1.084 12.02 3.556 12.052 ;
  LAYER M2 ;
        RECT 1.084 11.956 3.556 11.988 ;
  LAYER M2 ;
        RECT 1.084 11.892 3.556 11.924 ;
  LAYER M2 ;
        RECT 1.084 11.828 3.556 11.86 ;
  LAYER M2 ;
        RECT 1.084 11.764 3.556 11.796 ;
  LAYER M2 ;
        RECT 1.084 11.7 3.556 11.732 ;
  LAYER M2 ;
        RECT 1.084 11.636 3.556 11.668 ;
  LAYER M2 ;
        RECT 1.084 11.572 3.556 11.604 ;
  LAYER M2 ;
        RECT 1.084 11.508 3.556 11.54 ;
  LAYER M2 ;
        RECT 1.084 11.444 3.556 11.476 ;
  LAYER M2 ;
        RECT 1.084 11.38 3.556 11.412 ;
  LAYER M2 ;
        RECT 1.084 11.316 3.556 11.348 ;
  LAYER M2 ;
        RECT 1.084 11.252 3.556 11.284 ;
  LAYER M2 ;
        RECT 1.084 11.188 3.556 11.22 ;
  LAYER M2 ;
        RECT 1.084 11.124 3.556 11.156 ;
  LAYER M2 ;
        RECT 1.084 11.06 3.556 11.092 ;
  LAYER M2 ;
        RECT 1.084 10.996 3.556 11.028 ;
  LAYER M2 ;
        RECT 1.084 10.932 3.556 10.964 ;
  LAYER M2 ;
        RECT 1.084 10.868 3.556 10.9 ;
  LAYER M3 ;
        RECT 1.104 10.716 1.136 13.224 ;
  LAYER M3 ;
        RECT 1.168 10.716 1.2 13.224 ;
  LAYER M3 ;
        RECT 1.232 10.716 1.264 13.224 ;
  LAYER M3 ;
        RECT 1.296 10.716 1.328 13.224 ;
  LAYER M3 ;
        RECT 1.36 10.716 1.392 13.224 ;
  LAYER M3 ;
        RECT 1.424 10.716 1.456 13.224 ;
  LAYER M3 ;
        RECT 1.488 10.716 1.52 13.224 ;
  LAYER M3 ;
        RECT 1.552 10.716 1.584 13.224 ;
  LAYER M3 ;
        RECT 1.616 10.716 1.648 13.224 ;
  LAYER M3 ;
        RECT 1.68 10.716 1.712 13.224 ;
  LAYER M3 ;
        RECT 1.744 10.716 1.776 13.224 ;
  LAYER M3 ;
        RECT 1.808 10.716 1.84 13.224 ;
  LAYER M3 ;
        RECT 1.872 10.716 1.904 13.224 ;
  LAYER M3 ;
        RECT 1.936 10.716 1.968 13.224 ;
  LAYER M3 ;
        RECT 2 10.716 2.032 13.224 ;
  LAYER M3 ;
        RECT 2.064 10.716 2.096 13.224 ;
  LAYER M3 ;
        RECT 2.128 10.716 2.16 13.224 ;
  LAYER M3 ;
        RECT 2.192 10.716 2.224 13.224 ;
  LAYER M3 ;
        RECT 2.256 10.716 2.288 13.224 ;
  LAYER M3 ;
        RECT 2.32 10.716 2.352 13.224 ;
  LAYER M3 ;
        RECT 2.384 10.716 2.416 13.224 ;
  LAYER M3 ;
        RECT 2.448 10.716 2.48 13.224 ;
  LAYER M3 ;
        RECT 2.512 10.716 2.544 13.224 ;
  LAYER M3 ;
        RECT 2.576 10.716 2.608 13.224 ;
  LAYER M3 ;
        RECT 2.64 10.716 2.672 13.224 ;
  LAYER M3 ;
        RECT 2.704 10.716 2.736 13.224 ;
  LAYER M3 ;
        RECT 2.768 10.716 2.8 13.224 ;
  LAYER M3 ;
        RECT 2.832 10.716 2.864 13.224 ;
  LAYER M3 ;
        RECT 2.896 10.716 2.928 13.224 ;
  LAYER M3 ;
        RECT 2.96 10.716 2.992 13.224 ;
  LAYER M3 ;
        RECT 3.024 10.716 3.056 13.224 ;
  LAYER M3 ;
        RECT 3.088 10.716 3.12 13.224 ;
  LAYER M3 ;
        RECT 3.152 10.716 3.184 13.224 ;
  LAYER M3 ;
        RECT 3.216 10.716 3.248 13.224 ;
  LAYER M3 ;
        RECT 3.28 10.716 3.312 13.224 ;
  LAYER M3 ;
        RECT 3.344 10.716 3.376 13.224 ;
  LAYER M3 ;
        RECT 3.408 10.716 3.44 13.224 ;
  LAYER M3 ;
        RECT 3.504 10.716 3.536 13.224 ;
  LAYER M1 ;
        RECT 1.119 10.752 1.121 13.188 ;
  LAYER M1 ;
        RECT 1.199 10.752 1.201 13.188 ;
  LAYER M1 ;
        RECT 1.279 10.752 1.281 13.188 ;
  LAYER M1 ;
        RECT 1.359 10.752 1.361 13.188 ;
  LAYER M1 ;
        RECT 1.439 10.752 1.441 13.188 ;
  LAYER M1 ;
        RECT 1.519 10.752 1.521 13.188 ;
  LAYER M1 ;
        RECT 1.599 10.752 1.601 13.188 ;
  LAYER M1 ;
        RECT 1.679 10.752 1.681 13.188 ;
  LAYER M1 ;
        RECT 1.759 10.752 1.761 13.188 ;
  LAYER M1 ;
        RECT 1.839 10.752 1.841 13.188 ;
  LAYER M1 ;
        RECT 1.919 10.752 1.921 13.188 ;
  LAYER M1 ;
        RECT 1.999 10.752 2.001 13.188 ;
  LAYER M1 ;
        RECT 2.079 10.752 2.081 13.188 ;
  LAYER M1 ;
        RECT 2.159 10.752 2.161 13.188 ;
  LAYER M1 ;
        RECT 2.239 10.752 2.241 13.188 ;
  LAYER M1 ;
        RECT 2.319 10.752 2.321 13.188 ;
  LAYER M1 ;
        RECT 2.399 10.752 2.401 13.188 ;
  LAYER M1 ;
        RECT 2.479 10.752 2.481 13.188 ;
  LAYER M1 ;
        RECT 2.559 10.752 2.561 13.188 ;
  LAYER M1 ;
        RECT 2.639 10.752 2.641 13.188 ;
  LAYER M1 ;
        RECT 2.719 10.752 2.721 13.188 ;
  LAYER M1 ;
        RECT 2.799 10.752 2.801 13.188 ;
  LAYER M1 ;
        RECT 2.879 10.752 2.881 13.188 ;
  LAYER M1 ;
        RECT 2.959 10.752 2.961 13.188 ;
  LAYER M1 ;
        RECT 3.039 10.752 3.041 13.188 ;
  LAYER M1 ;
        RECT 3.119 10.752 3.121 13.188 ;
  LAYER M1 ;
        RECT 3.199 10.752 3.201 13.188 ;
  LAYER M1 ;
        RECT 3.279 10.752 3.281 13.188 ;
  LAYER M1 ;
        RECT 3.359 10.752 3.361 13.188 ;
  LAYER M1 ;
        RECT 3.439 10.752 3.441 13.188 ;
  LAYER M2 ;
        RECT 1.12 13.187 3.52 13.189 ;
  LAYER M2 ;
        RECT 1.12 13.103 3.52 13.105 ;
  LAYER M2 ;
        RECT 1.12 13.019 3.52 13.021 ;
  LAYER M2 ;
        RECT 1.12 12.935 3.52 12.937 ;
  LAYER M2 ;
        RECT 1.12 12.851 3.52 12.853 ;
  LAYER M2 ;
        RECT 1.12 12.767 3.52 12.769 ;
  LAYER M2 ;
        RECT 1.12 12.683 3.52 12.685 ;
  LAYER M2 ;
        RECT 1.12 12.599 3.52 12.601 ;
  LAYER M2 ;
        RECT 1.12 12.515 3.52 12.517 ;
  LAYER M2 ;
        RECT 1.12 12.431 3.52 12.433 ;
  LAYER M2 ;
        RECT 1.12 12.347 3.52 12.349 ;
  LAYER M2 ;
        RECT 1.12 12.263 3.52 12.265 ;
  LAYER M2 ;
        RECT 1.12 12.1795 3.52 12.1815 ;
  LAYER M2 ;
        RECT 1.12 12.095 3.52 12.097 ;
  LAYER M2 ;
        RECT 1.12 12.011 3.52 12.013 ;
  LAYER M2 ;
        RECT 1.12 11.927 3.52 11.929 ;
  LAYER M2 ;
        RECT 1.12 11.843 3.52 11.845 ;
  LAYER M2 ;
        RECT 1.12 11.759 3.52 11.761 ;
  LAYER M2 ;
        RECT 1.12 11.675 3.52 11.677 ;
  LAYER M2 ;
        RECT 1.12 11.591 3.52 11.593 ;
  LAYER M2 ;
        RECT 1.12 11.507 3.52 11.509 ;
  LAYER M2 ;
        RECT 1.12 11.423 3.52 11.425 ;
  LAYER M2 ;
        RECT 1.12 11.339 3.52 11.341 ;
  LAYER M2 ;
        RECT 1.12 11.255 3.52 11.257 ;
  LAYER M2 ;
        RECT 1.12 11.171 3.52 11.173 ;
  LAYER M2 ;
        RECT 1.12 11.087 3.52 11.089 ;
  LAYER M2 ;
        RECT 1.12 11.003 3.52 11.005 ;
  LAYER M2 ;
        RECT 1.12 10.919 3.52 10.921 ;
  LAYER M2 ;
        RECT 1.12 10.835 3.52 10.837 ;
  LAYER M1 ;
        RECT 1.104 7.776 1.136 10.284 ;
  LAYER M1 ;
        RECT 1.168 7.776 1.2 10.284 ;
  LAYER M1 ;
        RECT 1.232 7.776 1.264 10.284 ;
  LAYER M1 ;
        RECT 1.296 7.776 1.328 10.284 ;
  LAYER M1 ;
        RECT 1.36 7.776 1.392 10.284 ;
  LAYER M1 ;
        RECT 1.424 7.776 1.456 10.284 ;
  LAYER M1 ;
        RECT 1.488 7.776 1.52 10.284 ;
  LAYER M1 ;
        RECT 1.552 7.776 1.584 10.284 ;
  LAYER M1 ;
        RECT 1.616 7.776 1.648 10.284 ;
  LAYER M1 ;
        RECT 1.68 7.776 1.712 10.284 ;
  LAYER M1 ;
        RECT 1.744 7.776 1.776 10.284 ;
  LAYER M1 ;
        RECT 1.808 7.776 1.84 10.284 ;
  LAYER M1 ;
        RECT 1.872 7.776 1.904 10.284 ;
  LAYER M1 ;
        RECT 1.936 7.776 1.968 10.284 ;
  LAYER M1 ;
        RECT 2 7.776 2.032 10.284 ;
  LAYER M1 ;
        RECT 2.064 7.776 2.096 10.284 ;
  LAYER M1 ;
        RECT 2.128 7.776 2.16 10.284 ;
  LAYER M1 ;
        RECT 2.192 7.776 2.224 10.284 ;
  LAYER M1 ;
        RECT 2.256 7.776 2.288 10.284 ;
  LAYER M1 ;
        RECT 2.32 7.776 2.352 10.284 ;
  LAYER M1 ;
        RECT 2.384 7.776 2.416 10.284 ;
  LAYER M1 ;
        RECT 2.448 7.776 2.48 10.284 ;
  LAYER M1 ;
        RECT 2.512 7.776 2.544 10.284 ;
  LAYER M1 ;
        RECT 2.576 7.776 2.608 10.284 ;
  LAYER M1 ;
        RECT 2.64 7.776 2.672 10.284 ;
  LAYER M1 ;
        RECT 2.704 7.776 2.736 10.284 ;
  LAYER M1 ;
        RECT 2.768 7.776 2.8 10.284 ;
  LAYER M1 ;
        RECT 2.832 7.776 2.864 10.284 ;
  LAYER M1 ;
        RECT 2.896 7.776 2.928 10.284 ;
  LAYER M1 ;
        RECT 2.96 7.776 2.992 10.284 ;
  LAYER M1 ;
        RECT 3.024 7.776 3.056 10.284 ;
  LAYER M1 ;
        RECT 3.088 7.776 3.12 10.284 ;
  LAYER M1 ;
        RECT 3.152 7.776 3.184 10.284 ;
  LAYER M1 ;
        RECT 3.216 7.776 3.248 10.284 ;
  LAYER M1 ;
        RECT 3.28 7.776 3.312 10.284 ;
  LAYER M1 ;
        RECT 3.344 7.776 3.376 10.284 ;
  LAYER M1 ;
        RECT 3.408 7.776 3.44 10.284 ;
  LAYER M2 ;
        RECT 1.084 10.168 3.556 10.2 ;
  LAYER M2 ;
        RECT 1.084 10.104 3.556 10.136 ;
  LAYER M2 ;
        RECT 1.084 10.04 3.556 10.072 ;
  LAYER M2 ;
        RECT 1.084 9.976 3.556 10.008 ;
  LAYER M2 ;
        RECT 1.084 9.912 3.556 9.944 ;
  LAYER M2 ;
        RECT 1.084 9.848 3.556 9.88 ;
  LAYER M2 ;
        RECT 1.084 9.784 3.556 9.816 ;
  LAYER M2 ;
        RECT 1.084 9.72 3.556 9.752 ;
  LAYER M2 ;
        RECT 1.084 9.656 3.556 9.688 ;
  LAYER M2 ;
        RECT 1.084 9.592 3.556 9.624 ;
  LAYER M2 ;
        RECT 1.084 9.528 3.556 9.56 ;
  LAYER M2 ;
        RECT 1.084 9.464 3.556 9.496 ;
  LAYER M2 ;
        RECT 1.084 9.4 3.556 9.432 ;
  LAYER M2 ;
        RECT 1.084 9.336 3.556 9.368 ;
  LAYER M2 ;
        RECT 1.084 9.272 3.556 9.304 ;
  LAYER M2 ;
        RECT 1.084 9.208 3.556 9.24 ;
  LAYER M2 ;
        RECT 1.084 9.144 3.556 9.176 ;
  LAYER M2 ;
        RECT 1.084 9.08 3.556 9.112 ;
  LAYER M2 ;
        RECT 1.084 9.016 3.556 9.048 ;
  LAYER M2 ;
        RECT 1.084 8.952 3.556 8.984 ;
  LAYER M2 ;
        RECT 1.084 8.888 3.556 8.92 ;
  LAYER M2 ;
        RECT 1.084 8.824 3.556 8.856 ;
  LAYER M2 ;
        RECT 1.084 8.76 3.556 8.792 ;
  LAYER M2 ;
        RECT 1.084 8.696 3.556 8.728 ;
  LAYER M2 ;
        RECT 1.084 8.632 3.556 8.664 ;
  LAYER M2 ;
        RECT 1.084 8.568 3.556 8.6 ;
  LAYER M2 ;
        RECT 1.084 8.504 3.556 8.536 ;
  LAYER M2 ;
        RECT 1.084 8.44 3.556 8.472 ;
  LAYER M2 ;
        RECT 1.084 8.376 3.556 8.408 ;
  LAYER M2 ;
        RECT 1.084 8.312 3.556 8.344 ;
  LAYER M2 ;
        RECT 1.084 8.248 3.556 8.28 ;
  LAYER M2 ;
        RECT 1.084 8.184 3.556 8.216 ;
  LAYER M2 ;
        RECT 1.084 8.12 3.556 8.152 ;
  LAYER M2 ;
        RECT 1.084 8.056 3.556 8.088 ;
  LAYER M2 ;
        RECT 1.084 7.992 3.556 8.024 ;
  LAYER M2 ;
        RECT 1.084 7.928 3.556 7.96 ;
  LAYER M3 ;
        RECT 1.104 7.776 1.136 10.284 ;
  LAYER M3 ;
        RECT 1.168 7.776 1.2 10.284 ;
  LAYER M3 ;
        RECT 1.232 7.776 1.264 10.284 ;
  LAYER M3 ;
        RECT 1.296 7.776 1.328 10.284 ;
  LAYER M3 ;
        RECT 1.36 7.776 1.392 10.284 ;
  LAYER M3 ;
        RECT 1.424 7.776 1.456 10.284 ;
  LAYER M3 ;
        RECT 1.488 7.776 1.52 10.284 ;
  LAYER M3 ;
        RECT 1.552 7.776 1.584 10.284 ;
  LAYER M3 ;
        RECT 1.616 7.776 1.648 10.284 ;
  LAYER M3 ;
        RECT 1.68 7.776 1.712 10.284 ;
  LAYER M3 ;
        RECT 1.744 7.776 1.776 10.284 ;
  LAYER M3 ;
        RECT 1.808 7.776 1.84 10.284 ;
  LAYER M3 ;
        RECT 1.872 7.776 1.904 10.284 ;
  LAYER M3 ;
        RECT 1.936 7.776 1.968 10.284 ;
  LAYER M3 ;
        RECT 2 7.776 2.032 10.284 ;
  LAYER M3 ;
        RECT 2.064 7.776 2.096 10.284 ;
  LAYER M3 ;
        RECT 2.128 7.776 2.16 10.284 ;
  LAYER M3 ;
        RECT 2.192 7.776 2.224 10.284 ;
  LAYER M3 ;
        RECT 2.256 7.776 2.288 10.284 ;
  LAYER M3 ;
        RECT 2.32 7.776 2.352 10.284 ;
  LAYER M3 ;
        RECT 2.384 7.776 2.416 10.284 ;
  LAYER M3 ;
        RECT 2.448 7.776 2.48 10.284 ;
  LAYER M3 ;
        RECT 2.512 7.776 2.544 10.284 ;
  LAYER M3 ;
        RECT 2.576 7.776 2.608 10.284 ;
  LAYER M3 ;
        RECT 2.64 7.776 2.672 10.284 ;
  LAYER M3 ;
        RECT 2.704 7.776 2.736 10.284 ;
  LAYER M3 ;
        RECT 2.768 7.776 2.8 10.284 ;
  LAYER M3 ;
        RECT 2.832 7.776 2.864 10.284 ;
  LAYER M3 ;
        RECT 2.896 7.776 2.928 10.284 ;
  LAYER M3 ;
        RECT 2.96 7.776 2.992 10.284 ;
  LAYER M3 ;
        RECT 3.024 7.776 3.056 10.284 ;
  LAYER M3 ;
        RECT 3.088 7.776 3.12 10.284 ;
  LAYER M3 ;
        RECT 3.152 7.776 3.184 10.284 ;
  LAYER M3 ;
        RECT 3.216 7.776 3.248 10.284 ;
  LAYER M3 ;
        RECT 3.28 7.776 3.312 10.284 ;
  LAYER M3 ;
        RECT 3.344 7.776 3.376 10.284 ;
  LAYER M3 ;
        RECT 3.408 7.776 3.44 10.284 ;
  LAYER M3 ;
        RECT 3.504 7.776 3.536 10.284 ;
  LAYER M1 ;
        RECT 1.119 7.812 1.121 10.248 ;
  LAYER M1 ;
        RECT 1.199 7.812 1.201 10.248 ;
  LAYER M1 ;
        RECT 1.279 7.812 1.281 10.248 ;
  LAYER M1 ;
        RECT 1.359 7.812 1.361 10.248 ;
  LAYER M1 ;
        RECT 1.439 7.812 1.441 10.248 ;
  LAYER M1 ;
        RECT 1.519 7.812 1.521 10.248 ;
  LAYER M1 ;
        RECT 1.599 7.812 1.601 10.248 ;
  LAYER M1 ;
        RECT 1.679 7.812 1.681 10.248 ;
  LAYER M1 ;
        RECT 1.759 7.812 1.761 10.248 ;
  LAYER M1 ;
        RECT 1.839 7.812 1.841 10.248 ;
  LAYER M1 ;
        RECT 1.919 7.812 1.921 10.248 ;
  LAYER M1 ;
        RECT 1.999 7.812 2.001 10.248 ;
  LAYER M1 ;
        RECT 2.079 7.812 2.081 10.248 ;
  LAYER M1 ;
        RECT 2.159 7.812 2.161 10.248 ;
  LAYER M1 ;
        RECT 2.239 7.812 2.241 10.248 ;
  LAYER M1 ;
        RECT 2.319 7.812 2.321 10.248 ;
  LAYER M1 ;
        RECT 2.399 7.812 2.401 10.248 ;
  LAYER M1 ;
        RECT 2.479 7.812 2.481 10.248 ;
  LAYER M1 ;
        RECT 2.559 7.812 2.561 10.248 ;
  LAYER M1 ;
        RECT 2.639 7.812 2.641 10.248 ;
  LAYER M1 ;
        RECT 2.719 7.812 2.721 10.248 ;
  LAYER M1 ;
        RECT 2.799 7.812 2.801 10.248 ;
  LAYER M1 ;
        RECT 2.879 7.812 2.881 10.248 ;
  LAYER M1 ;
        RECT 2.959 7.812 2.961 10.248 ;
  LAYER M1 ;
        RECT 3.039 7.812 3.041 10.248 ;
  LAYER M1 ;
        RECT 3.119 7.812 3.121 10.248 ;
  LAYER M1 ;
        RECT 3.199 7.812 3.201 10.248 ;
  LAYER M1 ;
        RECT 3.279 7.812 3.281 10.248 ;
  LAYER M1 ;
        RECT 3.359 7.812 3.361 10.248 ;
  LAYER M1 ;
        RECT 3.439 7.812 3.441 10.248 ;
  LAYER M2 ;
        RECT 1.12 10.247 3.52 10.249 ;
  LAYER M2 ;
        RECT 1.12 10.163 3.52 10.165 ;
  LAYER M2 ;
        RECT 1.12 10.079 3.52 10.081 ;
  LAYER M2 ;
        RECT 1.12 9.995 3.52 9.997 ;
  LAYER M2 ;
        RECT 1.12 9.911 3.52 9.913 ;
  LAYER M2 ;
        RECT 1.12 9.827 3.52 9.829 ;
  LAYER M2 ;
        RECT 1.12 9.743 3.52 9.745 ;
  LAYER M2 ;
        RECT 1.12 9.659 3.52 9.661 ;
  LAYER M2 ;
        RECT 1.12 9.575 3.52 9.577 ;
  LAYER M2 ;
        RECT 1.12 9.491 3.52 9.493 ;
  LAYER M2 ;
        RECT 1.12 9.407 3.52 9.409 ;
  LAYER M2 ;
        RECT 1.12 9.323 3.52 9.325 ;
  LAYER M2 ;
        RECT 1.12 9.2395 3.52 9.2415 ;
  LAYER M2 ;
        RECT 1.12 9.155 3.52 9.157 ;
  LAYER M2 ;
        RECT 1.12 9.071 3.52 9.073 ;
  LAYER M2 ;
        RECT 1.12 8.987 3.52 8.989 ;
  LAYER M2 ;
        RECT 1.12 8.903 3.52 8.905 ;
  LAYER M2 ;
        RECT 1.12 8.819 3.52 8.821 ;
  LAYER M2 ;
        RECT 1.12 8.735 3.52 8.737 ;
  LAYER M2 ;
        RECT 1.12 8.651 3.52 8.653 ;
  LAYER M2 ;
        RECT 1.12 8.567 3.52 8.569 ;
  LAYER M2 ;
        RECT 1.12 8.483 3.52 8.485 ;
  LAYER M2 ;
        RECT 1.12 8.399 3.52 8.401 ;
  LAYER M2 ;
        RECT 1.12 8.315 3.52 8.317 ;
  LAYER M2 ;
        RECT 1.12 8.231 3.52 8.233 ;
  LAYER M2 ;
        RECT 1.12 8.147 3.52 8.149 ;
  LAYER M2 ;
        RECT 1.12 8.063 3.52 8.065 ;
  LAYER M2 ;
        RECT 1.12 7.979 3.52 7.981 ;
  LAYER M2 ;
        RECT 1.12 7.895 3.52 7.897 ;
  LAYER M1 ;
        RECT 1.104 4.836 1.136 7.344 ;
  LAYER M1 ;
        RECT 1.168 4.836 1.2 7.344 ;
  LAYER M1 ;
        RECT 1.232 4.836 1.264 7.344 ;
  LAYER M1 ;
        RECT 1.296 4.836 1.328 7.344 ;
  LAYER M1 ;
        RECT 1.36 4.836 1.392 7.344 ;
  LAYER M1 ;
        RECT 1.424 4.836 1.456 7.344 ;
  LAYER M1 ;
        RECT 1.488 4.836 1.52 7.344 ;
  LAYER M1 ;
        RECT 1.552 4.836 1.584 7.344 ;
  LAYER M1 ;
        RECT 1.616 4.836 1.648 7.344 ;
  LAYER M1 ;
        RECT 1.68 4.836 1.712 7.344 ;
  LAYER M1 ;
        RECT 1.744 4.836 1.776 7.344 ;
  LAYER M1 ;
        RECT 1.808 4.836 1.84 7.344 ;
  LAYER M1 ;
        RECT 1.872 4.836 1.904 7.344 ;
  LAYER M1 ;
        RECT 1.936 4.836 1.968 7.344 ;
  LAYER M1 ;
        RECT 2 4.836 2.032 7.344 ;
  LAYER M1 ;
        RECT 2.064 4.836 2.096 7.344 ;
  LAYER M1 ;
        RECT 2.128 4.836 2.16 7.344 ;
  LAYER M1 ;
        RECT 2.192 4.836 2.224 7.344 ;
  LAYER M1 ;
        RECT 2.256 4.836 2.288 7.344 ;
  LAYER M1 ;
        RECT 2.32 4.836 2.352 7.344 ;
  LAYER M1 ;
        RECT 2.384 4.836 2.416 7.344 ;
  LAYER M1 ;
        RECT 2.448 4.836 2.48 7.344 ;
  LAYER M1 ;
        RECT 2.512 4.836 2.544 7.344 ;
  LAYER M1 ;
        RECT 2.576 4.836 2.608 7.344 ;
  LAYER M1 ;
        RECT 2.64 4.836 2.672 7.344 ;
  LAYER M1 ;
        RECT 2.704 4.836 2.736 7.344 ;
  LAYER M1 ;
        RECT 2.768 4.836 2.8 7.344 ;
  LAYER M1 ;
        RECT 2.832 4.836 2.864 7.344 ;
  LAYER M1 ;
        RECT 2.896 4.836 2.928 7.344 ;
  LAYER M1 ;
        RECT 2.96 4.836 2.992 7.344 ;
  LAYER M1 ;
        RECT 3.024 4.836 3.056 7.344 ;
  LAYER M1 ;
        RECT 3.088 4.836 3.12 7.344 ;
  LAYER M1 ;
        RECT 3.152 4.836 3.184 7.344 ;
  LAYER M1 ;
        RECT 3.216 4.836 3.248 7.344 ;
  LAYER M1 ;
        RECT 3.28 4.836 3.312 7.344 ;
  LAYER M1 ;
        RECT 3.344 4.836 3.376 7.344 ;
  LAYER M1 ;
        RECT 3.408 4.836 3.44 7.344 ;
  LAYER M2 ;
        RECT 1.084 7.228 3.556 7.26 ;
  LAYER M2 ;
        RECT 1.084 7.164 3.556 7.196 ;
  LAYER M2 ;
        RECT 1.084 7.1 3.556 7.132 ;
  LAYER M2 ;
        RECT 1.084 7.036 3.556 7.068 ;
  LAYER M2 ;
        RECT 1.084 6.972 3.556 7.004 ;
  LAYER M2 ;
        RECT 1.084 6.908 3.556 6.94 ;
  LAYER M2 ;
        RECT 1.084 6.844 3.556 6.876 ;
  LAYER M2 ;
        RECT 1.084 6.78 3.556 6.812 ;
  LAYER M2 ;
        RECT 1.084 6.716 3.556 6.748 ;
  LAYER M2 ;
        RECT 1.084 6.652 3.556 6.684 ;
  LAYER M2 ;
        RECT 1.084 6.588 3.556 6.62 ;
  LAYER M2 ;
        RECT 1.084 6.524 3.556 6.556 ;
  LAYER M2 ;
        RECT 1.084 6.46 3.556 6.492 ;
  LAYER M2 ;
        RECT 1.084 6.396 3.556 6.428 ;
  LAYER M2 ;
        RECT 1.084 6.332 3.556 6.364 ;
  LAYER M2 ;
        RECT 1.084 6.268 3.556 6.3 ;
  LAYER M2 ;
        RECT 1.084 6.204 3.556 6.236 ;
  LAYER M2 ;
        RECT 1.084 6.14 3.556 6.172 ;
  LAYER M2 ;
        RECT 1.084 6.076 3.556 6.108 ;
  LAYER M2 ;
        RECT 1.084 6.012 3.556 6.044 ;
  LAYER M2 ;
        RECT 1.084 5.948 3.556 5.98 ;
  LAYER M2 ;
        RECT 1.084 5.884 3.556 5.916 ;
  LAYER M2 ;
        RECT 1.084 5.82 3.556 5.852 ;
  LAYER M2 ;
        RECT 1.084 5.756 3.556 5.788 ;
  LAYER M2 ;
        RECT 1.084 5.692 3.556 5.724 ;
  LAYER M2 ;
        RECT 1.084 5.628 3.556 5.66 ;
  LAYER M2 ;
        RECT 1.084 5.564 3.556 5.596 ;
  LAYER M2 ;
        RECT 1.084 5.5 3.556 5.532 ;
  LAYER M2 ;
        RECT 1.084 5.436 3.556 5.468 ;
  LAYER M2 ;
        RECT 1.084 5.372 3.556 5.404 ;
  LAYER M2 ;
        RECT 1.084 5.308 3.556 5.34 ;
  LAYER M2 ;
        RECT 1.084 5.244 3.556 5.276 ;
  LAYER M2 ;
        RECT 1.084 5.18 3.556 5.212 ;
  LAYER M2 ;
        RECT 1.084 5.116 3.556 5.148 ;
  LAYER M2 ;
        RECT 1.084 5.052 3.556 5.084 ;
  LAYER M2 ;
        RECT 1.084 4.988 3.556 5.02 ;
  LAYER M3 ;
        RECT 1.104 4.836 1.136 7.344 ;
  LAYER M3 ;
        RECT 1.168 4.836 1.2 7.344 ;
  LAYER M3 ;
        RECT 1.232 4.836 1.264 7.344 ;
  LAYER M3 ;
        RECT 1.296 4.836 1.328 7.344 ;
  LAYER M3 ;
        RECT 1.36 4.836 1.392 7.344 ;
  LAYER M3 ;
        RECT 1.424 4.836 1.456 7.344 ;
  LAYER M3 ;
        RECT 1.488 4.836 1.52 7.344 ;
  LAYER M3 ;
        RECT 1.552 4.836 1.584 7.344 ;
  LAYER M3 ;
        RECT 1.616 4.836 1.648 7.344 ;
  LAYER M3 ;
        RECT 1.68 4.836 1.712 7.344 ;
  LAYER M3 ;
        RECT 1.744 4.836 1.776 7.344 ;
  LAYER M3 ;
        RECT 1.808 4.836 1.84 7.344 ;
  LAYER M3 ;
        RECT 1.872 4.836 1.904 7.344 ;
  LAYER M3 ;
        RECT 1.936 4.836 1.968 7.344 ;
  LAYER M3 ;
        RECT 2 4.836 2.032 7.344 ;
  LAYER M3 ;
        RECT 2.064 4.836 2.096 7.344 ;
  LAYER M3 ;
        RECT 2.128 4.836 2.16 7.344 ;
  LAYER M3 ;
        RECT 2.192 4.836 2.224 7.344 ;
  LAYER M3 ;
        RECT 2.256 4.836 2.288 7.344 ;
  LAYER M3 ;
        RECT 2.32 4.836 2.352 7.344 ;
  LAYER M3 ;
        RECT 2.384 4.836 2.416 7.344 ;
  LAYER M3 ;
        RECT 2.448 4.836 2.48 7.344 ;
  LAYER M3 ;
        RECT 2.512 4.836 2.544 7.344 ;
  LAYER M3 ;
        RECT 2.576 4.836 2.608 7.344 ;
  LAYER M3 ;
        RECT 2.64 4.836 2.672 7.344 ;
  LAYER M3 ;
        RECT 2.704 4.836 2.736 7.344 ;
  LAYER M3 ;
        RECT 2.768 4.836 2.8 7.344 ;
  LAYER M3 ;
        RECT 2.832 4.836 2.864 7.344 ;
  LAYER M3 ;
        RECT 2.896 4.836 2.928 7.344 ;
  LAYER M3 ;
        RECT 2.96 4.836 2.992 7.344 ;
  LAYER M3 ;
        RECT 3.024 4.836 3.056 7.344 ;
  LAYER M3 ;
        RECT 3.088 4.836 3.12 7.344 ;
  LAYER M3 ;
        RECT 3.152 4.836 3.184 7.344 ;
  LAYER M3 ;
        RECT 3.216 4.836 3.248 7.344 ;
  LAYER M3 ;
        RECT 3.28 4.836 3.312 7.344 ;
  LAYER M3 ;
        RECT 3.344 4.836 3.376 7.344 ;
  LAYER M3 ;
        RECT 3.408 4.836 3.44 7.344 ;
  LAYER M3 ;
        RECT 3.504 4.836 3.536 7.344 ;
  LAYER M1 ;
        RECT 1.119 4.872 1.121 7.308 ;
  LAYER M1 ;
        RECT 1.199 4.872 1.201 7.308 ;
  LAYER M1 ;
        RECT 1.279 4.872 1.281 7.308 ;
  LAYER M1 ;
        RECT 1.359 4.872 1.361 7.308 ;
  LAYER M1 ;
        RECT 1.439 4.872 1.441 7.308 ;
  LAYER M1 ;
        RECT 1.519 4.872 1.521 7.308 ;
  LAYER M1 ;
        RECT 1.599 4.872 1.601 7.308 ;
  LAYER M1 ;
        RECT 1.679 4.872 1.681 7.308 ;
  LAYER M1 ;
        RECT 1.759 4.872 1.761 7.308 ;
  LAYER M1 ;
        RECT 1.839 4.872 1.841 7.308 ;
  LAYER M1 ;
        RECT 1.919 4.872 1.921 7.308 ;
  LAYER M1 ;
        RECT 1.999 4.872 2.001 7.308 ;
  LAYER M1 ;
        RECT 2.079 4.872 2.081 7.308 ;
  LAYER M1 ;
        RECT 2.159 4.872 2.161 7.308 ;
  LAYER M1 ;
        RECT 2.239 4.872 2.241 7.308 ;
  LAYER M1 ;
        RECT 2.319 4.872 2.321 7.308 ;
  LAYER M1 ;
        RECT 2.399 4.872 2.401 7.308 ;
  LAYER M1 ;
        RECT 2.479 4.872 2.481 7.308 ;
  LAYER M1 ;
        RECT 2.559 4.872 2.561 7.308 ;
  LAYER M1 ;
        RECT 2.639 4.872 2.641 7.308 ;
  LAYER M1 ;
        RECT 2.719 4.872 2.721 7.308 ;
  LAYER M1 ;
        RECT 2.799 4.872 2.801 7.308 ;
  LAYER M1 ;
        RECT 2.879 4.872 2.881 7.308 ;
  LAYER M1 ;
        RECT 2.959 4.872 2.961 7.308 ;
  LAYER M1 ;
        RECT 3.039 4.872 3.041 7.308 ;
  LAYER M1 ;
        RECT 3.119 4.872 3.121 7.308 ;
  LAYER M1 ;
        RECT 3.199 4.872 3.201 7.308 ;
  LAYER M1 ;
        RECT 3.279 4.872 3.281 7.308 ;
  LAYER M1 ;
        RECT 3.359 4.872 3.361 7.308 ;
  LAYER M1 ;
        RECT 3.439 4.872 3.441 7.308 ;
  LAYER M2 ;
        RECT 1.12 7.307 3.52 7.309 ;
  LAYER M2 ;
        RECT 1.12 7.223 3.52 7.225 ;
  LAYER M2 ;
        RECT 1.12 7.139 3.52 7.141 ;
  LAYER M2 ;
        RECT 1.12 7.055 3.52 7.057 ;
  LAYER M2 ;
        RECT 1.12 6.971 3.52 6.973 ;
  LAYER M2 ;
        RECT 1.12 6.887 3.52 6.889 ;
  LAYER M2 ;
        RECT 1.12 6.803 3.52 6.805 ;
  LAYER M2 ;
        RECT 1.12 6.719 3.52 6.721 ;
  LAYER M2 ;
        RECT 1.12 6.635 3.52 6.637 ;
  LAYER M2 ;
        RECT 1.12 6.551 3.52 6.553 ;
  LAYER M2 ;
        RECT 1.12 6.467 3.52 6.469 ;
  LAYER M2 ;
        RECT 1.12 6.383 3.52 6.385 ;
  LAYER M2 ;
        RECT 1.12 6.2995 3.52 6.3015 ;
  LAYER M2 ;
        RECT 1.12 6.215 3.52 6.217 ;
  LAYER M2 ;
        RECT 1.12 6.131 3.52 6.133 ;
  LAYER M2 ;
        RECT 1.12 6.047 3.52 6.049 ;
  LAYER M2 ;
        RECT 1.12 5.963 3.52 5.965 ;
  LAYER M2 ;
        RECT 1.12 5.879 3.52 5.881 ;
  LAYER M2 ;
        RECT 1.12 5.795 3.52 5.797 ;
  LAYER M2 ;
        RECT 1.12 5.711 3.52 5.713 ;
  LAYER M2 ;
        RECT 1.12 5.627 3.52 5.629 ;
  LAYER M2 ;
        RECT 1.12 5.543 3.52 5.545 ;
  LAYER M2 ;
        RECT 1.12 5.459 3.52 5.461 ;
  LAYER M2 ;
        RECT 1.12 5.375 3.52 5.377 ;
  LAYER M2 ;
        RECT 1.12 5.291 3.52 5.293 ;
  LAYER M2 ;
        RECT 1.12 5.207 3.52 5.209 ;
  LAYER M2 ;
        RECT 1.12 5.123 3.52 5.125 ;
  LAYER M2 ;
        RECT 1.12 5.039 3.52 5.041 ;
  LAYER M2 ;
        RECT 1.12 4.955 3.52 4.957 ;
  LAYER M1 ;
        RECT 1.104 1.896 1.136 4.404 ;
  LAYER M1 ;
        RECT 1.168 1.896 1.2 4.404 ;
  LAYER M1 ;
        RECT 1.232 1.896 1.264 4.404 ;
  LAYER M1 ;
        RECT 1.296 1.896 1.328 4.404 ;
  LAYER M1 ;
        RECT 1.36 1.896 1.392 4.404 ;
  LAYER M1 ;
        RECT 1.424 1.896 1.456 4.404 ;
  LAYER M1 ;
        RECT 1.488 1.896 1.52 4.404 ;
  LAYER M1 ;
        RECT 1.552 1.896 1.584 4.404 ;
  LAYER M1 ;
        RECT 1.616 1.896 1.648 4.404 ;
  LAYER M1 ;
        RECT 1.68 1.896 1.712 4.404 ;
  LAYER M1 ;
        RECT 1.744 1.896 1.776 4.404 ;
  LAYER M1 ;
        RECT 1.808 1.896 1.84 4.404 ;
  LAYER M1 ;
        RECT 1.872 1.896 1.904 4.404 ;
  LAYER M1 ;
        RECT 1.936 1.896 1.968 4.404 ;
  LAYER M1 ;
        RECT 2 1.896 2.032 4.404 ;
  LAYER M1 ;
        RECT 2.064 1.896 2.096 4.404 ;
  LAYER M1 ;
        RECT 2.128 1.896 2.16 4.404 ;
  LAYER M1 ;
        RECT 2.192 1.896 2.224 4.404 ;
  LAYER M1 ;
        RECT 2.256 1.896 2.288 4.404 ;
  LAYER M1 ;
        RECT 2.32 1.896 2.352 4.404 ;
  LAYER M1 ;
        RECT 2.384 1.896 2.416 4.404 ;
  LAYER M1 ;
        RECT 2.448 1.896 2.48 4.404 ;
  LAYER M1 ;
        RECT 2.512 1.896 2.544 4.404 ;
  LAYER M1 ;
        RECT 2.576 1.896 2.608 4.404 ;
  LAYER M1 ;
        RECT 2.64 1.896 2.672 4.404 ;
  LAYER M1 ;
        RECT 2.704 1.896 2.736 4.404 ;
  LAYER M1 ;
        RECT 2.768 1.896 2.8 4.404 ;
  LAYER M1 ;
        RECT 2.832 1.896 2.864 4.404 ;
  LAYER M1 ;
        RECT 2.896 1.896 2.928 4.404 ;
  LAYER M1 ;
        RECT 2.96 1.896 2.992 4.404 ;
  LAYER M1 ;
        RECT 3.024 1.896 3.056 4.404 ;
  LAYER M1 ;
        RECT 3.088 1.896 3.12 4.404 ;
  LAYER M1 ;
        RECT 3.152 1.896 3.184 4.404 ;
  LAYER M1 ;
        RECT 3.216 1.896 3.248 4.404 ;
  LAYER M1 ;
        RECT 3.28 1.896 3.312 4.404 ;
  LAYER M1 ;
        RECT 3.344 1.896 3.376 4.404 ;
  LAYER M1 ;
        RECT 3.408 1.896 3.44 4.404 ;
  LAYER M2 ;
        RECT 1.084 4.288 3.556 4.32 ;
  LAYER M2 ;
        RECT 1.084 4.224 3.556 4.256 ;
  LAYER M2 ;
        RECT 1.084 4.16 3.556 4.192 ;
  LAYER M2 ;
        RECT 1.084 4.096 3.556 4.128 ;
  LAYER M2 ;
        RECT 1.084 4.032 3.556 4.064 ;
  LAYER M2 ;
        RECT 1.084 3.968 3.556 4 ;
  LAYER M2 ;
        RECT 1.084 3.904 3.556 3.936 ;
  LAYER M2 ;
        RECT 1.084 3.84 3.556 3.872 ;
  LAYER M2 ;
        RECT 1.084 3.776 3.556 3.808 ;
  LAYER M2 ;
        RECT 1.084 3.712 3.556 3.744 ;
  LAYER M2 ;
        RECT 1.084 3.648 3.556 3.68 ;
  LAYER M2 ;
        RECT 1.084 3.584 3.556 3.616 ;
  LAYER M2 ;
        RECT 1.084 3.52 3.556 3.552 ;
  LAYER M2 ;
        RECT 1.084 3.456 3.556 3.488 ;
  LAYER M2 ;
        RECT 1.084 3.392 3.556 3.424 ;
  LAYER M2 ;
        RECT 1.084 3.328 3.556 3.36 ;
  LAYER M2 ;
        RECT 1.084 3.264 3.556 3.296 ;
  LAYER M2 ;
        RECT 1.084 3.2 3.556 3.232 ;
  LAYER M2 ;
        RECT 1.084 3.136 3.556 3.168 ;
  LAYER M2 ;
        RECT 1.084 3.072 3.556 3.104 ;
  LAYER M2 ;
        RECT 1.084 3.008 3.556 3.04 ;
  LAYER M2 ;
        RECT 1.084 2.944 3.556 2.976 ;
  LAYER M2 ;
        RECT 1.084 2.88 3.556 2.912 ;
  LAYER M2 ;
        RECT 1.084 2.816 3.556 2.848 ;
  LAYER M2 ;
        RECT 1.084 2.752 3.556 2.784 ;
  LAYER M2 ;
        RECT 1.084 2.688 3.556 2.72 ;
  LAYER M2 ;
        RECT 1.084 2.624 3.556 2.656 ;
  LAYER M2 ;
        RECT 1.084 2.56 3.556 2.592 ;
  LAYER M2 ;
        RECT 1.084 2.496 3.556 2.528 ;
  LAYER M2 ;
        RECT 1.084 2.432 3.556 2.464 ;
  LAYER M2 ;
        RECT 1.084 2.368 3.556 2.4 ;
  LAYER M2 ;
        RECT 1.084 2.304 3.556 2.336 ;
  LAYER M2 ;
        RECT 1.084 2.24 3.556 2.272 ;
  LAYER M2 ;
        RECT 1.084 2.176 3.556 2.208 ;
  LAYER M2 ;
        RECT 1.084 2.112 3.556 2.144 ;
  LAYER M2 ;
        RECT 1.084 2.048 3.556 2.08 ;
  LAYER M3 ;
        RECT 1.104 1.896 1.136 4.404 ;
  LAYER M3 ;
        RECT 1.168 1.896 1.2 4.404 ;
  LAYER M3 ;
        RECT 1.232 1.896 1.264 4.404 ;
  LAYER M3 ;
        RECT 1.296 1.896 1.328 4.404 ;
  LAYER M3 ;
        RECT 1.36 1.896 1.392 4.404 ;
  LAYER M3 ;
        RECT 1.424 1.896 1.456 4.404 ;
  LAYER M3 ;
        RECT 1.488 1.896 1.52 4.404 ;
  LAYER M3 ;
        RECT 1.552 1.896 1.584 4.404 ;
  LAYER M3 ;
        RECT 1.616 1.896 1.648 4.404 ;
  LAYER M3 ;
        RECT 1.68 1.896 1.712 4.404 ;
  LAYER M3 ;
        RECT 1.744 1.896 1.776 4.404 ;
  LAYER M3 ;
        RECT 1.808 1.896 1.84 4.404 ;
  LAYER M3 ;
        RECT 1.872 1.896 1.904 4.404 ;
  LAYER M3 ;
        RECT 1.936 1.896 1.968 4.404 ;
  LAYER M3 ;
        RECT 2 1.896 2.032 4.404 ;
  LAYER M3 ;
        RECT 2.064 1.896 2.096 4.404 ;
  LAYER M3 ;
        RECT 2.128 1.896 2.16 4.404 ;
  LAYER M3 ;
        RECT 2.192 1.896 2.224 4.404 ;
  LAYER M3 ;
        RECT 2.256 1.896 2.288 4.404 ;
  LAYER M3 ;
        RECT 2.32 1.896 2.352 4.404 ;
  LAYER M3 ;
        RECT 2.384 1.896 2.416 4.404 ;
  LAYER M3 ;
        RECT 2.448 1.896 2.48 4.404 ;
  LAYER M3 ;
        RECT 2.512 1.896 2.544 4.404 ;
  LAYER M3 ;
        RECT 2.576 1.896 2.608 4.404 ;
  LAYER M3 ;
        RECT 2.64 1.896 2.672 4.404 ;
  LAYER M3 ;
        RECT 2.704 1.896 2.736 4.404 ;
  LAYER M3 ;
        RECT 2.768 1.896 2.8 4.404 ;
  LAYER M3 ;
        RECT 2.832 1.896 2.864 4.404 ;
  LAYER M3 ;
        RECT 2.896 1.896 2.928 4.404 ;
  LAYER M3 ;
        RECT 2.96 1.896 2.992 4.404 ;
  LAYER M3 ;
        RECT 3.024 1.896 3.056 4.404 ;
  LAYER M3 ;
        RECT 3.088 1.896 3.12 4.404 ;
  LAYER M3 ;
        RECT 3.152 1.896 3.184 4.404 ;
  LAYER M3 ;
        RECT 3.216 1.896 3.248 4.404 ;
  LAYER M3 ;
        RECT 3.28 1.896 3.312 4.404 ;
  LAYER M3 ;
        RECT 3.344 1.896 3.376 4.404 ;
  LAYER M3 ;
        RECT 3.408 1.896 3.44 4.404 ;
  LAYER M3 ;
        RECT 3.504 1.896 3.536 4.404 ;
  LAYER M1 ;
        RECT 1.119 1.932 1.121 4.368 ;
  LAYER M1 ;
        RECT 1.199 1.932 1.201 4.368 ;
  LAYER M1 ;
        RECT 1.279 1.932 1.281 4.368 ;
  LAYER M1 ;
        RECT 1.359 1.932 1.361 4.368 ;
  LAYER M1 ;
        RECT 1.439 1.932 1.441 4.368 ;
  LAYER M1 ;
        RECT 1.519 1.932 1.521 4.368 ;
  LAYER M1 ;
        RECT 1.599 1.932 1.601 4.368 ;
  LAYER M1 ;
        RECT 1.679 1.932 1.681 4.368 ;
  LAYER M1 ;
        RECT 1.759 1.932 1.761 4.368 ;
  LAYER M1 ;
        RECT 1.839 1.932 1.841 4.368 ;
  LAYER M1 ;
        RECT 1.919 1.932 1.921 4.368 ;
  LAYER M1 ;
        RECT 1.999 1.932 2.001 4.368 ;
  LAYER M1 ;
        RECT 2.079 1.932 2.081 4.368 ;
  LAYER M1 ;
        RECT 2.159 1.932 2.161 4.368 ;
  LAYER M1 ;
        RECT 2.239 1.932 2.241 4.368 ;
  LAYER M1 ;
        RECT 2.319 1.932 2.321 4.368 ;
  LAYER M1 ;
        RECT 2.399 1.932 2.401 4.368 ;
  LAYER M1 ;
        RECT 2.479 1.932 2.481 4.368 ;
  LAYER M1 ;
        RECT 2.559 1.932 2.561 4.368 ;
  LAYER M1 ;
        RECT 2.639 1.932 2.641 4.368 ;
  LAYER M1 ;
        RECT 2.719 1.932 2.721 4.368 ;
  LAYER M1 ;
        RECT 2.799 1.932 2.801 4.368 ;
  LAYER M1 ;
        RECT 2.879 1.932 2.881 4.368 ;
  LAYER M1 ;
        RECT 2.959 1.932 2.961 4.368 ;
  LAYER M1 ;
        RECT 3.039 1.932 3.041 4.368 ;
  LAYER M1 ;
        RECT 3.119 1.932 3.121 4.368 ;
  LAYER M1 ;
        RECT 3.199 1.932 3.201 4.368 ;
  LAYER M1 ;
        RECT 3.279 1.932 3.281 4.368 ;
  LAYER M1 ;
        RECT 3.359 1.932 3.361 4.368 ;
  LAYER M1 ;
        RECT 3.439 1.932 3.441 4.368 ;
  LAYER M2 ;
        RECT 1.12 4.367 3.52 4.369 ;
  LAYER M2 ;
        RECT 1.12 4.283 3.52 4.285 ;
  LAYER M2 ;
        RECT 1.12 4.199 3.52 4.201 ;
  LAYER M2 ;
        RECT 1.12 4.115 3.52 4.117 ;
  LAYER M2 ;
        RECT 1.12 4.031 3.52 4.033 ;
  LAYER M2 ;
        RECT 1.12 3.947 3.52 3.949 ;
  LAYER M2 ;
        RECT 1.12 3.863 3.52 3.865 ;
  LAYER M2 ;
        RECT 1.12 3.779 3.52 3.781 ;
  LAYER M2 ;
        RECT 1.12 3.695 3.52 3.697 ;
  LAYER M2 ;
        RECT 1.12 3.611 3.52 3.613 ;
  LAYER M2 ;
        RECT 1.12 3.527 3.52 3.529 ;
  LAYER M2 ;
        RECT 1.12 3.443 3.52 3.445 ;
  LAYER M2 ;
        RECT 1.12 3.3595 3.52 3.3615 ;
  LAYER M2 ;
        RECT 1.12 3.275 3.52 3.277 ;
  LAYER M2 ;
        RECT 1.12 3.191 3.52 3.193 ;
  LAYER M2 ;
        RECT 1.12 3.107 3.52 3.109 ;
  LAYER M2 ;
        RECT 1.12 3.023 3.52 3.025 ;
  LAYER M2 ;
        RECT 1.12 2.939 3.52 2.941 ;
  LAYER M2 ;
        RECT 1.12 2.855 3.52 2.857 ;
  LAYER M2 ;
        RECT 1.12 2.771 3.52 2.773 ;
  LAYER M2 ;
        RECT 1.12 2.687 3.52 2.689 ;
  LAYER M2 ;
        RECT 1.12 2.603 3.52 2.605 ;
  LAYER M2 ;
        RECT 1.12 2.519 3.52 2.521 ;
  LAYER M2 ;
        RECT 1.12 2.435 3.52 2.437 ;
  LAYER M2 ;
        RECT 1.12 2.351 3.52 2.353 ;
  LAYER M2 ;
        RECT 1.12 2.267 3.52 2.269 ;
  LAYER M2 ;
        RECT 1.12 2.183 3.52 2.185 ;
  LAYER M2 ;
        RECT 1.12 2.099 3.52 2.101 ;
  LAYER M2 ;
        RECT 1.12 2.015 3.52 2.017 ;
  LAYER M1 ;
        RECT 3.984 13.656 4.016 16.164 ;
  LAYER M1 ;
        RECT 4.048 13.656 4.08 16.164 ;
  LAYER M1 ;
        RECT 4.112 13.656 4.144 16.164 ;
  LAYER M1 ;
        RECT 4.176 13.656 4.208 16.164 ;
  LAYER M1 ;
        RECT 4.24 13.656 4.272 16.164 ;
  LAYER M1 ;
        RECT 4.304 13.656 4.336 16.164 ;
  LAYER M1 ;
        RECT 4.368 13.656 4.4 16.164 ;
  LAYER M1 ;
        RECT 4.432 13.656 4.464 16.164 ;
  LAYER M1 ;
        RECT 4.496 13.656 4.528 16.164 ;
  LAYER M1 ;
        RECT 4.56 13.656 4.592 16.164 ;
  LAYER M1 ;
        RECT 4.624 13.656 4.656 16.164 ;
  LAYER M1 ;
        RECT 4.688 13.656 4.72 16.164 ;
  LAYER M1 ;
        RECT 4.752 13.656 4.784 16.164 ;
  LAYER M1 ;
        RECT 4.816 13.656 4.848 16.164 ;
  LAYER M1 ;
        RECT 4.88 13.656 4.912 16.164 ;
  LAYER M1 ;
        RECT 4.944 13.656 4.976 16.164 ;
  LAYER M1 ;
        RECT 5.008 13.656 5.04 16.164 ;
  LAYER M1 ;
        RECT 5.072 13.656 5.104 16.164 ;
  LAYER M1 ;
        RECT 5.136 13.656 5.168 16.164 ;
  LAYER M1 ;
        RECT 5.2 13.656 5.232 16.164 ;
  LAYER M1 ;
        RECT 5.264 13.656 5.296 16.164 ;
  LAYER M1 ;
        RECT 5.328 13.656 5.36 16.164 ;
  LAYER M1 ;
        RECT 5.392 13.656 5.424 16.164 ;
  LAYER M1 ;
        RECT 5.456 13.656 5.488 16.164 ;
  LAYER M1 ;
        RECT 5.52 13.656 5.552 16.164 ;
  LAYER M1 ;
        RECT 5.584 13.656 5.616 16.164 ;
  LAYER M1 ;
        RECT 5.648 13.656 5.68 16.164 ;
  LAYER M1 ;
        RECT 5.712 13.656 5.744 16.164 ;
  LAYER M1 ;
        RECT 5.776 13.656 5.808 16.164 ;
  LAYER M1 ;
        RECT 5.84 13.656 5.872 16.164 ;
  LAYER M1 ;
        RECT 5.904 13.656 5.936 16.164 ;
  LAYER M1 ;
        RECT 5.968 13.656 6 16.164 ;
  LAYER M1 ;
        RECT 6.032 13.656 6.064 16.164 ;
  LAYER M1 ;
        RECT 6.096 13.656 6.128 16.164 ;
  LAYER M1 ;
        RECT 6.16 13.656 6.192 16.164 ;
  LAYER M1 ;
        RECT 6.224 13.656 6.256 16.164 ;
  LAYER M1 ;
        RECT 6.288 13.656 6.32 16.164 ;
  LAYER M2 ;
        RECT 3.964 16.048 6.436 16.08 ;
  LAYER M2 ;
        RECT 3.964 15.984 6.436 16.016 ;
  LAYER M2 ;
        RECT 3.964 15.92 6.436 15.952 ;
  LAYER M2 ;
        RECT 3.964 15.856 6.436 15.888 ;
  LAYER M2 ;
        RECT 3.964 15.792 6.436 15.824 ;
  LAYER M2 ;
        RECT 3.964 15.728 6.436 15.76 ;
  LAYER M2 ;
        RECT 3.964 15.664 6.436 15.696 ;
  LAYER M2 ;
        RECT 3.964 15.6 6.436 15.632 ;
  LAYER M2 ;
        RECT 3.964 15.536 6.436 15.568 ;
  LAYER M2 ;
        RECT 3.964 15.472 6.436 15.504 ;
  LAYER M2 ;
        RECT 3.964 15.408 6.436 15.44 ;
  LAYER M2 ;
        RECT 3.964 15.344 6.436 15.376 ;
  LAYER M2 ;
        RECT 3.964 15.28 6.436 15.312 ;
  LAYER M2 ;
        RECT 3.964 15.216 6.436 15.248 ;
  LAYER M2 ;
        RECT 3.964 15.152 6.436 15.184 ;
  LAYER M2 ;
        RECT 3.964 15.088 6.436 15.12 ;
  LAYER M2 ;
        RECT 3.964 15.024 6.436 15.056 ;
  LAYER M2 ;
        RECT 3.964 14.96 6.436 14.992 ;
  LAYER M2 ;
        RECT 3.964 14.896 6.436 14.928 ;
  LAYER M2 ;
        RECT 3.964 14.832 6.436 14.864 ;
  LAYER M2 ;
        RECT 3.964 14.768 6.436 14.8 ;
  LAYER M2 ;
        RECT 3.964 14.704 6.436 14.736 ;
  LAYER M2 ;
        RECT 3.964 14.64 6.436 14.672 ;
  LAYER M2 ;
        RECT 3.964 14.576 6.436 14.608 ;
  LAYER M2 ;
        RECT 3.964 14.512 6.436 14.544 ;
  LAYER M2 ;
        RECT 3.964 14.448 6.436 14.48 ;
  LAYER M2 ;
        RECT 3.964 14.384 6.436 14.416 ;
  LAYER M2 ;
        RECT 3.964 14.32 6.436 14.352 ;
  LAYER M2 ;
        RECT 3.964 14.256 6.436 14.288 ;
  LAYER M2 ;
        RECT 3.964 14.192 6.436 14.224 ;
  LAYER M2 ;
        RECT 3.964 14.128 6.436 14.16 ;
  LAYER M2 ;
        RECT 3.964 14.064 6.436 14.096 ;
  LAYER M2 ;
        RECT 3.964 14 6.436 14.032 ;
  LAYER M2 ;
        RECT 3.964 13.936 6.436 13.968 ;
  LAYER M2 ;
        RECT 3.964 13.872 6.436 13.904 ;
  LAYER M2 ;
        RECT 3.964 13.808 6.436 13.84 ;
  LAYER M3 ;
        RECT 3.984 13.656 4.016 16.164 ;
  LAYER M3 ;
        RECT 4.048 13.656 4.08 16.164 ;
  LAYER M3 ;
        RECT 4.112 13.656 4.144 16.164 ;
  LAYER M3 ;
        RECT 4.176 13.656 4.208 16.164 ;
  LAYER M3 ;
        RECT 4.24 13.656 4.272 16.164 ;
  LAYER M3 ;
        RECT 4.304 13.656 4.336 16.164 ;
  LAYER M3 ;
        RECT 4.368 13.656 4.4 16.164 ;
  LAYER M3 ;
        RECT 4.432 13.656 4.464 16.164 ;
  LAYER M3 ;
        RECT 4.496 13.656 4.528 16.164 ;
  LAYER M3 ;
        RECT 4.56 13.656 4.592 16.164 ;
  LAYER M3 ;
        RECT 4.624 13.656 4.656 16.164 ;
  LAYER M3 ;
        RECT 4.688 13.656 4.72 16.164 ;
  LAYER M3 ;
        RECT 4.752 13.656 4.784 16.164 ;
  LAYER M3 ;
        RECT 4.816 13.656 4.848 16.164 ;
  LAYER M3 ;
        RECT 4.88 13.656 4.912 16.164 ;
  LAYER M3 ;
        RECT 4.944 13.656 4.976 16.164 ;
  LAYER M3 ;
        RECT 5.008 13.656 5.04 16.164 ;
  LAYER M3 ;
        RECT 5.072 13.656 5.104 16.164 ;
  LAYER M3 ;
        RECT 5.136 13.656 5.168 16.164 ;
  LAYER M3 ;
        RECT 5.2 13.656 5.232 16.164 ;
  LAYER M3 ;
        RECT 5.264 13.656 5.296 16.164 ;
  LAYER M3 ;
        RECT 5.328 13.656 5.36 16.164 ;
  LAYER M3 ;
        RECT 5.392 13.656 5.424 16.164 ;
  LAYER M3 ;
        RECT 5.456 13.656 5.488 16.164 ;
  LAYER M3 ;
        RECT 5.52 13.656 5.552 16.164 ;
  LAYER M3 ;
        RECT 5.584 13.656 5.616 16.164 ;
  LAYER M3 ;
        RECT 5.648 13.656 5.68 16.164 ;
  LAYER M3 ;
        RECT 5.712 13.656 5.744 16.164 ;
  LAYER M3 ;
        RECT 5.776 13.656 5.808 16.164 ;
  LAYER M3 ;
        RECT 5.84 13.656 5.872 16.164 ;
  LAYER M3 ;
        RECT 5.904 13.656 5.936 16.164 ;
  LAYER M3 ;
        RECT 5.968 13.656 6 16.164 ;
  LAYER M3 ;
        RECT 6.032 13.656 6.064 16.164 ;
  LAYER M3 ;
        RECT 6.096 13.656 6.128 16.164 ;
  LAYER M3 ;
        RECT 6.16 13.656 6.192 16.164 ;
  LAYER M3 ;
        RECT 6.224 13.656 6.256 16.164 ;
  LAYER M3 ;
        RECT 6.288 13.656 6.32 16.164 ;
  LAYER M3 ;
        RECT 6.384 13.656 6.416 16.164 ;
  LAYER M1 ;
        RECT 3.999 13.692 4.001 16.128 ;
  LAYER M1 ;
        RECT 4.079 13.692 4.081 16.128 ;
  LAYER M1 ;
        RECT 4.159 13.692 4.161 16.128 ;
  LAYER M1 ;
        RECT 4.239 13.692 4.241 16.128 ;
  LAYER M1 ;
        RECT 4.319 13.692 4.321 16.128 ;
  LAYER M1 ;
        RECT 4.399 13.692 4.401 16.128 ;
  LAYER M1 ;
        RECT 4.479 13.692 4.481 16.128 ;
  LAYER M1 ;
        RECT 4.559 13.692 4.561 16.128 ;
  LAYER M1 ;
        RECT 4.639 13.692 4.641 16.128 ;
  LAYER M1 ;
        RECT 4.719 13.692 4.721 16.128 ;
  LAYER M1 ;
        RECT 4.799 13.692 4.801 16.128 ;
  LAYER M1 ;
        RECT 4.879 13.692 4.881 16.128 ;
  LAYER M1 ;
        RECT 4.959 13.692 4.961 16.128 ;
  LAYER M1 ;
        RECT 5.039 13.692 5.041 16.128 ;
  LAYER M1 ;
        RECT 5.119 13.692 5.121 16.128 ;
  LAYER M1 ;
        RECT 5.199 13.692 5.201 16.128 ;
  LAYER M1 ;
        RECT 5.279 13.692 5.281 16.128 ;
  LAYER M1 ;
        RECT 5.359 13.692 5.361 16.128 ;
  LAYER M1 ;
        RECT 5.439 13.692 5.441 16.128 ;
  LAYER M1 ;
        RECT 5.519 13.692 5.521 16.128 ;
  LAYER M1 ;
        RECT 5.599 13.692 5.601 16.128 ;
  LAYER M1 ;
        RECT 5.679 13.692 5.681 16.128 ;
  LAYER M1 ;
        RECT 5.759 13.692 5.761 16.128 ;
  LAYER M1 ;
        RECT 5.839 13.692 5.841 16.128 ;
  LAYER M1 ;
        RECT 5.919 13.692 5.921 16.128 ;
  LAYER M1 ;
        RECT 5.999 13.692 6.001 16.128 ;
  LAYER M1 ;
        RECT 6.079 13.692 6.081 16.128 ;
  LAYER M1 ;
        RECT 6.159 13.692 6.161 16.128 ;
  LAYER M1 ;
        RECT 6.239 13.692 6.241 16.128 ;
  LAYER M1 ;
        RECT 6.319 13.692 6.321 16.128 ;
  LAYER M2 ;
        RECT 4 16.127 6.4 16.129 ;
  LAYER M2 ;
        RECT 4 16.043 6.4 16.045 ;
  LAYER M2 ;
        RECT 4 15.959 6.4 15.961 ;
  LAYER M2 ;
        RECT 4 15.875 6.4 15.877 ;
  LAYER M2 ;
        RECT 4 15.791 6.4 15.793 ;
  LAYER M2 ;
        RECT 4 15.707 6.4 15.709 ;
  LAYER M2 ;
        RECT 4 15.623 6.4 15.625 ;
  LAYER M2 ;
        RECT 4 15.539 6.4 15.541 ;
  LAYER M2 ;
        RECT 4 15.455 6.4 15.457 ;
  LAYER M2 ;
        RECT 4 15.371 6.4 15.373 ;
  LAYER M2 ;
        RECT 4 15.287 6.4 15.289 ;
  LAYER M2 ;
        RECT 4 15.203 6.4 15.205 ;
  LAYER M2 ;
        RECT 4 15.1195 6.4 15.1215 ;
  LAYER M2 ;
        RECT 4 15.035 6.4 15.037 ;
  LAYER M2 ;
        RECT 4 14.951 6.4 14.953 ;
  LAYER M2 ;
        RECT 4 14.867 6.4 14.869 ;
  LAYER M2 ;
        RECT 4 14.783 6.4 14.785 ;
  LAYER M2 ;
        RECT 4 14.699 6.4 14.701 ;
  LAYER M2 ;
        RECT 4 14.615 6.4 14.617 ;
  LAYER M2 ;
        RECT 4 14.531 6.4 14.533 ;
  LAYER M2 ;
        RECT 4 14.447 6.4 14.449 ;
  LAYER M2 ;
        RECT 4 14.363 6.4 14.365 ;
  LAYER M2 ;
        RECT 4 14.279 6.4 14.281 ;
  LAYER M2 ;
        RECT 4 14.195 6.4 14.197 ;
  LAYER M2 ;
        RECT 4 14.111 6.4 14.113 ;
  LAYER M2 ;
        RECT 4 14.027 6.4 14.029 ;
  LAYER M2 ;
        RECT 4 13.943 6.4 13.945 ;
  LAYER M2 ;
        RECT 4 13.859 6.4 13.861 ;
  LAYER M2 ;
        RECT 4 13.775 6.4 13.777 ;
  LAYER M1 ;
        RECT 3.984 10.716 4.016 13.224 ;
  LAYER M1 ;
        RECT 4.048 10.716 4.08 13.224 ;
  LAYER M1 ;
        RECT 4.112 10.716 4.144 13.224 ;
  LAYER M1 ;
        RECT 4.176 10.716 4.208 13.224 ;
  LAYER M1 ;
        RECT 4.24 10.716 4.272 13.224 ;
  LAYER M1 ;
        RECT 4.304 10.716 4.336 13.224 ;
  LAYER M1 ;
        RECT 4.368 10.716 4.4 13.224 ;
  LAYER M1 ;
        RECT 4.432 10.716 4.464 13.224 ;
  LAYER M1 ;
        RECT 4.496 10.716 4.528 13.224 ;
  LAYER M1 ;
        RECT 4.56 10.716 4.592 13.224 ;
  LAYER M1 ;
        RECT 4.624 10.716 4.656 13.224 ;
  LAYER M1 ;
        RECT 4.688 10.716 4.72 13.224 ;
  LAYER M1 ;
        RECT 4.752 10.716 4.784 13.224 ;
  LAYER M1 ;
        RECT 4.816 10.716 4.848 13.224 ;
  LAYER M1 ;
        RECT 4.88 10.716 4.912 13.224 ;
  LAYER M1 ;
        RECT 4.944 10.716 4.976 13.224 ;
  LAYER M1 ;
        RECT 5.008 10.716 5.04 13.224 ;
  LAYER M1 ;
        RECT 5.072 10.716 5.104 13.224 ;
  LAYER M1 ;
        RECT 5.136 10.716 5.168 13.224 ;
  LAYER M1 ;
        RECT 5.2 10.716 5.232 13.224 ;
  LAYER M1 ;
        RECT 5.264 10.716 5.296 13.224 ;
  LAYER M1 ;
        RECT 5.328 10.716 5.36 13.224 ;
  LAYER M1 ;
        RECT 5.392 10.716 5.424 13.224 ;
  LAYER M1 ;
        RECT 5.456 10.716 5.488 13.224 ;
  LAYER M1 ;
        RECT 5.52 10.716 5.552 13.224 ;
  LAYER M1 ;
        RECT 5.584 10.716 5.616 13.224 ;
  LAYER M1 ;
        RECT 5.648 10.716 5.68 13.224 ;
  LAYER M1 ;
        RECT 5.712 10.716 5.744 13.224 ;
  LAYER M1 ;
        RECT 5.776 10.716 5.808 13.224 ;
  LAYER M1 ;
        RECT 5.84 10.716 5.872 13.224 ;
  LAYER M1 ;
        RECT 5.904 10.716 5.936 13.224 ;
  LAYER M1 ;
        RECT 5.968 10.716 6 13.224 ;
  LAYER M1 ;
        RECT 6.032 10.716 6.064 13.224 ;
  LAYER M1 ;
        RECT 6.096 10.716 6.128 13.224 ;
  LAYER M1 ;
        RECT 6.16 10.716 6.192 13.224 ;
  LAYER M1 ;
        RECT 6.224 10.716 6.256 13.224 ;
  LAYER M1 ;
        RECT 6.288 10.716 6.32 13.224 ;
  LAYER M2 ;
        RECT 3.964 13.108 6.436 13.14 ;
  LAYER M2 ;
        RECT 3.964 13.044 6.436 13.076 ;
  LAYER M2 ;
        RECT 3.964 12.98 6.436 13.012 ;
  LAYER M2 ;
        RECT 3.964 12.916 6.436 12.948 ;
  LAYER M2 ;
        RECT 3.964 12.852 6.436 12.884 ;
  LAYER M2 ;
        RECT 3.964 12.788 6.436 12.82 ;
  LAYER M2 ;
        RECT 3.964 12.724 6.436 12.756 ;
  LAYER M2 ;
        RECT 3.964 12.66 6.436 12.692 ;
  LAYER M2 ;
        RECT 3.964 12.596 6.436 12.628 ;
  LAYER M2 ;
        RECT 3.964 12.532 6.436 12.564 ;
  LAYER M2 ;
        RECT 3.964 12.468 6.436 12.5 ;
  LAYER M2 ;
        RECT 3.964 12.404 6.436 12.436 ;
  LAYER M2 ;
        RECT 3.964 12.34 6.436 12.372 ;
  LAYER M2 ;
        RECT 3.964 12.276 6.436 12.308 ;
  LAYER M2 ;
        RECT 3.964 12.212 6.436 12.244 ;
  LAYER M2 ;
        RECT 3.964 12.148 6.436 12.18 ;
  LAYER M2 ;
        RECT 3.964 12.084 6.436 12.116 ;
  LAYER M2 ;
        RECT 3.964 12.02 6.436 12.052 ;
  LAYER M2 ;
        RECT 3.964 11.956 6.436 11.988 ;
  LAYER M2 ;
        RECT 3.964 11.892 6.436 11.924 ;
  LAYER M2 ;
        RECT 3.964 11.828 6.436 11.86 ;
  LAYER M2 ;
        RECT 3.964 11.764 6.436 11.796 ;
  LAYER M2 ;
        RECT 3.964 11.7 6.436 11.732 ;
  LAYER M2 ;
        RECT 3.964 11.636 6.436 11.668 ;
  LAYER M2 ;
        RECT 3.964 11.572 6.436 11.604 ;
  LAYER M2 ;
        RECT 3.964 11.508 6.436 11.54 ;
  LAYER M2 ;
        RECT 3.964 11.444 6.436 11.476 ;
  LAYER M2 ;
        RECT 3.964 11.38 6.436 11.412 ;
  LAYER M2 ;
        RECT 3.964 11.316 6.436 11.348 ;
  LAYER M2 ;
        RECT 3.964 11.252 6.436 11.284 ;
  LAYER M2 ;
        RECT 3.964 11.188 6.436 11.22 ;
  LAYER M2 ;
        RECT 3.964 11.124 6.436 11.156 ;
  LAYER M2 ;
        RECT 3.964 11.06 6.436 11.092 ;
  LAYER M2 ;
        RECT 3.964 10.996 6.436 11.028 ;
  LAYER M2 ;
        RECT 3.964 10.932 6.436 10.964 ;
  LAYER M2 ;
        RECT 3.964 10.868 6.436 10.9 ;
  LAYER M3 ;
        RECT 3.984 10.716 4.016 13.224 ;
  LAYER M3 ;
        RECT 4.048 10.716 4.08 13.224 ;
  LAYER M3 ;
        RECT 4.112 10.716 4.144 13.224 ;
  LAYER M3 ;
        RECT 4.176 10.716 4.208 13.224 ;
  LAYER M3 ;
        RECT 4.24 10.716 4.272 13.224 ;
  LAYER M3 ;
        RECT 4.304 10.716 4.336 13.224 ;
  LAYER M3 ;
        RECT 4.368 10.716 4.4 13.224 ;
  LAYER M3 ;
        RECT 4.432 10.716 4.464 13.224 ;
  LAYER M3 ;
        RECT 4.496 10.716 4.528 13.224 ;
  LAYER M3 ;
        RECT 4.56 10.716 4.592 13.224 ;
  LAYER M3 ;
        RECT 4.624 10.716 4.656 13.224 ;
  LAYER M3 ;
        RECT 4.688 10.716 4.72 13.224 ;
  LAYER M3 ;
        RECT 4.752 10.716 4.784 13.224 ;
  LAYER M3 ;
        RECT 4.816 10.716 4.848 13.224 ;
  LAYER M3 ;
        RECT 4.88 10.716 4.912 13.224 ;
  LAYER M3 ;
        RECT 4.944 10.716 4.976 13.224 ;
  LAYER M3 ;
        RECT 5.008 10.716 5.04 13.224 ;
  LAYER M3 ;
        RECT 5.072 10.716 5.104 13.224 ;
  LAYER M3 ;
        RECT 5.136 10.716 5.168 13.224 ;
  LAYER M3 ;
        RECT 5.2 10.716 5.232 13.224 ;
  LAYER M3 ;
        RECT 5.264 10.716 5.296 13.224 ;
  LAYER M3 ;
        RECT 5.328 10.716 5.36 13.224 ;
  LAYER M3 ;
        RECT 5.392 10.716 5.424 13.224 ;
  LAYER M3 ;
        RECT 5.456 10.716 5.488 13.224 ;
  LAYER M3 ;
        RECT 5.52 10.716 5.552 13.224 ;
  LAYER M3 ;
        RECT 5.584 10.716 5.616 13.224 ;
  LAYER M3 ;
        RECT 5.648 10.716 5.68 13.224 ;
  LAYER M3 ;
        RECT 5.712 10.716 5.744 13.224 ;
  LAYER M3 ;
        RECT 5.776 10.716 5.808 13.224 ;
  LAYER M3 ;
        RECT 5.84 10.716 5.872 13.224 ;
  LAYER M3 ;
        RECT 5.904 10.716 5.936 13.224 ;
  LAYER M3 ;
        RECT 5.968 10.716 6 13.224 ;
  LAYER M3 ;
        RECT 6.032 10.716 6.064 13.224 ;
  LAYER M3 ;
        RECT 6.096 10.716 6.128 13.224 ;
  LAYER M3 ;
        RECT 6.16 10.716 6.192 13.224 ;
  LAYER M3 ;
        RECT 6.224 10.716 6.256 13.224 ;
  LAYER M3 ;
        RECT 6.288 10.716 6.32 13.224 ;
  LAYER M3 ;
        RECT 6.384 10.716 6.416 13.224 ;
  LAYER M1 ;
        RECT 3.999 10.752 4.001 13.188 ;
  LAYER M1 ;
        RECT 4.079 10.752 4.081 13.188 ;
  LAYER M1 ;
        RECT 4.159 10.752 4.161 13.188 ;
  LAYER M1 ;
        RECT 4.239 10.752 4.241 13.188 ;
  LAYER M1 ;
        RECT 4.319 10.752 4.321 13.188 ;
  LAYER M1 ;
        RECT 4.399 10.752 4.401 13.188 ;
  LAYER M1 ;
        RECT 4.479 10.752 4.481 13.188 ;
  LAYER M1 ;
        RECT 4.559 10.752 4.561 13.188 ;
  LAYER M1 ;
        RECT 4.639 10.752 4.641 13.188 ;
  LAYER M1 ;
        RECT 4.719 10.752 4.721 13.188 ;
  LAYER M1 ;
        RECT 4.799 10.752 4.801 13.188 ;
  LAYER M1 ;
        RECT 4.879 10.752 4.881 13.188 ;
  LAYER M1 ;
        RECT 4.959 10.752 4.961 13.188 ;
  LAYER M1 ;
        RECT 5.039 10.752 5.041 13.188 ;
  LAYER M1 ;
        RECT 5.119 10.752 5.121 13.188 ;
  LAYER M1 ;
        RECT 5.199 10.752 5.201 13.188 ;
  LAYER M1 ;
        RECT 5.279 10.752 5.281 13.188 ;
  LAYER M1 ;
        RECT 5.359 10.752 5.361 13.188 ;
  LAYER M1 ;
        RECT 5.439 10.752 5.441 13.188 ;
  LAYER M1 ;
        RECT 5.519 10.752 5.521 13.188 ;
  LAYER M1 ;
        RECT 5.599 10.752 5.601 13.188 ;
  LAYER M1 ;
        RECT 5.679 10.752 5.681 13.188 ;
  LAYER M1 ;
        RECT 5.759 10.752 5.761 13.188 ;
  LAYER M1 ;
        RECT 5.839 10.752 5.841 13.188 ;
  LAYER M1 ;
        RECT 5.919 10.752 5.921 13.188 ;
  LAYER M1 ;
        RECT 5.999 10.752 6.001 13.188 ;
  LAYER M1 ;
        RECT 6.079 10.752 6.081 13.188 ;
  LAYER M1 ;
        RECT 6.159 10.752 6.161 13.188 ;
  LAYER M1 ;
        RECT 6.239 10.752 6.241 13.188 ;
  LAYER M1 ;
        RECT 6.319 10.752 6.321 13.188 ;
  LAYER M2 ;
        RECT 4 13.187 6.4 13.189 ;
  LAYER M2 ;
        RECT 4 13.103 6.4 13.105 ;
  LAYER M2 ;
        RECT 4 13.019 6.4 13.021 ;
  LAYER M2 ;
        RECT 4 12.935 6.4 12.937 ;
  LAYER M2 ;
        RECT 4 12.851 6.4 12.853 ;
  LAYER M2 ;
        RECT 4 12.767 6.4 12.769 ;
  LAYER M2 ;
        RECT 4 12.683 6.4 12.685 ;
  LAYER M2 ;
        RECT 4 12.599 6.4 12.601 ;
  LAYER M2 ;
        RECT 4 12.515 6.4 12.517 ;
  LAYER M2 ;
        RECT 4 12.431 6.4 12.433 ;
  LAYER M2 ;
        RECT 4 12.347 6.4 12.349 ;
  LAYER M2 ;
        RECT 4 12.263 6.4 12.265 ;
  LAYER M2 ;
        RECT 4 12.1795 6.4 12.1815 ;
  LAYER M2 ;
        RECT 4 12.095 6.4 12.097 ;
  LAYER M2 ;
        RECT 4 12.011 6.4 12.013 ;
  LAYER M2 ;
        RECT 4 11.927 6.4 11.929 ;
  LAYER M2 ;
        RECT 4 11.843 6.4 11.845 ;
  LAYER M2 ;
        RECT 4 11.759 6.4 11.761 ;
  LAYER M2 ;
        RECT 4 11.675 6.4 11.677 ;
  LAYER M2 ;
        RECT 4 11.591 6.4 11.593 ;
  LAYER M2 ;
        RECT 4 11.507 6.4 11.509 ;
  LAYER M2 ;
        RECT 4 11.423 6.4 11.425 ;
  LAYER M2 ;
        RECT 4 11.339 6.4 11.341 ;
  LAYER M2 ;
        RECT 4 11.255 6.4 11.257 ;
  LAYER M2 ;
        RECT 4 11.171 6.4 11.173 ;
  LAYER M2 ;
        RECT 4 11.087 6.4 11.089 ;
  LAYER M2 ;
        RECT 4 11.003 6.4 11.005 ;
  LAYER M2 ;
        RECT 4 10.919 6.4 10.921 ;
  LAYER M2 ;
        RECT 4 10.835 6.4 10.837 ;
  LAYER M1 ;
        RECT 3.984 7.776 4.016 10.284 ;
  LAYER M1 ;
        RECT 4.048 7.776 4.08 10.284 ;
  LAYER M1 ;
        RECT 4.112 7.776 4.144 10.284 ;
  LAYER M1 ;
        RECT 4.176 7.776 4.208 10.284 ;
  LAYER M1 ;
        RECT 4.24 7.776 4.272 10.284 ;
  LAYER M1 ;
        RECT 4.304 7.776 4.336 10.284 ;
  LAYER M1 ;
        RECT 4.368 7.776 4.4 10.284 ;
  LAYER M1 ;
        RECT 4.432 7.776 4.464 10.284 ;
  LAYER M1 ;
        RECT 4.496 7.776 4.528 10.284 ;
  LAYER M1 ;
        RECT 4.56 7.776 4.592 10.284 ;
  LAYER M1 ;
        RECT 4.624 7.776 4.656 10.284 ;
  LAYER M1 ;
        RECT 4.688 7.776 4.72 10.284 ;
  LAYER M1 ;
        RECT 4.752 7.776 4.784 10.284 ;
  LAYER M1 ;
        RECT 4.816 7.776 4.848 10.284 ;
  LAYER M1 ;
        RECT 4.88 7.776 4.912 10.284 ;
  LAYER M1 ;
        RECT 4.944 7.776 4.976 10.284 ;
  LAYER M1 ;
        RECT 5.008 7.776 5.04 10.284 ;
  LAYER M1 ;
        RECT 5.072 7.776 5.104 10.284 ;
  LAYER M1 ;
        RECT 5.136 7.776 5.168 10.284 ;
  LAYER M1 ;
        RECT 5.2 7.776 5.232 10.284 ;
  LAYER M1 ;
        RECT 5.264 7.776 5.296 10.284 ;
  LAYER M1 ;
        RECT 5.328 7.776 5.36 10.284 ;
  LAYER M1 ;
        RECT 5.392 7.776 5.424 10.284 ;
  LAYER M1 ;
        RECT 5.456 7.776 5.488 10.284 ;
  LAYER M1 ;
        RECT 5.52 7.776 5.552 10.284 ;
  LAYER M1 ;
        RECT 5.584 7.776 5.616 10.284 ;
  LAYER M1 ;
        RECT 5.648 7.776 5.68 10.284 ;
  LAYER M1 ;
        RECT 5.712 7.776 5.744 10.284 ;
  LAYER M1 ;
        RECT 5.776 7.776 5.808 10.284 ;
  LAYER M1 ;
        RECT 5.84 7.776 5.872 10.284 ;
  LAYER M1 ;
        RECT 5.904 7.776 5.936 10.284 ;
  LAYER M1 ;
        RECT 5.968 7.776 6 10.284 ;
  LAYER M1 ;
        RECT 6.032 7.776 6.064 10.284 ;
  LAYER M1 ;
        RECT 6.096 7.776 6.128 10.284 ;
  LAYER M1 ;
        RECT 6.16 7.776 6.192 10.284 ;
  LAYER M1 ;
        RECT 6.224 7.776 6.256 10.284 ;
  LAYER M1 ;
        RECT 6.288 7.776 6.32 10.284 ;
  LAYER M2 ;
        RECT 3.964 10.168 6.436 10.2 ;
  LAYER M2 ;
        RECT 3.964 10.104 6.436 10.136 ;
  LAYER M2 ;
        RECT 3.964 10.04 6.436 10.072 ;
  LAYER M2 ;
        RECT 3.964 9.976 6.436 10.008 ;
  LAYER M2 ;
        RECT 3.964 9.912 6.436 9.944 ;
  LAYER M2 ;
        RECT 3.964 9.848 6.436 9.88 ;
  LAYER M2 ;
        RECT 3.964 9.784 6.436 9.816 ;
  LAYER M2 ;
        RECT 3.964 9.72 6.436 9.752 ;
  LAYER M2 ;
        RECT 3.964 9.656 6.436 9.688 ;
  LAYER M2 ;
        RECT 3.964 9.592 6.436 9.624 ;
  LAYER M2 ;
        RECT 3.964 9.528 6.436 9.56 ;
  LAYER M2 ;
        RECT 3.964 9.464 6.436 9.496 ;
  LAYER M2 ;
        RECT 3.964 9.4 6.436 9.432 ;
  LAYER M2 ;
        RECT 3.964 9.336 6.436 9.368 ;
  LAYER M2 ;
        RECT 3.964 9.272 6.436 9.304 ;
  LAYER M2 ;
        RECT 3.964 9.208 6.436 9.24 ;
  LAYER M2 ;
        RECT 3.964 9.144 6.436 9.176 ;
  LAYER M2 ;
        RECT 3.964 9.08 6.436 9.112 ;
  LAYER M2 ;
        RECT 3.964 9.016 6.436 9.048 ;
  LAYER M2 ;
        RECT 3.964 8.952 6.436 8.984 ;
  LAYER M2 ;
        RECT 3.964 8.888 6.436 8.92 ;
  LAYER M2 ;
        RECT 3.964 8.824 6.436 8.856 ;
  LAYER M2 ;
        RECT 3.964 8.76 6.436 8.792 ;
  LAYER M2 ;
        RECT 3.964 8.696 6.436 8.728 ;
  LAYER M2 ;
        RECT 3.964 8.632 6.436 8.664 ;
  LAYER M2 ;
        RECT 3.964 8.568 6.436 8.6 ;
  LAYER M2 ;
        RECT 3.964 8.504 6.436 8.536 ;
  LAYER M2 ;
        RECT 3.964 8.44 6.436 8.472 ;
  LAYER M2 ;
        RECT 3.964 8.376 6.436 8.408 ;
  LAYER M2 ;
        RECT 3.964 8.312 6.436 8.344 ;
  LAYER M2 ;
        RECT 3.964 8.248 6.436 8.28 ;
  LAYER M2 ;
        RECT 3.964 8.184 6.436 8.216 ;
  LAYER M2 ;
        RECT 3.964 8.12 6.436 8.152 ;
  LAYER M2 ;
        RECT 3.964 8.056 6.436 8.088 ;
  LAYER M2 ;
        RECT 3.964 7.992 6.436 8.024 ;
  LAYER M2 ;
        RECT 3.964 7.928 6.436 7.96 ;
  LAYER M3 ;
        RECT 3.984 7.776 4.016 10.284 ;
  LAYER M3 ;
        RECT 4.048 7.776 4.08 10.284 ;
  LAYER M3 ;
        RECT 4.112 7.776 4.144 10.284 ;
  LAYER M3 ;
        RECT 4.176 7.776 4.208 10.284 ;
  LAYER M3 ;
        RECT 4.24 7.776 4.272 10.284 ;
  LAYER M3 ;
        RECT 4.304 7.776 4.336 10.284 ;
  LAYER M3 ;
        RECT 4.368 7.776 4.4 10.284 ;
  LAYER M3 ;
        RECT 4.432 7.776 4.464 10.284 ;
  LAYER M3 ;
        RECT 4.496 7.776 4.528 10.284 ;
  LAYER M3 ;
        RECT 4.56 7.776 4.592 10.284 ;
  LAYER M3 ;
        RECT 4.624 7.776 4.656 10.284 ;
  LAYER M3 ;
        RECT 4.688 7.776 4.72 10.284 ;
  LAYER M3 ;
        RECT 4.752 7.776 4.784 10.284 ;
  LAYER M3 ;
        RECT 4.816 7.776 4.848 10.284 ;
  LAYER M3 ;
        RECT 4.88 7.776 4.912 10.284 ;
  LAYER M3 ;
        RECT 4.944 7.776 4.976 10.284 ;
  LAYER M3 ;
        RECT 5.008 7.776 5.04 10.284 ;
  LAYER M3 ;
        RECT 5.072 7.776 5.104 10.284 ;
  LAYER M3 ;
        RECT 5.136 7.776 5.168 10.284 ;
  LAYER M3 ;
        RECT 5.2 7.776 5.232 10.284 ;
  LAYER M3 ;
        RECT 5.264 7.776 5.296 10.284 ;
  LAYER M3 ;
        RECT 5.328 7.776 5.36 10.284 ;
  LAYER M3 ;
        RECT 5.392 7.776 5.424 10.284 ;
  LAYER M3 ;
        RECT 5.456 7.776 5.488 10.284 ;
  LAYER M3 ;
        RECT 5.52 7.776 5.552 10.284 ;
  LAYER M3 ;
        RECT 5.584 7.776 5.616 10.284 ;
  LAYER M3 ;
        RECT 5.648 7.776 5.68 10.284 ;
  LAYER M3 ;
        RECT 5.712 7.776 5.744 10.284 ;
  LAYER M3 ;
        RECT 5.776 7.776 5.808 10.284 ;
  LAYER M3 ;
        RECT 5.84 7.776 5.872 10.284 ;
  LAYER M3 ;
        RECT 5.904 7.776 5.936 10.284 ;
  LAYER M3 ;
        RECT 5.968 7.776 6 10.284 ;
  LAYER M3 ;
        RECT 6.032 7.776 6.064 10.284 ;
  LAYER M3 ;
        RECT 6.096 7.776 6.128 10.284 ;
  LAYER M3 ;
        RECT 6.16 7.776 6.192 10.284 ;
  LAYER M3 ;
        RECT 6.224 7.776 6.256 10.284 ;
  LAYER M3 ;
        RECT 6.288 7.776 6.32 10.284 ;
  LAYER M3 ;
        RECT 6.384 7.776 6.416 10.284 ;
  LAYER M1 ;
        RECT 3.999 7.812 4.001 10.248 ;
  LAYER M1 ;
        RECT 4.079 7.812 4.081 10.248 ;
  LAYER M1 ;
        RECT 4.159 7.812 4.161 10.248 ;
  LAYER M1 ;
        RECT 4.239 7.812 4.241 10.248 ;
  LAYER M1 ;
        RECT 4.319 7.812 4.321 10.248 ;
  LAYER M1 ;
        RECT 4.399 7.812 4.401 10.248 ;
  LAYER M1 ;
        RECT 4.479 7.812 4.481 10.248 ;
  LAYER M1 ;
        RECT 4.559 7.812 4.561 10.248 ;
  LAYER M1 ;
        RECT 4.639 7.812 4.641 10.248 ;
  LAYER M1 ;
        RECT 4.719 7.812 4.721 10.248 ;
  LAYER M1 ;
        RECT 4.799 7.812 4.801 10.248 ;
  LAYER M1 ;
        RECT 4.879 7.812 4.881 10.248 ;
  LAYER M1 ;
        RECT 4.959 7.812 4.961 10.248 ;
  LAYER M1 ;
        RECT 5.039 7.812 5.041 10.248 ;
  LAYER M1 ;
        RECT 5.119 7.812 5.121 10.248 ;
  LAYER M1 ;
        RECT 5.199 7.812 5.201 10.248 ;
  LAYER M1 ;
        RECT 5.279 7.812 5.281 10.248 ;
  LAYER M1 ;
        RECT 5.359 7.812 5.361 10.248 ;
  LAYER M1 ;
        RECT 5.439 7.812 5.441 10.248 ;
  LAYER M1 ;
        RECT 5.519 7.812 5.521 10.248 ;
  LAYER M1 ;
        RECT 5.599 7.812 5.601 10.248 ;
  LAYER M1 ;
        RECT 5.679 7.812 5.681 10.248 ;
  LAYER M1 ;
        RECT 5.759 7.812 5.761 10.248 ;
  LAYER M1 ;
        RECT 5.839 7.812 5.841 10.248 ;
  LAYER M1 ;
        RECT 5.919 7.812 5.921 10.248 ;
  LAYER M1 ;
        RECT 5.999 7.812 6.001 10.248 ;
  LAYER M1 ;
        RECT 6.079 7.812 6.081 10.248 ;
  LAYER M1 ;
        RECT 6.159 7.812 6.161 10.248 ;
  LAYER M1 ;
        RECT 6.239 7.812 6.241 10.248 ;
  LAYER M1 ;
        RECT 6.319 7.812 6.321 10.248 ;
  LAYER M2 ;
        RECT 4 10.247 6.4 10.249 ;
  LAYER M2 ;
        RECT 4 10.163 6.4 10.165 ;
  LAYER M2 ;
        RECT 4 10.079 6.4 10.081 ;
  LAYER M2 ;
        RECT 4 9.995 6.4 9.997 ;
  LAYER M2 ;
        RECT 4 9.911 6.4 9.913 ;
  LAYER M2 ;
        RECT 4 9.827 6.4 9.829 ;
  LAYER M2 ;
        RECT 4 9.743 6.4 9.745 ;
  LAYER M2 ;
        RECT 4 9.659 6.4 9.661 ;
  LAYER M2 ;
        RECT 4 9.575 6.4 9.577 ;
  LAYER M2 ;
        RECT 4 9.491 6.4 9.493 ;
  LAYER M2 ;
        RECT 4 9.407 6.4 9.409 ;
  LAYER M2 ;
        RECT 4 9.323 6.4 9.325 ;
  LAYER M2 ;
        RECT 4 9.2395 6.4 9.2415 ;
  LAYER M2 ;
        RECT 4 9.155 6.4 9.157 ;
  LAYER M2 ;
        RECT 4 9.071 6.4 9.073 ;
  LAYER M2 ;
        RECT 4 8.987 6.4 8.989 ;
  LAYER M2 ;
        RECT 4 8.903 6.4 8.905 ;
  LAYER M2 ;
        RECT 4 8.819 6.4 8.821 ;
  LAYER M2 ;
        RECT 4 8.735 6.4 8.737 ;
  LAYER M2 ;
        RECT 4 8.651 6.4 8.653 ;
  LAYER M2 ;
        RECT 4 8.567 6.4 8.569 ;
  LAYER M2 ;
        RECT 4 8.483 6.4 8.485 ;
  LAYER M2 ;
        RECT 4 8.399 6.4 8.401 ;
  LAYER M2 ;
        RECT 4 8.315 6.4 8.317 ;
  LAYER M2 ;
        RECT 4 8.231 6.4 8.233 ;
  LAYER M2 ;
        RECT 4 8.147 6.4 8.149 ;
  LAYER M2 ;
        RECT 4 8.063 6.4 8.065 ;
  LAYER M2 ;
        RECT 4 7.979 6.4 7.981 ;
  LAYER M2 ;
        RECT 4 7.895 6.4 7.897 ;
  LAYER M1 ;
        RECT 3.984 4.836 4.016 7.344 ;
  LAYER M1 ;
        RECT 4.048 4.836 4.08 7.344 ;
  LAYER M1 ;
        RECT 4.112 4.836 4.144 7.344 ;
  LAYER M1 ;
        RECT 4.176 4.836 4.208 7.344 ;
  LAYER M1 ;
        RECT 4.24 4.836 4.272 7.344 ;
  LAYER M1 ;
        RECT 4.304 4.836 4.336 7.344 ;
  LAYER M1 ;
        RECT 4.368 4.836 4.4 7.344 ;
  LAYER M1 ;
        RECT 4.432 4.836 4.464 7.344 ;
  LAYER M1 ;
        RECT 4.496 4.836 4.528 7.344 ;
  LAYER M1 ;
        RECT 4.56 4.836 4.592 7.344 ;
  LAYER M1 ;
        RECT 4.624 4.836 4.656 7.344 ;
  LAYER M1 ;
        RECT 4.688 4.836 4.72 7.344 ;
  LAYER M1 ;
        RECT 4.752 4.836 4.784 7.344 ;
  LAYER M1 ;
        RECT 4.816 4.836 4.848 7.344 ;
  LAYER M1 ;
        RECT 4.88 4.836 4.912 7.344 ;
  LAYER M1 ;
        RECT 4.944 4.836 4.976 7.344 ;
  LAYER M1 ;
        RECT 5.008 4.836 5.04 7.344 ;
  LAYER M1 ;
        RECT 5.072 4.836 5.104 7.344 ;
  LAYER M1 ;
        RECT 5.136 4.836 5.168 7.344 ;
  LAYER M1 ;
        RECT 5.2 4.836 5.232 7.344 ;
  LAYER M1 ;
        RECT 5.264 4.836 5.296 7.344 ;
  LAYER M1 ;
        RECT 5.328 4.836 5.36 7.344 ;
  LAYER M1 ;
        RECT 5.392 4.836 5.424 7.344 ;
  LAYER M1 ;
        RECT 5.456 4.836 5.488 7.344 ;
  LAYER M1 ;
        RECT 5.52 4.836 5.552 7.344 ;
  LAYER M1 ;
        RECT 5.584 4.836 5.616 7.344 ;
  LAYER M1 ;
        RECT 5.648 4.836 5.68 7.344 ;
  LAYER M1 ;
        RECT 5.712 4.836 5.744 7.344 ;
  LAYER M1 ;
        RECT 5.776 4.836 5.808 7.344 ;
  LAYER M1 ;
        RECT 5.84 4.836 5.872 7.344 ;
  LAYER M1 ;
        RECT 5.904 4.836 5.936 7.344 ;
  LAYER M1 ;
        RECT 5.968 4.836 6 7.344 ;
  LAYER M1 ;
        RECT 6.032 4.836 6.064 7.344 ;
  LAYER M1 ;
        RECT 6.096 4.836 6.128 7.344 ;
  LAYER M1 ;
        RECT 6.16 4.836 6.192 7.344 ;
  LAYER M1 ;
        RECT 6.224 4.836 6.256 7.344 ;
  LAYER M1 ;
        RECT 6.288 4.836 6.32 7.344 ;
  LAYER M2 ;
        RECT 3.964 7.228 6.436 7.26 ;
  LAYER M2 ;
        RECT 3.964 7.164 6.436 7.196 ;
  LAYER M2 ;
        RECT 3.964 7.1 6.436 7.132 ;
  LAYER M2 ;
        RECT 3.964 7.036 6.436 7.068 ;
  LAYER M2 ;
        RECT 3.964 6.972 6.436 7.004 ;
  LAYER M2 ;
        RECT 3.964 6.908 6.436 6.94 ;
  LAYER M2 ;
        RECT 3.964 6.844 6.436 6.876 ;
  LAYER M2 ;
        RECT 3.964 6.78 6.436 6.812 ;
  LAYER M2 ;
        RECT 3.964 6.716 6.436 6.748 ;
  LAYER M2 ;
        RECT 3.964 6.652 6.436 6.684 ;
  LAYER M2 ;
        RECT 3.964 6.588 6.436 6.62 ;
  LAYER M2 ;
        RECT 3.964 6.524 6.436 6.556 ;
  LAYER M2 ;
        RECT 3.964 6.46 6.436 6.492 ;
  LAYER M2 ;
        RECT 3.964 6.396 6.436 6.428 ;
  LAYER M2 ;
        RECT 3.964 6.332 6.436 6.364 ;
  LAYER M2 ;
        RECT 3.964 6.268 6.436 6.3 ;
  LAYER M2 ;
        RECT 3.964 6.204 6.436 6.236 ;
  LAYER M2 ;
        RECT 3.964 6.14 6.436 6.172 ;
  LAYER M2 ;
        RECT 3.964 6.076 6.436 6.108 ;
  LAYER M2 ;
        RECT 3.964 6.012 6.436 6.044 ;
  LAYER M2 ;
        RECT 3.964 5.948 6.436 5.98 ;
  LAYER M2 ;
        RECT 3.964 5.884 6.436 5.916 ;
  LAYER M2 ;
        RECT 3.964 5.82 6.436 5.852 ;
  LAYER M2 ;
        RECT 3.964 5.756 6.436 5.788 ;
  LAYER M2 ;
        RECT 3.964 5.692 6.436 5.724 ;
  LAYER M2 ;
        RECT 3.964 5.628 6.436 5.66 ;
  LAYER M2 ;
        RECT 3.964 5.564 6.436 5.596 ;
  LAYER M2 ;
        RECT 3.964 5.5 6.436 5.532 ;
  LAYER M2 ;
        RECT 3.964 5.436 6.436 5.468 ;
  LAYER M2 ;
        RECT 3.964 5.372 6.436 5.404 ;
  LAYER M2 ;
        RECT 3.964 5.308 6.436 5.34 ;
  LAYER M2 ;
        RECT 3.964 5.244 6.436 5.276 ;
  LAYER M2 ;
        RECT 3.964 5.18 6.436 5.212 ;
  LAYER M2 ;
        RECT 3.964 5.116 6.436 5.148 ;
  LAYER M2 ;
        RECT 3.964 5.052 6.436 5.084 ;
  LAYER M2 ;
        RECT 3.964 4.988 6.436 5.02 ;
  LAYER M3 ;
        RECT 3.984 4.836 4.016 7.344 ;
  LAYER M3 ;
        RECT 4.048 4.836 4.08 7.344 ;
  LAYER M3 ;
        RECT 4.112 4.836 4.144 7.344 ;
  LAYER M3 ;
        RECT 4.176 4.836 4.208 7.344 ;
  LAYER M3 ;
        RECT 4.24 4.836 4.272 7.344 ;
  LAYER M3 ;
        RECT 4.304 4.836 4.336 7.344 ;
  LAYER M3 ;
        RECT 4.368 4.836 4.4 7.344 ;
  LAYER M3 ;
        RECT 4.432 4.836 4.464 7.344 ;
  LAYER M3 ;
        RECT 4.496 4.836 4.528 7.344 ;
  LAYER M3 ;
        RECT 4.56 4.836 4.592 7.344 ;
  LAYER M3 ;
        RECT 4.624 4.836 4.656 7.344 ;
  LAYER M3 ;
        RECT 4.688 4.836 4.72 7.344 ;
  LAYER M3 ;
        RECT 4.752 4.836 4.784 7.344 ;
  LAYER M3 ;
        RECT 4.816 4.836 4.848 7.344 ;
  LAYER M3 ;
        RECT 4.88 4.836 4.912 7.344 ;
  LAYER M3 ;
        RECT 4.944 4.836 4.976 7.344 ;
  LAYER M3 ;
        RECT 5.008 4.836 5.04 7.344 ;
  LAYER M3 ;
        RECT 5.072 4.836 5.104 7.344 ;
  LAYER M3 ;
        RECT 5.136 4.836 5.168 7.344 ;
  LAYER M3 ;
        RECT 5.2 4.836 5.232 7.344 ;
  LAYER M3 ;
        RECT 5.264 4.836 5.296 7.344 ;
  LAYER M3 ;
        RECT 5.328 4.836 5.36 7.344 ;
  LAYER M3 ;
        RECT 5.392 4.836 5.424 7.344 ;
  LAYER M3 ;
        RECT 5.456 4.836 5.488 7.344 ;
  LAYER M3 ;
        RECT 5.52 4.836 5.552 7.344 ;
  LAYER M3 ;
        RECT 5.584 4.836 5.616 7.344 ;
  LAYER M3 ;
        RECT 5.648 4.836 5.68 7.344 ;
  LAYER M3 ;
        RECT 5.712 4.836 5.744 7.344 ;
  LAYER M3 ;
        RECT 5.776 4.836 5.808 7.344 ;
  LAYER M3 ;
        RECT 5.84 4.836 5.872 7.344 ;
  LAYER M3 ;
        RECT 5.904 4.836 5.936 7.344 ;
  LAYER M3 ;
        RECT 5.968 4.836 6 7.344 ;
  LAYER M3 ;
        RECT 6.032 4.836 6.064 7.344 ;
  LAYER M3 ;
        RECT 6.096 4.836 6.128 7.344 ;
  LAYER M3 ;
        RECT 6.16 4.836 6.192 7.344 ;
  LAYER M3 ;
        RECT 6.224 4.836 6.256 7.344 ;
  LAYER M3 ;
        RECT 6.288 4.836 6.32 7.344 ;
  LAYER M3 ;
        RECT 6.384 4.836 6.416 7.344 ;
  LAYER M1 ;
        RECT 3.999 4.872 4.001 7.308 ;
  LAYER M1 ;
        RECT 4.079 4.872 4.081 7.308 ;
  LAYER M1 ;
        RECT 4.159 4.872 4.161 7.308 ;
  LAYER M1 ;
        RECT 4.239 4.872 4.241 7.308 ;
  LAYER M1 ;
        RECT 4.319 4.872 4.321 7.308 ;
  LAYER M1 ;
        RECT 4.399 4.872 4.401 7.308 ;
  LAYER M1 ;
        RECT 4.479 4.872 4.481 7.308 ;
  LAYER M1 ;
        RECT 4.559 4.872 4.561 7.308 ;
  LAYER M1 ;
        RECT 4.639 4.872 4.641 7.308 ;
  LAYER M1 ;
        RECT 4.719 4.872 4.721 7.308 ;
  LAYER M1 ;
        RECT 4.799 4.872 4.801 7.308 ;
  LAYER M1 ;
        RECT 4.879 4.872 4.881 7.308 ;
  LAYER M1 ;
        RECT 4.959 4.872 4.961 7.308 ;
  LAYER M1 ;
        RECT 5.039 4.872 5.041 7.308 ;
  LAYER M1 ;
        RECT 5.119 4.872 5.121 7.308 ;
  LAYER M1 ;
        RECT 5.199 4.872 5.201 7.308 ;
  LAYER M1 ;
        RECT 5.279 4.872 5.281 7.308 ;
  LAYER M1 ;
        RECT 5.359 4.872 5.361 7.308 ;
  LAYER M1 ;
        RECT 5.439 4.872 5.441 7.308 ;
  LAYER M1 ;
        RECT 5.519 4.872 5.521 7.308 ;
  LAYER M1 ;
        RECT 5.599 4.872 5.601 7.308 ;
  LAYER M1 ;
        RECT 5.679 4.872 5.681 7.308 ;
  LAYER M1 ;
        RECT 5.759 4.872 5.761 7.308 ;
  LAYER M1 ;
        RECT 5.839 4.872 5.841 7.308 ;
  LAYER M1 ;
        RECT 5.919 4.872 5.921 7.308 ;
  LAYER M1 ;
        RECT 5.999 4.872 6.001 7.308 ;
  LAYER M1 ;
        RECT 6.079 4.872 6.081 7.308 ;
  LAYER M1 ;
        RECT 6.159 4.872 6.161 7.308 ;
  LAYER M1 ;
        RECT 6.239 4.872 6.241 7.308 ;
  LAYER M1 ;
        RECT 6.319 4.872 6.321 7.308 ;
  LAYER M2 ;
        RECT 4 7.307 6.4 7.309 ;
  LAYER M2 ;
        RECT 4 7.223 6.4 7.225 ;
  LAYER M2 ;
        RECT 4 7.139 6.4 7.141 ;
  LAYER M2 ;
        RECT 4 7.055 6.4 7.057 ;
  LAYER M2 ;
        RECT 4 6.971 6.4 6.973 ;
  LAYER M2 ;
        RECT 4 6.887 6.4 6.889 ;
  LAYER M2 ;
        RECT 4 6.803 6.4 6.805 ;
  LAYER M2 ;
        RECT 4 6.719 6.4 6.721 ;
  LAYER M2 ;
        RECT 4 6.635 6.4 6.637 ;
  LAYER M2 ;
        RECT 4 6.551 6.4 6.553 ;
  LAYER M2 ;
        RECT 4 6.467 6.4 6.469 ;
  LAYER M2 ;
        RECT 4 6.383 6.4 6.385 ;
  LAYER M2 ;
        RECT 4 6.2995 6.4 6.3015 ;
  LAYER M2 ;
        RECT 4 6.215 6.4 6.217 ;
  LAYER M2 ;
        RECT 4 6.131 6.4 6.133 ;
  LAYER M2 ;
        RECT 4 6.047 6.4 6.049 ;
  LAYER M2 ;
        RECT 4 5.963 6.4 5.965 ;
  LAYER M2 ;
        RECT 4 5.879 6.4 5.881 ;
  LAYER M2 ;
        RECT 4 5.795 6.4 5.797 ;
  LAYER M2 ;
        RECT 4 5.711 6.4 5.713 ;
  LAYER M2 ;
        RECT 4 5.627 6.4 5.629 ;
  LAYER M2 ;
        RECT 4 5.543 6.4 5.545 ;
  LAYER M2 ;
        RECT 4 5.459 6.4 5.461 ;
  LAYER M2 ;
        RECT 4 5.375 6.4 5.377 ;
  LAYER M2 ;
        RECT 4 5.291 6.4 5.293 ;
  LAYER M2 ;
        RECT 4 5.207 6.4 5.209 ;
  LAYER M2 ;
        RECT 4 5.123 6.4 5.125 ;
  LAYER M2 ;
        RECT 4 5.039 6.4 5.041 ;
  LAYER M2 ;
        RECT 4 4.955 6.4 4.957 ;
  LAYER M1 ;
        RECT 3.984 1.896 4.016 4.404 ;
  LAYER M1 ;
        RECT 4.048 1.896 4.08 4.404 ;
  LAYER M1 ;
        RECT 4.112 1.896 4.144 4.404 ;
  LAYER M1 ;
        RECT 4.176 1.896 4.208 4.404 ;
  LAYER M1 ;
        RECT 4.24 1.896 4.272 4.404 ;
  LAYER M1 ;
        RECT 4.304 1.896 4.336 4.404 ;
  LAYER M1 ;
        RECT 4.368 1.896 4.4 4.404 ;
  LAYER M1 ;
        RECT 4.432 1.896 4.464 4.404 ;
  LAYER M1 ;
        RECT 4.496 1.896 4.528 4.404 ;
  LAYER M1 ;
        RECT 4.56 1.896 4.592 4.404 ;
  LAYER M1 ;
        RECT 4.624 1.896 4.656 4.404 ;
  LAYER M1 ;
        RECT 4.688 1.896 4.72 4.404 ;
  LAYER M1 ;
        RECT 4.752 1.896 4.784 4.404 ;
  LAYER M1 ;
        RECT 4.816 1.896 4.848 4.404 ;
  LAYER M1 ;
        RECT 4.88 1.896 4.912 4.404 ;
  LAYER M1 ;
        RECT 4.944 1.896 4.976 4.404 ;
  LAYER M1 ;
        RECT 5.008 1.896 5.04 4.404 ;
  LAYER M1 ;
        RECT 5.072 1.896 5.104 4.404 ;
  LAYER M1 ;
        RECT 5.136 1.896 5.168 4.404 ;
  LAYER M1 ;
        RECT 5.2 1.896 5.232 4.404 ;
  LAYER M1 ;
        RECT 5.264 1.896 5.296 4.404 ;
  LAYER M1 ;
        RECT 5.328 1.896 5.36 4.404 ;
  LAYER M1 ;
        RECT 5.392 1.896 5.424 4.404 ;
  LAYER M1 ;
        RECT 5.456 1.896 5.488 4.404 ;
  LAYER M1 ;
        RECT 5.52 1.896 5.552 4.404 ;
  LAYER M1 ;
        RECT 5.584 1.896 5.616 4.404 ;
  LAYER M1 ;
        RECT 5.648 1.896 5.68 4.404 ;
  LAYER M1 ;
        RECT 5.712 1.896 5.744 4.404 ;
  LAYER M1 ;
        RECT 5.776 1.896 5.808 4.404 ;
  LAYER M1 ;
        RECT 5.84 1.896 5.872 4.404 ;
  LAYER M1 ;
        RECT 5.904 1.896 5.936 4.404 ;
  LAYER M1 ;
        RECT 5.968 1.896 6 4.404 ;
  LAYER M1 ;
        RECT 6.032 1.896 6.064 4.404 ;
  LAYER M1 ;
        RECT 6.096 1.896 6.128 4.404 ;
  LAYER M1 ;
        RECT 6.16 1.896 6.192 4.404 ;
  LAYER M1 ;
        RECT 6.224 1.896 6.256 4.404 ;
  LAYER M1 ;
        RECT 6.288 1.896 6.32 4.404 ;
  LAYER M2 ;
        RECT 3.964 4.288 6.436 4.32 ;
  LAYER M2 ;
        RECT 3.964 4.224 6.436 4.256 ;
  LAYER M2 ;
        RECT 3.964 4.16 6.436 4.192 ;
  LAYER M2 ;
        RECT 3.964 4.096 6.436 4.128 ;
  LAYER M2 ;
        RECT 3.964 4.032 6.436 4.064 ;
  LAYER M2 ;
        RECT 3.964 3.968 6.436 4 ;
  LAYER M2 ;
        RECT 3.964 3.904 6.436 3.936 ;
  LAYER M2 ;
        RECT 3.964 3.84 6.436 3.872 ;
  LAYER M2 ;
        RECT 3.964 3.776 6.436 3.808 ;
  LAYER M2 ;
        RECT 3.964 3.712 6.436 3.744 ;
  LAYER M2 ;
        RECT 3.964 3.648 6.436 3.68 ;
  LAYER M2 ;
        RECT 3.964 3.584 6.436 3.616 ;
  LAYER M2 ;
        RECT 3.964 3.52 6.436 3.552 ;
  LAYER M2 ;
        RECT 3.964 3.456 6.436 3.488 ;
  LAYER M2 ;
        RECT 3.964 3.392 6.436 3.424 ;
  LAYER M2 ;
        RECT 3.964 3.328 6.436 3.36 ;
  LAYER M2 ;
        RECT 3.964 3.264 6.436 3.296 ;
  LAYER M2 ;
        RECT 3.964 3.2 6.436 3.232 ;
  LAYER M2 ;
        RECT 3.964 3.136 6.436 3.168 ;
  LAYER M2 ;
        RECT 3.964 3.072 6.436 3.104 ;
  LAYER M2 ;
        RECT 3.964 3.008 6.436 3.04 ;
  LAYER M2 ;
        RECT 3.964 2.944 6.436 2.976 ;
  LAYER M2 ;
        RECT 3.964 2.88 6.436 2.912 ;
  LAYER M2 ;
        RECT 3.964 2.816 6.436 2.848 ;
  LAYER M2 ;
        RECT 3.964 2.752 6.436 2.784 ;
  LAYER M2 ;
        RECT 3.964 2.688 6.436 2.72 ;
  LAYER M2 ;
        RECT 3.964 2.624 6.436 2.656 ;
  LAYER M2 ;
        RECT 3.964 2.56 6.436 2.592 ;
  LAYER M2 ;
        RECT 3.964 2.496 6.436 2.528 ;
  LAYER M2 ;
        RECT 3.964 2.432 6.436 2.464 ;
  LAYER M2 ;
        RECT 3.964 2.368 6.436 2.4 ;
  LAYER M2 ;
        RECT 3.964 2.304 6.436 2.336 ;
  LAYER M2 ;
        RECT 3.964 2.24 6.436 2.272 ;
  LAYER M2 ;
        RECT 3.964 2.176 6.436 2.208 ;
  LAYER M2 ;
        RECT 3.964 2.112 6.436 2.144 ;
  LAYER M2 ;
        RECT 3.964 2.048 6.436 2.08 ;
  LAYER M3 ;
        RECT 3.984 1.896 4.016 4.404 ;
  LAYER M3 ;
        RECT 4.048 1.896 4.08 4.404 ;
  LAYER M3 ;
        RECT 4.112 1.896 4.144 4.404 ;
  LAYER M3 ;
        RECT 4.176 1.896 4.208 4.404 ;
  LAYER M3 ;
        RECT 4.24 1.896 4.272 4.404 ;
  LAYER M3 ;
        RECT 4.304 1.896 4.336 4.404 ;
  LAYER M3 ;
        RECT 4.368 1.896 4.4 4.404 ;
  LAYER M3 ;
        RECT 4.432 1.896 4.464 4.404 ;
  LAYER M3 ;
        RECT 4.496 1.896 4.528 4.404 ;
  LAYER M3 ;
        RECT 4.56 1.896 4.592 4.404 ;
  LAYER M3 ;
        RECT 4.624 1.896 4.656 4.404 ;
  LAYER M3 ;
        RECT 4.688 1.896 4.72 4.404 ;
  LAYER M3 ;
        RECT 4.752 1.896 4.784 4.404 ;
  LAYER M3 ;
        RECT 4.816 1.896 4.848 4.404 ;
  LAYER M3 ;
        RECT 4.88 1.896 4.912 4.404 ;
  LAYER M3 ;
        RECT 4.944 1.896 4.976 4.404 ;
  LAYER M3 ;
        RECT 5.008 1.896 5.04 4.404 ;
  LAYER M3 ;
        RECT 5.072 1.896 5.104 4.404 ;
  LAYER M3 ;
        RECT 5.136 1.896 5.168 4.404 ;
  LAYER M3 ;
        RECT 5.2 1.896 5.232 4.404 ;
  LAYER M3 ;
        RECT 5.264 1.896 5.296 4.404 ;
  LAYER M3 ;
        RECT 5.328 1.896 5.36 4.404 ;
  LAYER M3 ;
        RECT 5.392 1.896 5.424 4.404 ;
  LAYER M3 ;
        RECT 5.456 1.896 5.488 4.404 ;
  LAYER M3 ;
        RECT 5.52 1.896 5.552 4.404 ;
  LAYER M3 ;
        RECT 5.584 1.896 5.616 4.404 ;
  LAYER M3 ;
        RECT 5.648 1.896 5.68 4.404 ;
  LAYER M3 ;
        RECT 5.712 1.896 5.744 4.404 ;
  LAYER M3 ;
        RECT 5.776 1.896 5.808 4.404 ;
  LAYER M3 ;
        RECT 5.84 1.896 5.872 4.404 ;
  LAYER M3 ;
        RECT 5.904 1.896 5.936 4.404 ;
  LAYER M3 ;
        RECT 5.968 1.896 6 4.404 ;
  LAYER M3 ;
        RECT 6.032 1.896 6.064 4.404 ;
  LAYER M3 ;
        RECT 6.096 1.896 6.128 4.404 ;
  LAYER M3 ;
        RECT 6.16 1.896 6.192 4.404 ;
  LAYER M3 ;
        RECT 6.224 1.896 6.256 4.404 ;
  LAYER M3 ;
        RECT 6.288 1.896 6.32 4.404 ;
  LAYER M3 ;
        RECT 6.384 1.896 6.416 4.404 ;
  LAYER M1 ;
        RECT 3.999 1.932 4.001 4.368 ;
  LAYER M1 ;
        RECT 4.079 1.932 4.081 4.368 ;
  LAYER M1 ;
        RECT 4.159 1.932 4.161 4.368 ;
  LAYER M1 ;
        RECT 4.239 1.932 4.241 4.368 ;
  LAYER M1 ;
        RECT 4.319 1.932 4.321 4.368 ;
  LAYER M1 ;
        RECT 4.399 1.932 4.401 4.368 ;
  LAYER M1 ;
        RECT 4.479 1.932 4.481 4.368 ;
  LAYER M1 ;
        RECT 4.559 1.932 4.561 4.368 ;
  LAYER M1 ;
        RECT 4.639 1.932 4.641 4.368 ;
  LAYER M1 ;
        RECT 4.719 1.932 4.721 4.368 ;
  LAYER M1 ;
        RECT 4.799 1.932 4.801 4.368 ;
  LAYER M1 ;
        RECT 4.879 1.932 4.881 4.368 ;
  LAYER M1 ;
        RECT 4.959 1.932 4.961 4.368 ;
  LAYER M1 ;
        RECT 5.039 1.932 5.041 4.368 ;
  LAYER M1 ;
        RECT 5.119 1.932 5.121 4.368 ;
  LAYER M1 ;
        RECT 5.199 1.932 5.201 4.368 ;
  LAYER M1 ;
        RECT 5.279 1.932 5.281 4.368 ;
  LAYER M1 ;
        RECT 5.359 1.932 5.361 4.368 ;
  LAYER M1 ;
        RECT 5.439 1.932 5.441 4.368 ;
  LAYER M1 ;
        RECT 5.519 1.932 5.521 4.368 ;
  LAYER M1 ;
        RECT 5.599 1.932 5.601 4.368 ;
  LAYER M1 ;
        RECT 5.679 1.932 5.681 4.368 ;
  LAYER M1 ;
        RECT 5.759 1.932 5.761 4.368 ;
  LAYER M1 ;
        RECT 5.839 1.932 5.841 4.368 ;
  LAYER M1 ;
        RECT 5.919 1.932 5.921 4.368 ;
  LAYER M1 ;
        RECT 5.999 1.932 6.001 4.368 ;
  LAYER M1 ;
        RECT 6.079 1.932 6.081 4.368 ;
  LAYER M1 ;
        RECT 6.159 1.932 6.161 4.368 ;
  LAYER M1 ;
        RECT 6.239 1.932 6.241 4.368 ;
  LAYER M1 ;
        RECT 6.319 1.932 6.321 4.368 ;
  LAYER M2 ;
        RECT 4 4.367 6.4 4.369 ;
  LAYER M2 ;
        RECT 4 4.283 6.4 4.285 ;
  LAYER M2 ;
        RECT 4 4.199 6.4 4.201 ;
  LAYER M2 ;
        RECT 4 4.115 6.4 4.117 ;
  LAYER M2 ;
        RECT 4 4.031 6.4 4.033 ;
  LAYER M2 ;
        RECT 4 3.947 6.4 3.949 ;
  LAYER M2 ;
        RECT 4 3.863 6.4 3.865 ;
  LAYER M2 ;
        RECT 4 3.779 6.4 3.781 ;
  LAYER M2 ;
        RECT 4 3.695 6.4 3.697 ;
  LAYER M2 ;
        RECT 4 3.611 6.4 3.613 ;
  LAYER M2 ;
        RECT 4 3.527 6.4 3.529 ;
  LAYER M2 ;
        RECT 4 3.443 6.4 3.445 ;
  LAYER M2 ;
        RECT 4 3.3595 6.4 3.3615 ;
  LAYER M2 ;
        RECT 4 3.275 6.4 3.277 ;
  LAYER M2 ;
        RECT 4 3.191 6.4 3.193 ;
  LAYER M2 ;
        RECT 4 3.107 6.4 3.109 ;
  LAYER M2 ;
        RECT 4 3.023 6.4 3.025 ;
  LAYER M2 ;
        RECT 4 2.939 6.4 2.941 ;
  LAYER M2 ;
        RECT 4 2.855 6.4 2.857 ;
  LAYER M2 ;
        RECT 4 2.771 6.4 2.773 ;
  LAYER M2 ;
        RECT 4 2.687 6.4 2.689 ;
  LAYER M2 ;
        RECT 4 2.603 6.4 2.605 ;
  LAYER M2 ;
        RECT 4 2.519 6.4 2.521 ;
  LAYER M2 ;
        RECT 4 2.435 6.4 2.437 ;
  LAYER M2 ;
        RECT 4 2.351 6.4 2.353 ;
  LAYER M2 ;
        RECT 4 2.267 6.4 2.269 ;
  LAYER M2 ;
        RECT 4 2.183 6.4 2.185 ;
  LAYER M2 ;
        RECT 4 2.099 6.4 2.101 ;
  LAYER M2 ;
        RECT 4 2.015 6.4 2.017 ;
  LAYER M1 ;
        RECT 6.864 13.656 6.896 16.164 ;
  LAYER M1 ;
        RECT 6.928 13.656 6.96 16.164 ;
  LAYER M1 ;
        RECT 6.992 13.656 7.024 16.164 ;
  LAYER M1 ;
        RECT 7.056 13.656 7.088 16.164 ;
  LAYER M1 ;
        RECT 7.12 13.656 7.152 16.164 ;
  LAYER M1 ;
        RECT 7.184 13.656 7.216 16.164 ;
  LAYER M1 ;
        RECT 7.248 13.656 7.28 16.164 ;
  LAYER M1 ;
        RECT 7.312 13.656 7.344 16.164 ;
  LAYER M1 ;
        RECT 7.376 13.656 7.408 16.164 ;
  LAYER M1 ;
        RECT 7.44 13.656 7.472 16.164 ;
  LAYER M1 ;
        RECT 7.504 13.656 7.536 16.164 ;
  LAYER M1 ;
        RECT 7.568 13.656 7.6 16.164 ;
  LAYER M1 ;
        RECT 7.632 13.656 7.664 16.164 ;
  LAYER M1 ;
        RECT 7.696 13.656 7.728 16.164 ;
  LAYER M1 ;
        RECT 7.76 13.656 7.792 16.164 ;
  LAYER M1 ;
        RECT 7.824 13.656 7.856 16.164 ;
  LAYER M1 ;
        RECT 7.888 13.656 7.92 16.164 ;
  LAYER M1 ;
        RECT 7.952 13.656 7.984 16.164 ;
  LAYER M1 ;
        RECT 8.016 13.656 8.048 16.164 ;
  LAYER M1 ;
        RECT 8.08 13.656 8.112 16.164 ;
  LAYER M1 ;
        RECT 8.144 13.656 8.176 16.164 ;
  LAYER M1 ;
        RECT 8.208 13.656 8.24 16.164 ;
  LAYER M1 ;
        RECT 8.272 13.656 8.304 16.164 ;
  LAYER M1 ;
        RECT 8.336 13.656 8.368 16.164 ;
  LAYER M1 ;
        RECT 8.4 13.656 8.432 16.164 ;
  LAYER M1 ;
        RECT 8.464 13.656 8.496 16.164 ;
  LAYER M1 ;
        RECT 8.528 13.656 8.56 16.164 ;
  LAYER M1 ;
        RECT 8.592 13.656 8.624 16.164 ;
  LAYER M1 ;
        RECT 8.656 13.656 8.688 16.164 ;
  LAYER M1 ;
        RECT 8.72 13.656 8.752 16.164 ;
  LAYER M1 ;
        RECT 8.784 13.656 8.816 16.164 ;
  LAYER M1 ;
        RECT 8.848 13.656 8.88 16.164 ;
  LAYER M1 ;
        RECT 8.912 13.656 8.944 16.164 ;
  LAYER M1 ;
        RECT 8.976 13.656 9.008 16.164 ;
  LAYER M1 ;
        RECT 9.04 13.656 9.072 16.164 ;
  LAYER M1 ;
        RECT 9.104 13.656 9.136 16.164 ;
  LAYER M1 ;
        RECT 9.168 13.656 9.2 16.164 ;
  LAYER M2 ;
        RECT 6.844 16.048 9.316 16.08 ;
  LAYER M2 ;
        RECT 6.844 15.984 9.316 16.016 ;
  LAYER M2 ;
        RECT 6.844 15.92 9.316 15.952 ;
  LAYER M2 ;
        RECT 6.844 15.856 9.316 15.888 ;
  LAYER M2 ;
        RECT 6.844 15.792 9.316 15.824 ;
  LAYER M2 ;
        RECT 6.844 15.728 9.316 15.76 ;
  LAYER M2 ;
        RECT 6.844 15.664 9.316 15.696 ;
  LAYER M2 ;
        RECT 6.844 15.6 9.316 15.632 ;
  LAYER M2 ;
        RECT 6.844 15.536 9.316 15.568 ;
  LAYER M2 ;
        RECT 6.844 15.472 9.316 15.504 ;
  LAYER M2 ;
        RECT 6.844 15.408 9.316 15.44 ;
  LAYER M2 ;
        RECT 6.844 15.344 9.316 15.376 ;
  LAYER M2 ;
        RECT 6.844 15.28 9.316 15.312 ;
  LAYER M2 ;
        RECT 6.844 15.216 9.316 15.248 ;
  LAYER M2 ;
        RECT 6.844 15.152 9.316 15.184 ;
  LAYER M2 ;
        RECT 6.844 15.088 9.316 15.12 ;
  LAYER M2 ;
        RECT 6.844 15.024 9.316 15.056 ;
  LAYER M2 ;
        RECT 6.844 14.96 9.316 14.992 ;
  LAYER M2 ;
        RECT 6.844 14.896 9.316 14.928 ;
  LAYER M2 ;
        RECT 6.844 14.832 9.316 14.864 ;
  LAYER M2 ;
        RECT 6.844 14.768 9.316 14.8 ;
  LAYER M2 ;
        RECT 6.844 14.704 9.316 14.736 ;
  LAYER M2 ;
        RECT 6.844 14.64 9.316 14.672 ;
  LAYER M2 ;
        RECT 6.844 14.576 9.316 14.608 ;
  LAYER M2 ;
        RECT 6.844 14.512 9.316 14.544 ;
  LAYER M2 ;
        RECT 6.844 14.448 9.316 14.48 ;
  LAYER M2 ;
        RECT 6.844 14.384 9.316 14.416 ;
  LAYER M2 ;
        RECT 6.844 14.32 9.316 14.352 ;
  LAYER M2 ;
        RECT 6.844 14.256 9.316 14.288 ;
  LAYER M2 ;
        RECT 6.844 14.192 9.316 14.224 ;
  LAYER M2 ;
        RECT 6.844 14.128 9.316 14.16 ;
  LAYER M2 ;
        RECT 6.844 14.064 9.316 14.096 ;
  LAYER M2 ;
        RECT 6.844 14 9.316 14.032 ;
  LAYER M2 ;
        RECT 6.844 13.936 9.316 13.968 ;
  LAYER M2 ;
        RECT 6.844 13.872 9.316 13.904 ;
  LAYER M2 ;
        RECT 6.844 13.808 9.316 13.84 ;
  LAYER M3 ;
        RECT 6.864 13.656 6.896 16.164 ;
  LAYER M3 ;
        RECT 6.928 13.656 6.96 16.164 ;
  LAYER M3 ;
        RECT 6.992 13.656 7.024 16.164 ;
  LAYER M3 ;
        RECT 7.056 13.656 7.088 16.164 ;
  LAYER M3 ;
        RECT 7.12 13.656 7.152 16.164 ;
  LAYER M3 ;
        RECT 7.184 13.656 7.216 16.164 ;
  LAYER M3 ;
        RECT 7.248 13.656 7.28 16.164 ;
  LAYER M3 ;
        RECT 7.312 13.656 7.344 16.164 ;
  LAYER M3 ;
        RECT 7.376 13.656 7.408 16.164 ;
  LAYER M3 ;
        RECT 7.44 13.656 7.472 16.164 ;
  LAYER M3 ;
        RECT 7.504 13.656 7.536 16.164 ;
  LAYER M3 ;
        RECT 7.568 13.656 7.6 16.164 ;
  LAYER M3 ;
        RECT 7.632 13.656 7.664 16.164 ;
  LAYER M3 ;
        RECT 7.696 13.656 7.728 16.164 ;
  LAYER M3 ;
        RECT 7.76 13.656 7.792 16.164 ;
  LAYER M3 ;
        RECT 7.824 13.656 7.856 16.164 ;
  LAYER M3 ;
        RECT 7.888 13.656 7.92 16.164 ;
  LAYER M3 ;
        RECT 7.952 13.656 7.984 16.164 ;
  LAYER M3 ;
        RECT 8.016 13.656 8.048 16.164 ;
  LAYER M3 ;
        RECT 8.08 13.656 8.112 16.164 ;
  LAYER M3 ;
        RECT 8.144 13.656 8.176 16.164 ;
  LAYER M3 ;
        RECT 8.208 13.656 8.24 16.164 ;
  LAYER M3 ;
        RECT 8.272 13.656 8.304 16.164 ;
  LAYER M3 ;
        RECT 8.336 13.656 8.368 16.164 ;
  LAYER M3 ;
        RECT 8.4 13.656 8.432 16.164 ;
  LAYER M3 ;
        RECT 8.464 13.656 8.496 16.164 ;
  LAYER M3 ;
        RECT 8.528 13.656 8.56 16.164 ;
  LAYER M3 ;
        RECT 8.592 13.656 8.624 16.164 ;
  LAYER M3 ;
        RECT 8.656 13.656 8.688 16.164 ;
  LAYER M3 ;
        RECT 8.72 13.656 8.752 16.164 ;
  LAYER M3 ;
        RECT 8.784 13.656 8.816 16.164 ;
  LAYER M3 ;
        RECT 8.848 13.656 8.88 16.164 ;
  LAYER M3 ;
        RECT 8.912 13.656 8.944 16.164 ;
  LAYER M3 ;
        RECT 8.976 13.656 9.008 16.164 ;
  LAYER M3 ;
        RECT 9.04 13.656 9.072 16.164 ;
  LAYER M3 ;
        RECT 9.104 13.656 9.136 16.164 ;
  LAYER M3 ;
        RECT 9.168 13.656 9.2 16.164 ;
  LAYER M3 ;
        RECT 9.264 13.656 9.296 16.164 ;
  LAYER M1 ;
        RECT 6.879 13.692 6.881 16.128 ;
  LAYER M1 ;
        RECT 6.959 13.692 6.961 16.128 ;
  LAYER M1 ;
        RECT 7.039 13.692 7.041 16.128 ;
  LAYER M1 ;
        RECT 7.119 13.692 7.121 16.128 ;
  LAYER M1 ;
        RECT 7.199 13.692 7.201 16.128 ;
  LAYER M1 ;
        RECT 7.279 13.692 7.281 16.128 ;
  LAYER M1 ;
        RECT 7.359 13.692 7.361 16.128 ;
  LAYER M1 ;
        RECT 7.439 13.692 7.441 16.128 ;
  LAYER M1 ;
        RECT 7.519 13.692 7.521 16.128 ;
  LAYER M1 ;
        RECT 7.599 13.692 7.601 16.128 ;
  LAYER M1 ;
        RECT 7.679 13.692 7.681 16.128 ;
  LAYER M1 ;
        RECT 7.759 13.692 7.761 16.128 ;
  LAYER M1 ;
        RECT 7.839 13.692 7.841 16.128 ;
  LAYER M1 ;
        RECT 7.919 13.692 7.921 16.128 ;
  LAYER M1 ;
        RECT 7.999 13.692 8.001 16.128 ;
  LAYER M1 ;
        RECT 8.079 13.692 8.081 16.128 ;
  LAYER M1 ;
        RECT 8.159 13.692 8.161 16.128 ;
  LAYER M1 ;
        RECT 8.239 13.692 8.241 16.128 ;
  LAYER M1 ;
        RECT 8.319 13.692 8.321 16.128 ;
  LAYER M1 ;
        RECT 8.399 13.692 8.401 16.128 ;
  LAYER M1 ;
        RECT 8.479 13.692 8.481 16.128 ;
  LAYER M1 ;
        RECT 8.559 13.692 8.561 16.128 ;
  LAYER M1 ;
        RECT 8.639 13.692 8.641 16.128 ;
  LAYER M1 ;
        RECT 8.719 13.692 8.721 16.128 ;
  LAYER M1 ;
        RECT 8.799 13.692 8.801 16.128 ;
  LAYER M1 ;
        RECT 8.879 13.692 8.881 16.128 ;
  LAYER M1 ;
        RECT 8.959 13.692 8.961 16.128 ;
  LAYER M1 ;
        RECT 9.039 13.692 9.041 16.128 ;
  LAYER M1 ;
        RECT 9.119 13.692 9.121 16.128 ;
  LAYER M1 ;
        RECT 9.199 13.692 9.201 16.128 ;
  LAYER M2 ;
        RECT 6.88 16.127 9.28 16.129 ;
  LAYER M2 ;
        RECT 6.88 16.043 9.28 16.045 ;
  LAYER M2 ;
        RECT 6.88 15.959 9.28 15.961 ;
  LAYER M2 ;
        RECT 6.88 15.875 9.28 15.877 ;
  LAYER M2 ;
        RECT 6.88 15.791 9.28 15.793 ;
  LAYER M2 ;
        RECT 6.88 15.707 9.28 15.709 ;
  LAYER M2 ;
        RECT 6.88 15.623 9.28 15.625 ;
  LAYER M2 ;
        RECT 6.88 15.539 9.28 15.541 ;
  LAYER M2 ;
        RECT 6.88 15.455 9.28 15.457 ;
  LAYER M2 ;
        RECT 6.88 15.371 9.28 15.373 ;
  LAYER M2 ;
        RECT 6.88 15.287 9.28 15.289 ;
  LAYER M2 ;
        RECT 6.88 15.203 9.28 15.205 ;
  LAYER M2 ;
        RECT 6.88 15.1195 9.28 15.1215 ;
  LAYER M2 ;
        RECT 6.88 15.035 9.28 15.037 ;
  LAYER M2 ;
        RECT 6.88 14.951 9.28 14.953 ;
  LAYER M2 ;
        RECT 6.88 14.867 9.28 14.869 ;
  LAYER M2 ;
        RECT 6.88 14.783 9.28 14.785 ;
  LAYER M2 ;
        RECT 6.88 14.699 9.28 14.701 ;
  LAYER M2 ;
        RECT 6.88 14.615 9.28 14.617 ;
  LAYER M2 ;
        RECT 6.88 14.531 9.28 14.533 ;
  LAYER M2 ;
        RECT 6.88 14.447 9.28 14.449 ;
  LAYER M2 ;
        RECT 6.88 14.363 9.28 14.365 ;
  LAYER M2 ;
        RECT 6.88 14.279 9.28 14.281 ;
  LAYER M2 ;
        RECT 6.88 14.195 9.28 14.197 ;
  LAYER M2 ;
        RECT 6.88 14.111 9.28 14.113 ;
  LAYER M2 ;
        RECT 6.88 14.027 9.28 14.029 ;
  LAYER M2 ;
        RECT 6.88 13.943 9.28 13.945 ;
  LAYER M2 ;
        RECT 6.88 13.859 9.28 13.861 ;
  LAYER M2 ;
        RECT 6.88 13.775 9.28 13.777 ;
  LAYER M1 ;
        RECT 6.864 10.716 6.896 13.224 ;
  LAYER M1 ;
        RECT 6.928 10.716 6.96 13.224 ;
  LAYER M1 ;
        RECT 6.992 10.716 7.024 13.224 ;
  LAYER M1 ;
        RECT 7.056 10.716 7.088 13.224 ;
  LAYER M1 ;
        RECT 7.12 10.716 7.152 13.224 ;
  LAYER M1 ;
        RECT 7.184 10.716 7.216 13.224 ;
  LAYER M1 ;
        RECT 7.248 10.716 7.28 13.224 ;
  LAYER M1 ;
        RECT 7.312 10.716 7.344 13.224 ;
  LAYER M1 ;
        RECT 7.376 10.716 7.408 13.224 ;
  LAYER M1 ;
        RECT 7.44 10.716 7.472 13.224 ;
  LAYER M1 ;
        RECT 7.504 10.716 7.536 13.224 ;
  LAYER M1 ;
        RECT 7.568 10.716 7.6 13.224 ;
  LAYER M1 ;
        RECT 7.632 10.716 7.664 13.224 ;
  LAYER M1 ;
        RECT 7.696 10.716 7.728 13.224 ;
  LAYER M1 ;
        RECT 7.76 10.716 7.792 13.224 ;
  LAYER M1 ;
        RECT 7.824 10.716 7.856 13.224 ;
  LAYER M1 ;
        RECT 7.888 10.716 7.92 13.224 ;
  LAYER M1 ;
        RECT 7.952 10.716 7.984 13.224 ;
  LAYER M1 ;
        RECT 8.016 10.716 8.048 13.224 ;
  LAYER M1 ;
        RECT 8.08 10.716 8.112 13.224 ;
  LAYER M1 ;
        RECT 8.144 10.716 8.176 13.224 ;
  LAYER M1 ;
        RECT 8.208 10.716 8.24 13.224 ;
  LAYER M1 ;
        RECT 8.272 10.716 8.304 13.224 ;
  LAYER M1 ;
        RECT 8.336 10.716 8.368 13.224 ;
  LAYER M1 ;
        RECT 8.4 10.716 8.432 13.224 ;
  LAYER M1 ;
        RECT 8.464 10.716 8.496 13.224 ;
  LAYER M1 ;
        RECT 8.528 10.716 8.56 13.224 ;
  LAYER M1 ;
        RECT 8.592 10.716 8.624 13.224 ;
  LAYER M1 ;
        RECT 8.656 10.716 8.688 13.224 ;
  LAYER M1 ;
        RECT 8.72 10.716 8.752 13.224 ;
  LAYER M1 ;
        RECT 8.784 10.716 8.816 13.224 ;
  LAYER M1 ;
        RECT 8.848 10.716 8.88 13.224 ;
  LAYER M1 ;
        RECT 8.912 10.716 8.944 13.224 ;
  LAYER M1 ;
        RECT 8.976 10.716 9.008 13.224 ;
  LAYER M1 ;
        RECT 9.04 10.716 9.072 13.224 ;
  LAYER M1 ;
        RECT 9.104 10.716 9.136 13.224 ;
  LAYER M1 ;
        RECT 9.168 10.716 9.2 13.224 ;
  LAYER M2 ;
        RECT 6.844 13.108 9.316 13.14 ;
  LAYER M2 ;
        RECT 6.844 13.044 9.316 13.076 ;
  LAYER M2 ;
        RECT 6.844 12.98 9.316 13.012 ;
  LAYER M2 ;
        RECT 6.844 12.916 9.316 12.948 ;
  LAYER M2 ;
        RECT 6.844 12.852 9.316 12.884 ;
  LAYER M2 ;
        RECT 6.844 12.788 9.316 12.82 ;
  LAYER M2 ;
        RECT 6.844 12.724 9.316 12.756 ;
  LAYER M2 ;
        RECT 6.844 12.66 9.316 12.692 ;
  LAYER M2 ;
        RECT 6.844 12.596 9.316 12.628 ;
  LAYER M2 ;
        RECT 6.844 12.532 9.316 12.564 ;
  LAYER M2 ;
        RECT 6.844 12.468 9.316 12.5 ;
  LAYER M2 ;
        RECT 6.844 12.404 9.316 12.436 ;
  LAYER M2 ;
        RECT 6.844 12.34 9.316 12.372 ;
  LAYER M2 ;
        RECT 6.844 12.276 9.316 12.308 ;
  LAYER M2 ;
        RECT 6.844 12.212 9.316 12.244 ;
  LAYER M2 ;
        RECT 6.844 12.148 9.316 12.18 ;
  LAYER M2 ;
        RECT 6.844 12.084 9.316 12.116 ;
  LAYER M2 ;
        RECT 6.844 12.02 9.316 12.052 ;
  LAYER M2 ;
        RECT 6.844 11.956 9.316 11.988 ;
  LAYER M2 ;
        RECT 6.844 11.892 9.316 11.924 ;
  LAYER M2 ;
        RECT 6.844 11.828 9.316 11.86 ;
  LAYER M2 ;
        RECT 6.844 11.764 9.316 11.796 ;
  LAYER M2 ;
        RECT 6.844 11.7 9.316 11.732 ;
  LAYER M2 ;
        RECT 6.844 11.636 9.316 11.668 ;
  LAYER M2 ;
        RECT 6.844 11.572 9.316 11.604 ;
  LAYER M2 ;
        RECT 6.844 11.508 9.316 11.54 ;
  LAYER M2 ;
        RECT 6.844 11.444 9.316 11.476 ;
  LAYER M2 ;
        RECT 6.844 11.38 9.316 11.412 ;
  LAYER M2 ;
        RECT 6.844 11.316 9.316 11.348 ;
  LAYER M2 ;
        RECT 6.844 11.252 9.316 11.284 ;
  LAYER M2 ;
        RECT 6.844 11.188 9.316 11.22 ;
  LAYER M2 ;
        RECT 6.844 11.124 9.316 11.156 ;
  LAYER M2 ;
        RECT 6.844 11.06 9.316 11.092 ;
  LAYER M2 ;
        RECT 6.844 10.996 9.316 11.028 ;
  LAYER M2 ;
        RECT 6.844 10.932 9.316 10.964 ;
  LAYER M2 ;
        RECT 6.844 10.868 9.316 10.9 ;
  LAYER M3 ;
        RECT 6.864 10.716 6.896 13.224 ;
  LAYER M3 ;
        RECT 6.928 10.716 6.96 13.224 ;
  LAYER M3 ;
        RECT 6.992 10.716 7.024 13.224 ;
  LAYER M3 ;
        RECT 7.056 10.716 7.088 13.224 ;
  LAYER M3 ;
        RECT 7.12 10.716 7.152 13.224 ;
  LAYER M3 ;
        RECT 7.184 10.716 7.216 13.224 ;
  LAYER M3 ;
        RECT 7.248 10.716 7.28 13.224 ;
  LAYER M3 ;
        RECT 7.312 10.716 7.344 13.224 ;
  LAYER M3 ;
        RECT 7.376 10.716 7.408 13.224 ;
  LAYER M3 ;
        RECT 7.44 10.716 7.472 13.224 ;
  LAYER M3 ;
        RECT 7.504 10.716 7.536 13.224 ;
  LAYER M3 ;
        RECT 7.568 10.716 7.6 13.224 ;
  LAYER M3 ;
        RECT 7.632 10.716 7.664 13.224 ;
  LAYER M3 ;
        RECT 7.696 10.716 7.728 13.224 ;
  LAYER M3 ;
        RECT 7.76 10.716 7.792 13.224 ;
  LAYER M3 ;
        RECT 7.824 10.716 7.856 13.224 ;
  LAYER M3 ;
        RECT 7.888 10.716 7.92 13.224 ;
  LAYER M3 ;
        RECT 7.952 10.716 7.984 13.224 ;
  LAYER M3 ;
        RECT 8.016 10.716 8.048 13.224 ;
  LAYER M3 ;
        RECT 8.08 10.716 8.112 13.224 ;
  LAYER M3 ;
        RECT 8.144 10.716 8.176 13.224 ;
  LAYER M3 ;
        RECT 8.208 10.716 8.24 13.224 ;
  LAYER M3 ;
        RECT 8.272 10.716 8.304 13.224 ;
  LAYER M3 ;
        RECT 8.336 10.716 8.368 13.224 ;
  LAYER M3 ;
        RECT 8.4 10.716 8.432 13.224 ;
  LAYER M3 ;
        RECT 8.464 10.716 8.496 13.224 ;
  LAYER M3 ;
        RECT 8.528 10.716 8.56 13.224 ;
  LAYER M3 ;
        RECT 8.592 10.716 8.624 13.224 ;
  LAYER M3 ;
        RECT 8.656 10.716 8.688 13.224 ;
  LAYER M3 ;
        RECT 8.72 10.716 8.752 13.224 ;
  LAYER M3 ;
        RECT 8.784 10.716 8.816 13.224 ;
  LAYER M3 ;
        RECT 8.848 10.716 8.88 13.224 ;
  LAYER M3 ;
        RECT 8.912 10.716 8.944 13.224 ;
  LAYER M3 ;
        RECT 8.976 10.716 9.008 13.224 ;
  LAYER M3 ;
        RECT 9.04 10.716 9.072 13.224 ;
  LAYER M3 ;
        RECT 9.104 10.716 9.136 13.224 ;
  LAYER M3 ;
        RECT 9.168 10.716 9.2 13.224 ;
  LAYER M3 ;
        RECT 9.264 10.716 9.296 13.224 ;
  LAYER M1 ;
        RECT 6.879 10.752 6.881 13.188 ;
  LAYER M1 ;
        RECT 6.959 10.752 6.961 13.188 ;
  LAYER M1 ;
        RECT 7.039 10.752 7.041 13.188 ;
  LAYER M1 ;
        RECT 7.119 10.752 7.121 13.188 ;
  LAYER M1 ;
        RECT 7.199 10.752 7.201 13.188 ;
  LAYER M1 ;
        RECT 7.279 10.752 7.281 13.188 ;
  LAYER M1 ;
        RECT 7.359 10.752 7.361 13.188 ;
  LAYER M1 ;
        RECT 7.439 10.752 7.441 13.188 ;
  LAYER M1 ;
        RECT 7.519 10.752 7.521 13.188 ;
  LAYER M1 ;
        RECT 7.599 10.752 7.601 13.188 ;
  LAYER M1 ;
        RECT 7.679 10.752 7.681 13.188 ;
  LAYER M1 ;
        RECT 7.759 10.752 7.761 13.188 ;
  LAYER M1 ;
        RECT 7.839 10.752 7.841 13.188 ;
  LAYER M1 ;
        RECT 7.919 10.752 7.921 13.188 ;
  LAYER M1 ;
        RECT 7.999 10.752 8.001 13.188 ;
  LAYER M1 ;
        RECT 8.079 10.752 8.081 13.188 ;
  LAYER M1 ;
        RECT 8.159 10.752 8.161 13.188 ;
  LAYER M1 ;
        RECT 8.239 10.752 8.241 13.188 ;
  LAYER M1 ;
        RECT 8.319 10.752 8.321 13.188 ;
  LAYER M1 ;
        RECT 8.399 10.752 8.401 13.188 ;
  LAYER M1 ;
        RECT 8.479 10.752 8.481 13.188 ;
  LAYER M1 ;
        RECT 8.559 10.752 8.561 13.188 ;
  LAYER M1 ;
        RECT 8.639 10.752 8.641 13.188 ;
  LAYER M1 ;
        RECT 8.719 10.752 8.721 13.188 ;
  LAYER M1 ;
        RECT 8.799 10.752 8.801 13.188 ;
  LAYER M1 ;
        RECT 8.879 10.752 8.881 13.188 ;
  LAYER M1 ;
        RECT 8.959 10.752 8.961 13.188 ;
  LAYER M1 ;
        RECT 9.039 10.752 9.041 13.188 ;
  LAYER M1 ;
        RECT 9.119 10.752 9.121 13.188 ;
  LAYER M1 ;
        RECT 9.199 10.752 9.201 13.188 ;
  LAYER M2 ;
        RECT 6.88 13.187 9.28 13.189 ;
  LAYER M2 ;
        RECT 6.88 13.103 9.28 13.105 ;
  LAYER M2 ;
        RECT 6.88 13.019 9.28 13.021 ;
  LAYER M2 ;
        RECT 6.88 12.935 9.28 12.937 ;
  LAYER M2 ;
        RECT 6.88 12.851 9.28 12.853 ;
  LAYER M2 ;
        RECT 6.88 12.767 9.28 12.769 ;
  LAYER M2 ;
        RECT 6.88 12.683 9.28 12.685 ;
  LAYER M2 ;
        RECT 6.88 12.599 9.28 12.601 ;
  LAYER M2 ;
        RECT 6.88 12.515 9.28 12.517 ;
  LAYER M2 ;
        RECT 6.88 12.431 9.28 12.433 ;
  LAYER M2 ;
        RECT 6.88 12.347 9.28 12.349 ;
  LAYER M2 ;
        RECT 6.88 12.263 9.28 12.265 ;
  LAYER M2 ;
        RECT 6.88 12.1795 9.28 12.1815 ;
  LAYER M2 ;
        RECT 6.88 12.095 9.28 12.097 ;
  LAYER M2 ;
        RECT 6.88 12.011 9.28 12.013 ;
  LAYER M2 ;
        RECT 6.88 11.927 9.28 11.929 ;
  LAYER M2 ;
        RECT 6.88 11.843 9.28 11.845 ;
  LAYER M2 ;
        RECT 6.88 11.759 9.28 11.761 ;
  LAYER M2 ;
        RECT 6.88 11.675 9.28 11.677 ;
  LAYER M2 ;
        RECT 6.88 11.591 9.28 11.593 ;
  LAYER M2 ;
        RECT 6.88 11.507 9.28 11.509 ;
  LAYER M2 ;
        RECT 6.88 11.423 9.28 11.425 ;
  LAYER M2 ;
        RECT 6.88 11.339 9.28 11.341 ;
  LAYER M2 ;
        RECT 6.88 11.255 9.28 11.257 ;
  LAYER M2 ;
        RECT 6.88 11.171 9.28 11.173 ;
  LAYER M2 ;
        RECT 6.88 11.087 9.28 11.089 ;
  LAYER M2 ;
        RECT 6.88 11.003 9.28 11.005 ;
  LAYER M2 ;
        RECT 6.88 10.919 9.28 10.921 ;
  LAYER M2 ;
        RECT 6.88 10.835 9.28 10.837 ;
  LAYER M1 ;
        RECT 6.864 7.776 6.896 10.284 ;
  LAYER M1 ;
        RECT 6.928 7.776 6.96 10.284 ;
  LAYER M1 ;
        RECT 6.992 7.776 7.024 10.284 ;
  LAYER M1 ;
        RECT 7.056 7.776 7.088 10.284 ;
  LAYER M1 ;
        RECT 7.12 7.776 7.152 10.284 ;
  LAYER M1 ;
        RECT 7.184 7.776 7.216 10.284 ;
  LAYER M1 ;
        RECT 7.248 7.776 7.28 10.284 ;
  LAYER M1 ;
        RECT 7.312 7.776 7.344 10.284 ;
  LAYER M1 ;
        RECT 7.376 7.776 7.408 10.284 ;
  LAYER M1 ;
        RECT 7.44 7.776 7.472 10.284 ;
  LAYER M1 ;
        RECT 7.504 7.776 7.536 10.284 ;
  LAYER M1 ;
        RECT 7.568 7.776 7.6 10.284 ;
  LAYER M1 ;
        RECT 7.632 7.776 7.664 10.284 ;
  LAYER M1 ;
        RECT 7.696 7.776 7.728 10.284 ;
  LAYER M1 ;
        RECT 7.76 7.776 7.792 10.284 ;
  LAYER M1 ;
        RECT 7.824 7.776 7.856 10.284 ;
  LAYER M1 ;
        RECT 7.888 7.776 7.92 10.284 ;
  LAYER M1 ;
        RECT 7.952 7.776 7.984 10.284 ;
  LAYER M1 ;
        RECT 8.016 7.776 8.048 10.284 ;
  LAYER M1 ;
        RECT 8.08 7.776 8.112 10.284 ;
  LAYER M1 ;
        RECT 8.144 7.776 8.176 10.284 ;
  LAYER M1 ;
        RECT 8.208 7.776 8.24 10.284 ;
  LAYER M1 ;
        RECT 8.272 7.776 8.304 10.284 ;
  LAYER M1 ;
        RECT 8.336 7.776 8.368 10.284 ;
  LAYER M1 ;
        RECT 8.4 7.776 8.432 10.284 ;
  LAYER M1 ;
        RECT 8.464 7.776 8.496 10.284 ;
  LAYER M1 ;
        RECT 8.528 7.776 8.56 10.284 ;
  LAYER M1 ;
        RECT 8.592 7.776 8.624 10.284 ;
  LAYER M1 ;
        RECT 8.656 7.776 8.688 10.284 ;
  LAYER M1 ;
        RECT 8.72 7.776 8.752 10.284 ;
  LAYER M1 ;
        RECT 8.784 7.776 8.816 10.284 ;
  LAYER M1 ;
        RECT 8.848 7.776 8.88 10.284 ;
  LAYER M1 ;
        RECT 8.912 7.776 8.944 10.284 ;
  LAYER M1 ;
        RECT 8.976 7.776 9.008 10.284 ;
  LAYER M1 ;
        RECT 9.04 7.776 9.072 10.284 ;
  LAYER M1 ;
        RECT 9.104 7.776 9.136 10.284 ;
  LAYER M1 ;
        RECT 9.168 7.776 9.2 10.284 ;
  LAYER M2 ;
        RECT 6.844 10.168 9.316 10.2 ;
  LAYER M2 ;
        RECT 6.844 10.104 9.316 10.136 ;
  LAYER M2 ;
        RECT 6.844 10.04 9.316 10.072 ;
  LAYER M2 ;
        RECT 6.844 9.976 9.316 10.008 ;
  LAYER M2 ;
        RECT 6.844 9.912 9.316 9.944 ;
  LAYER M2 ;
        RECT 6.844 9.848 9.316 9.88 ;
  LAYER M2 ;
        RECT 6.844 9.784 9.316 9.816 ;
  LAYER M2 ;
        RECT 6.844 9.72 9.316 9.752 ;
  LAYER M2 ;
        RECT 6.844 9.656 9.316 9.688 ;
  LAYER M2 ;
        RECT 6.844 9.592 9.316 9.624 ;
  LAYER M2 ;
        RECT 6.844 9.528 9.316 9.56 ;
  LAYER M2 ;
        RECT 6.844 9.464 9.316 9.496 ;
  LAYER M2 ;
        RECT 6.844 9.4 9.316 9.432 ;
  LAYER M2 ;
        RECT 6.844 9.336 9.316 9.368 ;
  LAYER M2 ;
        RECT 6.844 9.272 9.316 9.304 ;
  LAYER M2 ;
        RECT 6.844 9.208 9.316 9.24 ;
  LAYER M2 ;
        RECT 6.844 9.144 9.316 9.176 ;
  LAYER M2 ;
        RECT 6.844 9.08 9.316 9.112 ;
  LAYER M2 ;
        RECT 6.844 9.016 9.316 9.048 ;
  LAYER M2 ;
        RECT 6.844 8.952 9.316 8.984 ;
  LAYER M2 ;
        RECT 6.844 8.888 9.316 8.92 ;
  LAYER M2 ;
        RECT 6.844 8.824 9.316 8.856 ;
  LAYER M2 ;
        RECT 6.844 8.76 9.316 8.792 ;
  LAYER M2 ;
        RECT 6.844 8.696 9.316 8.728 ;
  LAYER M2 ;
        RECT 6.844 8.632 9.316 8.664 ;
  LAYER M2 ;
        RECT 6.844 8.568 9.316 8.6 ;
  LAYER M2 ;
        RECT 6.844 8.504 9.316 8.536 ;
  LAYER M2 ;
        RECT 6.844 8.44 9.316 8.472 ;
  LAYER M2 ;
        RECT 6.844 8.376 9.316 8.408 ;
  LAYER M2 ;
        RECT 6.844 8.312 9.316 8.344 ;
  LAYER M2 ;
        RECT 6.844 8.248 9.316 8.28 ;
  LAYER M2 ;
        RECT 6.844 8.184 9.316 8.216 ;
  LAYER M2 ;
        RECT 6.844 8.12 9.316 8.152 ;
  LAYER M2 ;
        RECT 6.844 8.056 9.316 8.088 ;
  LAYER M2 ;
        RECT 6.844 7.992 9.316 8.024 ;
  LAYER M2 ;
        RECT 6.844 7.928 9.316 7.96 ;
  LAYER M3 ;
        RECT 6.864 7.776 6.896 10.284 ;
  LAYER M3 ;
        RECT 6.928 7.776 6.96 10.284 ;
  LAYER M3 ;
        RECT 6.992 7.776 7.024 10.284 ;
  LAYER M3 ;
        RECT 7.056 7.776 7.088 10.284 ;
  LAYER M3 ;
        RECT 7.12 7.776 7.152 10.284 ;
  LAYER M3 ;
        RECT 7.184 7.776 7.216 10.284 ;
  LAYER M3 ;
        RECT 7.248 7.776 7.28 10.284 ;
  LAYER M3 ;
        RECT 7.312 7.776 7.344 10.284 ;
  LAYER M3 ;
        RECT 7.376 7.776 7.408 10.284 ;
  LAYER M3 ;
        RECT 7.44 7.776 7.472 10.284 ;
  LAYER M3 ;
        RECT 7.504 7.776 7.536 10.284 ;
  LAYER M3 ;
        RECT 7.568 7.776 7.6 10.284 ;
  LAYER M3 ;
        RECT 7.632 7.776 7.664 10.284 ;
  LAYER M3 ;
        RECT 7.696 7.776 7.728 10.284 ;
  LAYER M3 ;
        RECT 7.76 7.776 7.792 10.284 ;
  LAYER M3 ;
        RECT 7.824 7.776 7.856 10.284 ;
  LAYER M3 ;
        RECT 7.888 7.776 7.92 10.284 ;
  LAYER M3 ;
        RECT 7.952 7.776 7.984 10.284 ;
  LAYER M3 ;
        RECT 8.016 7.776 8.048 10.284 ;
  LAYER M3 ;
        RECT 8.08 7.776 8.112 10.284 ;
  LAYER M3 ;
        RECT 8.144 7.776 8.176 10.284 ;
  LAYER M3 ;
        RECT 8.208 7.776 8.24 10.284 ;
  LAYER M3 ;
        RECT 8.272 7.776 8.304 10.284 ;
  LAYER M3 ;
        RECT 8.336 7.776 8.368 10.284 ;
  LAYER M3 ;
        RECT 8.4 7.776 8.432 10.284 ;
  LAYER M3 ;
        RECT 8.464 7.776 8.496 10.284 ;
  LAYER M3 ;
        RECT 8.528 7.776 8.56 10.284 ;
  LAYER M3 ;
        RECT 8.592 7.776 8.624 10.284 ;
  LAYER M3 ;
        RECT 8.656 7.776 8.688 10.284 ;
  LAYER M3 ;
        RECT 8.72 7.776 8.752 10.284 ;
  LAYER M3 ;
        RECT 8.784 7.776 8.816 10.284 ;
  LAYER M3 ;
        RECT 8.848 7.776 8.88 10.284 ;
  LAYER M3 ;
        RECT 8.912 7.776 8.944 10.284 ;
  LAYER M3 ;
        RECT 8.976 7.776 9.008 10.284 ;
  LAYER M3 ;
        RECT 9.04 7.776 9.072 10.284 ;
  LAYER M3 ;
        RECT 9.104 7.776 9.136 10.284 ;
  LAYER M3 ;
        RECT 9.168 7.776 9.2 10.284 ;
  LAYER M3 ;
        RECT 9.264 7.776 9.296 10.284 ;
  LAYER M1 ;
        RECT 6.879 7.812 6.881 10.248 ;
  LAYER M1 ;
        RECT 6.959 7.812 6.961 10.248 ;
  LAYER M1 ;
        RECT 7.039 7.812 7.041 10.248 ;
  LAYER M1 ;
        RECT 7.119 7.812 7.121 10.248 ;
  LAYER M1 ;
        RECT 7.199 7.812 7.201 10.248 ;
  LAYER M1 ;
        RECT 7.279 7.812 7.281 10.248 ;
  LAYER M1 ;
        RECT 7.359 7.812 7.361 10.248 ;
  LAYER M1 ;
        RECT 7.439 7.812 7.441 10.248 ;
  LAYER M1 ;
        RECT 7.519 7.812 7.521 10.248 ;
  LAYER M1 ;
        RECT 7.599 7.812 7.601 10.248 ;
  LAYER M1 ;
        RECT 7.679 7.812 7.681 10.248 ;
  LAYER M1 ;
        RECT 7.759 7.812 7.761 10.248 ;
  LAYER M1 ;
        RECT 7.839 7.812 7.841 10.248 ;
  LAYER M1 ;
        RECT 7.919 7.812 7.921 10.248 ;
  LAYER M1 ;
        RECT 7.999 7.812 8.001 10.248 ;
  LAYER M1 ;
        RECT 8.079 7.812 8.081 10.248 ;
  LAYER M1 ;
        RECT 8.159 7.812 8.161 10.248 ;
  LAYER M1 ;
        RECT 8.239 7.812 8.241 10.248 ;
  LAYER M1 ;
        RECT 8.319 7.812 8.321 10.248 ;
  LAYER M1 ;
        RECT 8.399 7.812 8.401 10.248 ;
  LAYER M1 ;
        RECT 8.479 7.812 8.481 10.248 ;
  LAYER M1 ;
        RECT 8.559 7.812 8.561 10.248 ;
  LAYER M1 ;
        RECT 8.639 7.812 8.641 10.248 ;
  LAYER M1 ;
        RECT 8.719 7.812 8.721 10.248 ;
  LAYER M1 ;
        RECT 8.799 7.812 8.801 10.248 ;
  LAYER M1 ;
        RECT 8.879 7.812 8.881 10.248 ;
  LAYER M1 ;
        RECT 8.959 7.812 8.961 10.248 ;
  LAYER M1 ;
        RECT 9.039 7.812 9.041 10.248 ;
  LAYER M1 ;
        RECT 9.119 7.812 9.121 10.248 ;
  LAYER M1 ;
        RECT 9.199 7.812 9.201 10.248 ;
  LAYER M2 ;
        RECT 6.88 10.247 9.28 10.249 ;
  LAYER M2 ;
        RECT 6.88 10.163 9.28 10.165 ;
  LAYER M2 ;
        RECT 6.88 10.079 9.28 10.081 ;
  LAYER M2 ;
        RECT 6.88 9.995 9.28 9.997 ;
  LAYER M2 ;
        RECT 6.88 9.911 9.28 9.913 ;
  LAYER M2 ;
        RECT 6.88 9.827 9.28 9.829 ;
  LAYER M2 ;
        RECT 6.88 9.743 9.28 9.745 ;
  LAYER M2 ;
        RECT 6.88 9.659 9.28 9.661 ;
  LAYER M2 ;
        RECT 6.88 9.575 9.28 9.577 ;
  LAYER M2 ;
        RECT 6.88 9.491 9.28 9.493 ;
  LAYER M2 ;
        RECT 6.88 9.407 9.28 9.409 ;
  LAYER M2 ;
        RECT 6.88 9.323 9.28 9.325 ;
  LAYER M2 ;
        RECT 6.88 9.2395 9.28 9.2415 ;
  LAYER M2 ;
        RECT 6.88 9.155 9.28 9.157 ;
  LAYER M2 ;
        RECT 6.88 9.071 9.28 9.073 ;
  LAYER M2 ;
        RECT 6.88 8.987 9.28 8.989 ;
  LAYER M2 ;
        RECT 6.88 8.903 9.28 8.905 ;
  LAYER M2 ;
        RECT 6.88 8.819 9.28 8.821 ;
  LAYER M2 ;
        RECT 6.88 8.735 9.28 8.737 ;
  LAYER M2 ;
        RECT 6.88 8.651 9.28 8.653 ;
  LAYER M2 ;
        RECT 6.88 8.567 9.28 8.569 ;
  LAYER M2 ;
        RECT 6.88 8.483 9.28 8.485 ;
  LAYER M2 ;
        RECT 6.88 8.399 9.28 8.401 ;
  LAYER M2 ;
        RECT 6.88 8.315 9.28 8.317 ;
  LAYER M2 ;
        RECT 6.88 8.231 9.28 8.233 ;
  LAYER M2 ;
        RECT 6.88 8.147 9.28 8.149 ;
  LAYER M2 ;
        RECT 6.88 8.063 9.28 8.065 ;
  LAYER M2 ;
        RECT 6.88 7.979 9.28 7.981 ;
  LAYER M2 ;
        RECT 6.88 7.895 9.28 7.897 ;
  LAYER M1 ;
        RECT 6.864 4.836 6.896 7.344 ;
  LAYER M1 ;
        RECT 6.928 4.836 6.96 7.344 ;
  LAYER M1 ;
        RECT 6.992 4.836 7.024 7.344 ;
  LAYER M1 ;
        RECT 7.056 4.836 7.088 7.344 ;
  LAYER M1 ;
        RECT 7.12 4.836 7.152 7.344 ;
  LAYER M1 ;
        RECT 7.184 4.836 7.216 7.344 ;
  LAYER M1 ;
        RECT 7.248 4.836 7.28 7.344 ;
  LAYER M1 ;
        RECT 7.312 4.836 7.344 7.344 ;
  LAYER M1 ;
        RECT 7.376 4.836 7.408 7.344 ;
  LAYER M1 ;
        RECT 7.44 4.836 7.472 7.344 ;
  LAYER M1 ;
        RECT 7.504 4.836 7.536 7.344 ;
  LAYER M1 ;
        RECT 7.568 4.836 7.6 7.344 ;
  LAYER M1 ;
        RECT 7.632 4.836 7.664 7.344 ;
  LAYER M1 ;
        RECT 7.696 4.836 7.728 7.344 ;
  LAYER M1 ;
        RECT 7.76 4.836 7.792 7.344 ;
  LAYER M1 ;
        RECT 7.824 4.836 7.856 7.344 ;
  LAYER M1 ;
        RECT 7.888 4.836 7.92 7.344 ;
  LAYER M1 ;
        RECT 7.952 4.836 7.984 7.344 ;
  LAYER M1 ;
        RECT 8.016 4.836 8.048 7.344 ;
  LAYER M1 ;
        RECT 8.08 4.836 8.112 7.344 ;
  LAYER M1 ;
        RECT 8.144 4.836 8.176 7.344 ;
  LAYER M1 ;
        RECT 8.208 4.836 8.24 7.344 ;
  LAYER M1 ;
        RECT 8.272 4.836 8.304 7.344 ;
  LAYER M1 ;
        RECT 8.336 4.836 8.368 7.344 ;
  LAYER M1 ;
        RECT 8.4 4.836 8.432 7.344 ;
  LAYER M1 ;
        RECT 8.464 4.836 8.496 7.344 ;
  LAYER M1 ;
        RECT 8.528 4.836 8.56 7.344 ;
  LAYER M1 ;
        RECT 8.592 4.836 8.624 7.344 ;
  LAYER M1 ;
        RECT 8.656 4.836 8.688 7.344 ;
  LAYER M1 ;
        RECT 8.72 4.836 8.752 7.344 ;
  LAYER M1 ;
        RECT 8.784 4.836 8.816 7.344 ;
  LAYER M1 ;
        RECT 8.848 4.836 8.88 7.344 ;
  LAYER M1 ;
        RECT 8.912 4.836 8.944 7.344 ;
  LAYER M1 ;
        RECT 8.976 4.836 9.008 7.344 ;
  LAYER M1 ;
        RECT 9.04 4.836 9.072 7.344 ;
  LAYER M1 ;
        RECT 9.104 4.836 9.136 7.344 ;
  LAYER M1 ;
        RECT 9.168 4.836 9.2 7.344 ;
  LAYER M2 ;
        RECT 6.844 7.228 9.316 7.26 ;
  LAYER M2 ;
        RECT 6.844 7.164 9.316 7.196 ;
  LAYER M2 ;
        RECT 6.844 7.1 9.316 7.132 ;
  LAYER M2 ;
        RECT 6.844 7.036 9.316 7.068 ;
  LAYER M2 ;
        RECT 6.844 6.972 9.316 7.004 ;
  LAYER M2 ;
        RECT 6.844 6.908 9.316 6.94 ;
  LAYER M2 ;
        RECT 6.844 6.844 9.316 6.876 ;
  LAYER M2 ;
        RECT 6.844 6.78 9.316 6.812 ;
  LAYER M2 ;
        RECT 6.844 6.716 9.316 6.748 ;
  LAYER M2 ;
        RECT 6.844 6.652 9.316 6.684 ;
  LAYER M2 ;
        RECT 6.844 6.588 9.316 6.62 ;
  LAYER M2 ;
        RECT 6.844 6.524 9.316 6.556 ;
  LAYER M2 ;
        RECT 6.844 6.46 9.316 6.492 ;
  LAYER M2 ;
        RECT 6.844 6.396 9.316 6.428 ;
  LAYER M2 ;
        RECT 6.844 6.332 9.316 6.364 ;
  LAYER M2 ;
        RECT 6.844 6.268 9.316 6.3 ;
  LAYER M2 ;
        RECT 6.844 6.204 9.316 6.236 ;
  LAYER M2 ;
        RECT 6.844 6.14 9.316 6.172 ;
  LAYER M2 ;
        RECT 6.844 6.076 9.316 6.108 ;
  LAYER M2 ;
        RECT 6.844 6.012 9.316 6.044 ;
  LAYER M2 ;
        RECT 6.844 5.948 9.316 5.98 ;
  LAYER M2 ;
        RECT 6.844 5.884 9.316 5.916 ;
  LAYER M2 ;
        RECT 6.844 5.82 9.316 5.852 ;
  LAYER M2 ;
        RECT 6.844 5.756 9.316 5.788 ;
  LAYER M2 ;
        RECT 6.844 5.692 9.316 5.724 ;
  LAYER M2 ;
        RECT 6.844 5.628 9.316 5.66 ;
  LAYER M2 ;
        RECT 6.844 5.564 9.316 5.596 ;
  LAYER M2 ;
        RECT 6.844 5.5 9.316 5.532 ;
  LAYER M2 ;
        RECT 6.844 5.436 9.316 5.468 ;
  LAYER M2 ;
        RECT 6.844 5.372 9.316 5.404 ;
  LAYER M2 ;
        RECT 6.844 5.308 9.316 5.34 ;
  LAYER M2 ;
        RECT 6.844 5.244 9.316 5.276 ;
  LAYER M2 ;
        RECT 6.844 5.18 9.316 5.212 ;
  LAYER M2 ;
        RECT 6.844 5.116 9.316 5.148 ;
  LAYER M2 ;
        RECT 6.844 5.052 9.316 5.084 ;
  LAYER M2 ;
        RECT 6.844 4.988 9.316 5.02 ;
  LAYER M3 ;
        RECT 6.864 4.836 6.896 7.344 ;
  LAYER M3 ;
        RECT 6.928 4.836 6.96 7.344 ;
  LAYER M3 ;
        RECT 6.992 4.836 7.024 7.344 ;
  LAYER M3 ;
        RECT 7.056 4.836 7.088 7.344 ;
  LAYER M3 ;
        RECT 7.12 4.836 7.152 7.344 ;
  LAYER M3 ;
        RECT 7.184 4.836 7.216 7.344 ;
  LAYER M3 ;
        RECT 7.248 4.836 7.28 7.344 ;
  LAYER M3 ;
        RECT 7.312 4.836 7.344 7.344 ;
  LAYER M3 ;
        RECT 7.376 4.836 7.408 7.344 ;
  LAYER M3 ;
        RECT 7.44 4.836 7.472 7.344 ;
  LAYER M3 ;
        RECT 7.504 4.836 7.536 7.344 ;
  LAYER M3 ;
        RECT 7.568 4.836 7.6 7.344 ;
  LAYER M3 ;
        RECT 7.632 4.836 7.664 7.344 ;
  LAYER M3 ;
        RECT 7.696 4.836 7.728 7.344 ;
  LAYER M3 ;
        RECT 7.76 4.836 7.792 7.344 ;
  LAYER M3 ;
        RECT 7.824 4.836 7.856 7.344 ;
  LAYER M3 ;
        RECT 7.888 4.836 7.92 7.344 ;
  LAYER M3 ;
        RECT 7.952 4.836 7.984 7.344 ;
  LAYER M3 ;
        RECT 8.016 4.836 8.048 7.344 ;
  LAYER M3 ;
        RECT 8.08 4.836 8.112 7.344 ;
  LAYER M3 ;
        RECT 8.144 4.836 8.176 7.344 ;
  LAYER M3 ;
        RECT 8.208 4.836 8.24 7.344 ;
  LAYER M3 ;
        RECT 8.272 4.836 8.304 7.344 ;
  LAYER M3 ;
        RECT 8.336 4.836 8.368 7.344 ;
  LAYER M3 ;
        RECT 8.4 4.836 8.432 7.344 ;
  LAYER M3 ;
        RECT 8.464 4.836 8.496 7.344 ;
  LAYER M3 ;
        RECT 8.528 4.836 8.56 7.344 ;
  LAYER M3 ;
        RECT 8.592 4.836 8.624 7.344 ;
  LAYER M3 ;
        RECT 8.656 4.836 8.688 7.344 ;
  LAYER M3 ;
        RECT 8.72 4.836 8.752 7.344 ;
  LAYER M3 ;
        RECT 8.784 4.836 8.816 7.344 ;
  LAYER M3 ;
        RECT 8.848 4.836 8.88 7.344 ;
  LAYER M3 ;
        RECT 8.912 4.836 8.944 7.344 ;
  LAYER M3 ;
        RECT 8.976 4.836 9.008 7.344 ;
  LAYER M3 ;
        RECT 9.04 4.836 9.072 7.344 ;
  LAYER M3 ;
        RECT 9.104 4.836 9.136 7.344 ;
  LAYER M3 ;
        RECT 9.168 4.836 9.2 7.344 ;
  LAYER M3 ;
        RECT 9.264 4.836 9.296 7.344 ;
  LAYER M1 ;
        RECT 6.879 4.872 6.881 7.308 ;
  LAYER M1 ;
        RECT 6.959 4.872 6.961 7.308 ;
  LAYER M1 ;
        RECT 7.039 4.872 7.041 7.308 ;
  LAYER M1 ;
        RECT 7.119 4.872 7.121 7.308 ;
  LAYER M1 ;
        RECT 7.199 4.872 7.201 7.308 ;
  LAYER M1 ;
        RECT 7.279 4.872 7.281 7.308 ;
  LAYER M1 ;
        RECT 7.359 4.872 7.361 7.308 ;
  LAYER M1 ;
        RECT 7.439 4.872 7.441 7.308 ;
  LAYER M1 ;
        RECT 7.519 4.872 7.521 7.308 ;
  LAYER M1 ;
        RECT 7.599 4.872 7.601 7.308 ;
  LAYER M1 ;
        RECT 7.679 4.872 7.681 7.308 ;
  LAYER M1 ;
        RECT 7.759 4.872 7.761 7.308 ;
  LAYER M1 ;
        RECT 7.839 4.872 7.841 7.308 ;
  LAYER M1 ;
        RECT 7.919 4.872 7.921 7.308 ;
  LAYER M1 ;
        RECT 7.999 4.872 8.001 7.308 ;
  LAYER M1 ;
        RECT 8.079 4.872 8.081 7.308 ;
  LAYER M1 ;
        RECT 8.159 4.872 8.161 7.308 ;
  LAYER M1 ;
        RECT 8.239 4.872 8.241 7.308 ;
  LAYER M1 ;
        RECT 8.319 4.872 8.321 7.308 ;
  LAYER M1 ;
        RECT 8.399 4.872 8.401 7.308 ;
  LAYER M1 ;
        RECT 8.479 4.872 8.481 7.308 ;
  LAYER M1 ;
        RECT 8.559 4.872 8.561 7.308 ;
  LAYER M1 ;
        RECT 8.639 4.872 8.641 7.308 ;
  LAYER M1 ;
        RECT 8.719 4.872 8.721 7.308 ;
  LAYER M1 ;
        RECT 8.799 4.872 8.801 7.308 ;
  LAYER M1 ;
        RECT 8.879 4.872 8.881 7.308 ;
  LAYER M1 ;
        RECT 8.959 4.872 8.961 7.308 ;
  LAYER M1 ;
        RECT 9.039 4.872 9.041 7.308 ;
  LAYER M1 ;
        RECT 9.119 4.872 9.121 7.308 ;
  LAYER M1 ;
        RECT 9.199 4.872 9.201 7.308 ;
  LAYER M2 ;
        RECT 6.88 7.307 9.28 7.309 ;
  LAYER M2 ;
        RECT 6.88 7.223 9.28 7.225 ;
  LAYER M2 ;
        RECT 6.88 7.139 9.28 7.141 ;
  LAYER M2 ;
        RECT 6.88 7.055 9.28 7.057 ;
  LAYER M2 ;
        RECT 6.88 6.971 9.28 6.973 ;
  LAYER M2 ;
        RECT 6.88 6.887 9.28 6.889 ;
  LAYER M2 ;
        RECT 6.88 6.803 9.28 6.805 ;
  LAYER M2 ;
        RECT 6.88 6.719 9.28 6.721 ;
  LAYER M2 ;
        RECT 6.88 6.635 9.28 6.637 ;
  LAYER M2 ;
        RECT 6.88 6.551 9.28 6.553 ;
  LAYER M2 ;
        RECT 6.88 6.467 9.28 6.469 ;
  LAYER M2 ;
        RECT 6.88 6.383 9.28 6.385 ;
  LAYER M2 ;
        RECT 6.88 6.2995 9.28 6.3015 ;
  LAYER M2 ;
        RECT 6.88 6.215 9.28 6.217 ;
  LAYER M2 ;
        RECT 6.88 6.131 9.28 6.133 ;
  LAYER M2 ;
        RECT 6.88 6.047 9.28 6.049 ;
  LAYER M2 ;
        RECT 6.88 5.963 9.28 5.965 ;
  LAYER M2 ;
        RECT 6.88 5.879 9.28 5.881 ;
  LAYER M2 ;
        RECT 6.88 5.795 9.28 5.797 ;
  LAYER M2 ;
        RECT 6.88 5.711 9.28 5.713 ;
  LAYER M2 ;
        RECT 6.88 5.627 9.28 5.629 ;
  LAYER M2 ;
        RECT 6.88 5.543 9.28 5.545 ;
  LAYER M2 ;
        RECT 6.88 5.459 9.28 5.461 ;
  LAYER M2 ;
        RECT 6.88 5.375 9.28 5.377 ;
  LAYER M2 ;
        RECT 6.88 5.291 9.28 5.293 ;
  LAYER M2 ;
        RECT 6.88 5.207 9.28 5.209 ;
  LAYER M2 ;
        RECT 6.88 5.123 9.28 5.125 ;
  LAYER M2 ;
        RECT 6.88 5.039 9.28 5.041 ;
  LAYER M2 ;
        RECT 6.88 4.955 9.28 4.957 ;
  LAYER M1 ;
        RECT 6.864 1.896 6.896 4.404 ;
  LAYER M1 ;
        RECT 6.928 1.896 6.96 4.404 ;
  LAYER M1 ;
        RECT 6.992 1.896 7.024 4.404 ;
  LAYER M1 ;
        RECT 7.056 1.896 7.088 4.404 ;
  LAYER M1 ;
        RECT 7.12 1.896 7.152 4.404 ;
  LAYER M1 ;
        RECT 7.184 1.896 7.216 4.404 ;
  LAYER M1 ;
        RECT 7.248 1.896 7.28 4.404 ;
  LAYER M1 ;
        RECT 7.312 1.896 7.344 4.404 ;
  LAYER M1 ;
        RECT 7.376 1.896 7.408 4.404 ;
  LAYER M1 ;
        RECT 7.44 1.896 7.472 4.404 ;
  LAYER M1 ;
        RECT 7.504 1.896 7.536 4.404 ;
  LAYER M1 ;
        RECT 7.568 1.896 7.6 4.404 ;
  LAYER M1 ;
        RECT 7.632 1.896 7.664 4.404 ;
  LAYER M1 ;
        RECT 7.696 1.896 7.728 4.404 ;
  LAYER M1 ;
        RECT 7.76 1.896 7.792 4.404 ;
  LAYER M1 ;
        RECT 7.824 1.896 7.856 4.404 ;
  LAYER M1 ;
        RECT 7.888 1.896 7.92 4.404 ;
  LAYER M1 ;
        RECT 7.952 1.896 7.984 4.404 ;
  LAYER M1 ;
        RECT 8.016 1.896 8.048 4.404 ;
  LAYER M1 ;
        RECT 8.08 1.896 8.112 4.404 ;
  LAYER M1 ;
        RECT 8.144 1.896 8.176 4.404 ;
  LAYER M1 ;
        RECT 8.208 1.896 8.24 4.404 ;
  LAYER M1 ;
        RECT 8.272 1.896 8.304 4.404 ;
  LAYER M1 ;
        RECT 8.336 1.896 8.368 4.404 ;
  LAYER M1 ;
        RECT 8.4 1.896 8.432 4.404 ;
  LAYER M1 ;
        RECT 8.464 1.896 8.496 4.404 ;
  LAYER M1 ;
        RECT 8.528 1.896 8.56 4.404 ;
  LAYER M1 ;
        RECT 8.592 1.896 8.624 4.404 ;
  LAYER M1 ;
        RECT 8.656 1.896 8.688 4.404 ;
  LAYER M1 ;
        RECT 8.72 1.896 8.752 4.404 ;
  LAYER M1 ;
        RECT 8.784 1.896 8.816 4.404 ;
  LAYER M1 ;
        RECT 8.848 1.896 8.88 4.404 ;
  LAYER M1 ;
        RECT 8.912 1.896 8.944 4.404 ;
  LAYER M1 ;
        RECT 8.976 1.896 9.008 4.404 ;
  LAYER M1 ;
        RECT 9.04 1.896 9.072 4.404 ;
  LAYER M1 ;
        RECT 9.104 1.896 9.136 4.404 ;
  LAYER M1 ;
        RECT 9.168 1.896 9.2 4.404 ;
  LAYER M2 ;
        RECT 6.844 4.288 9.316 4.32 ;
  LAYER M2 ;
        RECT 6.844 4.224 9.316 4.256 ;
  LAYER M2 ;
        RECT 6.844 4.16 9.316 4.192 ;
  LAYER M2 ;
        RECT 6.844 4.096 9.316 4.128 ;
  LAYER M2 ;
        RECT 6.844 4.032 9.316 4.064 ;
  LAYER M2 ;
        RECT 6.844 3.968 9.316 4 ;
  LAYER M2 ;
        RECT 6.844 3.904 9.316 3.936 ;
  LAYER M2 ;
        RECT 6.844 3.84 9.316 3.872 ;
  LAYER M2 ;
        RECT 6.844 3.776 9.316 3.808 ;
  LAYER M2 ;
        RECT 6.844 3.712 9.316 3.744 ;
  LAYER M2 ;
        RECT 6.844 3.648 9.316 3.68 ;
  LAYER M2 ;
        RECT 6.844 3.584 9.316 3.616 ;
  LAYER M2 ;
        RECT 6.844 3.52 9.316 3.552 ;
  LAYER M2 ;
        RECT 6.844 3.456 9.316 3.488 ;
  LAYER M2 ;
        RECT 6.844 3.392 9.316 3.424 ;
  LAYER M2 ;
        RECT 6.844 3.328 9.316 3.36 ;
  LAYER M2 ;
        RECT 6.844 3.264 9.316 3.296 ;
  LAYER M2 ;
        RECT 6.844 3.2 9.316 3.232 ;
  LAYER M2 ;
        RECT 6.844 3.136 9.316 3.168 ;
  LAYER M2 ;
        RECT 6.844 3.072 9.316 3.104 ;
  LAYER M2 ;
        RECT 6.844 3.008 9.316 3.04 ;
  LAYER M2 ;
        RECT 6.844 2.944 9.316 2.976 ;
  LAYER M2 ;
        RECT 6.844 2.88 9.316 2.912 ;
  LAYER M2 ;
        RECT 6.844 2.816 9.316 2.848 ;
  LAYER M2 ;
        RECT 6.844 2.752 9.316 2.784 ;
  LAYER M2 ;
        RECT 6.844 2.688 9.316 2.72 ;
  LAYER M2 ;
        RECT 6.844 2.624 9.316 2.656 ;
  LAYER M2 ;
        RECT 6.844 2.56 9.316 2.592 ;
  LAYER M2 ;
        RECT 6.844 2.496 9.316 2.528 ;
  LAYER M2 ;
        RECT 6.844 2.432 9.316 2.464 ;
  LAYER M2 ;
        RECT 6.844 2.368 9.316 2.4 ;
  LAYER M2 ;
        RECT 6.844 2.304 9.316 2.336 ;
  LAYER M2 ;
        RECT 6.844 2.24 9.316 2.272 ;
  LAYER M2 ;
        RECT 6.844 2.176 9.316 2.208 ;
  LAYER M2 ;
        RECT 6.844 2.112 9.316 2.144 ;
  LAYER M2 ;
        RECT 6.844 2.048 9.316 2.08 ;
  LAYER M3 ;
        RECT 6.864 1.896 6.896 4.404 ;
  LAYER M3 ;
        RECT 6.928 1.896 6.96 4.404 ;
  LAYER M3 ;
        RECT 6.992 1.896 7.024 4.404 ;
  LAYER M3 ;
        RECT 7.056 1.896 7.088 4.404 ;
  LAYER M3 ;
        RECT 7.12 1.896 7.152 4.404 ;
  LAYER M3 ;
        RECT 7.184 1.896 7.216 4.404 ;
  LAYER M3 ;
        RECT 7.248 1.896 7.28 4.404 ;
  LAYER M3 ;
        RECT 7.312 1.896 7.344 4.404 ;
  LAYER M3 ;
        RECT 7.376 1.896 7.408 4.404 ;
  LAYER M3 ;
        RECT 7.44 1.896 7.472 4.404 ;
  LAYER M3 ;
        RECT 7.504 1.896 7.536 4.404 ;
  LAYER M3 ;
        RECT 7.568 1.896 7.6 4.404 ;
  LAYER M3 ;
        RECT 7.632 1.896 7.664 4.404 ;
  LAYER M3 ;
        RECT 7.696 1.896 7.728 4.404 ;
  LAYER M3 ;
        RECT 7.76 1.896 7.792 4.404 ;
  LAYER M3 ;
        RECT 7.824 1.896 7.856 4.404 ;
  LAYER M3 ;
        RECT 7.888 1.896 7.92 4.404 ;
  LAYER M3 ;
        RECT 7.952 1.896 7.984 4.404 ;
  LAYER M3 ;
        RECT 8.016 1.896 8.048 4.404 ;
  LAYER M3 ;
        RECT 8.08 1.896 8.112 4.404 ;
  LAYER M3 ;
        RECT 8.144 1.896 8.176 4.404 ;
  LAYER M3 ;
        RECT 8.208 1.896 8.24 4.404 ;
  LAYER M3 ;
        RECT 8.272 1.896 8.304 4.404 ;
  LAYER M3 ;
        RECT 8.336 1.896 8.368 4.404 ;
  LAYER M3 ;
        RECT 8.4 1.896 8.432 4.404 ;
  LAYER M3 ;
        RECT 8.464 1.896 8.496 4.404 ;
  LAYER M3 ;
        RECT 8.528 1.896 8.56 4.404 ;
  LAYER M3 ;
        RECT 8.592 1.896 8.624 4.404 ;
  LAYER M3 ;
        RECT 8.656 1.896 8.688 4.404 ;
  LAYER M3 ;
        RECT 8.72 1.896 8.752 4.404 ;
  LAYER M3 ;
        RECT 8.784 1.896 8.816 4.404 ;
  LAYER M3 ;
        RECT 8.848 1.896 8.88 4.404 ;
  LAYER M3 ;
        RECT 8.912 1.896 8.944 4.404 ;
  LAYER M3 ;
        RECT 8.976 1.896 9.008 4.404 ;
  LAYER M3 ;
        RECT 9.04 1.896 9.072 4.404 ;
  LAYER M3 ;
        RECT 9.104 1.896 9.136 4.404 ;
  LAYER M3 ;
        RECT 9.168 1.896 9.2 4.404 ;
  LAYER M3 ;
        RECT 9.264 1.896 9.296 4.404 ;
  LAYER M1 ;
        RECT 6.879 1.932 6.881 4.368 ;
  LAYER M1 ;
        RECT 6.959 1.932 6.961 4.368 ;
  LAYER M1 ;
        RECT 7.039 1.932 7.041 4.368 ;
  LAYER M1 ;
        RECT 7.119 1.932 7.121 4.368 ;
  LAYER M1 ;
        RECT 7.199 1.932 7.201 4.368 ;
  LAYER M1 ;
        RECT 7.279 1.932 7.281 4.368 ;
  LAYER M1 ;
        RECT 7.359 1.932 7.361 4.368 ;
  LAYER M1 ;
        RECT 7.439 1.932 7.441 4.368 ;
  LAYER M1 ;
        RECT 7.519 1.932 7.521 4.368 ;
  LAYER M1 ;
        RECT 7.599 1.932 7.601 4.368 ;
  LAYER M1 ;
        RECT 7.679 1.932 7.681 4.368 ;
  LAYER M1 ;
        RECT 7.759 1.932 7.761 4.368 ;
  LAYER M1 ;
        RECT 7.839 1.932 7.841 4.368 ;
  LAYER M1 ;
        RECT 7.919 1.932 7.921 4.368 ;
  LAYER M1 ;
        RECT 7.999 1.932 8.001 4.368 ;
  LAYER M1 ;
        RECT 8.079 1.932 8.081 4.368 ;
  LAYER M1 ;
        RECT 8.159 1.932 8.161 4.368 ;
  LAYER M1 ;
        RECT 8.239 1.932 8.241 4.368 ;
  LAYER M1 ;
        RECT 8.319 1.932 8.321 4.368 ;
  LAYER M1 ;
        RECT 8.399 1.932 8.401 4.368 ;
  LAYER M1 ;
        RECT 8.479 1.932 8.481 4.368 ;
  LAYER M1 ;
        RECT 8.559 1.932 8.561 4.368 ;
  LAYER M1 ;
        RECT 8.639 1.932 8.641 4.368 ;
  LAYER M1 ;
        RECT 8.719 1.932 8.721 4.368 ;
  LAYER M1 ;
        RECT 8.799 1.932 8.801 4.368 ;
  LAYER M1 ;
        RECT 8.879 1.932 8.881 4.368 ;
  LAYER M1 ;
        RECT 8.959 1.932 8.961 4.368 ;
  LAYER M1 ;
        RECT 9.039 1.932 9.041 4.368 ;
  LAYER M1 ;
        RECT 9.119 1.932 9.121 4.368 ;
  LAYER M1 ;
        RECT 9.199 1.932 9.201 4.368 ;
  LAYER M2 ;
        RECT 6.88 4.367 9.28 4.369 ;
  LAYER M2 ;
        RECT 6.88 4.283 9.28 4.285 ;
  LAYER M2 ;
        RECT 6.88 4.199 9.28 4.201 ;
  LAYER M2 ;
        RECT 6.88 4.115 9.28 4.117 ;
  LAYER M2 ;
        RECT 6.88 4.031 9.28 4.033 ;
  LAYER M2 ;
        RECT 6.88 3.947 9.28 3.949 ;
  LAYER M2 ;
        RECT 6.88 3.863 9.28 3.865 ;
  LAYER M2 ;
        RECT 6.88 3.779 9.28 3.781 ;
  LAYER M2 ;
        RECT 6.88 3.695 9.28 3.697 ;
  LAYER M2 ;
        RECT 6.88 3.611 9.28 3.613 ;
  LAYER M2 ;
        RECT 6.88 3.527 9.28 3.529 ;
  LAYER M2 ;
        RECT 6.88 3.443 9.28 3.445 ;
  LAYER M2 ;
        RECT 6.88 3.3595 9.28 3.3615 ;
  LAYER M2 ;
        RECT 6.88 3.275 9.28 3.277 ;
  LAYER M2 ;
        RECT 6.88 3.191 9.28 3.193 ;
  LAYER M2 ;
        RECT 6.88 3.107 9.28 3.109 ;
  LAYER M2 ;
        RECT 6.88 3.023 9.28 3.025 ;
  LAYER M2 ;
        RECT 6.88 2.939 9.28 2.941 ;
  LAYER M2 ;
        RECT 6.88 2.855 9.28 2.857 ;
  LAYER M2 ;
        RECT 6.88 2.771 9.28 2.773 ;
  LAYER M2 ;
        RECT 6.88 2.687 9.28 2.689 ;
  LAYER M2 ;
        RECT 6.88 2.603 9.28 2.605 ;
  LAYER M2 ;
        RECT 6.88 2.519 9.28 2.521 ;
  LAYER M2 ;
        RECT 6.88 2.435 9.28 2.437 ;
  LAYER M2 ;
        RECT 6.88 2.351 9.28 2.353 ;
  LAYER M2 ;
        RECT 6.88 2.267 9.28 2.269 ;
  LAYER M2 ;
        RECT 6.88 2.183 9.28 2.185 ;
  LAYER M2 ;
        RECT 6.88 2.099 9.28 2.101 ;
  LAYER M2 ;
        RECT 6.88 2.015 9.28 2.017 ;
  LAYER M1 ;
        RECT 9.744 13.656 9.776 16.164 ;
  LAYER M1 ;
        RECT 9.808 13.656 9.84 16.164 ;
  LAYER M1 ;
        RECT 9.872 13.656 9.904 16.164 ;
  LAYER M1 ;
        RECT 9.936 13.656 9.968 16.164 ;
  LAYER M1 ;
        RECT 10 13.656 10.032 16.164 ;
  LAYER M1 ;
        RECT 10.064 13.656 10.096 16.164 ;
  LAYER M1 ;
        RECT 10.128 13.656 10.16 16.164 ;
  LAYER M1 ;
        RECT 10.192 13.656 10.224 16.164 ;
  LAYER M1 ;
        RECT 10.256 13.656 10.288 16.164 ;
  LAYER M1 ;
        RECT 10.32 13.656 10.352 16.164 ;
  LAYER M1 ;
        RECT 10.384 13.656 10.416 16.164 ;
  LAYER M1 ;
        RECT 10.448 13.656 10.48 16.164 ;
  LAYER M1 ;
        RECT 10.512 13.656 10.544 16.164 ;
  LAYER M1 ;
        RECT 10.576 13.656 10.608 16.164 ;
  LAYER M1 ;
        RECT 10.64 13.656 10.672 16.164 ;
  LAYER M1 ;
        RECT 10.704 13.656 10.736 16.164 ;
  LAYER M1 ;
        RECT 10.768 13.656 10.8 16.164 ;
  LAYER M1 ;
        RECT 10.832 13.656 10.864 16.164 ;
  LAYER M1 ;
        RECT 10.896 13.656 10.928 16.164 ;
  LAYER M1 ;
        RECT 10.96 13.656 10.992 16.164 ;
  LAYER M1 ;
        RECT 11.024 13.656 11.056 16.164 ;
  LAYER M1 ;
        RECT 11.088 13.656 11.12 16.164 ;
  LAYER M1 ;
        RECT 11.152 13.656 11.184 16.164 ;
  LAYER M1 ;
        RECT 11.216 13.656 11.248 16.164 ;
  LAYER M1 ;
        RECT 11.28 13.656 11.312 16.164 ;
  LAYER M1 ;
        RECT 11.344 13.656 11.376 16.164 ;
  LAYER M1 ;
        RECT 11.408 13.656 11.44 16.164 ;
  LAYER M1 ;
        RECT 11.472 13.656 11.504 16.164 ;
  LAYER M1 ;
        RECT 11.536 13.656 11.568 16.164 ;
  LAYER M1 ;
        RECT 11.6 13.656 11.632 16.164 ;
  LAYER M1 ;
        RECT 11.664 13.656 11.696 16.164 ;
  LAYER M1 ;
        RECT 11.728 13.656 11.76 16.164 ;
  LAYER M1 ;
        RECT 11.792 13.656 11.824 16.164 ;
  LAYER M1 ;
        RECT 11.856 13.656 11.888 16.164 ;
  LAYER M1 ;
        RECT 11.92 13.656 11.952 16.164 ;
  LAYER M1 ;
        RECT 11.984 13.656 12.016 16.164 ;
  LAYER M1 ;
        RECT 12.048 13.656 12.08 16.164 ;
  LAYER M2 ;
        RECT 9.724 16.048 12.196 16.08 ;
  LAYER M2 ;
        RECT 9.724 15.984 12.196 16.016 ;
  LAYER M2 ;
        RECT 9.724 15.92 12.196 15.952 ;
  LAYER M2 ;
        RECT 9.724 15.856 12.196 15.888 ;
  LAYER M2 ;
        RECT 9.724 15.792 12.196 15.824 ;
  LAYER M2 ;
        RECT 9.724 15.728 12.196 15.76 ;
  LAYER M2 ;
        RECT 9.724 15.664 12.196 15.696 ;
  LAYER M2 ;
        RECT 9.724 15.6 12.196 15.632 ;
  LAYER M2 ;
        RECT 9.724 15.536 12.196 15.568 ;
  LAYER M2 ;
        RECT 9.724 15.472 12.196 15.504 ;
  LAYER M2 ;
        RECT 9.724 15.408 12.196 15.44 ;
  LAYER M2 ;
        RECT 9.724 15.344 12.196 15.376 ;
  LAYER M2 ;
        RECT 9.724 15.28 12.196 15.312 ;
  LAYER M2 ;
        RECT 9.724 15.216 12.196 15.248 ;
  LAYER M2 ;
        RECT 9.724 15.152 12.196 15.184 ;
  LAYER M2 ;
        RECT 9.724 15.088 12.196 15.12 ;
  LAYER M2 ;
        RECT 9.724 15.024 12.196 15.056 ;
  LAYER M2 ;
        RECT 9.724 14.96 12.196 14.992 ;
  LAYER M2 ;
        RECT 9.724 14.896 12.196 14.928 ;
  LAYER M2 ;
        RECT 9.724 14.832 12.196 14.864 ;
  LAYER M2 ;
        RECT 9.724 14.768 12.196 14.8 ;
  LAYER M2 ;
        RECT 9.724 14.704 12.196 14.736 ;
  LAYER M2 ;
        RECT 9.724 14.64 12.196 14.672 ;
  LAYER M2 ;
        RECT 9.724 14.576 12.196 14.608 ;
  LAYER M2 ;
        RECT 9.724 14.512 12.196 14.544 ;
  LAYER M2 ;
        RECT 9.724 14.448 12.196 14.48 ;
  LAYER M2 ;
        RECT 9.724 14.384 12.196 14.416 ;
  LAYER M2 ;
        RECT 9.724 14.32 12.196 14.352 ;
  LAYER M2 ;
        RECT 9.724 14.256 12.196 14.288 ;
  LAYER M2 ;
        RECT 9.724 14.192 12.196 14.224 ;
  LAYER M2 ;
        RECT 9.724 14.128 12.196 14.16 ;
  LAYER M2 ;
        RECT 9.724 14.064 12.196 14.096 ;
  LAYER M2 ;
        RECT 9.724 14 12.196 14.032 ;
  LAYER M2 ;
        RECT 9.724 13.936 12.196 13.968 ;
  LAYER M2 ;
        RECT 9.724 13.872 12.196 13.904 ;
  LAYER M2 ;
        RECT 9.724 13.808 12.196 13.84 ;
  LAYER M3 ;
        RECT 9.744 13.656 9.776 16.164 ;
  LAYER M3 ;
        RECT 9.808 13.656 9.84 16.164 ;
  LAYER M3 ;
        RECT 9.872 13.656 9.904 16.164 ;
  LAYER M3 ;
        RECT 9.936 13.656 9.968 16.164 ;
  LAYER M3 ;
        RECT 10 13.656 10.032 16.164 ;
  LAYER M3 ;
        RECT 10.064 13.656 10.096 16.164 ;
  LAYER M3 ;
        RECT 10.128 13.656 10.16 16.164 ;
  LAYER M3 ;
        RECT 10.192 13.656 10.224 16.164 ;
  LAYER M3 ;
        RECT 10.256 13.656 10.288 16.164 ;
  LAYER M3 ;
        RECT 10.32 13.656 10.352 16.164 ;
  LAYER M3 ;
        RECT 10.384 13.656 10.416 16.164 ;
  LAYER M3 ;
        RECT 10.448 13.656 10.48 16.164 ;
  LAYER M3 ;
        RECT 10.512 13.656 10.544 16.164 ;
  LAYER M3 ;
        RECT 10.576 13.656 10.608 16.164 ;
  LAYER M3 ;
        RECT 10.64 13.656 10.672 16.164 ;
  LAYER M3 ;
        RECT 10.704 13.656 10.736 16.164 ;
  LAYER M3 ;
        RECT 10.768 13.656 10.8 16.164 ;
  LAYER M3 ;
        RECT 10.832 13.656 10.864 16.164 ;
  LAYER M3 ;
        RECT 10.896 13.656 10.928 16.164 ;
  LAYER M3 ;
        RECT 10.96 13.656 10.992 16.164 ;
  LAYER M3 ;
        RECT 11.024 13.656 11.056 16.164 ;
  LAYER M3 ;
        RECT 11.088 13.656 11.12 16.164 ;
  LAYER M3 ;
        RECT 11.152 13.656 11.184 16.164 ;
  LAYER M3 ;
        RECT 11.216 13.656 11.248 16.164 ;
  LAYER M3 ;
        RECT 11.28 13.656 11.312 16.164 ;
  LAYER M3 ;
        RECT 11.344 13.656 11.376 16.164 ;
  LAYER M3 ;
        RECT 11.408 13.656 11.44 16.164 ;
  LAYER M3 ;
        RECT 11.472 13.656 11.504 16.164 ;
  LAYER M3 ;
        RECT 11.536 13.656 11.568 16.164 ;
  LAYER M3 ;
        RECT 11.6 13.656 11.632 16.164 ;
  LAYER M3 ;
        RECT 11.664 13.656 11.696 16.164 ;
  LAYER M3 ;
        RECT 11.728 13.656 11.76 16.164 ;
  LAYER M3 ;
        RECT 11.792 13.656 11.824 16.164 ;
  LAYER M3 ;
        RECT 11.856 13.656 11.888 16.164 ;
  LAYER M3 ;
        RECT 11.92 13.656 11.952 16.164 ;
  LAYER M3 ;
        RECT 11.984 13.656 12.016 16.164 ;
  LAYER M3 ;
        RECT 12.048 13.656 12.08 16.164 ;
  LAYER M3 ;
        RECT 12.144 13.656 12.176 16.164 ;
  LAYER M1 ;
        RECT 9.759 13.692 9.761 16.128 ;
  LAYER M1 ;
        RECT 9.839 13.692 9.841 16.128 ;
  LAYER M1 ;
        RECT 9.919 13.692 9.921 16.128 ;
  LAYER M1 ;
        RECT 9.999 13.692 10.001 16.128 ;
  LAYER M1 ;
        RECT 10.079 13.692 10.081 16.128 ;
  LAYER M1 ;
        RECT 10.159 13.692 10.161 16.128 ;
  LAYER M1 ;
        RECT 10.239 13.692 10.241 16.128 ;
  LAYER M1 ;
        RECT 10.319 13.692 10.321 16.128 ;
  LAYER M1 ;
        RECT 10.399 13.692 10.401 16.128 ;
  LAYER M1 ;
        RECT 10.479 13.692 10.481 16.128 ;
  LAYER M1 ;
        RECT 10.559 13.692 10.561 16.128 ;
  LAYER M1 ;
        RECT 10.639 13.692 10.641 16.128 ;
  LAYER M1 ;
        RECT 10.719 13.692 10.721 16.128 ;
  LAYER M1 ;
        RECT 10.799 13.692 10.801 16.128 ;
  LAYER M1 ;
        RECT 10.879 13.692 10.881 16.128 ;
  LAYER M1 ;
        RECT 10.959 13.692 10.961 16.128 ;
  LAYER M1 ;
        RECT 11.039 13.692 11.041 16.128 ;
  LAYER M1 ;
        RECT 11.119 13.692 11.121 16.128 ;
  LAYER M1 ;
        RECT 11.199 13.692 11.201 16.128 ;
  LAYER M1 ;
        RECT 11.279 13.692 11.281 16.128 ;
  LAYER M1 ;
        RECT 11.359 13.692 11.361 16.128 ;
  LAYER M1 ;
        RECT 11.439 13.692 11.441 16.128 ;
  LAYER M1 ;
        RECT 11.519 13.692 11.521 16.128 ;
  LAYER M1 ;
        RECT 11.599 13.692 11.601 16.128 ;
  LAYER M1 ;
        RECT 11.679 13.692 11.681 16.128 ;
  LAYER M1 ;
        RECT 11.759 13.692 11.761 16.128 ;
  LAYER M1 ;
        RECT 11.839 13.692 11.841 16.128 ;
  LAYER M1 ;
        RECT 11.919 13.692 11.921 16.128 ;
  LAYER M1 ;
        RECT 11.999 13.692 12.001 16.128 ;
  LAYER M1 ;
        RECT 12.079 13.692 12.081 16.128 ;
  LAYER M2 ;
        RECT 9.76 16.127 12.16 16.129 ;
  LAYER M2 ;
        RECT 9.76 16.043 12.16 16.045 ;
  LAYER M2 ;
        RECT 9.76 15.959 12.16 15.961 ;
  LAYER M2 ;
        RECT 9.76 15.875 12.16 15.877 ;
  LAYER M2 ;
        RECT 9.76 15.791 12.16 15.793 ;
  LAYER M2 ;
        RECT 9.76 15.707 12.16 15.709 ;
  LAYER M2 ;
        RECT 9.76 15.623 12.16 15.625 ;
  LAYER M2 ;
        RECT 9.76 15.539 12.16 15.541 ;
  LAYER M2 ;
        RECT 9.76 15.455 12.16 15.457 ;
  LAYER M2 ;
        RECT 9.76 15.371 12.16 15.373 ;
  LAYER M2 ;
        RECT 9.76 15.287 12.16 15.289 ;
  LAYER M2 ;
        RECT 9.76 15.203 12.16 15.205 ;
  LAYER M2 ;
        RECT 9.76 15.1195 12.16 15.1215 ;
  LAYER M2 ;
        RECT 9.76 15.035 12.16 15.037 ;
  LAYER M2 ;
        RECT 9.76 14.951 12.16 14.953 ;
  LAYER M2 ;
        RECT 9.76 14.867 12.16 14.869 ;
  LAYER M2 ;
        RECT 9.76 14.783 12.16 14.785 ;
  LAYER M2 ;
        RECT 9.76 14.699 12.16 14.701 ;
  LAYER M2 ;
        RECT 9.76 14.615 12.16 14.617 ;
  LAYER M2 ;
        RECT 9.76 14.531 12.16 14.533 ;
  LAYER M2 ;
        RECT 9.76 14.447 12.16 14.449 ;
  LAYER M2 ;
        RECT 9.76 14.363 12.16 14.365 ;
  LAYER M2 ;
        RECT 9.76 14.279 12.16 14.281 ;
  LAYER M2 ;
        RECT 9.76 14.195 12.16 14.197 ;
  LAYER M2 ;
        RECT 9.76 14.111 12.16 14.113 ;
  LAYER M2 ;
        RECT 9.76 14.027 12.16 14.029 ;
  LAYER M2 ;
        RECT 9.76 13.943 12.16 13.945 ;
  LAYER M2 ;
        RECT 9.76 13.859 12.16 13.861 ;
  LAYER M2 ;
        RECT 9.76 13.775 12.16 13.777 ;
  LAYER M1 ;
        RECT 9.744 10.716 9.776 13.224 ;
  LAYER M1 ;
        RECT 9.808 10.716 9.84 13.224 ;
  LAYER M1 ;
        RECT 9.872 10.716 9.904 13.224 ;
  LAYER M1 ;
        RECT 9.936 10.716 9.968 13.224 ;
  LAYER M1 ;
        RECT 10 10.716 10.032 13.224 ;
  LAYER M1 ;
        RECT 10.064 10.716 10.096 13.224 ;
  LAYER M1 ;
        RECT 10.128 10.716 10.16 13.224 ;
  LAYER M1 ;
        RECT 10.192 10.716 10.224 13.224 ;
  LAYER M1 ;
        RECT 10.256 10.716 10.288 13.224 ;
  LAYER M1 ;
        RECT 10.32 10.716 10.352 13.224 ;
  LAYER M1 ;
        RECT 10.384 10.716 10.416 13.224 ;
  LAYER M1 ;
        RECT 10.448 10.716 10.48 13.224 ;
  LAYER M1 ;
        RECT 10.512 10.716 10.544 13.224 ;
  LAYER M1 ;
        RECT 10.576 10.716 10.608 13.224 ;
  LAYER M1 ;
        RECT 10.64 10.716 10.672 13.224 ;
  LAYER M1 ;
        RECT 10.704 10.716 10.736 13.224 ;
  LAYER M1 ;
        RECT 10.768 10.716 10.8 13.224 ;
  LAYER M1 ;
        RECT 10.832 10.716 10.864 13.224 ;
  LAYER M1 ;
        RECT 10.896 10.716 10.928 13.224 ;
  LAYER M1 ;
        RECT 10.96 10.716 10.992 13.224 ;
  LAYER M1 ;
        RECT 11.024 10.716 11.056 13.224 ;
  LAYER M1 ;
        RECT 11.088 10.716 11.12 13.224 ;
  LAYER M1 ;
        RECT 11.152 10.716 11.184 13.224 ;
  LAYER M1 ;
        RECT 11.216 10.716 11.248 13.224 ;
  LAYER M1 ;
        RECT 11.28 10.716 11.312 13.224 ;
  LAYER M1 ;
        RECT 11.344 10.716 11.376 13.224 ;
  LAYER M1 ;
        RECT 11.408 10.716 11.44 13.224 ;
  LAYER M1 ;
        RECT 11.472 10.716 11.504 13.224 ;
  LAYER M1 ;
        RECT 11.536 10.716 11.568 13.224 ;
  LAYER M1 ;
        RECT 11.6 10.716 11.632 13.224 ;
  LAYER M1 ;
        RECT 11.664 10.716 11.696 13.224 ;
  LAYER M1 ;
        RECT 11.728 10.716 11.76 13.224 ;
  LAYER M1 ;
        RECT 11.792 10.716 11.824 13.224 ;
  LAYER M1 ;
        RECT 11.856 10.716 11.888 13.224 ;
  LAYER M1 ;
        RECT 11.92 10.716 11.952 13.224 ;
  LAYER M1 ;
        RECT 11.984 10.716 12.016 13.224 ;
  LAYER M1 ;
        RECT 12.048 10.716 12.08 13.224 ;
  LAYER M2 ;
        RECT 9.724 13.108 12.196 13.14 ;
  LAYER M2 ;
        RECT 9.724 13.044 12.196 13.076 ;
  LAYER M2 ;
        RECT 9.724 12.98 12.196 13.012 ;
  LAYER M2 ;
        RECT 9.724 12.916 12.196 12.948 ;
  LAYER M2 ;
        RECT 9.724 12.852 12.196 12.884 ;
  LAYER M2 ;
        RECT 9.724 12.788 12.196 12.82 ;
  LAYER M2 ;
        RECT 9.724 12.724 12.196 12.756 ;
  LAYER M2 ;
        RECT 9.724 12.66 12.196 12.692 ;
  LAYER M2 ;
        RECT 9.724 12.596 12.196 12.628 ;
  LAYER M2 ;
        RECT 9.724 12.532 12.196 12.564 ;
  LAYER M2 ;
        RECT 9.724 12.468 12.196 12.5 ;
  LAYER M2 ;
        RECT 9.724 12.404 12.196 12.436 ;
  LAYER M2 ;
        RECT 9.724 12.34 12.196 12.372 ;
  LAYER M2 ;
        RECT 9.724 12.276 12.196 12.308 ;
  LAYER M2 ;
        RECT 9.724 12.212 12.196 12.244 ;
  LAYER M2 ;
        RECT 9.724 12.148 12.196 12.18 ;
  LAYER M2 ;
        RECT 9.724 12.084 12.196 12.116 ;
  LAYER M2 ;
        RECT 9.724 12.02 12.196 12.052 ;
  LAYER M2 ;
        RECT 9.724 11.956 12.196 11.988 ;
  LAYER M2 ;
        RECT 9.724 11.892 12.196 11.924 ;
  LAYER M2 ;
        RECT 9.724 11.828 12.196 11.86 ;
  LAYER M2 ;
        RECT 9.724 11.764 12.196 11.796 ;
  LAYER M2 ;
        RECT 9.724 11.7 12.196 11.732 ;
  LAYER M2 ;
        RECT 9.724 11.636 12.196 11.668 ;
  LAYER M2 ;
        RECT 9.724 11.572 12.196 11.604 ;
  LAYER M2 ;
        RECT 9.724 11.508 12.196 11.54 ;
  LAYER M2 ;
        RECT 9.724 11.444 12.196 11.476 ;
  LAYER M2 ;
        RECT 9.724 11.38 12.196 11.412 ;
  LAYER M2 ;
        RECT 9.724 11.316 12.196 11.348 ;
  LAYER M2 ;
        RECT 9.724 11.252 12.196 11.284 ;
  LAYER M2 ;
        RECT 9.724 11.188 12.196 11.22 ;
  LAYER M2 ;
        RECT 9.724 11.124 12.196 11.156 ;
  LAYER M2 ;
        RECT 9.724 11.06 12.196 11.092 ;
  LAYER M2 ;
        RECT 9.724 10.996 12.196 11.028 ;
  LAYER M2 ;
        RECT 9.724 10.932 12.196 10.964 ;
  LAYER M2 ;
        RECT 9.724 10.868 12.196 10.9 ;
  LAYER M3 ;
        RECT 9.744 10.716 9.776 13.224 ;
  LAYER M3 ;
        RECT 9.808 10.716 9.84 13.224 ;
  LAYER M3 ;
        RECT 9.872 10.716 9.904 13.224 ;
  LAYER M3 ;
        RECT 9.936 10.716 9.968 13.224 ;
  LAYER M3 ;
        RECT 10 10.716 10.032 13.224 ;
  LAYER M3 ;
        RECT 10.064 10.716 10.096 13.224 ;
  LAYER M3 ;
        RECT 10.128 10.716 10.16 13.224 ;
  LAYER M3 ;
        RECT 10.192 10.716 10.224 13.224 ;
  LAYER M3 ;
        RECT 10.256 10.716 10.288 13.224 ;
  LAYER M3 ;
        RECT 10.32 10.716 10.352 13.224 ;
  LAYER M3 ;
        RECT 10.384 10.716 10.416 13.224 ;
  LAYER M3 ;
        RECT 10.448 10.716 10.48 13.224 ;
  LAYER M3 ;
        RECT 10.512 10.716 10.544 13.224 ;
  LAYER M3 ;
        RECT 10.576 10.716 10.608 13.224 ;
  LAYER M3 ;
        RECT 10.64 10.716 10.672 13.224 ;
  LAYER M3 ;
        RECT 10.704 10.716 10.736 13.224 ;
  LAYER M3 ;
        RECT 10.768 10.716 10.8 13.224 ;
  LAYER M3 ;
        RECT 10.832 10.716 10.864 13.224 ;
  LAYER M3 ;
        RECT 10.896 10.716 10.928 13.224 ;
  LAYER M3 ;
        RECT 10.96 10.716 10.992 13.224 ;
  LAYER M3 ;
        RECT 11.024 10.716 11.056 13.224 ;
  LAYER M3 ;
        RECT 11.088 10.716 11.12 13.224 ;
  LAYER M3 ;
        RECT 11.152 10.716 11.184 13.224 ;
  LAYER M3 ;
        RECT 11.216 10.716 11.248 13.224 ;
  LAYER M3 ;
        RECT 11.28 10.716 11.312 13.224 ;
  LAYER M3 ;
        RECT 11.344 10.716 11.376 13.224 ;
  LAYER M3 ;
        RECT 11.408 10.716 11.44 13.224 ;
  LAYER M3 ;
        RECT 11.472 10.716 11.504 13.224 ;
  LAYER M3 ;
        RECT 11.536 10.716 11.568 13.224 ;
  LAYER M3 ;
        RECT 11.6 10.716 11.632 13.224 ;
  LAYER M3 ;
        RECT 11.664 10.716 11.696 13.224 ;
  LAYER M3 ;
        RECT 11.728 10.716 11.76 13.224 ;
  LAYER M3 ;
        RECT 11.792 10.716 11.824 13.224 ;
  LAYER M3 ;
        RECT 11.856 10.716 11.888 13.224 ;
  LAYER M3 ;
        RECT 11.92 10.716 11.952 13.224 ;
  LAYER M3 ;
        RECT 11.984 10.716 12.016 13.224 ;
  LAYER M3 ;
        RECT 12.048 10.716 12.08 13.224 ;
  LAYER M3 ;
        RECT 12.144 10.716 12.176 13.224 ;
  LAYER M1 ;
        RECT 9.759 10.752 9.761 13.188 ;
  LAYER M1 ;
        RECT 9.839 10.752 9.841 13.188 ;
  LAYER M1 ;
        RECT 9.919 10.752 9.921 13.188 ;
  LAYER M1 ;
        RECT 9.999 10.752 10.001 13.188 ;
  LAYER M1 ;
        RECT 10.079 10.752 10.081 13.188 ;
  LAYER M1 ;
        RECT 10.159 10.752 10.161 13.188 ;
  LAYER M1 ;
        RECT 10.239 10.752 10.241 13.188 ;
  LAYER M1 ;
        RECT 10.319 10.752 10.321 13.188 ;
  LAYER M1 ;
        RECT 10.399 10.752 10.401 13.188 ;
  LAYER M1 ;
        RECT 10.479 10.752 10.481 13.188 ;
  LAYER M1 ;
        RECT 10.559 10.752 10.561 13.188 ;
  LAYER M1 ;
        RECT 10.639 10.752 10.641 13.188 ;
  LAYER M1 ;
        RECT 10.719 10.752 10.721 13.188 ;
  LAYER M1 ;
        RECT 10.799 10.752 10.801 13.188 ;
  LAYER M1 ;
        RECT 10.879 10.752 10.881 13.188 ;
  LAYER M1 ;
        RECT 10.959 10.752 10.961 13.188 ;
  LAYER M1 ;
        RECT 11.039 10.752 11.041 13.188 ;
  LAYER M1 ;
        RECT 11.119 10.752 11.121 13.188 ;
  LAYER M1 ;
        RECT 11.199 10.752 11.201 13.188 ;
  LAYER M1 ;
        RECT 11.279 10.752 11.281 13.188 ;
  LAYER M1 ;
        RECT 11.359 10.752 11.361 13.188 ;
  LAYER M1 ;
        RECT 11.439 10.752 11.441 13.188 ;
  LAYER M1 ;
        RECT 11.519 10.752 11.521 13.188 ;
  LAYER M1 ;
        RECT 11.599 10.752 11.601 13.188 ;
  LAYER M1 ;
        RECT 11.679 10.752 11.681 13.188 ;
  LAYER M1 ;
        RECT 11.759 10.752 11.761 13.188 ;
  LAYER M1 ;
        RECT 11.839 10.752 11.841 13.188 ;
  LAYER M1 ;
        RECT 11.919 10.752 11.921 13.188 ;
  LAYER M1 ;
        RECT 11.999 10.752 12.001 13.188 ;
  LAYER M1 ;
        RECT 12.079 10.752 12.081 13.188 ;
  LAYER M2 ;
        RECT 9.76 13.187 12.16 13.189 ;
  LAYER M2 ;
        RECT 9.76 13.103 12.16 13.105 ;
  LAYER M2 ;
        RECT 9.76 13.019 12.16 13.021 ;
  LAYER M2 ;
        RECT 9.76 12.935 12.16 12.937 ;
  LAYER M2 ;
        RECT 9.76 12.851 12.16 12.853 ;
  LAYER M2 ;
        RECT 9.76 12.767 12.16 12.769 ;
  LAYER M2 ;
        RECT 9.76 12.683 12.16 12.685 ;
  LAYER M2 ;
        RECT 9.76 12.599 12.16 12.601 ;
  LAYER M2 ;
        RECT 9.76 12.515 12.16 12.517 ;
  LAYER M2 ;
        RECT 9.76 12.431 12.16 12.433 ;
  LAYER M2 ;
        RECT 9.76 12.347 12.16 12.349 ;
  LAYER M2 ;
        RECT 9.76 12.263 12.16 12.265 ;
  LAYER M2 ;
        RECT 9.76 12.1795 12.16 12.1815 ;
  LAYER M2 ;
        RECT 9.76 12.095 12.16 12.097 ;
  LAYER M2 ;
        RECT 9.76 12.011 12.16 12.013 ;
  LAYER M2 ;
        RECT 9.76 11.927 12.16 11.929 ;
  LAYER M2 ;
        RECT 9.76 11.843 12.16 11.845 ;
  LAYER M2 ;
        RECT 9.76 11.759 12.16 11.761 ;
  LAYER M2 ;
        RECT 9.76 11.675 12.16 11.677 ;
  LAYER M2 ;
        RECT 9.76 11.591 12.16 11.593 ;
  LAYER M2 ;
        RECT 9.76 11.507 12.16 11.509 ;
  LAYER M2 ;
        RECT 9.76 11.423 12.16 11.425 ;
  LAYER M2 ;
        RECT 9.76 11.339 12.16 11.341 ;
  LAYER M2 ;
        RECT 9.76 11.255 12.16 11.257 ;
  LAYER M2 ;
        RECT 9.76 11.171 12.16 11.173 ;
  LAYER M2 ;
        RECT 9.76 11.087 12.16 11.089 ;
  LAYER M2 ;
        RECT 9.76 11.003 12.16 11.005 ;
  LAYER M2 ;
        RECT 9.76 10.919 12.16 10.921 ;
  LAYER M2 ;
        RECT 9.76 10.835 12.16 10.837 ;
  LAYER M1 ;
        RECT 9.744 7.776 9.776 10.284 ;
  LAYER M1 ;
        RECT 9.808 7.776 9.84 10.284 ;
  LAYER M1 ;
        RECT 9.872 7.776 9.904 10.284 ;
  LAYER M1 ;
        RECT 9.936 7.776 9.968 10.284 ;
  LAYER M1 ;
        RECT 10 7.776 10.032 10.284 ;
  LAYER M1 ;
        RECT 10.064 7.776 10.096 10.284 ;
  LAYER M1 ;
        RECT 10.128 7.776 10.16 10.284 ;
  LAYER M1 ;
        RECT 10.192 7.776 10.224 10.284 ;
  LAYER M1 ;
        RECT 10.256 7.776 10.288 10.284 ;
  LAYER M1 ;
        RECT 10.32 7.776 10.352 10.284 ;
  LAYER M1 ;
        RECT 10.384 7.776 10.416 10.284 ;
  LAYER M1 ;
        RECT 10.448 7.776 10.48 10.284 ;
  LAYER M1 ;
        RECT 10.512 7.776 10.544 10.284 ;
  LAYER M1 ;
        RECT 10.576 7.776 10.608 10.284 ;
  LAYER M1 ;
        RECT 10.64 7.776 10.672 10.284 ;
  LAYER M1 ;
        RECT 10.704 7.776 10.736 10.284 ;
  LAYER M1 ;
        RECT 10.768 7.776 10.8 10.284 ;
  LAYER M1 ;
        RECT 10.832 7.776 10.864 10.284 ;
  LAYER M1 ;
        RECT 10.896 7.776 10.928 10.284 ;
  LAYER M1 ;
        RECT 10.96 7.776 10.992 10.284 ;
  LAYER M1 ;
        RECT 11.024 7.776 11.056 10.284 ;
  LAYER M1 ;
        RECT 11.088 7.776 11.12 10.284 ;
  LAYER M1 ;
        RECT 11.152 7.776 11.184 10.284 ;
  LAYER M1 ;
        RECT 11.216 7.776 11.248 10.284 ;
  LAYER M1 ;
        RECT 11.28 7.776 11.312 10.284 ;
  LAYER M1 ;
        RECT 11.344 7.776 11.376 10.284 ;
  LAYER M1 ;
        RECT 11.408 7.776 11.44 10.284 ;
  LAYER M1 ;
        RECT 11.472 7.776 11.504 10.284 ;
  LAYER M1 ;
        RECT 11.536 7.776 11.568 10.284 ;
  LAYER M1 ;
        RECT 11.6 7.776 11.632 10.284 ;
  LAYER M1 ;
        RECT 11.664 7.776 11.696 10.284 ;
  LAYER M1 ;
        RECT 11.728 7.776 11.76 10.284 ;
  LAYER M1 ;
        RECT 11.792 7.776 11.824 10.284 ;
  LAYER M1 ;
        RECT 11.856 7.776 11.888 10.284 ;
  LAYER M1 ;
        RECT 11.92 7.776 11.952 10.284 ;
  LAYER M1 ;
        RECT 11.984 7.776 12.016 10.284 ;
  LAYER M1 ;
        RECT 12.048 7.776 12.08 10.284 ;
  LAYER M2 ;
        RECT 9.724 10.168 12.196 10.2 ;
  LAYER M2 ;
        RECT 9.724 10.104 12.196 10.136 ;
  LAYER M2 ;
        RECT 9.724 10.04 12.196 10.072 ;
  LAYER M2 ;
        RECT 9.724 9.976 12.196 10.008 ;
  LAYER M2 ;
        RECT 9.724 9.912 12.196 9.944 ;
  LAYER M2 ;
        RECT 9.724 9.848 12.196 9.88 ;
  LAYER M2 ;
        RECT 9.724 9.784 12.196 9.816 ;
  LAYER M2 ;
        RECT 9.724 9.72 12.196 9.752 ;
  LAYER M2 ;
        RECT 9.724 9.656 12.196 9.688 ;
  LAYER M2 ;
        RECT 9.724 9.592 12.196 9.624 ;
  LAYER M2 ;
        RECT 9.724 9.528 12.196 9.56 ;
  LAYER M2 ;
        RECT 9.724 9.464 12.196 9.496 ;
  LAYER M2 ;
        RECT 9.724 9.4 12.196 9.432 ;
  LAYER M2 ;
        RECT 9.724 9.336 12.196 9.368 ;
  LAYER M2 ;
        RECT 9.724 9.272 12.196 9.304 ;
  LAYER M2 ;
        RECT 9.724 9.208 12.196 9.24 ;
  LAYER M2 ;
        RECT 9.724 9.144 12.196 9.176 ;
  LAYER M2 ;
        RECT 9.724 9.08 12.196 9.112 ;
  LAYER M2 ;
        RECT 9.724 9.016 12.196 9.048 ;
  LAYER M2 ;
        RECT 9.724 8.952 12.196 8.984 ;
  LAYER M2 ;
        RECT 9.724 8.888 12.196 8.92 ;
  LAYER M2 ;
        RECT 9.724 8.824 12.196 8.856 ;
  LAYER M2 ;
        RECT 9.724 8.76 12.196 8.792 ;
  LAYER M2 ;
        RECT 9.724 8.696 12.196 8.728 ;
  LAYER M2 ;
        RECT 9.724 8.632 12.196 8.664 ;
  LAYER M2 ;
        RECT 9.724 8.568 12.196 8.6 ;
  LAYER M2 ;
        RECT 9.724 8.504 12.196 8.536 ;
  LAYER M2 ;
        RECT 9.724 8.44 12.196 8.472 ;
  LAYER M2 ;
        RECT 9.724 8.376 12.196 8.408 ;
  LAYER M2 ;
        RECT 9.724 8.312 12.196 8.344 ;
  LAYER M2 ;
        RECT 9.724 8.248 12.196 8.28 ;
  LAYER M2 ;
        RECT 9.724 8.184 12.196 8.216 ;
  LAYER M2 ;
        RECT 9.724 8.12 12.196 8.152 ;
  LAYER M2 ;
        RECT 9.724 8.056 12.196 8.088 ;
  LAYER M2 ;
        RECT 9.724 7.992 12.196 8.024 ;
  LAYER M2 ;
        RECT 9.724 7.928 12.196 7.96 ;
  LAYER M3 ;
        RECT 9.744 7.776 9.776 10.284 ;
  LAYER M3 ;
        RECT 9.808 7.776 9.84 10.284 ;
  LAYER M3 ;
        RECT 9.872 7.776 9.904 10.284 ;
  LAYER M3 ;
        RECT 9.936 7.776 9.968 10.284 ;
  LAYER M3 ;
        RECT 10 7.776 10.032 10.284 ;
  LAYER M3 ;
        RECT 10.064 7.776 10.096 10.284 ;
  LAYER M3 ;
        RECT 10.128 7.776 10.16 10.284 ;
  LAYER M3 ;
        RECT 10.192 7.776 10.224 10.284 ;
  LAYER M3 ;
        RECT 10.256 7.776 10.288 10.284 ;
  LAYER M3 ;
        RECT 10.32 7.776 10.352 10.284 ;
  LAYER M3 ;
        RECT 10.384 7.776 10.416 10.284 ;
  LAYER M3 ;
        RECT 10.448 7.776 10.48 10.284 ;
  LAYER M3 ;
        RECT 10.512 7.776 10.544 10.284 ;
  LAYER M3 ;
        RECT 10.576 7.776 10.608 10.284 ;
  LAYER M3 ;
        RECT 10.64 7.776 10.672 10.284 ;
  LAYER M3 ;
        RECT 10.704 7.776 10.736 10.284 ;
  LAYER M3 ;
        RECT 10.768 7.776 10.8 10.284 ;
  LAYER M3 ;
        RECT 10.832 7.776 10.864 10.284 ;
  LAYER M3 ;
        RECT 10.896 7.776 10.928 10.284 ;
  LAYER M3 ;
        RECT 10.96 7.776 10.992 10.284 ;
  LAYER M3 ;
        RECT 11.024 7.776 11.056 10.284 ;
  LAYER M3 ;
        RECT 11.088 7.776 11.12 10.284 ;
  LAYER M3 ;
        RECT 11.152 7.776 11.184 10.284 ;
  LAYER M3 ;
        RECT 11.216 7.776 11.248 10.284 ;
  LAYER M3 ;
        RECT 11.28 7.776 11.312 10.284 ;
  LAYER M3 ;
        RECT 11.344 7.776 11.376 10.284 ;
  LAYER M3 ;
        RECT 11.408 7.776 11.44 10.284 ;
  LAYER M3 ;
        RECT 11.472 7.776 11.504 10.284 ;
  LAYER M3 ;
        RECT 11.536 7.776 11.568 10.284 ;
  LAYER M3 ;
        RECT 11.6 7.776 11.632 10.284 ;
  LAYER M3 ;
        RECT 11.664 7.776 11.696 10.284 ;
  LAYER M3 ;
        RECT 11.728 7.776 11.76 10.284 ;
  LAYER M3 ;
        RECT 11.792 7.776 11.824 10.284 ;
  LAYER M3 ;
        RECT 11.856 7.776 11.888 10.284 ;
  LAYER M3 ;
        RECT 11.92 7.776 11.952 10.284 ;
  LAYER M3 ;
        RECT 11.984 7.776 12.016 10.284 ;
  LAYER M3 ;
        RECT 12.048 7.776 12.08 10.284 ;
  LAYER M3 ;
        RECT 12.144 7.776 12.176 10.284 ;
  LAYER M1 ;
        RECT 9.759 7.812 9.761 10.248 ;
  LAYER M1 ;
        RECT 9.839 7.812 9.841 10.248 ;
  LAYER M1 ;
        RECT 9.919 7.812 9.921 10.248 ;
  LAYER M1 ;
        RECT 9.999 7.812 10.001 10.248 ;
  LAYER M1 ;
        RECT 10.079 7.812 10.081 10.248 ;
  LAYER M1 ;
        RECT 10.159 7.812 10.161 10.248 ;
  LAYER M1 ;
        RECT 10.239 7.812 10.241 10.248 ;
  LAYER M1 ;
        RECT 10.319 7.812 10.321 10.248 ;
  LAYER M1 ;
        RECT 10.399 7.812 10.401 10.248 ;
  LAYER M1 ;
        RECT 10.479 7.812 10.481 10.248 ;
  LAYER M1 ;
        RECT 10.559 7.812 10.561 10.248 ;
  LAYER M1 ;
        RECT 10.639 7.812 10.641 10.248 ;
  LAYER M1 ;
        RECT 10.719 7.812 10.721 10.248 ;
  LAYER M1 ;
        RECT 10.799 7.812 10.801 10.248 ;
  LAYER M1 ;
        RECT 10.879 7.812 10.881 10.248 ;
  LAYER M1 ;
        RECT 10.959 7.812 10.961 10.248 ;
  LAYER M1 ;
        RECT 11.039 7.812 11.041 10.248 ;
  LAYER M1 ;
        RECT 11.119 7.812 11.121 10.248 ;
  LAYER M1 ;
        RECT 11.199 7.812 11.201 10.248 ;
  LAYER M1 ;
        RECT 11.279 7.812 11.281 10.248 ;
  LAYER M1 ;
        RECT 11.359 7.812 11.361 10.248 ;
  LAYER M1 ;
        RECT 11.439 7.812 11.441 10.248 ;
  LAYER M1 ;
        RECT 11.519 7.812 11.521 10.248 ;
  LAYER M1 ;
        RECT 11.599 7.812 11.601 10.248 ;
  LAYER M1 ;
        RECT 11.679 7.812 11.681 10.248 ;
  LAYER M1 ;
        RECT 11.759 7.812 11.761 10.248 ;
  LAYER M1 ;
        RECT 11.839 7.812 11.841 10.248 ;
  LAYER M1 ;
        RECT 11.919 7.812 11.921 10.248 ;
  LAYER M1 ;
        RECT 11.999 7.812 12.001 10.248 ;
  LAYER M1 ;
        RECT 12.079 7.812 12.081 10.248 ;
  LAYER M2 ;
        RECT 9.76 10.247 12.16 10.249 ;
  LAYER M2 ;
        RECT 9.76 10.163 12.16 10.165 ;
  LAYER M2 ;
        RECT 9.76 10.079 12.16 10.081 ;
  LAYER M2 ;
        RECT 9.76 9.995 12.16 9.997 ;
  LAYER M2 ;
        RECT 9.76 9.911 12.16 9.913 ;
  LAYER M2 ;
        RECT 9.76 9.827 12.16 9.829 ;
  LAYER M2 ;
        RECT 9.76 9.743 12.16 9.745 ;
  LAYER M2 ;
        RECT 9.76 9.659 12.16 9.661 ;
  LAYER M2 ;
        RECT 9.76 9.575 12.16 9.577 ;
  LAYER M2 ;
        RECT 9.76 9.491 12.16 9.493 ;
  LAYER M2 ;
        RECT 9.76 9.407 12.16 9.409 ;
  LAYER M2 ;
        RECT 9.76 9.323 12.16 9.325 ;
  LAYER M2 ;
        RECT 9.76 9.2395 12.16 9.2415 ;
  LAYER M2 ;
        RECT 9.76 9.155 12.16 9.157 ;
  LAYER M2 ;
        RECT 9.76 9.071 12.16 9.073 ;
  LAYER M2 ;
        RECT 9.76 8.987 12.16 8.989 ;
  LAYER M2 ;
        RECT 9.76 8.903 12.16 8.905 ;
  LAYER M2 ;
        RECT 9.76 8.819 12.16 8.821 ;
  LAYER M2 ;
        RECT 9.76 8.735 12.16 8.737 ;
  LAYER M2 ;
        RECT 9.76 8.651 12.16 8.653 ;
  LAYER M2 ;
        RECT 9.76 8.567 12.16 8.569 ;
  LAYER M2 ;
        RECT 9.76 8.483 12.16 8.485 ;
  LAYER M2 ;
        RECT 9.76 8.399 12.16 8.401 ;
  LAYER M2 ;
        RECT 9.76 8.315 12.16 8.317 ;
  LAYER M2 ;
        RECT 9.76 8.231 12.16 8.233 ;
  LAYER M2 ;
        RECT 9.76 8.147 12.16 8.149 ;
  LAYER M2 ;
        RECT 9.76 8.063 12.16 8.065 ;
  LAYER M2 ;
        RECT 9.76 7.979 12.16 7.981 ;
  LAYER M2 ;
        RECT 9.76 7.895 12.16 7.897 ;
  LAYER M1 ;
        RECT 9.744 4.836 9.776 7.344 ;
  LAYER M1 ;
        RECT 9.808 4.836 9.84 7.344 ;
  LAYER M1 ;
        RECT 9.872 4.836 9.904 7.344 ;
  LAYER M1 ;
        RECT 9.936 4.836 9.968 7.344 ;
  LAYER M1 ;
        RECT 10 4.836 10.032 7.344 ;
  LAYER M1 ;
        RECT 10.064 4.836 10.096 7.344 ;
  LAYER M1 ;
        RECT 10.128 4.836 10.16 7.344 ;
  LAYER M1 ;
        RECT 10.192 4.836 10.224 7.344 ;
  LAYER M1 ;
        RECT 10.256 4.836 10.288 7.344 ;
  LAYER M1 ;
        RECT 10.32 4.836 10.352 7.344 ;
  LAYER M1 ;
        RECT 10.384 4.836 10.416 7.344 ;
  LAYER M1 ;
        RECT 10.448 4.836 10.48 7.344 ;
  LAYER M1 ;
        RECT 10.512 4.836 10.544 7.344 ;
  LAYER M1 ;
        RECT 10.576 4.836 10.608 7.344 ;
  LAYER M1 ;
        RECT 10.64 4.836 10.672 7.344 ;
  LAYER M1 ;
        RECT 10.704 4.836 10.736 7.344 ;
  LAYER M1 ;
        RECT 10.768 4.836 10.8 7.344 ;
  LAYER M1 ;
        RECT 10.832 4.836 10.864 7.344 ;
  LAYER M1 ;
        RECT 10.896 4.836 10.928 7.344 ;
  LAYER M1 ;
        RECT 10.96 4.836 10.992 7.344 ;
  LAYER M1 ;
        RECT 11.024 4.836 11.056 7.344 ;
  LAYER M1 ;
        RECT 11.088 4.836 11.12 7.344 ;
  LAYER M1 ;
        RECT 11.152 4.836 11.184 7.344 ;
  LAYER M1 ;
        RECT 11.216 4.836 11.248 7.344 ;
  LAYER M1 ;
        RECT 11.28 4.836 11.312 7.344 ;
  LAYER M1 ;
        RECT 11.344 4.836 11.376 7.344 ;
  LAYER M1 ;
        RECT 11.408 4.836 11.44 7.344 ;
  LAYER M1 ;
        RECT 11.472 4.836 11.504 7.344 ;
  LAYER M1 ;
        RECT 11.536 4.836 11.568 7.344 ;
  LAYER M1 ;
        RECT 11.6 4.836 11.632 7.344 ;
  LAYER M1 ;
        RECT 11.664 4.836 11.696 7.344 ;
  LAYER M1 ;
        RECT 11.728 4.836 11.76 7.344 ;
  LAYER M1 ;
        RECT 11.792 4.836 11.824 7.344 ;
  LAYER M1 ;
        RECT 11.856 4.836 11.888 7.344 ;
  LAYER M1 ;
        RECT 11.92 4.836 11.952 7.344 ;
  LAYER M1 ;
        RECT 11.984 4.836 12.016 7.344 ;
  LAYER M1 ;
        RECT 12.048 4.836 12.08 7.344 ;
  LAYER M2 ;
        RECT 9.724 7.228 12.196 7.26 ;
  LAYER M2 ;
        RECT 9.724 7.164 12.196 7.196 ;
  LAYER M2 ;
        RECT 9.724 7.1 12.196 7.132 ;
  LAYER M2 ;
        RECT 9.724 7.036 12.196 7.068 ;
  LAYER M2 ;
        RECT 9.724 6.972 12.196 7.004 ;
  LAYER M2 ;
        RECT 9.724 6.908 12.196 6.94 ;
  LAYER M2 ;
        RECT 9.724 6.844 12.196 6.876 ;
  LAYER M2 ;
        RECT 9.724 6.78 12.196 6.812 ;
  LAYER M2 ;
        RECT 9.724 6.716 12.196 6.748 ;
  LAYER M2 ;
        RECT 9.724 6.652 12.196 6.684 ;
  LAYER M2 ;
        RECT 9.724 6.588 12.196 6.62 ;
  LAYER M2 ;
        RECT 9.724 6.524 12.196 6.556 ;
  LAYER M2 ;
        RECT 9.724 6.46 12.196 6.492 ;
  LAYER M2 ;
        RECT 9.724 6.396 12.196 6.428 ;
  LAYER M2 ;
        RECT 9.724 6.332 12.196 6.364 ;
  LAYER M2 ;
        RECT 9.724 6.268 12.196 6.3 ;
  LAYER M2 ;
        RECT 9.724 6.204 12.196 6.236 ;
  LAYER M2 ;
        RECT 9.724 6.14 12.196 6.172 ;
  LAYER M2 ;
        RECT 9.724 6.076 12.196 6.108 ;
  LAYER M2 ;
        RECT 9.724 6.012 12.196 6.044 ;
  LAYER M2 ;
        RECT 9.724 5.948 12.196 5.98 ;
  LAYER M2 ;
        RECT 9.724 5.884 12.196 5.916 ;
  LAYER M2 ;
        RECT 9.724 5.82 12.196 5.852 ;
  LAYER M2 ;
        RECT 9.724 5.756 12.196 5.788 ;
  LAYER M2 ;
        RECT 9.724 5.692 12.196 5.724 ;
  LAYER M2 ;
        RECT 9.724 5.628 12.196 5.66 ;
  LAYER M2 ;
        RECT 9.724 5.564 12.196 5.596 ;
  LAYER M2 ;
        RECT 9.724 5.5 12.196 5.532 ;
  LAYER M2 ;
        RECT 9.724 5.436 12.196 5.468 ;
  LAYER M2 ;
        RECT 9.724 5.372 12.196 5.404 ;
  LAYER M2 ;
        RECT 9.724 5.308 12.196 5.34 ;
  LAYER M2 ;
        RECT 9.724 5.244 12.196 5.276 ;
  LAYER M2 ;
        RECT 9.724 5.18 12.196 5.212 ;
  LAYER M2 ;
        RECT 9.724 5.116 12.196 5.148 ;
  LAYER M2 ;
        RECT 9.724 5.052 12.196 5.084 ;
  LAYER M2 ;
        RECT 9.724 4.988 12.196 5.02 ;
  LAYER M3 ;
        RECT 9.744 4.836 9.776 7.344 ;
  LAYER M3 ;
        RECT 9.808 4.836 9.84 7.344 ;
  LAYER M3 ;
        RECT 9.872 4.836 9.904 7.344 ;
  LAYER M3 ;
        RECT 9.936 4.836 9.968 7.344 ;
  LAYER M3 ;
        RECT 10 4.836 10.032 7.344 ;
  LAYER M3 ;
        RECT 10.064 4.836 10.096 7.344 ;
  LAYER M3 ;
        RECT 10.128 4.836 10.16 7.344 ;
  LAYER M3 ;
        RECT 10.192 4.836 10.224 7.344 ;
  LAYER M3 ;
        RECT 10.256 4.836 10.288 7.344 ;
  LAYER M3 ;
        RECT 10.32 4.836 10.352 7.344 ;
  LAYER M3 ;
        RECT 10.384 4.836 10.416 7.344 ;
  LAYER M3 ;
        RECT 10.448 4.836 10.48 7.344 ;
  LAYER M3 ;
        RECT 10.512 4.836 10.544 7.344 ;
  LAYER M3 ;
        RECT 10.576 4.836 10.608 7.344 ;
  LAYER M3 ;
        RECT 10.64 4.836 10.672 7.344 ;
  LAYER M3 ;
        RECT 10.704 4.836 10.736 7.344 ;
  LAYER M3 ;
        RECT 10.768 4.836 10.8 7.344 ;
  LAYER M3 ;
        RECT 10.832 4.836 10.864 7.344 ;
  LAYER M3 ;
        RECT 10.896 4.836 10.928 7.344 ;
  LAYER M3 ;
        RECT 10.96 4.836 10.992 7.344 ;
  LAYER M3 ;
        RECT 11.024 4.836 11.056 7.344 ;
  LAYER M3 ;
        RECT 11.088 4.836 11.12 7.344 ;
  LAYER M3 ;
        RECT 11.152 4.836 11.184 7.344 ;
  LAYER M3 ;
        RECT 11.216 4.836 11.248 7.344 ;
  LAYER M3 ;
        RECT 11.28 4.836 11.312 7.344 ;
  LAYER M3 ;
        RECT 11.344 4.836 11.376 7.344 ;
  LAYER M3 ;
        RECT 11.408 4.836 11.44 7.344 ;
  LAYER M3 ;
        RECT 11.472 4.836 11.504 7.344 ;
  LAYER M3 ;
        RECT 11.536 4.836 11.568 7.344 ;
  LAYER M3 ;
        RECT 11.6 4.836 11.632 7.344 ;
  LAYER M3 ;
        RECT 11.664 4.836 11.696 7.344 ;
  LAYER M3 ;
        RECT 11.728 4.836 11.76 7.344 ;
  LAYER M3 ;
        RECT 11.792 4.836 11.824 7.344 ;
  LAYER M3 ;
        RECT 11.856 4.836 11.888 7.344 ;
  LAYER M3 ;
        RECT 11.92 4.836 11.952 7.344 ;
  LAYER M3 ;
        RECT 11.984 4.836 12.016 7.344 ;
  LAYER M3 ;
        RECT 12.048 4.836 12.08 7.344 ;
  LAYER M3 ;
        RECT 12.144 4.836 12.176 7.344 ;
  LAYER M1 ;
        RECT 9.759 4.872 9.761 7.308 ;
  LAYER M1 ;
        RECT 9.839 4.872 9.841 7.308 ;
  LAYER M1 ;
        RECT 9.919 4.872 9.921 7.308 ;
  LAYER M1 ;
        RECT 9.999 4.872 10.001 7.308 ;
  LAYER M1 ;
        RECT 10.079 4.872 10.081 7.308 ;
  LAYER M1 ;
        RECT 10.159 4.872 10.161 7.308 ;
  LAYER M1 ;
        RECT 10.239 4.872 10.241 7.308 ;
  LAYER M1 ;
        RECT 10.319 4.872 10.321 7.308 ;
  LAYER M1 ;
        RECT 10.399 4.872 10.401 7.308 ;
  LAYER M1 ;
        RECT 10.479 4.872 10.481 7.308 ;
  LAYER M1 ;
        RECT 10.559 4.872 10.561 7.308 ;
  LAYER M1 ;
        RECT 10.639 4.872 10.641 7.308 ;
  LAYER M1 ;
        RECT 10.719 4.872 10.721 7.308 ;
  LAYER M1 ;
        RECT 10.799 4.872 10.801 7.308 ;
  LAYER M1 ;
        RECT 10.879 4.872 10.881 7.308 ;
  LAYER M1 ;
        RECT 10.959 4.872 10.961 7.308 ;
  LAYER M1 ;
        RECT 11.039 4.872 11.041 7.308 ;
  LAYER M1 ;
        RECT 11.119 4.872 11.121 7.308 ;
  LAYER M1 ;
        RECT 11.199 4.872 11.201 7.308 ;
  LAYER M1 ;
        RECT 11.279 4.872 11.281 7.308 ;
  LAYER M1 ;
        RECT 11.359 4.872 11.361 7.308 ;
  LAYER M1 ;
        RECT 11.439 4.872 11.441 7.308 ;
  LAYER M1 ;
        RECT 11.519 4.872 11.521 7.308 ;
  LAYER M1 ;
        RECT 11.599 4.872 11.601 7.308 ;
  LAYER M1 ;
        RECT 11.679 4.872 11.681 7.308 ;
  LAYER M1 ;
        RECT 11.759 4.872 11.761 7.308 ;
  LAYER M1 ;
        RECT 11.839 4.872 11.841 7.308 ;
  LAYER M1 ;
        RECT 11.919 4.872 11.921 7.308 ;
  LAYER M1 ;
        RECT 11.999 4.872 12.001 7.308 ;
  LAYER M1 ;
        RECT 12.079 4.872 12.081 7.308 ;
  LAYER M2 ;
        RECT 9.76 7.307 12.16 7.309 ;
  LAYER M2 ;
        RECT 9.76 7.223 12.16 7.225 ;
  LAYER M2 ;
        RECT 9.76 7.139 12.16 7.141 ;
  LAYER M2 ;
        RECT 9.76 7.055 12.16 7.057 ;
  LAYER M2 ;
        RECT 9.76 6.971 12.16 6.973 ;
  LAYER M2 ;
        RECT 9.76 6.887 12.16 6.889 ;
  LAYER M2 ;
        RECT 9.76 6.803 12.16 6.805 ;
  LAYER M2 ;
        RECT 9.76 6.719 12.16 6.721 ;
  LAYER M2 ;
        RECT 9.76 6.635 12.16 6.637 ;
  LAYER M2 ;
        RECT 9.76 6.551 12.16 6.553 ;
  LAYER M2 ;
        RECT 9.76 6.467 12.16 6.469 ;
  LAYER M2 ;
        RECT 9.76 6.383 12.16 6.385 ;
  LAYER M2 ;
        RECT 9.76 6.2995 12.16 6.3015 ;
  LAYER M2 ;
        RECT 9.76 6.215 12.16 6.217 ;
  LAYER M2 ;
        RECT 9.76 6.131 12.16 6.133 ;
  LAYER M2 ;
        RECT 9.76 6.047 12.16 6.049 ;
  LAYER M2 ;
        RECT 9.76 5.963 12.16 5.965 ;
  LAYER M2 ;
        RECT 9.76 5.879 12.16 5.881 ;
  LAYER M2 ;
        RECT 9.76 5.795 12.16 5.797 ;
  LAYER M2 ;
        RECT 9.76 5.711 12.16 5.713 ;
  LAYER M2 ;
        RECT 9.76 5.627 12.16 5.629 ;
  LAYER M2 ;
        RECT 9.76 5.543 12.16 5.545 ;
  LAYER M2 ;
        RECT 9.76 5.459 12.16 5.461 ;
  LAYER M2 ;
        RECT 9.76 5.375 12.16 5.377 ;
  LAYER M2 ;
        RECT 9.76 5.291 12.16 5.293 ;
  LAYER M2 ;
        RECT 9.76 5.207 12.16 5.209 ;
  LAYER M2 ;
        RECT 9.76 5.123 12.16 5.125 ;
  LAYER M2 ;
        RECT 9.76 5.039 12.16 5.041 ;
  LAYER M2 ;
        RECT 9.76 4.955 12.16 4.957 ;
  LAYER M1 ;
        RECT 9.744 1.896 9.776 4.404 ;
  LAYER M1 ;
        RECT 9.808 1.896 9.84 4.404 ;
  LAYER M1 ;
        RECT 9.872 1.896 9.904 4.404 ;
  LAYER M1 ;
        RECT 9.936 1.896 9.968 4.404 ;
  LAYER M1 ;
        RECT 10 1.896 10.032 4.404 ;
  LAYER M1 ;
        RECT 10.064 1.896 10.096 4.404 ;
  LAYER M1 ;
        RECT 10.128 1.896 10.16 4.404 ;
  LAYER M1 ;
        RECT 10.192 1.896 10.224 4.404 ;
  LAYER M1 ;
        RECT 10.256 1.896 10.288 4.404 ;
  LAYER M1 ;
        RECT 10.32 1.896 10.352 4.404 ;
  LAYER M1 ;
        RECT 10.384 1.896 10.416 4.404 ;
  LAYER M1 ;
        RECT 10.448 1.896 10.48 4.404 ;
  LAYER M1 ;
        RECT 10.512 1.896 10.544 4.404 ;
  LAYER M1 ;
        RECT 10.576 1.896 10.608 4.404 ;
  LAYER M1 ;
        RECT 10.64 1.896 10.672 4.404 ;
  LAYER M1 ;
        RECT 10.704 1.896 10.736 4.404 ;
  LAYER M1 ;
        RECT 10.768 1.896 10.8 4.404 ;
  LAYER M1 ;
        RECT 10.832 1.896 10.864 4.404 ;
  LAYER M1 ;
        RECT 10.896 1.896 10.928 4.404 ;
  LAYER M1 ;
        RECT 10.96 1.896 10.992 4.404 ;
  LAYER M1 ;
        RECT 11.024 1.896 11.056 4.404 ;
  LAYER M1 ;
        RECT 11.088 1.896 11.12 4.404 ;
  LAYER M1 ;
        RECT 11.152 1.896 11.184 4.404 ;
  LAYER M1 ;
        RECT 11.216 1.896 11.248 4.404 ;
  LAYER M1 ;
        RECT 11.28 1.896 11.312 4.404 ;
  LAYER M1 ;
        RECT 11.344 1.896 11.376 4.404 ;
  LAYER M1 ;
        RECT 11.408 1.896 11.44 4.404 ;
  LAYER M1 ;
        RECT 11.472 1.896 11.504 4.404 ;
  LAYER M1 ;
        RECT 11.536 1.896 11.568 4.404 ;
  LAYER M1 ;
        RECT 11.6 1.896 11.632 4.404 ;
  LAYER M1 ;
        RECT 11.664 1.896 11.696 4.404 ;
  LAYER M1 ;
        RECT 11.728 1.896 11.76 4.404 ;
  LAYER M1 ;
        RECT 11.792 1.896 11.824 4.404 ;
  LAYER M1 ;
        RECT 11.856 1.896 11.888 4.404 ;
  LAYER M1 ;
        RECT 11.92 1.896 11.952 4.404 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 4.404 ;
  LAYER M1 ;
        RECT 12.048 1.896 12.08 4.404 ;
  LAYER M2 ;
        RECT 9.724 4.288 12.196 4.32 ;
  LAYER M2 ;
        RECT 9.724 4.224 12.196 4.256 ;
  LAYER M2 ;
        RECT 9.724 4.16 12.196 4.192 ;
  LAYER M2 ;
        RECT 9.724 4.096 12.196 4.128 ;
  LAYER M2 ;
        RECT 9.724 4.032 12.196 4.064 ;
  LAYER M2 ;
        RECT 9.724 3.968 12.196 4 ;
  LAYER M2 ;
        RECT 9.724 3.904 12.196 3.936 ;
  LAYER M2 ;
        RECT 9.724 3.84 12.196 3.872 ;
  LAYER M2 ;
        RECT 9.724 3.776 12.196 3.808 ;
  LAYER M2 ;
        RECT 9.724 3.712 12.196 3.744 ;
  LAYER M2 ;
        RECT 9.724 3.648 12.196 3.68 ;
  LAYER M2 ;
        RECT 9.724 3.584 12.196 3.616 ;
  LAYER M2 ;
        RECT 9.724 3.52 12.196 3.552 ;
  LAYER M2 ;
        RECT 9.724 3.456 12.196 3.488 ;
  LAYER M2 ;
        RECT 9.724 3.392 12.196 3.424 ;
  LAYER M2 ;
        RECT 9.724 3.328 12.196 3.36 ;
  LAYER M2 ;
        RECT 9.724 3.264 12.196 3.296 ;
  LAYER M2 ;
        RECT 9.724 3.2 12.196 3.232 ;
  LAYER M2 ;
        RECT 9.724 3.136 12.196 3.168 ;
  LAYER M2 ;
        RECT 9.724 3.072 12.196 3.104 ;
  LAYER M2 ;
        RECT 9.724 3.008 12.196 3.04 ;
  LAYER M2 ;
        RECT 9.724 2.944 12.196 2.976 ;
  LAYER M2 ;
        RECT 9.724 2.88 12.196 2.912 ;
  LAYER M2 ;
        RECT 9.724 2.816 12.196 2.848 ;
  LAYER M2 ;
        RECT 9.724 2.752 12.196 2.784 ;
  LAYER M2 ;
        RECT 9.724 2.688 12.196 2.72 ;
  LAYER M2 ;
        RECT 9.724 2.624 12.196 2.656 ;
  LAYER M2 ;
        RECT 9.724 2.56 12.196 2.592 ;
  LAYER M2 ;
        RECT 9.724 2.496 12.196 2.528 ;
  LAYER M2 ;
        RECT 9.724 2.432 12.196 2.464 ;
  LAYER M2 ;
        RECT 9.724 2.368 12.196 2.4 ;
  LAYER M2 ;
        RECT 9.724 2.304 12.196 2.336 ;
  LAYER M2 ;
        RECT 9.724 2.24 12.196 2.272 ;
  LAYER M2 ;
        RECT 9.724 2.176 12.196 2.208 ;
  LAYER M2 ;
        RECT 9.724 2.112 12.196 2.144 ;
  LAYER M2 ;
        RECT 9.724 2.048 12.196 2.08 ;
  LAYER M3 ;
        RECT 9.744 1.896 9.776 4.404 ;
  LAYER M3 ;
        RECT 9.808 1.896 9.84 4.404 ;
  LAYER M3 ;
        RECT 9.872 1.896 9.904 4.404 ;
  LAYER M3 ;
        RECT 9.936 1.896 9.968 4.404 ;
  LAYER M3 ;
        RECT 10 1.896 10.032 4.404 ;
  LAYER M3 ;
        RECT 10.064 1.896 10.096 4.404 ;
  LAYER M3 ;
        RECT 10.128 1.896 10.16 4.404 ;
  LAYER M3 ;
        RECT 10.192 1.896 10.224 4.404 ;
  LAYER M3 ;
        RECT 10.256 1.896 10.288 4.404 ;
  LAYER M3 ;
        RECT 10.32 1.896 10.352 4.404 ;
  LAYER M3 ;
        RECT 10.384 1.896 10.416 4.404 ;
  LAYER M3 ;
        RECT 10.448 1.896 10.48 4.404 ;
  LAYER M3 ;
        RECT 10.512 1.896 10.544 4.404 ;
  LAYER M3 ;
        RECT 10.576 1.896 10.608 4.404 ;
  LAYER M3 ;
        RECT 10.64 1.896 10.672 4.404 ;
  LAYER M3 ;
        RECT 10.704 1.896 10.736 4.404 ;
  LAYER M3 ;
        RECT 10.768 1.896 10.8 4.404 ;
  LAYER M3 ;
        RECT 10.832 1.896 10.864 4.404 ;
  LAYER M3 ;
        RECT 10.896 1.896 10.928 4.404 ;
  LAYER M3 ;
        RECT 10.96 1.896 10.992 4.404 ;
  LAYER M3 ;
        RECT 11.024 1.896 11.056 4.404 ;
  LAYER M3 ;
        RECT 11.088 1.896 11.12 4.404 ;
  LAYER M3 ;
        RECT 11.152 1.896 11.184 4.404 ;
  LAYER M3 ;
        RECT 11.216 1.896 11.248 4.404 ;
  LAYER M3 ;
        RECT 11.28 1.896 11.312 4.404 ;
  LAYER M3 ;
        RECT 11.344 1.896 11.376 4.404 ;
  LAYER M3 ;
        RECT 11.408 1.896 11.44 4.404 ;
  LAYER M3 ;
        RECT 11.472 1.896 11.504 4.404 ;
  LAYER M3 ;
        RECT 11.536 1.896 11.568 4.404 ;
  LAYER M3 ;
        RECT 11.6 1.896 11.632 4.404 ;
  LAYER M3 ;
        RECT 11.664 1.896 11.696 4.404 ;
  LAYER M3 ;
        RECT 11.728 1.896 11.76 4.404 ;
  LAYER M3 ;
        RECT 11.792 1.896 11.824 4.404 ;
  LAYER M3 ;
        RECT 11.856 1.896 11.888 4.404 ;
  LAYER M3 ;
        RECT 11.92 1.896 11.952 4.404 ;
  LAYER M3 ;
        RECT 11.984 1.896 12.016 4.404 ;
  LAYER M3 ;
        RECT 12.048 1.896 12.08 4.404 ;
  LAYER M3 ;
        RECT 12.144 1.896 12.176 4.404 ;
  LAYER M1 ;
        RECT 9.759 1.932 9.761 4.368 ;
  LAYER M1 ;
        RECT 9.839 1.932 9.841 4.368 ;
  LAYER M1 ;
        RECT 9.919 1.932 9.921 4.368 ;
  LAYER M1 ;
        RECT 9.999 1.932 10.001 4.368 ;
  LAYER M1 ;
        RECT 10.079 1.932 10.081 4.368 ;
  LAYER M1 ;
        RECT 10.159 1.932 10.161 4.368 ;
  LAYER M1 ;
        RECT 10.239 1.932 10.241 4.368 ;
  LAYER M1 ;
        RECT 10.319 1.932 10.321 4.368 ;
  LAYER M1 ;
        RECT 10.399 1.932 10.401 4.368 ;
  LAYER M1 ;
        RECT 10.479 1.932 10.481 4.368 ;
  LAYER M1 ;
        RECT 10.559 1.932 10.561 4.368 ;
  LAYER M1 ;
        RECT 10.639 1.932 10.641 4.368 ;
  LAYER M1 ;
        RECT 10.719 1.932 10.721 4.368 ;
  LAYER M1 ;
        RECT 10.799 1.932 10.801 4.368 ;
  LAYER M1 ;
        RECT 10.879 1.932 10.881 4.368 ;
  LAYER M1 ;
        RECT 10.959 1.932 10.961 4.368 ;
  LAYER M1 ;
        RECT 11.039 1.932 11.041 4.368 ;
  LAYER M1 ;
        RECT 11.119 1.932 11.121 4.368 ;
  LAYER M1 ;
        RECT 11.199 1.932 11.201 4.368 ;
  LAYER M1 ;
        RECT 11.279 1.932 11.281 4.368 ;
  LAYER M1 ;
        RECT 11.359 1.932 11.361 4.368 ;
  LAYER M1 ;
        RECT 11.439 1.932 11.441 4.368 ;
  LAYER M1 ;
        RECT 11.519 1.932 11.521 4.368 ;
  LAYER M1 ;
        RECT 11.599 1.932 11.601 4.368 ;
  LAYER M1 ;
        RECT 11.679 1.932 11.681 4.368 ;
  LAYER M1 ;
        RECT 11.759 1.932 11.761 4.368 ;
  LAYER M1 ;
        RECT 11.839 1.932 11.841 4.368 ;
  LAYER M1 ;
        RECT 11.919 1.932 11.921 4.368 ;
  LAYER M1 ;
        RECT 11.999 1.932 12.001 4.368 ;
  LAYER M1 ;
        RECT 12.079 1.932 12.081 4.368 ;
  LAYER M2 ;
        RECT 9.76 4.367 12.16 4.369 ;
  LAYER M2 ;
        RECT 9.76 4.283 12.16 4.285 ;
  LAYER M2 ;
        RECT 9.76 4.199 12.16 4.201 ;
  LAYER M2 ;
        RECT 9.76 4.115 12.16 4.117 ;
  LAYER M2 ;
        RECT 9.76 4.031 12.16 4.033 ;
  LAYER M2 ;
        RECT 9.76 3.947 12.16 3.949 ;
  LAYER M2 ;
        RECT 9.76 3.863 12.16 3.865 ;
  LAYER M2 ;
        RECT 9.76 3.779 12.16 3.781 ;
  LAYER M2 ;
        RECT 9.76 3.695 12.16 3.697 ;
  LAYER M2 ;
        RECT 9.76 3.611 12.16 3.613 ;
  LAYER M2 ;
        RECT 9.76 3.527 12.16 3.529 ;
  LAYER M2 ;
        RECT 9.76 3.443 12.16 3.445 ;
  LAYER M2 ;
        RECT 9.76 3.3595 12.16 3.3615 ;
  LAYER M2 ;
        RECT 9.76 3.275 12.16 3.277 ;
  LAYER M2 ;
        RECT 9.76 3.191 12.16 3.193 ;
  LAYER M2 ;
        RECT 9.76 3.107 12.16 3.109 ;
  LAYER M2 ;
        RECT 9.76 3.023 12.16 3.025 ;
  LAYER M2 ;
        RECT 9.76 2.939 12.16 2.941 ;
  LAYER M2 ;
        RECT 9.76 2.855 12.16 2.857 ;
  LAYER M2 ;
        RECT 9.76 2.771 12.16 2.773 ;
  LAYER M2 ;
        RECT 9.76 2.687 12.16 2.689 ;
  LAYER M2 ;
        RECT 9.76 2.603 12.16 2.605 ;
  LAYER M2 ;
        RECT 9.76 2.519 12.16 2.521 ;
  LAYER M2 ;
        RECT 9.76 2.435 12.16 2.437 ;
  LAYER M2 ;
        RECT 9.76 2.351 12.16 2.353 ;
  LAYER M2 ;
        RECT 9.76 2.267 12.16 2.269 ;
  LAYER M2 ;
        RECT 9.76 2.183 12.16 2.185 ;
  LAYER M2 ;
        RECT 9.76 2.099 12.16 2.101 ;
  LAYER M2 ;
        RECT 9.76 2.015 12.16 2.017 ;
  LAYER M1 ;
        RECT 12.624 13.656 12.656 16.164 ;
  LAYER M1 ;
        RECT 12.688 13.656 12.72 16.164 ;
  LAYER M1 ;
        RECT 12.752 13.656 12.784 16.164 ;
  LAYER M1 ;
        RECT 12.816 13.656 12.848 16.164 ;
  LAYER M1 ;
        RECT 12.88 13.656 12.912 16.164 ;
  LAYER M1 ;
        RECT 12.944 13.656 12.976 16.164 ;
  LAYER M1 ;
        RECT 13.008 13.656 13.04 16.164 ;
  LAYER M1 ;
        RECT 13.072 13.656 13.104 16.164 ;
  LAYER M1 ;
        RECT 13.136 13.656 13.168 16.164 ;
  LAYER M1 ;
        RECT 13.2 13.656 13.232 16.164 ;
  LAYER M1 ;
        RECT 13.264 13.656 13.296 16.164 ;
  LAYER M1 ;
        RECT 13.328 13.656 13.36 16.164 ;
  LAYER M1 ;
        RECT 13.392 13.656 13.424 16.164 ;
  LAYER M1 ;
        RECT 13.456 13.656 13.488 16.164 ;
  LAYER M1 ;
        RECT 13.52 13.656 13.552 16.164 ;
  LAYER M1 ;
        RECT 13.584 13.656 13.616 16.164 ;
  LAYER M1 ;
        RECT 13.648 13.656 13.68 16.164 ;
  LAYER M1 ;
        RECT 13.712 13.656 13.744 16.164 ;
  LAYER M1 ;
        RECT 13.776 13.656 13.808 16.164 ;
  LAYER M1 ;
        RECT 13.84 13.656 13.872 16.164 ;
  LAYER M1 ;
        RECT 13.904 13.656 13.936 16.164 ;
  LAYER M1 ;
        RECT 13.968 13.656 14 16.164 ;
  LAYER M1 ;
        RECT 14.032 13.656 14.064 16.164 ;
  LAYER M1 ;
        RECT 14.096 13.656 14.128 16.164 ;
  LAYER M1 ;
        RECT 14.16 13.656 14.192 16.164 ;
  LAYER M1 ;
        RECT 14.224 13.656 14.256 16.164 ;
  LAYER M1 ;
        RECT 14.288 13.656 14.32 16.164 ;
  LAYER M1 ;
        RECT 14.352 13.656 14.384 16.164 ;
  LAYER M1 ;
        RECT 14.416 13.656 14.448 16.164 ;
  LAYER M1 ;
        RECT 14.48 13.656 14.512 16.164 ;
  LAYER M1 ;
        RECT 14.544 13.656 14.576 16.164 ;
  LAYER M1 ;
        RECT 14.608 13.656 14.64 16.164 ;
  LAYER M1 ;
        RECT 14.672 13.656 14.704 16.164 ;
  LAYER M1 ;
        RECT 14.736 13.656 14.768 16.164 ;
  LAYER M1 ;
        RECT 14.8 13.656 14.832 16.164 ;
  LAYER M1 ;
        RECT 14.864 13.656 14.896 16.164 ;
  LAYER M1 ;
        RECT 14.928 13.656 14.96 16.164 ;
  LAYER M2 ;
        RECT 12.604 16.048 15.076 16.08 ;
  LAYER M2 ;
        RECT 12.604 15.984 15.076 16.016 ;
  LAYER M2 ;
        RECT 12.604 15.92 15.076 15.952 ;
  LAYER M2 ;
        RECT 12.604 15.856 15.076 15.888 ;
  LAYER M2 ;
        RECT 12.604 15.792 15.076 15.824 ;
  LAYER M2 ;
        RECT 12.604 15.728 15.076 15.76 ;
  LAYER M2 ;
        RECT 12.604 15.664 15.076 15.696 ;
  LAYER M2 ;
        RECT 12.604 15.6 15.076 15.632 ;
  LAYER M2 ;
        RECT 12.604 15.536 15.076 15.568 ;
  LAYER M2 ;
        RECT 12.604 15.472 15.076 15.504 ;
  LAYER M2 ;
        RECT 12.604 15.408 15.076 15.44 ;
  LAYER M2 ;
        RECT 12.604 15.344 15.076 15.376 ;
  LAYER M2 ;
        RECT 12.604 15.28 15.076 15.312 ;
  LAYER M2 ;
        RECT 12.604 15.216 15.076 15.248 ;
  LAYER M2 ;
        RECT 12.604 15.152 15.076 15.184 ;
  LAYER M2 ;
        RECT 12.604 15.088 15.076 15.12 ;
  LAYER M2 ;
        RECT 12.604 15.024 15.076 15.056 ;
  LAYER M2 ;
        RECT 12.604 14.96 15.076 14.992 ;
  LAYER M2 ;
        RECT 12.604 14.896 15.076 14.928 ;
  LAYER M2 ;
        RECT 12.604 14.832 15.076 14.864 ;
  LAYER M2 ;
        RECT 12.604 14.768 15.076 14.8 ;
  LAYER M2 ;
        RECT 12.604 14.704 15.076 14.736 ;
  LAYER M2 ;
        RECT 12.604 14.64 15.076 14.672 ;
  LAYER M2 ;
        RECT 12.604 14.576 15.076 14.608 ;
  LAYER M2 ;
        RECT 12.604 14.512 15.076 14.544 ;
  LAYER M2 ;
        RECT 12.604 14.448 15.076 14.48 ;
  LAYER M2 ;
        RECT 12.604 14.384 15.076 14.416 ;
  LAYER M2 ;
        RECT 12.604 14.32 15.076 14.352 ;
  LAYER M2 ;
        RECT 12.604 14.256 15.076 14.288 ;
  LAYER M2 ;
        RECT 12.604 14.192 15.076 14.224 ;
  LAYER M2 ;
        RECT 12.604 14.128 15.076 14.16 ;
  LAYER M2 ;
        RECT 12.604 14.064 15.076 14.096 ;
  LAYER M2 ;
        RECT 12.604 14 15.076 14.032 ;
  LAYER M2 ;
        RECT 12.604 13.936 15.076 13.968 ;
  LAYER M2 ;
        RECT 12.604 13.872 15.076 13.904 ;
  LAYER M2 ;
        RECT 12.604 13.808 15.076 13.84 ;
  LAYER M3 ;
        RECT 12.624 13.656 12.656 16.164 ;
  LAYER M3 ;
        RECT 12.688 13.656 12.72 16.164 ;
  LAYER M3 ;
        RECT 12.752 13.656 12.784 16.164 ;
  LAYER M3 ;
        RECT 12.816 13.656 12.848 16.164 ;
  LAYER M3 ;
        RECT 12.88 13.656 12.912 16.164 ;
  LAYER M3 ;
        RECT 12.944 13.656 12.976 16.164 ;
  LAYER M3 ;
        RECT 13.008 13.656 13.04 16.164 ;
  LAYER M3 ;
        RECT 13.072 13.656 13.104 16.164 ;
  LAYER M3 ;
        RECT 13.136 13.656 13.168 16.164 ;
  LAYER M3 ;
        RECT 13.2 13.656 13.232 16.164 ;
  LAYER M3 ;
        RECT 13.264 13.656 13.296 16.164 ;
  LAYER M3 ;
        RECT 13.328 13.656 13.36 16.164 ;
  LAYER M3 ;
        RECT 13.392 13.656 13.424 16.164 ;
  LAYER M3 ;
        RECT 13.456 13.656 13.488 16.164 ;
  LAYER M3 ;
        RECT 13.52 13.656 13.552 16.164 ;
  LAYER M3 ;
        RECT 13.584 13.656 13.616 16.164 ;
  LAYER M3 ;
        RECT 13.648 13.656 13.68 16.164 ;
  LAYER M3 ;
        RECT 13.712 13.656 13.744 16.164 ;
  LAYER M3 ;
        RECT 13.776 13.656 13.808 16.164 ;
  LAYER M3 ;
        RECT 13.84 13.656 13.872 16.164 ;
  LAYER M3 ;
        RECT 13.904 13.656 13.936 16.164 ;
  LAYER M3 ;
        RECT 13.968 13.656 14 16.164 ;
  LAYER M3 ;
        RECT 14.032 13.656 14.064 16.164 ;
  LAYER M3 ;
        RECT 14.096 13.656 14.128 16.164 ;
  LAYER M3 ;
        RECT 14.16 13.656 14.192 16.164 ;
  LAYER M3 ;
        RECT 14.224 13.656 14.256 16.164 ;
  LAYER M3 ;
        RECT 14.288 13.656 14.32 16.164 ;
  LAYER M3 ;
        RECT 14.352 13.656 14.384 16.164 ;
  LAYER M3 ;
        RECT 14.416 13.656 14.448 16.164 ;
  LAYER M3 ;
        RECT 14.48 13.656 14.512 16.164 ;
  LAYER M3 ;
        RECT 14.544 13.656 14.576 16.164 ;
  LAYER M3 ;
        RECT 14.608 13.656 14.64 16.164 ;
  LAYER M3 ;
        RECT 14.672 13.656 14.704 16.164 ;
  LAYER M3 ;
        RECT 14.736 13.656 14.768 16.164 ;
  LAYER M3 ;
        RECT 14.8 13.656 14.832 16.164 ;
  LAYER M3 ;
        RECT 14.864 13.656 14.896 16.164 ;
  LAYER M3 ;
        RECT 14.928 13.656 14.96 16.164 ;
  LAYER M3 ;
        RECT 15.024 13.656 15.056 16.164 ;
  LAYER M1 ;
        RECT 12.639 13.692 12.641 16.128 ;
  LAYER M1 ;
        RECT 12.719 13.692 12.721 16.128 ;
  LAYER M1 ;
        RECT 12.799 13.692 12.801 16.128 ;
  LAYER M1 ;
        RECT 12.879 13.692 12.881 16.128 ;
  LAYER M1 ;
        RECT 12.959 13.692 12.961 16.128 ;
  LAYER M1 ;
        RECT 13.039 13.692 13.041 16.128 ;
  LAYER M1 ;
        RECT 13.119 13.692 13.121 16.128 ;
  LAYER M1 ;
        RECT 13.199 13.692 13.201 16.128 ;
  LAYER M1 ;
        RECT 13.279 13.692 13.281 16.128 ;
  LAYER M1 ;
        RECT 13.359 13.692 13.361 16.128 ;
  LAYER M1 ;
        RECT 13.439 13.692 13.441 16.128 ;
  LAYER M1 ;
        RECT 13.519 13.692 13.521 16.128 ;
  LAYER M1 ;
        RECT 13.599 13.692 13.601 16.128 ;
  LAYER M1 ;
        RECT 13.679 13.692 13.681 16.128 ;
  LAYER M1 ;
        RECT 13.759 13.692 13.761 16.128 ;
  LAYER M1 ;
        RECT 13.839 13.692 13.841 16.128 ;
  LAYER M1 ;
        RECT 13.919 13.692 13.921 16.128 ;
  LAYER M1 ;
        RECT 13.999 13.692 14.001 16.128 ;
  LAYER M1 ;
        RECT 14.079 13.692 14.081 16.128 ;
  LAYER M1 ;
        RECT 14.159 13.692 14.161 16.128 ;
  LAYER M1 ;
        RECT 14.239 13.692 14.241 16.128 ;
  LAYER M1 ;
        RECT 14.319 13.692 14.321 16.128 ;
  LAYER M1 ;
        RECT 14.399 13.692 14.401 16.128 ;
  LAYER M1 ;
        RECT 14.479 13.692 14.481 16.128 ;
  LAYER M1 ;
        RECT 14.559 13.692 14.561 16.128 ;
  LAYER M1 ;
        RECT 14.639 13.692 14.641 16.128 ;
  LAYER M1 ;
        RECT 14.719 13.692 14.721 16.128 ;
  LAYER M1 ;
        RECT 14.799 13.692 14.801 16.128 ;
  LAYER M1 ;
        RECT 14.879 13.692 14.881 16.128 ;
  LAYER M1 ;
        RECT 14.959 13.692 14.961 16.128 ;
  LAYER M2 ;
        RECT 12.64 16.127 15.04 16.129 ;
  LAYER M2 ;
        RECT 12.64 16.043 15.04 16.045 ;
  LAYER M2 ;
        RECT 12.64 15.959 15.04 15.961 ;
  LAYER M2 ;
        RECT 12.64 15.875 15.04 15.877 ;
  LAYER M2 ;
        RECT 12.64 15.791 15.04 15.793 ;
  LAYER M2 ;
        RECT 12.64 15.707 15.04 15.709 ;
  LAYER M2 ;
        RECT 12.64 15.623 15.04 15.625 ;
  LAYER M2 ;
        RECT 12.64 15.539 15.04 15.541 ;
  LAYER M2 ;
        RECT 12.64 15.455 15.04 15.457 ;
  LAYER M2 ;
        RECT 12.64 15.371 15.04 15.373 ;
  LAYER M2 ;
        RECT 12.64 15.287 15.04 15.289 ;
  LAYER M2 ;
        RECT 12.64 15.203 15.04 15.205 ;
  LAYER M2 ;
        RECT 12.64 15.1195 15.04 15.1215 ;
  LAYER M2 ;
        RECT 12.64 15.035 15.04 15.037 ;
  LAYER M2 ;
        RECT 12.64 14.951 15.04 14.953 ;
  LAYER M2 ;
        RECT 12.64 14.867 15.04 14.869 ;
  LAYER M2 ;
        RECT 12.64 14.783 15.04 14.785 ;
  LAYER M2 ;
        RECT 12.64 14.699 15.04 14.701 ;
  LAYER M2 ;
        RECT 12.64 14.615 15.04 14.617 ;
  LAYER M2 ;
        RECT 12.64 14.531 15.04 14.533 ;
  LAYER M2 ;
        RECT 12.64 14.447 15.04 14.449 ;
  LAYER M2 ;
        RECT 12.64 14.363 15.04 14.365 ;
  LAYER M2 ;
        RECT 12.64 14.279 15.04 14.281 ;
  LAYER M2 ;
        RECT 12.64 14.195 15.04 14.197 ;
  LAYER M2 ;
        RECT 12.64 14.111 15.04 14.113 ;
  LAYER M2 ;
        RECT 12.64 14.027 15.04 14.029 ;
  LAYER M2 ;
        RECT 12.64 13.943 15.04 13.945 ;
  LAYER M2 ;
        RECT 12.64 13.859 15.04 13.861 ;
  LAYER M2 ;
        RECT 12.64 13.775 15.04 13.777 ;
  LAYER M1 ;
        RECT 12.624 10.716 12.656 13.224 ;
  LAYER M1 ;
        RECT 12.688 10.716 12.72 13.224 ;
  LAYER M1 ;
        RECT 12.752 10.716 12.784 13.224 ;
  LAYER M1 ;
        RECT 12.816 10.716 12.848 13.224 ;
  LAYER M1 ;
        RECT 12.88 10.716 12.912 13.224 ;
  LAYER M1 ;
        RECT 12.944 10.716 12.976 13.224 ;
  LAYER M1 ;
        RECT 13.008 10.716 13.04 13.224 ;
  LAYER M1 ;
        RECT 13.072 10.716 13.104 13.224 ;
  LAYER M1 ;
        RECT 13.136 10.716 13.168 13.224 ;
  LAYER M1 ;
        RECT 13.2 10.716 13.232 13.224 ;
  LAYER M1 ;
        RECT 13.264 10.716 13.296 13.224 ;
  LAYER M1 ;
        RECT 13.328 10.716 13.36 13.224 ;
  LAYER M1 ;
        RECT 13.392 10.716 13.424 13.224 ;
  LAYER M1 ;
        RECT 13.456 10.716 13.488 13.224 ;
  LAYER M1 ;
        RECT 13.52 10.716 13.552 13.224 ;
  LAYER M1 ;
        RECT 13.584 10.716 13.616 13.224 ;
  LAYER M1 ;
        RECT 13.648 10.716 13.68 13.224 ;
  LAYER M1 ;
        RECT 13.712 10.716 13.744 13.224 ;
  LAYER M1 ;
        RECT 13.776 10.716 13.808 13.224 ;
  LAYER M1 ;
        RECT 13.84 10.716 13.872 13.224 ;
  LAYER M1 ;
        RECT 13.904 10.716 13.936 13.224 ;
  LAYER M1 ;
        RECT 13.968 10.716 14 13.224 ;
  LAYER M1 ;
        RECT 14.032 10.716 14.064 13.224 ;
  LAYER M1 ;
        RECT 14.096 10.716 14.128 13.224 ;
  LAYER M1 ;
        RECT 14.16 10.716 14.192 13.224 ;
  LAYER M1 ;
        RECT 14.224 10.716 14.256 13.224 ;
  LAYER M1 ;
        RECT 14.288 10.716 14.32 13.224 ;
  LAYER M1 ;
        RECT 14.352 10.716 14.384 13.224 ;
  LAYER M1 ;
        RECT 14.416 10.716 14.448 13.224 ;
  LAYER M1 ;
        RECT 14.48 10.716 14.512 13.224 ;
  LAYER M1 ;
        RECT 14.544 10.716 14.576 13.224 ;
  LAYER M1 ;
        RECT 14.608 10.716 14.64 13.224 ;
  LAYER M1 ;
        RECT 14.672 10.716 14.704 13.224 ;
  LAYER M1 ;
        RECT 14.736 10.716 14.768 13.224 ;
  LAYER M1 ;
        RECT 14.8 10.716 14.832 13.224 ;
  LAYER M1 ;
        RECT 14.864 10.716 14.896 13.224 ;
  LAYER M1 ;
        RECT 14.928 10.716 14.96 13.224 ;
  LAYER M2 ;
        RECT 12.604 13.108 15.076 13.14 ;
  LAYER M2 ;
        RECT 12.604 13.044 15.076 13.076 ;
  LAYER M2 ;
        RECT 12.604 12.98 15.076 13.012 ;
  LAYER M2 ;
        RECT 12.604 12.916 15.076 12.948 ;
  LAYER M2 ;
        RECT 12.604 12.852 15.076 12.884 ;
  LAYER M2 ;
        RECT 12.604 12.788 15.076 12.82 ;
  LAYER M2 ;
        RECT 12.604 12.724 15.076 12.756 ;
  LAYER M2 ;
        RECT 12.604 12.66 15.076 12.692 ;
  LAYER M2 ;
        RECT 12.604 12.596 15.076 12.628 ;
  LAYER M2 ;
        RECT 12.604 12.532 15.076 12.564 ;
  LAYER M2 ;
        RECT 12.604 12.468 15.076 12.5 ;
  LAYER M2 ;
        RECT 12.604 12.404 15.076 12.436 ;
  LAYER M2 ;
        RECT 12.604 12.34 15.076 12.372 ;
  LAYER M2 ;
        RECT 12.604 12.276 15.076 12.308 ;
  LAYER M2 ;
        RECT 12.604 12.212 15.076 12.244 ;
  LAYER M2 ;
        RECT 12.604 12.148 15.076 12.18 ;
  LAYER M2 ;
        RECT 12.604 12.084 15.076 12.116 ;
  LAYER M2 ;
        RECT 12.604 12.02 15.076 12.052 ;
  LAYER M2 ;
        RECT 12.604 11.956 15.076 11.988 ;
  LAYER M2 ;
        RECT 12.604 11.892 15.076 11.924 ;
  LAYER M2 ;
        RECT 12.604 11.828 15.076 11.86 ;
  LAYER M2 ;
        RECT 12.604 11.764 15.076 11.796 ;
  LAYER M2 ;
        RECT 12.604 11.7 15.076 11.732 ;
  LAYER M2 ;
        RECT 12.604 11.636 15.076 11.668 ;
  LAYER M2 ;
        RECT 12.604 11.572 15.076 11.604 ;
  LAYER M2 ;
        RECT 12.604 11.508 15.076 11.54 ;
  LAYER M2 ;
        RECT 12.604 11.444 15.076 11.476 ;
  LAYER M2 ;
        RECT 12.604 11.38 15.076 11.412 ;
  LAYER M2 ;
        RECT 12.604 11.316 15.076 11.348 ;
  LAYER M2 ;
        RECT 12.604 11.252 15.076 11.284 ;
  LAYER M2 ;
        RECT 12.604 11.188 15.076 11.22 ;
  LAYER M2 ;
        RECT 12.604 11.124 15.076 11.156 ;
  LAYER M2 ;
        RECT 12.604 11.06 15.076 11.092 ;
  LAYER M2 ;
        RECT 12.604 10.996 15.076 11.028 ;
  LAYER M2 ;
        RECT 12.604 10.932 15.076 10.964 ;
  LAYER M2 ;
        RECT 12.604 10.868 15.076 10.9 ;
  LAYER M3 ;
        RECT 12.624 10.716 12.656 13.224 ;
  LAYER M3 ;
        RECT 12.688 10.716 12.72 13.224 ;
  LAYER M3 ;
        RECT 12.752 10.716 12.784 13.224 ;
  LAYER M3 ;
        RECT 12.816 10.716 12.848 13.224 ;
  LAYER M3 ;
        RECT 12.88 10.716 12.912 13.224 ;
  LAYER M3 ;
        RECT 12.944 10.716 12.976 13.224 ;
  LAYER M3 ;
        RECT 13.008 10.716 13.04 13.224 ;
  LAYER M3 ;
        RECT 13.072 10.716 13.104 13.224 ;
  LAYER M3 ;
        RECT 13.136 10.716 13.168 13.224 ;
  LAYER M3 ;
        RECT 13.2 10.716 13.232 13.224 ;
  LAYER M3 ;
        RECT 13.264 10.716 13.296 13.224 ;
  LAYER M3 ;
        RECT 13.328 10.716 13.36 13.224 ;
  LAYER M3 ;
        RECT 13.392 10.716 13.424 13.224 ;
  LAYER M3 ;
        RECT 13.456 10.716 13.488 13.224 ;
  LAYER M3 ;
        RECT 13.52 10.716 13.552 13.224 ;
  LAYER M3 ;
        RECT 13.584 10.716 13.616 13.224 ;
  LAYER M3 ;
        RECT 13.648 10.716 13.68 13.224 ;
  LAYER M3 ;
        RECT 13.712 10.716 13.744 13.224 ;
  LAYER M3 ;
        RECT 13.776 10.716 13.808 13.224 ;
  LAYER M3 ;
        RECT 13.84 10.716 13.872 13.224 ;
  LAYER M3 ;
        RECT 13.904 10.716 13.936 13.224 ;
  LAYER M3 ;
        RECT 13.968 10.716 14 13.224 ;
  LAYER M3 ;
        RECT 14.032 10.716 14.064 13.224 ;
  LAYER M3 ;
        RECT 14.096 10.716 14.128 13.224 ;
  LAYER M3 ;
        RECT 14.16 10.716 14.192 13.224 ;
  LAYER M3 ;
        RECT 14.224 10.716 14.256 13.224 ;
  LAYER M3 ;
        RECT 14.288 10.716 14.32 13.224 ;
  LAYER M3 ;
        RECT 14.352 10.716 14.384 13.224 ;
  LAYER M3 ;
        RECT 14.416 10.716 14.448 13.224 ;
  LAYER M3 ;
        RECT 14.48 10.716 14.512 13.224 ;
  LAYER M3 ;
        RECT 14.544 10.716 14.576 13.224 ;
  LAYER M3 ;
        RECT 14.608 10.716 14.64 13.224 ;
  LAYER M3 ;
        RECT 14.672 10.716 14.704 13.224 ;
  LAYER M3 ;
        RECT 14.736 10.716 14.768 13.224 ;
  LAYER M3 ;
        RECT 14.8 10.716 14.832 13.224 ;
  LAYER M3 ;
        RECT 14.864 10.716 14.896 13.224 ;
  LAYER M3 ;
        RECT 14.928 10.716 14.96 13.224 ;
  LAYER M3 ;
        RECT 15.024 10.716 15.056 13.224 ;
  LAYER M1 ;
        RECT 12.639 10.752 12.641 13.188 ;
  LAYER M1 ;
        RECT 12.719 10.752 12.721 13.188 ;
  LAYER M1 ;
        RECT 12.799 10.752 12.801 13.188 ;
  LAYER M1 ;
        RECT 12.879 10.752 12.881 13.188 ;
  LAYER M1 ;
        RECT 12.959 10.752 12.961 13.188 ;
  LAYER M1 ;
        RECT 13.039 10.752 13.041 13.188 ;
  LAYER M1 ;
        RECT 13.119 10.752 13.121 13.188 ;
  LAYER M1 ;
        RECT 13.199 10.752 13.201 13.188 ;
  LAYER M1 ;
        RECT 13.279 10.752 13.281 13.188 ;
  LAYER M1 ;
        RECT 13.359 10.752 13.361 13.188 ;
  LAYER M1 ;
        RECT 13.439 10.752 13.441 13.188 ;
  LAYER M1 ;
        RECT 13.519 10.752 13.521 13.188 ;
  LAYER M1 ;
        RECT 13.599 10.752 13.601 13.188 ;
  LAYER M1 ;
        RECT 13.679 10.752 13.681 13.188 ;
  LAYER M1 ;
        RECT 13.759 10.752 13.761 13.188 ;
  LAYER M1 ;
        RECT 13.839 10.752 13.841 13.188 ;
  LAYER M1 ;
        RECT 13.919 10.752 13.921 13.188 ;
  LAYER M1 ;
        RECT 13.999 10.752 14.001 13.188 ;
  LAYER M1 ;
        RECT 14.079 10.752 14.081 13.188 ;
  LAYER M1 ;
        RECT 14.159 10.752 14.161 13.188 ;
  LAYER M1 ;
        RECT 14.239 10.752 14.241 13.188 ;
  LAYER M1 ;
        RECT 14.319 10.752 14.321 13.188 ;
  LAYER M1 ;
        RECT 14.399 10.752 14.401 13.188 ;
  LAYER M1 ;
        RECT 14.479 10.752 14.481 13.188 ;
  LAYER M1 ;
        RECT 14.559 10.752 14.561 13.188 ;
  LAYER M1 ;
        RECT 14.639 10.752 14.641 13.188 ;
  LAYER M1 ;
        RECT 14.719 10.752 14.721 13.188 ;
  LAYER M1 ;
        RECT 14.799 10.752 14.801 13.188 ;
  LAYER M1 ;
        RECT 14.879 10.752 14.881 13.188 ;
  LAYER M1 ;
        RECT 14.959 10.752 14.961 13.188 ;
  LAYER M2 ;
        RECT 12.64 13.187 15.04 13.189 ;
  LAYER M2 ;
        RECT 12.64 13.103 15.04 13.105 ;
  LAYER M2 ;
        RECT 12.64 13.019 15.04 13.021 ;
  LAYER M2 ;
        RECT 12.64 12.935 15.04 12.937 ;
  LAYER M2 ;
        RECT 12.64 12.851 15.04 12.853 ;
  LAYER M2 ;
        RECT 12.64 12.767 15.04 12.769 ;
  LAYER M2 ;
        RECT 12.64 12.683 15.04 12.685 ;
  LAYER M2 ;
        RECT 12.64 12.599 15.04 12.601 ;
  LAYER M2 ;
        RECT 12.64 12.515 15.04 12.517 ;
  LAYER M2 ;
        RECT 12.64 12.431 15.04 12.433 ;
  LAYER M2 ;
        RECT 12.64 12.347 15.04 12.349 ;
  LAYER M2 ;
        RECT 12.64 12.263 15.04 12.265 ;
  LAYER M2 ;
        RECT 12.64 12.1795 15.04 12.1815 ;
  LAYER M2 ;
        RECT 12.64 12.095 15.04 12.097 ;
  LAYER M2 ;
        RECT 12.64 12.011 15.04 12.013 ;
  LAYER M2 ;
        RECT 12.64 11.927 15.04 11.929 ;
  LAYER M2 ;
        RECT 12.64 11.843 15.04 11.845 ;
  LAYER M2 ;
        RECT 12.64 11.759 15.04 11.761 ;
  LAYER M2 ;
        RECT 12.64 11.675 15.04 11.677 ;
  LAYER M2 ;
        RECT 12.64 11.591 15.04 11.593 ;
  LAYER M2 ;
        RECT 12.64 11.507 15.04 11.509 ;
  LAYER M2 ;
        RECT 12.64 11.423 15.04 11.425 ;
  LAYER M2 ;
        RECT 12.64 11.339 15.04 11.341 ;
  LAYER M2 ;
        RECT 12.64 11.255 15.04 11.257 ;
  LAYER M2 ;
        RECT 12.64 11.171 15.04 11.173 ;
  LAYER M2 ;
        RECT 12.64 11.087 15.04 11.089 ;
  LAYER M2 ;
        RECT 12.64 11.003 15.04 11.005 ;
  LAYER M2 ;
        RECT 12.64 10.919 15.04 10.921 ;
  LAYER M2 ;
        RECT 12.64 10.835 15.04 10.837 ;
  LAYER M1 ;
        RECT 12.624 7.776 12.656 10.284 ;
  LAYER M1 ;
        RECT 12.688 7.776 12.72 10.284 ;
  LAYER M1 ;
        RECT 12.752 7.776 12.784 10.284 ;
  LAYER M1 ;
        RECT 12.816 7.776 12.848 10.284 ;
  LAYER M1 ;
        RECT 12.88 7.776 12.912 10.284 ;
  LAYER M1 ;
        RECT 12.944 7.776 12.976 10.284 ;
  LAYER M1 ;
        RECT 13.008 7.776 13.04 10.284 ;
  LAYER M1 ;
        RECT 13.072 7.776 13.104 10.284 ;
  LAYER M1 ;
        RECT 13.136 7.776 13.168 10.284 ;
  LAYER M1 ;
        RECT 13.2 7.776 13.232 10.284 ;
  LAYER M1 ;
        RECT 13.264 7.776 13.296 10.284 ;
  LAYER M1 ;
        RECT 13.328 7.776 13.36 10.284 ;
  LAYER M1 ;
        RECT 13.392 7.776 13.424 10.284 ;
  LAYER M1 ;
        RECT 13.456 7.776 13.488 10.284 ;
  LAYER M1 ;
        RECT 13.52 7.776 13.552 10.284 ;
  LAYER M1 ;
        RECT 13.584 7.776 13.616 10.284 ;
  LAYER M1 ;
        RECT 13.648 7.776 13.68 10.284 ;
  LAYER M1 ;
        RECT 13.712 7.776 13.744 10.284 ;
  LAYER M1 ;
        RECT 13.776 7.776 13.808 10.284 ;
  LAYER M1 ;
        RECT 13.84 7.776 13.872 10.284 ;
  LAYER M1 ;
        RECT 13.904 7.776 13.936 10.284 ;
  LAYER M1 ;
        RECT 13.968 7.776 14 10.284 ;
  LAYER M1 ;
        RECT 14.032 7.776 14.064 10.284 ;
  LAYER M1 ;
        RECT 14.096 7.776 14.128 10.284 ;
  LAYER M1 ;
        RECT 14.16 7.776 14.192 10.284 ;
  LAYER M1 ;
        RECT 14.224 7.776 14.256 10.284 ;
  LAYER M1 ;
        RECT 14.288 7.776 14.32 10.284 ;
  LAYER M1 ;
        RECT 14.352 7.776 14.384 10.284 ;
  LAYER M1 ;
        RECT 14.416 7.776 14.448 10.284 ;
  LAYER M1 ;
        RECT 14.48 7.776 14.512 10.284 ;
  LAYER M1 ;
        RECT 14.544 7.776 14.576 10.284 ;
  LAYER M1 ;
        RECT 14.608 7.776 14.64 10.284 ;
  LAYER M1 ;
        RECT 14.672 7.776 14.704 10.284 ;
  LAYER M1 ;
        RECT 14.736 7.776 14.768 10.284 ;
  LAYER M1 ;
        RECT 14.8 7.776 14.832 10.284 ;
  LAYER M1 ;
        RECT 14.864 7.776 14.896 10.284 ;
  LAYER M1 ;
        RECT 14.928 7.776 14.96 10.284 ;
  LAYER M2 ;
        RECT 12.604 10.168 15.076 10.2 ;
  LAYER M2 ;
        RECT 12.604 10.104 15.076 10.136 ;
  LAYER M2 ;
        RECT 12.604 10.04 15.076 10.072 ;
  LAYER M2 ;
        RECT 12.604 9.976 15.076 10.008 ;
  LAYER M2 ;
        RECT 12.604 9.912 15.076 9.944 ;
  LAYER M2 ;
        RECT 12.604 9.848 15.076 9.88 ;
  LAYER M2 ;
        RECT 12.604 9.784 15.076 9.816 ;
  LAYER M2 ;
        RECT 12.604 9.72 15.076 9.752 ;
  LAYER M2 ;
        RECT 12.604 9.656 15.076 9.688 ;
  LAYER M2 ;
        RECT 12.604 9.592 15.076 9.624 ;
  LAYER M2 ;
        RECT 12.604 9.528 15.076 9.56 ;
  LAYER M2 ;
        RECT 12.604 9.464 15.076 9.496 ;
  LAYER M2 ;
        RECT 12.604 9.4 15.076 9.432 ;
  LAYER M2 ;
        RECT 12.604 9.336 15.076 9.368 ;
  LAYER M2 ;
        RECT 12.604 9.272 15.076 9.304 ;
  LAYER M2 ;
        RECT 12.604 9.208 15.076 9.24 ;
  LAYER M2 ;
        RECT 12.604 9.144 15.076 9.176 ;
  LAYER M2 ;
        RECT 12.604 9.08 15.076 9.112 ;
  LAYER M2 ;
        RECT 12.604 9.016 15.076 9.048 ;
  LAYER M2 ;
        RECT 12.604 8.952 15.076 8.984 ;
  LAYER M2 ;
        RECT 12.604 8.888 15.076 8.92 ;
  LAYER M2 ;
        RECT 12.604 8.824 15.076 8.856 ;
  LAYER M2 ;
        RECT 12.604 8.76 15.076 8.792 ;
  LAYER M2 ;
        RECT 12.604 8.696 15.076 8.728 ;
  LAYER M2 ;
        RECT 12.604 8.632 15.076 8.664 ;
  LAYER M2 ;
        RECT 12.604 8.568 15.076 8.6 ;
  LAYER M2 ;
        RECT 12.604 8.504 15.076 8.536 ;
  LAYER M2 ;
        RECT 12.604 8.44 15.076 8.472 ;
  LAYER M2 ;
        RECT 12.604 8.376 15.076 8.408 ;
  LAYER M2 ;
        RECT 12.604 8.312 15.076 8.344 ;
  LAYER M2 ;
        RECT 12.604 8.248 15.076 8.28 ;
  LAYER M2 ;
        RECT 12.604 8.184 15.076 8.216 ;
  LAYER M2 ;
        RECT 12.604 8.12 15.076 8.152 ;
  LAYER M2 ;
        RECT 12.604 8.056 15.076 8.088 ;
  LAYER M2 ;
        RECT 12.604 7.992 15.076 8.024 ;
  LAYER M2 ;
        RECT 12.604 7.928 15.076 7.96 ;
  LAYER M3 ;
        RECT 12.624 7.776 12.656 10.284 ;
  LAYER M3 ;
        RECT 12.688 7.776 12.72 10.284 ;
  LAYER M3 ;
        RECT 12.752 7.776 12.784 10.284 ;
  LAYER M3 ;
        RECT 12.816 7.776 12.848 10.284 ;
  LAYER M3 ;
        RECT 12.88 7.776 12.912 10.284 ;
  LAYER M3 ;
        RECT 12.944 7.776 12.976 10.284 ;
  LAYER M3 ;
        RECT 13.008 7.776 13.04 10.284 ;
  LAYER M3 ;
        RECT 13.072 7.776 13.104 10.284 ;
  LAYER M3 ;
        RECT 13.136 7.776 13.168 10.284 ;
  LAYER M3 ;
        RECT 13.2 7.776 13.232 10.284 ;
  LAYER M3 ;
        RECT 13.264 7.776 13.296 10.284 ;
  LAYER M3 ;
        RECT 13.328 7.776 13.36 10.284 ;
  LAYER M3 ;
        RECT 13.392 7.776 13.424 10.284 ;
  LAYER M3 ;
        RECT 13.456 7.776 13.488 10.284 ;
  LAYER M3 ;
        RECT 13.52 7.776 13.552 10.284 ;
  LAYER M3 ;
        RECT 13.584 7.776 13.616 10.284 ;
  LAYER M3 ;
        RECT 13.648 7.776 13.68 10.284 ;
  LAYER M3 ;
        RECT 13.712 7.776 13.744 10.284 ;
  LAYER M3 ;
        RECT 13.776 7.776 13.808 10.284 ;
  LAYER M3 ;
        RECT 13.84 7.776 13.872 10.284 ;
  LAYER M3 ;
        RECT 13.904 7.776 13.936 10.284 ;
  LAYER M3 ;
        RECT 13.968 7.776 14 10.284 ;
  LAYER M3 ;
        RECT 14.032 7.776 14.064 10.284 ;
  LAYER M3 ;
        RECT 14.096 7.776 14.128 10.284 ;
  LAYER M3 ;
        RECT 14.16 7.776 14.192 10.284 ;
  LAYER M3 ;
        RECT 14.224 7.776 14.256 10.284 ;
  LAYER M3 ;
        RECT 14.288 7.776 14.32 10.284 ;
  LAYER M3 ;
        RECT 14.352 7.776 14.384 10.284 ;
  LAYER M3 ;
        RECT 14.416 7.776 14.448 10.284 ;
  LAYER M3 ;
        RECT 14.48 7.776 14.512 10.284 ;
  LAYER M3 ;
        RECT 14.544 7.776 14.576 10.284 ;
  LAYER M3 ;
        RECT 14.608 7.776 14.64 10.284 ;
  LAYER M3 ;
        RECT 14.672 7.776 14.704 10.284 ;
  LAYER M3 ;
        RECT 14.736 7.776 14.768 10.284 ;
  LAYER M3 ;
        RECT 14.8 7.776 14.832 10.284 ;
  LAYER M3 ;
        RECT 14.864 7.776 14.896 10.284 ;
  LAYER M3 ;
        RECT 14.928 7.776 14.96 10.284 ;
  LAYER M3 ;
        RECT 15.024 7.776 15.056 10.284 ;
  LAYER M1 ;
        RECT 12.639 7.812 12.641 10.248 ;
  LAYER M1 ;
        RECT 12.719 7.812 12.721 10.248 ;
  LAYER M1 ;
        RECT 12.799 7.812 12.801 10.248 ;
  LAYER M1 ;
        RECT 12.879 7.812 12.881 10.248 ;
  LAYER M1 ;
        RECT 12.959 7.812 12.961 10.248 ;
  LAYER M1 ;
        RECT 13.039 7.812 13.041 10.248 ;
  LAYER M1 ;
        RECT 13.119 7.812 13.121 10.248 ;
  LAYER M1 ;
        RECT 13.199 7.812 13.201 10.248 ;
  LAYER M1 ;
        RECT 13.279 7.812 13.281 10.248 ;
  LAYER M1 ;
        RECT 13.359 7.812 13.361 10.248 ;
  LAYER M1 ;
        RECT 13.439 7.812 13.441 10.248 ;
  LAYER M1 ;
        RECT 13.519 7.812 13.521 10.248 ;
  LAYER M1 ;
        RECT 13.599 7.812 13.601 10.248 ;
  LAYER M1 ;
        RECT 13.679 7.812 13.681 10.248 ;
  LAYER M1 ;
        RECT 13.759 7.812 13.761 10.248 ;
  LAYER M1 ;
        RECT 13.839 7.812 13.841 10.248 ;
  LAYER M1 ;
        RECT 13.919 7.812 13.921 10.248 ;
  LAYER M1 ;
        RECT 13.999 7.812 14.001 10.248 ;
  LAYER M1 ;
        RECT 14.079 7.812 14.081 10.248 ;
  LAYER M1 ;
        RECT 14.159 7.812 14.161 10.248 ;
  LAYER M1 ;
        RECT 14.239 7.812 14.241 10.248 ;
  LAYER M1 ;
        RECT 14.319 7.812 14.321 10.248 ;
  LAYER M1 ;
        RECT 14.399 7.812 14.401 10.248 ;
  LAYER M1 ;
        RECT 14.479 7.812 14.481 10.248 ;
  LAYER M1 ;
        RECT 14.559 7.812 14.561 10.248 ;
  LAYER M1 ;
        RECT 14.639 7.812 14.641 10.248 ;
  LAYER M1 ;
        RECT 14.719 7.812 14.721 10.248 ;
  LAYER M1 ;
        RECT 14.799 7.812 14.801 10.248 ;
  LAYER M1 ;
        RECT 14.879 7.812 14.881 10.248 ;
  LAYER M1 ;
        RECT 14.959 7.812 14.961 10.248 ;
  LAYER M2 ;
        RECT 12.64 10.247 15.04 10.249 ;
  LAYER M2 ;
        RECT 12.64 10.163 15.04 10.165 ;
  LAYER M2 ;
        RECT 12.64 10.079 15.04 10.081 ;
  LAYER M2 ;
        RECT 12.64 9.995 15.04 9.997 ;
  LAYER M2 ;
        RECT 12.64 9.911 15.04 9.913 ;
  LAYER M2 ;
        RECT 12.64 9.827 15.04 9.829 ;
  LAYER M2 ;
        RECT 12.64 9.743 15.04 9.745 ;
  LAYER M2 ;
        RECT 12.64 9.659 15.04 9.661 ;
  LAYER M2 ;
        RECT 12.64 9.575 15.04 9.577 ;
  LAYER M2 ;
        RECT 12.64 9.491 15.04 9.493 ;
  LAYER M2 ;
        RECT 12.64 9.407 15.04 9.409 ;
  LAYER M2 ;
        RECT 12.64 9.323 15.04 9.325 ;
  LAYER M2 ;
        RECT 12.64 9.2395 15.04 9.2415 ;
  LAYER M2 ;
        RECT 12.64 9.155 15.04 9.157 ;
  LAYER M2 ;
        RECT 12.64 9.071 15.04 9.073 ;
  LAYER M2 ;
        RECT 12.64 8.987 15.04 8.989 ;
  LAYER M2 ;
        RECT 12.64 8.903 15.04 8.905 ;
  LAYER M2 ;
        RECT 12.64 8.819 15.04 8.821 ;
  LAYER M2 ;
        RECT 12.64 8.735 15.04 8.737 ;
  LAYER M2 ;
        RECT 12.64 8.651 15.04 8.653 ;
  LAYER M2 ;
        RECT 12.64 8.567 15.04 8.569 ;
  LAYER M2 ;
        RECT 12.64 8.483 15.04 8.485 ;
  LAYER M2 ;
        RECT 12.64 8.399 15.04 8.401 ;
  LAYER M2 ;
        RECT 12.64 8.315 15.04 8.317 ;
  LAYER M2 ;
        RECT 12.64 8.231 15.04 8.233 ;
  LAYER M2 ;
        RECT 12.64 8.147 15.04 8.149 ;
  LAYER M2 ;
        RECT 12.64 8.063 15.04 8.065 ;
  LAYER M2 ;
        RECT 12.64 7.979 15.04 7.981 ;
  LAYER M2 ;
        RECT 12.64 7.895 15.04 7.897 ;
  LAYER M1 ;
        RECT 12.624 4.836 12.656 7.344 ;
  LAYER M1 ;
        RECT 12.688 4.836 12.72 7.344 ;
  LAYER M1 ;
        RECT 12.752 4.836 12.784 7.344 ;
  LAYER M1 ;
        RECT 12.816 4.836 12.848 7.344 ;
  LAYER M1 ;
        RECT 12.88 4.836 12.912 7.344 ;
  LAYER M1 ;
        RECT 12.944 4.836 12.976 7.344 ;
  LAYER M1 ;
        RECT 13.008 4.836 13.04 7.344 ;
  LAYER M1 ;
        RECT 13.072 4.836 13.104 7.344 ;
  LAYER M1 ;
        RECT 13.136 4.836 13.168 7.344 ;
  LAYER M1 ;
        RECT 13.2 4.836 13.232 7.344 ;
  LAYER M1 ;
        RECT 13.264 4.836 13.296 7.344 ;
  LAYER M1 ;
        RECT 13.328 4.836 13.36 7.344 ;
  LAYER M1 ;
        RECT 13.392 4.836 13.424 7.344 ;
  LAYER M1 ;
        RECT 13.456 4.836 13.488 7.344 ;
  LAYER M1 ;
        RECT 13.52 4.836 13.552 7.344 ;
  LAYER M1 ;
        RECT 13.584 4.836 13.616 7.344 ;
  LAYER M1 ;
        RECT 13.648 4.836 13.68 7.344 ;
  LAYER M1 ;
        RECT 13.712 4.836 13.744 7.344 ;
  LAYER M1 ;
        RECT 13.776 4.836 13.808 7.344 ;
  LAYER M1 ;
        RECT 13.84 4.836 13.872 7.344 ;
  LAYER M1 ;
        RECT 13.904 4.836 13.936 7.344 ;
  LAYER M1 ;
        RECT 13.968 4.836 14 7.344 ;
  LAYER M1 ;
        RECT 14.032 4.836 14.064 7.344 ;
  LAYER M1 ;
        RECT 14.096 4.836 14.128 7.344 ;
  LAYER M1 ;
        RECT 14.16 4.836 14.192 7.344 ;
  LAYER M1 ;
        RECT 14.224 4.836 14.256 7.344 ;
  LAYER M1 ;
        RECT 14.288 4.836 14.32 7.344 ;
  LAYER M1 ;
        RECT 14.352 4.836 14.384 7.344 ;
  LAYER M1 ;
        RECT 14.416 4.836 14.448 7.344 ;
  LAYER M1 ;
        RECT 14.48 4.836 14.512 7.344 ;
  LAYER M1 ;
        RECT 14.544 4.836 14.576 7.344 ;
  LAYER M1 ;
        RECT 14.608 4.836 14.64 7.344 ;
  LAYER M1 ;
        RECT 14.672 4.836 14.704 7.344 ;
  LAYER M1 ;
        RECT 14.736 4.836 14.768 7.344 ;
  LAYER M1 ;
        RECT 14.8 4.836 14.832 7.344 ;
  LAYER M1 ;
        RECT 14.864 4.836 14.896 7.344 ;
  LAYER M1 ;
        RECT 14.928 4.836 14.96 7.344 ;
  LAYER M2 ;
        RECT 12.604 7.228 15.076 7.26 ;
  LAYER M2 ;
        RECT 12.604 7.164 15.076 7.196 ;
  LAYER M2 ;
        RECT 12.604 7.1 15.076 7.132 ;
  LAYER M2 ;
        RECT 12.604 7.036 15.076 7.068 ;
  LAYER M2 ;
        RECT 12.604 6.972 15.076 7.004 ;
  LAYER M2 ;
        RECT 12.604 6.908 15.076 6.94 ;
  LAYER M2 ;
        RECT 12.604 6.844 15.076 6.876 ;
  LAYER M2 ;
        RECT 12.604 6.78 15.076 6.812 ;
  LAYER M2 ;
        RECT 12.604 6.716 15.076 6.748 ;
  LAYER M2 ;
        RECT 12.604 6.652 15.076 6.684 ;
  LAYER M2 ;
        RECT 12.604 6.588 15.076 6.62 ;
  LAYER M2 ;
        RECT 12.604 6.524 15.076 6.556 ;
  LAYER M2 ;
        RECT 12.604 6.46 15.076 6.492 ;
  LAYER M2 ;
        RECT 12.604 6.396 15.076 6.428 ;
  LAYER M2 ;
        RECT 12.604 6.332 15.076 6.364 ;
  LAYER M2 ;
        RECT 12.604 6.268 15.076 6.3 ;
  LAYER M2 ;
        RECT 12.604 6.204 15.076 6.236 ;
  LAYER M2 ;
        RECT 12.604 6.14 15.076 6.172 ;
  LAYER M2 ;
        RECT 12.604 6.076 15.076 6.108 ;
  LAYER M2 ;
        RECT 12.604 6.012 15.076 6.044 ;
  LAYER M2 ;
        RECT 12.604 5.948 15.076 5.98 ;
  LAYER M2 ;
        RECT 12.604 5.884 15.076 5.916 ;
  LAYER M2 ;
        RECT 12.604 5.82 15.076 5.852 ;
  LAYER M2 ;
        RECT 12.604 5.756 15.076 5.788 ;
  LAYER M2 ;
        RECT 12.604 5.692 15.076 5.724 ;
  LAYER M2 ;
        RECT 12.604 5.628 15.076 5.66 ;
  LAYER M2 ;
        RECT 12.604 5.564 15.076 5.596 ;
  LAYER M2 ;
        RECT 12.604 5.5 15.076 5.532 ;
  LAYER M2 ;
        RECT 12.604 5.436 15.076 5.468 ;
  LAYER M2 ;
        RECT 12.604 5.372 15.076 5.404 ;
  LAYER M2 ;
        RECT 12.604 5.308 15.076 5.34 ;
  LAYER M2 ;
        RECT 12.604 5.244 15.076 5.276 ;
  LAYER M2 ;
        RECT 12.604 5.18 15.076 5.212 ;
  LAYER M2 ;
        RECT 12.604 5.116 15.076 5.148 ;
  LAYER M2 ;
        RECT 12.604 5.052 15.076 5.084 ;
  LAYER M2 ;
        RECT 12.604 4.988 15.076 5.02 ;
  LAYER M3 ;
        RECT 12.624 4.836 12.656 7.344 ;
  LAYER M3 ;
        RECT 12.688 4.836 12.72 7.344 ;
  LAYER M3 ;
        RECT 12.752 4.836 12.784 7.344 ;
  LAYER M3 ;
        RECT 12.816 4.836 12.848 7.344 ;
  LAYER M3 ;
        RECT 12.88 4.836 12.912 7.344 ;
  LAYER M3 ;
        RECT 12.944 4.836 12.976 7.344 ;
  LAYER M3 ;
        RECT 13.008 4.836 13.04 7.344 ;
  LAYER M3 ;
        RECT 13.072 4.836 13.104 7.344 ;
  LAYER M3 ;
        RECT 13.136 4.836 13.168 7.344 ;
  LAYER M3 ;
        RECT 13.2 4.836 13.232 7.344 ;
  LAYER M3 ;
        RECT 13.264 4.836 13.296 7.344 ;
  LAYER M3 ;
        RECT 13.328 4.836 13.36 7.344 ;
  LAYER M3 ;
        RECT 13.392 4.836 13.424 7.344 ;
  LAYER M3 ;
        RECT 13.456 4.836 13.488 7.344 ;
  LAYER M3 ;
        RECT 13.52 4.836 13.552 7.344 ;
  LAYER M3 ;
        RECT 13.584 4.836 13.616 7.344 ;
  LAYER M3 ;
        RECT 13.648 4.836 13.68 7.344 ;
  LAYER M3 ;
        RECT 13.712 4.836 13.744 7.344 ;
  LAYER M3 ;
        RECT 13.776 4.836 13.808 7.344 ;
  LAYER M3 ;
        RECT 13.84 4.836 13.872 7.344 ;
  LAYER M3 ;
        RECT 13.904 4.836 13.936 7.344 ;
  LAYER M3 ;
        RECT 13.968 4.836 14 7.344 ;
  LAYER M3 ;
        RECT 14.032 4.836 14.064 7.344 ;
  LAYER M3 ;
        RECT 14.096 4.836 14.128 7.344 ;
  LAYER M3 ;
        RECT 14.16 4.836 14.192 7.344 ;
  LAYER M3 ;
        RECT 14.224 4.836 14.256 7.344 ;
  LAYER M3 ;
        RECT 14.288 4.836 14.32 7.344 ;
  LAYER M3 ;
        RECT 14.352 4.836 14.384 7.344 ;
  LAYER M3 ;
        RECT 14.416 4.836 14.448 7.344 ;
  LAYER M3 ;
        RECT 14.48 4.836 14.512 7.344 ;
  LAYER M3 ;
        RECT 14.544 4.836 14.576 7.344 ;
  LAYER M3 ;
        RECT 14.608 4.836 14.64 7.344 ;
  LAYER M3 ;
        RECT 14.672 4.836 14.704 7.344 ;
  LAYER M3 ;
        RECT 14.736 4.836 14.768 7.344 ;
  LAYER M3 ;
        RECT 14.8 4.836 14.832 7.344 ;
  LAYER M3 ;
        RECT 14.864 4.836 14.896 7.344 ;
  LAYER M3 ;
        RECT 14.928 4.836 14.96 7.344 ;
  LAYER M3 ;
        RECT 15.024 4.836 15.056 7.344 ;
  LAYER M1 ;
        RECT 12.639 4.872 12.641 7.308 ;
  LAYER M1 ;
        RECT 12.719 4.872 12.721 7.308 ;
  LAYER M1 ;
        RECT 12.799 4.872 12.801 7.308 ;
  LAYER M1 ;
        RECT 12.879 4.872 12.881 7.308 ;
  LAYER M1 ;
        RECT 12.959 4.872 12.961 7.308 ;
  LAYER M1 ;
        RECT 13.039 4.872 13.041 7.308 ;
  LAYER M1 ;
        RECT 13.119 4.872 13.121 7.308 ;
  LAYER M1 ;
        RECT 13.199 4.872 13.201 7.308 ;
  LAYER M1 ;
        RECT 13.279 4.872 13.281 7.308 ;
  LAYER M1 ;
        RECT 13.359 4.872 13.361 7.308 ;
  LAYER M1 ;
        RECT 13.439 4.872 13.441 7.308 ;
  LAYER M1 ;
        RECT 13.519 4.872 13.521 7.308 ;
  LAYER M1 ;
        RECT 13.599 4.872 13.601 7.308 ;
  LAYER M1 ;
        RECT 13.679 4.872 13.681 7.308 ;
  LAYER M1 ;
        RECT 13.759 4.872 13.761 7.308 ;
  LAYER M1 ;
        RECT 13.839 4.872 13.841 7.308 ;
  LAYER M1 ;
        RECT 13.919 4.872 13.921 7.308 ;
  LAYER M1 ;
        RECT 13.999 4.872 14.001 7.308 ;
  LAYER M1 ;
        RECT 14.079 4.872 14.081 7.308 ;
  LAYER M1 ;
        RECT 14.159 4.872 14.161 7.308 ;
  LAYER M1 ;
        RECT 14.239 4.872 14.241 7.308 ;
  LAYER M1 ;
        RECT 14.319 4.872 14.321 7.308 ;
  LAYER M1 ;
        RECT 14.399 4.872 14.401 7.308 ;
  LAYER M1 ;
        RECT 14.479 4.872 14.481 7.308 ;
  LAYER M1 ;
        RECT 14.559 4.872 14.561 7.308 ;
  LAYER M1 ;
        RECT 14.639 4.872 14.641 7.308 ;
  LAYER M1 ;
        RECT 14.719 4.872 14.721 7.308 ;
  LAYER M1 ;
        RECT 14.799 4.872 14.801 7.308 ;
  LAYER M1 ;
        RECT 14.879 4.872 14.881 7.308 ;
  LAYER M1 ;
        RECT 14.959 4.872 14.961 7.308 ;
  LAYER M2 ;
        RECT 12.64 7.307 15.04 7.309 ;
  LAYER M2 ;
        RECT 12.64 7.223 15.04 7.225 ;
  LAYER M2 ;
        RECT 12.64 7.139 15.04 7.141 ;
  LAYER M2 ;
        RECT 12.64 7.055 15.04 7.057 ;
  LAYER M2 ;
        RECT 12.64 6.971 15.04 6.973 ;
  LAYER M2 ;
        RECT 12.64 6.887 15.04 6.889 ;
  LAYER M2 ;
        RECT 12.64 6.803 15.04 6.805 ;
  LAYER M2 ;
        RECT 12.64 6.719 15.04 6.721 ;
  LAYER M2 ;
        RECT 12.64 6.635 15.04 6.637 ;
  LAYER M2 ;
        RECT 12.64 6.551 15.04 6.553 ;
  LAYER M2 ;
        RECT 12.64 6.467 15.04 6.469 ;
  LAYER M2 ;
        RECT 12.64 6.383 15.04 6.385 ;
  LAYER M2 ;
        RECT 12.64 6.2995 15.04 6.3015 ;
  LAYER M2 ;
        RECT 12.64 6.215 15.04 6.217 ;
  LAYER M2 ;
        RECT 12.64 6.131 15.04 6.133 ;
  LAYER M2 ;
        RECT 12.64 6.047 15.04 6.049 ;
  LAYER M2 ;
        RECT 12.64 5.963 15.04 5.965 ;
  LAYER M2 ;
        RECT 12.64 5.879 15.04 5.881 ;
  LAYER M2 ;
        RECT 12.64 5.795 15.04 5.797 ;
  LAYER M2 ;
        RECT 12.64 5.711 15.04 5.713 ;
  LAYER M2 ;
        RECT 12.64 5.627 15.04 5.629 ;
  LAYER M2 ;
        RECT 12.64 5.543 15.04 5.545 ;
  LAYER M2 ;
        RECT 12.64 5.459 15.04 5.461 ;
  LAYER M2 ;
        RECT 12.64 5.375 15.04 5.377 ;
  LAYER M2 ;
        RECT 12.64 5.291 15.04 5.293 ;
  LAYER M2 ;
        RECT 12.64 5.207 15.04 5.209 ;
  LAYER M2 ;
        RECT 12.64 5.123 15.04 5.125 ;
  LAYER M2 ;
        RECT 12.64 5.039 15.04 5.041 ;
  LAYER M2 ;
        RECT 12.64 4.955 15.04 4.957 ;
  LAYER M1 ;
        RECT 12.624 1.896 12.656 4.404 ;
  LAYER M1 ;
        RECT 12.688 1.896 12.72 4.404 ;
  LAYER M1 ;
        RECT 12.752 1.896 12.784 4.404 ;
  LAYER M1 ;
        RECT 12.816 1.896 12.848 4.404 ;
  LAYER M1 ;
        RECT 12.88 1.896 12.912 4.404 ;
  LAYER M1 ;
        RECT 12.944 1.896 12.976 4.404 ;
  LAYER M1 ;
        RECT 13.008 1.896 13.04 4.404 ;
  LAYER M1 ;
        RECT 13.072 1.896 13.104 4.404 ;
  LAYER M1 ;
        RECT 13.136 1.896 13.168 4.404 ;
  LAYER M1 ;
        RECT 13.2 1.896 13.232 4.404 ;
  LAYER M1 ;
        RECT 13.264 1.896 13.296 4.404 ;
  LAYER M1 ;
        RECT 13.328 1.896 13.36 4.404 ;
  LAYER M1 ;
        RECT 13.392 1.896 13.424 4.404 ;
  LAYER M1 ;
        RECT 13.456 1.896 13.488 4.404 ;
  LAYER M1 ;
        RECT 13.52 1.896 13.552 4.404 ;
  LAYER M1 ;
        RECT 13.584 1.896 13.616 4.404 ;
  LAYER M1 ;
        RECT 13.648 1.896 13.68 4.404 ;
  LAYER M1 ;
        RECT 13.712 1.896 13.744 4.404 ;
  LAYER M1 ;
        RECT 13.776 1.896 13.808 4.404 ;
  LAYER M1 ;
        RECT 13.84 1.896 13.872 4.404 ;
  LAYER M1 ;
        RECT 13.904 1.896 13.936 4.404 ;
  LAYER M1 ;
        RECT 13.968 1.896 14 4.404 ;
  LAYER M1 ;
        RECT 14.032 1.896 14.064 4.404 ;
  LAYER M1 ;
        RECT 14.096 1.896 14.128 4.404 ;
  LAYER M1 ;
        RECT 14.16 1.896 14.192 4.404 ;
  LAYER M1 ;
        RECT 14.224 1.896 14.256 4.404 ;
  LAYER M1 ;
        RECT 14.288 1.896 14.32 4.404 ;
  LAYER M1 ;
        RECT 14.352 1.896 14.384 4.404 ;
  LAYER M1 ;
        RECT 14.416 1.896 14.448 4.404 ;
  LAYER M1 ;
        RECT 14.48 1.896 14.512 4.404 ;
  LAYER M1 ;
        RECT 14.544 1.896 14.576 4.404 ;
  LAYER M1 ;
        RECT 14.608 1.896 14.64 4.404 ;
  LAYER M1 ;
        RECT 14.672 1.896 14.704 4.404 ;
  LAYER M1 ;
        RECT 14.736 1.896 14.768 4.404 ;
  LAYER M1 ;
        RECT 14.8 1.896 14.832 4.404 ;
  LAYER M1 ;
        RECT 14.864 1.896 14.896 4.404 ;
  LAYER M1 ;
        RECT 14.928 1.896 14.96 4.404 ;
  LAYER M2 ;
        RECT 12.604 4.288 15.076 4.32 ;
  LAYER M2 ;
        RECT 12.604 4.224 15.076 4.256 ;
  LAYER M2 ;
        RECT 12.604 4.16 15.076 4.192 ;
  LAYER M2 ;
        RECT 12.604 4.096 15.076 4.128 ;
  LAYER M2 ;
        RECT 12.604 4.032 15.076 4.064 ;
  LAYER M2 ;
        RECT 12.604 3.968 15.076 4 ;
  LAYER M2 ;
        RECT 12.604 3.904 15.076 3.936 ;
  LAYER M2 ;
        RECT 12.604 3.84 15.076 3.872 ;
  LAYER M2 ;
        RECT 12.604 3.776 15.076 3.808 ;
  LAYER M2 ;
        RECT 12.604 3.712 15.076 3.744 ;
  LAYER M2 ;
        RECT 12.604 3.648 15.076 3.68 ;
  LAYER M2 ;
        RECT 12.604 3.584 15.076 3.616 ;
  LAYER M2 ;
        RECT 12.604 3.52 15.076 3.552 ;
  LAYER M2 ;
        RECT 12.604 3.456 15.076 3.488 ;
  LAYER M2 ;
        RECT 12.604 3.392 15.076 3.424 ;
  LAYER M2 ;
        RECT 12.604 3.328 15.076 3.36 ;
  LAYER M2 ;
        RECT 12.604 3.264 15.076 3.296 ;
  LAYER M2 ;
        RECT 12.604 3.2 15.076 3.232 ;
  LAYER M2 ;
        RECT 12.604 3.136 15.076 3.168 ;
  LAYER M2 ;
        RECT 12.604 3.072 15.076 3.104 ;
  LAYER M2 ;
        RECT 12.604 3.008 15.076 3.04 ;
  LAYER M2 ;
        RECT 12.604 2.944 15.076 2.976 ;
  LAYER M2 ;
        RECT 12.604 2.88 15.076 2.912 ;
  LAYER M2 ;
        RECT 12.604 2.816 15.076 2.848 ;
  LAYER M2 ;
        RECT 12.604 2.752 15.076 2.784 ;
  LAYER M2 ;
        RECT 12.604 2.688 15.076 2.72 ;
  LAYER M2 ;
        RECT 12.604 2.624 15.076 2.656 ;
  LAYER M2 ;
        RECT 12.604 2.56 15.076 2.592 ;
  LAYER M2 ;
        RECT 12.604 2.496 15.076 2.528 ;
  LAYER M2 ;
        RECT 12.604 2.432 15.076 2.464 ;
  LAYER M2 ;
        RECT 12.604 2.368 15.076 2.4 ;
  LAYER M2 ;
        RECT 12.604 2.304 15.076 2.336 ;
  LAYER M2 ;
        RECT 12.604 2.24 15.076 2.272 ;
  LAYER M2 ;
        RECT 12.604 2.176 15.076 2.208 ;
  LAYER M2 ;
        RECT 12.604 2.112 15.076 2.144 ;
  LAYER M2 ;
        RECT 12.604 2.048 15.076 2.08 ;
  LAYER M3 ;
        RECT 12.624 1.896 12.656 4.404 ;
  LAYER M3 ;
        RECT 12.688 1.896 12.72 4.404 ;
  LAYER M3 ;
        RECT 12.752 1.896 12.784 4.404 ;
  LAYER M3 ;
        RECT 12.816 1.896 12.848 4.404 ;
  LAYER M3 ;
        RECT 12.88 1.896 12.912 4.404 ;
  LAYER M3 ;
        RECT 12.944 1.896 12.976 4.404 ;
  LAYER M3 ;
        RECT 13.008 1.896 13.04 4.404 ;
  LAYER M3 ;
        RECT 13.072 1.896 13.104 4.404 ;
  LAYER M3 ;
        RECT 13.136 1.896 13.168 4.404 ;
  LAYER M3 ;
        RECT 13.2 1.896 13.232 4.404 ;
  LAYER M3 ;
        RECT 13.264 1.896 13.296 4.404 ;
  LAYER M3 ;
        RECT 13.328 1.896 13.36 4.404 ;
  LAYER M3 ;
        RECT 13.392 1.896 13.424 4.404 ;
  LAYER M3 ;
        RECT 13.456 1.896 13.488 4.404 ;
  LAYER M3 ;
        RECT 13.52 1.896 13.552 4.404 ;
  LAYER M3 ;
        RECT 13.584 1.896 13.616 4.404 ;
  LAYER M3 ;
        RECT 13.648 1.896 13.68 4.404 ;
  LAYER M3 ;
        RECT 13.712 1.896 13.744 4.404 ;
  LAYER M3 ;
        RECT 13.776 1.896 13.808 4.404 ;
  LAYER M3 ;
        RECT 13.84 1.896 13.872 4.404 ;
  LAYER M3 ;
        RECT 13.904 1.896 13.936 4.404 ;
  LAYER M3 ;
        RECT 13.968 1.896 14 4.404 ;
  LAYER M3 ;
        RECT 14.032 1.896 14.064 4.404 ;
  LAYER M3 ;
        RECT 14.096 1.896 14.128 4.404 ;
  LAYER M3 ;
        RECT 14.16 1.896 14.192 4.404 ;
  LAYER M3 ;
        RECT 14.224 1.896 14.256 4.404 ;
  LAYER M3 ;
        RECT 14.288 1.896 14.32 4.404 ;
  LAYER M3 ;
        RECT 14.352 1.896 14.384 4.404 ;
  LAYER M3 ;
        RECT 14.416 1.896 14.448 4.404 ;
  LAYER M3 ;
        RECT 14.48 1.896 14.512 4.404 ;
  LAYER M3 ;
        RECT 14.544 1.896 14.576 4.404 ;
  LAYER M3 ;
        RECT 14.608 1.896 14.64 4.404 ;
  LAYER M3 ;
        RECT 14.672 1.896 14.704 4.404 ;
  LAYER M3 ;
        RECT 14.736 1.896 14.768 4.404 ;
  LAYER M3 ;
        RECT 14.8 1.896 14.832 4.404 ;
  LAYER M3 ;
        RECT 14.864 1.896 14.896 4.404 ;
  LAYER M3 ;
        RECT 14.928 1.896 14.96 4.404 ;
  LAYER M3 ;
        RECT 15.024 1.896 15.056 4.404 ;
  LAYER M1 ;
        RECT 12.639 1.932 12.641 4.368 ;
  LAYER M1 ;
        RECT 12.719 1.932 12.721 4.368 ;
  LAYER M1 ;
        RECT 12.799 1.932 12.801 4.368 ;
  LAYER M1 ;
        RECT 12.879 1.932 12.881 4.368 ;
  LAYER M1 ;
        RECT 12.959 1.932 12.961 4.368 ;
  LAYER M1 ;
        RECT 13.039 1.932 13.041 4.368 ;
  LAYER M1 ;
        RECT 13.119 1.932 13.121 4.368 ;
  LAYER M1 ;
        RECT 13.199 1.932 13.201 4.368 ;
  LAYER M1 ;
        RECT 13.279 1.932 13.281 4.368 ;
  LAYER M1 ;
        RECT 13.359 1.932 13.361 4.368 ;
  LAYER M1 ;
        RECT 13.439 1.932 13.441 4.368 ;
  LAYER M1 ;
        RECT 13.519 1.932 13.521 4.368 ;
  LAYER M1 ;
        RECT 13.599 1.932 13.601 4.368 ;
  LAYER M1 ;
        RECT 13.679 1.932 13.681 4.368 ;
  LAYER M1 ;
        RECT 13.759 1.932 13.761 4.368 ;
  LAYER M1 ;
        RECT 13.839 1.932 13.841 4.368 ;
  LAYER M1 ;
        RECT 13.919 1.932 13.921 4.368 ;
  LAYER M1 ;
        RECT 13.999 1.932 14.001 4.368 ;
  LAYER M1 ;
        RECT 14.079 1.932 14.081 4.368 ;
  LAYER M1 ;
        RECT 14.159 1.932 14.161 4.368 ;
  LAYER M1 ;
        RECT 14.239 1.932 14.241 4.368 ;
  LAYER M1 ;
        RECT 14.319 1.932 14.321 4.368 ;
  LAYER M1 ;
        RECT 14.399 1.932 14.401 4.368 ;
  LAYER M1 ;
        RECT 14.479 1.932 14.481 4.368 ;
  LAYER M1 ;
        RECT 14.559 1.932 14.561 4.368 ;
  LAYER M1 ;
        RECT 14.639 1.932 14.641 4.368 ;
  LAYER M1 ;
        RECT 14.719 1.932 14.721 4.368 ;
  LAYER M1 ;
        RECT 14.799 1.932 14.801 4.368 ;
  LAYER M1 ;
        RECT 14.879 1.932 14.881 4.368 ;
  LAYER M1 ;
        RECT 14.959 1.932 14.961 4.368 ;
  LAYER M2 ;
        RECT 12.64 4.367 15.04 4.369 ;
  LAYER M2 ;
        RECT 12.64 4.283 15.04 4.285 ;
  LAYER M2 ;
        RECT 12.64 4.199 15.04 4.201 ;
  LAYER M2 ;
        RECT 12.64 4.115 15.04 4.117 ;
  LAYER M2 ;
        RECT 12.64 4.031 15.04 4.033 ;
  LAYER M2 ;
        RECT 12.64 3.947 15.04 3.949 ;
  LAYER M2 ;
        RECT 12.64 3.863 15.04 3.865 ;
  LAYER M2 ;
        RECT 12.64 3.779 15.04 3.781 ;
  LAYER M2 ;
        RECT 12.64 3.695 15.04 3.697 ;
  LAYER M2 ;
        RECT 12.64 3.611 15.04 3.613 ;
  LAYER M2 ;
        RECT 12.64 3.527 15.04 3.529 ;
  LAYER M2 ;
        RECT 12.64 3.443 15.04 3.445 ;
  LAYER M2 ;
        RECT 12.64 3.3595 15.04 3.3615 ;
  LAYER M2 ;
        RECT 12.64 3.275 15.04 3.277 ;
  LAYER M2 ;
        RECT 12.64 3.191 15.04 3.193 ;
  LAYER M2 ;
        RECT 12.64 3.107 15.04 3.109 ;
  LAYER M2 ;
        RECT 12.64 3.023 15.04 3.025 ;
  LAYER M2 ;
        RECT 12.64 2.939 15.04 2.941 ;
  LAYER M2 ;
        RECT 12.64 2.855 15.04 2.857 ;
  LAYER M2 ;
        RECT 12.64 2.771 15.04 2.773 ;
  LAYER M2 ;
        RECT 12.64 2.687 15.04 2.689 ;
  LAYER M2 ;
        RECT 12.64 2.603 15.04 2.605 ;
  LAYER M2 ;
        RECT 12.64 2.519 15.04 2.521 ;
  LAYER M2 ;
        RECT 12.64 2.435 15.04 2.437 ;
  LAYER M2 ;
        RECT 12.64 2.351 15.04 2.353 ;
  LAYER M2 ;
        RECT 12.64 2.267 15.04 2.269 ;
  LAYER M2 ;
        RECT 12.64 2.183 15.04 2.185 ;
  LAYER M2 ;
        RECT 12.64 2.099 15.04 2.101 ;
  LAYER M2 ;
        RECT 12.64 2.015 15.04 2.017 ;
  END 
END switched_capacitor_combination
