MACRO CKT_OBS_LEF
  ORIGIN 0 0 ;
  FOREIGN CKT_OBS_LEF 0 0 ;
  SIZE 1.542 BY 3.84 ;
  PIN VOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.294 1.15 1.218 1.19 ;
      LAYER M2 ;
        RECT 0.186 0.79 1.326 0.83 ;
      LAYER M2 ;
        RECT 0.294 1.78 1.218 1.82 ;
      LAYER M2 ;
        RECT 0.186 1.42 1.326 1.46 ;
      LAYER M2 ;
        RECT 0.186 2.95 1.326 2.99 ;
      LAYER M2 ;
        RECT 0.186 2.32 1.326 2.36 ;
      LAYER M3 ;
        RECT 0.618 2.32 0.678 2.99 ;
      LAYER M2 ;
        RECT 0.618 1.78 0.678 1.82 ;
      LAYER M3 ;
        RECT 0.618 1.8 0.678 2.34 ;
    END
  END VOP
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.294 2.59 1.218 2.63 ;
      LAYER M2 ;
        RECT 0.294 1.96 1.218 2 ;
      LAYER M3 ;
        RECT 0.726 1.96 0.786 2.63 ;
    END
  END VIN
  OBS 
  LAYER M1 ;
        RECT 0.186 0.07 0.246 1.64 ;
  LAYER M1 ;
        RECT 0.402 0.07 0.462 1.64 ;
  LAYER M1 ;
        RECT 0.618 0.07 0.678 1.64 ;
  LAYER M1 ;
        RECT 0.834 0.07 0.894 1.64 ;
  LAYER M1 ;
        RECT 1.05 0.07 1.11 1.64 ;
  LAYER M1 ;
        RECT 1.266 0.07 1.326 1.64 ;
  LAYER M1 ;
        RECT 0.294 0.7 0.354 1.82 ;
  LAYER M1 ;
        RECT 0.51 0.7 0.57 1.82 ;
  LAYER M1 ;
        RECT 0.942 0.7 1.002 1.82 ;
  LAYER M1 ;
        RECT 1.158 0.7 1.218 1.82 ;
  LAYER M2 ;
        RECT 0.294 1.15 1.218 1.19 ;
  LAYER M2 ;
        RECT 0.186 0.79 1.326 0.83 ;
  LAYER M2 ;
        RECT 0.294 1.78 1.218 1.82 ;
  LAYER M2 ;
        RECT 0.186 1.42 1.326 1.46 ;
  LAYER M2 ;
        RECT 0.186 0.34 1.326 0.38 ;
  LAYER M2 ;
        RECT 0.186 0.97 1.326 1.01 ;
  LAYER M2 ;
        RECT 0.186 1.6 1.326 1.64 ;
  LAYER M1 ;
        RECT 0.186 2.14 0.246 3.71 ;
  LAYER M1 ;
        RECT 0.402 2.14 0.462 3.71 ;
  LAYER M1 ;
        RECT 0.618 2.14 0.678 3.71 ;
  LAYER M1 ;
        RECT 0.834 2.14 0.894 3.71 ;
  LAYER M1 ;
        RECT 1.05 2.14 1.11 3.71 ;
  LAYER M1 ;
        RECT 1.266 2.14 1.326 3.71 ;
  LAYER M1 ;
        RECT 0.294 2.77 0.354 3.08 ;
  LAYER M1 ;
        RECT 0.294 2.59 0.354 2.72 ;
  LAYER M1 ;
        RECT 0.294 2.14 0.354 2.45 ;
  LAYER M1 ;
        RECT 0.294 1.96 0.354 2.09 ;
  LAYER M1 ;
        RECT 0.51 2.77 0.57 3.08 ;
  LAYER M1 ;
        RECT 0.51 2.59 0.57 2.72 ;
  LAYER M1 ;
        RECT 0.51 2.14 0.57 2.45 ;
  LAYER M1 ;
        RECT 0.51 1.96 0.57 2.09 ;
  LAYER M1 ;
        RECT 0.942 2.77 1.002 3.08 ;
  LAYER M1 ;
        RECT 0.942 2.59 1.002 2.72 ;
  LAYER M1 ;
        RECT 0.942 2.14 1.002 2.45 ;
  LAYER M1 ;
        RECT 0.942 1.96 1.002 2.09 ;
  LAYER M1 ;
        RECT 1.158 2.77 1.218 3.08 ;
  LAYER M1 ;
        RECT 1.158 2.59 1.218 2.72 ;
  LAYER M1 ;
        RECT 1.158 2.14 1.218 2.45 ;
  LAYER M1 ;
        RECT 1.158 1.96 1.218 2.09 ;
  LAYER M2 ;
        RECT 0.186 2.95 1.326 2.99 ;
  LAYER M2 ;
        RECT 0.186 2.32 1.326 2.36 ;
  LAYER M3 ;
        RECT 0.618 2.32 0.678 2.99 ;
  LAYER M2 ;
        RECT 0.294 2.59 1.218 2.63 ;
  LAYER M2 ;
        RECT 0.294 1.96 1.218 2 ;
  LAYER M3 ;
        RECT 0.726 1.96 0.786 2.63 ;
  LAYER M2 ;
        RECT 0.186 3.58 1.326 3.62 ;
  LAYER M2 ;
        RECT 0.186 2.77 1.326 2.81 ;
  LAYER M2 ;
        RECT 0.186 2.14 1.326 2.18 ;
  END 
  OBS
    LAYER Poly ;
      RECT 0 0 1.512 1.89 ;
    LAYER Poly ;
      RECT -0.0399 -0.0399 1.5818 3.8798 ;
    LAYER Boundary ;
      RECT 0 0 0.108 0.63 ;
    LAYER Boundary ;
      RECT 0.108 0 0.756 0.63 ;
    LAYER Boundary ;
      RECT 0.756 0 1.404 0.63 ;
    LAYER Boundary ;
      RECT 1.404 0 1.512 0.63 ;
    LAYER Boundary ;
      RECT 0 0.63 0.108 1.26 ;
    LAYER Boundary ;
      RECT 0.108 0.63 0.756 1.26 ;
    LAYER Boundary ;
      RECT 0.756 0.63 1.404 1.26 ;
    LAYER Boundary ;
      RECT 1.404 0.63 1.512 1.26 ;
    LAYER Boundary ;
      RECT 0 1.26 0.108 1.89 ;
    LAYER Boundary ;
      RECT 0.108 1.26 0.756 1.89 ;
    LAYER Boundary ;
      RECT 0.756 1.26 1.404 1.89 ;
    LAYER Boundary ;
      RECT 1.404 1.26 1.512 1.89 ;
    LAYER Boundary ;
      RECT 0 0 0.108 0.63 ;
    LAYER Boundary ;
      RECT 0.108 0 0.756 0.63 ;
    LAYER Boundary ;
      RECT 0.756 0 1.404 0.63 ;
    LAYER Boundary ;
      RECT 1.404 0 1.512 0.63 ;
    LAYER Boundary ;
      RECT 0 0.63 0.108 1.26 ;
    LAYER Boundary ;
      RECT 0.108 0.63 0.756 1.26 ;
    LAYER Boundary ;
      RECT 0.756 0.63 1.404 1.26 ;
    LAYER Boundary ;
      RECT 1.404 0.63 1.512 1.26 ;
    LAYER Boundary ;
      RECT 0 1.26 0.108 1.89 ;
    LAYER Boundary ;
      RECT 0.108 1.26 0.756 1.89 ;
    LAYER Boundary ;
      RECT 0.756 1.26 1.404 1.89 ;
    LAYER Boundary ;
      RECT 1.404 1.26 1.512 1.89 ;
    LAYER M1 ;
      RECT 0.186 0.07 0.246 1.64 ;
    LAYER M1 ;
      RECT 0.402 0.07 0.462 1.64 ;
    LAYER M1 ;
      RECT 0.618 0.07 0.678 1.64 ;
    LAYER M1 ;
      RECT 0.834 0.07 0.894 1.64 ;
    LAYER M1 ;
      RECT 1.05 0.07 1.11 1.64 ;
    LAYER M1 ;
      RECT 1.266 0.07 1.326 1.64 ;
    LAYER M1 ;
      RECT 0.294 0.7 0.354 1.82 ;
    LAYER M1 ;
      RECT 0.51 0.7 0.57 1.82 ;
    LAYER M1 ;
      RECT 0.942 0.7 1.002 1.82 ;
    LAYER M1 ;
      RECT 1.158 0.7 1.218 1.82 ;
    LAYER M1 ;
      RECT 0.186 0.07 0.246 1.64 ;
    LAYER M1 ;
      RECT 0.402 0.07 0.462 1.64 ;
    LAYER M1 ;
      RECT 0.618 0.07 0.678 1.64 ;
    LAYER M1 ;
      RECT 0.834 0.07 0.894 1.64 ;
    LAYER M1 ;
      RECT 1.05 0.07 1.11 1.64 ;
    LAYER M1 ;
      RECT 1.266 0.07 1.326 1.64 ;
    LAYER M1 ;
      RECT 0.294 0.7 0.354 1.01 ;
    LAYER M1 ;
      RECT 0.294 1.06 0.354 1.19 ;
    LAYER M1 ;
      RECT 0.294 1.33 0.354 1.64 ;
    LAYER M1 ;
      RECT 0.294 1.69 0.354 1.82 ;
    LAYER M1 ;
      RECT 0.51 0.7 0.57 1.01 ;
    LAYER M1 ;
      RECT 0.51 1.06 0.57 1.19 ;
    LAYER M1 ;
      RECT 0.51 1.33 0.57 1.64 ;
    LAYER M1 ;
      RECT 0.51 1.69 0.57 1.82 ;
    LAYER M1 ;
      RECT 0.942 0.7 1.002 1.01 ;
    LAYER M1 ;
      RECT 0.942 1.06 1.002 1.19 ;
    LAYER M1 ;
      RECT 0.942 1.33 1.002 1.64 ;
    LAYER M1 ;
      RECT 0.942 1.69 1.002 1.82 ;
    LAYER M1 ;
      RECT 1.158 0.7 1.218 1.01 ;
    LAYER M1 ;
      RECT 1.158 1.06 1.218 1.19 ;
    LAYER M1 ;
      RECT 1.158 1.33 1.218 1.64 ;
    LAYER M1 ;
      RECT 1.158 1.69 1.218 1.82 ;
    LAYER M2 ;
      RECT 0.186 0.34 1.326 0.38 ;
    LAYER M2 ;
      RECT 0.186 0.97 1.326 1.01 ;
    LAYER M2 ;
      RECT 0.186 1.6 1.326 1.64 ;
    LAYER M2 ;
      RECT 0.186 0.16 1.326 0.2 ;
    LAYER M2 ;
      RECT 0.186 0.97 1.326 1.01 ;
    LAYER M2 ;
      RECT 0.186 1.6 1.326 1.64 ;
    LAYER M2 ;
      RECT 0.2352 0.92 0.9744 0.952 ;
    LAYER M2 ;
      RECT 0.2352 2.072 0.9744 2.104 ;
    LAYER M2 ;
      RECT 0.2352 0.92 0.9744 0.952 ;
    LAYER M2 ;
      RECT 0.1488 0.632 1.0608 0.664 ;
    LAYER M2 ;
      RECT 0.1488 0.272 1.0608 0.304 ;
    LAYER M2 ;
      RECT 0.1488 1.28 1.0608 1.312 ;
    LAYER M2 ;
      RECT 0.1488 2.36 1.0608 2.392 ;
    LAYER M2 ;
      RECT 0.1488 1.856 1.0608 1.888 ;
    LAYER M2 ;
      RECT 0.2352 2.072 0.9744 2.104 ;
    LAYER M2 ;
      RECT 0.2352 1.568 0.9744 1.6 ;
    LAYER M2 ;
      RECT 0.1488 2.864 1.0608 2.896 ;
    LAYER M2 ;
      RECT 0.1488 2.216 1.0608 2.248 ;
    LAYER M2 ;
      RECT 0.1488 1.712 1.0608 1.744 ;
    LAYER M2 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER M2 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER M2 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER M2 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER V1 ;
      RECT 0.186 0.34 0.246 0.38 ;
    LAYER V1 ;
      RECT 0.186 0.97 0.246 1.01 ;
    LAYER V1 ;
      RECT 0.186 1.6 0.246 1.64 ;
    LAYER V1 ;
      RECT 0.402 0.34 0.462 0.38 ;
    LAYER V1 ;
      RECT 0.402 0.97 0.462 1.01 ;
    LAYER V1 ;
      RECT 0.402 1.6 0.462 1.64 ;
    LAYER V1 ;
      RECT 0.618 0.34 0.678 0.38 ;
    LAYER V1 ;
      RECT 0.618 0.97 0.678 1.01 ;
    LAYER V1 ;
      RECT 0.618 1.6 0.678 1.64 ;
    LAYER V1 ;
      RECT 0.834 0.34 0.894 0.38 ;
    LAYER V1 ;
      RECT 0.834 0.97 0.894 1.01 ;
    LAYER V1 ;
      RECT 0.834 1.6 0.894 1.64 ;
    LAYER V1 ;
      RECT 1.05 0.34 1.11 0.38 ;
    LAYER V1 ;
      RECT 1.05 0.97 1.11 1.01 ;
    LAYER V1 ;
      RECT 1.05 1.6 1.11 1.64 ;
    LAYER V1 ;
      RECT 1.266 0.34 1.326 0.38 ;
    LAYER V1 ;
      RECT 1.266 0.97 1.326 1.01 ;
    LAYER V1 ;
      RECT 1.266 1.6 1.326 1.64 ;
    LAYER V1 ;
      RECT 0.294 0.79 0.354 0.83 ;
    LAYER V1 ;
      RECT 0.294 1.15 0.354 1.19 ;
    LAYER V1 ;
      RECT 0.294 1.42 0.354 1.46 ;
    LAYER V1 ;
      RECT 0.294 1.78 0.354 1.82 ;
    LAYER V1 ;
      RECT 0.51 0.79 0.57 0.83 ;
    LAYER V1 ;
      RECT 0.51 1.15 0.57 1.19 ;
    LAYER V1 ;
      RECT 0.51 1.42 0.57 1.46 ;
    LAYER V1 ;
      RECT 0.51 1.78 0.57 1.82 ;
    LAYER V1 ;
      RECT 0.942 0.79 1.002 0.83 ;
    LAYER V1 ;
      RECT 0.942 1.15 1.002 1.19 ;
    LAYER V1 ;
      RECT 0.942 1.42 1.002 1.46 ;
    LAYER V1 ;
      RECT 0.942 1.78 1.002 1.82 ;
    LAYER V1 ;
      RECT 1.158 0.79 1.218 0.83 ;
    LAYER V1 ;
      RECT 1.158 1.15 1.218 1.19 ;
    LAYER V1 ;
      RECT 1.158 1.42 1.218 1.46 ;
    LAYER V1 ;
      RECT 1.158 1.78 1.218 1.82 ;
    LAYER V1 ;
      RECT 0.186 0.16 0.246 0.2 ;
    LAYER V1 ;
      RECT 0.186 0.97 0.246 1.01 ;
    LAYER V1 ;
      RECT 0.186 1.6 0.246 1.64 ;
    LAYER V1 ;
      RECT 0.402 0.16 0.462 0.2 ;
    LAYER V1 ;
      RECT 0.402 0.97 0.462 1.01 ;
    LAYER V1 ;
      RECT 0.402 1.6 0.462 1.64 ;
    LAYER V1 ;
      RECT 0.618 0.16 0.678 0.2 ;
    LAYER V1 ;
      RECT 0.618 0.97 0.678 1.01 ;
    LAYER V1 ;
      RECT 0.618 1.6 0.678 1.64 ;
    LAYER V1 ;
      RECT 0.834 0.16 0.894 0.2 ;
    LAYER V1 ;
      RECT 0.834 0.97 0.894 1.01 ;
    LAYER V1 ;
      RECT 0.834 1.6 0.894 1.64 ;
    LAYER V1 ;
      RECT 1.05 0.16 1.11 0.2 ;
    LAYER V1 ;
      RECT 1.05 0.97 1.11 1.01 ;
    LAYER V1 ;
      RECT 1.05 1.6 1.11 1.64 ;
    LAYER V1 ;
      RECT 1.266 0.16 1.326 0.2 ;
    LAYER V1 ;
      RECT 1.266 0.97 1.326 1.01 ;
    LAYER V1 ;
      RECT 1.266 1.6 1.326 1.64 ;
    LAYER V1 ;
      RECT 0.294 0.79 0.354 0.83 ;
    LAYER V1 ;
      RECT 0.294 1.15 0.354 1.19 ;
    LAYER V1 ;
      RECT 0.294 1.42 0.354 1.46 ;
    LAYER V1 ;
      RECT 0.294 1.78 0.354 1.82 ;
    LAYER V1 ;
      RECT 0.51 0.79 0.57 0.83 ;
    LAYER V1 ;
      RECT 0.51 1.15 0.57 1.19 ;
    LAYER V1 ;
      RECT 0.51 1.42 0.57 1.46 ;
    LAYER V1 ;
      RECT 0.51 1.78 0.57 1.82 ;
    LAYER V1 ;
      RECT 0.942 0.79 1.002 0.83 ;
    LAYER V1 ;
      RECT 0.942 1.15 1.002 1.19 ;
    LAYER V1 ;
      RECT 0.942 1.42 1.002 1.46 ;
    LAYER V1 ;
      RECT 0.942 1.78 1.002 1.82 ;
    LAYER V1 ;
      RECT 1.158 0.79 1.218 0.83 ;
    LAYER V1 ;
      RECT 1.158 1.15 1.218 1.19 ;
    LAYER V1 ;
      RECT 1.158 1.42 1.218 1.46 ;
    LAYER V1 ;
      RECT 1.158 1.78 1.218 1.82 ;
    LAYER Bbox ;
      RECT 0 0 1.512 1.89 ;
    LAYER Bbox ;
      RECT 0 0 1.512 1.89 ;
    LAYER M3 ;
      RECT 0.618 0.79 0.678 1.46 ;
    LAYER M3 ;
      RECT 0.726 1.15 0.786 1.82 ;
    LAYER M3 ;
      RECT 0.4944 1.856 0.5424 2.392 ;
    LAYER M3 ;
      RECT 0.1859 1.8899 0.2459 2.1599 ;
    LAYER M3 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER M3 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER M3 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER M3 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER M3 ;
      RECT 0.1859 0.9899 0.2459 1.2599 ;
    LAYER M3 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER M3 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER M3 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER M3 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER V2 ;
      RECT 0.726 1.15 0.786 1.19 ;
    LAYER V2 ;
      RECT 0.726 1.78 0.786 1.82 ;
    LAYER V2 ;
      RECT 0.618 0.79 0.678 0.83 ;
    LAYER V2 ;
      RECT 0.618 1.42 0.678 1.46 ;
    LAYER V2 ;
      RECT 0.6179 1.7799 0.6779 1.8199 ;
    LAYER V2 ;
      RECT 0.6179 1.7799 0.6779 1.8199 ;
    LAYER V2 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER V2 ;
      RECT 0.1859 2.1399 0.2459 2.1799 ;
    LAYER V2 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER V2 ;
      RECT 0.1859 0.9699 0.2459 1.0099 ;
    LAYER V3 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER V3 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER V3 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER V3 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER M4 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER M4 ;
      RECT 0.1859 1.8699 0.2459 1.9099 ;
    LAYER M4 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER M4 ;
      RECT 0.1859 1.2399 0.2459 1.2799 ;
    LAYER M4 ;
      RECT -0.0199 -0.0199 0.8839 0.0199 ;
    LAYER M4 ;
      RECT -0.0199 1.2399 0.8839 1.2799 ;
    LAYER M4 ;
      RECT -0.0199 2.4999 0.8839 2.5399 ;
    LAYER M4 ;
      RECT -0.0199 3.7599 0.8839 3.7999 ;
    LAYER M4 ;
      RECT 0.8339 -0.0199 0.8939 0.0199 ;
    LAYER M4 ;
      RECT 0.8339 1.2399 0.8939 1.2799 ;
    LAYER M4 ;
      RECT 0.8339 2.4999 0.8939 2.5399 ;
    LAYER M4 ;
      RECT 0.8339 3.7599 0.8939 3.7999 ;
    LAYER M4 ;
      RECT -0.0199 0.6099 0.8839 0.6499 ;
    LAYER M4 ;
      RECT -0.0199 1.8699 0.8839 1.9099 ;
    LAYER M4 ;
      RECT -0.0199 3.1299 0.8839 3.1699 ;
    LAYER M4 ;
      RECT -0.0299 0.6099 0.0299 0.6499 ;
    LAYER M4 ;
      RECT -0.0299 1.8699 0.0299 1.9099 ;
    LAYER M4 ;
      RECT -0.0299 3.1299 0.0299 3.1699 ;
    LAYER M5 ;
      RECT 0.8339 -0.0299 0.8939 0.6599 ;
    LAYER M5 ;
      RECT 0.8339 0.5999 0.8939 1.2899 ;
    LAYER M5 ;
      RECT 0.8339 1.2299 0.8939 1.9199 ;
    LAYER M5 ;
      RECT 0.8339 1.8599 0.8939 2.5499 ;
    LAYER M5 ;
      RECT 0.8339 2.4899 0.8939 3.1799 ;
    LAYER M5 ;
      RECT 0.8339 3.1199 0.8939 3.8099 ;
    LAYER M5 ;
      RECT 0.8339 -0.0199 0.8939 0.0199 ;
    LAYER M5 ;
      RECT 0.8339 1.2399 0.8939 1.2799 ;
    LAYER M5 ;
      RECT 0.8339 2.4999 0.8939 2.5399 ;
    LAYER M5 ;
      RECT 0.8339 3.7599 0.8939 3.7999 ;
    LAYER M5 ;
      RECT -0.0299 -0.0299 0.0299 0.6599 ;
    LAYER M5 ;
      RECT -0.0299 0.5999 0.0299 1.2899 ;
    LAYER M5 ;
      RECT -0.0299 1.2299 0.0299 1.9199 ;
    LAYER M5 ;
      RECT -0.0299 1.8599 0.0299 2.5499 ;
    LAYER M5 ;
      RECT -0.0299 2.4899 0.0299 3.1799 ;
    LAYER M5 ;
      RECT -0.0299 3.1199 0.0299 3.8099 ;
    LAYER M5 ;
      RECT -0.0299 0.6099 0.0299 0.6499 ;
    LAYER M5 ;
      RECT -0.0299 1.8699 0.0299 1.9099 ;
    LAYER M5 ;
      RECT -0.0299 3.1299 0.0299 3.1699 ;
    LAYER V4 ;
      RECT 0.8339 -0.0199 0.8939 0.0199 ;
    LAYER V4 ;
      RECT 0.8339 1.2399 0.8939 1.2799 ;
    LAYER V4 ;
      RECT 0.8339 2.4999 0.8939 2.5399 ;
    LAYER V4 ;
      RECT 0.8339 3.7599 0.8939 3.7999 ;
    LAYER V4 ;
      RECT -0.0299 0.6099 0.0299 0.6499 ;
    LAYER V4 ;
      RECT -0.0299 1.8699 0.0299 1.9099 ;
    LAYER V4 ;
      RECT -0.0299 3.1299 0.0299 3.1699 ;
  END
END CKT_OBS_LEF
