MACRO Switch_NMOS_n12_X3_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y2 0 0 ;
  SIZE 1.296 BY 1.080 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.040 0.099 1.148 0.117 ;
      LAYER M2 ;
        RECT 0.040 0.153 1.148 0.171 ;
      LAYER M2 ;
        RECT 0.040 0.207 1.148 0.225 ;
      LAYER M2 ;
        RECT 0.040 0.639 1.148 0.657 ;
      LAYER M2 ;
        RECT 0.040 0.693 1.148 0.711 ;
      LAYER M2 ;
        RECT 0.040 0.747 1.148 0.765 ;
      LAYER M3 ;
        RECT 0.585 0.094 0.603 0.770 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.261 1.256 0.279 ;
      LAYER M2 ;
        RECT 0.148 0.801 1.256 0.819 ;
      LAYER M3 ;
        RECT 0.639 0.256 0.657 0.824 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.315 1.202 0.333 ;
      LAYER M2 ;
        RECT 0.094 0.855 1.202 0.873 ;
      LAYER M3 ;
        RECT 0.531 0.310 0.549 0.878 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.099 0.580 0.117 1.040 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.580 0.333 1.040 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.580 0.549 1.040 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.580 0.765 1.040 ;
    LAYER M1 ;
      RECT 0.963 0.040 0.981 0.500 ;
    LAYER M1 ;
      RECT 0.963 0.580 0.981 1.040 ;
    LAYER M1 ;
      RECT 1.179 0.040 1.197 0.500 ;
    LAYER M1 ;
      RECT 1.179 0.580 1.197 1.040 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.580 0.063 1.040 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.580 0.279 1.040 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.580 0.495 1.040 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.580 0.711 1.040 ;
    LAYER M1 ;
      RECT 0.909 0.040 0.927 0.500 ;
    LAYER M1 ;
      RECT 0.909 0.580 0.927 1.040 ;
    LAYER M1 ;
      RECT 1.125 0.040 1.143 0.500 ;
    LAYER M1 ;
      RECT 1.125 0.580 1.143 1.040 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.580 0.171 1.040 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.580 0.387 1.040 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.580 0.603 1.040 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.580 0.819 1.040 ;
    LAYER M1 ;
      RECT 1.017 0.040 1.035 0.500 ;
    LAYER M1 ;
      RECT 1.017 0.580 1.035 1.040 ;
    LAYER M1 ;
      RECT 1.233 0.040 1.251 0.500 ;
    LAYER M1 ;
      RECT 1.233 0.580 1.251 1.040 ;
  END
END Switch_NMOS_n12_X3_Y2
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.432 BY 0.540 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.040 0.099 0.284 0.117 ;
      LAYER M2 ;
        RECT 0.040 0.153 0.284 0.171 ;
      LAYER M2 ;
        RECT 0.040 0.207 0.284 0.225 ;
      LAYER M3 ;
        RECT 0.153 0.094 0.171 0.446 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.261 0.392 0.279 ;
      LAYER M3 ;
        RECT 0.207 0.094 0.225 0.446 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.315 0.338 0.333 ;
      LAYER M3 ;
        RECT 0.099 0.094 0.117 0.446 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X3_Y1 0 0 ;
  SIZE 1.296 BY 0.540 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.040 0.099 1.148 0.117 ;
      LAYER M2 ;
        RECT 0.040 0.153 1.148 0.171 ;
      LAYER M2 ;
        RECT 0.040 0.207 1.148 0.225 ;
      LAYER M3 ;
        RECT 0.585 0.094 0.603 0.446 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.261 1.256 0.279 ;
      LAYER M3 ;
        RECT 0.639 0.094 0.657 0.446 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.315 1.202 0.333 ;
      LAYER M3 ;
        RECT 0.531 0.094 0.549 0.446 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.963 0.040 0.981 0.500 ;
    LAYER M1 ;
      RECT 1.179 0.040 1.197 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.909 0.040 0.927 0.500 ;
    LAYER M1 ;
      RECT 1.125 0.040 1.143 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 1.017 0.040 1.035 0.500 ;
    LAYER M1 ;
      RECT 1.233 0.040 1.251 0.500 ;
  END
END Switch_PMOS_n12_X3_Y1
