MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 11.68 BY 15.708 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 15.42 3.136 15.492 ;
      LAYER M2 ;
        RECT 3.084 15.44 3.156 15.472 ;
      LAYER M1 ;
        RECT 8.864 15.42 8.896 15.492 ;
      LAYER M2 ;
        RECT 8.844 15.44 8.916 15.472 ;
      LAYER M2 ;
        RECT 3.12 15.44 8.88 15.472 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
      LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.664 6.6 5.696 6.672 ;
  LAYER M2 ;
        RECT 5.644 6.62 5.716 6.652 ;
  LAYER M1 ;
        RECT 5.664 6.468 5.696 6.636 ;
  LAYER M1 ;
        RECT 5.664 6.432 5.696 6.504 ;
  LAYER M2 ;
        RECT 5.644 6.452 5.716 6.484 ;
  LAYER M2 ;
        RECT 5.68 6.452 5.84 6.484 ;
  LAYER M1 ;
        RECT 5.824 6.432 5.856 6.504 ;
  LAYER M2 ;
        RECT 5.804 6.452 5.876 6.484 ;
  LAYER M1 ;
        RECT 8.544 6.6 8.576 6.672 ;
  LAYER M2 ;
        RECT 8.524 6.62 8.596 6.652 ;
  LAYER M2 ;
        RECT 5.84 6.62 8.56 6.652 ;
  LAYER M1 ;
        RECT 5.824 6.6 5.856 6.672 ;
  LAYER M2 ;
        RECT 5.804 6.62 5.876 6.652 ;
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M1 ;
        RECT 5.664 9.408 5.696 9.576 ;
  LAYER M1 ;
        RECT 5.664 9.372 5.696 9.444 ;
  LAYER M2 ;
        RECT 5.644 9.392 5.716 9.424 ;
  LAYER M2 ;
        RECT 5.68 9.392 5.84 9.424 ;
  LAYER M1 ;
        RECT 5.824 9.372 5.856 9.444 ;
  LAYER M2 ;
        RECT 5.804 9.392 5.876 9.424 ;
  LAYER M1 ;
        RECT 8.544 3.66 8.576 3.732 ;
  LAYER M2 ;
        RECT 8.524 3.68 8.596 3.712 ;
  LAYER M2 ;
        RECT 5.84 3.68 8.56 3.712 ;
  LAYER M1 ;
        RECT 5.824 3.66 5.856 3.732 ;
  LAYER M2 ;
        RECT 5.804 3.68 5.876 3.712 ;
  LAYER M1 ;
        RECT 5.664 3.66 5.696 3.732 ;
  LAYER M2 ;
        RECT 5.644 3.68 5.716 3.712 ;
  LAYER M1 ;
        RECT 5.664 3.528 5.696 3.696 ;
  LAYER M1 ;
        RECT 5.664 3.492 5.696 3.564 ;
  LAYER M2 ;
        RECT 5.644 3.512 5.716 3.544 ;
  LAYER M2 ;
        RECT 5.68 3.512 5.84 3.544 ;
  LAYER M1 ;
        RECT 5.824 3.492 5.856 3.564 ;
  LAYER M2 ;
        RECT 5.804 3.512 5.876 3.544 ;
  LAYER M1 ;
        RECT 8.544 9.54 8.576 9.612 ;
  LAYER M2 ;
        RECT 8.524 9.56 8.596 9.592 ;
  LAYER M2 ;
        RECT 5.84 9.56 8.56 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
  LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
  LAYER M1 ;
        RECT 5.824 0.252 5.856 0.42 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 9.576 ;
  LAYER M1 ;
        RECT 2.784 0.72 2.816 0.792 ;
  LAYER M2 ;
        RECT 2.764 0.74 2.836 0.772 ;
  LAYER M1 ;
        RECT 2.784 0.588 2.816 0.756 ;
  LAYER M1 ;
        RECT 2.784 0.552 2.816 0.624 ;
  LAYER M2 ;
        RECT 2.764 0.572 2.836 0.604 ;
  LAYER M2 ;
        RECT 2.8 0.572 2.96 0.604 ;
  LAYER M1 ;
        RECT 2.944 0.552 2.976 0.624 ;
  LAYER M2 ;
        RECT 2.924 0.572 2.996 0.604 ;
  LAYER M1 ;
        RECT 2.784 3.66 2.816 3.732 ;
  LAYER M2 ;
        RECT 2.764 3.68 2.836 3.712 ;
  LAYER M1 ;
        RECT 2.784 3.528 2.816 3.696 ;
  LAYER M1 ;
        RECT 2.784 3.492 2.816 3.564 ;
  LAYER M2 ;
        RECT 2.764 3.512 2.836 3.544 ;
  LAYER M2 ;
        RECT 2.8 3.512 2.96 3.544 ;
  LAYER M1 ;
        RECT 2.944 3.492 2.976 3.564 ;
  LAYER M2 ;
        RECT 2.924 3.512 2.996 3.544 ;
  LAYER M1 ;
        RECT 2.784 6.6 2.816 6.672 ;
  LAYER M2 ;
        RECT 2.764 6.62 2.836 6.652 ;
  LAYER M1 ;
        RECT 2.784 6.468 2.816 6.636 ;
  LAYER M1 ;
        RECT 2.784 6.432 2.816 6.504 ;
  LAYER M2 ;
        RECT 2.764 6.452 2.836 6.484 ;
  LAYER M2 ;
        RECT 2.8 6.452 2.96 6.484 ;
  LAYER M1 ;
        RECT 2.944 6.432 2.976 6.504 ;
  LAYER M2 ;
        RECT 2.924 6.452 2.996 6.484 ;
  LAYER M1 ;
        RECT 2.784 9.54 2.816 9.612 ;
  LAYER M2 ;
        RECT 2.764 9.56 2.836 9.592 ;
  LAYER M1 ;
        RECT 2.784 9.408 2.816 9.576 ;
  LAYER M1 ;
        RECT 2.784 9.372 2.816 9.444 ;
  LAYER M2 ;
        RECT 2.764 9.392 2.836 9.424 ;
  LAYER M2 ;
        RECT 2.8 9.392 2.96 9.424 ;
  LAYER M1 ;
        RECT 2.944 9.372 2.976 9.444 ;
  LAYER M2 ;
        RECT 2.924 9.392 2.996 9.424 ;
  LAYER M1 ;
        RECT 2.784 12.48 2.816 12.552 ;
  LAYER M2 ;
        RECT 2.764 12.5 2.836 12.532 ;
  LAYER M1 ;
        RECT 2.784 12.348 2.816 12.516 ;
  LAYER M1 ;
        RECT 2.784 12.312 2.816 12.384 ;
  LAYER M2 ;
        RECT 2.764 12.332 2.836 12.364 ;
  LAYER M2 ;
        RECT 2.8 12.332 2.96 12.364 ;
  LAYER M1 ;
        RECT 2.944 12.312 2.976 12.384 ;
  LAYER M2 ;
        RECT 2.924 12.332 2.996 12.364 ;
  LAYER M1 ;
        RECT 5.664 0.72 5.696 0.792 ;
  LAYER M2 ;
        RECT 5.644 0.74 5.716 0.772 ;
  LAYER M2 ;
        RECT 2.96 0.74 5.68 0.772 ;
  LAYER M1 ;
        RECT 2.944 0.72 2.976 0.792 ;
  LAYER M2 ;
        RECT 2.924 0.74 2.996 0.772 ;
  LAYER M1 ;
        RECT 5.664 12.48 5.696 12.552 ;
  LAYER M2 ;
        RECT 5.644 12.5 5.716 12.532 ;
  LAYER M2 ;
        RECT 2.96 12.5 5.68 12.532 ;
  LAYER M1 ;
        RECT 2.944 12.48 2.976 12.552 ;
  LAYER M2 ;
        RECT 2.924 12.5 2.996 12.532 ;
  LAYER M1 ;
        RECT 2.944 0.048 2.976 0.12 ;
  LAYER M2 ;
        RECT 2.924 0.068 2.996 0.1 ;
  LAYER M1 ;
        RECT 2.944 0.084 2.976 0.42 ;
  LAYER M1 ;
        RECT 2.944 0.42 2.976 12.516 ;
  LAYER M1 ;
        RECT 8.544 0.72 8.576 0.792 ;
  LAYER M2 ;
        RECT 8.524 0.74 8.596 0.772 ;
  LAYER M1 ;
        RECT 8.544 0.588 8.576 0.756 ;
  LAYER M1 ;
        RECT 8.544 0.552 8.576 0.624 ;
  LAYER M2 ;
        RECT 8.524 0.572 8.596 0.604 ;
  LAYER M2 ;
        RECT 8.56 0.572 8.72 0.604 ;
  LAYER M1 ;
        RECT 8.704 0.552 8.736 0.624 ;
  LAYER M2 ;
        RECT 8.684 0.572 8.756 0.604 ;
  LAYER M1 ;
        RECT 8.544 12.48 8.576 12.552 ;
  LAYER M2 ;
        RECT 8.524 12.5 8.596 12.532 ;
  LAYER M1 ;
        RECT 8.544 12.348 8.576 12.516 ;
  LAYER M1 ;
        RECT 8.544 12.312 8.576 12.384 ;
  LAYER M2 ;
        RECT 8.524 12.332 8.596 12.364 ;
  LAYER M2 ;
        RECT 8.56 12.332 8.72 12.364 ;
  LAYER M1 ;
        RECT 8.704 12.312 8.736 12.384 ;
  LAYER M2 ;
        RECT 8.684 12.332 8.756 12.364 ;
  LAYER M1 ;
        RECT 11.424 0.72 11.456 0.792 ;
  LAYER M2 ;
        RECT 11.404 0.74 11.476 0.772 ;
  LAYER M2 ;
        RECT 8.72 0.74 11.44 0.772 ;
  LAYER M1 ;
        RECT 8.704 0.72 8.736 0.792 ;
  LAYER M2 ;
        RECT 8.684 0.74 8.756 0.772 ;
  LAYER M1 ;
        RECT 11.424 3.66 11.456 3.732 ;
  LAYER M2 ;
        RECT 11.404 3.68 11.476 3.712 ;
  LAYER M2 ;
        RECT 8.72 3.68 11.44 3.712 ;
  LAYER M1 ;
        RECT 8.704 3.66 8.736 3.732 ;
  LAYER M2 ;
        RECT 8.684 3.68 8.756 3.712 ;
  LAYER M1 ;
        RECT 11.424 6.6 11.456 6.672 ;
  LAYER M2 ;
        RECT 11.404 6.62 11.476 6.652 ;
  LAYER M2 ;
        RECT 8.72 6.62 11.44 6.652 ;
  LAYER M1 ;
        RECT 8.704 6.6 8.736 6.672 ;
  LAYER M2 ;
        RECT 8.684 6.62 8.756 6.652 ;
  LAYER M1 ;
        RECT 11.424 9.54 11.456 9.612 ;
  LAYER M2 ;
        RECT 11.404 9.56 11.476 9.592 ;
  LAYER M2 ;
        RECT 8.72 9.56 11.44 9.592 ;
  LAYER M1 ;
        RECT 8.704 9.54 8.736 9.612 ;
  LAYER M2 ;
        RECT 8.684 9.56 8.756 9.592 ;
  LAYER M1 ;
        RECT 11.424 12.48 11.456 12.552 ;
  LAYER M2 ;
        RECT 11.404 12.5 11.476 12.532 ;
  LAYER M2 ;
        RECT 8.72 12.5 11.44 12.532 ;
  LAYER M1 ;
        RECT 8.704 12.48 8.736 12.552 ;
  LAYER M2 ;
        RECT 8.684 12.5 8.756 12.532 ;
  LAYER M1 ;
        RECT 8.704 0.048 8.736 0.12 ;
  LAYER M2 ;
        RECT 8.684 0.068 8.756 0.1 ;
  LAYER M1 ;
        RECT 8.704 0.084 8.736 0.42 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 12.516 ;
  LAYER M2 ;
        RECT 2.96 0.068 8.72 0.1 ;
  LAYER M1 ;
        RECT 3.264 9.036 3.296 9.108 ;
  LAYER M2 ;
        RECT 3.244 9.056 3.316 9.088 ;
  LAYER M2 ;
        RECT 3.12 9.056 3.28 9.088 ;
  LAYER M1 ;
        RECT 3.104 9.036 3.136 9.108 ;
  LAYER M2 ;
        RECT 3.084 9.056 3.156 9.088 ;
  LAYER M1 ;
        RECT 3.264 11.976 3.296 12.048 ;
  LAYER M2 ;
        RECT 3.244 11.996 3.316 12.028 ;
  LAYER M2 ;
        RECT 3.12 11.996 3.28 12.028 ;
  LAYER M1 ;
        RECT 3.104 11.976 3.136 12.048 ;
  LAYER M2 ;
        RECT 3.084 11.996 3.156 12.028 ;
  LAYER M1 ;
        RECT 3.264 6.096 3.296 6.168 ;
  LAYER M2 ;
        RECT 3.244 6.116 3.316 6.148 ;
  LAYER M2 ;
        RECT 3.12 6.116 3.28 6.148 ;
  LAYER M1 ;
        RECT 3.104 6.096 3.136 6.168 ;
  LAYER M2 ;
        RECT 3.084 6.116 3.156 6.148 ;
  LAYER M1 ;
        RECT 3.104 15.42 3.136 15.492 ;
  LAYER M2 ;
        RECT 3.084 15.44 3.156 15.472 ;
  LAYER M1 ;
        RECT 3.104 15.288 3.136 15.456 ;
  LAYER M1 ;
        RECT 3.104 6.132 3.136 15.288 ;
  LAYER M1 ;
        RECT 6.144 9.036 6.176 9.108 ;
  LAYER M2 ;
        RECT 6.124 9.056 6.196 9.088 ;
  LAYER M1 ;
        RECT 6.144 9.072 6.176 9.24 ;
  LAYER M1 ;
        RECT 6.144 9.204 6.176 9.276 ;
  LAYER M2 ;
        RECT 6.124 9.224 6.196 9.256 ;
  LAYER M2 ;
        RECT 6.16 9.224 8.88 9.256 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M1 ;
        RECT 6.144 6.096 6.176 6.168 ;
  LAYER M2 ;
        RECT 6.124 6.116 6.196 6.148 ;
  LAYER M1 ;
        RECT 6.144 6.132 6.176 6.3 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M2 ;
        RECT 6.16 6.284 8.88 6.316 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M1 ;
        RECT 6.144 11.976 6.176 12.048 ;
  LAYER M2 ;
        RECT 6.124 11.996 6.196 12.028 ;
  LAYER M1 ;
        RECT 6.144 12.012 6.176 12.18 ;
  LAYER M1 ;
        RECT 6.144 12.144 6.176 12.216 ;
  LAYER M2 ;
        RECT 6.124 12.164 6.196 12.196 ;
  LAYER M2 ;
        RECT 6.16 12.164 8.88 12.196 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M1 ;
        RECT 8.864 15.42 8.896 15.492 ;
  LAYER M2 ;
        RECT 8.844 15.44 8.916 15.472 ;
  LAYER M1 ;
        RECT 8.864 15.288 8.896 15.456 ;
  LAYER M1 ;
        RECT 8.864 6.3 8.896 15.288 ;
  LAYER M2 ;
        RECT 3.12 15.44 8.88 15.472 ;
  LAYER M1 ;
        RECT 0.384 3.156 0.416 3.228 ;
  LAYER M2 ;
        RECT 0.364 3.176 0.436 3.208 ;
  LAYER M2 ;
        RECT 0.08 3.176 0.4 3.208 ;
  LAYER M1 ;
        RECT 0.064 3.156 0.096 3.228 ;
  LAYER M2 ;
        RECT 0.044 3.176 0.116 3.208 ;
  LAYER M1 ;
        RECT 0.384 6.096 0.416 6.168 ;
  LAYER M2 ;
        RECT 0.364 6.116 0.436 6.148 ;
  LAYER M2 ;
        RECT 0.08 6.116 0.4 6.148 ;
  LAYER M1 ;
        RECT 0.064 6.096 0.096 6.168 ;
  LAYER M2 ;
        RECT 0.044 6.116 0.116 6.148 ;
  LAYER M1 ;
        RECT 0.384 9.036 0.416 9.108 ;
  LAYER M2 ;
        RECT 0.364 9.056 0.436 9.088 ;
  LAYER M2 ;
        RECT 0.08 9.056 0.4 9.088 ;
  LAYER M1 ;
        RECT 0.064 9.036 0.096 9.108 ;
  LAYER M2 ;
        RECT 0.044 9.056 0.116 9.088 ;
  LAYER M1 ;
        RECT 0.384 11.976 0.416 12.048 ;
  LAYER M2 ;
        RECT 0.364 11.996 0.436 12.028 ;
  LAYER M2 ;
        RECT 0.08 11.996 0.4 12.028 ;
  LAYER M1 ;
        RECT 0.064 11.976 0.096 12.048 ;
  LAYER M2 ;
        RECT 0.044 11.996 0.116 12.028 ;
  LAYER M1 ;
        RECT 0.384 14.916 0.416 14.988 ;
  LAYER M2 ;
        RECT 0.364 14.936 0.436 14.968 ;
  LAYER M2 ;
        RECT 0.08 14.936 0.4 14.968 ;
  LAYER M1 ;
        RECT 0.064 14.916 0.096 14.988 ;
  LAYER M2 ;
        RECT 0.044 14.936 0.116 14.968 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.288 0.096 15.624 ;
  LAYER M1 ;
        RECT 0.064 3.192 0.096 15.288 ;
  LAYER M1 ;
        RECT 9.024 3.156 9.056 3.228 ;
  LAYER M2 ;
        RECT 9.004 3.176 9.076 3.208 ;
  LAYER M1 ;
        RECT 9.024 3.192 9.056 3.36 ;
  LAYER M1 ;
        RECT 9.024 3.324 9.056 3.396 ;
  LAYER M2 ;
        RECT 9.004 3.344 9.076 3.376 ;
  LAYER M2 ;
        RECT 9.04 3.344 11.6 3.376 ;
  LAYER M1 ;
        RECT 11.584 3.324 11.616 3.396 ;
  LAYER M2 ;
        RECT 11.564 3.344 11.636 3.376 ;
  LAYER M1 ;
        RECT 9.024 6.096 9.056 6.168 ;
  LAYER M2 ;
        RECT 9.004 6.116 9.076 6.148 ;
  LAYER M1 ;
        RECT 9.024 6.132 9.056 6.3 ;
  LAYER M1 ;
        RECT 9.024 6.264 9.056 6.336 ;
  LAYER M2 ;
        RECT 9.004 6.284 9.076 6.316 ;
  LAYER M2 ;
        RECT 9.04 6.284 11.6 6.316 ;
  LAYER M1 ;
        RECT 11.584 6.264 11.616 6.336 ;
  LAYER M2 ;
        RECT 11.564 6.284 11.636 6.316 ;
  LAYER M1 ;
        RECT 9.024 9.036 9.056 9.108 ;
  LAYER M2 ;
        RECT 9.004 9.056 9.076 9.088 ;
  LAYER M1 ;
        RECT 9.024 9.072 9.056 9.24 ;
  LAYER M1 ;
        RECT 9.024 9.204 9.056 9.276 ;
  LAYER M2 ;
        RECT 9.004 9.224 9.076 9.256 ;
  LAYER M2 ;
        RECT 9.04 9.224 11.6 9.256 ;
  LAYER M1 ;
        RECT 11.584 9.204 11.616 9.276 ;
  LAYER M2 ;
        RECT 11.564 9.224 11.636 9.256 ;
  LAYER M1 ;
        RECT 9.024 11.976 9.056 12.048 ;
  LAYER M2 ;
        RECT 9.004 11.996 9.076 12.028 ;
  LAYER M1 ;
        RECT 9.024 12.012 9.056 12.18 ;
  LAYER M1 ;
        RECT 9.024 12.144 9.056 12.216 ;
  LAYER M2 ;
        RECT 9.004 12.164 9.076 12.196 ;
  LAYER M2 ;
        RECT 9.04 12.164 11.6 12.196 ;
  LAYER M1 ;
        RECT 11.584 12.144 11.616 12.216 ;
  LAYER M2 ;
        RECT 11.564 12.164 11.636 12.196 ;
  LAYER M1 ;
        RECT 9.024 14.916 9.056 14.988 ;
  LAYER M2 ;
        RECT 9.004 14.936 9.076 14.968 ;
  LAYER M1 ;
        RECT 9.024 14.952 9.056 15.12 ;
  LAYER M1 ;
        RECT 9.024 15.084 9.056 15.156 ;
  LAYER M2 ;
        RECT 9.004 15.104 9.076 15.136 ;
  LAYER M2 ;
        RECT 9.04 15.104 11.6 15.136 ;
  LAYER M1 ;
        RECT 11.584 15.084 11.616 15.156 ;
  LAYER M2 ;
        RECT 11.564 15.104 11.636 15.136 ;
  LAYER M1 ;
        RECT 11.584 15.588 11.616 15.66 ;
  LAYER M2 ;
        RECT 11.564 15.608 11.636 15.64 ;
  LAYER M1 ;
        RECT 11.584 15.288 11.616 15.624 ;
  LAYER M1 ;
        RECT 11.584 3.36 11.616 15.288 ;
  LAYER M2 ;
        RECT 0.08 15.608 11.6 15.64 ;
  LAYER M1 ;
        RECT 3.264 3.156 3.296 3.228 ;
  LAYER M2 ;
        RECT 3.244 3.176 3.316 3.208 ;
  LAYER M2 ;
        RECT 0.4 3.176 3.28 3.208 ;
  LAYER M1 ;
        RECT 0.384 3.156 0.416 3.228 ;
  LAYER M2 ;
        RECT 0.364 3.176 0.436 3.208 ;
  LAYER M1 ;
        RECT 3.264 14.916 3.296 14.988 ;
  LAYER M2 ;
        RECT 3.244 14.936 3.316 14.968 ;
  LAYER M2 ;
        RECT 0.4 14.936 3.28 14.968 ;
  LAYER M1 ;
        RECT 0.384 14.916 0.416 14.988 ;
  LAYER M2 ;
        RECT 0.364 14.936 0.436 14.968 ;
  LAYER M1 ;
        RECT 6.144 14.916 6.176 14.988 ;
  LAYER M2 ;
        RECT 6.124 14.936 6.196 14.968 ;
  LAYER M2 ;
        RECT 3.28 14.936 6.16 14.968 ;
  LAYER M1 ;
        RECT 3.264 14.916 3.296 14.988 ;
  LAYER M2 ;
        RECT 3.244 14.936 3.316 14.968 ;
  LAYER M1 ;
        RECT 6.144 3.156 6.176 3.228 ;
  LAYER M2 ;
        RECT 6.124 3.176 6.196 3.208 ;
  LAYER M2 ;
        RECT 6.16 3.176 9.04 3.208 ;
  LAYER M1 ;
        RECT 9.024 3.156 9.056 3.228 ;
  LAYER M2 ;
        RECT 9.004 3.176 9.076 3.208 ;
  LAYER M1 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M3 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M1 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M2 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M3 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M1 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M2 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M3 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M1 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M2 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M3 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M1 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M2 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M3 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M1 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M2 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M3 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M1 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M2 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M3 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M1 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M2 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M3 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M1 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M2 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M3 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M1 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M2 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M3 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M1 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M2 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M3 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M1 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M2 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M3 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M1 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M2 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M3 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M1 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M2 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M3 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M1 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M2 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M3 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M1 ;
        RECT 9.04 0.756 11.44 3.192 ;
  LAYER M2 ;
        RECT 9.04 0.756 11.44 3.192 ;
  LAYER M3 ;
        RECT 9.04 0.756 11.44 3.192 ;
  LAYER M1 ;
        RECT 9.04 3.696 11.44 6.132 ;
  LAYER M2 ;
        RECT 9.04 3.696 11.44 6.132 ;
  LAYER M3 ;
        RECT 9.04 3.696 11.44 6.132 ;
  LAYER M1 ;
        RECT 9.04 6.636 11.44 9.072 ;
  LAYER M2 ;
        RECT 9.04 6.636 11.44 9.072 ;
  LAYER M3 ;
        RECT 9.04 6.636 11.44 9.072 ;
  LAYER M1 ;
        RECT 9.04 9.576 11.44 12.012 ;
  LAYER M2 ;
        RECT 9.04 9.576 11.44 12.012 ;
  LAYER M3 ;
        RECT 9.04 9.576 11.44 12.012 ;
  LAYER M1 ;
        RECT 9.04 12.516 11.44 14.952 ;
  LAYER M2 ;
        RECT 9.04 12.516 11.44 14.952 ;
  LAYER M3 ;
        RECT 9.04 12.516 11.44 14.952 ;
  END 
END Cap_60fF
