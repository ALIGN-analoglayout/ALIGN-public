MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 10.16 BY 26.208 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.68 25.752 3.712 25.824 ;
      LAYER M2 ;
        RECT 3.66 25.772 3.732 25.804 ;
      LAYER M1 ;
        RECT 6.976 25.752 7.008 25.824 ;
      LAYER M2 ;
        RECT 6.956 25.772 7.028 25.804 ;
      LAYER M2 ;
        RECT 3.696 25.772 6.992 25.804 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
      LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
      LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
      LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
      LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.84 25.92 3.872 25.992 ;
      LAYER M2 ;
        RECT 3.82 25.94 3.892 25.972 ;
      LAYER M1 ;
        RECT 7.136 25.92 7.168 25.992 ;
      LAYER M2 ;
        RECT 7.116 25.94 7.188 25.972 ;
      LAYER M2 ;
        RECT 3.856 25.94 7.152 25.972 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
      LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
      LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
      LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
      LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M2 ;
        RECT 3.376 13.424 6.448 13.456 ;
  LAYER M1 ;
        RECT 3.36 13.404 3.392 13.476 ;
  LAYER M2 ;
        RECT 3.34 13.424 3.412 13.456 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M2 ;
        RECT 3.376 7.208 6.448 7.24 ;
  LAYER M1 ;
        RECT 3.36 7.188 3.392 7.26 ;
  LAYER M2 ;
        RECT 3.34 7.208 3.412 7.24 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M2 ;
        RECT 3.376 16.532 6.448 16.564 ;
  LAYER M1 ;
        RECT 3.36 16.512 3.392 16.584 ;
  LAYER M2 ;
        RECT 3.34 16.532 3.412 16.564 ;
  LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
  LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
  LAYER M1 ;
        RECT 3.36 0.42 3.392 0.672 ;
  LAYER M1 ;
        RECT 3.36 0.672 3.392 16.548 ;
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M1 ;
        RECT 6.432 13.272 6.464 13.44 ;
  LAYER M1 ;
        RECT 6.432 13.236 6.464 13.308 ;
  LAYER M2 ;
        RECT 6.412 13.256 6.484 13.288 ;
  LAYER M2 ;
        RECT 6.448 13.256 6.672 13.288 ;
  LAYER M1 ;
        RECT 6.656 13.236 6.688 13.308 ;
  LAYER M2 ;
        RECT 6.636 13.256 6.708 13.288 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M1 ;
        RECT 6.432 7.056 6.464 7.224 ;
  LAYER M1 ;
        RECT 6.432 7.02 6.464 7.092 ;
  LAYER M2 ;
        RECT 6.412 7.04 6.484 7.072 ;
  LAYER M2 ;
        RECT 6.448 7.04 6.672 7.072 ;
  LAYER M1 ;
        RECT 6.656 7.02 6.688 7.092 ;
  LAYER M2 ;
        RECT 6.636 7.04 6.708 7.072 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M1 ;
        RECT 6.432 16.38 6.464 16.548 ;
  LAYER M1 ;
        RECT 6.432 16.344 6.464 16.416 ;
  LAYER M2 ;
        RECT 6.412 16.364 6.484 16.396 ;
  LAYER M2 ;
        RECT 6.448 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 16.416 ;
  LAYER M2 ;
        RECT 6.636 16.364 6.708 16.396 ;
  LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
  LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
  LAYER M1 ;
        RECT 6.656 0.42 6.688 0.672 ;
  LAYER M1 ;
        RECT 6.656 0.672 6.688 16.38 ;
  LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M2 ;
        RECT 3.536 10.316 6.448 10.348 ;
  LAYER M1 ;
        RECT 3.52 10.296 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.5 10.316 3.572 10.348 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M2 ;
        RECT 3.536 4.1 6.448 4.132 ;
  LAYER M1 ;
        RECT 3.52 4.08 3.552 4.152 ;
  LAYER M2 ;
        RECT 3.5 4.1 3.572 4.132 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M2 ;
        RECT 3.536 19.64 6.448 19.672 ;
  LAYER M1 ;
        RECT 3.52 19.62 3.552 19.692 ;
  LAYER M2 ;
        RECT 3.5 19.64 3.572 19.672 ;
  LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
  LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
  LAYER M1 ;
        RECT 3.52 0.252 3.552 0.672 ;
  LAYER M1 ;
        RECT 3.52 0.672 3.552 19.656 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M1 ;
        RECT 6.432 10.164 6.464 10.332 ;
  LAYER M1 ;
        RECT 6.432 10.128 6.464 10.2 ;
  LAYER M2 ;
        RECT 6.412 10.148 6.484 10.18 ;
  LAYER M2 ;
        RECT 6.448 10.148 6.832 10.18 ;
  LAYER M1 ;
        RECT 6.816 10.128 6.848 10.2 ;
  LAYER M2 ;
        RECT 6.796 10.148 6.868 10.18 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M1 ;
        RECT 6.432 3.948 6.464 4.116 ;
  LAYER M1 ;
        RECT 6.432 3.912 6.464 3.984 ;
  LAYER M2 ;
        RECT 6.412 3.932 6.484 3.964 ;
  LAYER M2 ;
        RECT 6.448 3.932 6.832 3.964 ;
  LAYER M1 ;
        RECT 6.816 3.912 6.848 3.984 ;
  LAYER M2 ;
        RECT 6.796 3.932 6.868 3.964 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M1 ;
        RECT 6.432 19.488 6.464 19.656 ;
  LAYER M1 ;
        RECT 6.432 19.452 6.464 19.524 ;
  LAYER M2 ;
        RECT 6.412 19.472 6.484 19.504 ;
  LAYER M2 ;
        RECT 6.448 19.472 6.832 19.504 ;
  LAYER M1 ;
        RECT 6.816 19.452 6.848 19.524 ;
  LAYER M2 ;
        RECT 6.796 19.472 6.868 19.504 ;
  LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
  LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
  LAYER M1 ;
        RECT 6.816 0.252 6.848 0.672 ;
  LAYER M1 ;
        RECT 6.816 0.672 6.848 19.488 ;
  LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 3.152 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 3.136 4.08 3.168 4.152 ;
  LAYER M2 ;
        RECT 3.116 4.1 3.188 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 3.152 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 3.136 7.188 3.168 7.26 ;
  LAYER M2 ;
        RECT 3.116 7.208 3.188 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 3.152 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 3.136 10.296 3.168 10.368 ;
  LAYER M2 ;
        RECT 3.116 10.316 3.188 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 3.152 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 3.136 13.404 3.168 13.476 ;
  LAYER M2 ;
        RECT 3.116 13.424 3.188 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 3.152 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 3.136 16.512 3.168 16.584 ;
  LAYER M2 ;
        RECT 3.116 16.532 3.188 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 3.152 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 3.136 19.62 3.168 19.692 ;
  LAYER M2 ;
        RECT 3.116 19.64 3.188 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 3.152 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 22.8 ;
  LAYER M2 ;
        RECT 3.116 22.748 3.188 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 3.152 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 22.764 ;
  LAYER M1 ;
        RECT 9.728 0.972 9.76 1.044 ;
  LAYER M2 ;
        RECT 9.708 0.992 9.78 1.024 ;
  LAYER M1 ;
        RECT 9.728 0.84 9.76 1.008 ;
  LAYER M1 ;
        RECT 9.728 0.804 9.76 0.876 ;
  LAYER M2 ;
        RECT 9.708 0.824 9.78 0.856 ;
  LAYER M2 ;
        RECT 9.744 0.824 9.968 0.856 ;
  LAYER M1 ;
        RECT 9.952 0.804 9.984 0.876 ;
  LAYER M2 ;
        RECT 9.932 0.824 10.004 0.856 ;
  LAYER M1 ;
        RECT 9.728 4.08 9.76 4.152 ;
  LAYER M2 ;
        RECT 9.708 4.1 9.78 4.132 ;
  LAYER M1 ;
        RECT 9.728 3.948 9.76 4.116 ;
  LAYER M1 ;
        RECT 9.728 3.912 9.76 3.984 ;
  LAYER M2 ;
        RECT 9.708 3.932 9.78 3.964 ;
  LAYER M2 ;
        RECT 9.744 3.932 9.968 3.964 ;
  LAYER M1 ;
        RECT 9.952 3.912 9.984 3.984 ;
  LAYER M2 ;
        RECT 9.932 3.932 10.004 3.964 ;
  LAYER M1 ;
        RECT 9.728 7.188 9.76 7.26 ;
  LAYER M2 ;
        RECT 9.708 7.208 9.78 7.24 ;
  LAYER M1 ;
        RECT 9.728 7.056 9.76 7.224 ;
  LAYER M1 ;
        RECT 9.728 7.02 9.76 7.092 ;
  LAYER M2 ;
        RECT 9.708 7.04 9.78 7.072 ;
  LAYER M2 ;
        RECT 9.744 7.04 9.968 7.072 ;
  LAYER M1 ;
        RECT 9.952 7.02 9.984 7.092 ;
  LAYER M2 ;
        RECT 9.932 7.04 10.004 7.072 ;
  LAYER M1 ;
        RECT 9.728 10.296 9.76 10.368 ;
  LAYER M2 ;
        RECT 9.708 10.316 9.78 10.348 ;
  LAYER M1 ;
        RECT 9.728 10.164 9.76 10.332 ;
  LAYER M1 ;
        RECT 9.728 10.128 9.76 10.2 ;
  LAYER M2 ;
        RECT 9.708 10.148 9.78 10.18 ;
  LAYER M2 ;
        RECT 9.744 10.148 9.968 10.18 ;
  LAYER M1 ;
        RECT 9.952 10.128 9.984 10.2 ;
  LAYER M2 ;
        RECT 9.932 10.148 10.004 10.18 ;
  LAYER M1 ;
        RECT 9.728 13.404 9.76 13.476 ;
  LAYER M2 ;
        RECT 9.708 13.424 9.78 13.456 ;
  LAYER M1 ;
        RECT 9.728 13.272 9.76 13.44 ;
  LAYER M1 ;
        RECT 9.728 13.236 9.76 13.308 ;
  LAYER M2 ;
        RECT 9.708 13.256 9.78 13.288 ;
  LAYER M2 ;
        RECT 9.744 13.256 9.968 13.288 ;
  LAYER M1 ;
        RECT 9.952 13.236 9.984 13.308 ;
  LAYER M2 ;
        RECT 9.932 13.256 10.004 13.288 ;
  LAYER M1 ;
        RECT 9.728 16.512 9.76 16.584 ;
  LAYER M2 ;
        RECT 9.708 16.532 9.78 16.564 ;
  LAYER M1 ;
        RECT 9.728 16.38 9.76 16.548 ;
  LAYER M1 ;
        RECT 9.728 16.344 9.76 16.416 ;
  LAYER M2 ;
        RECT 9.708 16.364 9.78 16.396 ;
  LAYER M2 ;
        RECT 9.744 16.364 9.968 16.396 ;
  LAYER M1 ;
        RECT 9.952 16.344 9.984 16.416 ;
  LAYER M2 ;
        RECT 9.932 16.364 10.004 16.396 ;
  LAYER M1 ;
        RECT 9.728 19.62 9.76 19.692 ;
  LAYER M2 ;
        RECT 9.708 19.64 9.78 19.672 ;
  LAYER M1 ;
        RECT 9.728 19.488 9.76 19.656 ;
  LAYER M1 ;
        RECT 9.728 19.452 9.76 19.524 ;
  LAYER M2 ;
        RECT 9.708 19.472 9.78 19.504 ;
  LAYER M2 ;
        RECT 9.744 19.472 9.968 19.504 ;
  LAYER M1 ;
        RECT 9.952 19.452 9.984 19.524 ;
  LAYER M2 ;
        RECT 9.932 19.472 10.004 19.504 ;
  LAYER M1 ;
        RECT 9.728 22.728 9.76 22.8 ;
  LAYER M2 ;
        RECT 9.708 22.748 9.78 22.78 ;
  LAYER M1 ;
        RECT 9.728 22.596 9.76 22.764 ;
  LAYER M1 ;
        RECT 9.728 22.56 9.76 22.632 ;
  LAYER M2 ;
        RECT 9.708 22.58 9.78 22.612 ;
  LAYER M2 ;
        RECT 9.744 22.58 9.968 22.612 ;
  LAYER M1 ;
        RECT 9.952 22.56 9.984 22.632 ;
  LAYER M2 ;
        RECT 9.932 22.58 10.004 22.612 ;
  LAYER M1 ;
        RECT 9.952 0.048 9.984 0.12 ;
  LAYER M2 ;
        RECT 9.932 0.068 10.004 0.1 ;
  LAYER M1 ;
        RECT 9.952 0.084 9.984 0.672 ;
  LAYER M1 ;
        RECT 9.952 0.672 9.984 22.596 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.968 0.1 ;
  LAYER M1 ;
        RECT 6.432 0.972 6.464 1.044 ;
  LAYER M2 ;
        RECT 6.412 0.992 6.484 1.024 ;
  LAYER M2 ;
        RECT 3.152 0.992 6.448 1.024 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M1 ;
        RECT 6.432 22.728 6.464 22.8 ;
  LAYER M2 ;
        RECT 6.412 22.748 6.484 22.78 ;
  LAYER M2 ;
        RECT 3.152 22.748 6.448 22.78 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 22.8 ;
  LAYER M2 ;
        RECT 3.116 22.748 3.188 22.78 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M2 ;
        RECT 3.696 15.86 4.08 15.892 ;
  LAYER M1 ;
        RECT 3.68 15.84 3.712 15.912 ;
  LAYER M2 ;
        RECT 3.66 15.86 3.732 15.892 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M2 ;
        RECT 3.696 9.644 4.08 9.676 ;
  LAYER M1 ;
        RECT 3.68 9.624 3.712 9.696 ;
  LAYER M2 ;
        RECT 3.66 9.644 3.732 9.676 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M2 ;
        RECT 3.696 18.968 4.08 19 ;
  LAYER M1 ;
        RECT 3.68 18.948 3.712 19.02 ;
  LAYER M2 ;
        RECT 3.66 18.968 3.732 19 ;
  LAYER M1 ;
        RECT 3.68 25.752 3.712 25.824 ;
  LAYER M2 ;
        RECT 3.66 25.772 3.732 25.804 ;
  LAYER M1 ;
        RECT 3.68 25.536 3.712 25.788 ;
  LAYER M1 ;
        RECT 3.68 9.66 3.712 25.536 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M1 ;
        RECT 4.064 15.876 4.096 16.044 ;
  LAYER M1 ;
        RECT 4.064 16.008 4.096 16.08 ;
  LAYER M2 ;
        RECT 4.044 16.028 4.116 16.06 ;
  LAYER M2 ;
        RECT 4.08 16.028 6.992 16.06 ;
  LAYER M1 ;
        RECT 6.976 16.008 7.008 16.08 ;
  LAYER M2 ;
        RECT 6.956 16.028 7.028 16.06 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M1 ;
        RECT 4.064 9.66 4.096 9.828 ;
  LAYER M1 ;
        RECT 4.064 9.792 4.096 9.864 ;
  LAYER M2 ;
        RECT 4.044 9.812 4.116 9.844 ;
  LAYER M2 ;
        RECT 4.08 9.812 6.992 9.844 ;
  LAYER M1 ;
        RECT 6.976 9.792 7.008 9.864 ;
  LAYER M2 ;
        RECT 6.956 9.812 7.028 9.844 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M1 ;
        RECT 4.064 18.984 4.096 19.152 ;
  LAYER M1 ;
        RECT 4.064 19.116 4.096 19.188 ;
  LAYER M2 ;
        RECT 4.044 19.136 4.116 19.168 ;
  LAYER M2 ;
        RECT 4.08 19.136 6.992 19.168 ;
  LAYER M1 ;
        RECT 6.976 19.116 7.008 19.188 ;
  LAYER M2 ;
        RECT 6.956 19.136 7.028 19.168 ;
  LAYER M1 ;
        RECT 6.976 25.752 7.008 25.824 ;
  LAYER M2 ;
        RECT 6.956 25.772 7.028 25.804 ;
  LAYER M1 ;
        RECT 6.976 25.536 7.008 25.788 ;
  LAYER M1 ;
        RECT 6.976 9.828 7.008 25.536 ;
  LAYER M2 ;
        RECT 3.696 25.772 6.992 25.804 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M2 ;
        RECT 3.856 12.752 4.08 12.784 ;
  LAYER M1 ;
        RECT 3.84 12.732 3.872 12.804 ;
  LAYER M2 ;
        RECT 3.82 12.752 3.892 12.784 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M2 ;
        RECT 3.856 6.536 4.08 6.568 ;
  LAYER M1 ;
        RECT 3.84 6.516 3.872 6.588 ;
  LAYER M2 ;
        RECT 3.82 6.536 3.892 6.568 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M2 ;
        RECT 3.856 22.076 4.08 22.108 ;
  LAYER M1 ;
        RECT 3.84 22.056 3.872 22.128 ;
  LAYER M2 ;
        RECT 3.82 22.076 3.892 22.108 ;
  LAYER M1 ;
        RECT 3.84 25.92 3.872 25.992 ;
  LAYER M2 ;
        RECT 3.82 25.94 3.892 25.972 ;
  LAYER M1 ;
        RECT 3.84 25.536 3.872 25.956 ;
  LAYER M1 ;
        RECT 3.84 6.552 3.872 25.536 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M1 ;
        RECT 4.064 12.768 4.096 12.936 ;
  LAYER M1 ;
        RECT 4.064 12.9 4.096 12.972 ;
  LAYER M2 ;
        RECT 4.044 12.92 4.116 12.952 ;
  LAYER M2 ;
        RECT 4.08 12.92 7.152 12.952 ;
  LAYER M1 ;
        RECT 7.136 12.9 7.168 12.972 ;
  LAYER M2 ;
        RECT 7.116 12.92 7.188 12.952 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M1 ;
        RECT 4.064 6.552 4.096 6.72 ;
  LAYER M1 ;
        RECT 4.064 6.684 4.096 6.756 ;
  LAYER M2 ;
        RECT 4.044 6.704 4.116 6.736 ;
  LAYER M2 ;
        RECT 4.08 6.704 7.152 6.736 ;
  LAYER M1 ;
        RECT 7.136 6.684 7.168 6.756 ;
  LAYER M2 ;
        RECT 7.116 6.704 7.188 6.736 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M1 ;
        RECT 4.064 22.092 4.096 22.26 ;
  LAYER M1 ;
        RECT 4.064 22.224 4.096 22.296 ;
  LAYER M2 ;
        RECT 4.044 22.244 4.116 22.276 ;
  LAYER M2 ;
        RECT 4.08 22.244 7.152 22.276 ;
  LAYER M1 ;
        RECT 7.136 22.224 7.168 22.296 ;
  LAYER M2 ;
        RECT 7.116 22.244 7.188 22.276 ;
  LAYER M1 ;
        RECT 7.136 25.92 7.168 25.992 ;
  LAYER M2 ;
        RECT 7.116 25.94 7.188 25.972 ;
  LAYER M1 ;
        RECT 7.136 25.536 7.168 25.956 ;
  LAYER M1 ;
        RECT 7.136 6.72 7.168 25.536 ;
  LAYER M2 ;
        RECT 3.856 25.94 7.152 25.972 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.784 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.768 6.516 0.8 6.588 ;
  LAYER M2 ;
        RECT 0.748 6.536 0.82 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.784 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.768 9.624 0.8 9.696 ;
  LAYER M2 ;
        RECT 0.748 9.644 0.82 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.784 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.768 12.732 0.8 12.804 ;
  LAYER M2 ;
        RECT 0.748 12.752 0.82 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.784 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.768 15.84 0.8 15.912 ;
  LAYER M2 ;
        RECT 0.748 15.86 0.82 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.784 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.768 18.948 0.8 19.02 ;
  LAYER M2 ;
        RECT 0.748 18.968 0.82 19 ;
  LAYER M2 ;
        RECT 0.24 18.968 0.784 19 ;
  LAYER M1 ;
        RECT 0.224 18.948 0.256 19.02 ;
  LAYER M2 ;
        RECT 0.204 18.968 0.276 19 ;
  LAYER M1 ;
        RECT 0.768 22.056 0.8 22.128 ;
  LAYER M2 ;
        RECT 0.748 22.076 0.82 22.108 ;
  LAYER M2 ;
        RECT 0.24 22.076 0.784 22.108 ;
  LAYER M1 ;
        RECT 0.224 22.056 0.256 22.128 ;
  LAYER M2 ;
        RECT 0.204 22.076 0.276 22.108 ;
  LAYER M1 ;
        RECT 0.768 25.164 0.8 25.236 ;
  LAYER M2 ;
        RECT 0.748 25.184 0.82 25.216 ;
  LAYER M2 ;
        RECT 0.24 25.184 0.784 25.216 ;
  LAYER M1 ;
        RECT 0.224 25.164 0.256 25.236 ;
  LAYER M2 ;
        RECT 0.204 25.184 0.276 25.216 ;
  LAYER M1 ;
        RECT 0.224 26.088 0.256 26.16 ;
  LAYER M2 ;
        RECT 0.204 26.108 0.276 26.14 ;
  LAYER M1 ;
        RECT 0.224 25.536 0.256 26.124 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 25.536 ;
  LAYER M1 ;
        RECT 7.36 3.408 7.392 3.48 ;
  LAYER M2 ;
        RECT 7.34 3.428 7.412 3.46 ;
  LAYER M1 ;
        RECT 7.36 3.444 7.392 3.612 ;
  LAYER M1 ;
        RECT 7.36 3.576 7.392 3.648 ;
  LAYER M2 ;
        RECT 7.34 3.596 7.412 3.628 ;
  LAYER M2 ;
        RECT 7.376 3.596 10.128 3.628 ;
  LAYER M1 ;
        RECT 10.112 3.576 10.144 3.648 ;
  LAYER M2 ;
        RECT 10.092 3.596 10.164 3.628 ;
  LAYER M1 ;
        RECT 7.36 6.516 7.392 6.588 ;
  LAYER M2 ;
        RECT 7.34 6.536 7.412 6.568 ;
  LAYER M1 ;
        RECT 7.36 6.552 7.392 6.72 ;
  LAYER M1 ;
        RECT 7.36 6.684 7.392 6.756 ;
  LAYER M2 ;
        RECT 7.34 6.704 7.412 6.736 ;
  LAYER M2 ;
        RECT 7.376 6.704 10.128 6.736 ;
  LAYER M1 ;
        RECT 10.112 6.684 10.144 6.756 ;
  LAYER M2 ;
        RECT 10.092 6.704 10.164 6.736 ;
  LAYER M1 ;
        RECT 7.36 9.624 7.392 9.696 ;
  LAYER M2 ;
        RECT 7.34 9.644 7.412 9.676 ;
  LAYER M1 ;
        RECT 7.36 9.66 7.392 9.828 ;
  LAYER M1 ;
        RECT 7.36 9.792 7.392 9.864 ;
  LAYER M2 ;
        RECT 7.34 9.812 7.412 9.844 ;
  LAYER M2 ;
        RECT 7.376 9.812 10.128 9.844 ;
  LAYER M1 ;
        RECT 10.112 9.792 10.144 9.864 ;
  LAYER M2 ;
        RECT 10.092 9.812 10.164 9.844 ;
  LAYER M1 ;
        RECT 7.36 12.732 7.392 12.804 ;
  LAYER M2 ;
        RECT 7.34 12.752 7.412 12.784 ;
  LAYER M1 ;
        RECT 7.36 12.768 7.392 12.936 ;
  LAYER M1 ;
        RECT 7.36 12.9 7.392 12.972 ;
  LAYER M2 ;
        RECT 7.34 12.92 7.412 12.952 ;
  LAYER M2 ;
        RECT 7.376 12.92 10.128 12.952 ;
  LAYER M1 ;
        RECT 10.112 12.9 10.144 12.972 ;
  LAYER M2 ;
        RECT 10.092 12.92 10.164 12.952 ;
  LAYER M1 ;
        RECT 7.36 15.84 7.392 15.912 ;
  LAYER M2 ;
        RECT 7.34 15.86 7.412 15.892 ;
  LAYER M1 ;
        RECT 7.36 15.876 7.392 16.044 ;
  LAYER M1 ;
        RECT 7.36 16.008 7.392 16.08 ;
  LAYER M2 ;
        RECT 7.34 16.028 7.412 16.06 ;
  LAYER M2 ;
        RECT 7.376 16.028 10.128 16.06 ;
  LAYER M1 ;
        RECT 10.112 16.008 10.144 16.08 ;
  LAYER M2 ;
        RECT 10.092 16.028 10.164 16.06 ;
  LAYER M1 ;
        RECT 7.36 18.948 7.392 19.02 ;
  LAYER M2 ;
        RECT 7.34 18.968 7.412 19 ;
  LAYER M1 ;
        RECT 7.36 18.984 7.392 19.152 ;
  LAYER M1 ;
        RECT 7.36 19.116 7.392 19.188 ;
  LAYER M2 ;
        RECT 7.34 19.136 7.412 19.168 ;
  LAYER M2 ;
        RECT 7.376 19.136 10.128 19.168 ;
  LAYER M1 ;
        RECT 10.112 19.116 10.144 19.188 ;
  LAYER M2 ;
        RECT 10.092 19.136 10.164 19.168 ;
  LAYER M1 ;
        RECT 7.36 22.056 7.392 22.128 ;
  LAYER M2 ;
        RECT 7.34 22.076 7.412 22.108 ;
  LAYER M1 ;
        RECT 7.36 22.092 7.392 22.26 ;
  LAYER M1 ;
        RECT 7.36 22.224 7.392 22.296 ;
  LAYER M2 ;
        RECT 7.34 22.244 7.412 22.276 ;
  LAYER M2 ;
        RECT 7.376 22.244 10.128 22.276 ;
  LAYER M1 ;
        RECT 10.112 22.224 10.144 22.296 ;
  LAYER M2 ;
        RECT 10.092 22.244 10.164 22.276 ;
  LAYER M1 ;
        RECT 7.36 25.164 7.392 25.236 ;
  LAYER M2 ;
        RECT 7.34 25.184 7.412 25.216 ;
  LAYER M1 ;
        RECT 7.36 25.2 7.392 25.368 ;
  LAYER M1 ;
        RECT 7.36 25.332 7.392 25.404 ;
  LAYER M2 ;
        RECT 7.34 25.352 7.412 25.384 ;
  LAYER M2 ;
        RECT 7.376 25.352 10.128 25.384 ;
  LAYER M1 ;
        RECT 10.112 25.332 10.144 25.404 ;
  LAYER M2 ;
        RECT 10.092 25.352 10.164 25.384 ;
  LAYER M1 ;
        RECT 10.112 26.088 10.144 26.16 ;
  LAYER M2 ;
        RECT 10.092 26.108 10.164 26.14 ;
  LAYER M1 ;
        RECT 10.112 25.536 10.144 26.124 ;
  LAYER M1 ;
        RECT 10.112 3.612 10.144 25.536 ;
  LAYER M2 ;
        RECT 0.24 26.108 10.128 26.14 ;
  LAYER M1 ;
        RECT 4.064 3.408 4.096 3.48 ;
  LAYER M2 ;
        RECT 4.044 3.428 4.116 3.46 ;
  LAYER M2 ;
        RECT 0.784 3.428 4.08 3.46 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M1 ;
        RECT 4.064 25.164 4.096 25.236 ;
  LAYER M2 ;
        RECT 4.044 25.184 4.116 25.216 ;
  LAYER M2 ;
        RECT 0.784 25.184 4.08 25.216 ;
  LAYER M1 ;
        RECT 0.768 25.164 0.8 25.236 ;
  LAYER M2 ;
        RECT 0.748 25.184 0.82 25.216 ;
  LAYER M1 ;
        RECT 0.768 0.972 0.8 3.48 ;
  LAYER M3 ;
        RECT 0.768 3.428 0.8 3.46 ;
  LAYER M1 ;
        RECT 0.832 0.972 0.864 3.48 ;
  LAYER M3 ;
        RECT 0.832 0.992 0.864 1.024 ;
  LAYER M1 ;
        RECT 0.896 0.972 0.928 3.48 ;
  LAYER M3 ;
        RECT 0.896 3.428 0.928 3.46 ;
  LAYER M1 ;
        RECT 0.96 0.972 0.992 3.48 ;
  LAYER M3 ;
        RECT 0.96 0.992 0.992 1.024 ;
  LAYER M1 ;
        RECT 1.024 0.972 1.056 3.48 ;
  LAYER M3 ;
        RECT 1.024 3.428 1.056 3.46 ;
  LAYER M1 ;
        RECT 1.088 0.972 1.12 3.48 ;
  LAYER M3 ;
        RECT 1.088 0.992 1.12 1.024 ;
  LAYER M1 ;
        RECT 1.152 0.972 1.184 3.48 ;
  LAYER M3 ;
        RECT 1.152 3.428 1.184 3.46 ;
  LAYER M1 ;
        RECT 1.216 0.972 1.248 3.48 ;
  LAYER M3 ;
        RECT 1.216 0.992 1.248 1.024 ;
  LAYER M1 ;
        RECT 1.28 0.972 1.312 3.48 ;
  LAYER M3 ;
        RECT 1.28 3.428 1.312 3.46 ;
  LAYER M1 ;
        RECT 1.344 0.972 1.376 3.48 ;
  LAYER M3 ;
        RECT 1.344 0.992 1.376 1.024 ;
  LAYER M1 ;
        RECT 1.408 0.972 1.44 3.48 ;
  LAYER M3 ;
        RECT 1.408 3.428 1.44 3.46 ;
  LAYER M1 ;
        RECT 1.472 0.972 1.504 3.48 ;
  LAYER M3 ;
        RECT 1.472 0.992 1.504 1.024 ;
  LAYER M1 ;
        RECT 1.536 0.972 1.568 3.48 ;
  LAYER M3 ;
        RECT 1.536 3.428 1.568 3.46 ;
  LAYER M1 ;
        RECT 1.6 0.972 1.632 3.48 ;
  LAYER M3 ;
        RECT 1.6 0.992 1.632 1.024 ;
  LAYER M1 ;
        RECT 1.664 0.972 1.696 3.48 ;
  LAYER M3 ;
        RECT 1.664 3.428 1.696 3.46 ;
  LAYER M1 ;
        RECT 1.728 0.972 1.76 3.48 ;
  LAYER M3 ;
        RECT 1.728 0.992 1.76 1.024 ;
  LAYER M1 ;
        RECT 1.792 0.972 1.824 3.48 ;
  LAYER M3 ;
        RECT 1.792 3.428 1.824 3.46 ;
  LAYER M1 ;
        RECT 1.856 0.972 1.888 3.48 ;
  LAYER M3 ;
        RECT 1.856 0.992 1.888 1.024 ;
  LAYER M1 ;
        RECT 1.92 0.972 1.952 3.48 ;
  LAYER M3 ;
        RECT 1.92 3.428 1.952 3.46 ;
  LAYER M1 ;
        RECT 1.984 0.972 2.016 3.48 ;
  LAYER M3 ;
        RECT 1.984 0.992 2.016 1.024 ;
  LAYER M1 ;
        RECT 2.048 0.972 2.08 3.48 ;
  LAYER M3 ;
        RECT 2.048 3.428 2.08 3.46 ;
  LAYER M1 ;
        RECT 2.112 0.972 2.144 3.48 ;
  LAYER M3 ;
        RECT 2.112 0.992 2.144 1.024 ;
  LAYER M1 ;
        RECT 2.176 0.972 2.208 3.48 ;
  LAYER M3 ;
        RECT 2.176 3.428 2.208 3.46 ;
  LAYER M1 ;
        RECT 2.24 0.972 2.272 3.48 ;
  LAYER M3 ;
        RECT 2.24 0.992 2.272 1.024 ;
  LAYER M1 ;
        RECT 2.304 0.972 2.336 3.48 ;
  LAYER M3 ;
        RECT 2.304 3.428 2.336 3.46 ;
  LAYER M1 ;
        RECT 2.368 0.972 2.4 3.48 ;
  LAYER M3 ;
        RECT 2.368 0.992 2.4 1.024 ;
  LAYER M1 ;
        RECT 2.432 0.972 2.464 3.48 ;
  LAYER M3 ;
        RECT 2.432 3.428 2.464 3.46 ;
  LAYER M1 ;
        RECT 2.496 0.972 2.528 3.48 ;
  LAYER M3 ;
        RECT 2.496 0.992 2.528 1.024 ;
  LAYER M1 ;
        RECT 2.56 0.972 2.592 3.48 ;
  LAYER M3 ;
        RECT 2.56 3.428 2.592 3.46 ;
  LAYER M1 ;
        RECT 2.624 0.972 2.656 3.48 ;
  LAYER M3 ;
        RECT 2.624 0.992 2.656 1.024 ;
  LAYER M1 ;
        RECT 2.688 0.972 2.72 3.48 ;
  LAYER M3 ;
        RECT 2.688 3.428 2.72 3.46 ;
  LAYER M1 ;
        RECT 2.752 0.972 2.784 3.48 ;
  LAYER M3 ;
        RECT 2.752 0.992 2.784 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 3.48 ;
  LAYER M3 ;
        RECT 2.816 3.428 2.848 3.46 ;
  LAYER M1 ;
        RECT 2.88 0.972 2.912 3.48 ;
  LAYER M3 ;
        RECT 2.88 0.992 2.912 1.024 ;
  LAYER M1 ;
        RECT 2.944 0.972 2.976 3.48 ;
  LAYER M3 ;
        RECT 2.944 3.428 2.976 3.46 ;
  LAYER M1 ;
        RECT 3.008 0.972 3.04 3.48 ;
  LAYER M3 ;
        RECT 3.008 0.992 3.04 1.024 ;
  LAYER M1 ;
        RECT 3.072 0.972 3.104 3.48 ;
  LAYER M3 ;
        RECT 3.072 3.428 3.104 3.46 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 3.48 ;
  LAYER M3 ;
        RECT 0.768 1.056 0.8 1.088 ;
  LAYER M2 ;
        RECT 3.136 1.12 3.168 1.152 ;
  LAYER M2 ;
        RECT 0.768 1.184 0.8 1.216 ;
  LAYER M2 ;
        RECT 3.136 1.248 3.168 1.28 ;
  LAYER M2 ;
        RECT 0.768 1.312 0.8 1.344 ;
  LAYER M2 ;
        RECT 3.136 1.376 3.168 1.408 ;
  LAYER M2 ;
        RECT 0.768 1.44 0.8 1.472 ;
  LAYER M2 ;
        RECT 3.136 1.504 3.168 1.536 ;
  LAYER M2 ;
        RECT 0.768 1.568 0.8 1.6 ;
  LAYER M2 ;
        RECT 3.136 1.632 3.168 1.664 ;
  LAYER M2 ;
        RECT 0.768 1.696 0.8 1.728 ;
  LAYER M2 ;
        RECT 3.136 1.76 3.168 1.792 ;
  LAYER M2 ;
        RECT 0.768 1.824 0.8 1.856 ;
  LAYER M2 ;
        RECT 3.136 1.888 3.168 1.92 ;
  LAYER M2 ;
        RECT 0.768 1.952 0.8 1.984 ;
  LAYER M2 ;
        RECT 3.136 2.016 3.168 2.048 ;
  LAYER M2 ;
        RECT 0.768 2.08 0.8 2.112 ;
  LAYER M2 ;
        RECT 3.136 2.144 3.168 2.176 ;
  LAYER M2 ;
        RECT 0.768 2.208 0.8 2.24 ;
  LAYER M2 ;
        RECT 3.136 2.272 3.168 2.304 ;
  LAYER M2 ;
        RECT 0.768 2.336 0.8 2.368 ;
  LAYER M2 ;
        RECT 3.136 2.4 3.168 2.432 ;
  LAYER M2 ;
        RECT 0.768 2.464 0.8 2.496 ;
  LAYER M2 ;
        RECT 3.136 2.528 3.168 2.56 ;
  LAYER M2 ;
        RECT 0.768 2.592 0.8 2.624 ;
  LAYER M2 ;
        RECT 3.136 2.656 3.168 2.688 ;
  LAYER M2 ;
        RECT 0.768 2.72 0.8 2.752 ;
  LAYER M2 ;
        RECT 3.136 2.784 3.168 2.816 ;
  LAYER M2 ;
        RECT 0.768 2.848 0.8 2.88 ;
  LAYER M2 ;
        RECT 3.136 2.912 3.168 2.944 ;
  LAYER M2 ;
        RECT 0.768 2.976 0.8 3.008 ;
  LAYER M2 ;
        RECT 3.136 3.04 3.168 3.072 ;
  LAYER M2 ;
        RECT 0.768 3.104 0.8 3.136 ;
  LAYER M2 ;
        RECT 3.136 3.168 3.168 3.2 ;
  LAYER M2 ;
        RECT 0.768 3.232 0.8 3.264 ;
  LAYER M2 ;
        RECT 3.136 3.296 3.168 3.328 ;
  LAYER M2 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M1 ;
        RECT 0.768 4.08 0.8 6.588 ;
  LAYER M3 ;
        RECT 0.768 6.536 0.8 6.568 ;
  LAYER M1 ;
        RECT 0.832 4.08 0.864 6.588 ;
  LAYER M3 ;
        RECT 0.832 4.1 0.864 4.132 ;
  LAYER M1 ;
        RECT 0.896 4.08 0.928 6.588 ;
  LAYER M3 ;
        RECT 0.896 6.536 0.928 6.568 ;
  LAYER M1 ;
        RECT 0.96 4.08 0.992 6.588 ;
  LAYER M3 ;
        RECT 0.96 4.1 0.992 4.132 ;
  LAYER M1 ;
        RECT 1.024 4.08 1.056 6.588 ;
  LAYER M3 ;
        RECT 1.024 6.536 1.056 6.568 ;
  LAYER M1 ;
        RECT 1.088 4.08 1.12 6.588 ;
  LAYER M3 ;
        RECT 1.088 4.1 1.12 4.132 ;
  LAYER M1 ;
        RECT 1.152 4.08 1.184 6.588 ;
  LAYER M3 ;
        RECT 1.152 6.536 1.184 6.568 ;
  LAYER M1 ;
        RECT 1.216 4.08 1.248 6.588 ;
  LAYER M3 ;
        RECT 1.216 4.1 1.248 4.132 ;
  LAYER M1 ;
        RECT 1.28 4.08 1.312 6.588 ;
  LAYER M3 ;
        RECT 1.28 6.536 1.312 6.568 ;
  LAYER M1 ;
        RECT 1.344 4.08 1.376 6.588 ;
  LAYER M3 ;
        RECT 1.344 4.1 1.376 4.132 ;
  LAYER M1 ;
        RECT 1.408 4.08 1.44 6.588 ;
  LAYER M3 ;
        RECT 1.408 6.536 1.44 6.568 ;
  LAYER M1 ;
        RECT 1.472 4.08 1.504 6.588 ;
  LAYER M3 ;
        RECT 1.472 4.1 1.504 4.132 ;
  LAYER M1 ;
        RECT 1.536 4.08 1.568 6.588 ;
  LAYER M3 ;
        RECT 1.536 6.536 1.568 6.568 ;
  LAYER M1 ;
        RECT 1.6 4.08 1.632 6.588 ;
  LAYER M3 ;
        RECT 1.6 4.1 1.632 4.132 ;
  LAYER M1 ;
        RECT 1.664 4.08 1.696 6.588 ;
  LAYER M3 ;
        RECT 1.664 6.536 1.696 6.568 ;
  LAYER M1 ;
        RECT 1.728 4.08 1.76 6.588 ;
  LAYER M3 ;
        RECT 1.728 4.1 1.76 4.132 ;
  LAYER M1 ;
        RECT 1.792 4.08 1.824 6.588 ;
  LAYER M3 ;
        RECT 1.792 6.536 1.824 6.568 ;
  LAYER M1 ;
        RECT 1.856 4.08 1.888 6.588 ;
  LAYER M3 ;
        RECT 1.856 4.1 1.888 4.132 ;
  LAYER M1 ;
        RECT 1.92 4.08 1.952 6.588 ;
  LAYER M3 ;
        RECT 1.92 6.536 1.952 6.568 ;
  LAYER M1 ;
        RECT 1.984 4.08 2.016 6.588 ;
  LAYER M3 ;
        RECT 1.984 4.1 2.016 4.132 ;
  LAYER M1 ;
        RECT 2.048 4.08 2.08 6.588 ;
  LAYER M3 ;
        RECT 2.048 6.536 2.08 6.568 ;
  LAYER M1 ;
        RECT 2.112 4.08 2.144 6.588 ;
  LAYER M3 ;
        RECT 2.112 4.1 2.144 4.132 ;
  LAYER M1 ;
        RECT 2.176 4.08 2.208 6.588 ;
  LAYER M3 ;
        RECT 2.176 6.536 2.208 6.568 ;
  LAYER M1 ;
        RECT 2.24 4.08 2.272 6.588 ;
  LAYER M3 ;
        RECT 2.24 4.1 2.272 4.132 ;
  LAYER M1 ;
        RECT 2.304 4.08 2.336 6.588 ;
  LAYER M3 ;
        RECT 2.304 6.536 2.336 6.568 ;
  LAYER M1 ;
        RECT 2.368 4.08 2.4 6.588 ;
  LAYER M3 ;
        RECT 2.368 4.1 2.4 4.132 ;
  LAYER M1 ;
        RECT 2.432 4.08 2.464 6.588 ;
  LAYER M3 ;
        RECT 2.432 6.536 2.464 6.568 ;
  LAYER M1 ;
        RECT 2.496 4.08 2.528 6.588 ;
  LAYER M3 ;
        RECT 2.496 4.1 2.528 4.132 ;
  LAYER M1 ;
        RECT 2.56 4.08 2.592 6.588 ;
  LAYER M3 ;
        RECT 2.56 6.536 2.592 6.568 ;
  LAYER M1 ;
        RECT 2.624 4.08 2.656 6.588 ;
  LAYER M3 ;
        RECT 2.624 4.1 2.656 4.132 ;
  LAYER M1 ;
        RECT 2.688 4.08 2.72 6.588 ;
  LAYER M3 ;
        RECT 2.688 6.536 2.72 6.568 ;
  LAYER M1 ;
        RECT 2.752 4.08 2.784 6.588 ;
  LAYER M3 ;
        RECT 2.752 4.1 2.784 4.132 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 6.588 ;
  LAYER M3 ;
        RECT 2.816 6.536 2.848 6.568 ;
  LAYER M1 ;
        RECT 2.88 4.08 2.912 6.588 ;
  LAYER M3 ;
        RECT 2.88 4.1 2.912 4.132 ;
  LAYER M1 ;
        RECT 2.944 4.08 2.976 6.588 ;
  LAYER M3 ;
        RECT 2.944 6.536 2.976 6.568 ;
  LAYER M1 ;
        RECT 3.008 4.08 3.04 6.588 ;
  LAYER M3 ;
        RECT 3.008 4.1 3.04 4.132 ;
  LAYER M1 ;
        RECT 3.072 4.08 3.104 6.588 ;
  LAYER M3 ;
        RECT 3.072 6.536 3.104 6.568 ;
  LAYER M1 ;
        RECT 3.136 4.08 3.168 6.588 ;
  LAYER M3 ;
        RECT 0.768 4.164 0.8 4.196 ;
  LAYER M2 ;
        RECT 3.136 4.228 3.168 4.26 ;
  LAYER M2 ;
        RECT 0.768 4.292 0.8 4.324 ;
  LAYER M2 ;
        RECT 3.136 4.356 3.168 4.388 ;
  LAYER M2 ;
        RECT 0.768 4.42 0.8 4.452 ;
  LAYER M2 ;
        RECT 3.136 4.484 3.168 4.516 ;
  LAYER M2 ;
        RECT 0.768 4.548 0.8 4.58 ;
  LAYER M2 ;
        RECT 3.136 4.612 3.168 4.644 ;
  LAYER M2 ;
        RECT 0.768 4.676 0.8 4.708 ;
  LAYER M2 ;
        RECT 3.136 4.74 3.168 4.772 ;
  LAYER M2 ;
        RECT 0.768 4.804 0.8 4.836 ;
  LAYER M2 ;
        RECT 3.136 4.868 3.168 4.9 ;
  LAYER M2 ;
        RECT 0.768 4.932 0.8 4.964 ;
  LAYER M2 ;
        RECT 3.136 4.996 3.168 5.028 ;
  LAYER M2 ;
        RECT 0.768 5.06 0.8 5.092 ;
  LAYER M2 ;
        RECT 3.136 5.124 3.168 5.156 ;
  LAYER M2 ;
        RECT 0.768 5.188 0.8 5.22 ;
  LAYER M2 ;
        RECT 3.136 5.252 3.168 5.284 ;
  LAYER M2 ;
        RECT 0.768 5.316 0.8 5.348 ;
  LAYER M2 ;
        RECT 3.136 5.38 3.168 5.412 ;
  LAYER M2 ;
        RECT 0.768 5.444 0.8 5.476 ;
  LAYER M2 ;
        RECT 3.136 5.508 3.168 5.54 ;
  LAYER M2 ;
        RECT 0.768 5.572 0.8 5.604 ;
  LAYER M2 ;
        RECT 3.136 5.636 3.168 5.668 ;
  LAYER M2 ;
        RECT 0.768 5.7 0.8 5.732 ;
  LAYER M2 ;
        RECT 3.136 5.764 3.168 5.796 ;
  LAYER M2 ;
        RECT 0.768 5.828 0.8 5.86 ;
  LAYER M2 ;
        RECT 3.136 5.892 3.168 5.924 ;
  LAYER M2 ;
        RECT 0.768 5.956 0.8 5.988 ;
  LAYER M2 ;
        RECT 3.136 6.02 3.168 6.052 ;
  LAYER M2 ;
        RECT 0.768 6.084 0.8 6.116 ;
  LAYER M2 ;
        RECT 3.136 6.148 3.168 6.18 ;
  LAYER M2 ;
        RECT 0.768 6.212 0.8 6.244 ;
  LAYER M2 ;
        RECT 3.136 6.276 3.168 6.308 ;
  LAYER M2 ;
        RECT 0.768 6.34 0.8 6.372 ;
  LAYER M2 ;
        RECT 3.136 6.404 3.168 6.436 ;
  LAYER M2 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M1 ;
        RECT 0.768 7.188 0.8 9.696 ;
  LAYER M3 ;
        RECT 0.768 9.644 0.8 9.676 ;
  LAYER M1 ;
        RECT 0.832 7.188 0.864 9.696 ;
  LAYER M3 ;
        RECT 0.832 7.208 0.864 7.24 ;
  LAYER M1 ;
        RECT 0.896 7.188 0.928 9.696 ;
  LAYER M3 ;
        RECT 0.896 9.644 0.928 9.676 ;
  LAYER M1 ;
        RECT 0.96 7.188 0.992 9.696 ;
  LAYER M3 ;
        RECT 0.96 7.208 0.992 7.24 ;
  LAYER M1 ;
        RECT 1.024 7.188 1.056 9.696 ;
  LAYER M3 ;
        RECT 1.024 9.644 1.056 9.676 ;
  LAYER M1 ;
        RECT 1.088 7.188 1.12 9.696 ;
  LAYER M3 ;
        RECT 1.088 7.208 1.12 7.24 ;
  LAYER M1 ;
        RECT 1.152 7.188 1.184 9.696 ;
  LAYER M3 ;
        RECT 1.152 9.644 1.184 9.676 ;
  LAYER M1 ;
        RECT 1.216 7.188 1.248 9.696 ;
  LAYER M3 ;
        RECT 1.216 7.208 1.248 7.24 ;
  LAYER M1 ;
        RECT 1.28 7.188 1.312 9.696 ;
  LAYER M3 ;
        RECT 1.28 9.644 1.312 9.676 ;
  LAYER M1 ;
        RECT 1.344 7.188 1.376 9.696 ;
  LAYER M3 ;
        RECT 1.344 7.208 1.376 7.24 ;
  LAYER M1 ;
        RECT 1.408 7.188 1.44 9.696 ;
  LAYER M3 ;
        RECT 1.408 9.644 1.44 9.676 ;
  LAYER M1 ;
        RECT 1.472 7.188 1.504 9.696 ;
  LAYER M3 ;
        RECT 1.472 7.208 1.504 7.24 ;
  LAYER M1 ;
        RECT 1.536 7.188 1.568 9.696 ;
  LAYER M3 ;
        RECT 1.536 9.644 1.568 9.676 ;
  LAYER M1 ;
        RECT 1.6 7.188 1.632 9.696 ;
  LAYER M3 ;
        RECT 1.6 7.208 1.632 7.24 ;
  LAYER M1 ;
        RECT 1.664 7.188 1.696 9.696 ;
  LAYER M3 ;
        RECT 1.664 9.644 1.696 9.676 ;
  LAYER M1 ;
        RECT 1.728 7.188 1.76 9.696 ;
  LAYER M3 ;
        RECT 1.728 7.208 1.76 7.24 ;
  LAYER M1 ;
        RECT 1.792 7.188 1.824 9.696 ;
  LAYER M3 ;
        RECT 1.792 9.644 1.824 9.676 ;
  LAYER M1 ;
        RECT 1.856 7.188 1.888 9.696 ;
  LAYER M3 ;
        RECT 1.856 7.208 1.888 7.24 ;
  LAYER M1 ;
        RECT 1.92 7.188 1.952 9.696 ;
  LAYER M3 ;
        RECT 1.92 9.644 1.952 9.676 ;
  LAYER M1 ;
        RECT 1.984 7.188 2.016 9.696 ;
  LAYER M3 ;
        RECT 1.984 7.208 2.016 7.24 ;
  LAYER M1 ;
        RECT 2.048 7.188 2.08 9.696 ;
  LAYER M3 ;
        RECT 2.048 9.644 2.08 9.676 ;
  LAYER M1 ;
        RECT 2.112 7.188 2.144 9.696 ;
  LAYER M3 ;
        RECT 2.112 7.208 2.144 7.24 ;
  LAYER M1 ;
        RECT 2.176 7.188 2.208 9.696 ;
  LAYER M3 ;
        RECT 2.176 9.644 2.208 9.676 ;
  LAYER M1 ;
        RECT 2.24 7.188 2.272 9.696 ;
  LAYER M3 ;
        RECT 2.24 7.208 2.272 7.24 ;
  LAYER M1 ;
        RECT 2.304 7.188 2.336 9.696 ;
  LAYER M3 ;
        RECT 2.304 9.644 2.336 9.676 ;
  LAYER M1 ;
        RECT 2.368 7.188 2.4 9.696 ;
  LAYER M3 ;
        RECT 2.368 7.208 2.4 7.24 ;
  LAYER M1 ;
        RECT 2.432 7.188 2.464 9.696 ;
  LAYER M3 ;
        RECT 2.432 9.644 2.464 9.676 ;
  LAYER M1 ;
        RECT 2.496 7.188 2.528 9.696 ;
  LAYER M3 ;
        RECT 2.496 7.208 2.528 7.24 ;
  LAYER M1 ;
        RECT 2.56 7.188 2.592 9.696 ;
  LAYER M3 ;
        RECT 2.56 9.644 2.592 9.676 ;
  LAYER M1 ;
        RECT 2.624 7.188 2.656 9.696 ;
  LAYER M3 ;
        RECT 2.624 7.208 2.656 7.24 ;
  LAYER M1 ;
        RECT 2.688 7.188 2.72 9.696 ;
  LAYER M3 ;
        RECT 2.688 9.644 2.72 9.676 ;
  LAYER M1 ;
        RECT 2.752 7.188 2.784 9.696 ;
  LAYER M3 ;
        RECT 2.752 7.208 2.784 7.24 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 9.696 ;
  LAYER M3 ;
        RECT 2.816 9.644 2.848 9.676 ;
  LAYER M1 ;
        RECT 2.88 7.188 2.912 9.696 ;
  LAYER M3 ;
        RECT 2.88 7.208 2.912 7.24 ;
  LAYER M1 ;
        RECT 2.944 7.188 2.976 9.696 ;
  LAYER M3 ;
        RECT 2.944 9.644 2.976 9.676 ;
  LAYER M1 ;
        RECT 3.008 7.188 3.04 9.696 ;
  LAYER M3 ;
        RECT 3.008 7.208 3.04 7.24 ;
  LAYER M1 ;
        RECT 3.072 7.188 3.104 9.696 ;
  LAYER M3 ;
        RECT 3.072 9.644 3.104 9.676 ;
  LAYER M1 ;
        RECT 3.136 7.188 3.168 9.696 ;
  LAYER M3 ;
        RECT 0.768 7.272 0.8 7.304 ;
  LAYER M2 ;
        RECT 3.136 7.336 3.168 7.368 ;
  LAYER M2 ;
        RECT 0.768 7.4 0.8 7.432 ;
  LAYER M2 ;
        RECT 3.136 7.464 3.168 7.496 ;
  LAYER M2 ;
        RECT 0.768 7.528 0.8 7.56 ;
  LAYER M2 ;
        RECT 3.136 7.592 3.168 7.624 ;
  LAYER M2 ;
        RECT 0.768 7.656 0.8 7.688 ;
  LAYER M2 ;
        RECT 3.136 7.72 3.168 7.752 ;
  LAYER M2 ;
        RECT 0.768 7.784 0.8 7.816 ;
  LAYER M2 ;
        RECT 3.136 7.848 3.168 7.88 ;
  LAYER M2 ;
        RECT 0.768 7.912 0.8 7.944 ;
  LAYER M2 ;
        RECT 3.136 7.976 3.168 8.008 ;
  LAYER M2 ;
        RECT 0.768 8.04 0.8 8.072 ;
  LAYER M2 ;
        RECT 3.136 8.104 3.168 8.136 ;
  LAYER M2 ;
        RECT 0.768 8.168 0.8 8.2 ;
  LAYER M2 ;
        RECT 3.136 8.232 3.168 8.264 ;
  LAYER M2 ;
        RECT 0.768 8.296 0.8 8.328 ;
  LAYER M2 ;
        RECT 3.136 8.36 3.168 8.392 ;
  LAYER M2 ;
        RECT 0.768 8.424 0.8 8.456 ;
  LAYER M2 ;
        RECT 3.136 8.488 3.168 8.52 ;
  LAYER M2 ;
        RECT 0.768 8.552 0.8 8.584 ;
  LAYER M2 ;
        RECT 3.136 8.616 3.168 8.648 ;
  LAYER M2 ;
        RECT 0.768 8.68 0.8 8.712 ;
  LAYER M2 ;
        RECT 3.136 8.744 3.168 8.776 ;
  LAYER M2 ;
        RECT 0.768 8.808 0.8 8.84 ;
  LAYER M2 ;
        RECT 3.136 8.872 3.168 8.904 ;
  LAYER M2 ;
        RECT 0.768 8.936 0.8 8.968 ;
  LAYER M2 ;
        RECT 3.136 9 3.168 9.032 ;
  LAYER M2 ;
        RECT 0.768 9.064 0.8 9.096 ;
  LAYER M2 ;
        RECT 3.136 9.128 3.168 9.16 ;
  LAYER M2 ;
        RECT 0.768 9.192 0.8 9.224 ;
  LAYER M2 ;
        RECT 3.136 9.256 3.168 9.288 ;
  LAYER M2 ;
        RECT 0.768 9.32 0.8 9.352 ;
  LAYER M2 ;
        RECT 3.136 9.384 3.168 9.416 ;
  LAYER M2 ;
        RECT 0.768 9.448 0.8 9.48 ;
  LAYER M2 ;
        RECT 3.136 9.512 3.168 9.544 ;
  LAYER M2 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M1 ;
        RECT 0.768 10.296 0.8 12.804 ;
  LAYER M3 ;
        RECT 0.768 12.752 0.8 12.784 ;
  LAYER M1 ;
        RECT 0.832 10.296 0.864 12.804 ;
  LAYER M3 ;
        RECT 0.832 10.316 0.864 10.348 ;
  LAYER M1 ;
        RECT 0.896 10.296 0.928 12.804 ;
  LAYER M3 ;
        RECT 0.896 12.752 0.928 12.784 ;
  LAYER M1 ;
        RECT 0.96 10.296 0.992 12.804 ;
  LAYER M3 ;
        RECT 0.96 10.316 0.992 10.348 ;
  LAYER M1 ;
        RECT 1.024 10.296 1.056 12.804 ;
  LAYER M3 ;
        RECT 1.024 12.752 1.056 12.784 ;
  LAYER M1 ;
        RECT 1.088 10.296 1.12 12.804 ;
  LAYER M3 ;
        RECT 1.088 10.316 1.12 10.348 ;
  LAYER M1 ;
        RECT 1.152 10.296 1.184 12.804 ;
  LAYER M3 ;
        RECT 1.152 12.752 1.184 12.784 ;
  LAYER M1 ;
        RECT 1.216 10.296 1.248 12.804 ;
  LAYER M3 ;
        RECT 1.216 10.316 1.248 10.348 ;
  LAYER M1 ;
        RECT 1.28 10.296 1.312 12.804 ;
  LAYER M3 ;
        RECT 1.28 12.752 1.312 12.784 ;
  LAYER M1 ;
        RECT 1.344 10.296 1.376 12.804 ;
  LAYER M3 ;
        RECT 1.344 10.316 1.376 10.348 ;
  LAYER M1 ;
        RECT 1.408 10.296 1.44 12.804 ;
  LAYER M3 ;
        RECT 1.408 12.752 1.44 12.784 ;
  LAYER M1 ;
        RECT 1.472 10.296 1.504 12.804 ;
  LAYER M3 ;
        RECT 1.472 10.316 1.504 10.348 ;
  LAYER M1 ;
        RECT 1.536 10.296 1.568 12.804 ;
  LAYER M3 ;
        RECT 1.536 12.752 1.568 12.784 ;
  LAYER M1 ;
        RECT 1.6 10.296 1.632 12.804 ;
  LAYER M3 ;
        RECT 1.6 10.316 1.632 10.348 ;
  LAYER M1 ;
        RECT 1.664 10.296 1.696 12.804 ;
  LAYER M3 ;
        RECT 1.664 12.752 1.696 12.784 ;
  LAYER M1 ;
        RECT 1.728 10.296 1.76 12.804 ;
  LAYER M3 ;
        RECT 1.728 10.316 1.76 10.348 ;
  LAYER M1 ;
        RECT 1.792 10.296 1.824 12.804 ;
  LAYER M3 ;
        RECT 1.792 12.752 1.824 12.784 ;
  LAYER M1 ;
        RECT 1.856 10.296 1.888 12.804 ;
  LAYER M3 ;
        RECT 1.856 10.316 1.888 10.348 ;
  LAYER M1 ;
        RECT 1.92 10.296 1.952 12.804 ;
  LAYER M3 ;
        RECT 1.92 12.752 1.952 12.784 ;
  LAYER M1 ;
        RECT 1.984 10.296 2.016 12.804 ;
  LAYER M3 ;
        RECT 1.984 10.316 2.016 10.348 ;
  LAYER M1 ;
        RECT 2.048 10.296 2.08 12.804 ;
  LAYER M3 ;
        RECT 2.048 12.752 2.08 12.784 ;
  LAYER M1 ;
        RECT 2.112 10.296 2.144 12.804 ;
  LAYER M3 ;
        RECT 2.112 10.316 2.144 10.348 ;
  LAYER M1 ;
        RECT 2.176 10.296 2.208 12.804 ;
  LAYER M3 ;
        RECT 2.176 12.752 2.208 12.784 ;
  LAYER M1 ;
        RECT 2.24 10.296 2.272 12.804 ;
  LAYER M3 ;
        RECT 2.24 10.316 2.272 10.348 ;
  LAYER M1 ;
        RECT 2.304 10.296 2.336 12.804 ;
  LAYER M3 ;
        RECT 2.304 12.752 2.336 12.784 ;
  LAYER M1 ;
        RECT 2.368 10.296 2.4 12.804 ;
  LAYER M3 ;
        RECT 2.368 10.316 2.4 10.348 ;
  LAYER M1 ;
        RECT 2.432 10.296 2.464 12.804 ;
  LAYER M3 ;
        RECT 2.432 12.752 2.464 12.784 ;
  LAYER M1 ;
        RECT 2.496 10.296 2.528 12.804 ;
  LAYER M3 ;
        RECT 2.496 10.316 2.528 10.348 ;
  LAYER M1 ;
        RECT 2.56 10.296 2.592 12.804 ;
  LAYER M3 ;
        RECT 2.56 12.752 2.592 12.784 ;
  LAYER M1 ;
        RECT 2.624 10.296 2.656 12.804 ;
  LAYER M3 ;
        RECT 2.624 10.316 2.656 10.348 ;
  LAYER M1 ;
        RECT 2.688 10.296 2.72 12.804 ;
  LAYER M3 ;
        RECT 2.688 12.752 2.72 12.784 ;
  LAYER M1 ;
        RECT 2.752 10.296 2.784 12.804 ;
  LAYER M3 ;
        RECT 2.752 10.316 2.784 10.348 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 12.804 ;
  LAYER M3 ;
        RECT 2.816 12.752 2.848 12.784 ;
  LAYER M1 ;
        RECT 2.88 10.296 2.912 12.804 ;
  LAYER M3 ;
        RECT 2.88 10.316 2.912 10.348 ;
  LAYER M1 ;
        RECT 2.944 10.296 2.976 12.804 ;
  LAYER M3 ;
        RECT 2.944 12.752 2.976 12.784 ;
  LAYER M1 ;
        RECT 3.008 10.296 3.04 12.804 ;
  LAYER M3 ;
        RECT 3.008 10.316 3.04 10.348 ;
  LAYER M1 ;
        RECT 3.072 10.296 3.104 12.804 ;
  LAYER M3 ;
        RECT 3.072 12.752 3.104 12.784 ;
  LAYER M1 ;
        RECT 3.136 10.296 3.168 12.804 ;
  LAYER M3 ;
        RECT 0.768 10.38 0.8 10.412 ;
  LAYER M2 ;
        RECT 3.136 10.444 3.168 10.476 ;
  LAYER M2 ;
        RECT 0.768 10.508 0.8 10.54 ;
  LAYER M2 ;
        RECT 3.136 10.572 3.168 10.604 ;
  LAYER M2 ;
        RECT 0.768 10.636 0.8 10.668 ;
  LAYER M2 ;
        RECT 3.136 10.7 3.168 10.732 ;
  LAYER M2 ;
        RECT 0.768 10.764 0.8 10.796 ;
  LAYER M2 ;
        RECT 3.136 10.828 3.168 10.86 ;
  LAYER M2 ;
        RECT 0.768 10.892 0.8 10.924 ;
  LAYER M2 ;
        RECT 3.136 10.956 3.168 10.988 ;
  LAYER M2 ;
        RECT 0.768 11.02 0.8 11.052 ;
  LAYER M2 ;
        RECT 3.136 11.084 3.168 11.116 ;
  LAYER M2 ;
        RECT 0.768 11.148 0.8 11.18 ;
  LAYER M2 ;
        RECT 3.136 11.212 3.168 11.244 ;
  LAYER M2 ;
        RECT 0.768 11.276 0.8 11.308 ;
  LAYER M2 ;
        RECT 3.136 11.34 3.168 11.372 ;
  LAYER M2 ;
        RECT 0.768 11.404 0.8 11.436 ;
  LAYER M2 ;
        RECT 3.136 11.468 3.168 11.5 ;
  LAYER M2 ;
        RECT 0.768 11.532 0.8 11.564 ;
  LAYER M2 ;
        RECT 3.136 11.596 3.168 11.628 ;
  LAYER M2 ;
        RECT 0.768 11.66 0.8 11.692 ;
  LAYER M2 ;
        RECT 3.136 11.724 3.168 11.756 ;
  LAYER M2 ;
        RECT 0.768 11.788 0.8 11.82 ;
  LAYER M2 ;
        RECT 3.136 11.852 3.168 11.884 ;
  LAYER M2 ;
        RECT 0.768 11.916 0.8 11.948 ;
  LAYER M2 ;
        RECT 3.136 11.98 3.168 12.012 ;
  LAYER M2 ;
        RECT 0.768 12.044 0.8 12.076 ;
  LAYER M2 ;
        RECT 3.136 12.108 3.168 12.14 ;
  LAYER M2 ;
        RECT 0.768 12.172 0.8 12.204 ;
  LAYER M2 ;
        RECT 3.136 12.236 3.168 12.268 ;
  LAYER M2 ;
        RECT 0.768 12.3 0.8 12.332 ;
  LAYER M2 ;
        RECT 3.136 12.364 3.168 12.396 ;
  LAYER M2 ;
        RECT 0.768 12.428 0.8 12.46 ;
  LAYER M2 ;
        RECT 3.136 12.492 3.168 12.524 ;
  LAYER M2 ;
        RECT 0.768 12.556 0.8 12.588 ;
  LAYER M2 ;
        RECT 3.136 12.62 3.168 12.652 ;
  LAYER M2 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M1 ;
        RECT 0.768 13.404 0.8 15.912 ;
  LAYER M3 ;
        RECT 0.768 15.86 0.8 15.892 ;
  LAYER M1 ;
        RECT 0.832 13.404 0.864 15.912 ;
  LAYER M3 ;
        RECT 0.832 13.424 0.864 13.456 ;
  LAYER M1 ;
        RECT 0.896 13.404 0.928 15.912 ;
  LAYER M3 ;
        RECT 0.896 15.86 0.928 15.892 ;
  LAYER M1 ;
        RECT 0.96 13.404 0.992 15.912 ;
  LAYER M3 ;
        RECT 0.96 13.424 0.992 13.456 ;
  LAYER M1 ;
        RECT 1.024 13.404 1.056 15.912 ;
  LAYER M3 ;
        RECT 1.024 15.86 1.056 15.892 ;
  LAYER M1 ;
        RECT 1.088 13.404 1.12 15.912 ;
  LAYER M3 ;
        RECT 1.088 13.424 1.12 13.456 ;
  LAYER M1 ;
        RECT 1.152 13.404 1.184 15.912 ;
  LAYER M3 ;
        RECT 1.152 15.86 1.184 15.892 ;
  LAYER M1 ;
        RECT 1.216 13.404 1.248 15.912 ;
  LAYER M3 ;
        RECT 1.216 13.424 1.248 13.456 ;
  LAYER M1 ;
        RECT 1.28 13.404 1.312 15.912 ;
  LAYER M3 ;
        RECT 1.28 15.86 1.312 15.892 ;
  LAYER M1 ;
        RECT 1.344 13.404 1.376 15.912 ;
  LAYER M3 ;
        RECT 1.344 13.424 1.376 13.456 ;
  LAYER M1 ;
        RECT 1.408 13.404 1.44 15.912 ;
  LAYER M3 ;
        RECT 1.408 15.86 1.44 15.892 ;
  LAYER M1 ;
        RECT 1.472 13.404 1.504 15.912 ;
  LAYER M3 ;
        RECT 1.472 13.424 1.504 13.456 ;
  LAYER M1 ;
        RECT 1.536 13.404 1.568 15.912 ;
  LAYER M3 ;
        RECT 1.536 15.86 1.568 15.892 ;
  LAYER M1 ;
        RECT 1.6 13.404 1.632 15.912 ;
  LAYER M3 ;
        RECT 1.6 13.424 1.632 13.456 ;
  LAYER M1 ;
        RECT 1.664 13.404 1.696 15.912 ;
  LAYER M3 ;
        RECT 1.664 15.86 1.696 15.892 ;
  LAYER M1 ;
        RECT 1.728 13.404 1.76 15.912 ;
  LAYER M3 ;
        RECT 1.728 13.424 1.76 13.456 ;
  LAYER M1 ;
        RECT 1.792 13.404 1.824 15.912 ;
  LAYER M3 ;
        RECT 1.792 15.86 1.824 15.892 ;
  LAYER M1 ;
        RECT 1.856 13.404 1.888 15.912 ;
  LAYER M3 ;
        RECT 1.856 13.424 1.888 13.456 ;
  LAYER M1 ;
        RECT 1.92 13.404 1.952 15.912 ;
  LAYER M3 ;
        RECT 1.92 15.86 1.952 15.892 ;
  LAYER M1 ;
        RECT 1.984 13.404 2.016 15.912 ;
  LAYER M3 ;
        RECT 1.984 13.424 2.016 13.456 ;
  LAYER M1 ;
        RECT 2.048 13.404 2.08 15.912 ;
  LAYER M3 ;
        RECT 2.048 15.86 2.08 15.892 ;
  LAYER M1 ;
        RECT 2.112 13.404 2.144 15.912 ;
  LAYER M3 ;
        RECT 2.112 13.424 2.144 13.456 ;
  LAYER M1 ;
        RECT 2.176 13.404 2.208 15.912 ;
  LAYER M3 ;
        RECT 2.176 15.86 2.208 15.892 ;
  LAYER M1 ;
        RECT 2.24 13.404 2.272 15.912 ;
  LAYER M3 ;
        RECT 2.24 13.424 2.272 13.456 ;
  LAYER M1 ;
        RECT 2.304 13.404 2.336 15.912 ;
  LAYER M3 ;
        RECT 2.304 15.86 2.336 15.892 ;
  LAYER M1 ;
        RECT 2.368 13.404 2.4 15.912 ;
  LAYER M3 ;
        RECT 2.368 13.424 2.4 13.456 ;
  LAYER M1 ;
        RECT 2.432 13.404 2.464 15.912 ;
  LAYER M3 ;
        RECT 2.432 15.86 2.464 15.892 ;
  LAYER M1 ;
        RECT 2.496 13.404 2.528 15.912 ;
  LAYER M3 ;
        RECT 2.496 13.424 2.528 13.456 ;
  LAYER M1 ;
        RECT 2.56 13.404 2.592 15.912 ;
  LAYER M3 ;
        RECT 2.56 15.86 2.592 15.892 ;
  LAYER M1 ;
        RECT 2.624 13.404 2.656 15.912 ;
  LAYER M3 ;
        RECT 2.624 13.424 2.656 13.456 ;
  LAYER M1 ;
        RECT 2.688 13.404 2.72 15.912 ;
  LAYER M3 ;
        RECT 2.688 15.86 2.72 15.892 ;
  LAYER M1 ;
        RECT 2.752 13.404 2.784 15.912 ;
  LAYER M3 ;
        RECT 2.752 13.424 2.784 13.456 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 15.912 ;
  LAYER M3 ;
        RECT 2.816 15.86 2.848 15.892 ;
  LAYER M1 ;
        RECT 2.88 13.404 2.912 15.912 ;
  LAYER M3 ;
        RECT 2.88 13.424 2.912 13.456 ;
  LAYER M1 ;
        RECT 2.944 13.404 2.976 15.912 ;
  LAYER M3 ;
        RECT 2.944 15.86 2.976 15.892 ;
  LAYER M1 ;
        RECT 3.008 13.404 3.04 15.912 ;
  LAYER M3 ;
        RECT 3.008 13.424 3.04 13.456 ;
  LAYER M1 ;
        RECT 3.072 13.404 3.104 15.912 ;
  LAYER M3 ;
        RECT 3.072 15.86 3.104 15.892 ;
  LAYER M1 ;
        RECT 3.136 13.404 3.168 15.912 ;
  LAYER M3 ;
        RECT 0.768 13.488 0.8 13.52 ;
  LAYER M2 ;
        RECT 3.136 13.552 3.168 13.584 ;
  LAYER M2 ;
        RECT 0.768 13.616 0.8 13.648 ;
  LAYER M2 ;
        RECT 3.136 13.68 3.168 13.712 ;
  LAYER M2 ;
        RECT 0.768 13.744 0.8 13.776 ;
  LAYER M2 ;
        RECT 3.136 13.808 3.168 13.84 ;
  LAYER M2 ;
        RECT 0.768 13.872 0.8 13.904 ;
  LAYER M2 ;
        RECT 3.136 13.936 3.168 13.968 ;
  LAYER M2 ;
        RECT 0.768 14 0.8 14.032 ;
  LAYER M2 ;
        RECT 3.136 14.064 3.168 14.096 ;
  LAYER M2 ;
        RECT 0.768 14.128 0.8 14.16 ;
  LAYER M2 ;
        RECT 3.136 14.192 3.168 14.224 ;
  LAYER M2 ;
        RECT 0.768 14.256 0.8 14.288 ;
  LAYER M2 ;
        RECT 3.136 14.32 3.168 14.352 ;
  LAYER M2 ;
        RECT 0.768 14.384 0.8 14.416 ;
  LAYER M2 ;
        RECT 3.136 14.448 3.168 14.48 ;
  LAYER M2 ;
        RECT 0.768 14.512 0.8 14.544 ;
  LAYER M2 ;
        RECT 3.136 14.576 3.168 14.608 ;
  LAYER M2 ;
        RECT 0.768 14.64 0.8 14.672 ;
  LAYER M2 ;
        RECT 3.136 14.704 3.168 14.736 ;
  LAYER M2 ;
        RECT 0.768 14.768 0.8 14.8 ;
  LAYER M2 ;
        RECT 3.136 14.832 3.168 14.864 ;
  LAYER M2 ;
        RECT 0.768 14.896 0.8 14.928 ;
  LAYER M2 ;
        RECT 3.136 14.96 3.168 14.992 ;
  LAYER M2 ;
        RECT 0.768 15.024 0.8 15.056 ;
  LAYER M2 ;
        RECT 3.136 15.088 3.168 15.12 ;
  LAYER M2 ;
        RECT 0.768 15.152 0.8 15.184 ;
  LAYER M2 ;
        RECT 3.136 15.216 3.168 15.248 ;
  LAYER M2 ;
        RECT 0.768 15.28 0.8 15.312 ;
  LAYER M2 ;
        RECT 3.136 15.344 3.168 15.376 ;
  LAYER M2 ;
        RECT 0.768 15.408 0.8 15.44 ;
  LAYER M2 ;
        RECT 3.136 15.472 3.168 15.504 ;
  LAYER M2 ;
        RECT 0.768 15.536 0.8 15.568 ;
  LAYER M2 ;
        RECT 3.136 15.6 3.168 15.632 ;
  LAYER M2 ;
        RECT 0.768 15.664 0.8 15.696 ;
  LAYER M2 ;
        RECT 3.136 15.728 3.168 15.76 ;
  LAYER M2 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M1 ;
        RECT 0.768 16.512 0.8 19.02 ;
  LAYER M3 ;
        RECT 0.768 18.968 0.8 19 ;
  LAYER M1 ;
        RECT 0.832 16.512 0.864 19.02 ;
  LAYER M3 ;
        RECT 0.832 16.532 0.864 16.564 ;
  LAYER M1 ;
        RECT 0.896 16.512 0.928 19.02 ;
  LAYER M3 ;
        RECT 0.896 18.968 0.928 19 ;
  LAYER M1 ;
        RECT 0.96 16.512 0.992 19.02 ;
  LAYER M3 ;
        RECT 0.96 16.532 0.992 16.564 ;
  LAYER M1 ;
        RECT 1.024 16.512 1.056 19.02 ;
  LAYER M3 ;
        RECT 1.024 18.968 1.056 19 ;
  LAYER M1 ;
        RECT 1.088 16.512 1.12 19.02 ;
  LAYER M3 ;
        RECT 1.088 16.532 1.12 16.564 ;
  LAYER M1 ;
        RECT 1.152 16.512 1.184 19.02 ;
  LAYER M3 ;
        RECT 1.152 18.968 1.184 19 ;
  LAYER M1 ;
        RECT 1.216 16.512 1.248 19.02 ;
  LAYER M3 ;
        RECT 1.216 16.532 1.248 16.564 ;
  LAYER M1 ;
        RECT 1.28 16.512 1.312 19.02 ;
  LAYER M3 ;
        RECT 1.28 18.968 1.312 19 ;
  LAYER M1 ;
        RECT 1.344 16.512 1.376 19.02 ;
  LAYER M3 ;
        RECT 1.344 16.532 1.376 16.564 ;
  LAYER M1 ;
        RECT 1.408 16.512 1.44 19.02 ;
  LAYER M3 ;
        RECT 1.408 18.968 1.44 19 ;
  LAYER M1 ;
        RECT 1.472 16.512 1.504 19.02 ;
  LAYER M3 ;
        RECT 1.472 16.532 1.504 16.564 ;
  LAYER M1 ;
        RECT 1.536 16.512 1.568 19.02 ;
  LAYER M3 ;
        RECT 1.536 18.968 1.568 19 ;
  LAYER M1 ;
        RECT 1.6 16.512 1.632 19.02 ;
  LAYER M3 ;
        RECT 1.6 16.532 1.632 16.564 ;
  LAYER M1 ;
        RECT 1.664 16.512 1.696 19.02 ;
  LAYER M3 ;
        RECT 1.664 18.968 1.696 19 ;
  LAYER M1 ;
        RECT 1.728 16.512 1.76 19.02 ;
  LAYER M3 ;
        RECT 1.728 16.532 1.76 16.564 ;
  LAYER M1 ;
        RECT 1.792 16.512 1.824 19.02 ;
  LAYER M3 ;
        RECT 1.792 18.968 1.824 19 ;
  LAYER M1 ;
        RECT 1.856 16.512 1.888 19.02 ;
  LAYER M3 ;
        RECT 1.856 16.532 1.888 16.564 ;
  LAYER M1 ;
        RECT 1.92 16.512 1.952 19.02 ;
  LAYER M3 ;
        RECT 1.92 18.968 1.952 19 ;
  LAYER M1 ;
        RECT 1.984 16.512 2.016 19.02 ;
  LAYER M3 ;
        RECT 1.984 16.532 2.016 16.564 ;
  LAYER M1 ;
        RECT 2.048 16.512 2.08 19.02 ;
  LAYER M3 ;
        RECT 2.048 18.968 2.08 19 ;
  LAYER M1 ;
        RECT 2.112 16.512 2.144 19.02 ;
  LAYER M3 ;
        RECT 2.112 16.532 2.144 16.564 ;
  LAYER M1 ;
        RECT 2.176 16.512 2.208 19.02 ;
  LAYER M3 ;
        RECT 2.176 18.968 2.208 19 ;
  LAYER M1 ;
        RECT 2.24 16.512 2.272 19.02 ;
  LAYER M3 ;
        RECT 2.24 16.532 2.272 16.564 ;
  LAYER M1 ;
        RECT 2.304 16.512 2.336 19.02 ;
  LAYER M3 ;
        RECT 2.304 18.968 2.336 19 ;
  LAYER M1 ;
        RECT 2.368 16.512 2.4 19.02 ;
  LAYER M3 ;
        RECT 2.368 16.532 2.4 16.564 ;
  LAYER M1 ;
        RECT 2.432 16.512 2.464 19.02 ;
  LAYER M3 ;
        RECT 2.432 18.968 2.464 19 ;
  LAYER M1 ;
        RECT 2.496 16.512 2.528 19.02 ;
  LAYER M3 ;
        RECT 2.496 16.532 2.528 16.564 ;
  LAYER M1 ;
        RECT 2.56 16.512 2.592 19.02 ;
  LAYER M3 ;
        RECT 2.56 18.968 2.592 19 ;
  LAYER M1 ;
        RECT 2.624 16.512 2.656 19.02 ;
  LAYER M3 ;
        RECT 2.624 16.532 2.656 16.564 ;
  LAYER M1 ;
        RECT 2.688 16.512 2.72 19.02 ;
  LAYER M3 ;
        RECT 2.688 18.968 2.72 19 ;
  LAYER M1 ;
        RECT 2.752 16.512 2.784 19.02 ;
  LAYER M3 ;
        RECT 2.752 16.532 2.784 16.564 ;
  LAYER M1 ;
        RECT 2.816 16.512 2.848 19.02 ;
  LAYER M3 ;
        RECT 2.816 18.968 2.848 19 ;
  LAYER M1 ;
        RECT 2.88 16.512 2.912 19.02 ;
  LAYER M3 ;
        RECT 2.88 16.532 2.912 16.564 ;
  LAYER M1 ;
        RECT 2.944 16.512 2.976 19.02 ;
  LAYER M3 ;
        RECT 2.944 18.968 2.976 19 ;
  LAYER M1 ;
        RECT 3.008 16.512 3.04 19.02 ;
  LAYER M3 ;
        RECT 3.008 16.532 3.04 16.564 ;
  LAYER M1 ;
        RECT 3.072 16.512 3.104 19.02 ;
  LAYER M3 ;
        RECT 3.072 18.968 3.104 19 ;
  LAYER M1 ;
        RECT 3.136 16.512 3.168 19.02 ;
  LAYER M3 ;
        RECT 0.768 16.596 0.8 16.628 ;
  LAYER M2 ;
        RECT 3.136 16.66 3.168 16.692 ;
  LAYER M2 ;
        RECT 0.768 16.724 0.8 16.756 ;
  LAYER M2 ;
        RECT 3.136 16.788 3.168 16.82 ;
  LAYER M2 ;
        RECT 0.768 16.852 0.8 16.884 ;
  LAYER M2 ;
        RECT 3.136 16.916 3.168 16.948 ;
  LAYER M2 ;
        RECT 0.768 16.98 0.8 17.012 ;
  LAYER M2 ;
        RECT 3.136 17.044 3.168 17.076 ;
  LAYER M2 ;
        RECT 0.768 17.108 0.8 17.14 ;
  LAYER M2 ;
        RECT 3.136 17.172 3.168 17.204 ;
  LAYER M2 ;
        RECT 0.768 17.236 0.8 17.268 ;
  LAYER M2 ;
        RECT 3.136 17.3 3.168 17.332 ;
  LAYER M2 ;
        RECT 0.768 17.364 0.8 17.396 ;
  LAYER M2 ;
        RECT 3.136 17.428 3.168 17.46 ;
  LAYER M2 ;
        RECT 0.768 17.492 0.8 17.524 ;
  LAYER M2 ;
        RECT 3.136 17.556 3.168 17.588 ;
  LAYER M2 ;
        RECT 0.768 17.62 0.8 17.652 ;
  LAYER M2 ;
        RECT 3.136 17.684 3.168 17.716 ;
  LAYER M2 ;
        RECT 0.768 17.748 0.8 17.78 ;
  LAYER M2 ;
        RECT 3.136 17.812 3.168 17.844 ;
  LAYER M2 ;
        RECT 0.768 17.876 0.8 17.908 ;
  LAYER M2 ;
        RECT 3.136 17.94 3.168 17.972 ;
  LAYER M2 ;
        RECT 0.768 18.004 0.8 18.036 ;
  LAYER M2 ;
        RECT 3.136 18.068 3.168 18.1 ;
  LAYER M2 ;
        RECT 0.768 18.132 0.8 18.164 ;
  LAYER M2 ;
        RECT 3.136 18.196 3.168 18.228 ;
  LAYER M2 ;
        RECT 0.768 18.26 0.8 18.292 ;
  LAYER M2 ;
        RECT 3.136 18.324 3.168 18.356 ;
  LAYER M2 ;
        RECT 0.768 18.388 0.8 18.42 ;
  LAYER M2 ;
        RECT 3.136 18.452 3.168 18.484 ;
  LAYER M2 ;
        RECT 0.768 18.516 0.8 18.548 ;
  LAYER M2 ;
        RECT 3.136 18.58 3.168 18.612 ;
  LAYER M2 ;
        RECT 0.768 18.644 0.8 18.676 ;
  LAYER M2 ;
        RECT 3.136 18.708 3.168 18.74 ;
  LAYER M2 ;
        RECT 0.768 18.772 0.8 18.804 ;
  LAYER M2 ;
        RECT 3.136 18.836 3.168 18.868 ;
  LAYER M2 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M1 ;
        RECT 0.768 19.62 0.8 22.128 ;
  LAYER M3 ;
        RECT 0.768 22.076 0.8 22.108 ;
  LAYER M1 ;
        RECT 0.832 19.62 0.864 22.128 ;
  LAYER M3 ;
        RECT 0.832 19.64 0.864 19.672 ;
  LAYER M1 ;
        RECT 0.896 19.62 0.928 22.128 ;
  LAYER M3 ;
        RECT 0.896 22.076 0.928 22.108 ;
  LAYER M1 ;
        RECT 0.96 19.62 0.992 22.128 ;
  LAYER M3 ;
        RECT 0.96 19.64 0.992 19.672 ;
  LAYER M1 ;
        RECT 1.024 19.62 1.056 22.128 ;
  LAYER M3 ;
        RECT 1.024 22.076 1.056 22.108 ;
  LAYER M1 ;
        RECT 1.088 19.62 1.12 22.128 ;
  LAYER M3 ;
        RECT 1.088 19.64 1.12 19.672 ;
  LAYER M1 ;
        RECT 1.152 19.62 1.184 22.128 ;
  LAYER M3 ;
        RECT 1.152 22.076 1.184 22.108 ;
  LAYER M1 ;
        RECT 1.216 19.62 1.248 22.128 ;
  LAYER M3 ;
        RECT 1.216 19.64 1.248 19.672 ;
  LAYER M1 ;
        RECT 1.28 19.62 1.312 22.128 ;
  LAYER M3 ;
        RECT 1.28 22.076 1.312 22.108 ;
  LAYER M1 ;
        RECT 1.344 19.62 1.376 22.128 ;
  LAYER M3 ;
        RECT 1.344 19.64 1.376 19.672 ;
  LAYER M1 ;
        RECT 1.408 19.62 1.44 22.128 ;
  LAYER M3 ;
        RECT 1.408 22.076 1.44 22.108 ;
  LAYER M1 ;
        RECT 1.472 19.62 1.504 22.128 ;
  LAYER M3 ;
        RECT 1.472 19.64 1.504 19.672 ;
  LAYER M1 ;
        RECT 1.536 19.62 1.568 22.128 ;
  LAYER M3 ;
        RECT 1.536 22.076 1.568 22.108 ;
  LAYER M1 ;
        RECT 1.6 19.62 1.632 22.128 ;
  LAYER M3 ;
        RECT 1.6 19.64 1.632 19.672 ;
  LAYER M1 ;
        RECT 1.664 19.62 1.696 22.128 ;
  LAYER M3 ;
        RECT 1.664 22.076 1.696 22.108 ;
  LAYER M1 ;
        RECT 1.728 19.62 1.76 22.128 ;
  LAYER M3 ;
        RECT 1.728 19.64 1.76 19.672 ;
  LAYER M1 ;
        RECT 1.792 19.62 1.824 22.128 ;
  LAYER M3 ;
        RECT 1.792 22.076 1.824 22.108 ;
  LAYER M1 ;
        RECT 1.856 19.62 1.888 22.128 ;
  LAYER M3 ;
        RECT 1.856 19.64 1.888 19.672 ;
  LAYER M1 ;
        RECT 1.92 19.62 1.952 22.128 ;
  LAYER M3 ;
        RECT 1.92 22.076 1.952 22.108 ;
  LAYER M1 ;
        RECT 1.984 19.62 2.016 22.128 ;
  LAYER M3 ;
        RECT 1.984 19.64 2.016 19.672 ;
  LAYER M1 ;
        RECT 2.048 19.62 2.08 22.128 ;
  LAYER M3 ;
        RECT 2.048 22.076 2.08 22.108 ;
  LAYER M1 ;
        RECT 2.112 19.62 2.144 22.128 ;
  LAYER M3 ;
        RECT 2.112 19.64 2.144 19.672 ;
  LAYER M1 ;
        RECT 2.176 19.62 2.208 22.128 ;
  LAYER M3 ;
        RECT 2.176 22.076 2.208 22.108 ;
  LAYER M1 ;
        RECT 2.24 19.62 2.272 22.128 ;
  LAYER M3 ;
        RECT 2.24 19.64 2.272 19.672 ;
  LAYER M1 ;
        RECT 2.304 19.62 2.336 22.128 ;
  LAYER M3 ;
        RECT 2.304 22.076 2.336 22.108 ;
  LAYER M1 ;
        RECT 2.368 19.62 2.4 22.128 ;
  LAYER M3 ;
        RECT 2.368 19.64 2.4 19.672 ;
  LAYER M1 ;
        RECT 2.432 19.62 2.464 22.128 ;
  LAYER M3 ;
        RECT 2.432 22.076 2.464 22.108 ;
  LAYER M1 ;
        RECT 2.496 19.62 2.528 22.128 ;
  LAYER M3 ;
        RECT 2.496 19.64 2.528 19.672 ;
  LAYER M1 ;
        RECT 2.56 19.62 2.592 22.128 ;
  LAYER M3 ;
        RECT 2.56 22.076 2.592 22.108 ;
  LAYER M1 ;
        RECT 2.624 19.62 2.656 22.128 ;
  LAYER M3 ;
        RECT 2.624 19.64 2.656 19.672 ;
  LAYER M1 ;
        RECT 2.688 19.62 2.72 22.128 ;
  LAYER M3 ;
        RECT 2.688 22.076 2.72 22.108 ;
  LAYER M1 ;
        RECT 2.752 19.62 2.784 22.128 ;
  LAYER M3 ;
        RECT 2.752 19.64 2.784 19.672 ;
  LAYER M1 ;
        RECT 2.816 19.62 2.848 22.128 ;
  LAYER M3 ;
        RECT 2.816 22.076 2.848 22.108 ;
  LAYER M1 ;
        RECT 2.88 19.62 2.912 22.128 ;
  LAYER M3 ;
        RECT 2.88 19.64 2.912 19.672 ;
  LAYER M1 ;
        RECT 2.944 19.62 2.976 22.128 ;
  LAYER M3 ;
        RECT 2.944 22.076 2.976 22.108 ;
  LAYER M1 ;
        RECT 3.008 19.62 3.04 22.128 ;
  LAYER M3 ;
        RECT 3.008 19.64 3.04 19.672 ;
  LAYER M1 ;
        RECT 3.072 19.62 3.104 22.128 ;
  LAYER M3 ;
        RECT 3.072 22.076 3.104 22.108 ;
  LAYER M1 ;
        RECT 3.136 19.62 3.168 22.128 ;
  LAYER M3 ;
        RECT 0.768 19.704 0.8 19.736 ;
  LAYER M2 ;
        RECT 3.136 19.768 3.168 19.8 ;
  LAYER M2 ;
        RECT 0.768 19.832 0.8 19.864 ;
  LAYER M2 ;
        RECT 3.136 19.896 3.168 19.928 ;
  LAYER M2 ;
        RECT 0.768 19.96 0.8 19.992 ;
  LAYER M2 ;
        RECT 3.136 20.024 3.168 20.056 ;
  LAYER M2 ;
        RECT 0.768 20.088 0.8 20.12 ;
  LAYER M2 ;
        RECT 3.136 20.152 3.168 20.184 ;
  LAYER M2 ;
        RECT 0.768 20.216 0.8 20.248 ;
  LAYER M2 ;
        RECT 3.136 20.28 3.168 20.312 ;
  LAYER M2 ;
        RECT 0.768 20.344 0.8 20.376 ;
  LAYER M2 ;
        RECT 3.136 20.408 3.168 20.44 ;
  LAYER M2 ;
        RECT 0.768 20.472 0.8 20.504 ;
  LAYER M2 ;
        RECT 3.136 20.536 3.168 20.568 ;
  LAYER M2 ;
        RECT 0.768 20.6 0.8 20.632 ;
  LAYER M2 ;
        RECT 3.136 20.664 3.168 20.696 ;
  LAYER M2 ;
        RECT 0.768 20.728 0.8 20.76 ;
  LAYER M2 ;
        RECT 3.136 20.792 3.168 20.824 ;
  LAYER M2 ;
        RECT 0.768 20.856 0.8 20.888 ;
  LAYER M2 ;
        RECT 3.136 20.92 3.168 20.952 ;
  LAYER M2 ;
        RECT 0.768 20.984 0.8 21.016 ;
  LAYER M2 ;
        RECT 3.136 21.048 3.168 21.08 ;
  LAYER M2 ;
        RECT 0.768 21.112 0.8 21.144 ;
  LAYER M2 ;
        RECT 3.136 21.176 3.168 21.208 ;
  LAYER M2 ;
        RECT 0.768 21.24 0.8 21.272 ;
  LAYER M2 ;
        RECT 3.136 21.304 3.168 21.336 ;
  LAYER M2 ;
        RECT 0.768 21.368 0.8 21.4 ;
  LAYER M2 ;
        RECT 3.136 21.432 3.168 21.464 ;
  LAYER M2 ;
        RECT 0.768 21.496 0.8 21.528 ;
  LAYER M2 ;
        RECT 3.136 21.56 3.168 21.592 ;
  LAYER M2 ;
        RECT 0.768 21.624 0.8 21.656 ;
  LAYER M2 ;
        RECT 3.136 21.688 3.168 21.72 ;
  LAYER M2 ;
        RECT 0.768 21.752 0.8 21.784 ;
  LAYER M2 ;
        RECT 3.136 21.816 3.168 21.848 ;
  LAYER M2 ;
        RECT 0.768 21.88 0.8 21.912 ;
  LAYER M2 ;
        RECT 3.136 21.944 3.168 21.976 ;
  LAYER M2 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M1 ;
        RECT 0.768 22.728 0.8 25.236 ;
  LAYER M3 ;
        RECT 0.768 25.184 0.8 25.216 ;
  LAYER M1 ;
        RECT 0.832 22.728 0.864 25.236 ;
  LAYER M3 ;
        RECT 0.832 22.748 0.864 22.78 ;
  LAYER M1 ;
        RECT 0.896 22.728 0.928 25.236 ;
  LAYER M3 ;
        RECT 0.896 25.184 0.928 25.216 ;
  LAYER M1 ;
        RECT 0.96 22.728 0.992 25.236 ;
  LAYER M3 ;
        RECT 0.96 22.748 0.992 22.78 ;
  LAYER M1 ;
        RECT 1.024 22.728 1.056 25.236 ;
  LAYER M3 ;
        RECT 1.024 25.184 1.056 25.216 ;
  LAYER M1 ;
        RECT 1.088 22.728 1.12 25.236 ;
  LAYER M3 ;
        RECT 1.088 22.748 1.12 22.78 ;
  LAYER M1 ;
        RECT 1.152 22.728 1.184 25.236 ;
  LAYER M3 ;
        RECT 1.152 25.184 1.184 25.216 ;
  LAYER M1 ;
        RECT 1.216 22.728 1.248 25.236 ;
  LAYER M3 ;
        RECT 1.216 22.748 1.248 22.78 ;
  LAYER M1 ;
        RECT 1.28 22.728 1.312 25.236 ;
  LAYER M3 ;
        RECT 1.28 25.184 1.312 25.216 ;
  LAYER M1 ;
        RECT 1.344 22.728 1.376 25.236 ;
  LAYER M3 ;
        RECT 1.344 22.748 1.376 22.78 ;
  LAYER M1 ;
        RECT 1.408 22.728 1.44 25.236 ;
  LAYER M3 ;
        RECT 1.408 25.184 1.44 25.216 ;
  LAYER M1 ;
        RECT 1.472 22.728 1.504 25.236 ;
  LAYER M3 ;
        RECT 1.472 22.748 1.504 22.78 ;
  LAYER M1 ;
        RECT 1.536 22.728 1.568 25.236 ;
  LAYER M3 ;
        RECT 1.536 25.184 1.568 25.216 ;
  LAYER M1 ;
        RECT 1.6 22.728 1.632 25.236 ;
  LAYER M3 ;
        RECT 1.6 22.748 1.632 22.78 ;
  LAYER M1 ;
        RECT 1.664 22.728 1.696 25.236 ;
  LAYER M3 ;
        RECT 1.664 25.184 1.696 25.216 ;
  LAYER M1 ;
        RECT 1.728 22.728 1.76 25.236 ;
  LAYER M3 ;
        RECT 1.728 22.748 1.76 22.78 ;
  LAYER M1 ;
        RECT 1.792 22.728 1.824 25.236 ;
  LAYER M3 ;
        RECT 1.792 25.184 1.824 25.216 ;
  LAYER M1 ;
        RECT 1.856 22.728 1.888 25.236 ;
  LAYER M3 ;
        RECT 1.856 22.748 1.888 22.78 ;
  LAYER M1 ;
        RECT 1.92 22.728 1.952 25.236 ;
  LAYER M3 ;
        RECT 1.92 25.184 1.952 25.216 ;
  LAYER M1 ;
        RECT 1.984 22.728 2.016 25.236 ;
  LAYER M3 ;
        RECT 1.984 22.748 2.016 22.78 ;
  LAYER M1 ;
        RECT 2.048 22.728 2.08 25.236 ;
  LAYER M3 ;
        RECT 2.048 25.184 2.08 25.216 ;
  LAYER M1 ;
        RECT 2.112 22.728 2.144 25.236 ;
  LAYER M3 ;
        RECT 2.112 22.748 2.144 22.78 ;
  LAYER M1 ;
        RECT 2.176 22.728 2.208 25.236 ;
  LAYER M3 ;
        RECT 2.176 25.184 2.208 25.216 ;
  LAYER M1 ;
        RECT 2.24 22.728 2.272 25.236 ;
  LAYER M3 ;
        RECT 2.24 22.748 2.272 22.78 ;
  LAYER M1 ;
        RECT 2.304 22.728 2.336 25.236 ;
  LAYER M3 ;
        RECT 2.304 25.184 2.336 25.216 ;
  LAYER M1 ;
        RECT 2.368 22.728 2.4 25.236 ;
  LAYER M3 ;
        RECT 2.368 22.748 2.4 22.78 ;
  LAYER M1 ;
        RECT 2.432 22.728 2.464 25.236 ;
  LAYER M3 ;
        RECT 2.432 25.184 2.464 25.216 ;
  LAYER M1 ;
        RECT 2.496 22.728 2.528 25.236 ;
  LAYER M3 ;
        RECT 2.496 22.748 2.528 22.78 ;
  LAYER M1 ;
        RECT 2.56 22.728 2.592 25.236 ;
  LAYER M3 ;
        RECT 2.56 25.184 2.592 25.216 ;
  LAYER M1 ;
        RECT 2.624 22.728 2.656 25.236 ;
  LAYER M3 ;
        RECT 2.624 22.748 2.656 22.78 ;
  LAYER M1 ;
        RECT 2.688 22.728 2.72 25.236 ;
  LAYER M3 ;
        RECT 2.688 25.184 2.72 25.216 ;
  LAYER M1 ;
        RECT 2.752 22.728 2.784 25.236 ;
  LAYER M3 ;
        RECT 2.752 22.748 2.784 22.78 ;
  LAYER M1 ;
        RECT 2.816 22.728 2.848 25.236 ;
  LAYER M3 ;
        RECT 2.816 25.184 2.848 25.216 ;
  LAYER M1 ;
        RECT 2.88 22.728 2.912 25.236 ;
  LAYER M3 ;
        RECT 2.88 22.748 2.912 22.78 ;
  LAYER M1 ;
        RECT 2.944 22.728 2.976 25.236 ;
  LAYER M3 ;
        RECT 2.944 25.184 2.976 25.216 ;
  LAYER M1 ;
        RECT 3.008 22.728 3.04 25.236 ;
  LAYER M3 ;
        RECT 3.008 22.748 3.04 22.78 ;
  LAYER M1 ;
        RECT 3.072 22.728 3.104 25.236 ;
  LAYER M3 ;
        RECT 3.072 25.184 3.104 25.216 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 25.236 ;
  LAYER M3 ;
        RECT 0.768 22.812 0.8 22.844 ;
  LAYER M2 ;
        RECT 3.136 22.876 3.168 22.908 ;
  LAYER M2 ;
        RECT 0.768 22.94 0.8 22.972 ;
  LAYER M2 ;
        RECT 3.136 23.004 3.168 23.036 ;
  LAYER M2 ;
        RECT 0.768 23.068 0.8 23.1 ;
  LAYER M2 ;
        RECT 3.136 23.132 3.168 23.164 ;
  LAYER M2 ;
        RECT 0.768 23.196 0.8 23.228 ;
  LAYER M2 ;
        RECT 3.136 23.26 3.168 23.292 ;
  LAYER M2 ;
        RECT 0.768 23.324 0.8 23.356 ;
  LAYER M2 ;
        RECT 3.136 23.388 3.168 23.42 ;
  LAYER M2 ;
        RECT 0.768 23.452 0.8 23.484 ;
  LAYER M2 ;
        RECT 3.136 23.516 3.168 23.548 ;
  LAYER M2 ;
        RECT 0.768 23.58 0.8 23.612 ;
  LAYER M2 ;
        RECT 3.136 23.644 3.168 23.676 ;
  LAYER M2 ;
        RECT 0.768 23.708 0.8 23.74 ;
  LAYER M2 ;
        RECT 3.136 23.772 3.168 23.804 ;
  LAYER M2 ;
        RECT 0.768 23.836 0.8 23.868 ;
  LAYER M2 ;
        RECT 3.136 23.9 3.168 23.932 ;
  LAYER M2 ;
        RECT 0.768 23.964 0.8 23.996 ;
  LAYER M2 ;
        RECT 3.136 24.028 3.168 24.06 ;
  LAYER M2 ;
        RECT 0.768 24.092 0.8 24.124 ;
  LAYER M2 ;
        RECT 3.136 24.156 3.168 24.188 ;
  LAYER M2 ;
        RECT 0.768 24.22 0.8 24.252 ;
  LAYER M2 ;
        RECT 3.136 24.284 3.168 24.316 ;
  LAYER M2 ;
        RECT 0.768 24.348 0.8 24.38 ;
  LAYER M2 ;
        RECT 3.136 24.412 3.168 24.444 ;
  LAYER M2 ;
        RECT 0.768 24.476 0.8 24.508 ;
  LAYER M2 ;
        RECT 3.136 24.54 3.168 24.572 ;
  LAYER M2 ;
        RECT 0.768 24.604 0.8 24.636 ;
  LAYER M2 ;
        RECT 3.136 24.668 3.168 24.7 ;
  LAYER M2 ;
        RECT 0.768 24.732 0.8 24.764 ;
  LAYER M2 ;
        RECT 3.136 24.796 3.168 24.828 ;
  LAYER M2 ;
        RECT 0.768 24.86 0.8 24.892 ;
  LAYER M2 ;
        RECT 3.136 24.924 3.168 24.956 ;
  LAYER M2 ;
        RECT 0.768 24.988 0.8 25.02 ;
  LAYER M2 ;
        RECT 3.136 25.052 3.168 25.084 ;
  LAYER M2 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M1 ;
        RECT 4.064 0.972 4.096 3.48 ;
  LAYER M3 ;
        RECT 4.064 3.428 4.096 3.46 ;
  LAYER M1 ;
        RECT 4.128 0.972 4.16 3.48 ;
  LAYER M3 ;
        RECT 4.128 0.992 4.16 1.024 ;
  LAYER M1 ;
        RECT 4.192 0.972 4.224 3.48 ;
  LAYER M3 ;
        RECT 4.192 3.428 4.224 3.46 ;
  LAYER M1 ;
        RECT 4.256 0.972 4.288 3.48 ;
  LAYER M3 ;
        RECT 4.256 0.992 4.288 1.024 ;
  LAYER M1 ;
        RECT 4.32 0.972 4.352 3.48 ;
  LAYER M3 ;
        RECT 4.32 3.428 4.352 3.46 ;
  LAYER M1 ;
        RECT 4.384 0.972 4.416 3.48 ;
  LAYER M3 ;
        RECT 4.384 0.992 4.416 1.024 ;
  LAYER M1 ;
        RECT 4.448 0.972 4.48 3.48 ;
  LAYER M3 ;
        RECT 4.448 3.428 4.48 3.46 ;
  LAYER M1 ;
        RECT 4.512 0.972 4.544 3.48 ;
  LAYER M3 ;
        RECT 4.512 0.992 4.544 1.024 ;
  LAYER M1 ;
        RECT 4.576 0.972 4.608 3.48 ;
  LAYER M3 ;
        RECT 4.576 3.428 4.608 3.46 ;
  LAYER M1 ;
        RECT 4.64 0.972 4.672 3.48 ;
  LAYER M3 ;
        RECT 4.64 0.992 4.672 1.024 ;
  LAYER M1 ;
        RECT 4.704 0.972 4.736 3.48 ;
  LAYER M3 ;
        RECT 4.704 3.428 4.736 3.46 ;
  LAYER M1 ;
        RECT 4.768 0.972 4.8 3.48 ;
  LAYER M3 ;
        RECT 4.768 0.992 4.8 1.024 ;
  LAYER M1 ;
        RECT 4.832 0.972 4.864 3.48 ;
  LAYER M3 ;
        RECT 4.832 3.428 4.864 3.46 ;
  LAYER M1 ;
        RECT 4.896 0.972 4.928 3.48 ;
  LAYER M3 ;
        RECT 4.896 0.992 4.928 1.024 ;
  LAYER M1 ;
        RECT 4.96 0.972 4.992 3.48 ;
  LAYER M3 ;
        RECT 4.96 3.428 4.992 3.46 ;
  LAYER M1 ;
        RECT 5.024 0.972 5.056 3.48 ;
  LAYER M3 ;
        RECT 5.024 0.992 5.056 1.024 ;
  LAYER M1 ;
        RECT 5.088 0.972 5.12 3.48 ;
  LAYER M3 ;
        RECT 5.088 3.428 5.12 3.46 ;
  LAYER M1 ;
        RECT 5.152 0.972 5.184 3.48 ;
  LAYER M3 ;
        RECT 5.152 0.992 5.184 1.024 ;
  LAYER M1 ;
        RECT 5.216 0.972 5.248 3.48 ;
  LAYER M3 ;
        RECT 5.216 3.428 5.248 3.46 ;
  LAYER M1 ;
        RECT 5.28 0.972 5.312 3.48 ;
  LAYER M3 ;
        RECT 5.28 0.992 5.312 1.024 ;
  LAYER M1 ;
        RECT 5.344 0.972 5.376 3.48 ;
  LAYER M3 ;
        RECT 5.344 3.428 5.376 3.46 ;
  LAYER M1 ;
        RECT 5.408 0.972 5.44 3.48 ;
  LAYER M3 ;
        RECT 5.408 0.992 5.44 1.024 ;
  LAYER M1 ;
        RECT 5.472 0.972 5.504 3.48 ;
  LAYER M3 ;
        RECT 5.472 3.428 5.504 3.46 ;
  LAYER M1 ;
        RECT 5.536 0.972 5.568 3.48 ;
  LAYER M3 ;
        RECT 5.536 0.992 5.568 1.024 ;
  LAYER M1 ;
        RECT 5.6 0.972 5.632 3.48 ;
  LAYER M3 ;
        RECT 5.6 3.428 5.632 3.46 ;
  LAYER M1 ;
        RECT 5.664 0.972 5.696 3.48 ;
  LAYER M3 ;
        RECT 5.664 0.992 5.696 1.024 ;
  LAYER M1 ;
        RECT 5.728 0.972 5.76 3.48 ;
  LAYER M3 ;
        RECT 5.728 3.428 5.76 3.46 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 3.48 ;
  LAYER M3 ;
        RECT 5.792 0.992 5.824 1.024 ;
  LAYER M1 ;
        RECT 5.856 0.972 5.888 3.48 ;
  LAYER M3 ;
        RECT 5.856 3.428 5.888 3.46 ;
  LAYER M1 ;
        RECT 5.92 0.972 5.952 3.48 ;
  LAYER M3 ;
        RECT 5.92 0.992 5.952 1.024 ;
  LAYER M1 ;
        RECT 5.984 0.972 6.016 3.48 ;
  LAYER M3 ;
        RECT 5.984 3.428 6.016 3.46 ;
  LAYER M1 ;
        RECT 6.048 0.972 6.08 3.48 ;
  LAYER M3 ;
        RECT 6.048 0.992 6.08 1.024 ;
  LAYER M1 ;
        RECT 6.112 0.972 6.144 3.48 ;
  LAYER M3 ;
        RECT 6.112 3.428 6.144 3.46 ;
  LAYER M1 ;
        RECT 6.176 0.972 6.208 3.48 ;
  LAYER M3 ;
        RECT 6.176 0.992 6.208 1.024 ;
  LAYER M1 ;
        RECT 6.24 0.972 6.272 3.48 ;
  LAYER M3 ;
        RECT 6.24 3.428 6.272 3.46 ;
  LAYER M1 ;
        RECT 6.304 0.972 6.336 3.48 ;
  LAYER M3 ;
        RECT 6.304 0.992 6.336 1.024 ;
  LAYER M1 ;
        RECT 6.368 0.972 6.4 3.48 ;
  LAYER M3 ;
        RECT 6.368 3.428 6.4 3.46 ;
  LAYER M1 ;
        RECT 6.432 0.972 6.464 3.48 ;
  LAYER M3 ;
        RECT 4.064 1.056 4.096 1.088 ;
  LAYER M2 ;
        RECT 6.432 1.12 6.464 1.152 ;
  LAYER M2 ;
        RECT 4.064 1.184 4.096 1.216 ;
  LAYER M2 ;
        RECT 6.432 1.248 6.464 1.28 ;
  LAYER M2 ;
        RECT 4.064 1.312 4.096 1.344 ;
  LAYER M2 ;
        RECT 6.432 1.376 6.464 1.408 ;
  LAYER M2 ;
        RECT 4.064 1.44 4.096 1.472 ;
  LAYER M2 ;
        RECT 6.432 1.504 6.464 1.536 ;
  LAYER M2 ;
        RECT 4.064 1.568 4.096 1.6 ;
  LAYER M2 ;
        RECT 6.432 1.632 6.464 1.664 ;
  LAYER M2 ;
        RECT 4.064 1.696 4.096 1.728 ;
  LAYER M2 ;
        RECT 6.432 1.76 6.464 1.792 ;
  LAYER M2 ;
        RECT 4.064 1.824 4.096 1.856 ;
  LAYER M2 ;
        RECT 6.432 1.888 6.464 1.92 ;
  LAYER M2 ;
        RECT 4.064 1.952 4.096 1.984 ;
  LAYER M2 ;
        RECT 6.432 2.016 6.464 2.048 ;
  LAYER M2 ;
        RECT 4.064 2.08 4.096 2.112 ;
  LAYER M2 ;
        RECT 6.432 2.144 6.464 2.176 ;
  LAYER M2 ;
        RECT 4.064 2.208 4.096 2.24 ;
  LAYER M2 ;
        RECT 6.432 2.272 6.464 2.304 ;
  LAYER M2 ;
        RECT 4.064 2.336 4.096 2.368 ;
  LAYER M2 ;
        RECT 6.432 2.4 6.464 2.432 ;
  LAYER M2 ;
        RECT 4.064 2.464 4.096 2.496 ;
  LAYER M2 ;
        RECT 6.432 2.528 6.464 2.56 ;
  LAYER M2 ;
        RECT 4.064 2.592 4.096 2.624 ;
  LAYER M2 ;
        RECT 6.432 2.656 6.464 2.688 ;
  LAYER M2 ;
        RECT 4.064 2.72 4.096 2.752 ;
  LAYER M2 ;
        RECT 6.432 2.784 6.464 2.816 ;
  LAYER M2 ;
        RECT 4.064 2.848 4.096 2.88 ;
  LAYER M2 ;
        RECT 6.432 2.912 6.464 2.944 ;
  LAYER M2 ;
        RECT 4.064 2.976 4.096 3.008 ;
  LAYER M2 ;
        RECT 6.432 3.04 6.464 3.072 ;
  LAYER M2 ;
        RECT 4.064 3.104 4.096 3.136 ;
  LAYER M2 ;
        RECT 6.432 3.168 6.464 3.2 ;
  LAYER M2 ;
        RECT 4.064 3.232 4.096 3.264 ;
  LAYER M2 ;
        RECT 6.432 3.296 6.464 3.328 ;
  LAYER M2 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M1 ;
        RECT 4.064 4.08 4.096 6.588 ;
  LAYER M3 ;
        RECT 4.064 6.536 4.096 6.568 ;
  LAYER M1 ;
        RECT 4.128 4.08 4.16 6.588 ;
  LAYER M3 ;
        RECT 4.128 4.1 4.16 4.132 ;
  LAYER M1 ;
        RECT 4.192 4.08 4.224 6.588 ;
  LAYER M3 ;
        RECT 4.192 6.536 4.224 6.568 ;
  LAYER M1 ;
        RECT 4.256 4.08 4.288 6.588 ;
  LAYER M3 ;
        RECT 4.256 4.1 4.288 4.132 ;
  LAYER M1 ;
        RECT 4.32 4.08 4.352 6.588 ;
  LAYER M3 ;
        RECT 4.32 6.536 4.352 6.568 ;
  LAYER M1 ;
        RECT 4.384 4.08 4.416 6.588 ;
  LAYER M3 ;
        RECT 4.384 4.1 4.416 4.132 ;
  LAYER M1 ;
        RECT 4.448 4.08 4.48 6.588 ;
  LAYER M3 ;
        RECT 4.448 6.536 4.48 6.568 ;
  LAYER M1 ;
        RECT 4.512 4.08 4.544 6.588 ;
  LAYER M3 ;
        RECT 4.512 4.1 4.544 4.132 ;
  LAYER M1 ;
        RECT 4.576 4.08 4.608 6.588 ;
  LAYER M3 ;
        RECT 4.576 6.536 4.608 6.568 ;
  LAYER M1 ;
        RECT 4.64 4.08 4.672 6.588 ;
  LAYER M3 ;
        RECT 4.64 4.1 4.672 4.132 ;
  LAYER M1 ;
        RECT 4.704 4.08 4.736 6.588 ;
  LAYER M3 ;
        RECT 4.704 6.536 4.736 6.568 ;
  LAYER M1 ;
        RECT 4.768 4.08 4.8 6.588 ;
  LAYER M3 ;
        RECT 4.768 4.1 4.8 4.132 ;
  LAYER M1 ;
        RECT 4.832 4.08 4.864 6.588 ;
  LAYER M3 ;
        RECT 4.832 6.536 4.864 6.568 ;
  LAYER M1 ;
        RECT 4.896 4.08 4.928 6.588 ;
  LAYER M3 ;
        RECT 4.896 4.1 4.928 4.132 ;
  LAYER M1 ;
        RECT 4.96 4.08 4.992 6.588 ;
  LAYER M3 ;
        RECT 4.96 6.536 4.992 6.568 ;
  LAYER M1 ;
        RECT 5.024 4.08 5.056 6.588 ;
  LAYER M3 ;
        RECT 5.024 4.1 5.056 4.132 ;
  LAYER M1 ;
        RECT 5.088 4.08 5.12 6.588 ;
  LAYER M3 ;
        RECT 5.088 6.536 5.12 6.568 ;
  LAYER M1 ;
        RECT 5.152 4.08 5.184 6.588 ;
  LAYER M3 ;
        RECT 5.152 4.1 5.184 4.132 ;
  LAYER M1 ;
        RECT 5.216 4.08 5.248 6.588 ;
  LAYER M3 ;
        RECT 5.216 6.536 5.248 6.568 ;
  LAYER M1 ;
        RECT 5.28 4.08 5.312 6.588 ;
  LAYER M3 ;
        RECT 5.28 4.1 5.312 4.132 ;
  LAYER M1 ;
        RECT 5.344 4.08 5.376 6.588 ;
  LAYER M3 ;
        RECT 5.344 6.536 5.376 6.568 ;
  LAYER M1 ;
        RECT 5.408 4.08 5.44 6.588 ;
  LAYER M3 ;
        RECT 5.408 4.1 5.44 4.132 ;
  LAYER M1 ;
        RECT 5.472 4.08 5.504 6.588 ;
  LAYER M3 ;
        RECT 5.472 6.536 5.504 6.568 ;
  LAYER M1 ;
        RECT 5.536 4.08 5.568 6.588 ;
  LAYER M3 ;
        RECT 5.536 4.1 5.568 4.132 ;
  LAYER M1 ;
        RECT 5.6 4.08 5.632 6.588 ;
  LAYER M3 ;
        RECT 5.6 6.536 5.632 6.568 ;
  LAYER M1 ;
        RECT 5.664 4.08 5.696 6.588 ;
  LAYER M3 ;
        RECT 5.664 4.1 5.696 4.132 ;
  LAYER M1 ;
        RECT 5.728 4.08 5.76 6.588 ;
  LAYER M3 ;
        RECT 5.728 6.536 5.76 6.568 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 6.588 ;
  LAYER M3 ;
        RECT 5.792 4.1 5.824 4.132 ;
  LAYER M1 ;
        RECT 5.856 4.08 5.888 6.588 ;
  LAYER M3 ;
        RECT 5.856 6.536 5.888 6.568 ;
  LAYER M1 ;
        RECT 5.92 4.08 5.952 6.588 ;
  LAYER M3 ;
        RECT 5.92 4.1 5.952 4.132 ;
  LAYER M1 ;
        RECT 5.984 4.08 6.016 6.588 ;
  LAYER M3 ;
        RECT 5.984 6.536 6.016 6.568 ;
  LAYER M1 ;
        RECT 6.048 4.08 6.08 6.588 ;
  LAYER M3 ;
        RECT 6.048 4.1 6.08 4.132 ;
  LAYER M1 ;
        RECT 6.112 4.08 6.144 6.588 ;
  LAYER M3 ;
        RECT 6.112 6.536 6.144 6.568 ;
  LAYER M1 ;
        RECT 6.176 4.08 6.208 6.588 ;
  LAYER M3 ;
        RECT 6.176 4.1 6.208 4.132 ;
  LAYER M1 ;
        RECT 6.24 4.08 6.272 6.588 ;
  LAYER M3 ;
        RECT 6.24 6.536 6.272 6.568 ;
  LAYER M1 ;
        RECT 6.304 4.08 6.336 6.588 ;
  LAYER M3 ;
        RECT 6.304 4.1 6.336 4.132 ;
  LAYER M1 ;
        RECT 6.368 4.08 6.4 6.588 ;
  LAYER M3 ;
        RECT 6.368 6.536 6.4 6.568 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 6.588 ;
  LAYER M3 ;
        RECT 4.064 4.164 4.096 4.196 ;
  LAYER M2 ;
        RECT 6.432 4.228 6.464 4.26 ;
  LAYER M2 ;
        RECT 4.064 4.292 4.096 4.324 ;
  LAYER M2 ;
        RECT 6.432 4.356 6.464 4.388 ;
  LAYER M2 ;
        RECT 4.064 4.42 4.096 4.452 ;
  LAYER M2 ;
        RECT 6.432 4.484 6.464 4.516 ;
  LAYER M2 ;
        RECT 4.064 4.548 4.096 4.58 ;
  LAYER M2 ;
        RECT 6.432 4.612 6.464 4.644 ;
  LAYER M2 ;
        RECT 4.064 4.676 4.096 4.708 ;
  LAYER M2 ;
        RECT 6.432 4.74 6.464 4.772 ;
  LAYER M2 ;
        RECT 4.064 4.804 4.096 4.836 ;
  LAYER M2 ;
        RECT 6.432 4.868 6.464 4.9 ;
  LAYER M2 ;
        RECT 4.064 4.932 4.096 4.964 ;
  LAYER M2 ;
        RECT 6.432 4.996 6.464 5.028 ;
  LAYER M2 ;
        RECT 4.064 5.06 4.096 5.092 ;
  LAYER M2 ;
        RECT 6.432 5.124 6.464 5.156 ;
  LAYER M2 ;
        RECT 4.064 5.188 4.096 5.22 ;
  LAYER M2 ;
        RECT 6.432 5.252 6.464 5.284 ;
  LAYER M2 ;
        RECT 4.064 5.316 4.096 5.348 ;
  LAYER M2 ;
        RECT 6.432 5.38 6.464 5.412 ;
  LAYER M2 ;
        RECT 4.064 5.444 4.096 5.476 ;
  LAYER M2 ;
        RECT 6.432 5.508 6.464 5.54 ;
  LAYER M2 ;
        RECT 4.064 5.572 4.096 5.604 ;
  LAYER M2 ;
        RECT 6.432 5.636 6.464 5.668 ;
  LAYER M2 ;
        RECT 4.064 5.7 4.096 5.732 ;
  LAYER M2 ;
        RECT 6.432 5.764 6.464 5.796 ;
  LAYER M2 ;
        RECT 4.064 5.828 4.096 5.86 ;
  LAYER M2 ;
        RECT 6.432 5.892 6.464 5.924 ;
  LAYER M2 ;
        RECT 4.064 5.956 4.096 5.988 ;
  LAYER M2 ;
        RECT 6.432 6.02 6.464 6.052 ;
  LAYER M2 ;
        RECT 4.064 6.084 4.096 6.116 ;
  LAYER M2 ;
        RECT 6.432 6.148 6.464 6.18 ;
  LAYER M2 ;
        RECT 4.064 6.212 4.096 6.244 ;
  LAYER M2 ;
        RECT 6.432 6.276 6.464 6.308 ;
  LAYER M2 ;
        RECT 4.064 6.34 4.096 6.372 ;
  LAYER M2 ;
        RECT 6.432 6.404 6.464 6.436 ;
  LAYER M2 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M1 ;
        RECT 4.064 7.188 4.096 9.696 ;
  LAYER M3 ;
        RECT 4.064 9.644 4.096 9.676 ;
  LAYER M1 ;
        RECT 4.128 7.188 4.16 9.696 ;
  LAYER M3 ;
        RECT 4.128 7.208 4.16 7.24 ;
  LAYER M1 ;
        RECT 4.192 7.188 4.224 9.696 ;
  LAYER M3 ;
        RECT 4.192 9.644 4.224 9.676 ;
  LAYER M1 ;
        RECT 4.256 7.188 4.288 9.696 ;
  LAYER M3 ;
        RECT 4.256 7.208 4.288 7.24 ;
  LAYER M1 ;
        RECT 4.32 7.188 4.352 9.696 ;
  LAYER M3 ;
        RECT 4.32 9.644 4.352 9.676 ;
  LAYER M1 ;
        RECT 4.384 7.188 4.416 9.696 ;
  LAYER M3 ;
        RECT 4.384 7.208 4.416 7.24 ;
  LAYER M1 ;
        RECT 4.448 7.188 4.48 9.696 ;
  LAYER M3 ;
        RECT 4.448 9.644 4.48 9.676 ;
  LAYER M1 ;
        RECT 4.512 7.188 4.544 9.696 ;
  LAYER M3 ;
        RECT 4.512 7.208 4.544 7.24 ;
  LAYER M1 ;
        RECT 4.576 7.188 4.608 9.696 ;
  LAYER M3 ;
        RECT 4.576 9.644 4.608 9.676 ;
  LAYER M1 ;
        RECT 4.64 7.188 4.672 9.696 ;
  LAYER M3 ;
        RECT 4.64 7.208 4.672 7.24 ;
  LAYER M1 ;
        RECT 4.704 7.188 4.736 9.696 ;
  LAYER M3 ;
        RECT 4.704 9.644 4.736 9.676 ;
  LAYER M1 ;
        RECT 4.768 7.188 4.8 9.696 ;
  LAYER M3 ;
        RECT 4.768 7.208 4.8 7.24 ;
  LAYER M1 ;
        RECT 4.832 7.188 4.864 9.696 ;
  LAYER M3 ;
        RECT 4.832 9.644 4.864 9.676 ;
  LAYER M1 ;
        RECT 4.896 7.188 4.928 9.696 ;
  LAYER M3 ;
        RECT 4.896 7.208 4.928 7.24 ;
  LAYER M1 ;
        RECT 4.96 7.188 4.992 9.696 ;
  LAYER M3 ;
        RECT 4.96 9.644 4.992 9.676 ;
  LAYER M1 ;
        RECT 5.024 7.188 5.056 9.696 ;
  LAYER M3 ;
        RECT 5.024 7.208 5.056 7.24 ;
  LAYER M1 ;
        RECT 5.088 7.188 5.12 9.696 ;
  LAYER M3 ;
        RECT 5.088 9.644 5.12 9.676 ;
  LAYER M1 ;
        RECT 5.152 7.188 5.184 9.696 ;
  LAYER M3 ;
        RECT 5.152 7.208 5.184 7.24 ;
  LAYER M1 ;
        RECT 5.216 7.188 5.248 9.696 ;
  LAYER M3 ;
        RECT 5.216 9.644 5.248 9.676 ;
  LAYER M1 ;
        RECT 5.28 7.188 5.312 9.696 ;
  LAYER M3 ;
        RECT 5.28 7.208 5.312 7.24 ;
  LAYER M1 ;
        RECT 5.344 7.188 5.376 9.696 ;
  LAYER M3 ;
        RECT 5.344 9.644 5.376 9.676 ;
  LAYER M1 ;
        RECT 5.408 7.188 5.44 9.696 ;
  LAYER M3 ;
        RECT 5.408 7.208 5.44 7.24 ;
  LAYER M1 ;
        RECT 5.472 7.188 5.504 9.696 ;
  LAYER M3 ;
        RECT 5.472 9.644 5.504 9.676 ;
  LAYER M1 ;
        RECT 5.536 7.188 5.568 9.696 ;
  LAYER M3 ;
        RECT 5.536 7.208 5.568 7.24 ;
  LAYER M1 ;
        RECT 5.6 7.188 5.632 9.696 ;
  LAYER M3 ;
        RECT 5.6 9.644 5.632 9.676 ;
  LAYER M1 ;
        RECT 5.664 7.188 5.696 9.696 ;
  LAYER M3 ;
        RECT 5.664 7.208 5.696 7.24 ;
  LAYER M1 ;
        RECT 5.728 7.188 5.76 9.696 ;
  LAYER M3 ;
        RECT 5.728 9.644 5.76 9.676 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 9.696 ;
  LAYER M3 ;
        RECT 5.792 7.208 5.824 7.24 ;
  LAYER M1 ;
        RECT 5.856 7.188 5.888 9.696 ;
  LAYER M3 ;
        RECT 5.856 9.644 5.888 9.676 ;
  LAYER M1 ;
        RECT 5.92 7.188 5.952 9.696 ;
  LAYER M3 ;
        RECT 5.92 7.208 5.952 7.24 ;
  LAYER M1 ;
        RECT 5.984 7.188 6.016 9.696 ;
  LAYER M3 ;
        RECT 5.984 9.644 6.016 9.676 ;
  LAYER M1 ;
        RECT 6.048 7.188 6.08 9.696 ;
  LAYER M3 ;
        RECT 6.048 7.208 6.08 7.24 ;
  LAYER M1 ;
        RECT 6.112 7.188 6.144 9.696 ;
  LAYER M3 ;
        RECT 6.112 9.644 6.144 9.676 ;
  LAYER M1 ;
        RECT 6.176 7.188 6.208 9.696 ;
  LAYER M3 ;
        RECT 6.176 7.208 6.208 7.24 ;
  LAYER M1 ;
        RECT 6.24 7.188 6.272 9.696 ;
  LAYER M3 ;
        RECT 6.24 9.644 6.272 9.676 ;
  LAYER M1 ;
        RECT 6.304 7.188 6.336 9.696 ;
  LAYER M3 ;
        RECT 6.304 7.208 6.336 7.24 ;
  LAYER M1 ;
        RECT 6.368 7.188 6.4 9.696 ;
  LAYER M3 ;
        RECT 6.368 9.644 6.4 9.676 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 9.696 ;
  LAYER M3 ;
        RECT 4.064 7.272 4.096 7.304 ;
  LAYER M2 ;
        RECT 6.432 7.336 6.464 7.368 ;
  LAYER M2 ;
        RECT 4.064 7.4 4.096 7.432 ;
  LAYER M2 ;
        RECT 6.432 7.464 6.464 7.496 ;
  LAYER M2 ;
        RECT 4.064 7.528 4.096 7.56 ;
  LAYER M2 ;
        RECT 6.432 7.592 6.464 7.624 ;
  LAYER M2 ;
        RECT 4.064 7.656 4.096 7.688 ;
  LAYER M2 ;
        RECT 6.432 7.72 6.464 7.752 ;
  LAYER M2 ;
        RECT 4.064 7.784 4.096 7.816 ;
  LAYER M2 ;
        RECT 6.432 7.848 6.464 7.88 ;
  LAYER M2 ;
        RECT 4.064 7.912 4.096 7.944 ;
  LAYER M2 ;
        RECT 6.432 7.976 6.464 8.008 ;
  LAYER M2 ;
        RECT 4.064 8.04 4.096 8.072 ;
  LAYER M2 ;
        RECT 6.432 8.104 6.464 8.136 ;
  LAYER M2 ;
        RECT 4.064 8.168 4.096 8.2 ;
  LAYER M2 ;
        RECT 6.432 8.232 6.464 8.264 ;
  LAYER M2 ;
        RECT 4.064 8.296 4.096 8.328 ;
  LAYER M2 ;
        RECT 6.432 8.36 6.464 8.392 ;
  LAYER M2 ;
        RECT 4.064 8.424 4.096 8.456 ;
  LAYER M2 ;
        RECT 6.432 8.488 6.464 8.52 ;
  LAYER M2 ;
        RECT 4.064 8.552 4.096 8.584 ;
  LAYER M2 ;
        RECT 6.432 8.616 6.464 8.648 ;
  LAYER M2 ;
        RECT 4.064 8.68 4.096 8.712 ;
  LAYER M2 ;
        RECT 6.432 8.744 6.464 8.776 ;
  LAYER M2 ;
        RECT 4.064 8.808 4.096 8.84 ;
  LAYER M2 ;
        RECT 6.432 8.872 6.464 8.904 ;
  LAYER M2 ;
        RECT 4.064 8.936 4.096 8.968 ;
  LAYER M2 ;
        RECT 6.432 9 6.464 9.032 ;
  LAYER M2 ;
        RECT 4.064 9.064 4.096 9.096 ;
  LAYER M2 ;
        RECT 6.432 9.128 6.464 9.16 ;
  LAYER M2 ;
        RECT 4.064 9.192 4.096 9.224 ;
  LAYER M2 ;
        RECT 6.432 9.256 6.464 9.288 ;
  LAYER M2 ;
        RECT 4.064 9.32 4.096 9.352 ;
  LAYER M2 ;
        RECT 6.432 9.384 6.464 9.416 ;
  LAYER M2 ;
        RECT 4.064 9.448 4.096 9.48 ;
  LAYER M2 ;
        RECT 6.432 9.512 6.464 9.544 ;
  LAYER M2 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M1 ;
        RECT 4.064 10.296 4.096 12.804 ;
  LAYER M3 ;
        RECT 4.064 12.752 4.096 12.784 ;
  LAYER M1 ;
        RECT 4.128 10.296 4.16 12.804 ;
  LAYER M3 ;
        RECT 4.128 10.316 4.16 10.348 ;
  LAYER M1 ;
        RECT 4.192 10.296 4.224 12.804 ;
  LAYER M3 ;
        RECT 4.192 12.752 4.224 12.784 ;
  LAYER M1 ;
        RECT 4.256 10.296 4.288 12.804 ;
  LAYER M3 ;
        RECT 4.256 10.316 4.288 10.348 ;
  LAYER M1 ;
        RECT 4.32 10.296 4.352 12.804 ;
  LAYER M3 ;
        RECT 4.32 12.752 4.352 12.784 ;
  LAYER M1 ;
        RECT 4.384 10.296 4.416 12.804 ;
  LAYER M3 ;
        RECT 4.384 10.316 4.416 10.348 ;
  LAYER M1 ;
        RECT 4.448 10.296 4.48 12.804 ;
  LAYER M3 ;
        RECT 4.448 12.752 4.48 12.784 ;
  LAYER M1 ;
        RECT 4.512 10.296 4.544 12.804 ;
  LAYER M3 ;
        RECT 4.512 10.316 4.544 10.348 ;
  LAYER M1 ;
        RECT 4.576 10.296 4.608 12.804 ;
  LAYER M3 ;
        RECT 4.576 12.752 4.608 12.784 ;
  LAYER M1 ;
        RECT 4.64 10.296 4.672 12.804 ;
  LAYER M3 ;
        RECT 4.64 10.316 4.672 10.348 ;
  LAYER M1 ;
        RECT 4.704 10.296 4.736 12.804 ;
  LAYER M3 ;
        RECT 4.704 12.752 4.736 12.784 ;
  LAYER M1 ;
        RECT 4.768 10.296 4.8 12.804 ;
  LAYER M3 ;
        RECT 4.768 10.316 4.8 10.348 ;
  LAYER M1 ;
        RECT 4.832 10.296 4.864 12.804 ;
  LAYER M3 ;
        RECT 4.832 12.752 4.864 12.784 ;
  LAYER M1 ;
        RECT 4.896 10.296 4.928 12.804 ;
  LAYER M3 ;
        RECT 4.896 10.316 4.928 10.348 ;
  LAYER M1 ;
        RECT 4.96 10.296 4.992 12.804 ;
  LAYER M3 ;
        RECT 4.96 12.752 4.992 12.784 ;
  LAYER M1 ;
        RECT 5.024 10.296 5.056 12.804 ;
  LAYER M3 ;
        RECT 5.024 10.316 5.056 10.348 ;
  LAYER M1 ;
        RECT 5.088 10.296 5.12 12.804 ;
  LAYER M3 ;
        RECT 5.088 12.752 5.12 12.784 ;
  LAYER M1 ;
        RECT 5.152 10.296 5.184 12.804 ;
  LAYER M3 ;
        RECT 5.152 10.316 5.184 10.348 ;
  LAYER M1 ;
        RECT 5.216 10.296 5.248 12.804 ;
  LAYER M3 ;
        RECT 5.216 12.752 5.248 12.784 ;
  LAYER M1 ;
        RECT 5.28 10.296 5.312 12.804 ;
  LAYER M3 ;
        RECT 5.28 10.316 5.312 10.348 ;
  LAYER M1 ;
        RECT 5.344 10.296 5.376 12.804 ;
  LAYER M3 ;
        RECT 5.344 12.752 5.376 12.784 ;
  LAYER M1 ;
        RECT 5.408 10.296 5.44 12.804 ;
  LAYER M3 ;
        RECT 5.408 10.316 5.44 10.348 ;
  LAYER M1 ;
        RECT 5.472 10.296 5.504 12.804 ;
  LAYER M3 ;
        RECT 5.472 12.752 5.504 12.784 ;
  LAYER M1 ;
        RECT 5.536 10.296 5.568 12.804 ;
  LAYER M3 ;
        RECT 5.536 10.316 5.568 10.348 ;
  LAYER M1 ;
        RECT 5.6 10.296 5.632 12.804 ;
  LAYER M3 ;
        RECT 5.6 12.752 5.632 12.784 ;
  LAYER M1 ;
        RECT 5.664 10.296 5.696 12.804 ;
  LAYER M3 ;
        RECT 5.664 10.316 5.696 10.348 ;
  LAYER M1 ;
        RECT 5.728 10.296 5.76 12.804 ;
  LAYER M3 ;
        RECT 5.728 12.752 5.76 12.784 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 12.804 ;
  LAYER M3 ;
        RECT 5.792 10.316 5.824 10.348 ;
  LAYER M1 ;
        RECT 5.856 10.296 5.888 12.804 ;
  LAYER M3 ;
        RECT 5.856 12.752 5.888 12.784 ;
  LAYER M1 ;
        RECT 5.92 10.296 5.952 12.804 ;
  LAYER M3 ;
        RECT 5.92 10.316 5.952 10.348 ;
  LAYER M1 ;
        RECT 5.984 10.296 6.016 12.804 ;
  LAYER M3 ;
        RECT 5.984 12.752 6.016 12.784 ;
  LAYER M1 ;
        RECT 6.048 10.296 6.08 12.804 ;
  LAYER M3 ;
        RECT 6.048 10.316 6.08 10.348 ;
  LAYER M1 ;
        RECT 6.112 10.296 6.144 12.804 ;
  LAYER M3 ;
        RECT 6.112 12.752 6.144 12.784 ;
  LAYER M1 ;
        RECT 6.176 10.296 6.208 12.804 ;
  LAYER M3 ;
        RECT 6.176 10.316 6.208 10.348 ;
  LAYER M1 ;
        RECT 6.24 10.296 6.272 12.804 ;
  LAYER M3 ;
        RECT 6.24 12.752 6.272 12.784 ;
  LAYER M1 ;
        RECT 6.304 10.296 6.336 12.804 ;
  LAYER M3 ;
        RECT 6.304 10.316 6.336 10.348 ;
  LAYER M1 ;
        RECT 6.368 10.296 6.4 12.804 ;
  LAYER M3 ;
        RECT 6.368 12.752 6.4 12.784 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 12.804 ;
  LAYER M3 ;
        RECT 4.064 10.38 4.096 10.412 ;
  LAYER M2 ;
        RECT 6.432 10.444 6.464 10.476 ;
  LAYER M2 ;
        RECT 4.064 10.508 4.096 10.54 ;
  LAYER M2 ;
        RECT 6.432 10.572 6.464 10.604 ;
  LAYER M2 ;
        RECT 4.064 10.636 4.096 10.668 ;
  LAYER M2 ;
        RECT 6.432 10.7 6.464 10.732 ;
  LAYER M2 ;
        RECT 4.064 10.764 4.096 10.796 ;
  LAYER M2 ;
        RECT 6.432 10.828 6.464 10.86 ;
  LAYER M2 ;
        RECT 4.064 10.892 4.096 10.924 ;
  LAYER M2 ;
        RECT 6.432 10.956 6.464 10.988 ;
  LAYER M2 ;
        RECT 4.064 11.02 4.096 11.052 ;
  LAYER M2 ;
        RECT 6.432 11.084 6.464 11.116 ;
  LAYER M2 ;
        RECT 4.064 11.148 4.096 11.18 ;
  LAYER M2 ;
        RECT 6.432 11.212 6.464 11.244 ;
  LAYER M2 ;
        RECT 4.064 11.276 4.096 11.308 ;
  LAYER M2 ;
        RECT 6.432 11.34 6.464 11.372 ;
  LAYER M2 ;
        RECT 4.064 11.404 4.096 11.436 ;
  LAYER M2 ;
        RECT 6.432 11.468 6.464 11.5 ;
  LAYER M2 ;
        RECT 4.064 11.532 4.096 11.564 ;
  LAYER M2 ;
        RECT 6.432 11.596 6.464 11.628 ;
  LAYER M2 ;
        RECT 4.064 11.66 4.096 11.692 ;
  LAYER M2 ;
        RECT 6.432 11.724 6.464 11.756 ;
  LAYER M2 ;
        RECT 4.064 11.788 4.096 11.82 ;
  LAYER M2 ;
        RECT 6.432 11.852 6.464 11.884 ;
  LAYER M2 ;
        RECT 4.064 11.916 4.096 11.948 ;
  LAYER M2 ;
        RECT 6.432 11.98 6.464 12.012 ;
  LAYER M2 ;
        RECT 4.064 12.044 4.096 12.076 ;
  LAYER M2 ;
        RECT 6.432 12.108 6.464 12.14 ;
  LAYER M2 ;
        RECT 4.064 12.172 4.096 12.204 ;
  LAYER M2 ;
        RECT 6.432 12.236 6.464 12.268 ;
  LAYER M2 ;
        RECT 4.064 12.3 4.096 12.332 ;
  LAYER M2 ;
        RECT 6.432 12.364 6.464 12.396 ;
  LAYER M2 ;
        RECT 4.064 12.428 4.096 12.46 ;
  LAYER M2 ;
        RECT 6.432 12.492 6.464 12.524 ;
  LAYER M2 ;
        RECT 4.064 12.556 4.096 12.588 ;
  LAYER M2 ;
        RECT 6.432 12.62 6.464 12.652 ;
  LAYER M2 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M1 ;
        RECT 4.064 13.404 4.096 15.912 ;
  LAYER M3 ;
        RECT 4.064 15.86 4.096 15.892 ;
  LAYER M1 ;
        RECT 4.128 13.404 4.16 15.912 ;
  LAYER M3 ;
        RECT 4.128 13.424 4.16 13.456 ;
  LAYER M1 ;
        RECT 4.192 13.404 4.224 15.912 ;
  LAYER M3 ;
        RECT 4.192 15.86 4.224 15.892 ;
  LAYER M1 ;
        RECT 4.256 13.404 4.288 15.912 ;
  LAYER M3 ;
        RECT 4.256 13.424 4.288 13.456 ;
  LAYER M1 ;
        RECT 4.32 13.404 4.352 15.912 ;
  LAYER M3 ;
        RECT 4.32 15.86 4.352 15.892 ;
  LAYER M1 ;
        RECT 4.384 13.404 4.416 15.912 ;
  LAYER M3 ;
        RECT 4.384 13.424 4.416 13.456 ;
  LAYER M1 ;
        RECT 4.448 13.404 4.48 15.912 ;
  LAYER M3 ;
        RECT 4.448 15.86 4.48 15.892 ;
  LAYER M1 ;
        RECT 4.512 13.404 4.544 15.912 ;
  LAYER M3 ;
        RECT 4.512 13.424 4.544 13.456 ;
  LAYER M1 ;
        RECT 4.576 13.404 4.608 15.912 ;
  LAYER M3 ;
        RECT 4.576 15.86 4.608 15.892 ;
  LAYER M1 ;
        RECT 4.64 13.404 4.672 15.912 ;
  LAYER M3 ;
        RECT 4.64 13.424 4.672 13.456 ;
  LAYER M1 ;
        RECT 4.704 13.404 4.736 15.912 ;
  LAYER M3 ;
        RECT 4.704 15.86 4.736 15.892 ;
  LAYER M1 ;
        RECT 4.768 13.404 4.8 15.912 ;
  LAYER M3 ;
        RECT 4.768 13.424 4.8 13.456 ;
  LAYER M1 ;
        RECT 4.832 13.404 4.864 15.912 ;
  LAYER M3 ;
        RECT 4.832 15.86 4.864 15.892 ;
  LAYER M1 ;
        RECT 4.896 13.404 4.928 15.912 ;
  LAYER M3 ;
        RECT 4.896 13.424 4.928 13.456 ;
  LAYER M1 ;
        RECT 4.96 13.404 4.992 15.912 ;
  LAYER M3 ;
        RECT 4.96 15.86 4.992 15.892 ;
  LAYER M1 ;
        RECT 5.024 13.404 5.056 15.912 ;
  LAYER M3 ;
        RECT 5.024 13.424 5.056 13.456 ;
  LAYER M1 ;
        RECT 5.088 13.404 5.12 15.912 ;
  LAYER M3 ;
        RECT 5.088 15.86 5.12 15.892 ;
  LAYER M1 ;
        RECT 5.152 13.404 5.184 15.912 ;
  LAYER M3 ;
        RECT 5.152 13.424 5.184 13.456 ;
  LAYER M1 ;
        RECT 5.216 13.404 5.248 15.912 ;
  LAYER M3 ;
        RECT 5.216 15.86 5.248 15.892 ;
  LAYER M1 ;
        RECT 5.28 13.404 5.312 15.912 ;
  LAYER M3 ;
        RECT 5.28 13.424 5.312 13.456 ;
  LAYER M1 ;
        RECT 5.344 13.404 5.376 15.912 ;
  LAYER M3 ;
        RECT 5.344 15.86 5.376 15.892 ;
  LAYER M1 ;
        RECT 5.408 13.404 5.44 15.912 ;
  LAYER M3 ;
        RECT 5.408 13.424 5.44 13.456 ;
  LAYER M1 ;
        RECT 5.472 13.404 5.504 15.912 ;
  LAYER M3 ;
        RECT 5.472 15.86 5.504 15.892 ;
  LAYER M1 ;
        RECT 5.536 13.404 5.568 15.912 ;
  LAYER M3 ;
        RECT 5.536 13.424 5.568 13.456 ;
  LAYER M1 ;
        RECT 5.6 13.404 5.632 15.912 ;
  LAYER M3 ;
        RECT 5.6 15.86 5.632 15.892 ;
  LAYER M1 ;
        RECT 5.664 13.404 5.696 15.912 ;
  LAYER M3 ;
        RECT 5.664 13.424 5.696 13.456 ;
  LAYER M1 ;
        RECT 5.728 13.404 5.76 15.912 ;
  LAYER M3 ;
        RECT 5.728 15.86 5.76 15.892 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 15.912 ;
  LAYER M3 ;
        RECT 5.792 13.424 5.824 13.456 ;
  LAYER M1 ;
        RECT 5.856 13.404 5.888 15.912 ;
  LAYER M3 ;
        RECT 5.856 15.86 5.888 15.892 ;
  LAYER M1 ;
        RECT 5.92 13.404 5.952 15.912 ;
  LAYER M3 ;
        RECT 5.92 13.424 5.952 13.456 ;
  LAYER M1 ;
        RECT 5.984 13.404 6.016 15.912 ;
  LAYER M3 ;
        RECT 5.984 15.86 6.016 15.892 ;
  LAYER M1 ;
        RECT 6.048 13.404 6.08 15.912 ;
  LAYER M3 ;
        RECT 6.048 13.424 6.08 13.456 ;
  LAYER M1 ;
        RECT 6.112 13.404 6.144 15.912 ;
  LAYER M3 ;
        RECT 6.112 15.86 6.144 15.892 ;
  LAYER M1 ;
        RECT 6.176 13.404 6.208 15.912 ;
  LAYER M3 ;
        RECT 6.176 13.424 6.208 13.456 ;
  LAYER M1 ;
        RECT 6.24 13.404 6.272 15.912 ;
  LAYER M3 ;
        RECT 6.24 15.86 6.272 15.892 ;
  LAYER M1 ;
        RECT 6.304 13.404 6.336 15.912 ;
  LAYER M3 ;
        RECT 6.304 13.424 6.336 13.456 ;
  LAYER M1 ;
        RECT 6.368 13.404 6.4 15.912 ;
  LAYER M3 ;
        RECT 6.368 15.86 6.4 15.892 ;
  LAYER M1 ;
        RECT 6.432 13.404 6.464 15.912 ;
  LAYER M3 ;
        RECT 4.064 13.488 4.096 13.52 ;
  LAYER M2 ;
        RECT 6.432 13.552 6.464 13.584 ;
  LAYER M2 ;
        RECT 4.064 13.616 4.096 13.648 ;
  LAYER M2 ;
        RECT 6.432 13.68 6.464 13.712 ;
  LAYER M2 ;
        RECT 4.064 13.744 4.096 13.776 ;
  LAYER M2 ;
        RECT 6.432 13.808 6.464 13.84 ;
  LAYER M2 ;
        RECT 4.064 13.872 4.096 13.904 ;
  LAYER M2 ;
        RECT 6.432 13.936 6.464 13.968 ;
  LAYER M2 ;
        RECT 4.064 14 4.096 14.032 ;
  LAYER M2 ;
        RECT 6.432 14.064 6.464 14.096 ;
  LAYER M2 ;
        RECT 4.064 14.128 4.096 14.16 ;
  LAYER M2 ;
        RECT 6.432 14.192 6.464 14.224 ;
  LAYER M2 ;
        RECT 4.064 14.256 4.096 14.288 ;
  LAYER M2 ;
        RECT 6.432 14.32 6.464 14.352 ;
  LAYER M2 ;
        RECT 4.064 14.384 4.096 14.416 ;
  LAYER M2 ;
        RECT 6.432 14.448 6.464 14.48 ;
  LAYER M2 ;
        RECT 4.064 14.512 4.096 14.544 ;
  LAYER M2 ;
        RECT 6.432 14.576 6.464 14.608 ;
  LAYER M2 ;
        RECT 4.064 14.64 4.096 14.672 ;
  LAYER M2 ;
        RECT 6.432 14.704 6.464 14.736 ;
  LAYER M2 ;
        RECT 4.064 14.768 4.096 14.8 ;
  LAYER M2 ;
        RECT 6.432 14.832 6.464 14.864 ;
  LAYER M2 ;
        RECT 4.064 14.896 4.096 14.928 ;
  LAYER M2 ;
        RECT 6.432 14.96 6.464 14.992 ;
  LAYER M2 ;
        RECT 4.064 15.024 4.096 15.056 ;
  LAYER M2 ;
        RECT 6.432 15.088 6.464 15.12 ;
  LAYER M2 ;
        RECT 4.064 15.152 4.096 15.184 ;
  LAYER M2 ;
        RECT 6.432 15.216 6.464 15.248 ;
  LAYER M2 ;
        RECT 4.064 15.28 4.096 15.312 ;
  LAYER M2 ;
        RECT 6.432 15.344 6.464 15.376 ;
  LAYER M2 ;
        RECT 4.064 15.408 4.096 15.44 ;
  LAYER M2 ;
        RECT 6.432 15.472 6.464 15.504 ;
  LAYER M2 ;
        RECT 4.064 15.536 4.096 15.568 ;
  LAYER M2 ;
        RECT 6.432 15.6 6.464 15.632 ;
  LAYER M2 ;
        RECT 4.064 15.664 4.096 15.696 ;
  LAYER M2 ;
        RECT 6.432 15.728 6.464 15.76 ;
  LAYER M2 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M1 ;
        RECT 4.064 16.512 4.096 19.02 ;
  LAYER M3 ;
        RECT 4.064 18.968 4.096 19 ;
  LAYER M1 ;
        RECT 4.128 16.512 4.16 19.02 ;
  LAYER M3 ;
        RECT 4.128 16.532 4.16 16.564 ;
  LAYER M1 ;
        RECT 4.192 16.512 4.224 19.02 ;
  LAYER M3 ;
        RECT 4.192 18.968 4.224 19 ;
  LAYER M1 ;
        RECT 4.256 16.512 4.288 19.02 ;
  LAYER M3 ;
        RECT 4.256 16.532 4.288 16.564 ;
  LAYER M1 ;
        RECT 4.32 16.512 4.352 19.02 ;
  LAYER M3 ;
        RECT 4.32 18.968 4.352 19 ;
  LAYER M1 ;
        RECT 4.384 16.512 4.416 19.02 ;
  LAYER M3 ;
        RECT 4.384 16.532 4.416 16.564 ;
  LAYER M1 ;
        RECT 4.448 16.512 4.48 19.02 ;
  LAYER M3 ;
        RECT 4.448 18.968 4.48 19 ;
  LAYER M1 ;
        RECT 4.512 16.512 4.544 19.02 ;
  LAYER M3 ;
        RECT 4.512 16.532 4.544 16.564 ;
  LAYER M1 ;
        RECT 4.576 16.512 4.608 19.02 ;
  LAYER M3 ;
        RECT 4.576 18.968 4.608 19 ;
  LAYER M1 ;
        RECT 4.64 16.512 4.672 19.02 ;
  LAYER M3 ;
        RECT 4.64 16.532 4.672 16.564 ;
  LAYER M1 ;
        RECT 4.704 16.512 4.736 19.02 ;
  LAYER M3 ;
        RECT 4.704 18.968 4.736 19 ;
  LAYER M1 ;
        RECT 4.768 16.512 4.8 19.02 ;
  LAYER M3 ;
        RECT 4.768 16.532 4.8 16.564 ;
  LAYER M1 ;
        RECT 4.832 16.512 4.864 19.02 ;
  LAYER M3 ;
        RECT 4.832 18.968 4.864 19 ;
  LAYER M1 ;
        RECT 4.896 16.512 4.928 19.02 ;
  LAYER M3 ;
        RECT 4.896 16.532 4.928 16.564 ;
  LAYER M1 ;
        RECT 4.96 16.512 4.992 19.02 ;
  LAYER M3 ;
        RECT 4.96 18.968 4.992 19 ;
  LAYER M1 ;
        RECT 5.024 16.512 5.056 19.02 ;
  LAYER M3 ;
        RECT 5.024 16.532 5.056 16.564 ;
  LAYER M1 ;
        RECT 5.088 16.512 5.12 19.02 ;
  LAYER M3 ;
        RECT 5.088 18.968 5.12 19 ;
  LAYER M1 ;
        RECT 5.152 16.512 5.184 19.02 ;
  LAYER M3 ;
        RECT 5.152 16.532 5.184 16.564 ;
  LAYER M1 ;
        RECT 5.216 16.512 5.248 19.02 ;
  LAYER M3 ;
        RECT 5.216 18.968 5.248 19 ;
  LAYER M1 ;
        RECT 5.28 16.512 5.312 19.02 ;
  LAYER M3 ;
        RECT 5.28 16.532 5.312 16.564 ;
  LAYER M1 ;
        RECT 5.344 16.512 5.376 19.02 ;
  LAYER M3 ;
        RECT 5.344 18.968 5.376 19 ;
  LAYER M1 ;
        RECT 5.408 16.512 5.44 19.02 ;
  LAYER M3 ;
        RECT 5.408 16.532 5.44 16.564 ;
  LAYER M1 ;
        RECT 5.472 16.512 5.504 19.02 ;
  LAYER M3 ;
        RECT 5.472 18.968 5.504 19 ;
  LAYER M1 ;
        RECT 5.536 16.512 5.568 19.02 ;
  LAYER M3 ;
        RECT 5.536 16.532 5.568 16.564 ;
  LAYER M1 ;
        RECT 5.6 16.512 5.632 19.02 ;
  LAYER M3 ;
        RECT 5.6 18.968 5.632 19 ;
  LAYER M1 ;
        RECT 5.664 16.512 5.696 19.02 ;
  LAYER M3 ;
        RECT 5.664 16.532 5.696 16.564 ;
  LAYER M1 ;
        RECT 5.728 16.512 5.76 19.02 ;
  LAYER M3 ;
        RECT 5.728 18.968 5.76 19 ;
  LAYER M1 ;
        RECT 5.792 16.512 5.824 19.02 ;
  LAYER M3 ;
        RECT 5.792 16.532 5.824 16.564 ;
  LAYER M1 ;
        RECT 5.856 16.512 5.888 19.02 ;
  LAYER M3 ;
        RECT 5.856 18.968 5.888 19 ;
  LAYER M1 ;
        RECT 5.92 16.512 5.952 19.02 ;
  LAYER M3 ;
        RECT 5.92 16.532 5.952 16.564 ;
  LAYER M1 ;
        RECT 5.984 16.512 6.016 19.02 ;
  LAYER M3 ;
        RECT 5.984 18.968 6.016 19 ;
  LAYER M1 ;
        RECT 6.048 16.512 6.08 19.02 ;
  LAYER M3 ;
        RECT 6.048 16.532 6.08 16.564 ;
  LAYER M1 ;
        RECT 6.112 16.512 6.144 19.02 ;
  LAYER M3 ;
        RECT 6.112 18.968 6.144 19 ;
  LAYER M1 ;
        RECT 6.176 16.512 6.208 19.02 ;
  LAYER M3 ;
        RECT 6.176 16.532 6.208 16.564 ;
  LAYER M1 ;
        RECT 6.24 16.512 6.272 19.02 ;
  LAYER M3 ;
        RECT 6.24 18.968 6.272 19 ;
  LAYER M1 ;
        RECT 6.304 16.512 6.336 19.02 ;
  LAYER M3 ;
        RECT 6.304 16.532 6.336 16.564 ;
  LAYER M1 ;
        RECT 6.368 16.512 6.4 19.02 ;
  LAYER M3 ;
        RECT 6.368 18.968 6.4 19 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 19.02 ;
  LAYER M3 ;
        RECT 4.064 16.596 4.096 16.628 ;
  LAYER M2 ;
        RECT 6.432 16.66 6.464 16.692 ;
  LAYER M2 ;
        RECT 4.064 16.724 4.096 16.756 ;
  LAYER M2 ;
        RECT 6.432 16.788 6.464 16.82 ;
  LAYER M2 ;
        RECT 4.064 16.852 4.096 16.884 ;
  LAYER M2 ;
        RECT 6.432 16.916 6.464 16.948 ;
  LAYER M2 ;
        RECT 4.064 16.98 4.096 17.012 ;
  LAYER M2 ;
        RECT 6.432 17.044 6.464 17.076 ;
  LAYER M2 ;
        RECT 4.064 17.108 4.096 17.14 ;
  LAYER M2 ;
        RECT 6.432 17.172 6.464 17.204 ;
  LAYER M2 ;
        RECT 4.064 17.236 4.096 17.268 ;
  LAYER M2 ;
        RECT 6.432 17.3 6.464 17.332 ;
  LAYER M2 ;
        RECT 4.064 17.364 4.096 17.396 ;
  LAYER M2 ;
        RECT 6.432 17.428 6.464 17.46 ;
  LAYER M2 ;
        RECT 4.064 17.492 4.096 17.524 ;
  LAYER M2 ;
        RECT 6.432 17.556 6.464 17.588 ;
  LAYER M2 ;
        RECT 4.064 17.62 4.096 17.652 ;
  LAYER M2 ;
        RECT 6.432 17.684 6.464 17.716 ;
  LAYER M2 ;
        RECT 4.064 17.748 4.096 17.78 ;
  LAYER M2 ;
        RECT 6.432 17.812 6.464 17.844 ;
  LAYER M2 ;
        RECT 4.064 17.876 4.096 17.908 ;
  LAYER M2 ;
        RECT 6.432 17.94 6.464 17.972 ;
  LAYER M2 ;
        RECT 4.064 18.004 4.096 18.036 ;
  LAYER M2 ;
        RECT 6.432 18.068 6.464 18.1 ;
  LAYER M2 ;
        RECT 4.064 18.132 4.096 18.164 ;
  LAYER M2 ;
        RECT 6.432 18.196 6.464 18.228 ;
  LAYER M2 ;
        RECT 4.064 18.26 4.096 18.292 ;
  LAYER M2 ;
        RECT 6.432 18.324 6.464 18.356 ;
  LAYER M2 ;
        RECT 4.064 18.388 4.096 18.42 ;
  LAYER M2 ;
        RECT 6.432 18.452 6.464 18.484 ;
  LAYER M2 ;
        RECT 4.064 18.516 4.096 18.548 ;
  LAYER M2 ;
        RECT 6.432 18.58 6.464 18.612 ;
  LAYER M2 ;
        RECT 4.064 18.644 4.096 18.676 ;
  LAYER M2 ;
        RECT 6.432 18.708 6.464 18.74 ;
  LAYER M2 ;
        RECT 4.064 18.772 4.096 18.804 ;
  LAYER M2 ;
        RECT 6.432 18.836 6.464 18.868 ;
  LAYER M2 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M1 ;
        RECT 4.064 19.62 4.096 22.128 ;
  LAYER M3 ;
        RECT 4.064 22.076 4.096 22.108 ;
  LAYER M1 ;
        RECT 4.128 19.62 4.16 22.128 ;
  LAYER M3 ;
        RECT 4.128 19.64 4.16 19.672 ;
  LAYER M1 ;
        RECT 4.192 19.62 4.224 22.128 ;
  LAYER M3 ;
        RECT 4.192 22.076 4.224 22.108 ;
  LAYER M1 ;
        RECT 4.256 19.62 4.288 22.128 ;
  LAYER M3 ;
        RECT 4.256 19.64 4.288 19.672 ;
  LAYER M1 ;
        RECT 4.32 19.62 4.352 22.128 ;
  LAYER M3 ;
        RECT 4.32 22.076 4.352 22.108 ;
  LAYER M1 ;
        RECT 4.384 19.62 4.416 22.128 ;
  LAYER M3 ;
        RECT 4.384 19.64 4.416 19.672 ;
  LAYER M1 ;
        RECT 4.448 19.62 4.48 22.128 ;
  LAYER M3 ;
        RECT 4.448 22.076 4.48 22.108 ;
  LAYER M1 ;
        RECT 4.512 19.62 4.544 22.128 ;
  LAYER M3 ;
        RECT 4.512 19.64 4.544 19.672 ;
  LAYER M1 ;
        RECT 4.576 19.62 4.608 22.128 ;
  LAYER M3 ;
        RECT 4.576 22.076 4.608 22.108 ;
  LAYER M1 ;
        RECT 4.64 19.62 4.672 22.128 ;
  LAYER M3 ;
        RECT 4.64 19.64 4.672 19.672 ;
  LAYER M1 ;
        RECT 4.704 19.62 4.736 22.128 ;
  LAYER M3 ;
        RECT 4.704 22.076 4.736 22.108 ;
  LAYER M1 ;
        RECT 4.768 19.62 4.8 22.128 ;
  LAYER M3 ;
        RECT 4.768 19.64 4.8 19.672 ;
  LAYER M1 ;
        RECT 4.832 19.62 4.864 22.128 ;
  LAYER M3 ;
        RECT 4.832 22.076 4.864 22.108 ;
  LAYER M1 ;
        RECT 4.896 19.62 4.928 22.128 ;
  LAYER M3 ;
        RECT 4.896 19.64 4.928 19.672 ;
  LAYER M1 ;
        RECT 4.96 19.62 4.992 22.128 ;
  LAYER M3 ;
        RECT 4.96 22.076 4.992 22.108 ;
  LAYER M1 ;
        RECT 5.024 19.62 5.056 22.128 ;
  LAYER M3 ;
        RECT 5.024 19.64 5.056 19.672 ;
  LAYER M1 ;
        RECT 5.088 19.62 5.12 22.128 ;
  LAYER M3 ;
        RECT 5.088 22.076 5.12 22.108 ;
  LAYER M1 ;
        RECT 5.152 19.62 5.184 22.128 ;
  LAYER M3 ;
        RECT 5.152 19.64 5.184 19.672 ;
  LAYER M1 ;
        RECT 5.216 19.62 5.248 22.128 ;
  LAYER M3 ;
        RECT 5.216 22.076 5.248 22.108 ;
  LAYER M1 ;
        RECT 5.28 19.62 5.312 22.128 ;
  LAYER M3 ;
        RECT 5.28 19.64 5.312 19.672 ;
  LAYER M1 ;
        RECT 5.344 19.62 5.376 22.128 ;
  LAYER M3 ;
        RECT 5.344 22.076 5.376 22.108 ;
  LAYER M1 ;
        RECT 5.408 19.62 5.44 22.128 ;
  LAYER M3 ;
        RECT 5.408 19.64 5.44 19.672 ;
  LAYER M1 ;
        RECT 5.472 19.62 5.504 22.128 ;
  LAYER M3 ;
        RECT 5.472 22.076 5.504 22.108 ;
  LAYER M1 ;
        RECT 5.536 19.62 5.568 22.128 ;
  LAYER M3 ;
        RECT 5.536 19.64 5.568 19.672 ;
  LAYER M1 ;
        RECT 5.6 19.62 5.632 22.128 ;
  LAYER M3 ;
        RECT 5.6 22.076 5.632 22.108 ;
  LAYER M1 ;
        RECT 5.664 19.62 5.696 22.128 ;
  LAYER M3 ;
        RECT 5.664 19.64 5.696 19.672 ;
  LAYER M1 ;
        RECT 5.728 19.62 5.76 22.128 ;
  LAYER M3 ;
        RECT 5.728 22.076 5.76 22.108 ;
  LAYER M1 ;
        RECT 5.792 19.62 5.824 22.128 ;
  LAYER M3 ;
        RECT 5.792 19.64 5.824 19.672 ;
  LAYER M1 ;
        RECT 5.856 19.62 5.888 22.128 ;
  LAYER M3 ;
        RECT 5.856 22.076 5.888 22.108 ;
  LAYER M1 ;
        RECT 5.92 19.62 5.952 22.128 ;
  LAYER M3 ;
        RECT 5.92 19.64 5.952 19.672 ;
  LAYER M1 ;
        RECT 5.984 19.62 6.016 22.128 ;
  LAYER M3 ;
        RECT 5.984 22.076 6.016 22.108 ;
  LAYER M1 ;
        RECT 6.048 19.62 6.08 22.128 ;
  LAYER M3 ;
        RECT 6.048 19.64 6.08 19.672 ;
  LAYER M1 ;
        RECT 6.112 19.62 6.144 22.128 ;
  LAYER M3 ;
        RECT 6.112 22.076 6.144 22.108 ;
  LAYER M1 ;
        RECT 6.176 19.62 6.208 22.128 ;
  LAYER M3 ;
        RECT 6.176 19.64 6.208 19.672 ;
  LAYER M1 ;
        RECT 6.24 19.62 6.272 22.128 ;
  LAYER M3 ;
        RECT 6.24 22.076 6.272 22.108 ;
  LAYER M1 ;
        RECT 6.304 19.62 6.336 22.128 ;
  LAYER M3 ;
        RECT 6.304 19.64 6.336 19.672 ;
  LAYER M1 ;
        RECT 6.368 19.62 6.4 22.128 ;
  LAYER M3 ;
        RECT 6.368 22.076 6.4 22.108 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 22.128 ;
  LAYER M3 ;
        RECT 4.064 19.704 4.096 19.736 ;
  LAYER M2 ;
        RECT 6.432 19.768 6.464 19.8 ;
  LAYER M2 ;
        RECT 4.064 19.832 4.096 19.864 ;
  LAYER M2 ;
        RECT 6.432 19.896 6.464 19.928 ;
  LAYER M2 ;
        RECT 4.064 19.96 4.096 19.992 ;
  LAYER M2 ;
        RECT 6.432 20.024 6.464 20.056 ;
  LAYER M2 ;
        RECT 4.064 20.088 4.096 20.12 ;
  LAYER M2 ;
        RECT 6.432 20.152 6.464 20.184 ;
  LAYER M2 ;
        RECT 4.064 20.216 4.096 20.248 ;
  LAYER M2 ;
        RECT 6.432 20.28 6.464 20.312 ;
  LAYER M2 ;
        RECT 4.064 20.344 4.096 20.376 ;
  LAYER M2 ;
        RECT 6.432 20.408 6.464 20.44 ;
  LAYER M2 ;
        RECT 4.064 20.472 4.096 20.504 ;
  LAYER M2 ;
        RECT 6.432 20.536 6.464 20.568 ;
  LAYER M2 ;
        RECT 4.064 20.6 4.096 20.632 ;
  LAYER M2 ;
        RECT 6.432 20.664 6.464 20.696 ;
  LAYER M2 ;
        RECT 4.064 20.728 4.096 20.76 ;
  LAYER M2 ;
        RECT 6.432 20.792 6.464 20.824 ;
  LAYER M2 ;
        RECT 4.064 20.856 4.096 20.888 ;
  LAYER M2 ;
        RECT 6.432 20.92 6.464 20.952 ;
  LAYER M2 ;
        RECT 4.064 20.984 4.096 21.016 ;
  LAYER M2 ;
        RECT 6.432 21.048 6.464 21.08 ;
  LAYER M2 ;
        RECT 4.064 21.112 4.096 21.144 ;
  LAYER M2 ;
        RECT 6.432 21.176 6.464 21.208 ;
  LAYER M2 ;
        RECT 4.064 21.24 4.096 21.272 ;
  LAYER M2 ;
        RECT 6.432 21.304 6.464 21.336 ;
  LAYER M2 ;
        RECT 4.064 21.368 4.096 21.4 ;
  LAYER M2 ;
        RECT 6.432 21.432 6.464 21.464 ;
  LAYER M2 ;
        RECT 4.064 21.496 4.096 21.528 ;
  LAYER M2 ;
        RECT 6.432 21.56 6.464 21.592 ;
  LAYER M2 ;
        RECT 4.064 21.624 4.096 21.656 ;
  LAYER M2 ;
        RECT 6.432 21.688 6.464 21.72 ;
  LAYER M2 ;
        RECT 4.064 21.752 4.096 21.784 ;
  LAYER M2 ;
        RECT 6.432 21.816 6.464 21.848 ;
  LAYER M2 ;
        RECT 4.064 21.88 4.096 21.912 ;
  LAYER M2 ;
        RECT 6.432 21.944 6.464 21.976 ;
  LAYER M2 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M1 ;
        RECT 4.064 22.728 4.096 25.236 ;
  LAYER M3 ;
        RECT 4.064 25.184 4.096 25.216 ;
  LAYER M1 ;
        RECT 4.128 22.728 4.16 25.236 ;
  LAYER M3 ;
        RECT 4.128 22.748 4.16 22.78 ;
  LAYER M1 ;
        RECT 4.192 22.728 4.224 25.236 ;
  LAYER M3 ;
        RECT 4.192 25.184 4.224 25.216 ;
  LAYER M1 ;
        RECT 4.256 22.728 4.288 25.236 ;
  LAYER M3 ;
        RECT 4.256 22.748 4.288 22.78 ;
  LAYER M1 ;
        RECT 4.32 22.728 4.352 25.236 ;
  LAYER M3 ;
        RECT 4.32 25.184 4.352 25.216 ;
  LAYER M1 ;
        RECT 4.384 22.728 4.416 25.236 ;
  LAYER M3 ;
        RECT 4.384 22.748 4.416 22.78 ;
  LAYER M1 ;
        RECT 4.448 22.728 4.48 25.236 ;
  LAYER M3 ;
        RECT 4.448 25.184 4.48 25.216 ;
  LAYER M1 ;
        RECT 4.512 22.728 4.544 25.236 ;
  LAYER M3 ;
        RECT 4.512 22.748 4.544 22.78 ;
  LAYER M1 ;
        RECT 4.576 22.728 4.608 25.236 ;
  LAYER M3 ;
        RECT 4.576 25.184 4.608 25.216 ;
  LAYER M1 ;
        RECT 4.64 22.728 4.672 25.236 ;
  LAYER M3 ;
        RECT 4.64 22.748 4.672 22.78 ;
  LAYER M1 ;
        RECT 4.704 22.728 4.736 25.236 ;
  LAYER M3 ;
        RECT 4.704 25.184 4.736 25.216 ;
  LAYER M1 ;
        RECT 4.768 22.728 4.8 25.236 ;
  LAYER M3 ;
        RECT 4.768 22.748 4.8 22.78 ;
  LAYER M1 ;
        RECT 4.832 22.728 4.864 25.236 ;
  LAYER M3 ;
        RECT 4.832 25.184 4.864 25.216 ;
  LAYER M1 ;
        RECT 4.896 22.728 4.928 25.236 ;
  LAYER M3 ;
        RECT 4.896 22.748 4.928 22.78 ;
  LAYER M1 ;
        RECT 4.96 22.728 4.992 25.236 ;
  LAYER M3 ;
        RECT 4.96 25.184 4.992 25.216 ;
  LAYER M1 ;
        RECT 5.024 22.728 5.056 25.236 ;
  LAYER M3 ;
        RECT 5.024 22.748 5.056 22.78 ;
  LAYER M1 ;
        RECT 5.088 22.728 5.12 25.236 ;
  LAYER M3 ;
        RECT 5.088 25.184 5.12 25.216 ;
  LAYER M1 ;
        RECT 5.152 22.728 5.184 25.236 ;
  LAYER M3 ;
        RECT 5.152 22.748 5.184 22.78 ;
  LAYER M1 ;
        RECT 5.216 22.728 5.248 25.236 ;
  LAYER M3 ;
        RECT 5.216 25.184 5.248 25.216 ;
  LAYER M1 ;
        RECT 5.28 22.728 5.312 25.236 ;
  LAYER M3 ;
        RECT 5.28 22.748 5.312 22.78 ;
  LAYER M1 ;
        RECT 5.344 22.728 5.376 25.236 ;
  LAYER M3 ;
        RECT 5.344 25.184 5.376 25.216 ;
  LAYER M1 ;
        RECT 5.408 22.728 5.44 25.236 ;
  LAYER M3 ;
        RECT 5.408 22.748 5.44 22.78 ;
  LAYER M1 ;
        RECT 5.472 22.728 5.504 25.236 ;
  LAYER M3 ;
        RECT 5.472 25.184 5.504 25.216 ;
  LAYER M1 ;
        RECT 5.536 22.728 5.568 25.236 ;
  LAYER M3 ;
        RECT 5.536 22.748 5.568 22.78 ;
  LAYER M1 ;
        RECT 5.6 22.728 5.632 25.236 ;
  LAYER M3 ;
        RECT 5.6 25.184 5.632 25.216 ;
  LAYER M1 ;
        RECT 5.664 22.728 5.696 25.236 ;
  LAYER M3 ;
        RECT 5.664 22.748 5.696 22.78 ;
  LAYER M1 ;
        RECT 5.728 22.728 5.76 25.236 ;
  LAYER M3 ;
        RECT 5.728 25.184 5.76 25.216 ;
  LAYER M1 ;
        RECT 5.792 22.728 5.824 25.236 ;
  LAYER M3 ;
        RECT 5.792 22.748 5.824 22.78 ;
  LAYER M1 ;
        RECT 5.856 22.728 5.888 25.236 ;
  LAYER M3 ;
        RECT 5.856 25.184 5.888 25.216 ;
  LAYER M1 ;
        RECT 5.92 22.728 5.952 25.236 ;
  LAYER M3 ;
        RECT 5.92 22.748 5.952 22.78 ;
  LAYER M1 ;
        RECT 5.984 22.728 6.016 25.236 ;
  LAYER M3 ;
        RECT 5.984 25.184 6.016 25.216 ;
  LAYER M1 ;
        RECT 6.048 22.728 6.08 25.236 ;
  LAYER M3 ;
        RECT 6.048 22.748 6.08 22.78 ;
  LAYER M1 ;
        RECT 6.112 22.728 6.144 25.236 ;
  LAYER M3 ;
        RECT 6.112 25.184 6.144 25.216 ;
  LAYER M1 ;
        RECT 6.176 22.728 6.208 25.236 ;
  LAYER M3 ;
        RECT 6.176 22.748 6.208 22.78 ;
  LAYER M1 ;
        RECT 6.24 22.728 6.272 25.236 ;
  LAYER M3 ;
        RECT 6.24 25.184 6.272 25.216 ;
  LAYER M1 ;
        RECT 6.304 22.728 6.336 25.236 ;
  LAYER M3 ;
        RECT 6.304 22.748 6.336 22.78 ;
  LAYER M1 ;
        RECT 6.368 22.728 6.4 25.236 ;
  LAYER M3 ;
        RECT 6.368 25.184 6.4 25.216 ;
  LAYER M1 ;
        RECT 6.432 22.728 6.464 25.236 ;
  LAYER M3 ;
        RECT 4.064 22.812 4.096 22.844 ;
  LAYER M2 ;
        RECT 6.432 22.876 6.464 22.908 ;
  LAYER M2 ;
        RECT 4.064 22.94 4.096 22.972 ;
  LAYER M2 ;
        RECT 6.432 23.004 6.464 23.036 ;
  LAYER M2 ;
        RECT 4.064 23.068 4.096 23.1 ;
  LAYER M2 ;
        RECT 6.432 23.132 6.464 23.164 ;
  LAYER M2 ;
        RECT 4.064 23.196 4.096 23.228 ;
  LAYER M2 ;
        RECT 6.432 23.26 6.464 23.292 ;
  LAYER M2 ;
        RECT 4.064 23.324 4.096 23.356 ;
  LAYER M2 ;
        RECT 6.432 23.388 6.464 23.42 ;
  LAYER M2 ;
        RECT 4.064 23.452 4.096 23.484 ;
  LAYER M2 ;
        RECT 6.432 23.516 6.464 23.548 ;
  LAYER M2 ;
        RECT 4.064 23.58 4.096 23.612 ;
  LAYER M2 ;
        RECT 6.432 23.644 6.464 23.676 ;
  LAYER M2 ;
        RECT 4.064 23.708 4.096 23.74 ;
  LAYER M2 ;
        RECT 6.432 23.772 6.464 23.804 ;
  LAYER M2 ;
        RECT 4.064 23.836 4.096 23.868 ;
  LAYER M2 ;
        RECT 6.432 23.9 6.464 23.932 ;
  LAYER M2 ;
        RECT 4.064 23.964 4.096 23.996 ;
  LAYER M2 ;
        RECT 6.432 24.028 6.464 24.06 ;
  LAYER M2 ;
        RECT 4.064 24.092 4.096 24.124 ;
  LAYER M2 ;
        RECT 6.432 24.156 6.464 24.188 ;
  LAYER M2 ;
        RECT 4.064 24.22 4.096 24.252 ;
  LAYER M2 ;
        RECT 6.432 24.284 6.464 24.316 ;
  LAYER M2 ;
        RECT 4.064 24.348 4.096 24.38 ;
  LAYER M2 ;
        RECT 6.432 24.412 6.464 24.444 ;
  LAYER M2 ;
        RECT 4.064 24.476 4.096 24.508 ;
  LAYER M2 ;
        RECT 6.432 24.54 6.464 24.572 ;
  LAYER M2 ;
        RECT 4.064 24.604 4.096 24.636 ;
  LAYER M2 ;
        RECT 6.432 24.668 6.464 24.7 ;
  LAYER M2 ;
        RECT 4.064 24.732 4.096 24.764 ;
  LAYER M2 ;
        RECT 6.432 24.796 6.464 24.828 ;
  LAYER M2 ;
        RECT 4.064 24.86 4.096 24.892 ;
  LAYER M2 ;
        RECT 6.432 24.924 6.464 24.956 ;
  LAYER M2 ;
        RECT 4.064 24.988 4.096 25.02 ;
  LAYER M2 ;
        RECT 6.432 25.052 6.464 25.084 ;
  LAYER M2 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M1 ;
        RECT 7.36 0.972 7.392 3.48 ;
  LAYER M3 ;
        RECT 7.36 3.428 7.392 3.46 ;
  LAYER M1 ;
        RECT 7.424 0.972 7.456 3.48 ;
  LAYER M3 ;
        RECT 7.424 0.992 7.456 1.024 ;
  LAYER M1 ;
        RECT 7.488 0.972 7.52 3.48 ;
  LAYER M3 ;
        RECT 7.488 3.428 7.52 3.46 ;
  LAYER M1 ;
        RECT 7.552 0.972 7.584 3.48 ;
  LAYER M3 ;
        RECT 7.552 0.992 7.584 1.024 ;
  LAYER M1 ;
        RECT 7.616 0.972 7.648 3.48 ;
  LAYER M3 ;
        RECT 7.616 3.428 7.648 3.46 ;
  LAYER M1 ;
        RECT 7.68 0.972 7.712 3.48 ;
  LAYER M3 ;
        RECT 7.68 0.992 7.712 1.024 ;
  LAYER M1 ;
        RECT 7.744 0.972 7.776 3.48 ;
  LAYER M3 ;
        RECT 7.744 3.428 7.776 3.46 ;
  LAYER M1 ;
        RECT 7.808 0.972 7.84 3.48 ;
  LAYER M3 ;
        RECT 7.808 0.992 7.84 1.024 ;
  LAYER M1 ;
        RECT 7.872 0.972 7.904 3.48 ;
  LAYER M3 ;
        RECT 7.872 3.428 7.904 3.46 ;
  LAYER M1 ;
        RECT 7.936 0.972 7.968 3.48 ;
  LAYER M3 ;
        RECT 7.936 0.992 7.968 1.024 ;
  LAYER M1 ;
        RECT 8 0.972 8.032 3.48 ;
  LAYER M3 ;
        RECT 8 3.428 8.032 3.46 ;
  LAYER M1 ;
        RECT 8.064 0.972 8.096 3.48 ;
  LAYER M3 ;
        RECT 8.064 0.992 8.096 1.024 ;
  LAYER M1 ;
        RECT 8.128 0.972 8.16 3.48 ;
  LAYER M3 ;
        RECT 8.128 3.428 8.16 3.46 ;
  LAYER M1 ;
        RECT 8.192 0.972 8.224 3.48 ;
  LAYER M3 ;
        RECT 8.192 0.992 8.224 1.024 ;
  LAYER M1 ;
        RECT 8.256 0.972 8.288 3.48 ;
  LAYER M3 ;
        RECT 8.256 3.428 8.288 3.46 ;
  LAYER M1 ;
        RECT 8.32 0.972 8.352 3.48 ;
  LAYER M3 ;
        RECT 8.32 0.992 8.352 1.024 ;
  LAYER M1 ;
        RECT 8.384 0.972 8.416 3.48 ;
  LAYER M3 ;
        RECT 8.384 3.428 8.416 3.46 ;
  LAYER M1 ;
        RECT 8.448 0.972 8.48 3.48 ;
  LAYER M3 ;
        RECT 8.448 0.992 8.48 1.024 ;
  LAYER M1 ;
        RECT 8.512 0.972 8.544 3.48 ;
  LAYER M3 ;
        RECT 8.512 3.428 8.544 3.46 ;
  LAYER M1 ;
        RECT 8.576 0.972 8.608 3.48 ;
  LAYER M3 ;
        RECT 8.576 0.992 8.608 1.024 ;
  LAYER M1 ;
        RECT 8.64 0.972 8.672 3.48 ;
  LAYER M3 ;
        RECT 8.64 3.428 8.672 3.46 ;
  LAYER M1 ;
        RECT 8.704 0.972 8.736 3.48 ;
  LAYER M3 ;
        RECT 8.704 0.992 8.736 1.024 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 3.48 ;
  LAYER M3 ;
        RECT 8.768 3.428 8.8 3.46 ;
  LAYER M1 ;
        RECT 8.832 0.972 8.864 3.48 ;
  LAYER M3 ;
        RECT 8.832 0.992 8.864 1.024 ;
  LAYER M1 ;
        RECT 8.896 0.972 8.928 3.48 ;
  LAYER M3 ;
        RECT 8.896 3.428 8.928 3.46 ;
  LAYER M1 ;
        RECT 8.96 0.972 8.992 3.48 ;
  LAYER M3 ;
        RECT 8.96 0.992 8.992 1.024 ;
  LAYER M1 ;
        RECT 9.024 0.972 9.056 3.48 ;
  LAYER M3 ;
        RECT 9.024 3.428 9.056 3.46 ;
  LAYER M1 ;
        RECT 9.088 0.972 9.12 3.48 ;
  LAYER M3 ;
        RECT 9.088 0.992 9.12 1.024 ;
  LAYER M1 ;
        RECT 9.152 0.972 9.184 3.48 ;
  LAYER M3 ;
        RECT 9.152 3.428 9.184 3.46 ;
  LAYER M1 ;
        RECT 9.216 0.972 9.248 3.48 ;
  LAYER M3 ;
        RECT 9.216 0.992 9.248 1.024 ;
  LAYER M1 ;
        RECT 9.28 0.972 9.312 3.48 ;
  LAYER M3 ;
        RECT 9.28 3.428 9.312 3.46 ;
  LAYER M1 ;
        RECT 9.344 0.972 9.376 3.48 ;
  LAYER M3 ;
        RECT 9.344 0.992 9.376 1.024 ;
  LAYER M1 ;
        RECT 9.408 0.972 9.44 3.48 ;
  LAYER M3 ;
        RECT 9.408 3.428 9.44 3.46 ;
  LAYER M1 ;
        RECT 9.472 0.972 9.504 3.48 ;
  LAYER M3 ;
        RECT 9.472 0.992 9.504 1.024 ;
  LAYER M1 ;
        RECT 9.536 0.972 9.568 3.48 ;
  LAYER M3 ;
        RECT 9.536 3.428 9.568 3.46 ;
  LAYER M1 ;
        RECT 9.6 0.972 9.632 3.48 ;
  LAYER M3 ;
        RECT 9.6 0.992 9.632 1.024 ;
  LAYER M1 ;
        RECT 9.664 0.972 9.696 3.48 ;
  LAYER M3 ;
        RECT 9.664 3.428 9.696 3.46 ;
  LAYER M1 ;
        RECT 9.728 0.972 9.76 3.48 ;
  LAYER M3 ;
        RECT 7.36 1.056 7.392 1.088 ;
  LAYER M2 ;
        RECT 9.728 1.12 9.76 1.152 ;
  LAYER M2 ;
        RECT 7.36 1.184 7.392 1.216 ;
  LAYER M2 ;
        RECT 9.728 1.248 9.76 1.28 ;
  LAYER M2 ;
        RECT 7.36 1.312 7.392 1.344 ;
  LAYER M2 ;
        RECT 9.728 1.376 9.76 1.408 ;
  LAYER M2 ;
        RECT 7.36 1.44 7.392 1.472 ;
  LAYER M2 ;
        RECT 9.728 1.504 9.76 1.536 ;
  LAYER M2 ;
        RECT 7.36 1.568 7.392 1.6 ;
  LAYER M2 ;
        RECT 9.728 1.632 9.76 1.664 ;
  LAYER M2 ;
        RECT 7.36 1.696 7.392 1.728 ;
  LAYER M2 ;
        RECT 9.728 1.76 9.76 1.792 ;
  LAYER M2 ;
        RECT 7.36 1.824 7.392 1.856 ;
  LAYER M2 ;
        RECT 9.728 1.888 9.76 1.92 ;
  LAYER M2 ;
        RECT 7.36 1.952 7.392 1.984 ;
  LAYER M2 ;
        RECT 9.728 2.016 9.76 2.048 ;
  LAYER M2 ;
        RECT 7.36 2.08 7.392 2.112 ;
  LAYER M2 ;
        RECT 9.728 2.144 9.76 2.176 ;
  LAYER M2 ;
        RECT 7.36 2.208 7.392 2.24 ;
  LAYER M2 ;
        RECT 9.728 2.272 9.76 2.304 ;
  LAYER M2 ;
        RECT 7.36 2.336 7.392 2.368 ;
  LAYER M2 ;
        RECT 9.728 2.4 9.76 2.432 ;
  LAYER M2 ;
        RECT 7.36 2.464 7.392 2.496 ;
  LAYER M2 ;
        RECT 9.728 2.528 9.76 2.56 ;
  LAYER M2 ;
        RECT 7.36 2.592 7.392 2.624 ;
  LAYER M2 ;
        RECT 9.728 2.656 9.76 2.688 ;
  LAYER M2 ;
        RECT 7.36 2.72 7.392 2.752 ;
  LAYER M2 ;
        RECT 9.728 2.784 9.76 2.816 ;
  LAYER M2 ;
        RECT 7.36 2.848 7.392 2.88 ;
  LAYER M2 ;
        RECT 9.728 2.912 9.76 2.944 ;
  LAYER M2 ;
        RECT 7.36 2.976 7.392 3.008 ;
  LAYER M2 ;
        RECT 9.728 3.04 9.76 3.072 ;
  LAYER M2 ;
        RECT 7.36 3.104 7.392 3.136 ;
  LAYER M2 ;
        RECT 9.728 3.168 9.76 3.2 ;
  LAYER M2 ;
        RECT 7.36 3.232 7.392 3.264 ;
  LAYER M2 ;
        RECT 9.728 3.296 9.76 3.328 ;
  LAYER M2 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M1 ;
        RECT 7.36 4.08 7.392 6.588 ;
  LAYER M3 ;
        RECT 7.36 6.536 7.392 6.568 ;
  LAYER M1 ;
        RECT 7.424 4.08 7.456 6.588 ;
  LAYER M3 ;
        RECT 7.424 4.1 7.456 4.132 ;
  LAYER M1 ;
        RECT 7.488 4.08 7.52 6.588 ;
  LAYER M3 ;
        RECT 7.488 6.536 7.52 6.568 ;
  LAYER M1 ;
        RECT 7.552 4.08 7.584 6.588 ;
  LAYER M3 ;
        RECT 7.552 4.1 7.584 4.132 ;
  LAYER M1 ;
        RECT 7.616 4.08 7.648 6.588 ;
  LAYER M3 ;
        RECT 7.616 6.536 7.648 6.568 ;
  LAYER M1 ;
        RECT 7.68 4.08 7.712 6.588 ;
  LAYER M3 ;
        RECT 7.68 4.1 7.712 4.132 ;
  LAYER M1 ;
        RECT 7.744 4.08 7.776 6.588 ;
  LAYER M3 ;
        RECT 7.744 6.536 7.776 6.568 ;
  LAYER M1 ;
        RECT 7.808 4.08 7.84 6.588 ;
  LAYER M3 ;
        RECT 7.808 4.1 7.84 4.132 ;
  LAYER M1 ;
        RECT 7.872 4.08 7.904 6.588 ;
  LAYER M3 ;
        RECT 7.872 6.536 7.904 6.568 ;
  LAYER M1 ;
        RECT 7.936 4.08 7.968 6.588 ;
  LAYER M3 ;
        RECT 7.936 4.1 7.968 4.132 ;
  LAYER M1 ;
        RECT 8 4.08 8.032 6.588 ;
  LAYER M3 ;
        RECT 8 6.536 8.032 6.568 ;
  LAYER M1 ;
        RECT 8.064 4.08 8.096 6.588 ;
  LAYER M3 ;
        RECT 8.064 4.1 8.096 4.132 ;
  LAYER M1 ;
        RECT 8.128 4.08 8.16 6.588 ;
  LAYER M3 ;
        RECT 8.128 6.536 8.16 6.568 ;
  LAYER M1 ;
        RECT 8.192 4.08 8.224 6.588 ;
  LAYER M3 ;
        RECT 8.192 4.1 8.224 4.132 ;
  LAYER M1 ;
        RECT 8.256 4.08 8.288 6.588 ;
  LAYER M3 ;
        RECT 8.256 6.536 8.288 6.568 ;
  LAYER M1 ;
        RECT 8.32 4.08 8.352 6.588 ;
  LAYER M3 ;
        RECT 8.32 4.1 8.352 4.132 ;
  LAYER M1 ;
        RECT 8.384 4.08 8.416 6.588 ;
  LAYER M3 ;
        RECT 8.384 6.536 8.416 6.568 ;
  LAYER M1 ;
        RECT 8.448 4.08 8.48 6.588 ;
  LAYER M3 ;
        RECT 8.448 4.1 8.48 4.132 ;
  LAYER M1 ;
        RECT 8.512 4.08 8.544 6.588 ;
  LAYER M3 ;
        RECT 8.512 6.536 8.544 6.568 ;
  LAYER M1 ;
        RECT 8.576 4.08 8.608 6.588 ;
  LAYER M3 ;
        RECT 8.576 4.1 8.608 4.132 ;
  LAYER M1 ;
        RECT 8.64 4.08 8.672 6.588 ;
  LAYER M3 ;
        RECT 8.64 6.536 8.672 6.568 ;
  LAYER M1 ;
        RECT 8.704 4.08 8.736 6.588 ;
  LAYER M3 ;
        RECT 8.704 4.1 8.736 4.132 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 6.588 ;
  LAYER M3 ;
        RECT 8.768 6.536 8.8 6.568 ;
  LAYER M1 ;
        RECT 8.832 4.08 8.864 6.588 ;
  LAYER M3 ;
        RECT 8.832 4.1 8.864 4.132 ;
  LAYER M1 ;
        RECT 8.896 4.08 8.928 6.588 ;
  LAYER M3 ;
        RECT 8.896 6.536 8.928 6.568 ;
  LAYER M1 ;
        RECT 8.96 4.08 8.992 6.588 ;
  LAYER M3 ;
        RECT 8.96 4.1 8.992 4.132 ;
  LAYER M1 ;
        RECT 9.024 4.08 9.056 6.588 ;
  LAYER M3 ;
        RECT 9.024 6.536 9.056 6.568 ;
  LAYER M1 ;
        RECT 9.088 4.08 9.12 6.588 ;
  LAYER M3 ;
        RECT 9.088 4.1 9.12 4.132 ;
  LAYER M1 ;
        RECT 9.152 4.08 9.184 6.588 ;
  LAYER M3 ;
        RECT 9.152 6.536 9.184 6.568 ;
  LAYER M1 ;
        RECT 9.216 4.08 9.248 6.588 ;
  LAYER M3 ;
        RECT 9.216 4.1 9.248 4.132 ;
  LAYER M1 ;
        RECT 9.28 4.08 9.312 6.588 ;
  LAYER M3 ;
        RECT 9.28 6.536 9.312 6.568 ;
  LAYER M1 ;
        RECT 9.344 4.08 9.376 6.588 ;
  LAYER M3 ;
        RECT 9.344 4.1 9.376 4.132 ;
  LAYER M1 ;
        RECT 9.408 4.08 9.44 6.588 ;
  LAYER M3 ;
        RECT 9.408 6.536 9.44 6.568 ;
  LAYER M1 ;
        RECT 9.472 4.08 9.504 6.588 ;
  LAYER M3 ;
        RECT 9.472 4.1 9.504 4.132 ;
  LAYER M1 ;
        RECT 9.536 4.08 9.568 6.588 ;
  LAYER M3 ;
        RECT 9.536 6.536 9.568 6.568 ;
  LAYER M1 ;
        RECT 9.6 4.08 9.632 6.588 ;
  LAYER M3 ;
        RECT 9.6 4.1 9.632 4.132 ;
  LAYER M1 ;
        RECT 9.664 4.08 9.696 6.588 ;
  LAYER M3 ;
        RECT 9.664 6.536 9.696 6.568 ;
  LAYER M1 ;
        RECT 9.728 4.08 9.76 6.588 ;
  LAYER M3 ;
        RECT 7.36 4.164 7.392 4.196 ;
  LAYER M2 ;
        RECT 9.728 4.228 9.76 4.26 ;
  LAYER M2 ;
        RECT 7.36 4.292 7.392 4.324 ;
  LAYER M2 ;
        RECT 9.728 4.356 9.76 4.388 ;
  LAYER M2 ;
        RECT 7.36 4.42 7.392 4.452 ;
  LAYER M2 ;
        RECT 9.728 4.484 9.76 4.516 ;
  LAYER M2 ;
        RECT 7.36 4.548 7.392 4.58 ;
  LAYER M2 ;
        RECT 9.728 4.612 9.76 4.644 ;
  LAYER M2 ;
        RECT 7.36 4.676 7.392 4.708 ;
  LAYER M2 ;
        RECT 9.728 4.74 9.76 4.772 ;
  LAYER M2 ;
        RECT 7.36 4.804 7.392 4.836 ;
  LAYER M2 ;
        RECT 9.728 4.868 9.76 4.9 ;
  LAYER M2 ;
        RECT 7.36 4.932 7.392 4.964 ;
  LAYER M2 ;
        RECT 9.728 4.996 9.76 5.028 ;
  LAYER M2 ;
        RECT 7.36 5.06 7.392 5.092 ;
  LAYER M2 ;
        RECT 9.728 5.124 9.76 5.156 ;
  LAYER M2 ;
        RECT 7.36 5.188 7.392 5.22 ;
  LAYER M2 ;
        RECT 9.728 5.252 9.76 5.284 ;
  LAYER M2 ;
        RECT 7.36 5.316 7.392 5.348 ;
  LAYER M2 ;
        RECT 9.728 5.38 9.76 5.412 ;
  LAYER M2 ;
        RECT 7.36 5.444 7.392 5.476 ;
  LAYER M2 ;
        RECT 9.728 5.508 9.76 5.54 ;
  LAYER M2 ;
        RECT 7.36 5.572 7.392 5.604 ;
  LAYER M2 ;
        RECT 9.728 5.636 9.76 5.668 ;
  LAYER M2 ;
        RECT 7.36 5.7 7.392 5.732 ;
  LAYER M2 ;
        RECT 9.728 5.764 9.76 5.796 ;
  LAYER M2 ;
        RECT 7.36 5.828 7.392 5.86 ;
  LAYER M2 ;
        RECT 9.728 5.892 9.76 5.924 ;
  LAYER M2 ;
        RECT 7.36 5.956 7.392 5.988 ;
  LAYER M2 ;
        RECT 9.728 6.02 9.76 6.052 ;
  LAYER M2 ;
        RECT 7.36 6.084 7.392 6.116 ;
  LAYER M2 ;
        RECT 9.728 6.148 9.76 6.18 ;
  LAYER M2 ;
        RECT 7.36 6.212 7.392 6.244 ;
  LAYER M2 ;
        RECT 9.728 6.276 9.76 6.308 ;
  LAYER M2 ;
        RECT 7.36 6.34 7.392 6.372 ;
  LAYER M2 ;
        RECT 9.728 6.404 9.76 6.436 ;
  LAYER M2 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M1 ;
        RECT 7.36 7.188 7.392 9.696 ;
  LAYER M3 ;
        RECT 7.36 9.644 7.392 9.676 ;
  LAYER M1 ;
        RECT 7.424 7.188 7.456 9.696 ;
  LAYER M3 ;
        RECT 7.424 7.208 7.456 7.24 ;
  LAYER M1 ;
        RECT 7.488 7.188 7.52 9.696 ;
  LAYER M3 ;
        RECT 7.488 9.644 7.52 9.676 ;
  LAYER M1 ;
        RECT 7.552 7.188 7.584 9.696 ;
  LAYER M3 ;
        RECT 7.552 7.208 7.584 7.24 ;
  LAYER M1 ;
        RECT 7.616 7.188 7.648 9.696 ;
  LAYER M3 ;
        RECT 7.616 9.644 7.648 9.676 ;
  LAYER M1 ;
        RECT 7.68 7.188 7.712 9.696 ;
  LAYER M3 ;
        RECT 7.68 7.208 7.712 7.24 ;
  LAYER M1 ;
        RECT 7.744 7.188 7.776 9.696 ;
  LAYER M3 ;
        RECT 7.744 9.644 7.776 9.676 ;
  LAYER M1 ;
        RECT 7.808 7.188 7.84 9.696 ;
  LAYER M3 ;
        RECT 7.808 7.208 7.84 7.24 ;
  LAYER M1 ;
        RECT 7.872 7.188 7.904 9.696 ;
  LAYER M3 ;
        RECT 7.872 9.644 7.904 9.676 ;
  LAYER M1 ;
        RECT 7.936 7.188 7.968 9.696 ;
  LAYER M3 ;
        RECT 7.936 7.208 7.968 7.24 ;
  LAYER M1 ;
        RECT 8 7.188 8.032 9.696 ;
  LAYER M3 ;
        RECT 8 9.644 8.032 9.676 ;
  LAYER M1 ;
        RECT 8.064 7.188 8.096 9.696 ;
  LAYER M3 ;
        RECT 8.064 7.208 8.096 7.24 ;
  LAYER M1 ;
        RECT 8.128 7.188 8.16 9.696 ;
  LAYER M3 ;
        RECT 8.128 9.644 8.16 9.676 ;
  LAYER M1 ;
        RECT 8.192 7.188 8.224 9.696 ;
  LAYER M3 ;
        RECT 8.192 7.208 8.224 7.24 ;
  LAYER M1 ;
        RECT 8.256 7.188 8.288 9.696 ;
  LAYER M3 ;
        RECT 8.256 9.644 8.288 9.676 ;
  LAYER M1 ;
        RECT 8.32 7.188 8.352 9.696 ;
  LAYER M3 ;
        RECT 8.32 7.208 8.352 7.24 ;
  LAYER M1 ;
        RECT 8.384 7.188 8.416 9.696 ;
  LAYER M3 ;
        RECT 8.384 9.644 8.416 9.676 ;
  LAYER M1 ;
        RECT 8.448 7.188 8.48 9.696 ;
  LAYER M3 ;
        RECT 8.448 7.208 8.48 7.24 ;
  LAYER M1 ;
        RECT 8.512 7.188 8.544 9.696 ;
  LAYER M3 ;
        RECT 8.512 9.644 8.544 9.676 ;
  LAYER M1 ;
        RECT 8.576 7.188 8.608 9.696 ;
  LAYER M3 ;
        RECT 8.576 7.208 8.608 7.24 ;
  LAYER M1 ;
        RECT 8.64 7.188 8.672 9.696 ;
  LAYER M3 ;
        RECT 8.64 9.644 8.672 9.676 ;
  LAYER M1 ;
        RECT 8.704 7.188 8.736 9.696 ;
  LAYER M3 ;
        RECT 8.704 7.208 8.736 7.24 ;
  LAYER M1 ;
        RECT 8.768 7.188 8.8 9.696 ;
  LAYER M3 ;
        RECT 8.768 9.644 8.8 9.676 ;
  LAYER M1 ;
        RECT 8.832 7.188 8.864 9.696 ;
  LAYER M3 ;
        RECT 8.832 7.208 8.864 7.24 ;
  LAYER M1 ;
        RECT 8.896 7.188 8.928 9.696 ;
  LAYER M3 ;
        RECT 8.896 9.644 8.928 9.676 ;
  LAYER M1 ;
        RECT 8.96 7.188 8.992 9.696 ;
  LAYER M3 ;
        RECT 8.96 7.208 8.992 7.24 ;
  LAYER M1 ;
        RECT 9.024 7.188 9.056 9.696 ;
  LAYER M3 ;
        RECT 9.024 9.644 9.056 9.676 ;
  LAYER M1 ;
        RECT 9.088 7.188 9.12 9.696 ;
  LAYER M3 ;
        RECT 9.088 7.208 9.12 7.24 ;
  LAYER M1 ;
        RECT 9.152 7.188 9.184 9.696 ;
  LAYER M3 ;
        RECT 9.152 9.644 9.184 9.676 ;
  LAYER M1 ;
        RECT 9.216 7.188 9.248 9.696 ;
  LAYER M3 ;
        RECT 9.216 7.208 9.248 7.24 ;
  LAYER M1 ;
        RECT 9.28 7.188 9.312 9.696 ;
  LAYER M3 ;
        RECT 9.28 9.644 9.312 9.676 ;
  LAYER M1 ;
        RECT 9.344 7.188 9.376 9.696 ;
  LAYER M3 ;
        RECT 9.344 7.208 9.376 7.24 ;
  LAYER M1 ;
        RECT 9.408 7.188 9.44 9.696 ;
  LAYER M3 ;
        RECT 9.408 9.644 9.44 9.676 ;
  LAYER M1 ;
        RECT 9.472 7.188 9.504 9.696 ;
  LAYER M3 ;
        RECT 9.472 7.208 9.504 7.24 ;
  LAYER M1 ;
        RECT 9.536 7.188 9.568 9.696 ;
  LAYER M3 ;
        RECT 9.536 9.644 9.568 9.676 ;
  LAYER M1 ;
        RECT 9.6 7.188 9.632 9.696 ;
  LAYER M3 ;
        RECT 9.6 7.208 9.632 7.24 ;
  LAYER M1 ;
        RECT 9.664 7.188 9.696 9.696 ;
  LAYER M3 ;
        RECT 9.664 9.644 9.696 9.676 ;
  LAYER M1 ;
        RECT 9.728 7.188 9.76 9.696 ;
  LAYER M3 ;
        RECT 7.36 7.272 7.392 7.304 ;
  LAYER M2 ;
        RECT 9.728 7.336 9.76 7.368 ;
  LAYER M2 ;
        RECT 7.36 7.4 7.392 7.432 ;
  LAYER M2 ;
        RECT 9.728 7.464 9.76 7.496 ;
  LAYER M2 ;
        RECT 7.36 7.528 7.392 7.56 ;
  LAYER M2 ;
        RECT 9.728 7.592 9.76 7.624 ;
  LAYER M2 ;
        RECT 7.36 7.656 7.392 7.688 ;
  LAYER M2 ;
        RECT 9.728 7.72 9.76 7.752 ;
  LAYER M2 ;
        RECT 7.36 7.784 7.392 7.816 ;
  LAYER M2 ;
        RECT 9.728 7.848 9.76 7.88 ;
  LAYER M2 ;
        RECT 7.36 7.912 7.392 7.944 ;
  LAYER M2 ;
        RECT 9.728 7.976 9.76 8.008 ;
  LAYER M2 ;
        RECT 7.36 8.04 7.392 8.072 ;
  LAYER M2 ;
        RECT 9.728 8.104 9.76 8.136 ;
  LAYER M2 ;
        RECT 7.36 8.168 7.392 8.2 ;
  LAYER M2 ;
        RECT 9.728 8.232 9.76 8.264 ;
  LAYER M2 ;
        RECT 7.36 8.296 7.392 8.328 ;
  LAYER M2 ;
        RECT 9.728 8.36 9.76 8.392 ;
  LAYER M2 ;
        RECT 7.36 8.424 7.392 8.456 ;
  LAYER M2 ;
        RECT 9.728 8.488 9.76 8.52 ;
  LAYER M2 ;
        RECT 7.36 8.552 7.392 8.584 ;
  LAYER M2 ;
        RECT 9.728 8.616 9.76 8.648 ;
  LAYER M2 ;
        RECT 7.36 8.68 7.392 8.712 ;
  LAYER M2 ;
        RECT 9.728 8.744 9.76 8.776 ;
  LAYER M2 ;
        RECT 7.36 8.808 7.392 8.84 ;
  LAYER M2 ;
        RECT 9.728 8.872 9.76 8.904 ;
  LAYER M2 ;
        RECT 7.36 8.936 7.392 8.968 ;
  LAYER M2 ;
        RECT 9.728 9 9.76 9.032 ;
  LAYER M2 ;
        RECT 7.36 9.064 7.392 9.096 ;
  LAYER M2 ;
        RECT 9.728 9.128 9.76 9.16 ;
  LAYER M2 ;
        RECT 7.36 9.192 7.392 9.224 ;
  LAYER M2 ;
        RECT 9.728 9.256 9.76 9.288 ;
  LAYER M2 ;
        RECT 7.36 9.32 7.392 9.352 ;
  LAYER M2 ;
        RECT 9.728 9.384 9.76 9.416 ;
  LAYER M2 ;
        RECT 7.36 9.448 7.392 9.48 ;
  LAYER M2 ;
        RECT 9.728 9.512 9.76 9.544 ;
  LAYER M2 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M1 ;
        RECT 7.36 10.296 7.392 12.804 ;
  LAYER M3 ;
        RECT 7.36 12.752 7.392 12.784 ;
  LAYER M1 ;
        RECT 7.424 10.296 7.456 12.804 ;
  LAYER M3 ;
        RECT 7.424 10.316 7.456 10.348 ;
  LAYER M1 ;
        RECT 7.488 10.296 7.52 12.804 ;
  LAYER M3 ;
        RECT 7.488 12.752 7.52 12.784 ;
  LAYER M1 ;
        RECT 7.552 10.296 7.584 12.804 ;
  LAYER M3 ;
        RECT 7.552 10.316 7.584 10.348 ;
  LAYER M1 ;
        RECT 7.616 10.296 7.648 12.804 ;
  LAYER M3 ;
        RECT 7.616 12.752 7.648 12.784 ;
  LAYER M1 ;
        RECT 7.68 10.296 7.712 12.804 ;
  LAYER M3 ;
        RECT 7.68 10.316 7.712 10.348 ;
  LAYER M1 ;
        RECT 7.744 10.296 7.776 12.804 ;
  LAYER M3 ;
        RECT 7.744 12.752 7.776 12.784 ;
  LAYER M1 ;
        RECT 7.808 10.296 7.84 12.804 ;
  LAYER M3 ;
        RECT 7.808 10.316 7.84 10.348 ;
  LAYER M1 ;
        RECT 7.872 10.296 7.904 12.804 ;
  LAYER M3 ;
        RECT 7.872 12.752 7.904 12.784 ;
  LAYER M1 ;
        RECT 7.936 10.296 7.968 12.804 ;
  LAYER M3 ;
        RECT 7.936 10.316 7.968 10.348 ;
  LAYER M1 ;
        RECT 8 10.296 8.032 12.804 ;
  LAYER M3 ;
        RECT 8 12.752 8.032 12.784 ;
  LAYER M1 ;
        RECT 8.064 10.296 8.096 12.804 ;
  LAYER M3 ;
        RECT 8.064 10.316 8.096 10.348 ;
  LAYER M1 ;
        RECT 8.128 10.296 8.16 12.804 ;
  LAYER M3 ;
        RECT 8.128 12.752 8.16 12.784 ;
  LAYER M1 ;
        RECT 8.192 10.296 8.224 12.804 ;
  LAYER M3 ;
        RECT 8.192 10.316 8.224 10.348 ;
  LAYER M1 ;
        RECT 8.256 10.296 8.288 12.804 ;
  LAYER M3 ;
        RECT 8.256 12.752 8.288 12.784 ;
  LAYER M1 ;
        RECT 8.32 10.296 8.352 12.804 ;
  LAYER M3 ;
        RECT 8.32 10.316 8.352 10.348 ;
  LAYER M1 ;
        RECT 8.384 10.296 8.416 12.804 ;
  LAYER M3 ;
        RECT 8.384 12.752 8.416 12.784 ;
  LAYER M1 ;
        RECT 8.448 10.296 8.48 12.804 ;
  LAYER M3 ;
        RECT 8.448 10.316 8.48 10.348 ;
  LAYER M1 ;
        RECT 8.512 10.296 8.544 12.804 ;
  LAYER M3 ;
        RECT 8.512 12.752 8.544 12.784 ;
  LAYER M1 ;
        RECT 8.576 10.296 8.608 12.804 ;
  LAYER M3 ;
        RECT 8.576 10.316 8.608 10.348 ;
  LAYER M1 ;
        RECT 8.64 10.296 8.672 12.804 ;
  LAYER M3 ;
        RECT 8.64 12.752 8.672 12.784 ;
  LAYER M1 ;
        RECT 8.704 10.296 8.736 12.804 ;
  LAYER M3 ;
        RECT 8.704 10.316 8.736 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 12.804 ;
  LAYER M3 ;
        RECT 8.768 12.752 8.8 12.784 ;
  LAYER M1 ;
        RECT 8.832 10.296 8.864 12.804 ;
  LAYER M3 ;
        RECT 8.832 10.316 8.864 10.348 ;
  LAYER M1 ;
        RECT 8.896 10.296 8.928 12.804 ;
  LAYER M3 ;
        RECT 8.896 12.752 8.928 12.784 ;
  LAYER M1 ;
        RECT 8.96 10.296 8.992 12.804 ;
  LAYER M3 ;
        RECT 8.96 10.316 8.992 10.348 ;
  LAYER M1 ;
        RECT 9.024 10.296 9.056 12.804 ;
  LAYER M3 ;
        RECT 9.024 12.752 9.056 12.784 ;
  LAYER M1 ;
        RECT 9.088 10.296 9.12 12.804 ;
  LAYER M3 ;
        RECT 9.088 10.316 9.12 10.348 ;
  LAYER M1 ;
        RECT 9.152 10.296 9.184 12.804 ;
  LAYER M3 ;
        RECT 9.152 12.752 9.184 12.784 ;
  LAYER M1 ;
        RECT 9.216 10.296 9.248 12.804 ;
  LAYER M3 ;
        RECT 9.216 10.316 9.248 10.348 ;
  LAYER M1 ;
        RECT 9.28 10.296 9.312 12.804 ;
  LAYER M3 ;
        RECT 9.28 12.752 9.312 12.784 ;
  LAYER M1 ;
        RECT 9.344 10.296 9.376 12.804 ;
  LAYER M3 ;
        RECT 9.344 10.316 9.376 10.348 ;
  LAYER M1 ;
        RECT 9.408 10.296 9.44 12.804 ;
  LAYER M3 ;
        RECT 9.408 12.752 9.44 12.784 ;
  LAYER M1 ;
        RECT 9.472 10.296 9.504 12.804 ;
  LAYER M3 ;
        RECT 9.472 10.316 9.504 10.348 ;
  LAYER M1 ;
        RECT 9.536 10.296 9.568 12.804 ;
  LAYER M3 ;
        RECT 9.536 12.752 9.568 12.784 ;
  LAYER M1 ;
        RECT 9.6 10.296 9.632 12.804 ;
  LAYER M3 ;
        RECT 9.6 10.316 9.632 10.348 ;
  LAYER M1 ;
        RECT 9.664 10.296 9.696 12.804 ;
  LAYER M3 ;
        RECT 9.664 12.752 9.696 12.784 ;
  LAYER M1 ;
        RECT 9.728 10.296 9.76 12.804 ;
  LAYER M3 ;
        RECT 7.36 10.38 7.392 10.412 ;
  LAYER M2 ;
        RECT 9.728 10.444 9.76 10.476 ;
  LAYER M2 ;
        RECT 7.36 10.508 7.392 10.54 ;
  LAYER M2 ;
        RECT 9.728 10.572 9.76 10.604 ;
  LAYER M2 ;
        RECT 7.36 10.636 7.392 10.668 ;
  LAYER M2 ;
        RECT 9.728 10.7 9.76 10.732 ;
  LAYER M2 ;
        RECT 7.36 10.764 7.392 10.796 ;
  LAYER M2 ;
        RECT 9.728 10.828 9.76 10.86 ;
  LAYER M2 ;
        RECT 7.36 10.892 7.392 10.924 ;
  LAYER M2 ;
        RECT 9.728 10.956 9.76 10.988 ;
  LAYER M2 ;
        RECT 7.36 11.02 7.392 11.052 ;
  LAYER M2 ;
        RECT 9.728 11.084 9.76 11.116 ;
  LAYER M2 ;
        RECT 7.36 11.148 7.392 11.18 ;
  LAYER M2 ;
        RECT 9.728 11.212 9.76 11.244 ;
  LAYER M2 ;
        RECT 7.36 11.276 7.392 11.308 ;
  LAYER M2 ;
        RECT 9.728 11.34 9.76 11.372 ;
  LAYER M2 ;
        RECT 7.36 11.404 7.392 11.436 ;
  LAYER M2 ;
        RECT 9.728 11.468 9.76 11.5 ;
  LAYER M2 ;
        RECT 7.36 11.532 7.392 11.564 ;
  LAYER M2 ;
        RECT 9.728 11.596 9.76 11.628 ;
  LAYER M2 ;
        RECT 7.36 11.66 7.392 11.692 ;
  LAYER M2 ;
        RECT 9.728 11.724 9.76 11.756 ;
  LAYER M2 ;
        RECT 7.36 11.788 7.392 11.82 ;
  LAYER M2 ;
        RECT 9.728 11.852 9.76 11.884 ;
  LAYER M2 ;
        RECT 7.36 11.916 7.392 11.948 ;
  LAYER M2 ;
        RECT 9.728 11.98 9.76 12.012 ;
  LAYER M2 ;
        RECT 7.36 12.044 7.392 12.076 ;
  LAYER M2 ;
        RECT 9.728 12.108 9.76 12.14 ;
  LAYER M2 ;
        RECT 7.36 12.172 7.392 12.204 ;
  LAYER M2 ;
        RECT 9.728 12.236 9.76 12.268 ;
  LAYER M2 ;
        RECT 7.36 12.3 7.392 12.332 ;
  LAYER M2 ;
        RECT 9.728 12.364 9.76 12.396 ;
  LAYER M2 ;
        RECT 7.36 12.428 7.392 12.46 ;
  LAYER M2 ;
        RECT 9.728 12.492 9.76 12.524 ;
  LAYER M2 ;
        RECT 7.36 12.556 7.392 12.588 ;
  LAYER M2 ;
        RECT 9.728 12.62 9.76 12.652 ;
  LAYER M2 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M1 ;
        RECT 7.36 13.404 7.392 15.912 ;
  LAYER M3 ;
        RECT 7.36 15.86 7.392 15.892 ;
  LAYER M1 ;
        RECT 7.424 13.404 7.456 15.912 ;
  LAYER M3 ;
        RECT 7.424 13.424 7.456 13.456 ;
  LAYER M1 ;
        RECT 7.488 13.404 7.52 15.912 ;
  LAYER M3 ;
        RECT 7.488 15.86 7.52 15.892 ;
  LAYER M1 ;
        RECT 7.552 13.404 7.584 15.912 ;
  LAYER M3 ;
        RECT 7.552 13.424 7.584 13.456 ;
  LAYER M1 ;
        RECT 7.616 13.404 7.648 15.912 ;
  LAYER M3 ;
        RECT 7.616 15.86 7.648 15.892 ;
  LAYER M1 ;
        RECT 7.68 13.404 7.712 15.912 ;
  LAYER M3 ;
        RECT 7.68 13.424 7.712 13.456 ;
  LAYER M1 ;
        RECT 7.744 13.404 7.776 15.912 ;
  LAYER M3 ;
        RECT 7.744 15.86 7.776 15.892 ;
  LAYER M1 ;
        RECT 7.808 13.404 7.84 15.912 ;
  LAYER M3 ;
        RECT 7.808 13.424 7.84 13.456 ;
  LAYER M1 ;
        RECT 7.872 13.404 7.904 15.912 ;
  LAYER M3 ;
        RECT 7.872 15.86 7.904 15.892 ;
  LAYER M1 ;
        RECT 7.936 13.404 7.968 15.912 ;
  LAYER M3 ;
        RECT 7.936 13.424 7.968 13.456 ;
  LAYER M1 ;
        RECT 8 13.404 8.032 15.912 ;
  LAYER M3 ;
        RECT 8 15.86 8.032 15.892 ;
  LAYER M1 ;
        RECT 8.064 13.404 8.096 15.912 ;
  LAYER M3 ;
        RECT 8.064 13.424 8.096 13.456 ;
  LAYER M1 ;
        RECT 8.128 13.404 8.16 15.912 ;
  LAYER M3 ;
        RECT 8.128 15.86 8.16 15.892 ;
  LAYER M1 ;
        RECT 8.192 13.404 8.224 15.912 ;
  LAYER M3 ;
        RECT 8.192 13.424 8.224 13.456 ;
  LAYER M1 ;
        RECT 8.256 13.404 8.288 15.912 ;
  LAYER M3 ;
        RECT 8.256 15.86 8.288 15.892 ;
  LAYER M1 ;
        RECT 8.32 13.404 8.352 15.912 ;
  LAYER M3 ;
        RECT 8.32 13.424 8.352 13.456 ;
  LAYER M1 ;
        RECT 8.384 13.404 8.416 15.912 ;
  LAYER M3 ;
        RECT 8.384 15.86 8.416 15.892 ;
  LAYER M1 ;
        RECT 8.448 13.404 8.48 15.912 ;
  LAYER M3 ;
        RECT 8.448 13.424 8.48 13.456 ;
  LAYER M1 ;
        RECT 8.512 13.404 8.544 15.912 ;
  LAYER M3 ;
        RECT 8.512 15.86 8.544 15.892 ;
  LAYER M1 ;
        RECT 8.576 13.404 8.608 15.912 ;
  LAYER M3 ;
        RECT 8.576 13.424 8.608 13.456 ;
  LAYER M1 ;
        RECT 8.64 13.404 8.672 15.912 ;
  LAYER M3 ;
        RECT 8.64 15.86 8.672 15.892 ;
  LAYER M1 ;
        RECT 8.704 13.404 8.736 15.912 ;
  LAYER M3 ;
        RECT 8.704 13.424 8.736 13.456 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 15.912 ;
  LAYER M3 ;
        RECT 8.768 15.86 8.8 15.892 ;
  LAYER M1 ;
        RECT 8.832 13.404 8.864 15.912 ;
  LAYER M3 ;
        RECT 8.832 13.424 8.864 13.456 ;
  LAYER M1 ;
        RECT 8.896 13.404 8.928 15.912 ;
  LAYER M3 ;
        RECT 8.896 15.86 8.928 15.892 ;
  LAYER M1 ;
        RECT 8.96 13.404 8.992 15.912 ;
  LAYER M3 ;
        RECT 8.96 13.424 8.992 13.456 ;
  LAYER M1 ;
        RECT 9.024 13.404 9.056 15.912 ;
  LAYER M3 ;
        RECT 9.024 15.86 9.056 15.892 ;
  LAYER M1 ;
        RECT 9.088 13.404 9.12 15.912 ;
  LAYER M3 ;
        RECT 9.088 13.424 9.12 13.456 ;
  LAYER M1 ;
        RECT 9.152 13.404 9.184 15.912 ;
  LAYER M3 ;
        RECT 9.152 15.86 9.184 15.892 ;
  LAYER M1 ;
        RECT 9.216 13.404 9.248 15.912 ;
  LAYER M3 ;
        RECT 9.216 13.424 9.248 13.456 ;
  LAYER M1 ;
        RECT 9.28 13.404 9.312 15.912 ;
  LAYER M3 ;
        RECT 9.28 15.86 9.312 15.892 ;
  LAYER M1 ;
        RECT 9.344 13.404 9.376 15.912 ;
  LAYER M3 ;
        RECT 9.344 13.424 9.376 13.456 ;
  LAYER M1 ;
        RECT 9.408 13.404 9.44 15.912 ;
  LAYER M3 ;
        RECT 9.408 15.86 9.44 15.892 ;
  LAYER M1 ;
        RECT 9.472 13.404 9.504 15.912 ;
  LAYER M3 ;
        RECT 9.472 13.424 9.504 13.456 ;
  LAYER M1 ;
        RECT 9.536 13.404 9.568 15.912 ;
  LAYER M3 ;
        RECT 9.536 15.86 9.568 15.892 ;
  LAYER M1 ;
        RECT 9.6 13.404 9.632 15.912 ;
  LAYER M3 ;
        RECT 9.6 13.424 9.632 13.456 ;
  LAYER M1 ;
        RECT 9.664 13.404 9.696 15.912 ;
  LAYER M3 ;
        RECT 9.664 15.86 9.696 15.892 ;
  LAYER M1 ;
        RECT 9.728 13.404 9.76 15.912 ;
  LAYER M3 ;
        RECT 7.36 13.488 7.392 13.52 ;
  LAYER M2 ;
        RECT 9.728 13.552 9.76 13.584 ;
  LAYER M2 ;
        RECT 7.36 13.616 7.392 13.648 ;
  LAYER M2 ;
        RECT 9.728 13.68 9.76 13.712 ;
  LAYER M2 ;
        RECT 7.36 13.744 7.392 13.776 ;
  LAYER M2 ;
        RECT 9.728 13.808 9.76 13.84 ;
  LAYER M2 ;
        RECT 7.36 13.872 7.392 13.904 ;
  LAYER M2 ;
        RECT 9.728 13.936 9.76 13.968 ;
  LAYER M2 ;
        RECT 7.36 14 7.392 14.032 ;
  LAYER M2 ;
        RECT 9.728 14.064 9.76 14.096 ;
  LAYER M2 ;
        RECT 7.36 14.128 7.392 14.16 ;
  LAYER M2 ;
        RECT 9.728 14.192 9.76 14.224 ;
  LAYER M2 ;
        RECT 7.36 14.256 7.392 14.288 ;
  LAYER M2 ;
        RECT 9.728 14.32 9.76 14.352 ;
  LAYER M2 ;
        RECT 7.36 14.384 7.392 14.416 ;
  LAYER M2 ;
        RECT 9.728 14.448 9.76 14.48 ;
  LAYER M2 ;
        RECT 7.36 14.512 7.392 14.544 ;
  LAYER M2 ;
        RECT 9.728 14.576 9.76 14.608 ;
  LAYER M2 ;
        RECT 7.36 14.64 7.392 14.672 ;
  LAYER M2 ;
        RECT 9.728 14.704 9.76 14.736 ;
  LAYER M2 ;
        RECT 7.36 14.768 7.392 14.8 ;
  LAYER M2 ;
        RECT 9.728 14.832 9.76 14.864 ;
  LAYER M2 ;
        RECT 7.36 14.896 7.392 14.928 ;
  LAYER M2 ;
        RECT 9.728 14.96 9.76 14.992 ;
  LAYER M2 ;
        RECT 7.36 15.024 7.392 15.056 ;
  LAYER M2 ;
        RECT 9.728 15.088 9.76 15.12 ;
  LAYER M2 ;
        RECT 7.36 15.152 7.392 15.184 ;
  LAYER M2 ;
        RECT 9.728 15.216 9.76 15.248 ;
  LAYER M2 ;
        RECT 7.36 15.28 7.392 15.312 ;
  LAYER M2 ;
        RECT 9.728 15.344 9.76 15.376 ;
  LAYER M2 ;
        RECT 7.36 15.408 7.392 15.44 ;
  LAYER M2 ;
        RECT 9.728 15.472 9.76 15.504 ;
  LAYER M2 ;
        RECT 7.36 15.536 7.392 15.568 ;
  LAYER M2 ;
        RECT 9.728 15.6 9.76 15.632 ;
  LAYER M2 ;
        RECT 7.36 15.664 7.392 15.696 ;
  LAYER M2 ;
        RECT 9.728 15.728 9.76 15.76 ;
  LAYER M2 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M1 ;
        RECT 7.36 16.512 7.392 19.02 ;
  LAYER M3 ;
        RECT 7.36 18.968 7.392 19 ;
  LAYER M1 ;
        RECT 7.424 16.512 7.456 19.02 ;
  LAYER M3 ;
        RECT 7.424 16.532 7.456 16.564 ;
  LAYER M1 ;
        RECT 7.488 16.512 7.52 19.02 ;
  LAYER M3 ;
        RECT 7.488 18.968 7.52 19 ;
  LAYER M1 ;
        RECT 7.552 16.512 7.584 19.02 ;
  LAYER M3 ;
        RECT 7.552 16.532 7.584 16.564 ;
  LAYER M1 ;
        RECT 7.616 16.512 7.648 19.02 ;
  LAYER M3 ;
        RECT 7.616 18.968 7.648 19 ;
  LAYER M1 ;
        RECT 7.68 16.512 7.712 19.02 ;
  LAYER M3 ;
        RECT 7.68 16.532 7.712 16.564 ;
  LAYER M1 ;
        RECT 7.744 16.512 7.776 19.02 ;
  LAYER M3 ;
        RECT 7.744 18.968 7.776 19 ;
  LAYER M1 ;
        RECT 7.808 16.512 7.84 19.02 ;
  LAYER M3 ;
        RECT 7.808 16.532 7.84 16.564 ;
  LAYER M1 ;
        RECT 7.872 16.512 7.904 19.02 ;
  LAYER M3 ;
        RECT 7.872 18.968 7.904 19 ;
  LAYER M1 ;
        RECT 7.936 16.512 7.968 19.02 ;
  LAYER M3 ;
        RECT 7.936 16.532 7.968 16.564 ;
  LAYER M1 ;
        RECT 8 16.512 8.032 19.02 ;
  LAYER M3 ;
        RECT 8 18.968 8.032 19 ;
  LAYER M1 ;
        RECT 8.064 16.512 8.096 19.02 ;
  LAYER M3 ;
        RECT 8.064 16.532 8.096 16.564 ;
  LAYER M1 ;
        RECT 8.128 16.512 8.16 19.02 ;
  LAYER M3 ;
        RECT 8.128 18.968 8.16 19 ;
  LAYER M1 ;
        RECT 8.192 16.512 8.224 19.02 ;
  LAYER M3 ;
        RECT 8.192 16.532 8.224 16.564 ;
  LAYER M1 ;
        RECT 8.256 16.512 8.288 19.02 ;
  LAYER M3 ;
        RECT 8.256 18.968 8.288 19 ;
  LAYER M1 ;
        RECT 8.32 16.512 8.352 19.02 ;
  LAYER M3 ;
        RECT 8.32 16.532 8.352 16.564 ;
  LAYER M1 ;
        RECT 8.384 16.512 8.416 19.02 ;
  LAYER M3 ;
        RECT 8.384 18.968 8.416 19 ;
  LAYER M1 ;
        RECT 8.448 16.512 8.48 19.02 ;
  LAYER M3 ;
        RECT 8.448 16.532 8.48 16.564 ;
  LAYER M1 ;
        RECT 8.512 16.512 8.544 19.02 ;
  LAYER M3 ;
        RECT 8.512 18.968 8.544 19 ;
  LAYER M1 ;
        RECT 8.576 16.512 8.608 19.02 ;
  LAYER M3 ;
        RECT 8.576 16.532 8.608 16.564 ;
  LAYER M1 ;
        RECT 8.64 16.512 8.672 19.02 ;
  LAYER M3 ;
        RECT 8.64 18.968 8.672 19 ;
  LAYER M1 ;
        RECT 8.704 16.512 8.736 19.02 ;
  LAYER M3 ;
        RECT 8.704 16.532 8.736 16.564 ;
  LAYER M1 ;
        RECT 8.768 16.512 8.8 19.02 ;
  LAYER M3 ;
        RECT 8.768 18.968 8.8 19 ;
  LAYER M1 ;
        RECT 8.832 16.512 8.864 19.02 ;
  LAYER M3 ;
        RECT 8.832 16.532 8.864 16.564 ;
  LAYER M1 ;
        RECT 8.896 16.512 8.928 19.02 ;
  LAYER M3 ;
        RECT 8.896 18.968 8.928 19 ;
  LAYER M1 ;
        RECT 8.96 16.512 8.992 19.02 ;
  LAYER M3 ;
        RECT 8.96 16.532 8.992 16.564 ;
  LAYER M1 ;
        RECT 9.024 16.512 9.056 19.02 ;
  LAYER M3 ;
        RECT 9.024 18.968 9.056 19 ;
  LAYER M1 ;
        RECT 9.088 16.512 9.12 19.02 ;
  LAYER M3 ;
        RECT 9.088 16.532 9.12 16.564 ;
  LAYER M1 ;
        RECT 9.152 16.512 9.184 19.02 ;
  LAYER M3 ;
        RECT 9.152 18.968 9.184 19 ;
  LAYER M1 ;
        RECT 9.216 16.512 9.248 19.02 ;
  LAYER M3 ;
        RECT 9.216 16.532 9.248 16.564 ;
  LAYER M1 ;
        RECT 9.28 16.512 9.312 19.02 ;
  LAYER M3 ;
        RECT 9.28 18.968 9.312 19 ;
  LAYER M1 ;
        RECT 9.344 16.512 9.376 19.02 ;
  LAYER M3 ;
        RECT 9.344 16.532 9.376 16.564 ;
  LAYER M1 ;
        RECT 9.408 16.512 9.44 19.02 ;
  LAYER M3 ;
        RECT 9.408 18.968 9.44 19 ;
  LAYER M1 ;
        RECT 9.472 16.512 9.504 19.02 ;
  LAYER M3 ;
        RECT 9.472 16.532 9.504 16.564 ;
  LAYER M1 ;
        RECT 9.536 16.512 9.568 19.02 ;
  LAYER M3 ;
        RECT 9.536 18.968 9.568 19 ;
  LAYER M1 ;
        RECT 9.6 16.512 9.632 19.02 ;
  LAYER M3 ;
        RECT 9.6 16.532 9.632 16.564 ;
  LAYER M1 ;
        RECT 9.664 16.512 9.696 19.02 ;
  LAYER M3 ;
        RECT 9.664 18.968 9.696 19 ;
  LAYER M1 ;
        RECT 9.728 16.512 9.76 19.02 ;
  LAYER M3 ;
        RECT 7.36 16.596 7.392 16.628 ;
  LAYER M2 ;
        RECT 9.728 16.66 9.76 16.692 ;
  LAYER M2 ;
        RECT 7.36 16.724 7.392 16.756 ;
  LAYER M2 ;
        RECT 9.728 16.788 9.76 16.82 ;
  LAYER M2 ;
        RECT 7.36 16.852 7.392 16.884 ;
  LAYER M2 ;
        RECT 9.728 16.916 9.76 16.948 ;
  LAYER M2 ;
        RECT 7.36 16.98 7.392 17.012 ;
  LAYER M2 ;
        RECT 9.728 17.044 9.76 17.076 ;
  LAYER M2 ;
        RECT 7.36 17.108 7.392 17.14 ;
  LAYER M2 ;
        RECT 9.728 17.172 9.76 17.204 ;
  LAYER M2 ;
        RECT 7.36 17.236 7.392 17.268 ;
  LAYER M2 ;
        RECT 9.728 17.3 9.76 17.332 ;
  LAYER M2 ;
        RECT 7.36 17.364 7.392 17.396 ;
  LAYER M2 ;
        RECT 9.728 17.428 9.76 17.46 ;
  LAYER M2 ;
        RECT 7.36 17.492 7.392 17.524 ;
  LAYER M2 ;
        RECT 9.728 17.556 9.76 17.588 ;
  LAYER M2 ;
        RECT 7.36 17.62 7.392 17.652 ;
  LAYER M2 ;
        RECT 9.728 17.684 9.76 17.716 ;
  LAYER M2 ;
        RECT 7.36 17.748 7.392 17.78 ;
  LAYER M2 ;
        RECT 9.728 17.812 9.76 17.844 ;
  LAYER M2 ;
        RECT 7.36 17.876 7.392 17.908 ;
  LAYER M2 ;
        RECT 9.728 17.94 9.76 17.972 ;
  LAYER M2 ;
        RECT 7.36 18.004 7.392 18.036 ;
  LAYER M2 ;
        RECT 9.728 18.068 9.76 18.1 ;
  LAYER M2 ;
        RECT 7.36 18.132 7.392 18.164 ;
  LAYER M2 ;
        RECT 9.728 18.196 9.76 18.228 ;
  LAYER M2 ;
        RECT 7.36 18.26 7.392 18.292 ;
  LAYER M2 ;
        RECT 9.728 18.324 9.76 18.356 ;
  LAYER M2 ;
        RECT 7.36 18.388 7.392 18.42 ;
  LAYER M2 ;
        RECT 9.728 18.452 9.76 18.484 ;
  LAYER M2 ;
        RECT 7.36 18.516 7.392 18.548 ;
  LAYER M2 ;
        RECT 9.728 18.58 9.76 18.612 ;
  LAYER M2 ;
        RECT 7.36 18.644 7.392 18.676 ;
  LAYER M2 ;
        RECT 9.728 18.708 9.76 18.74 ;
  LAYER M2 ;
        RECT 7.36 18.772 7.392 18.804 ;
  LAYER M2 ;
        RECT 9.728 18.836 9.76 18.868 ;
  LAYER M2 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M1 ;
        RECT 7.36 19.62 7.392 22.128 ;
  LAYER M3 ;
        RECT 7.36 22.076 7.392 22.108 ;
  LAYER M1 ;
        RECT 7.424 19.62 7.456 22.128 ;
  LAYER M3 ;
        RECT 7.424 19.64 7.456 19.672 ;
  LAYER M1 ;
        RECT 7.488 19.62 7.52 22.128 ;
  LAYER M3 ;
        RECT 7.488 22.076 7.52 22.108 ;
  LAYER M1 ;
        RECT 7.552 19.62 7.584 22.128 ;
  LAYER M3 ;
        RECT 7.552 19.64 7.584 19.672 ;
  LAYER M1 ;
        RECT 7.616 19.62 7.648 22.128 ;
  LAYER M3 ;
        RECT 7.616 22.076 7.648 22.108 ;
  LAYER M1 ;
        RECT 7.68 19.62 7.712 22.128 ;
  LAYER M3 ;
        RECT 7.68 19.64 7.712 19.672 ;
  LAYER M1 ;
        RECT 7.744 19.62 7.776 22.128 ;
  LAYER M3 ;
        RECT 7.744 22.076 7.776 22.108 ;
  LAYER M1 ;
        RECT 7.808 19.62 7.84 22.128 ;
  LAYER M3 ;
        RECT 7.808 19.64 7.84 19.672 ;
  LAYER M1 ;
        RECT 7.872 19.62 7.904 22.128 ;
  LAYER M3 ;
        RECT 7.872 22.076 7.904 22.108 ;
  LAYER M1 ;
        RECT 7.936 19.62 7.968 22.128 ;
  LAYER M3 ;
        RECT 7.936 19.64 7.968 19.672 ;
  LAYER M1 ;
        RECT 8 19.62 8.032 22.128 ;
  LAYER M3 ;
        RECT 8 22.076 8.032 22.108 ;
  LAYER M1 ;
        RECT 8.064 19.62 8.096 22.128 ;
  LAYER M3 ;
        RECT 8.064 19.64 8.096 19.672 ;
  LAYER M1 ;
        RECT 8.128 19.62 8.16 22.128 ;
  LAYER M3 ;
        RECT 8.128 22.076 8.16 22.108 ;
  LAYER M1 ;
        RECT 8.192 19.62 8.224 22.128 ;
  LAYER M3 ;
        RECT 8.192 19.64 8.224 19.672 ;
  LAYER M1 ;
        RECT 8.256 19.62 8.288 22.128 ;
  LAYER M3 ;
        RECT 8.256 22.076 8.288 22.108 ;
  LAYER M1 ;
        RECT 8.32 19.62 8.352 22.128 ;
  LAYER M3 ;
        RECT 8.32 19.64 8.352 19.672 ;
  LAYER M1 ;
        RECT 8.384 19.62 8.416 22.128 ;
  LAYER M3 ;
        RECT 8.384 22.076 8.416 22.108 ;
  LAYER M1 ;
        RECT 8.448 19.62 8.48 22.128 ;
  LAYER M3 ;
        RECT 8.448 19.64 8.48 19.672 ;
  LAYER M1 ;
        RECT 8.512 19.62 8.544 22.128 ;
  LAYER M3 ;
        RECT 8.512 22.076 8.544 22.108 ;
  LAYER M1 ;
        RECT 8.576 19.62 8.608 22.128 ;
  LAYER M3 ;
        RECT 8.576 19.64 8.608 19.672 ;
  LAYER M1 ;
        RECT 8.64 19.62 8.672 22.128 ;
  LAYER M3 ;
        RECT 8.64 22.076 8.672 22.108 ;
  LAYER M1 ;
        RECT 8.704 19.62 8.736 22.128 ;
  LAYER M3 ;
        RECT 8.704 19.64 8.736 19.672 ;
  LAYER M1 ;
        RECT 8.768 19.62 8.8 22.128 ;
  LAYER M3 ;
        RECT 8.768 22.076 8.8 22.108 ;
  LAYER M1 ;
        RECT 8.832 19.62 8.864 22.128 ;
  LAYER M3 ;
        RECT 8.832 19.64 8.864 19.672 ;
  LAYER M1 ;
        RECT 8.896 19.62 8.928 22.128 ;
  LAYER M3 ;
        RECT 8.896 22.076 8.928 22.108 ;
  LAYER M1 ;
        RECT 8.96 19.62 8.992 22.128 ;
  LAYER M3 ;
        RECT 8.96 19.64 8.992 19.672 ;
  LAYER M1 ;
        RECT 9.024 19.62 9.056 22.128 ;
  LAYER M3 ;
        RECT 9.024 22.076 9.056 22.108 ;
  LAYER M1 ;
        RECT 9.088 19.62 9.12 22.128 ;
  LAYER M3 ;
        RECT 9.088 19.64 9.12 19.672 ;
  LAYER M1 ;
        RECT 9.152 19.62 9.184 22.128 ;
  LAYER M3 ;
        RECT 9.152 22.076 9.184 22.108 ;
  LAYER M1 ;
        RECT 9.216 19.62 9.248 22.128 ;
  LAYER M3 ;
        RECT 9.216 19.64 9.248 19.672 ;
  LAYER M1 ;
        RECT 9.28 19.62 9.312 22.128 ;
  LAYER M3 ;
        RECT 9.28 22.076 9.312 22.108 ;
  LAYER M1 ;
        RECT 9.344 19.62 9.376 22.128 ;
  LAYER M3 ;
        RECT 9.344 19.64 9.376 19.672 ;
  LAYER M1 ;
        RECT 9.408 19.62 9.44 22.128 ;
  LAYER M3 ;
        RECT 9.408 22.076 9.44 22.108 ;
  LAYER M1 ;
        RECT 9.472 19.62 9.504 22.128 ;
  LAYER M3 ;
        RECT 9.472 19.64 9.504 19.672 ;
  LAYER M1 ;
        RECT 9.536 19.62 9.568 22.128 ;
  LAYER M3 ;
        RECT 9.536 22.076 9.568 22.108 ;
  LAYER M1 ;
        RECT 9.6 19.62 9.632 22.128 ;
  LAYER M3 ;
        RECT 9.6 19.64 9.632 19.672 ;
  LAYER M1 ;
        RECT 9.664 19.62 9.696 22.128 ;
  LAYER M3 ;
        RECT 9.664 22.076 9.696 22.108 ;
  LAYER M1 ;
        RECT 9.728 19.62 9.76 22.128 ;
  LAYER M3 ;
        RECT 7.36 19.704 7.392 19.736 ;
  LAYER M2 ;
        RECT 9.728 19.768 9.76 19.8 ;
  LAYER M2 ;
        RECT 7.36 19.832 7.392 19.864 ;
  LAYER M2 ;
        RECT 9.728 19.896 9.76 19.928 ;
  LAYER M2 ;
        RECT 7.36 19.96 7.392 19.992 ;
  LAYER M2 ;
        RECT 9.728 20.024 9.76 20.056 ;
  LAYER M2 ;
        RECT 7.36 20.088 7.392 20.12 ;
  LAYER M2 ;
        RECT 9.728 20.152 9.76 20.184 ;
  LAYER M2 ;
        RECT 7.36 20.216 7.392 20.248 ;
  LAYER M2 ;
        RECT 9.728 20.28 9.76 20.312 ;
  LAYER M2 ;
        RECT 7.36 20.344 7.392 20.376 ;
  LAYER M2 ;
        RECT 9.728 20.408 9.76 20.44 ;
  LAYER M2 ;
        RECT 7.36 20.472 7.392 20.504 ;
  LAYER M2 ;
        RECT 9.728 20.536 9.76 20.568 ;
  LAYER M2 ;
        RECT 7.36 20.6 7.392 20.632 ;
  LAYER M2 ;
        RECT 9.728 20.664 9.76 20.696 ;
  LAYER M2 ;
        RECT 7.36 20.728 7.392 20.76 ;
  LAYER M2 ;
        RECT 9.728 20.792 9.76 20.824 ;
  LAYER M2 ;
        RECT 7.36 20.856 7.392 20.888 ;
  LAYER M2 ;
        RECT 9.728 20.92 9.76 20.952 ;
  LAYER M2 ;
        RECT 7.36 20.984 7.392 21.016 ;
  LAYER M2 ;
        RECT 9.728 21.048 9.76 21.08 ;
  LAYER M2 ;
        RECT 7.36 21.112 7.392 21.144 ;
  LAYER M2 ;
        RECT 9.728 21.176 9.76 21.208 ;
  LAYER M2 ;
        RECT 7.36 21.24 7.392 21.272 ;
  LAYER M2 ;
        RECT 9.728 21.304 9.76 21.336 ;
  LAYER M2 ;
        RECT 7.36 21.368 7.392 21.4 ;
  LAYER M2 ;
        RECT 9.728 21.432 9.76 21.464 ;
  LAYER M2 ;
        RECT 7.36 21.496 7.392 21.528 ;
  LAYER M2 ;
        RECT 9.728 21.56 9.76 21.592 ;
  LAYER M2 ;
        RECT 7.36 21.624 7.392 21.656 ;
  LAYER M2 ;
        RECT 9.728 21.688 9.76 21.72 ;
  LAYER M2 ;
        RECT 7.36 21.752 7.392 21.784 ;
  LAYER M2 ;
        RECT 9.728 21.816 9.76 21.848 ;
  LAYER M2 ;
        RECT 7.36 21.88 7.392 21.912 ;
  LAYER M2 ;
        RECT 9.728 21.944 9.76 21.976 ;
  LAYER M2 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M1 ;
        RECT 7.36 22.728 7.392 25.236 ;
  LAYER M3 ;
        RECT 7.36 25.184 7.392 25.216 ;
  LAYER M1 ;
        RECT 7.424 22.728 7.456 25.236 ;
  LAYER M3 ;
        RECT 7.424 22.748 7.456 22.78 ;
  LAYER M1 ;
        RECT 7.488 22.728 7.52 25.236 ;
  LAYER M3 ;
        RECT 7.488 25.184 7.52 25.216 ;
  LAYER M1 ;
        RECT 7.552 22.728 7.584 25.236 ;
  LAYER M3 ;
        RECT 7.552 22.748 7.584 22.78 ;
  LAYER M1 ;
        RECT 7.616 22.728 7.648 25.236 ;
  LAYER M3 ;
        RECT 7.616 25.184 7.648 25.216 ;
  LAYER M1 ;
        RECT 7.68 22.728 7.712 25.236 ;
  LAYER M3 ;
        RECT 7.68 22.748 7.712 22.78 ;
  LAYER M1 ;
        RECT 7.744 22.728 7.776 25.236 ;
  LAYER M3 ;
        RECT 7.744 25.184 7.776 25.216 ;
  LAYER M1 ;
        RECT 7.808 22.728 7.84 25.236 ;
  LAYER M3 ;
        RECT 7.808 22.748 7.84 22.78 ;
  LAYER M1 ;
        RECT 7.872 22.728 7.904 25.236 ;
  LAYER M3 ;
        RECT 7.872 25.184 7.904 25.216 ;
  LAYER M1 ;
        RECT 7.936 22.728 7.968 25.236 ;
  LAYER M3 ;
        RECT 7.936 22.748 7.968 22.78 ;
  LAYER M1 ;
        RECT 8 22.728 8.032 25.236 ;
  LAYER M3 ;
        RECT 8 25.184 8.032 25.216 ;
  LAYER M1 ;
        RECT 8.064 22.728 8.096 25.236 ;
  LAYER M3 ;
        RECT 8.064 22.748 8.096 22.78 ;
  LAYER M1 ;
        RECT 8.128 22.728 8.16 25.236 ;
  LAYER M3 ;
        RECT 8.128 25.184 8.16 25.216 ;
  LAYER M1 ;
        RECT 8.192 22.728 8.224 25.236 ;
  LAYER M3 ;
        RECT 8.192 22.748 8.224 22.78 ;
  LAYER M1 ;
        RECT 8.256 22.728 8.288 25.236 ;
  LAYER M3 ;
        RECT 8.256 25.184 8.288 25.216 ;
  LAYER M1 ;
        RECT 8.32 22.728 8.352 25.236 ;
  LAYER M3 ;
        RECT 8.32 22.748 8.352 22.78 ;
  LAYER M1 ;
        RECT 8.384 22.728 8.416 25.236 ;
  LAYER M3 ;
        RECT 8.384 25.184 8.416 25.216 ;
  LAYER M1 ;
        RECT 8.448 22.728 8.48 25.236 ;
  LAYER M3 ;
        RECT 8.448 22.748 8.48 22.78 ;
  LAYER M1 ;
        RECT 8.512 22.728 8.544 25.236 ;
  LAYER M3 ;
        RECT 8.512 25.184 8.544 25.216 ;
  LAYER M1 ;
        RECT 8.576 22.728 8.608 25.236 ;
  LAYER M3 ;
        RECT 8.576 22.748 8.608 22.78 ;
  LAYER M1 ;
        RECT 8.64 22.728 8.672 25.236 ;
  LAYER M3 ;
        RECT 8.64 25.184 8.672 25.216 ;
  LAYER M1 ;
        RECT 8.704 22.728 8.736 25.236 ;
  LAYER M3 ;
        RECT 8.704 22.748 8.736 22.78 ;
  LAYER M1 ;
        RECT 8.768 22.728 8.8 25.236 ;
  LAYER M3 ;
        RECT 8.768 25.184 8.8 25.216 ;
  LAYER M1 ;
        RECT 8.832 22.728 8.864 25.236 ;
  LAYER M3 ;
        RECT 8.832 22.748 8.864 22.78 ;
  LAYER M1 ;
        RECT 8.896 22.728 8.928 25.236 ;
  LAYER M3 ;
        RECT 8.896 25.184 8.928 25.216 ;
  LAYER M1 ;
        RECT 8.96 22.728 8.992 25.236 ;
  LAYER M3 ;
        RECT 8.96 22.748 8.992 22.78 ;
  LAYER M1 ;
        RECT 9.024 22.728 9.056 25.236 ;
  LAYER M3 ;
        RECT 9.024 25.184 9.056 25.216 ;
  LAYER M1 ;
        RECT 9.088 22.728 9.12 25.236 ;
  LAYER M3 ;
        RECT 9.088 22.748 9.12 22.78 ;
  LAYER M1 ;
        RECT 9.152 22.728 9.184 25.236 ;
  LAYER M3 ;
        RECT 9.152 25.184 9.184 25.216 ;
  LAYER M1 ;
        RECT 9.216 22.728 9.248 25.236 ;
  LAYER M3 ;
        RECT 9.216 22.748 9.248 22.78 ;
  LAYER M1 ;
        RECT 9.28 22.728 9.312 25.236 ;
  LAYER M3 ;
        RECT 9.28 25.184 9.312 25.216 ;
  LAYER M1 ;
        RECT 9.344 22.728 9.376 25.236 ;
  LAYER M3 ;
        RECT 9.344 22.748 9.376 22.78 ;
  LAYER M1 ;
        RECT 9.408 22.728 9.44 25.236 ;
  LAYER M3 ;
        RECT 9.408 25.184 9.44 25.216 ;
  LAYER M1 ;
        RECT 9.472 22.728 9.504 25.236 ;
  LAYER M3 ;
        RECT 9.472 22.748 9.504 22.78 ;
  LAYER M1 ;
        RECT 9.536 22.728 9.568 25.236 ;
  LAYER M3 ;
        RECT 9.536 25.184 9.568 25.216 ;
  LAYER M1 ;
        RECT 9.6 22.728 9.632 25.236 ;
  LAYER M3 ;
        RECT 9.6 22.748 9.632 22.78 ;
  LAYER M1 ;
        RECT 9.664 22.728 9.696 25.236 ;
  LAYER M3 ;
        RECT 9.664 25.184 9.696 25.216 ;
  LAYER M1 ;
        RECT 9.728 22.728 9.76 25.236 ;
  LAYER M3 ;
        RECT 7.36 22.812 7.392 22.844 ;
  LAYER M2 ;
        RECT 9.728 22.876 9.76 22.908 ;
  LAYER M2 ;
        RECT 7.36 22.94 7.392 22.972 ;
  LAYER M2 ;
        RECT 9.728 23.004 9.76 23.036 ;
  LAYER M2 ;
        RECT 7.36 23.068 7.392 23.1 ;
  LAYER M2 ;
        RECT 9.728 23.132 9.76 23.164 ;
  LAYER M2 ;
        RECT 7.36 23.196 7.392 23.228 ;
  LAYER M2 ;
        RECT 9.728 23.26 9.76 23.292 ;
  LAYER M2 ;
        RECT 7.36 23.324 7.392 23.356 ;
  LAYER M2 ;
        RECT 9.728 23.388 9.76 23.42 ;
  LAYER M2 ;
        RECT 7.36 23.452 7.392 23.484 ;
  LAYER M2 ;
        RECT 9.728 23.516 9.76 23.548 ;
  LAYER M2 ;
        RECT 7.36 23.58 7.392 23.612 ;
  LAYER M2 ;
        RECT 9.728 23.644 9.76 23.676 ;
  LAYER M2 ;
        RECT 7.36 23.708 7.392 23.74 ;
  LAYER M2 ;
        RECT 9.728 23.772 9.76 23.804 ;
  LAYER M2 ;
        RECT 7.36 23.836 7.392 23.868 ;
  LAYER M2 ;
        RECT 9.728 23.9 9.76 23.932 ;
  LAYER M2 ;
        RECT 7.36 23.964 7.392 23.996 ;
  LAYER M2 ;
        RECT 9.728 24.028 9.76 24.06 ;
  LAYER M2 ;
        RECT 7.36 24.092 7.392 24.124 ;
  LAYER M2 ;
        RECT 9.728 24.156 9.76 24.188 ;
  LAYER M2 ;
        RECT 7.36 24.22 7.392 24.252 ;
  LAYER M2 ;
        RECT 9.728 24.284 9.76 24.316 ;
  LAYER M2 ;
        RECT 7.36 24.348 7.392 24.38 ;
  LAYER M2 ;
        RECT 9.728 24.412 9.76 24.444 ;
  LAYER M2 ;
        RECT 7.36 24.476 7.392 24.508 ;
  LAYER M2 ;
        RECT 9.728 24.54 9.76 24.572 ;
  LAYER M2 ;
        RECT 7.36 24.604 7.392 24.636 ;
  LAYER M2 ;
        RECT 9.728 24.668 9.76 24.7 ;
  LAYER M2 ;
        RECT 7.36 24.732 7.392 24.764 ;
  LAYER M2 ;
        RECT 9.728 24.796 9.76 24.828 ;
  LAYER M2 ;
        RECT 7.36 24.86 7.392 24.892 ;
  LAYER M2 ;
        RECT 9.728 24.924 9.76 24.956 ;
  LAYER M2 ;
        RECT 7.36 24.988 7.392 25.02 ;
  LAYER M2 ;
        RECT 9.728 25.052 9.76 25.084 ;
  LAYER M2 ;
        RECT 7.312 22.68 9.808 25.284 ;
  END 
END Cap_30fF_Cap_30fF
