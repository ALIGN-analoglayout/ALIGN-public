VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DL1_NMOS_25_1x10
  ORIGIN 0 0 ;
  FOREIGN DL1_NMOS_25_1x10 0 0 ;
  SIZE 2.16 BY 0.402 ;
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.32 2.012 0.338 ;
    END
  END S2
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 2.16 0.018 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 2.16 0.402 ;
    END
  END VDD
  PIN G
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 2.066 0.082 ;
    END
  END G
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 1.904 0.146 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.192 2.12 0.21 ;
    END
  END D2
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 1.796 0.274 ;
    END
  END S1
  OBS
    LAYER M1 ;
      RECT 0 0 2.16 0.402 ;
  END
END DL1_NMOS_25_1x10

MACRO DL2_PMOS_10_1x4
  ORIGIN 0 0 ;
  FOREIGN DL2_PMOS_10_1x4 0 0 ;
  SIZE 0.864 BY 0.402 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.32 0.716 0.338 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.864 0.402 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
    END
  END VSS
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 0.77 0.082 ;
    END
  END G
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 0.824 0.146 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.192 0.608 0.21 ;
    END
  END D2
  OBS
    LAYER M1 ;
      RECT 0 0 0.864 0.402 ;
  END
END DL2_PMOS_10_1x4

MACRO DL1_PMOS_15_1x6
  ORIGIN 0 0 ;
  FOREIGN DL1_PMOS_15_1x6 0 0 ;
  SIZE 1.296 BY 0.402 ;
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.32 1.148 0.338 ;
    END
  END S2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 1.296 0.402 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
    END
  END VSS
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 1.202 0.082 ;
    END
  END G
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 1.04 0.146 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.192 1.256 0.21 ;
    END
  END D2
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 0.932 0.274 ;
    END
  END S1
  OBS
    LAYER M1 ;
      RECT 0 0 1.296 0.402 ;
  END
END DL1_PMOS_15_1x6

MACRO Cap_32f_1x1
  ORIGIN 0 0 ;
  FOREIGN Cap_32f_1x1 0 0 ;
  SIZE 4.024 BY 4.06 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.037 4.024 4.055 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 4.024 0.023 ;
    END
  END MINUS
END Cap_32f_1x1

MACRO Cap_50f_2x3
  ORIGIN 0 0 ;
  FOREIGN Cap_50f_2x3 0 0 ;
  SIZE 7.048 BY 4.7 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.677 4.672 4.695 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 7.048 0.023 ;
    END
  END MINUS
END Cap_50f_2x3

MACRO Cap_60f_2x3
  ORIGIN 0 0 ;
  FOREIGN Cap_60f_2x3 0 0 ;
  SIZE 7.048 BY 4.7 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.677 7.048 4.695 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 7.048 0.023 ;
    END
  END MINUS
END Cap_60f_2x3

MACRO DP_NMOS_75_3x10
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_75_3x10 0 0 ;
  SIZE 2.16 BY 1.298 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 1.152 2.012 1.17 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.148 0.576 2.12 0.594 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 2.012 0.274 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.896 2.16 0.914 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 0.832 2.16 0.85 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 0 2.16 0.018 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 1.28 2.16 1.298 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 0.448 2.16 0.466 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 0.384 2.16 0.402 ;
    END
  END VDD
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 1.024 1.904 1.042 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.256 0.704 2.012 0.722 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 1.904 0.146 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 1.088 2.12 1.106 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.04 0.64 1.796 0.658 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.364 0.192 2.12 0.21 ;
    END
  END D2
  PIN G1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.96 1.85 0.978 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.31 0.768 2.066 0.786 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 1.85 0.082 ;
    END
  END G1
  PIN G2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.31 1.216 2.066 1.234 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.094 0.512 1.85 0.53 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.31 0.32 2.066 0.338 ;
    END
  END G2
  OBS
    LAYER M1 ;
      RECT 0 0 2.16 0.402 ;
      RECT 0 0.402 2.16 0.85 ;
      RECT 0 0.85 2.16 1.298 ;
  END
END DP_NMOS_75_3x10

MACRO DiodeConnected_NMOS_5_1x1
  ORIGIN 0 0 ;
  FOREIGN DiodeConnected_NMOS_5_1x1 0 0 ;
  SIZE 0.216 BY 0.402 ;
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.216 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 0.176 0.082 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.068 0.146 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.216 0.402 ;
    END
  END VDD
END DiodeConnected_NMOS_5_1x1

MACRO DiodeConnected_PMOS_10_1x2
  ORIGIN 0 0 ;
  FOREIGN DiodeConnected_PMOS_10_1x2 0 0 ;
  SIZE 0.432 BY 0.402 ;
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 0.392 0.082 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.284 0.146 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.432 0.402 ;
    END
  END VDD
END DiodeConnected_PMOS_10_1x2

MACRO DiodeConnected_PMOS_20_1x4
  ORIGIN 0 0 ;
  FOREIGN DiodeConnected_PMOS_20_1x4 0 0 ;
  SIZE 0.864 BY 0.402 ;
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 0.824 0.082 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.716 0.146 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.864 0.402 ;
    END
  END VDD
END DiodeConnected_PMOS_20_1x4

MACRO SCM_NMOS_50_1x12
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_50_1x12 0 0 ;
  SIZE 2.592 BY 0.402 ;
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.228 0.192 1.472 0.21 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.444 0.192 1.472 0.21 ;
    END
  END D1
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 2.592 0.018 ;
    END
  END VSS
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 2.444 0.274 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 2.592 0.402 ;
    END
  END VDD
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 2.552 0.146 ;
    END
  END D2
  OBS
    LAYER M1 ;
      RECT 0 0 2.592 0.402 ;
  END
END SCM_NMOS_50_1x12

MACRO Switch_NMOS_10_1x1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_10_1x1 0 0 ;
  SIZE 0.432 BY 0.402 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.064 0.284 0.082 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.192 0.392 0.21 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.128 0.338 0.146 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.432 0.402 ;
    END
  END VDD
END Switch_NMOS_10_1x1

MACRO Switch_PMOS_10_1x1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_10_1x1 0 0 ;
  SIZE 0.432 BY 0.402 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.192 0.284 0.21 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.064 0.392 0.082 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.128 0.338 0.146 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.432 0.402 ;
    END
  END VDD
END Switch_PMOS_10_1x1

END LIBRARY
