.subckt powertrain vcc vg vout
mmp0 vout vg vcc vcc plplvt w=180n l=40n nfin=4 nf=8 m=20
.ends
