MACRO CMC_PMOS_S_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.3000 0.6600 0.7080 ;
      LAYER M3 ;
        RECT 0.9400 0.3000 0.9800 0.7080 ;
    END
  END G
  OBS
    LAYER M3 ;
      RECT 0.3800 0.0480 0.4200 0.4560 ;
    LAYER M3 ;
      RECT 0.7000 0.0480 0.7400 0.4560 ;
    LAYER M3 ;
      RECT 0.4600 0.1320 0.5000 0.5400 ;
    LAYER M3 ;
      RECT 0.7800 0.1320 0.8200 0.5400 ;
    LAYER M3 ;
      RECT 0.5400 0.2160 0.5800 0.6240 ;
    LAYER M3 ;
      RECT 0.8600 0.2160 0.9000 0.6240 ;
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 0.9160 0.4360 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.8360 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4880 0.8360 0.5200 ;
    LAYER M2 ;
      RECT 0.5240 0.2360 1.0760 0.2680 ;
    LAYER M2 ;
      RECT 0.5240 0.5720 1.0760 0.6040 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 0.9960 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.6560 0.9960 0.6880 ;
    LAYER pc ;
      RECT 0.2710 0.0680 0.3690 0.1000 ;
    LAYER pc ;
      RECT 0.9110 0.0680 1.0090 0.1000 ;
  END
END CMC_PMOS_S_n12_X1_Y1
