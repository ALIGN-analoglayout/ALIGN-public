MACRO DCL_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X1_Y1 0 0 ;
  SIZE 0.432 BY 0.648 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.153 0.094 0.171 0.446 ;
    END
  END S
  PIN BG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 0.585 0.432 0.603 ;
    END
  END BG
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.207 0.094 0.225 0.446 ;
    END
  END D
  OBS
    LAYER M2 ;
      RECT 0.094 0.261 0.392 0.279 ;
    LAYER M2 ;
      RECT 0.040 0.099 0.284 0.117 ;
    LAYER M2 ;
      RECT 0.040 0.153 0.284 0.171 ;
    LAYER M2 ;
      RECT 0.040 0.207 0.284 0.225 ;
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.000 0.585 0.432 0.603 ;   
  END
END DCL_NMOS_n12_X1_Y1
MACRO DCL_PMOS_n12_X5_Y2
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_n12_X5_Y2 0 0 ;
  SIZE 2.160 BY 1.188 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.017 0.094 1.035 0.770 ;
    END
  END S
  PIN BG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 1.125 2.160 1.143 ;
    END
  END BG
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.071 0.256 1.089 0.824 ;
    END
  END D
  OBS
    LAYER M2 ;
      RECT 0.094 0.261 2.120 0.279 ;
    LAYER M2 ;
      RECT 0.094 0.801 2.120 0.819 ;
    LAYER M2 ;
      RECT 0.040 0.099 2.012 0.117 ;
    LAYER M2 ;
      RECT 0.040 0.153 2.012 0.171 ;
    LAYER M2 ;
      RECT 0.040 0.207 2.012 0.225 ;
    LAYER M2 ;
      RECT 0.040 0.639 2.012 0.657 ;
    LAYER M2 ;
      RECT 0.040 0.693 2.012 0.711 ;
    LAYER M2 ;
      RECT 0.040 0.747 2.012 0.765 ;
    LAYER M1 ;
      RECT 0.000 1.125 2.160 1.143 ;
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.099 0.580 0.117 1.040 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.580 0.333 1.040 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.580 0.549 1.040 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.580 0.765 1.040 ;
    LAYER M1 ;
      RECT 0.963 0.040 0.981 0.500 ;
    LAYER M1 ;
      RECT 0.963 0.580 0.981 1.040 ;
    LAYER M1 ;
      RECT 1.179 0.040 1.197 0.500 ;
    LAYER M1 ;
      RECT 1.179 0.580 1.197 1.040 ;
    LAYER M1 ;
      RECT 1.395 0.040 1.413 0.500 ;
    LAYER M1 ;
      RECT 1.395 0.580 1.413 1.040 ;
    LAYER M1 ;
      RECT 1.611 0.040 1.629 0.500 ;
    LAYER M1 ;
      RECT 1.611 0.580 1.629 1.040 ;
    LAYER M1 ;
      RECT 1.827 0.040 1.845 0.500 ;
    LAYER M1 ;
      RECT 1.827 0.580 1.845 1.040 ;
    LAYER M1 ;
      RECT 2.043 0.040 2.061 0.500 ;
    LAYER M1 ;
      RECT 2.043 0.580 2.061 1.040 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.580 0.063 1.040 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.580 0.279 1.040 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.580 0.495 1.040 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.580 0.711 1.040 ;
    LAYER M1 ;
      RECT 0.909 0.040 0.927 0.500 ;
    LAYER M1 ;
      RECT 0.909 0.580 0.927 1.040 ;
    LAYER M1 ;
      RECT 1.125 0.040 1.143 0.500 ;
    LAYER M1 ;
      RECT 1.125 0.580 1.143 1.040 ;
    LAYER M1 ;
      RECT 1.341 0.040 1.359 0.500 ;
    LAYER M1 ;
      RECT 1.341 0.580 1.359 1.040 ;
    LAYER M1 ;
      RECT 1.557 0.040 1.575 0.500 ;
    LAYER M1 ;
      RECT 1.557 0.580 1.575 1.040 ;
    LAYER M1 ;
      RECT 1.773 0.040 1.791 0.500 ;
    LAYER M1 ;
      RECT 1.773 0.580 1.791 1.040 ;
    LAYER M1 ;
      RECT 1.989 0.040 2.007 0.500 ;
    LAYER M1 ;
      RECT 1.989 0.580 2.007 1.040 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.580 0.171 1.040 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.580 0.387 1.040 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.580 0.603 1.040 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.580 0.819 1.040 ;
    LAYER M1 ;
      RECT 1.017 0.040 1.035 0.500 ;
    LAYER M1 ;
      RECT 1.017 0.580 1.035 1.040 ;
    LAYER M1 ;
      RECT 1.233 0.040 1.251 0.500 ;
    LAYER M1 ;
      RECT 1.233 0.580 1.251 1.040 ;
    LAYER M1 ;
      RECT 1.449 0.040 1.467 0.500 ;
    LAYER M1 ;
      RECT 1.449 0.580 1.467 1.040 ;
    LAYER M1 ;
      RECT 1.665 0.040 1.683 0.500 ;
    LAYER M1 ;
      RECT 1.665 0.580 1.683 1.040 ;
    LAYER M1 ;
      RECT 1.881 0.040 1.899 0.500 ;
    LAYER M1 ;
      RECT 1.881 0.580 1.899 1.040 ;
    LAYER M1 ;
      RECT 2.097 0.040 2.115 0.500 ;
    LAYER M1 ;
      RECT 2.097 0.580 2.115 1.040 ;
  END
END DCL_PMOS_n12_X5_Y2
MACRO Switch_NMOS_n12_X2_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X2_Y2 0 0 ;
  SIZE 0.864 BY 1.188 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.369 0.094 0.387 0.770 ;
    END
  END S
  PIN BG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 1.125 0.864 1.143 ;
    END
  END BG
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.423 0.256 0.441 0.824 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.315 0.310 0.333 0.878 ;
    END
  END G
  OBS
    LAYER M2 ;
      RECT 0.094 0.315 0.770 0.333 ;
    LAYER M2 ;
      RECT 0.094 0.855 0.770 0.873 ;
    LAYER M2 ;
      RECT 0.148 0.261 0.824 0.279 ;
    LAYER M2 ;
      RECT 0.148 0.801 0.824 0.819 ;
    LAYER M2 ;
      RECT 0.040 0.099 0.716 0.117 ;
    LAYER M2 ;
      RECT 0.040 0.153 0.716 0.171 ;
    LAYER M2 ;
      RECT 0.040 0.207 0.716 0.225 ;
    LAYER M2 ;
      RECT 0.040 0.639 0.716 0.657 ;
    LAYER M2 ;
      RECT 0.040 0.693 0.716 0.711 ;
    LAYER M2 ;
      RECT 0.040 0.747 0.716 0.765 ;
    LAYER M1 ;
      RECT 0.000 1.125 0.864 1.143 ;
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.099 0.580 0.117 1.040 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.580 0.333 1.040 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.580 0.549 1.040 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.580 0.765 1.040 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.580 0.063 1.040 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.580 0.279 1.040 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.580 0.495 1.040 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.580 0.711 1.040 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.580 0.171 1.040 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.580 0.387 1.040 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.580 0.603 1.040 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.580 0.819 1.040 ;
  END
END Switch_NMOS_n12_X2_Y2
MACRO Switch_NMOS_n12_X4_Y4
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X4_Y4 0 0 ;
  SIZE 1.728 BY 2.268 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.801 0.094 0.819 1.850 ;
    END
  END S
  PIN BG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 2.205 1.728 2.223 ;
    END
  END BG
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.855 0.256 0.873 1.904 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.747 0.310 0.765 1.958 ;
    END
  END G
  OBS
    LAYER M2 ;
      RECT 0.094 0.315 1.634 0.333 ;
    LAYER M2 ;
      RECT 0.094 0.855 1.634 0.873 ;
    LAYER M2 ;
      RECT 0.094 1.395 1.634 1.413 ;
    LAYER M2 ;
      RECT 0.094 1.935 1.634 1.953 ;
    LAYER M2 ;
      RECT 0.148 0.261 1.688 0.279 ;
    LAYER M2 ;
      RECT 0.148 0.801 1.688 0.819 ;
    LAYER M2 ;
      RECT 0.148 1.341 1.688 1.359 ;
    LAYER M2 ;
      RECT 0.148 1.881 1.688 1.899 ;
    LAYER M2 ;
      RECT 0.040 0.099 1.580 0.117 ;
    LAYER M2 ;
      RECT 0.040 0.153 1.580 0.171 ;
    LAYER M2 ;
      RECT 0.040 0.207 1.580 0.225 ;
    LAYER M2 ;
      RECT 0.040 0.639 1.580 0.657 ;
    LAYER M2 ;
      RECT 0.040 0.693 1.580 0.711 ;
    LAYER M2 ;
      RECT 0.040 0.747 1.580 0.765 ;
    LAYER M2 ;
      RECT 0.040 1.179 1.580 1.197 ;
    LAYER M2 ;
      RECT 0.040 1.233 1.580 1.251 ;
    LAYER M2 ;
      RECT 0.040 1.287 1.580 1.305 ;
    LAYER M2 ;
      RECT 0.040 1.719 1.580 1.737 ;
    LAYER M2 ;
      RECT 0.040 1.773 1.580 1.791 ;
    LAYER M2 ;
      RECT 0.040 1.827 1.580 1.845 ;
    LAYER M1 ;
      RECT 0.000 2.205 1.728 2.223 ;
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.099 0.580 0.117 1.040 ;
    LAYER M1 ;
      RECT 0.099 1.120 0.117 1.580 ;
    LAYER M1 ;
      RECT 0.099 1.660 0.117 2.120 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.580 0.333 1.040 ;
    LAYER M1 ;
      RECT 0.315 1.120 0.333 1.580 ;
    LAYER M1 ;
      RECT 0.315 1.660 0.333 2.120 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.580 0.549 1.040 ;
    LAYER M1 ;
      RECT 0.531 1.120 0.549 1.580 ;
    LAYER M1 ;
      RECT 0.531 1.660 0.549 2.120 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.580 0.765 1.040 ;
    LAYER M1 ;
      RECT 0.747 1.120 0.765 1.580 ;
    LAYER M1 ;
      RECT 0.747 1.660 0.765 2.120 ;
    LAYER M1 ;
      RECT 0.963 0.040 0.981 0.500 ;
    LAYER M1 ;
      RECT 0.963 0.580 0.981 1.040 ;
    LAYER M1 ;
      RECT 0.963 1.120 0.981 1.580 ;
    LAYER M1 ;
      RECT 0.963 1.660 0.981 2.120 ;
    LAYER M1 ;
      RECT 1.179 0.040 1.197 0.500 ;
    LAYER M1 ;
      RECT 1.179 0.580 1.197 1.040 ;
    LAYER M1 ;
      RECT 1.179 1.120 1.197 1.580 ;
    LAYER M1 ;
      RECT 1.179 1.660 1.197 2.120 ;
    LAYER M1 ;
      RECT 1.395 0.040 1.413 0.500 ;
    LAYER M1 ;
      RECT 1.395 0.580 1.413 1.040 ;
    LAYER M1 ;
      RECT 1.395 1.120 1.413 1.580 ;
    LAYER M1 ;
      RECT 1.395 1.660 1.413 2.120 ;
    LAYER M1 ;
      RECT 1.611 0.040 1.629 0.500 ;
    LAYER M1 ;
      RECT 1.611 0.580 1.629 1.040 ;
    LAYER M1 ;
      RECT 1.611 1.120 1.629 1.580 ;
    LAYER M1 ;
      RECT 1.611 1.660 1.629 2.120 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.580 0.063 1.040 ;
    LAYER M1 ;
      RECT 0.045 1.120 0.063 1.580 ;
    LAYER M1 ;
      RECT 0.045 1.660 0.063 2.120 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.580 0.279 1.040 ;
    LAYER M1 ;
      RECT 0.261 1.120 0.279 1.580 ;
    LAYER M1 ;
      RECT 0.261 1.660 0.279 2.120 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.580 0.495 1.040 ;
    LAYER M1 ;
      RECT 0.477 1.120 0.495 1.580 ;
    LAYER M1 ;
      RECT 0.477 1.660 0.495 2.120 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.580 0.711 1.040 ;
    LAYER M1 ;
      RECT 0.693 1.120 0.711 1.580 ;
    LAYER M1 ;
      RECT 0.693 1.660 0.711 2.120 ;
    LAYER M1 ;
      RECT 0.909 0.040 0.927 0.500 ;
    LAYER M1 ;
      RECT 0.909 0.580 0.927 1.040 ;
    LAYER M1 ;
      RECT 0.909 1.120 0.927 1.580 ;
    LAYER M1 ;
      RECT 0.909 1.660 0.927 2.120 ;
    LAYER M1 ;
      RECT 1.125 0.040 1.143 0.500 ;
    LAYER M1 ;
      RECT 1.125 0.580 1.143 1.040 ;
    LAYER M1 ;
      RECT 1.125 1.120 1.143 1.580 ;
    LAYER M1 ;
      RECT 1.125 1.660 1.143 2.120 ;
    LAYER M1 ;
      RECT 1.341 0.040 1.359 0.500 ;
    LAYER M1 ;
      RECT 1.341 0.580 1.359 1.040 ;
    LAYER M1 ;
      RECT 1.341 1.120 1.359 1.580 ;
    LAYER M1 ;
      RECT 1.341 1.660 1.359 2.120 ;
    LAYER M1 ;
      RECT 1.557 0.040 1.575 0.500 ;
    LAYER M1 ;
      RECT 1.557 0.580 1.575 1.040 ;
    LAYER M1 ;
      RECT 1.557 1.120 1.575 1.580 ;
    LAYER M1 ;
      RECT 1.557 1.660 1.575 2.120 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.580 0.171 1.040 ;
    LAYER M1 ;
      RECT 0.153 1.120 0.171 1.580 ;
    LAYER M1 ;
      RECT 0.153 1.660 0.171 2.120 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.580 0.387 1.040 ;
    LAYER M1 ;
      RECT 0.369 1.120 0.387 1.580 ;
    LAYER M1 ;
      RECT 0.369 1.660 0.387 2.120 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.580 0.603 1.040 ;
    LAYER M1 ;
      RECT 0.585 1.120 0.603 1.580 ;
    LAYER M1 ;
      RECT 0.585 1.660 0.603 2.120 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.580 0.819 1.040 ;
    LAYER M1 ;
      RECT 0.801 1.120 0.819 1.580 ;
    LAYER M1 ;
      RECT 0.801 1.660 0.819 2.120 ;
    LAYER M1 ;
      RECT 1.017 0.040 1.035 0.500 ;
    LAYER M1 ;
      RECT 1.017 0.580 1.035 1.040 ;
    LAYER M1 ;
      RECT 1.017 1.120 1.035 1.580 ;
    LAYER M1 ;
      RECT 1.017 1.660 1.035 2.120 ;
    LAYER M1 ;
      RECT 1.233 0.040 1.251 0.500 ;
    LAYER M1 ;
      RECT 1.233 0.580 1.251 1.040 ;
    LAYER M1 ;
      RECT 1.233 1.120 1.251 1.580 ;
    LAYER M1 ;
      RECT 1.233 1.660 1.251 2.120 ;
    LAYER M1 ;
      RECT 1.449 0.040 1.467 0.500 ;
    LAYER M1 ;
      RECT 1.449 0.580 1.467 1.040 ;
    LAYER M1 ;
      RECT 1.449 1.120 1.467 1.580 ;
    LAYER M1 ;
      RECT 1.449 1.660 1.467 2.120 ;
    LAYER M1 ;
      RECT 1.665 0.040 1.683 0.500 ;
    LAYER M1 ;
      RECT 1.665 0.580 1.683 1.040 ;
    LAYER M1 ;
      RECT 1.665 1.120 1.683 1.580 ;
    LAYER M1 ;
      RECT 1.665 1.660 1.683 2.120 ;
  END
END Switch_NMOS_n12_X4_Y4
MACRO Switch_PMOS_n12_X5_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X5_Y2 0 0 ;
  SIZE 2.160 BY 1.188 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.017 0.094 1.035 0.770 ;
    END
  END S
  PIN BG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 1.125 2.160 1.143 ;
    END
  END BG
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.071 0.256 1.089 0.824 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.963 0.310 0.981 0.878 ;
    END
  END G
  OBS
    LAYER M2 ;
      RECT 0.094 0.315 2.066 0.333 ;
    LAYER M2 ;
      RECT 0.094 0.855 2.066 0.873 ;
    LAYER M2 ;
      RECT 0.148 0.261 2.120 0.279 ;
    LAYER M2 ;
      RECT 0.148 0.801 2.120 0.819 ;
    LAYER M2 ;
      RECT 0.040 0.099 2.012 0.117 ;
    LAYER M2 ;
      RECT 0.040 0.153 2.012 0.171 ;
    LAYER M2 ;
      RECT 0.040 0.207 2.012 0.225 ;
    LAYER M2 ;
      RECT 0.040 0.639 2.012 0.657 ;
    LAYER M2 ;
      RECT 0.040 0.693 2.012 0.711 ;
    LAYER M2 ;
      RECT 0.040 0.747 2.012 0.765 ;
    LAYER M1 ;
      RECT 0.000 1.125 2.160 1.143 ;
    LAYER M1 ;
      RECT 0.099 0.040 0.117 0.500 ;
    LAYER M1 ;
      RECT 0.099 0.580 0.117 1.040 ;
    LAYER M1 ;
      RECT 0.315 0.040 0.333 0.500 ;
    LAYER M1 ;
      RECT 0.315 0.580 0.333 1.040 ;
    LAYER M1 ;
      RECT 0.531 0.040 0.549 0.500 ;
    LAYER M1 ;
      RECT 0.531 0.580 0.549 1.040 ;
    LAYER M1 ;
      RECT 0.747 0.040 0.765 0.500 ;
    LAYER M1 ;
      RECT 0.747 0.580 0.765 1.040 ;
    LAYER M1 ;
      RECT 0.963 0.040 0.981 0.500 ;
    LAYER M1 ;
      RECT 0.963 0.580 0.981 1.040 ;
    LAYER M1 ;
      RECT 1.179 0.040 1.197 0.500 ;
    LAYER M1 ;
      RECT 1.179 0.580 1.197 1.040 ;
    LAYER M1 ;
      RECT 1.395 0.040 1.413 0.500 ;
    LAYER M1 ;
      RECT 1.395 0.580 1.413 1.040 ;
    LAYER M1 ;
      RECT 1.611 0.040 1.629 0.500 ;
    LAYER M1 ;
      RECT 1.611 0.580 1.629 1.040 ;
    LAYER M1 ;
      RECT 1.827 0.040 1.845 0.500 ;
    LAYER M1 ;
      RECT 1.827 0.580 1.845 1.040 ;
    LAYER M1 ;
      RECT 2.043 0.040 2.061 0.500 ;
    LAYER M1 ;
      RECT 2.043 0.580 2.061 1.040 ;
    LAYER M1 ;
      RECT 0.045 0.040 0.063 0.500 ;
    LAYER M1 ;
      RECT 0.045 0.580 0.063 1.040 ;
    LAYER M1 ;
      RECT 0.261 0.040 0.279 0.500 ;
    LAYER M1 ;
      RECT 0.261 0.580 0.279 1.040 ;
    LAYER M1 ;
      RECT 0.477 0.040 0.495 0.500 ;
    LAYER M1 ;
      RECT 0.477 0.580 0.495 1.040 ;
    LAYER M1 ;
      RECT 0.693 0.040 0.711 0.500 ;
    LAYER M1 ;
      RECT 0.693 0.580 0.711 1.040 ;
    LAYER M1 ;
      RECT 0.909 0.040 0.927 0.500 ;
    LAYER M1 ;
      RECT 0.909 0.580 0.927 1.040 ;
    LAYER M1 ;
      RECT 1.125 0.040 1.143 0.500 ;
    LAYER M1 ;
      RECT 1.125 0.580 1.143 1.040 ;
    LAYER M1 ;
      RECT 1.341 0.040 1.359 0.500 ;
    LAYER M1 ;
      RECT 1.341 0.580 1.359 1.040 ;
    LAYER M1 ;
      RECT 1.557 0.040 1.575 0.500 ;
    LAYER M1 ;
      RECT 1.557 0.580 1.575 1.040 ;
    LAYER M1 ;
      RECT 1.773 0.040 1.791 0.500 ;
    LAYER M1 ;
      RECT 1.773 0.580 1.791 1.040 ;
    LAYER M1 ;
      RECT 1.989 0.040 2.007 0.500 ;
    LAYER M1 ;
      RECT 1.989 0.580 2.007 1.040 ;
    LAYER M1 ;
      RECT 0.153 0.040 0.171 0.500 ;
    LAYER M1 ;
      RECT 0.153 0.580 0.171 1.040 ;
    LAYER M1 ;
      RECT 0.369 0.040 0.387 0.500 ;
    LAYER M1 ;
      RECT 0.369 0.580 0.387 1.040 ;
    LAYER M1 ;
      RECT 0.585 0.040 0.603 0.500 ;
    LAYER M1 ;
      RECT 0.585 0.580 0.603 1.040 ;
    LAYER M1 ;
      RECT 0.801 0.040 0.819 0.500 ;
    LAYER M1 ;
      RECT 0.801 0.580 0.819 1.040 ;
    LAYER M1 ;
      RECT 1.017 0.040 1.035 0.500 ;
    LAYER M1 ;
      RECT 1.017 0.580 1.035 1.040 ;
    LAYER M1 ;
      RECT 1.233 0.040 1.251 0.500 ;
    LAYER M1 ;
      RECT 1.233 0.580 1.251 1.040 ;
    LAYER M1 ;
      RECT 1.449 0.040 1.467 0.500 ;
    LAYER M1 ;
      RECT 1.449 0.580 1.467 1.040 ;
    LAYER M1 ;
      RECT 1.665 0.040 1.683 0.500 ;
    LAYER M1 ;
      RECT 1.665 0.580 1.683 1.040 ;
    LAYER M1 ;
      RECT 1.881 0.040 1.899 0.500 ;
    LAYER M1 ;
      RECT 1.881 0.580 1.899 1.040 ;
    LAYER M1 ;
      RECT 2.097 0.040 2.115 0.500 ;
    LAYER M1 ;
      RECT 2.097 0.580 2.115 1.040 ;
  END
END Switch_PMOS_n12_X5_Y2
