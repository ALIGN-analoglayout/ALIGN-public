MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 9.2 BY 25.872 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 25.584 3.232 25.656 ;
      LAYER M2 ;
        RECT 3.18 25.604 3.252 25.636 ;
      LAYER M1 ;
        RECT 6.176 25.584 6.208 25.656 ;
      LAYER M2 ;
        RECT 6.156 25.604 6.228 25.636 ;
      LAYER M2 ;
        RECT 3.216 25.604 6.192 25.636 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 3.056 10.148 5.808 10.18 ;
  LAYER M1 ;
        RECT 3.04 10.128 3.072 10.2 ;
  LAYER M2 ;
        RECT 3.02 10.148 3.092 10.18 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M2 ;
        RECT 3.056 13.256 5.808 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M2 ;
        RECT 3.056 7.04 5.808 7.072 ;
  LAYER M1 ;
        RECT 3.04 7.02 3.072 7.092 ;
  LAYER M2 ;
        RECT 3.02 7.04 3.092 7.072 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 16.416 ;
  LAYER M2 ;
        RECT 5.772 16.364 5.844 16.396 ;
  LAYER M2 ;
        RECT 3.056 16.364 5.808 16.396 ;
  LAYER M1 ;
        RECT 3.04 16.344 3.072 16.416 ;
  LAYER M2 ;
        RECT 3.02 16.364 3.092 16.396 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M2 ;
        RECT 3.056 3.932 5.808 3.964 ;
  LAYER M1 ;
        RECT 3.04 3.912 3.072 3.984 ;
  LAYER M2 ;
        RECT 3.02 3.932 3.092 3.964 ;
  LAYER M1 ;
        RECT 5.792 19.452 5.824 19.524 ;
  LAYER M2 ;
        RECT 5.772 19.472 5.844 19.504 ;
  LAYER M2 ;
        RECT 3.056 19.472 5.808 19.504 ;
  LAYER M1 ;
        RECT 3.04 19.452 3.072 19.524 ;
  LAYER M2 ;
        RECT 3.02 19.472 3.092 19.504 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.504 ;
  LAYER M1 ;
        RECT 3.04 0.504 3.072 19.488 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M1 ;
        RECT 5.792 9.996 5.824 10.164 ;
  LAYER M1 ;
        RECT 5.792 9.96 5.824 10.032 ;
  LAYER M2 ;
        RECT 5.772 9.98 5.844 10.012 ;
  LAYER M2 ;
        RECT 5.808 9.98 6.032 10.012 ;
  LAYER M1 ;
        RECT 6.016 9.96 6.048 10.032 ;
  LAYER M2 ;
        RECT 5.996 9.98 6.068 10.012 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M1 ;
        RECT 5.792 13.104 5.824 13.272 ;
  LAYER M1 ;
        RECT 5.792 13.068 5.824 13.14 ;
  LAYER M2 ;
        RECT 5.772 13.088 5.844 13.12 ;
  LAYER M2 ;
        RECT 5.808 13.088 6.032 13.12 ;
  LAYER M1 ;
        RECT 6.016 13.068 6.048 13.14 ;
  LAYER M2 ;
        RECT 5.996 13.088 6.068 13.12 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M1 ;
        RECT 5.792 6.888 5.824 7.056 ;
  LAYER M1 ;
        RECT 5.792 6.852 5.824 6.924 ;
  LAYER M2 ;
        RECT 5.772 6.872 5.844 6.904 ;
  LAYER M2 ;
        RECT 5.808 6.872 6.032 6.904 ;
  LAYER M1 ;
        RECT 6.016 6.852 6.048 6.924 ;
  LAYER M2 ;
        RECT 5.996 6.872 6.068 6.904 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 16.416 ;
  LAYER M2 ;
        RECT 5.772 16.364 5.844 16.396 ;
  LAYER M1 ;
        RECT 5.792 16.212 5.824 16.38 ;
  LAYER M1 ;
        RECT 5.792 16.176 5.824 16.248 ;
  LAYER M2 ;
        RECT 5.772 16.196 5.844 16.228 ;
  LAYER M2 ;
        RECT 5.808 16.196 6.032 16.228 ;
  LAYER M1 ;
        RECT 6.016 16.176 6.048 16.248 ;
  LAYER M2 ;
        RECT 5.996 16.196 6.068 16.228 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M1 ;
        RECT 5.792 3.78 5.824 3.948 ;
  LAYER M1 ;
        RECT 5.792 3.744 5.824 3.816 ;
  LAYER M2 ;
        RECT 5.772 3.764 5.844 3.796 ;
  LAYER M2 ;
        RECT 5.808 3.764 6.032 3.796 ;
  LAYER M1 ;
        RECT 6.016 3.744 6.048 3.816 ;
  LAYER M2 ;
        RECT 5.996 3.764 6.068 3.796 ;
  LAYER M1 ;
        RECT 5.792 19.452 5.824 19.524 ;
  LAYER M2 ;
        RECT 5.772 19.472 5.844 19.504 ;
  LAYER M1 ;
        RECT 5.792 19.32 5.824 19.488 ;
  LAYER M1 ;
        RECT 5.792 19.284 5.824 19.356 ;
  LAYER M2 ;
        RECT 5.772 19.304 5.844 19.336 ;
  LAYER M2 ;
        RECT 5.808 19.304 6.032 19.336 ;
  LAYER M1 ;
        RECT 6.016 19.284 6.048 19.356 ;
  LAYER M2 ;
        RECT 5.996 19.304 6.068 19.336 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.504 ;
  LAYER M1 ;
        RECT 6.016 0.504 6.048 19.32 ;
  LAYER M2 ;
        RECT 3.056 0.236 6.032 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M2 ;
        RECT 0.08 0.824 2.832 0.856 ;
  LAYER M1 ;
        RECT 0.064 0.804 0.096 0.876 ;
  LAYER M2 ;
        RECT 0.044 0.824 0.116 0.856 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M2 ;
        RECT 0.08 3.932 2.832 3.964 ;
  LAYER M1 ;
        RECT 0.064 3.912 0.096 3.984 ;
  LAYER M2 ;
        RECT 0.044 3.932 0.116 3.964 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M2 ;
        RECT 0.08 7.04 2.832 7.072 ;
  LAYER M1 ;
        RECT 0.064 7.02 0.096 7.092 ;
  LAYER M2 ;
        RECT 0.044 7.04 0.116 7.072 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M2 ;
        RECT 0.08 10.148 2.832 10.18 ;
  LAYER M1 ;
        RECT 0.064 10.128 0.096 10.2 ;
  LAYER M2 ;
        RECT 0.044 10.148 0.116 10.18 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 13.308 ;
  LAYER M2 ;
        RECT 2.796 13.256 2.868 13.288 ;
  LAYER M2 ;
        RECT 0.08 13.256 2.832 13.288 ;
  LAYER M1 ;
        RECT 0.064 13.236 0.096 13.308 ;
  LAYER M2 ;
        RECT 0.044 13.256 0.116 13.288 ;
  LAYER M1 ;
        RECT 2.816 16.344 2.848 16.416 ;
  LAYER M2 ;
        RECT 2.796 16.364 2.868 16.396 ;
  LAYER M2 ;
        RECT 0.08 16.364 2.832 16.396 ;
  LAYER M1 ;
        RECT 0.064 16.344 0.096 16.416 ;
  LAYER M2 ;
        RECT 0.044 16.364 0.116 16.396 ;
  LAYER M1 ;
        RECT 2.816 19.452 2.848 19.524 ;
  LAYER M2 ;
        RECT 2.796 19.472 2.868 19.504 ;
  LAYER M2 ;
        RECT 0.08 19.472 2.832 19.504 ;
  LAYER M1 ;
        RECT 0.064 19.452 0.096 19.524 ;
  LAYER M2 ;
        RECT 0.044 19.472 0.116 19.504 ;
  LAYER M1 ;
        RECT 2.816 22.56 2.848 22.632 ;
  LAYER M2 ;
        RECT 2.796 22.58 2.868 22.612 ;
  LAYER M2 ;
        RECT 0.08 22.58 2.832 22.612 ;
  LAYER M1 ;
        RECT 0.064 22.56 0.096 22.632 ;
  LAYER M2 ;
        RECT 0.044 22.58 0.116 22.612 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.504 ;
  LAYER M1 ;
        RECT 0.064 0.504 0.096 22.596 ;
  LAYER M1 ;
        RECT 8.768 0.804 8.8 0.876 ;
  LAYER M2 ;
        RECT 8.748 0.824 8.82 0.856 ;
  LAYER M1 ;
        RECT 8.768 0.672 8.8 0.84 ;
  LAYER M1 ;
        RECT 8.768 0.636 8.8 0.708 ;
  LAYER M2 ;
        RECT 8.748 0.656 8.82 0.688 ;
  LAYER M2 ;
        RECT 8.784 0.656 9.008 0.688 ;
  LAYER M1 ;
        RECT 8.992 0.636 9.024 0.708 ;
  LAYER M2 ;
        RECT 8.972 0.656 9.044 0.688 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M1 ;
        RECT 8.768 3.78 8.8 3.948 ;
  LAYER M1 ;
        RECT 8.768 3.744 8.8 3.816 ;
  LAYER M2 ;
        RECT 8.748 3.764 8.82 3.796 ;
  LAYER M2 ;
        RECT 8.784 3.764 9.008 3.796 ;
  LAYER M1 ;
        RECT 8.992 3.744 9.024 3.816 ;
  LAYER M2 ;
        RECT 8.972 3.764 9.044 3.796 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M1 ;
        RECT 8.768 6.888 8.8 7.056 ;
  LAYER M1 ;
        RECT 8.768 6.852 8.8 6.924 ;
  LAYER M2 ;
        RECT 8.748 6.872 8.82 6.904 ;
  LAYER M2 ;
        RECT 8.784 6.872 9.008 6.904 ;
  LAYER M1 ;
        RECT 8.992 6.852 9.024 6.924 ;
  LAYER M2 ;
        RECT 8.972 6.872 9.044 6.904 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M1 ;
        RECT 8.768 9.996 8.8 10.164 ;
  LAYER M1 ;
        RECT 8.768 9.96 8.8 10.032 ;
  LAYER M2 ;
        RECT 8.748 9.98 8.82 10.012 ;
  LAYER M2 ;
        RECT 8.784 9.98 9.008 10.012 ;
  LAYER M1 ;
        RECT 8.992 9.96 9.024 10.032 ;
  LAYER M2 ;
        RECT 8.972 9.98 9.044 10.012 ;
  LAYER M1 ;
        RECT 8.768 13.236 8.8 13.308 ;
  LAYER M2 ;
        RECT 8.748 13.256 8.82 13.288 ;
  LAYER M1 ;
        RECT 8.768 13.104 8.8 13.272 ;
  LAYER M1 ;
        RECT 8.768 13.068 8.8 13.14 ;
  LAYER M2 ;
        RECT 8.748 13.088 8.82 13.12 ;
  LAYER M2 ;
        RECT 8.784 13.088 9.008 13.12 ;
  LAYER M1 ;
        RECT 8.992 13.068 9.024 13.14 ;
  LAYER M2 ;
        RECT 8.972 13.088 9.044 13.12 ;
  LAYER M1 ;
        RECT 8.768 16.344 8.8 16.416 ;
  LAYER M2 ;
        RECT 8.748 16.364 8.82 16.396 ;
  LAYER M1 ;
        RECT 8.768 16.212 8.8 16.38 ;
  LAYER M1 ;
        RECT 8.768 16.176 8.8 16.248 ;
  LAYER M2 ;
        RECT 8.748 16.196 8.82 16.228 ;
  LAYER M2 ;
        RECT 8.784 16.196 9.008 16.228 ;
  LAYER M1 ;
        RECT 8.992 16.176 9.024 16.248 ;
  LAYER M2 ;
        RECT 8.972 16.196 9.044 16.228 ;
  LAYER M1 ;
        RECT 8.768 19.452 8.8 19.524 ;
  LAYER M2 ;
        RECT 8.748 19.472 8.82 19.504 ;
  LAYER M1 ;
        RECT 8.768 19.32 8.8 19.488 ;
  LAYER M1 ;
        RECT 8.768 19.284 8.8 19.356 ;
  LAYER M2 ;
        RECT 8.748 19.304 8.82 19.336 ;
  LAYER M2 ;
        RECT 8.784 19.304 9.008 19.336 ;
  LAYER M1 ;
        RECT 8.992 19.284 9.024 19.356 ;
  LAYER M2 ;
        RECT 8.972 19.304 9.044 19.336 ;
  LAYER M1 ;
        RECT 8.768 22.56 8.8 22.632 ;
  LAYER M2 ;
        RECT 8.748 22.58 8.82 22.612 ;
  LAYER M1 ;
        RECT 8.768 22.428 8.8 22.596 ;
  LAYER M1 ;
        RECT 8.768 22.392 8.8 22.464 ;
  LAYER M2 ;
        RECT 8.748 22.412 8.82 22.444 ;
  LAYER M2 ;
        RECT 8.784 22.412 9.008 22.444 ;
  LAYER M1 ;
        RECT 8.992 22.392 9.024 22.464 ;
  LAYER M2 ;
        RECT 8.972 22.412 9.044 22.444 ;
  LAYER M1 ;
        RECT 8.992 0.048 9.024 0.12 ;
  LAYER M2 ;
        RECT 8.972 0.068 9.044 0.1 ;
  LAYER M1 ;
        RECT 8.992 0.084 9.024 0.504 ;
  LAYER M1 ;
        RECT 8.992 0.504 9.024 22.428 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.008 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.804 5.824 0.876 ;
  LAYER M2 ;
        RECT 5.772 0.824 5.844 0.856 ;
  LAYER M2 ;
        RECT 2.832 0.824 5.808 0.856 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M1 ;
        RECT 5.792 22.56 5.824 22.632 ;
  LAYER M2 ;
        RECT 5.772 22.58 5.844 22.612 ;
  LAYER M2 ;
        RECT 2.832 22.58 5.808 22.612 ;
  LAYER M1 ;
        RECT 2.816 22.56 2.848 22.632 ;
  LAYER M2 ;
        RECT 2.796 22.58 2.868 22.612 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M2 ;
        RECT 3.216 12.584 3.44 12.616 ;
  LAYER M1 ;
        RECT 3.2 12.564 3.232 12.636 ;
  LAYER M2 ;
        RECT 3.18 12.584 3.252 12.616 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M2 ;
        RECT 3.216 15.692 3.44 15.724 ;
  LAYER M1 ;
        RECT 3.2 15.672 3.232 15.744 ;
  LAYER M2 ;
        RECT 3.18 15.692 3.252 15.724 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M2 ;
        RECT 3.216 9.476 3.44 9.508 ;
  LAYER M1 ;
        RECT 3.2 9.456 3.232 9.528 ;
  LAYER M2 ;
        RECT 3.18 9.476 3.252 9.508 ;
  LAYER M1 ;
        RECT 3.424 18.78 3.456 18.852 ;
  LAYER M2 ;
        RECT 3.404 18.8 3.476 18.832 ;
  LAYER M2 ;
        RECT 3.216 18.8 3.44 18.832 ;
  LAYER M1 ;
        RECT 3.2 18.78 3.232 18.852 ;
  LAYER M2 ;
        RECT 3.18 18.8 3.252 18.832 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M2 ;
        RECT 3.216 6.368 3.44 6.4 ;
  LAYER M1 ;
        RECT 3.2 6.348 3.232 6.42 ;
  LAYER M2 ;
        RECT 3.18 6.368 3.252 6.4 ;
  LAYER M1 ;
        RECT 3.424 21.888 3.456 21.96 ;
  LAYER M2 ;
        RECT 3.404 21.908 3.476 21.94 ;
  LAYER M2 ;
        RECT 3.216 21.908 3.44 21.94 ;
  LAYER M1 ;
        RECT 3.2 21.888 3.232 21.96 ;
  LAYER M2 ;
        RECT 3.18 21.908 3.252 21.94 ;
  LAYER M1 ;
        RECT 3.2 25.584 3.232 25.656 ;
  LAYER M2 ;
        RECT 3.18 25.604 3.252 25.636 ;
  LAYER M1 ;
        RECT 3.2 25.368 3.232 25.62 ;
  LAYER M1 ;
        RECT 3.2 6.384 3.232 25.368 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M1 ;
        RECT 3.424 12.6 3.456 12.768 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.44 12.752 6.192 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M1 ;
        RECT 3.424 15.708 3.456 15.876 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 3.44 15.86 6.192 15.892 ;
  LAYER M1 ;
        RECT 6.176 15.84 6.208 15.912 ;
  LAYER M2 ;
        RECT 6.156 15.86 6.228 15.892 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M1 ;
        RECT 3.424 9.492 3.456 9.66 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M2 ;
        RECT 3.44 9.644 6.192 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 3.424 18.78 3.456 18.852 ;
  LAYER M2 ;
        RECT 3.404 18.8 3.476 18.832 ;
  LAYER M1 ;
        RECT 3.424 18.816 3.456 18.984 ;
  LAYER M1 ;
        RECT 3.424 18.948 3.456 19.02 ;
  LAYER M2 ;
        RECT 3.404 18.968 3.476 19 ;
  LAYER M2 ;
        RECT 3.44 18.968 6.192 19 ;
  LAYER M1 ;
        RECT 6.176 18.948 6.208 19.02 ;
  LAYER M2 ;
        RECT 6.156 18.968 6.228 19 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M1 ;
        RECT 3.424 6.384 3.456 6.552 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M2 ;
        RECT 3.44 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 3.424 21.888 3.456 21.96 ;
  LAYER M2 ;
        RECT 3.404 21.908 3.476 21.94 ;
  LAYER M1 ;
        RECT 3.424 21.924 3.456 22.092 ;
  LAYER M1 ;
        RECT 3.424 22.056 3.456 22.128 ;
  LAYER M2 ;
        RECT 3.404 22.076 3.476 22.108 ;
  LAYER M2 ;
        RECT 3.44 22.076 6.192 22.108 ;
  LAYER M1 ;
        RECT 6.176 22.056 6.208 22.128 ;
  LAYER M2 ;
        RECT 6.156 22.076 6.228 22.108 ;
  LAYER M1 ;
        RECT 6.176 25.584 6.208 25.656 ;
  LAYER M2 ;
        RECT 6.156 25.604 6.228 25.636 ;
  LAYER M1 ;
        RECT 6.176 25.368 6.208 25.62 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 25.368 ;
  LAYER M2 ;
        RECT 3.216 25.604 6.192 25.636 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M2 ;
        RECT 0.24 3.26 0.464 3.292 ;
  LAYER M1 ;
        RECT 0.224 3.24 0.256 3.312 ;
  LAYER M2 ;
        RECT 0.204 3.26 0.276 3.292 ;
  LAYER M1 ;
        RECT 0.448 6.348 0.48 6.42 ;
  LAYER M2 ;
        RECT 0.428 6.368 0.5 6.4 ;
  LAYER M2 ;
        RECT 0.24 6.368 0.464 6.4 ;
  LAYER M1 ;
        RECT 0.224 6.348 0.256 6.42 ;
  LAYER M2 ;
        RECT 0.204 6.368 0.276 6.4 ;
  LAYER M1 ;
        RECT 0.448 9.456 0.48 9.528 ;
  LAYER M2 ;
        RECT 0.428 9.476 0.5 9.508 ;
  LAYER M2 ;
        RECT 0.24 9.476 0.464 9.508 ;
  LAYER M1 ;
        RECT 0.224 9.456 0.256 9.528 ;
  LAYER M2 ;
        RECT 0.204 9.476 0.276 9.508 ;
  LAYER M1 ;
        RECT 0.448 12.564 0.48 12.636 ;
  LAYER M2 ;
        RECT 0.428 12.584 0.5 12.616 ;
  LAYER M2 ;
        RECT 0.24 12.584 0.464 12.616 ;
  LAYER M1 ;
        RECT 0.224 12.564 0.256 12.636 ;
  LAYER M2 ;
        RECT 0.204 12.584 0.276 12.616 ;
  LAYER M1 ;
        RECT 0.448 15.672 0.48 15.744 ;
  LAYER M2 ;
        RECT 0.428 15.692 0.5 15.724 ;
  LAYER M2 ;
        RECT 0.24 15.692 0.464 15.724 ;
  LAYER M1 ;
        RECT 0.224 15.672 0.256 15.744 ;
  LAYER M2 ;
        RECT 0.204 15.692 0.276 15.724 ;
  LAYER M1 ;
        RECT 0.448 18.78 0.48 18.852 ;
  LAYER M2 ;
        RECT 0.428 18.8 0.5 18.832 ;
  LAYER M2 ;
        RECT 0.24 18.8 0.464 18.832 ;
  LAYER M1 ;
        RECT 0.224 18.78 0.256 18.852 ;
  LAYER M2 ;
        RECT 0.204 18.8 0.276 18.832 ;
  LAYER M1 ;
        RECT 0.448 21.888 0.48 21.96 ;
  LAYER M2 ;
        RECT 0.428 21.908 0.5 21.94 ;
  LAYER M2 ;
        RECT 0.24 21.908 0.464 21.94 ;
  LAYER M1 ;
        RECT 0.224 21.888 0.256 21.96 ;
  LAYER M2 ;
        RECT 0.204 21.908 0.276 21.94 ;
  LAYER M1 ;
        RECT 0.448 24.996 0.48 25.068 ;
  LAYER M2 ;
        RECT 0.428 25.016 0.5 25.048 ;
  LAYER M2 ;
        RECT 0.24 25.016 0.464 25.048 ;
  LAYER M1 ;
        RECT 0.224 24.996 0.256 25.068 ;
  LAYER M2 ;
        RECT 0.204 25.016 0.276 25.048 ;
  LAYER M1 ;
        RECT 0.224 25.752 0.256 25.824 ;
  LAYER M2 ;
        RECT 0.204 25.772 0.276 25.804 ;
  LAYER M1 ;
        RECT 0.224 25.368 0.256 25.788 ;
  LAYER M1 ;
        RECT 0.224 3.276 0.256 25.368 ;
  LAYER M1 ;
        RECT 6.4 3.24 6.432 3.312 ;
  LAYER M2 ;
        RECT 6.38 3.26 6.452 3.292 ;
  LAYER M1 ;
        RECT 6.4 3.276 6.432 3.444 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.168 3.46 ;
  LAYER M1 ;
        RECT 9.152 3.408 9.184 3.48 ;
  LAYER M2 ;
        RECT 9.132 3.428 9.204 3.46 ;
  LAYER M1 ;
        RECT 6.4 6.348 6.432 6.42 ;
  LAYER M2 ;
        RECT 6.38 6.368 6.452 6.4 ;
  LAYER M1 ;
        RECT 6.4 6.384 6.432 6.552 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.416 6.536 9.168 6.568 ;
  LAYER M1 ;
        RECT 9.152 6.516 9.184 6.588 ;
  LAYER M2 ;
        RECT 9.132 6.536 9.204 6.568 ;
  LAYER M1 ;
        RECT 6.4 9.456 6.432 9.528 ;
  LAYER M2 ;
        RECT 6.38 9.476 6.452 9.508 ;
  LAYER M1 ;
        RECT 6.4 9.492 6.432 9.66 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M2 ;
        RECT 6.416 9.644 9.168 9.676 ;
  LAYER M1 ;
        RECT 9.152 9.624 9.184 9.696 ;
  LAYER M2 ;
        RECT 9.132 9.644 9.204 9.676 ;
  LAYER M1 ;
        RECT 6.4 12.564 6.432 12.636 ;
  LAYER M2 ;
        RECT 6.38 12.584 6.452 12.616 ;
  LAYER M1 ;
        RECT 6.4 12.6 6.432 12.768 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 6.416 12.752 9.168 12.784 ;
  LAYER M1 ;
        RECT 9.152 12.732 9.184 12.804 ;
  LAYER M2 ;
        RECT 9.132 12.752 9.204 12.784 ;
  LAYER M1 ;
        RECT 6.4 15.672 6.432 15.744 ;
  LAYER M2 ;
        RECT 6.38 15.692 6.452 15.724 ;
  LAYER M1 ;
        RECT 6.4 15.708 6.432 15.876 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M2 ;
        RECT 6.416 15.86 9.168 15.892 ;
  LAYER M1 ;
        RECT 9.152 15.84 9.184 15.912 ;
  LAYER M2 ;
        RECT 9.132 15.86 9.204 15.892 ;
  LAYER M1 ;
        RECT 6.4 18.78 6.432 18.852 ;
  LAYER M2 ;
        RECT 6.38 18.8 6.452 18.832 ;
  LAYER M1 ;
        RECT 6.4 18.816 6.432 18.984 ;
  LAYER M1 ;
        RECT 6.4 18.948 6.432 19.02 ;
  LAYER M2 ;
        RECT 6.38 18.968 6.452 19 ;
  LAYER M2 ;
        RECT 6.416 18.968 9.168 19 ;
  LAYER M1 ;
        RECT 9.152 18.948 9.184 19.02 ;
  LAYER M2 ;
        RECT 9.132 18.968 9.204 19 ;
  LAYER M1 ;
        RECT 6.4 21.888 6.432 21.96 ;
  LAYER M2 ;
        RECT 6.38 21.908 6.452 21.94 ;
  LAYER M1 ;
        RECT 6.4 21.924 6.432 22.092 ;
  LAYER M1 ;
        RECT 6.4 22.056 6.432 22.128 ;
  LAYER M2 ;
        RECT 6.38 22.076 6.452 22.108 ;
  LAYER M2 ;
        RECT 6.416 22.076 9.168 22.108 ;
  LAYER M1 ;
        RECT 9.152 22.056 9.184 22.128 ;
  LAYER M2 ;
        RECT 9.132 22.076 9.204 22.108 ;
  LAYER M1 ;
        RECT 6.4 24.996 6.432 25.068 ;
  LAYER M2 ;
        RECT 6.38 25.016 6.452 25.048 ;
  LAYER M1 ;
        RECT 6.4 25.032 6.432 25.2 ;
  LAYER M1 ;
        RECT 6.4 25.164 6.432 25.236 ;
  LAYER M2 ;
        RECT 6.38 25.184 6.452 25.216 ;
  LAYER M2 ;
        RECT 6.416 25.184 9.168 25.216 ;
  LAYER M1 ;
        RECT 9.152 25.164 9.184 25.236 ;
  LAYER M2 ;
        RECT 9.132 25.184 9.204 25.216 ;
  LAYER M1 ;
        RECT 9.152 25.752 9.184 25.824 ;
  LAYER M2 ;
        RECT 9.132 25.772 9.204 25.804 ;
  LAYER M1 ;
        RECT 9.152 25.368 9.184 25.788 ;
  LAYER M1 ;
        RECT 9.152 3.444 9.184 25.368 ;
  LAYER M2 ;
        RECT 0.24 25.772 9.168 25.804 ;
  LAYER M1 ;
        RECT 3.424 3.24 3.456 3.312 ;
  LAYER M2 ;
        RECT 3.404 3.26 3.476 3.292 ;
  LAYER M2 ;
        RECT 0.464 3.26 3.44 3.292 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M1 ;
        RECT 3.424 24.996 3.456 25.068 ;
  LAYER M2 ;
        RECT 3.404 25.016 3.476 25.048 ;
  LAYER M2 ;
        RECT 0.464 25.016 3.44 25.048 ;
  LAYER M1 ;
        RECT 0.448 24.996 0.48 25.068 ;
  LAYER M2 ;
        RECT 0.428 25.016 0.5 25.048 ;
  LAYER M1 ;
        RECT 0.448 0.804 0.48 3.312 ;
  LAYER M3 ;
        RECT 0.448 3.26 0.48 3.292 ;
  LAYER M1 ;
        RECT 0.512 0.804 0.544 3.312 ;
  LAYER M3 ;
        RECT 0.512 0.824 0.544 0.856 ;
  LAYER M1 ;
        RECT 0.576 0.804 0.608 3.312 ;
  LAYER M3 ;
        RECT 0.576 3.26 0.608 3.292 ;
  LAYER M1 ;
        RECT 0.64 0.804 0.672 3.312 ;
  LAYER M3 ;
        RECT 0.64 0.824 0.672 0.856 ;
  LAYER M1 ;
        RECT 0.704 0.804 0.736 3.312 ;
  LAYER M3 ;
        RECT 0.704 3.26 0.736 3.292 ;
  LAYER M1 ;
        RECT 0.768 0.804 0.8 3.312 ;
  LAYER M3 ;
        RECT 0.768 0.824 0.8 0.856 ;
  LAYER M1 ;
        RECT 0.832 0.804 0.864 3.312 ;
  LAYER M3 ;
        RECT 0.832 3.26 0.864 3.292 ;
  LAYER M1 ;
        RECT 0.896 0.804 0.928 3.312 ;
  LAYER M3 ;
        RECT 0.896 0.824 0.928 0.856 ;
  LAYER M1 ;
        RECT 0.96 0.804 0.992 3.312 ;
  LAYER M3 ;
        RECT 0.96 3.26 0.992 3.292 ;
  LAYER M1 ;
        RECT 1.024 0.804 1.056 3.312 ;
  LAYER M3 ;
        RECT 1.024 0.824 1.056 0.856 ;
  LAYER M1 ;
        RECT 1.088 0.804 1.12 3.312 ;
  LAYER M3 ;
        RECT 1.088 3.26 1.12 3.292 ;
  LAYER M1 ;
        RECT 1.152 0.804 1.184 3.312 ;
  LAYER M3 ;
        RECT 1.152 0.824 1.184 0.856 ;
  LAYER M1 ;
        RECT 1.216 0.804 1.248 3.312 ;
  LAYER M3 ;
        RECT 1.216 3.26 1.248 3.292 ;
  LAYER M1 ;
        RECT 1.28 0.804 1.312 3.312 ;
  LAYER M3 ;
        RECT 1.28 0.824 1.312 0.856 ;
  LAYER M1 ;
        RECT 1.344 0.804 1.376 3.312 ;
  LAYER M3 ;
        RECT 1.344 3.26 1.376 3.292 ;
  LAYER M1 ;
        RECT 1.408 0.804 1.44 3.312 ;
  LAYER M3 ;
        RECT 1.408 0.824 1.44 0.856 ;
  LAYER M1 ;
        RECT 1.472 0.804 1.504 3.312 ;
  LAYER M3 ;
        RECT 1.472 3.26 1.504 3.292 ;
  LAYER M1 ;
        RECT 1.536 0.804 1.568 3.312 ;
  LAYER M3 ;
        RECT 1.536 0.824 1.568 0.856 ;
  LAYER M1 ;
        RECT 1.6 0.804 1.632 3.312 ;
  LAYER M3 ;
        RECT 1.6 3.26 1.632 3.292 ;
  LAYER M1 ;
        RECT 1.664 0.804 1.696 3.312 ;
  LAYER M3 ;
        RECT 1.664 0.824 1.696 0.856 ;
  LAYER M1 ;
        RECT 1.728 0.804 1.76 3.312 ;
  LAYER M3 ;
        RECT 1.728 3.26 1.76 3.292 ;
  LAYER M1 ;
        RECT 1.792 0.804 1.824 3.312 ;
  LAYER M3 ;
        RECT 1.792 0.824 1.824 0.856 ;
  LAYER M1 ;
        RECT 1.856 0.804 1.888 3.312 ;
  LAYER M3 ;
        RECT 1.856 3.26 1.888 3.292 ;
  LAYER M1 ;
        RECT 1.92 0.804 1.952 3.312 ;
  LAYER M3 ;
        RECT 1.92 0.824 1.952 0.856 ;
  LAYER M1 ;
        RECT 1.984 0.804 2.016 3.312 ;
  LAYER M3 ;
        RECT 1.984 3.26 2.016 3.292 ;
  LAYER M1 ;
        RECT 2.048 0.804 2.08 3.312 ;
  LAYER M3 ;
        RECT 2.048 0.824 2.08 0.856 ;
  LAYER M1 ;
        RECT 2.112 0.804 2.144 3.312 ;
  LAYER M3 ;
        RECT 2.112 3.26 2.144 3.292 ;
  LAYER M1 ;
        RECT 2.176 0.804 2.208 3.312 ;
  LAYER M3 ;
        RECT 2.176 0.824 2.208 0.856 ;
  LAYER M1 ;
        RECT 2.24 0.804 2.272 3.312 ;
  LAYER M3 ;
        RECT 2.24 3.26 2.272 3.292 ;
  LAYER M1 ;
        RECT 2.304 0.804 2.336 3.312 ;
  LAYER M3 ;
        RECT 2.304 0.824 2.336 0.856 ;
  LAYER M1 ;
        RECT 2.368 0.804 2.4 3.312 ;
  LAYER M3 ;
        RECT 2.368 3.26 2.4 3.292 ;
  LAYER M1 ;
        RECT 2.432 0.804 2.464 3.312 ;
  LAYER M3 ;
        RECT 2.432 0.824 2.464 0.856 ;
  LAYER M1 ;
        RECT 2.496 0.804 2.528 3.312 ;
  LAYER M3 ;
        RECT 2.496 3.26 2.528 3.292 ;
  LAYER M1 ;
        RECT 2.56 0.804 2.592 3.312 ;
  LAYER M3 ;
        RECT 2.56 0.824 2.592 0.856 ;
  LAYER M1 ;
        RECT 2.624 0.804 2.656 3.312 ;
  LAYER M3 ;
        RECT 2.624 3.26 2.656 3.292 ;
  LAYER M1 ;
        RECT 2.688 0.804 2.72 3.312 ;
  LAYER M3 ;
        RECT 2.688 0.824 2.72 0.856 ;
  LAYER M1 ;
        RECT 2.752 0.804 2.784 3.312 ;
  LAYER M3 ;
        RECT 2.752 3.26 2.784 3.292 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 3.312 ;
  LAYER M3 ;
        RECT 0.448 0.888 0.48 0.92 ;
  LAYER M2 ;
        RECT 2.816 0.952 2.848 0.984 ;
  LAYER M2 ;
        RECT 0.448 1.016 0.48 1.048 ;
  LAYER M2 ;
        RECT 2.816 1.08 2.848 1.112 ;
  LAYER M2 ;
        RECT 0.448 1.144 0.48 1.176 ;
  LAYER M2 ;
        RECT 2.816 1.208 2.848 1.24 ;
  LAYER M2 ;
        RECT 0.448 1.272 0.48 1.304 ;
  LAYER M2 ;
        RECT 2.816 1.336 2.848 1.368 ;
  LAYER M2 ;
        RECT 0.448 1.4 0.48 1.432 ;
  LAYER M2 ;
        RECT 2.816 1.464 2.848 1.496 ;
  LAYER M2 ;
        RECT 0.448 1.528 0.48 1.56 ;
  LAYER M2 ;
        RECT 2.816 1.592 2.848 1.624 ;
  LAYER M2 ;
        RECT 0.448 1.656 0.48 1.688 ;
  LAYER M2 ;
        RECT 2.816 1.72 2.848 1.752 ;
  LAYER M2 ;
        RECT 0.448 1.784 0.48 1.816 ;
  LAYER M2 ;
        RECT 2.816 1.848 2.848 1.88 ;
  LAYER M2 ;
        RECT 0.448 1.912 0.48 1.944 ;
  LAYER M2 ;
        RECT 2.816 1.976 2.848 2.008 ;
  LAYER M2 ;
        RECT 0.448 2.04 0.48 2.072 ;
  LAYER M2 ;
        RECT 2.816 2.104 2.848 2.136 ;
  LAYER M2 ;
        RECT 0.448 2.168 0.48 2.2 ;
  LAYER M2 ;
        RECT 2.816 2.232 2.848 2.264 ;
  LAYER M2 ;
        RECT 0.448 2.296 0.48 2.328 ;
  LAYER M2 ;
        RECT 2.816 2.36 2.848 2.392 ;
  LAYER M2 ;
        RECT 0.448 2.424 0.48 2.456 ;
  LAYER M2 ;
        RECT 2.816 2.488 2.848 2.52 ;
  LAYER M2 ;
        RECT 0.448 2.552 0.48 2.584 ;
  LAYER M2 ;
        RECT 2.816 2.616 2.848 2.648 ;
  LAYER M2 ;
        RECT 0.448 2.68 0.48 2.712 ;
  LAYER M2 ;
        RECT 2.816 2.744 2.848 2.776 ;
  LAYER M2 ;
        RECT 0.448 2.808 0.48 2.84 ;
  LAYER M2 ;
        RECT 2.816 2.872 2.848 2.904 ;
  LAYER M2 ;
        RECT 0.448 2.936 0.48 2.968 ;
  LAYER M2 ;
        RECT 2.816 3 2.848 3.032 ;
  LAYER M2 ;
        RECT 0.448 3.064 0.48 3.096 ;
  LAYER M2 ;
        RECT 2.816 3.128 2.848 3.16 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M1 ;
        RECT 0.448 3.912 0.48 6.42 ;
  LAYER M3 ;
        RECT 0.448 6.368 0.48 6.4 ;
  LAYER M1 ;
        RECT 0.512 3.912 0.544 6.42 ;
  LAYER M3 ;
        RECT 0.512 3.932 0.544 3.964 ;
  LAYER M1 ;
        RECT 0.576 3.912 0.608 6.42 ;
  LAYER M3 ;
        RECT 0.576 6.368 0.608 6.4 ;
  LAYER M1 ;
        RECT 0.64 3.912 0.672 6.42 ;
  LAYER M3 ;
        RECT 0.64 3.932 0.672 3.964 ;
  LAYER M1 ;
        RECT 0.704 3.912 0.736 6.42 ;
  LAYER M3 ;
        RECT 0.704 6.368 0.736 6.4 ;
  LAYER M1 ;
        RECT 0.768 3.912 0.8 6.42 ;
  LAYER M3 ;
        RECT 0.768 3.932 0.8 3.964 ;
  LAYER M1 ;
        RECT 0.832 3.912 0.864 6.42 ;
  LAYER M3 ;
        RECT 0.832 6.368 0.864 6.4 ;
  LAYER M1 ;
        RECT 0.896 3.912 0.928 6.42 ;
  LAYER M3 ;
        RECT 0.896 3.932 0.928 3.964 ;
  LAYER M1 ;
        RECT 0.96 3.912 0.992 6.42 ;
  LAYER M3 ;
        RECT 0.96 6.368 0.992 6.4 ;
  LAYER M1 ;
        RECT 1.024 3.912 1.056 6.42 ;
  LAYER M3 ;
        RECT 1.024 3.932 1.056 3.964 ;
  LAYER M1 ;
        RECT 1.088 3.912 1.12 6.42 ;
  LAYER M3 ;
        RECT 1.088 6.368 1.12 6.4 ;
  LAYER M1 ;
        RECT 1.152 3.912 1.184 6.42 ;
  LAYER M3 ;
        RECT 1.152 3.932 1.184 3.964 ;
  LAYER M1 ;
        RECT 1.216 3.912 1.248 6.42 ;
  LAYER M3 ;
        RECT 1.216 6.368 1.248 6.4 ;
  LAYER M1 ;
        RECT 1.28 3.912 1.312 6.42 ;
  LAYER M3 ;
        RECT 1.28 3.932 1.312 3.964 ;
  LAYER M1 ;
        RECT 1.344 3.912 1.376 6.42 ;
  LAYER M3 ;
        RECT 1.344 6.368 1.376 6.4 ;
  LAYER M1 ;
        RECT 1.408 3.912 1.44 6.42 ;
  LAYER M3 ;
        RECT 1.408 3.932 1.44 3.964 ;
  LAYER M1 ;
        RECT 1.472 3.912 1.504 6.42 ;
  LAYER M3 ;
        RECT 1.472 6.368 1.504 6.4 ;
  LAYER M1 ;
        RECT 1.536 3.912 1.568 6.42 ;
  LAYER M3 ;
        RECT 1.536 3.932 1.568 3.964 ;
  LAYER M1 ;
        RECT 1.6 3.912 1.632 6.42 ;
  LAYER M3 ;
        RECT 1.6 6.368 1.632 6.4 ;
  LAYER M1 ;
        RECT 1.664 3.912 1.696 6.42 ;
  LAYER M3 ;
        RECT 1.664 3.932 1.696 3.964 ;
  LAYER M1 ;
        RECT 1.728 3.912 1.76 6.42 ;
  LAYER M3 ;
        RECT 1.728 6.368 1.76 6.4 ;
  LAYER M1 ;
        RECT 1.792 3.912 1.824 6.42 ;
  LAYER M3 ;
        RECT 1.792 3.932 1.824 3.964 ;
  LAYER M1 ;
        RECT 1.856 3.912 1.888 6.42 ;
  LAYER M3 ;
        RECT 1.856 6.368 1.888 6.4 ;
  LAYER M1 ;
        RECT 1.92 3.912 1.952 6.42 ;
  LAYER M3 ;
        RECT 1.92 3.932 1.952 3.964 ;
  LAYER M1 ;
        RECT 1.984 3.912 2.016 6.42 ;
  LAYER M3 ;
        RECT 1.984 6.368 2.016 6.4 ;
  LAYER M1 ;
        RECT 2.048 3.912 2.08 6.42 ;
  LAYER M3 ;
        RECT 2.048 3.932 2.08 3.964 ;
  LAYER M1 ;
        RECT 2.112 3.912 2.144 6.42 ;
  LAYER M3 ;
        RECT 2.112 6.368 2.144 6.4 ;
  LAYER M1 ;
        RECT 2.176 3.912 2.208 6.42 ;
  LAYER M3 ;
        RECT 2.176 3.932 2.208 3.964 ;
  LAYER M1 ;
        RECT 2.24 3.912 2.272 6.42 ;
  LAYER M3 ;
        RECT 2.24 6.368 2.272 6.4 ;
  LAYER M1 ;
        RECT 2.304 3.912 2.336 6.42 ;
  LAYER M3 ;
        RECT 2.304 3.932 2.336 3.964 ;
  LAYER M1 ;
        RECT 2.368 3.912 2.4 6.42 ;
  LAYER M3 ;
        RECT 2.368 6.368 2.4 6.4 ;
  LAYER M1 ;
        RECT 2.432 3.912 2.464 6.42 ;
  LAYER M3 ;
        RECT 2.432 3.932 2.464 3.964 ;
  LAYER M1 ;
        RECT 2.496 3.912 2.528 6.42 ;
  LAYER M3 ;
        RECT 2.496 6.368 2.528 6.4 ;
  LAYER M1 ;
        RECT 2.56 3.912 2.592 6.42 ;
  LAYER M3 ;
        RECT 2.56 3.932 2.592 3.964 ;
  LAYER M1 ;
        RECT 2.624 3.912 2.656 6.42 ;
  LAYER M3 ;
        RECT 2.624 6.368 2.656 6.4 ;
  LAYER M1 ;
        RECT 2.688 3.912 2.72 6.42 ;
  LAYER M3 ;
        RECT 2.688 3.932 2.72 3.964 ;
  LAYER M1 ;
        RECT 2.752 3.912 2.784 6.42 ;
  LAYER M3 ;
        RECT 2.752 6.368 2.784 6.4 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 6.42 ;
  LAYER M3 ;
        RECT 0.448 3.996 0.48 4.028 ;
  LAYER M2 ;
        RECT 2.816 4.06 2.848 4.092 ;
  LAYER M2 ;
        RECT 0.448 4.124 0.48 4.156 ;
  LAYER M2 ;
        RECT 2.816 4.188 2.848 4.22 ;
  LAYER M2 ;
        RECT 0.448 4.252 0.48 4.284 ;
  LAYER M2 ;
        RECT 2.816 4.316 2.848 4.348 ;
  LAYER M2 ;
        RECT 0.448 4.38 0.48 4.412 ;
  LAYER M2 ;
        RECT 2.816 4.444 2.848 4.476 ;
  LAYER M2 ;
        RECT 0.448 4.508 0.48 4.54 ;
  LAYER M2 ;
        RECT 2.816 4.572 2.848 4.604 ;
  LAYER M2 ;
        RECT 0.448 4.636 0.48 4.668 ;
  LAYER M2 ;
        RECT 2.816 4.7 2.848 4.732 ;
  LAYER M2 ;
        RECT 0.448 4.764 0.48 4.796 ;
  LAYER M2 ;
        RECT 2.816 4.828 2.848 4.86 ;
  LAYER M2 ;
        RECT 0.448 4.892 0.48 4.924 ;
  LAYER M2 ;
        RECT 2.816 4.956 2.848 4.988 ;
  LAYER M2 ;
        RECT 0.448 5.02 0.48 5.052 ;
  LAYER M2 ;
        RECT 2.816 5.084 2.848 5.116 ;
  LAYER M2 ;
        RECT 0.448 5.148 0.48 5.18 ;
  LAYER M2 ;
        RECT 2.816 5.212 2.848 5.244 ;
  LAYER M2 ;
        RECT 0.448 5.276 0.48 5.308 ;
  LAYER M2 ;
        RECT 2.816 5.34 2.848 5.372 ;
  LAYER M2 ;
        RECT 0.448 5.404 0.48 5.436 ;
  LAYER M2 ;
        RECT 2.816 5.468 2.848 5.5 ;
  LAYER M2 ;
        RECT 0.448 5.532 0.48 5.564 ;
  LAYER M2 ;
        RECT 2.816 5.596 2.848 5.628 ;
  LAYER M2 ;
        RECT 0.448 5.66 0.48 5.692 ;
  LAYER M2 ;
        RECT 2.816 5.724 2.848 5.756 ;
  LAYER M2 ;
        RECT 0.448 5.788 0.48 5.82 ;
  LAYER M2 ;
        RECT 2.816 5.852 2.848 5.884 ;
  LAYER M2 ;
        RECT 0.448 5.916 0.48 5.948 ;
  LAYER M2 ;
        RECT 2.816 5.98 2.848 6.012 ;
  LAYER M2 ;
        RECT 0.448 6.044 0.48 6.076 ;
  LAYER M2 ;
        RECT 2.816 6.108 2.848 6.14 ;
  LAYER M2 ;
        RECT 0.448 6.172 0.48 6.204 ;
  LAYER M2 ;
        RECT 2.816 6.236 2.848 6.268 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M1 ;
        RECT 0.448 7.02 0.48 9.528 ;
  LAYER M3 ;
        RECT 0.448 9.476 0.48 9.508 ;
  LAYER M1 ;
        RECT 0.512 7.02 0.544 9.528 ;
  LAYER M3 ;
        RECT 0.512 7.04 0.544 7.072 ;
  LAYER M1 ;
        RECT 0.576 7.02 0.608 9.528 ;
  LAYER M3 ;
        RECT 0.576 9.476 0.608 9.508 ;
  LAYER M1 ;
        RECT 0.64 7.02 0.672 9.528 ;
  LAYER M3 ;
        RECT 0.64 7.04 0.672 7.072 ;
  LAYER M1 ;
        RECT 0.704 7.02 0.736 9.528 ;
  LAYER M3 ;
        RECT 0.704 9.476 0.736 9.508 ;
  LAYER M1 ;
        RECT 0.768 7.02 0.8 9.528 ;
  LAYER M3 ;
        RECT 0.768 7.04 0.8 7.072 ;
  LAYER M1 ;
        RECT 0.832 7.02 0.864 9.528 ;
  LAYER M3 ;
        RECT 0.832 9.476 0.864 9.508 ;
  LAYER M1 ;
        RECT 0.896 7.02 0.928 9.528 ;
  LAYER M3 ;
        RECT 0.896 7.04 0.928 7.072 ;
  LAYER M1 ;
        RECT 0.96 7.02 0.992 9.528 ;
  LAYER M3 ;
        RECT 0.96 9.476 0.992 9.508 ;
  LAYER M1 ;
        RECT 1.024 7.02 1.056 9.528 ;
  LAYER M3 ;
        RECT 1.024 7.04 1.056 7.072 ;
  LAYER M1 ;
        RECT 1.088 7.02 1.12 9.528 ;
  LAYER M3 ;
        RECT 1.088 9.476 1.12 9.508 ;
  LAYER M1 ;
        RECT 1.152 7.02 1.184 9.528 ;
  LAYER M3 ;
        RECT 1.152 7.04 1.184 7.072 ;
  LAYER M1 ;
        RECT 1.216 7.02 1.248 9.528 ;
  LAYER M3 ;
        RECT 1.216 9.476 1.248 9.508 ;
  LAYER M1 ;
        RECT 1.28 7.02 1.312 9.528 ;
  LAYER M3 ;
        RECT 1.28 7.04 1.312 7.072 ;
  LAYER M1 ;
        RECT 1.344 7.02 1.376 9.528 ;
  LAYER M3 ;
        RECT 1.344 9.476 1.376 9.508 ;
  LAYER M1 ;
        RECT 1.408 7.02 1.44 9.528 ;
  LAYER M3 ;
        RECT 1.408 7.04 1.44 7.072 ;
  LAYER M1 ;
        RECT 1.472 7.02 1.504 9.528 ;
  LAYER M3 ;
        RECT 1.472 9.476 1.504 9.508 ;
  LAYER M1 ;
        RECT 1.536 7.02 1.568 9.528 ;
  LAYER M3 ;
        RECT 1.536 7.04 1.568 7.072 ;
  LAYER M1 ;
        RECT 1.6 7.02 1.632 9.528 ;
  LAYER M3 ;
        RECT 1.6 9.476 1.632 9.508 ;
  LAYER M1 ;
        RECT 1.664 7.02 1.696 9.528 ;
  LAYER M3 ;
        RECT 1.664 7.04 1.696 7.072 ;
  LAYER M1 ;
        RECT 1.728 7.02 1.76 9.528 ;
  LAYER M3 ;
        RECT 1.728 9.476 1.76 9.508 ;
  LAYER M1 ;
        RECT 1.792 7.02 1.824 9.528 ;
  LAYER M3 ;
        RECT 1.792 7.04 1.824 7.072 ;
  LAYER M1 ;
        RECT 1.856 7.02 1.888 9.528 ;
  LAYER M3 ;
        RECT 1.856 9.476 1.888 9.508 ;
  LAYER M1 ;
        RECT 1.92 7.02 1.952 9.528 ;
  LAYER M3 ;
        RECT 1.92 7.04 1.952 7.072 ;
  LAYER M1 ;
        RECT 1.984 7.02 2.016 9.528 ;
  LAYER M3 ;
        RECT 1.984 9.476 2.016 9.508 ;
  LAYER M1 ;
        RECT 2.048 7.02 2.08 9.528 ;
  LAYER M3 ;
        RECT 2.048 7.04 2.08 7.072 ;
  LAYER M1 ;
        RECT 2.112 7.02 2.144 9.528 ;
  LAYER M3 ;
        RECT 2.112 9.476 2.144 9.508 ;
  LAYER M1 ;
        RECT 2.176 7.02 2.208 9.528 ;
  LAYER M3 ;
        RECT 2.176 7.04 2.208 7.072 ;
  LAYER M1 ;
        RECT 2.24 7.02 2.272 9.528 ;
  LAYER M3 ;
        RECT 2.24 9.476 2.272 9.508 ;
  LAYER M1 ;
        RECT 2.304 7.02 2.336 9.528 ;
  LAYER M3 ;
        RECT 2.304 7.04 2.336 7.072 ;
  LAYER M1 ;
        RECT 2.368 7.02 2.4 9.528 ;
  LAYER M3 ;
        RECT 2.368 9.476 2.4 9.508 ;
  LAYER M1 ;
        RECT 2.432 7.02 2.464 9.528 ;
  LAYER M3 ;
        RECT 2.432 7.04 2.464 7.072 ;
  LAYER M1 ;
        RECT 2.496 7.02 2.528 9.528 ;
  LAYER M3 ;
        RECT 2.496 9.476 2.528 9.508 ;
  LAYER M1 ;
        RECT 2.56 7.02 2.592 9.528 ;
  LAYER M3 ;
        RECT 2.56 7.04 2.592 7.072 ;
  LAYER M1 ;
        RECT 2.624 7.02 2.656 9.528 ;
  LAYER M3 ;
        RECT 2.624 9.476 2.656 9.508 ;
  LAYER M1 ;
        RECT 2.688 7.02 2.72 9.528 ;
  LAYER M3 ;
        RECT 2.688 7.04 2.72 7.072 ;
  LAYER M1 ;
        RECT 2.752 7.02 2.784 9.528 ;
  LAYER M3 ;
        RECT 2.752 9.476 2.784 9.508 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 9.528 ;
  LAYER M3 ;
        RECT 0.448 7.104 0.48 7.136 ;
  LAYER M2 ;
        RECT 2.816 7.168 2.848 7.2 ;
  LAYER M2 ;
        RECT 0.448 7.232 0.48 7.264 ;
  LAYER M2 ;
        RECT 2.816 7.296 2.848 7.328 ;
  LAYER M2 ;
        RECT 0.448 7.36 0.48 7.392 ;
  LAYER M2 ;
        RECT 2.816 7.424 2.848 7.456 ;
  LAYER M2 ;
        RECT 0.448 7.488 0.48 7.52 ;
  LAYER M2 ;
        RECT 2.816 7.552 2.848 7.584 ;
  LAYER M2 ;
        RECT 0.448 7.616 0.48 7.648 ;
  LAYER M2 ;
        RECT 2.816 7.68 2.848 7.712 ;
  LAYER M2 ;
        RECT 0.448 7.744 0.48 7.776 ;
  LAYER M2 ;
        RECT 2.816 7.808 2.848 7.84 ;
  LAYER M2 ;
        RECT 0.448 7.872 0.48 7.904 ;
  LAYER M2 ;
        RECT 2.816 7.936 2.848 7.968 ;
  LAYER M2 ;
        RECT 0.448 8 0.48 8.032 ;
  LAYER M2 ;
        RECT 2.816 8.064 2.848 8.096 ;
  LAYER M2 ;
        RECT 0.448 8.128 0.48 8.16 ;
  LAYER M2 ;
        RECT 2.816 8.192 2.848 8.224 ;
  LAYER M2 ;
        RECT 0.448 8.256 0.48 8.288 ;
  LAYER M2 ;
        RECT 2.816 8.32 2.848 8.352 ;
  LAYER M2 ;
        RECT 0.448 8.384 0.48 8.416 ;
  LAYER M2 ;
        RECT 2.816 8.448 2.848 8.48 ;
  LAYER M2 ;
        RECT 0.448 8.512 0.48 8.544 ;
  LAYER M2 ;
        RECT 2.816 8.576 2.848 8.608 ;
  LAYER M2 ;
        RECT 0.448 8.64 0.48 8.672 ;
  LAYER M2 ;
        RECT 2.816 8.704 2.848 8.736 ;
  LAYER M2 ;
        RECT 0.448 8.768 0.48 8.8 ;
  LAYER M2 ;
        RECT 2.816 8.832 2.848 8.864 ;
  LAYER M2 ;
        RECT 0.448 8.896 0.48 8.928 ;
  LAYER M2 ;
        RECT 2.816 8.96 2.848 8.992 ;
  LAYER M2 ;
        RECT 0.448 9.024 0.48 9.056 ;
  LAYER M2 ;
        RECT 2.816 9.088 2.848 9.12 ;
  LAYER M2 ;
        RECT 0.448 9.152 0.48 9.184 ;
  LAYER M2 ;
        RECT 2.816 9.216 2.848 9.248 ;
  LAYER M2 ;
        RECT 0.448 9.28 0.48 9.312 ;
  LAYER M2 ;
        RECT 2.816 9.344 2.848 9.376 ;
  LAYER M2 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M1 ;
        RECT 0.448 10.128 0.48 12.636 ;
  LAYER M3 ;
        RECT 0.448 12.584 0.48 12.616 ;
  LAYER M1 ;
        RECT 0.512 10.128 0.544 12.636 ;
  LAYER M3 ;
        RECT 0.512 10.148 0.544 10.18 ;
  LAYER M1 ;
        RECT 0.576 10.128 0.608 12.636 ;
  LAYER M3 ;
        RECT 0.576 12.584 0.608 12.616 ;
  LAYER M1 ;
        RECT 0.64 10.128 0.672 12.636 ;
  LAYER M3 ;
        RECT 0.64 10.148 0.672 10.18 ;
  LAYER M1 ;
        RECT 0.704 10.128 0.736 12.636 ;
  LAYER M3 ;
        RECT 0.704 12.584 0.736 12.616 ;
  LAYER M1 ;
        RECT 0.768 10.128 0.8 12.636 ;
  LAYER M3 ;
        RECT 0.768 10.148 0.8 10.18 ;
  LAYER M1 ;
        RECT 0.832 10.128 0.864 12.636 ;
  LAYER M3 ;
        RECT 0.832 12.584 0.864 12.616 ;
  LAYER M1 ;
        RECT 0.896 10.128 0.928 12.636 ;
  LAYER M3 ;
        RECT 0.896 10.148 0.928 10.18 ;
  LAYER M1 ;
        RECT 0.96 10.128 0.992 12.636 ;
  LAYER M3 ;
        RECT 0.96 12.584 0.992 12.616 ;
  LAYER M1 ;
        RECT 1.024 10.128 1.056 12.636 ;
  LAYER M3 ;
        RECT 1.024 10.148 1.056 10.18 ;
  LAYER M1 ;
        RECT 1.088 10.128 1.12 12.636 ;
  LAYER M3 ;
        RECT 1.088 12.584 1.12 12.616 ;
  LAYER M1 ;
        RECT 1.152 10.128 1.184 12.636 ;
  LAYER M3 ;
        RECT 1.152 10.148 1.184 10.18 ;
  LAYER M1 ;
        RECT 1.216 10.128 1.248 12.636 ;
  LAYER M3 ;
        RECT 1.216 12.584 1.248 12.616 ;
  LAYER M1 ;
        RECT 1.28 10.128 1.312 12.636 ;
  LAYER M3 ;
        RECT 1.28 10.148 1.312 10.18 ;
  LAYER M1 ;
        RECT 1.344 10.128 1.376 12.636 ;
  LAYER M3 ;
        RECT 1.344 12.584 1.376 12.616 ;
  LAYER M1 ;
        RECT 1.408 10.128 1.44 12.636 ;
  LAYER M3 ;
        RECT 1.408 10.148 1.44 10.18 ;
  LAYER M1 ;
        RECT 1.472 10.128 1.504 12.636 ;
  LAYER M3 ;
        RECT 1.472 12.584 1.504 12.616 ;
  LAYER M1 ;
        RECT 1.536 10.128 1.568 12.636 ;
  LAYER M3 ;
        RECT 1.536 10.148 1.568 10.18 ;
  LAYER M1 ;
        RECT 1.6 10.128 1.632 12.636 ;
  LAYER M3 ;
        RECT 1.6 12.584 1.632 12.616 ;
  LAYER M1 ;
        RECT 1.664 10.128 1.696 12.636 ;
  LAYER M3 ;
        RECT 1.664 10.148 1.696 10.18 ;
  LAYER M1 ;
        RECT 1.728 10.128 1.76 12.636 ;
  LAYER M3 ;
        RECT 1.728 12.584 1.76 12.616 ;
  LAYER M1 ;
        RECT 1.792 10.128 1.824 12.636 ;
  LAYER M3 ;
        RECT 1.792 10.148 1.824 10.18 ;
  LAYER M1 ;
        RECT 1.856 10.128 1.888 12.636 ;
  LAYER M3 ;
        RECT 1.856 12.584 1.888 12.616 ;
  LAYER M1 ;
        RECT 1.92 10.128 1.952 12.636 ;
  LAYER M3 ;
        RECT 1.92 10.148 1.952 10.18 ;
  LAYER M1 ;
        RECT 1.984 10.128 2.016 12.636 ;
  LAYER M3 ;
        RECT 1.984 12.584 2.016 12.616 ;
  LAYER M1 ;
        RECT 2.048 10.128 2.08 12.636 ;
  LAYER M3 ;
        RECT 2.048 10.148 2.08 10.18 ;
  LAYER M1 ;
        RECT 2.112 10.128 2.144 12.636 ;
  LAYER M3 ;
        RECT 2.112 12.584 2.144 12.616 ;
  LAYER M1 ;
        RECT 2.176 10.128 2.208 12.636 ;
  LAYER M3 ;
        RECT 2.176 10.148 2.208 10.18 ;
  LAYER M1 ;
        RECT 2.24 10.128 2.272 12.636 ;
  LAYER M3 ;
        RECT 2.24 12.584 2.272 12.616 ;
  LAYER M1 ;
        RECT 2.304 10.128 2.336 12.636 ;
  LAYER M3 ;
        RECT 2.304 10.148 2.336 10.18 ;
  LAYER M1 ;
        RECT 2.368 10.128 2.4 12.636 ;
  LAYER M3 ;
        RECT 2.368 12.584 2.4 12.616 ;
  LAYER M1 ;
        RECT 2.432 10.128 2.464 12.636 ;
  LAYER M3 ;
        RECT 2.432 10.148 2.464 10.18 ;
  LAYER M1 ;
        RECT 2.496 10.128 2.528 12.636 ;
  LAYER M3 ;
        RECT 2.496 12.584 2.528 12.616 ;
  LAYER M1 ;
        RECT 2.56 10.128 2.592 12.636 ;
  LAYER M3 ;
        RECT 2.56 10.148 2.592 10.18 ;
  LAYER M1 ;
        RECT 2.624 10.128 2.656 12.636 ;
  LAYER M3 ;
        RECT 2.624 12.584 2.656 12.616 ;
  LAYER M1 ;
        RECT 2.688 10.128 2.72 12.636 ;
  LAYER M3 ;
        RECT 2.688 10.148 2.72 10.18 ;
  LAYER M1 ;
        RECT 2.752 10.128 2.784 12.636 ;
  LAYER M3 ;
        RECT 2.752 12.584 2.784 12.616 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 12.636 ;
  LAYER M3 ;
        RECT 0.448 10.212 0.48 10.244 ;
  LAYER M2 ;
        RECT 2.816 10.276 2.848 10.308 ;
  LAYER M2 ;
        RECT 0.448 10.34 0.48 10.372 ;
  LAYER M2 ;
        RECT 2.816 10.404 2.848 10.436 ;
  LAYER M2 ;
        RECT 0.448 10.468 0.48 10.5 ;
  LAYER M2 ;
        RECT 2.816 10.532 2.848 10.564 ;
  LAYER M2 ;
        RECT 0.448 10.596 0.48 10.628 ;
  LAYER M2 ;
        RECT 2.816 10.66 2.848 10.692 ;
  LAYER M2 ;
        RECT 0.448 10.724 0.48 10.756 ;
  LAYER M2 ;
        RECT 2.816 10.788 2.848 10.82 ;
  LAYER M2 ;
        RECT 0.448 10.852 0.48 10.884 ;
  LAYER M2 ;
        RECT 2.816 10.916 2.848 10.948 ;
  LAYER M2 ;
        RECT 0.448 10.98 0.48 11.012 ;
  LAYER M2 ;
        RECT 2.816 11.044 2.848 11.076 ;
  LAYER M2 ;
        RECT 0.448 11.108 0.48 11.14 ;
  LAYER M2 ;
        RECT 2.816 11.172 2.848 11.204 ;
  LAYER M2 ;
        RECT 0.448 11.236 0.48 11.268 ;
  LAYER M2 ;
        RECT 2.816 11.3 2.848 11.332 ;
  LAYER M2 ;
        RECT 0.448 11.364 0.48 11.396 ;
  LAYER M2 ;
        RECT 2.816 11.428 2.848 11.46 ;
  LAYER M2 ;
        RECT 0.448 11.492 0.48 11.524 ;
  LAYER M2 ;
        RECT 2.816 11.556 2.848 11.588 ;
  LAYER M2 ;
        RECT 0.448 11.62 0.48 11.652 ;
  LAYER M2 ;
        RECT 2.816 11.684 2.848 11.716 ;
  LAYER M2 ;
        RECT 0.448 11.748 0.48 11.78 ;
  LAYER M2 ;
        RECT 2.816 11.812 2.848 11.844 ;
  LAYER M2 ;
        RECT 0.448 11.876 0.48 11.908 ;
  LAYER M2 ;
        RECT 2.816 11.94 2.848 11.972 ;
  LAYER M2 ;
        RECT 0.448 12.004 0.48 12.036 ;
  LAYER M2 ;
        RECT 2.816 12.068 2.848 12.1 ;
  LAYER M2 ;
        RECT 0.448 12.132 0.48 12.164 ;
  LAYER M2 ;
        RECT 2.816 12.196 2.848 12.228 ;
  LAYER M2 ;
        RECT 0.448 12.26 0.48 12.292 ;
  LAYER M2 ;
        RECT 2.816 12.324 2.848 12.356 ;
  LAYER M2 ;
        RECT 0.448 12.388 0.48 12.42 ;
  LAYER M2 ;
        RECT 2.816 12.452 2.848 12.484 ;
  LAYER M2 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M1 ;
        RECT 0.448 13.236 0.48 15.744 ;
  LAYER M3 ;
        RECT 0.448 15.692 0.48 15.724 ;
  LAYER M1 ;
        RECT 0.512 13.236 0.544 15.744 ;
  LAYER M3 ;
        RECT 0.512 13.256 0.544 13.288 ;
  LAYER M1 ;
        RECT 0.576 13.236 0.608 15.744 ;
  LAYER M3 ;
        RECT 0.576 15.692 0.608 15.724 ;
  LAYER M1 ;
        RECT 0.64 13.236 0.672 15.744 ;
  LAYER M3 ;
        RECT 0.64 13.256 0.672 13.288 ;
  LAYER M1 ;
        RECT 0.704 13.236 0.736 15.744 ;
  LAYER M3 ;
        RECT 0.704 15.692 0.736 15.724 ;
  LAYER M1 ;
        RECT 0.768 13.236 0.8 15.744 ;
  LAYER M3 ;
        RECT 0.768 13.256 0.8 13.288 ;
  LAYER M1 ;
        RECT 0.832 13.236 0.864 15.744 ;
  LAYER M3 ;
        RECT 0.832 15.692 0.864 15.724 ;
  LAYER M1 ;
        RECT 0.896 13.236 0.928 15.744 ;
  LAYER M3 ;
        RECT 0.896 13.256 0.928 13.288 ;
  LAYER M1 ;
        RECT 0.96 13.236 0.992 15.744 ;
  LAYER M3 ;
        RECT 0.96 15.692 0.992 15.724 ;
  LAYER M1 ;
        RECT 1.024 13.236 1.056 15.744 ;
  LAYER M3 ;
        RECT 1.024 13.256 1.056 13.288 ;
  LAYER M1 ;
        RECT 1.088 13.236 1.12 15.744 ;
  LAYER M3 ;
        RECT 1.088 15.692 1.12 15.724 ;
  LAYER M1 ;
        RECT 1.152 13.236 1.184 15.744 ;
  LAYER M3 ;
        RECT 1.152 13.256 1.184 13.288 ;
  LAYER M1 ;
        RECT 1.216 13.236 1.248 15.744 ;
  LAYER M3 ;
        RECT 1.216 15.692 1.248 15.724 ;
  LAYER M1 ;
        RECT 1.28 13.236 1.312 15.744 ;
  LAYER M3 ;
        RECT 1.28 13.256 1.312 13.288 ;
  LAYER M1 ;
        RECT 1.344 13.236 1.376 15.744 ;
  LAYER M3 ;
        RECT 1.344 15.692 1.376 15.724 ;
  LAYER M1 ;
        RECT 1.408 13.236 1.44 15.744 ;
  LAYER M3 ;
        RECT 1.408 13.256 1.44 13.288 ;
  LAYER M1 ;
        RECT 1.472 13.236 1.504 15.744 ;
  LAYER M3 ;
        RECT 1.472 15.692 1.504 15.724 ;
  LAYER M1 ;
        RECT 1.536 13.236 1.568 15.744 ;
  LAYER M3 ;
        RECT 1.536 13.256 1.568 13.288 ;
  LAYER M1 ;
        RECT 1.6 13.236 1.632 15.744 ;
  LAYER M3 ;
        RECT 1.6 15.692 1.632 15.724 ;
  LAYER M1 ;
        RECT 1.664 13.236 1.696 15.744 ;
  LAYER M3 ;
        RECT 1.664 13.256 1.696 13.288 ;
  LAYER M1 ;
        RECT 1.728 13.236 1.76 15.744 ;
  LAYER M3 ;
        RECT 1.728 15.692 1.76 15.724 ;
  LAYER M1 ;
        RECT 1.792 13.236 1.824 15.744 ;
  LAYER M3 ;
        RECT 1.792 13.256 1.824 13.288 ;
  LAYER M1 ;
        RECT 1.856 13.236 1.888 15.744 ;
  LAYER M3 ;
        RECT 1.856 15.692 1.888 15.724 ;
  LAYER M1 ;
        RECT 1.92 13.236 1.952 15.744 ;
  LAYER M3 ;
        RECT 1.92 13.256 1.952 13.288 ;
  LAYER M1 ;
        RECT 1.984 13.236 2.016 15.744 ;
  LAYER M3 ;
        RECT 1.984 15.692 2.016 15.724 ;
  LAYER M1 ;
        RECT 2.048 13.236 2.08 15.744 ;
  LAYER M3 ;
        RECT 2.048 13.256 2.08 13.288 ;
  LAYER M1 ;
        RECT 2.112 13.236 2.144 15.744 ;
  LAYER M3 ;
        RECT 2.112 15.692 2.144 15.724 ;
  LAYER M1 ;
        RECT 2.176 13.236 2.208 15.744 ;
  LAYER M3 ;
        RECT 2.176 13.256 2.208 13.288 ;
  LAYER M1 ;
        RECT 2.24 13.236 2.272 15.744 ;
  LAYER M3 ;
        RECT 2.24 15.692 2.272 15.724 ;
  LAYER M1 ;
        RECT 2.304 13.236 2.336 15.744 ;
  LAYER M3 ;
        RECT 2.304 13.256 2.336 13.288 ;
  LAYER M1 ;
        RECT 2.368 13.236 2.4 15.744 ;
  LAYER M3 ;
        RECT 2.368 15.692 2.4 15.724 ;
  LAYER M1 ;
        RECT 2.432 13.236 2.464 15.744 ;
  LAYER M3 ;
        RECT 2.432 13.256 2.464 13.288 ;
  LAYER M1 ;
        RECT 2.496 13.236 2.528 15.744 ;
  LAYER M3 ;
        RECT 2.496 15.692 2.528 15.724 ;
  LAYER M1 ;
        RECT 2.56 13.236 2.592 15.744 ;
  LAYER M3 ;
        RECT 2.56 13.256 2.592 13.288 ;
  LAYER M1 ;
        RECT 2.624 13.236 2.656 15.744 ;
  LAYER M3 ;
        RECT 2.624 15.692 2.656 15.724 ;
  LAYER M1 ;
        RECT 2.688 13.236 2.72 15.744 ;
  LAYER M3 ;
        RECT 2.688 13.256 2.72 13.288 ;
  LAYER M1 ;
        RECT 2.752 13.236 2.784 15.744 ;
  LAYER M3 ;
        RECT 2.752 15.692 2.784 15.724 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 15.744 ;
  LAYER M3 ;
        RECT 0.448 13.32 0.48 13.352 ;
  LAYER M2 ;
        RECT 2.816 13.384 2.848 13.416 ;
  LAYER M2 ;
        RECT 0.448 13.448 0.48 13.48 ;
  LAYER M2 ;
        RECT 2.816 13.512 2.848 13.544 ;
  LAYER M2 ;
        RECT 0.448 13.576 0.48 13.608 ;
  LAYER M2 ;
        RECT 2.816 13.64 2.848 13.672 ;
  LAYER M2 ;
        RECT 0.448 13.704 0.48 13.736 ;
  LAYER M2 ;
        RECT 2.816 13.768 2.848 13.8 ;
  LAYER M2 ;
        RECT 0.448 13.832 0.48 13.864 ;
  LAYER M2 ;
        RECT 2.816 13.896 2.848 13.928 ;
  LAYER M2 ;
        RECT 0.448 13.96 0.48 13.992 ;
  LAYER M2 ;
        RECT 2.816 14.024 2.848 14.056 ;
  LAYER M2 ;
        RECT 0.448 14.088 0.48 14.12 ;
  LAYER M2 ;
        RECT 2.816 14.152 2.848 14.184 ;
  LAYER M2 ;
        RECT 0.448 14.216 0.48 14.248 ;
  LAYER M2 ;
        RECT 2.816 14.28 2.848 14.312 ;
  LAYER M2 ;
        RECT 0.448 14.344 0.48 14.376 ;
  LAYER M2 ;
        RECT 2.816 14.408 2.848 14.44 ;
  LAYER M2 ;
        RECT 0.448 14.472 0.48 14.504 ;
  LAYER M2 ;
        RECT 2.816 14.536 2.848 14.568 ;
  LAYER M2 ;
        RECT 0.448 14.6 0.48 14.632 ;
  LAYER M2 ;
        RECT 2.816 14.664 2.848 14.696 ;
  LAYER M2 ;
        RECT 0.448 14.728 0.48 14.76 ;
  LAYER M2 ;
        RECT 2.816 14.792 2.848 14.824 ;
  LAYER M2 ;
        RECT 0.448 14.856 0.48 14.888 ;
  LAYER M2 ;
        RECT 2.816 14.92 2.848 14.952 ;
  LAYER M2 ;
        RECT 0.448 14.984 0.48 15.016 ;
  LAYER M2 ;
        RECT 2.816 15.048 2.848 15.08 ;
  LAYER M2 ;
        RECT 0.448 15.112 0.48 15.144 ;
  LAYER M2 ;
        RECT 2.816 15.176 2.848 15.208 ;
  LAYER M2 ;
        RECT 0.448 15.24 0.48 15.272 ;
  LAYER M2 ;
        RECT 2.816 15.304 2.848 15.336 ;
  LAYER M2 ;
        RECT 0.448 15.368 0.48 15.4 ;
  LAYER M2 ;
        RECT 2.816 15.432 2.848 15.464 ;
  LAYER M2 ;
        RECT 0.448 15.496 0.48 15.528 ;
  LAYER M2 ;
        RECT 2.816 15.56 2.848 15.592 ;
  LAYER M2 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M1 ;
        RECT 0.448 16.344 0.48 18.852 ;
  LAYER M3 ;
        RECT 0.448 18.8 0.48 18.832 ;
  LAYER M1 ;
        RECT 0.512 16.344 0.544 18.852 ;
  LAYER M3 ;
        RECT 0.512 16.364 0.544 16.396 ;
  LAYER M1 ;
        RECT 0.576 16.344 0.608 18.852 ;
  LAYER M3 ;
        RECT 0.576 18.8 0.608 18.832 ;
  LAYER M1 ;
        RECT 0.64 16.344 0.672 18.852 ;
  LAYER M3 ;
        RECT 0.64 16.364 0.672 16.396 ;
  LAYER M1 ;
        RECT 0.704 16.344 0.736 18.852 ;
  LAYER M3 ;
        RECT 0.704 18.8 0.736 18.832 ;
  LAYER M1 ;
        RECT 0.768 16.344 0.8 18.852 ;
  LAYER M3 ;
        RECT 0.768 16.364 0.8 16.396 ;
  LAYER M1 ;
        RECT 0.832 16.344 0.864 18.852 ;
  LAYER M3 ;
        RECT 0.832 18.8 0.864 18.832 ;
  LAYER M1 ;
        RECT 0.896 16.344 0.928 18.852 ;
  LAYER M3 ;
        RECT 0.896 16.364 0.928 16.396 ;
  LAYER M1 ;
        RECT 0.96 16.344 0.992 18.852 ;
  LAYER M3 ;
        RECT 0.96 18.8 0.992 18.832 ;
  LAYER M1 ;
        RECT 1.024 16.344 1.056 18.852 ;
  LAYER M3 ;
        RECT 1.024 16.364 1.056 16.396 ;
  LAYER M1 ;
        RECT 1.088 16.344 1.12 18.852 ;
  LAYER M3 ;
        RECT 1.088 18.8 1.12 18.832 ;
  LAYER M1 ;
        RECT 1.152 16.344 1.184 18.852 ;
  LAYER M3 ;
        RECT 1.152 16.364 1.184 16.396 ;
  LAYER M1 ;
        RECT 1.216 16.344 1.248 18.852 ;
  LAYER M3 ;
        RECT 1.216 18.8 1.248 18.832 ;
  LAYER M1 ;
        RECT 1.28 16.344 1.312 18.852 ;
  LAYER M3 ;
        RECT 1.28 16.364 1.312 16.396 ;
  LAYER M1 ;
        RECT 1.344 16.344 1.376 18.852 ;
  LAYER M3 ;
        RECT 1.344 18.8 1.376 18.832 ;
  LAYER M1 ;
        RECT 1.408 16.344 1.44 18.852 ;
  LAYER M3 ;
        RECT 1.408 16.364 1.44 16.396 ;
  LAYER M1 ;
        RECT 1.472 16.344 1.504 18.852 ;
  LAYER M3 ;
        RECT 1.472 18.8 1.504 18.832 ;
  LAYER M1 ;
        RECT 1.536 16.344 1.568 18.852 ;
  LAYER M3 ;
        RECT 1.536 16.364 1.568 16.396 ;
  LAYER M1 ;
        RECT 1.6 16.344 1.632 18.852 ;
  LAYER M3 ;
        RECT 1.6 18.8 1.632 18.832 ;
  LAYER M1 ;
        RECT 1.664 16.344 1.696 18.852 ;
  LAYER M3 ;
        RECT 1.664 16.364 1.696 16.396 ;
  LAYER M1 ;
        RECT 1.728 16.344 1.76 18.852 ;
  LAYER M3 ;
        RECT 1.728 18.8 1.76 18.832 ;
  LAYER M1 ;
        RECT 1.792 16.344 1.824 18.852 ;
  LAYER M3 ;
        RECT 1.792 16.364 1.824 16.396 ;
  LAYER M1 ;
        RECT 1.856 16.344 1.888 18.852 ;
  LAYER M3 ;
        RECT 1.856 18.8 1.888 18.832 ;
  LAYER M1 ;
        RECT 1.92 16.344 1.952 18.852 ;
  LAYER M3 ;
        RECT 1.92 16.364 1.952 16.396 ;
  LAYER M1 ;
        RECT 1.984 16.344 2.016 18.852 ;
  LAYER M3 ;
        RECT 1.984 18.8 2.016 18.832 ;
  LAYER M1 ;
        RECT 2.048 16.344 2.08 18.852 ;
  LAYER M3 ;
        RECT 2.048 16.364 2.08 16.396 ;
  LAYER M1 ;
        RECT 2.112 16.344 2.144 18.852 ;
  LAYER M3 ;
        RECT 2.112 18.8 2.144 18.832 ;
  LAYER M1 ;
        RECT 2.176 16.344 2.208 18.852 ;
  LAYER M3 ;
        RECT 2.176 16.364 2.208 16.396 ;
  LAYER M1 ;
        RECT 2.24 16.344 2.272 18.852 ;
  LAYER M3 ;
        RECT 2.24 18.8 2.272 18.832 ;
  LAYER M1 ;
        RECT 2.304 16.344 2.336 18.852 ;
  LAYER M3 ;
        RECT 2.304 16.364 2.336 16.396 ;
  LAYER M1 ;
        RECT 2.368 16.344 2.4 18.852 ;
  LAYER M3 ;
        RECT 2.368 18.8 2.4 18.832 ;
  LAYER M1 ;
        RECT 2.432 16.344 2.464 18.852 ;
  LAYER M3 ;
        RECT 2.432 16.364 2.464 16.396 ;
  LAYER M1 ;
        RECT 2.496 16.344 2.528 18.852 ;
  LAYER M3 ;
        RECT 2.496 18.8 2.528 18.832 ;
  LAYER M1 ;
        RECT 2.56 16.344 2.592 18.852 ;
  LAYER M3 ;
        RECT 2.56 16.364 2.592 16.396 ;
  LAYER M1 ;
        RECT 2.624 16.344 2.656 18.852 ;
  LAYER M3 ;
        RECT 2.624 18.8 2.656 18.832 ;
  LAYER M1 ;
        RECT 2.688 16.344 2.72 18.852 ;
  LAYER M3 ;
        RECT 2.688 16.364 2.72 16.396 ;
  LAYER M1 ;
        RECT 2.752 16.344 2.784 18.852 ;
  LAYER M3 ;
        RECT 2.752 18.8 2.784 18.832 ;
  LAYER M1 ;
        RECT 2.816 16.344 2.848 18.852 ;
  LAYER M3 ;
        RECT 0.448 16.428 0.48 16.46 ;
  LAYER M2 ;
        RECT 2.816 16.492 2.848 16.524 ;
  LAYER M2 ;
        RECT 0.448 16.556 0.48 16.588 ;
  LAYER M2 ;
        RECT 2.816 16.62 2.848 16.652 ;
  LAYER M2 ;
        RECT 0.448 16.684 0.48 16.716 ;
  LAYER M2 ;
        RECT 2.816 16.748 2.848 16.78 ;
  LAYER M2 ;
        RECT 0.448 16.812 0.48 16.844 ;
  LAYER M2 ;
        RECT 2.816 16.876 2.848 16.908 ;
  LAYER M2 ;
        RECT 0.448 16.94 0.48 16.972 ;
  LAYER M2 ;
        RECT 2.816 17.004 2.848 17.036 ;
  LAYER M2 ;
        RECT 0.448 17.068 0.48 17.1 ;
  LAYER M2 ;
        RECT 2.816 17.132 2.848 17.164 ;
  LAYER M2 ;
        RECT 0.448 17.196 0.48 17.228 ;
  LAYER M2 ;
        RECT 2.816 17.26 2.848 17.292 ;
  LAYER M2 ;
        RECT 0.448 17.324 0.48 17.356 ;
  LAYER M2 ;
        RECT 2.816 17.388 2.848 17.42 ;
  LAYER M2 ;
        RECT 0.448 17.452 0.48 17.484 ;
  LAYER M2 ;
        RECT 2.816 17.516 2.848 17.548 ;
  LAYER M2 ;
        RECT 0.448 17.58 0.48 17.612 ;
  LAYER M2 ;
        RECT 2.816 17.644 2.848 17.676 ;
  LAYER M2 ;
        RECT 0.448 17.708 0.48 17.74 ;
  LAYER M2 ;
        RECT 2.816 17.772 2.848 17.804 ;
  LAYER M2 ;
        RECT 0.448 17.836 0.48 17.868 ;
  LAYER M2 ;
        RECT 2.816 17.9 2.848 17.932 ;
  LAYER M2 ;
        RECT 0.448 17.964 0.48 17.996 ;
  LAYER M2 ;
        RECT 2.816 18.028 2.848 18.06 ;
  LAYER M2 ;
        RECT 0.448 18.092 0.48 18.124 ;
  LAYER M2 ;
        RECT 2.816 18.156 2.848 18.188 ;
  LAYER M2 ;
        RECT 0.448 18.22 0.48 18.252 ;
  LAYER M2 ;
        RECT 2.816 18.284 2.848 18.316 ;
  LAYER M2 ;
        RECT 0.448 18.348 0.48 18.38 ;
  LAYER M2 ;
        RECT 2.816 18.412 2.848 18.444 ;
  LAYER M2 ;
        RECT 0.448 18.476 0.48 18.508 ;
  LAYER M2 ;
        RECT 2.816 18.54 2.848 18.572 ;
  LAYER M2 ;
        RECT 0.448 18.604 0.48 18.636 ;
  LAYER M2 ;
        RECT 2.816 18.668 2.848 18.7 ;
  LAYER M2 ;
        RECT 0.4 16.296 2.896 18.9 ;
  LAYER M1 ;
        RECT 0.448 19.452 0.48 21.96 ;
  LAYER M3 ;
        RECT 0.448 21.908 0.48 21.94 ;
  LAYER M1 ;
        RECT 0.512 19.452 0.544 21.96 ;
  LAYER M3 ;
        RECT 0.512 19.472 0.544 19.504 ;
  LAYER M1 ;
        RECT 0.576 19.452 0.608 21.96 ;
  LAYER M3 ;
        RECT 0.576 21.908 0.608 21.94 ;
  LAYER M1 ;
        RECT 0.64 19.452 0.672 21.96 ;
  LAYER M3 ;
        RECT 0.64 19.472 0.672 19.504 ;
  LAYER M1 ;
        RECT 0.704 19.452 0.736 21.96 ;
  LAYER M3 ;
        RECT 0.704 21.908 0.736 21.94 ;
  LAYER M1 ;
        RECT 0.768 19.452 0.8 21.96 ;
  LAYER M3 ;
        RECT 0.768 19.472 0.8 19.504 ;
  LAYER M1 ;
        RECT 0.832 19.452 0.864 21.96 ;
  LAYER M3 ;
        RECT 0.832 21.908 0.864 21.94 ;
  LAYER M1 ;
        RECT 0.896 19.452 0.928 21.96 ;
  LAYER M3 ;
        RECT 0.896 19.472 0.928 19.504 ;
  LAYER M1 ;
        RECT 0.96 19.452 0.992 21.96 ;
  LAYER M3 ;
        RECT 0.96 21.908 0.992 21.94 ;
  LAYER M1 ;
        RECT 1.024 19.452 1.056 21.96 ;
  LAYER M3 ;
        RECT 1.024 19.472 1.056 19.504 ;
  LAYER M1 ;
        RECT 1.088 19.452 1.12 21.96 ;
  LAYER M3 ;
        RECT 1.088 21.908 1.12 21.94 ;
  LAYER M1 ;
        RECT 1.152 19.452 1.184 21.96 ;
  LAYER M3 ;
        RECT 1.152 19.472 1.184 19.504 ;
  LAYER M1 ;
        RECT 1.216 19.452 1.248 21.96 ;
  LAYER M3 ;
        RECT 1.216 21.908 1.248 21.94 ;
  LAYER M1 ;
        RECT 1.28 19.452 1.312 21.96 ;
  LAYER M3 ;
        RECT 1.28 19.472 1.312 19.504 ;
  LAYER M1 ;
        RECT 1.344 19.452 1.376 21.96 ;
  LAYER M3 ;
        RECT 1.344 21.908 1.376 21.94 ;
  LAYER M1 ;
        RECT 1.408 19.452 1.44 21.96 ;
  LAYER M3 ;
        RECT 1.408 19.472 1.44 19.504 ;
  LAYER M1 ;
        RECT 1.472 19.452 1.504 21.96 ;
  LAYER M3 ;
        RECT 1.472 21.908 1.504 21.94 ;
  LAYER M1 ;
        RECT 1.536 19.452 1.568 21.96 ;
  LAYER M3 ;
        RECT 1.536 19.472 1.568 19.504 ;
  LAYER M1 ;
        RECT 1.6 19.452 1.632 21.96 ;
  LAYER M3 ;
        RECT 1.6 21.908 1.632 21.94 ;
  LAYER M1 ;
        RECT 1.664 19.452 1.696 21.96 ;
  LAYER M3 ;
        RECT 1.664 19.472 1.696 19.504 ;
  LAYER M1 ;
        RECT 1.728 19.452 1.76 21.96 ;
  LAYER M3 ;
        RECT 1.728 21.908 1.76 21.94 ;
  LAYER M1 ;
        RECT 1.792 19.452 1.824 21.96 ;
  LAYER M3 ;
        RECT 1.792 19.472 1.824 19.504 ;
  LAYER M1 ;
        RECT 1.856 19.452 1.888 21.96 ;
  LAYER M3 ;
        RECT 1.856 21.908 1.888 21.94 ;
  LAYER M1 ;
        RECT 1.92 19.452 1.952 21.96 ;
  LAYER M3 ;
        RECT 1.92 19.472 1.952 19.504 ;
  LAYER M1 ;
        RECT 1.984 19.452 2.016 21.96 ;
  LAYER M3 ;
        RECT 1.984 21.908 2.016 21.94 ;
  LAYER M1 ;
        RECT 2.048 19.452 2.08 21.96 ;
  LAYER M3 ;
        RECT 2.048 19.472 2.08 19.504 ;
  LAYER M1 ;
        RECT 2.112 19.452 2.144 21.96 ;
  LAYER M3 ;
        RECT 2.112 21.908 2.144 21.94 ;
  LAYER M1 ;
        RECT 2.176 19.452 2.208 21.96 ;
  LAYER M3 ;
        RECT 2.176 19.472 2.208 19.504 ;
  LAYER M1 ;
        RECT 2.24 19.452 2.272 21.96 ;
  LAYER M3 ;
        RECT 2.24 21.908 2.272 21.94 ;
  LAYER M1 ;
        RECT 2.304 19.452 2.336 21.96 ;
  LAYER M3 ;
        RECT 2.304 19.472 2.336 19.504 ;
  LAYER M1 ;
        RECT 2.368 19.452 2.4 21.96 ;
  LAYER M3 ;
        RECT 2.368 21.908 2.4 21.94 ;
  LAYER M1 ;
        RECT 2.432 19.452 2.464 21.96 ;
  LAYER M3 ;
        RECT 2.432 19.472 2.464 19.504 ;
  LAYER M1 ;
        RECT 2.496 19.452 2.528 21.96 ;
  LAYER M3 ;
        RECT 2.496 21.908 2.528 21.94 ;
  LAYER M1 ;
        RECT 2.56 19.452 2.592 21.96 ;
  LAYER M3 ;
        RECT 2.56 19.472 2.592 19.504 ;
  LAYER M1 ;
        RECT 2.624 19.452 2.656 21.96 ;
  LAYER M3 ;
        RECT 2.624 21.908 2.656 21.94 ;
  LAYER M1 ;
        RECT 2.688 19.452 2.72 21.96 ;
  LAYER M3 ;
        RECT 2.688 19.472 2.72 19.504 ;
  LAYER M1 ;
        RECT 2.752 19.452 2.784 21.96 ;
  LAYER M3 ;
        RECT 2.752 21.908 2.784 21.94 ;
  LAYER M1 ;
        RECT 2.816 19.452 2.848 21.96 ;
  LAYER M3 ;
        RECT 0.448 19.536 0.48 19.568 ;
  LAYER M2 ;
        RECT 2.816 19.6 2.848 19.632 ;
  LAYER M2 ;
        RECT 0.448 19.664 0.48 19.696 ;
  LAYER M2 ;
        RECT 2.816 19.728 2.848 19.76 ;
  LAYER M2 ;
        RECT 0.448 19.792 0.48 19.824 ;
  LAYER M2 ;
        RECT 2.816 19.856 2.848 19.888 ;
  LAYER M2 ;
        RECT 0.448 19.92 0.48 19.952 ;
  LAYER M2 ;
        RECT 2.816 19.984 2.848 20.016 ;
  LAYER M2 ;
        RECT 0.448 20.048 0.48 20.08 ;
  LAYER M2 ;
        RECT 2.816 20.112 2.848 20.144 ;
  LAYER M2 ;
        RECT 0.448 20.176 0.48 20.208 ;
  LAYER M2 ;
        RECT 2.816 20.24 2.848 20.272 ;
  LAYER M2 ;
        RECT 0.448 20.304 0.48 20.336 ;
  LAYER M2 ;
        RECT 2.816 20.368 2.848 20.4 ;
  LAYER M2 ;
        RECT 0.448 20.432 0.48 20.464 ;
  LAYER M2 ;
        RECT 2.816 20.496 2.848 20.528 ;
  LAYER M2 ;
        RECT 0.448 20.56 0.48 20.592 ;
  LAYER M2 ;
        RECT 2.816 20.624 2.848 20.656 ;
  LAYER M2 ;
        RECT 0.448 20.688 0.48 20.72 ;
  LAYER M2 ;
        RECT 2.816 20.752 2.848 20.784 ;
  LAYER M2 ;
        RECT 0.448 20.816 0.48 20.848 ;
  LAYER M2 ;
        RECT 2.816 20.88 2.848 20.912 ;
  LAYER M2 ;
        RECT 0.448 20.944 0.48 20.976 ;
  LAYER M2 ;
        RECT 2.816 21.008 2.848 21.04 ;
  LAYER M2 ;
        RECT 0.448 21.072 0.48 21.104 ;
  LAYER M2 ;
        RECT 2.816 21.136 2.848 21.168 ;
  LAYER M2 ;
        RECT 0.448 21.2 0.48 21.232 ;
  LAYER M2 ;
        RECT 2.816 21.264 2.848 21.296 ;
  LAYER M2 ;
        RECT 0.448 21.328 0.48 21.36 ;
  LAYER M2 ;
        RECT 2.816 21.392 2.848 21.424 ;
  LAYER M2 ;
        RECT 0.448 21.456 0.48 21.488 ;
  LAYER M2 ;
        RECT 2.816 21.52 2.848 21.552 ;
  LAYER M2 ;
        RECT 0.448 21.584 0.48 21.616 ;
  LAYER M2 ;
        RECT 2.816 21.648 2.848 21.68 ;
  LAYER M2 ;
        RECT 0.448 21.712 0.48 21.744 ;
  LAYER M2 ;
        RECT 2.816 21.776 2.848 21.808 ;
  LAYER M2 ;
        RECT 0.4 19.404 2.896 22.008 ;
  LAYER M1 ;
        RECT 0.448 22.56 0.48 25.068 ;
  LAYER M3 ;
        RECT 0.448 25.016 0.48 25.048 ;
  LAYER M1 ;
        RECT 0.512 22.56 0.544 25.068 ;
  LAYER M3 ;
        RECT 0.512 22.58 0.544 22.612 ;
  LAYER M1 ;
        RECT 0.576 22.56 0.608 25.068 ;
  LAYER M3 ;
        RECT 0.576 25.016 0.608 25.048 ;
  LAYER M1 ;
        RECT 0.64 22.56 0.672 25.068 ;
  LAYER M3 ;
        RECT 0.64 22.58 0.672 22.612 ;
  LAYER M1 ;
        RECT 0.704 22.56 0.736 25.068 ;
  LAYER M3 ;
        RECT 0.704 25.016 0.736 25.048 ;
  LAYER M1 ;
        RECT 0.768 22.56 0.8 25.068 ;
  LAYER M3 ;
        RECT 0.768 22.58 0.8 22.612 ;
  LAYER M1 ;
        RECT 0.832 22.56 0.864 25.068 ;
  LAYER M3 ;
        RECT 0.832 25.016 0.864 25.048 ;
  LAYER M1 ;
        RECT 0.896 22.56 0.928 25.068 ;
  LAYER M3 ;
        RECT 0.896 22.58 0.928 22.612 ;
  LAYER M1 ;
        RECT 0.96 22.56 0.992 25.068 ;
  LAYER M3 ;
        RECT 0.96 25.016 0.992 25.048 ;
  LAYER M1 ;
        RECT 1.024 22.56 1.056 25.068 ;
  LAYER M3 ;
        RECT 1.024 22.58 1.056 22.612 ;
  LAYER M1 ;
        RECT 1.088 22.56 1.12 25.068 ;
  LAYER M3 ;
        RECT 1.088 25.016 1.12 25.048 ;
  LAYER M1 ;
        RECT 1.152 22.56 1.184 25.068 ;
  LAYER M3 ;
        RECT 1.152 22.58 1.184 22.612 ;
  LAYER M1 ;
        RECT 1.216 22.56 1.248 25.068 ;
  LAYER M3 ;
        RECT 1.216 25.016 1.248 25.048 ;
  LAYER M1 ;
        RECT 1.28 22.56 1.312 25.068 ;
  LAYER M3 ;
        RECT 1.28 22.58 1.312 22.612 ;
  LAYER M1 ;
        RECT 1.344 22.56 1.376 25.068 ;
  LAYER M3 ;
        RECT 1.344 25.016 1.376 25.048 ;
  LAYER M1 ;
        RECT 1.408 22.56 1.44 25.068 ;
  LAYER M3 ;
        RECT 1.408 22.58 1.44 22.612 ;
  LAYER M1 ;
        RECT 1.472 22.56 1.504 25.068 ;
  LAYER M3 ;
        RECT 1.472 25.016 1.504 25.048 ;
  LAYER M1 ;
        RECT 1.536 22.56 1.568 25.068 ;
  LAYER M3 ;
        RECT 1.536 22.58 1.568 22.612 ;
  LAYER M1 ;
        RECT 1.6 22.56 1.632 25.068 ;
  LAYER M3 ;
        RECT 1.6 25.016 1.632 25.048 ;
  LAYER M1 ;
        RECT 1.664 22.56 1.696 25.068 ;
  LAYER M3 ;
        RECT 1.664 22.58 1.696 22.612 ;
  LAYER M1 ;
        RECT 1.728 22.56 1.76 25.068 ;
  LAYER M3 ;
        RECT 1.728 25.016 1.76 25.048 ;
  LAYER M1 ;
        RECT 1.792 22.56 1.824 25.068 ;
  LAYER M3 ;
        RECT 1.792 22.58 1.824 22.612 ;
  LAYER M1 ;
        RECT 1.856 22.56 1.888 25.068 ;
  LAYER M3 ;
        RECT 1.856 25.016 1.888 25.048 ;
  LAYER M1 ;
        RECT 1.92 22.56 1.952 25.068 ;
  LAYER M3 ;
        RECT 1.92 22.58 1.952 22.612 ;
  LAYER M1 ;
        RECT 1.984 22.56 2.016 25.068 ;
  LAYER M3 ;
        RECT 1.984 25.016 2.016 25.048 ;
  LAYER M1 ;
        RECT 2.048 22.56 2.08 25.068 ;
  LAYER M3 ;
        RECT 2.048 22.58 2.08 22.612 ;
  LAYER M1 ;
        RECT 2.112 22.56 2.144 25.068 ;
  LAYER M3 ;
        RECT 2.112 25.016 2.144 25.048 ;
  LAYER M1 ;
        RECT 2.176 22.56 2.208 25.068 ;
  LAYER M3 ;
        RECT 2.176 22.58 2.208 22.612 ;
  LAYER M1 ;
        RECT 2.24 22.56 2.272 25.068 ;
  LAYER M3 ;
        RECT 2.24 25.016 2.272 25.048 ;
  LAYER M1 ;
        RECT 2.304 22.56 2.336 25.068 ;
  LAYER M3 ;
        RECT 2.304 22.58 2.336 22.612 ;
  LAYER M1 ;
        RECT 2.368 22.56 2.4 25.068 ;
  LAYER M3 ;
        RECT 2.368 25.016 2.4 25.048 ;
  LAYER M1 ;
        RECT 2.432 22.56 2.464 25.068 ;
  LAYER M3 ;
        RECT 2.432 22.58 2.464 22.612 ;
  LAYER M1 ;
        RECT 2.496 22.56 2.528 25.068 ;
  LAYER M3 ;
        RECT 2.496 25.016 2.528 25.048 ;
  LAYER M1 ;
        RECT 2.56 22.56 2.592 25.068 ;
  LAYER M3 ;
        RECT 2.56 22.58 2.592 22.612 ;
  LAYER M1 ;
        RECT 2.624 22.56 2.656 25.068 ;
  LAYER M3 ;
        RECT 2.624 25.016 2.656 25.048 ;
  LAYER M1 ;
        RECT 2.688 22.56 2.72 25.068 ;
  LAYER M3 ;
        RECT 2.688 22.58 2.72 22.612 ;
  LAYER M1 ;
        RECT 2.752 22.56 2.784 25.068 ;
  LAYER M3 ;
        RECT 2.752 25.016 2.784 25.048 ;
  LAYER M1 ;
        RECT 2.816 22.56 2.848 25.068 ;
  LAYER M3 ;
        RECT 0.448 22.644 0.48 22.676 ;
  LAYER M2 ;
        RECT 2.816 22.708 2.848 22.74 ;
  LAYER M2 ;
        RECT 0.448 22.772 0.48 22.804 ;
  LAYER M2 ;
        RECT 2.816 22.836 2.848 22.868 ;
  LAYER M2 ;
        RECT 0.448 22.9 0.48 22.932 ;
  LAYER M2 ;
        RECT 2.816 22.964 2.848 22.996 ;
  LAYER M2 ;
        RECT 0.448 23.028 0.48 23.06 ;
  LAYER M2 ;
        RECT 2.816 23.092 2.848 23.124 ;
  LAYER M2 ;
        RECT 0.448 23.156 0.48 23.188 ;
  LAYER M2 ;
        RECT 2.816 23.22 2.848 23.252 ;
  LAYER M2 ;
        RECT 0.448 23.284 0.48 23.316 ;
  LAYER M2 ;
        RECT 2.816 23.348 2.848 23.38 ;
  LAYER M2 ;
        RECT 0.448 23.412 0.48 23.444 ;
  LAYER M2 ;
        RECT 2.816 23.476 2.848 23.508 ;
  LAYER M2 ;
        RECT 0.448 23.54 0.48 23.572 ;
  LAYER M2 ;
        RECT 2.816 23.604 2.848 23.636 ;
  LAYER M2 ;
        RECT 0.448 23.668 0.48 23.7 ;
  LAYER M2 ;
        RECT 2.816 23.732 2.848 23.764 ;
  LAYER M2 ;
        RECT 0.448 23.796 0.48 23.828 ;
  LAYER M2 ;
        RECT 2.816 23.86 2.848 23.892 ;
  LAYER M2 ;
        RECT 0.448 23.924 0.48 23.956 ;
  LAYER M2 ;
        RECT 2.816 23.988 2.848 24.02 ;
  LAYER M2 ;
        RECT 0.448 24.052 0.48 24.084 ;
  LAYER M2 ;
        RECT 2.816 24.116 2.848 24.148 ;
  LAYER M2 ;
        RECT 0.448 24.18 0.48 24.212 ;
  LAYER M2 ;
        RECT 2.816 24.244 2.848 24.276 ;
  LAYER M2 ;
        RECT 0.448 24.308 0.48 24.34 ;
  LAYER M2 ;
        RECT 2.816 24.372 2.848 24.404 ;
  LAYER M2 ;
        RECT 0.448 24.436 0.48 24.468 ;
  LAYER M2 ;
        RECT 2.816 24.5 2.848 24.532 ;
  LAYER M2 ;
        RECT 0.448 24.564 0.48 24.596 ;
  LAYER M2 ;
        RECT 2.816 24.628 2.848 24.66 ;
  LAYER M2 ;
        RECT 0.448 24.692 0.48 24.724 ;
  LAYER M2 ;
        RECT 2.816 24.756 2.848 24.788 ;
  LAYER M2 ;
        RECT 0.448 24.82 0.48 24.852 ;
  LAYER M2 ;
        RECT 2.816 24.884 2.848 24.916 ;
  LAYER M2 ;
        RECT 0.4 22.512 2.896 25.116 ;
  LAYER M1 ;
        RECT 3.424 0.804 3.456 3.312 ;
  LAYER M3 ;
        RECT 3.424 3.26 3.456 3.292 ;
  LAYER M1 ;
        RECT 3.488 0.804 3.52 3.312 ;
  LAYER M3 ;
        RECT 3.488 0.824 3.52 0.856 ;
  LAYER M1 ;
        RECT 3.552 0.804 3.584 3.312 ;
  LAYER M3 ;
        RECT 3.552 3.26 3.584 3.292 ;
  LAYER M1 ;
        RECT 3.616 0.804 3.648 3.312 ;
  LAYER M3 ;
        RECT 3.616 0.824 3.648 0.856 ;
  LAYER M1 ;
        RECT 3.68 0.804 3.712 3.312 ;
  LAYER M3 ;
        RECT 3.68 3.26 3.712 3.292 ;
  LAYER M1 ;
        RECT 3.744 0.804 3.776 3.312 ;
  LAYER M3 ;
        RECT 3.744 0.824 3.776 0.856 ;
  LAYER M1 ;
        RECT 3.808 0.804 3.84 3.312 ;
  LAYER M3 ;
        RECT 3.808 3.26 3.84 3.292 ;
  LAYER M1 ;
        RECT 3.872 0.804 3.904 3.312 ;
  LAYER M3 ;
        RECT 3.872 0.824 3.904 0.856 ;
  LAYER M1 ;
        RECT 3.936 0.804 3.968 3.312 ;
  LAYER M3 ;
        RECT 3.936 3.26 3.968 3.292 ;
  LAYER M1 ;
        RECT 4 0.804 4.032 3.312 ;
  LAYER M3 ;
        RECT 4 0.824 4.032 0.856 ;
  LAYER M1 ;
        RECT 4.064 0.804 4.096 3.312 ;
  LAYER M3 ;
        RECT 4.064 3.26 4.096 3.292 ;
  LAYER M1 ;
        RECT 4.128 0.804 4.16 3.312 ;
  LAYER M3 ;
        RECT 4.128 0.824 4.16 0.856 ;
  LAYER M1 ;
        RECT 4.192 0.804 4.224 3.312 ;
  LAYER M3 ;
        RECT 4.192 3.26 4.224 3.292 ;
  LAYER M1 ;
        RECT 4.256 0.804 4.288 3.312 ;
  LAYER M3 ;
        RECT 4.256 0.824 4.288 0.856 ;
  LAYER M1 ;
        RECT 4.32 0.804 4.352 3.312 ;
  LAYER M3 ;
        RECT 4.32 3.26 4.352 3.292 ;
  LAYER M1 ;
        RECT 4.384 0.804 4.416 3.312 ;
  LAYER M3 ;
        RECT 4.384 0.824 4.416 0.856 ;
  LAYER M1 ;
        RECT 4.448 0.804 4.48 3.312 ;
  LAYER M3 ;
        RECT 4.448 3.26 4.48 3.292 ;
  LAYER M1 ;
        RECT 4.512 0.804 4.544 3.312 ;
  LAYER M3 ;
        RECT 4.512 0.824 4.544 0.856 ;
  LAYER M1 ;
        RECT 4.576 0.804 4.608 3.312 ;
  LAYER M3 ;
        RECT 4.576 3.26 4.608 3.292 ;
  LAYER M1 ;
        RECT 4.64 0.804 4.672 3.312 ;
  LAYER M3 ;
        RECT 4.64 0.824 4.672 0.856 ;
  LAYER M1 ;
        RECT 4.704 0.804 4.736 3.312 ;
  LAYER M3 ;
        RECT 4.704 3.26 4.736 3.292 ;
  LAYER M1 ;
        RECT 4.768 0.804 4.8 3.312 ;
  LAYER M3 ;
        RECT 4.768 0.824 4.8 0.856 ;
  LAYER M1 ;
        RECT 4.832 0.804 4.864 3.312 ;
  LAYER M3 ;
        RECT 4.832 3.26 4.864 3.292 ;
  LAYER M1 ;
        RECT 4.896 0.804 4.928 3.312 ;
  LAYER M3 ;
        RECT 4.896 0.824 4.928 0.856 ;
  LAYER M1 ;
        RECT 4.96 0.804 4.992 3.312 ;
  LAYER M3 ;
        RECT 4.96 3.26 4.992 3.292 ;
  LAYER M1 ;
        RECT 5.024 0.804 5.056 3.312 ;
  LAYER M3 ;
        RECT 5.024 0.824 5.056 0.856 ;
  LAYER M1 ;
        RECT 5.088 0.804 5.12 3.312 ;
  LAYER M3 ;
        RECT 5.088 3.26 5.12 3.292 ;
  LAYER M1 ;
        RECT 5.152 0.804 5.184 3.312 ;
  LAYER M3 ;
        RECT 5.152 0.824 5.184 0.856 ;
  LAYER M1 ;
        RECT 5.216 0.804 5.248 3.312 ;
  LAYER M3 ;
        RECT 5.216 3.26 5.248 3.292 ;
  LAYER M1 ;
        RECT 5.28 0.804 5.312 3.312 ;
  LAYER M3 ;
        RECT 5.28 0.824 5.312 0.856 ;
  LAYER M1 ;
        RECT 5.344 0.804 5.376 3.312 ;
  LAYER M3 ;
        RECT 5.344 3.26 5.376 3.292 ;
  LAYER M1 ;
        RECT 5.408 0.804 5.44 3.312 ;
  LAYER M3 ;
        RECT 5.408 0.824 5.44 0.856 ;
  LAYER M1 ;
        RECT 5.472 0.804 5.504 3.312 ;
  LAYER M3 ;
        RECT 5.472 3.26 5.504 3.292 ;
  LAYER M1 ;
        RECT 5.536 0.804 5.568 3.312 ;
  LAYER M3 ;
        RECT 5.536 0.824 5.568 0.856 ;
  LAYER M1 ;
        RECT 5.6 0.804 5.632 3.312 ;
  LAYER M3 ;
        RECT 5.6 3.26 5.632 3.292 ;
  LAYER M1 ;
        RECT 5.664 0.804 5.696 3.312 ;
  LAYER M3 ;
        RECT 5.664 0.824 5.696 0.856 ;
  LAYER M1 ;
        RECT 5.728 0.804 5.76 3.312 ;
  LAYER M3 ;
        RECT 5.728 3.26 5.76 3.292 ;
  LAYER M1 ;
        RECT 5.792 0.804 5.824 3.312 ;
  LAYER M3 ;
        RECT 3.424 0.888 3.456 0.92 ;
  LAYER M2 ;
        RECT 5.792 0.952 5.824 0.984 ;
  LAYER M2 ;
        RECT 3.424 1.016 3.456 1.048 ;
  LAYER M2 ;
        RECT 5.792 1.08 5.824 1.112 ;
  LAYER M2 ;
        RECT 3.424 1.144 3.456 1.176 ;
  LAYER M2 ;
        RECT 5.792 1.208 5.824 1.24 ;
  LAYER M2 ;
        RECT 3.424 1.272 3.456 1.304 ;
  LAYER M2 ;
        RECT 5.792 1.336 5.824 1.368 ;
  LAYER M2 ;
        RECT 3.424 1.4 3.456 1.432 ;
  LAYER M2 ;
        RECT 5.792 1.464 5.824 1.496 ;
  LAYER M2 ;
        RECT 3.424 1.528 3.456 1.56 ;
  LAYER M2 ;
        RECT 5.792 1.592 5.824 1.624 ;
  LAYER M2 ;
        RECT 3.424 1.656 3.456 1.688 ;
  LAYER M2 ;
        RECT 5.792 1.72 5.824 1.752 ;
  LAYER M2 ;
        RECT 3.424 1.784 3.456 1.816 ;
  LAYER M2 ;
        RECT 5.792 1.848 5.824 1.88 ;
  LAYER M2 ;
        RECT 3.424 1.912 3.456 1.944 ;
  LAYER M2 ;
        RECT 5.792 1.976 5.824 2.008 ;
  LAYER M2 ;
        RECT 3.424 2.04 3.456 2.072 ;
  LAYER M2 ;
        RECT 5.792 2.104 5.824 2.136 ;
  LAYER M2 ;
        RECT 3.424 2.168 3.456 2.2 ;
  LAYER M2 ;
        RECT 5.792 2.232 5.824 2.264 ;
  LAYER M2 ;
        RECT 3.424 2.296 3.456 2.328 ;
  LAYER M2 ;
        RECT 5.792 2.36 5.824 2.392 ;
  LAYER M2 ;
        RECT 3.424 2.424 3.456 2.456 ;
  LAYER M2 ;
        RECT 5.792 2.488 5.824 2.52 ;
  LAYER M2 ;
        RECT 3.424 2.552 3.456 2.584 ;
  LAYER M2 ;
        RECT 5.792 2.616 5.824 2.648 ;
  LAYER M2 ;
        RECT 3.424 2.68 3.456 2.712 ;
  LAYER M2 ;
        RECT 5.792 2.744 5.824 2.776 ;
  LAYER M2 ;
        RECT 3.424 2.808 3.456 2.84 ;
  LAYER M2 ;
        RECT 5.792 2.872 5.824 2.904 ;
  LAYER M2 ;
        RECT 3.424 2.936 3.456 2.968 ;
  LAYER M2 ;
        RECT 5.792 3 5.824 3.032 ;
  LAYER M2 ;
        RECT 3.424 3.064 3.456 3.096 ;
  LAYER M2 ;
        RECT 5.792 3.128 5.824 3.16 ;
  LAYER M2 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M1 ;
        RECT 3.424 3.912 3.456 6.42 ;
  LAYER M3 ;
        RECT 3.424 6.368 3.456 6.4 ;
  LAYER M1 ;
        RECT 3.488 3.912 3.52 6.42 ;
  LAYER M3 ;
        RECT 3.488 3.932 3.52 3.964 ;
  LAYER M1 ;
        RECT 3.552 3.912 3.584 6.42 ;
  LAYER M3 ;
        RECT 3.552 6.368 3.584 6.4 ;
  LAYER M1 ;
        RECT 3.616 3.912 3.648 6.42 ;
  LAYER M3 ;
        RECT 3.616 3.932 3.648 3.964 ;
  LAYER M1 ;
        RECT 3.68 3.912 3.712 6.42 ;
  LAYER M3 ;
        RECT 3.68 6.368 3.712 6.4 ;
  LAYER M1 ;
        RECT 3.744 3.912 3.776 6.42 ;
  LAYER M3 ;
        RECT 3.744 3.932 3.776 3.964 ;
  LAYER M1 ;
        RECT 3.808 3.912 3.84 6.42 ;
  LAYER M3 ;
        RECT 3.808 6.368 3.84 6.4 ;
  LAYER M1 ;
        RECT 3.872 3.912 3.904 6.42 ;
  LAYER M3 ;
        RECT 3.872 3.932 3.904 3.964 ;
  LAYER M1 ;
        RECT 3.936 3.912 3.968 6.42 ;
  LAYER M3 ;
        RECT 3.936 6.368 3.968 6.4 ;
  LAYER M1 ;
        RECT 4 3.912 4.032 6.42 ;
  LAYER M3 ;
        RECT 4 3.932 4.032 3.964 ;
  LAYER M1 ;
        RECT 4.064 3.912 4.096 6.42 ;
  LAYER M3 ;
        RECT 4.064 6.368 4.096 6.4 ;
  LAYER M1 ;
        RECT 4.128 3.912 4.16 6.42 ;
  LAYER M3 ;
        RECT 4.128 3.932 4.16 3.964 ;
  LAYER M1 ;
        RECT 4.192 3.912 4.224 6.42 ;
  LAYER M3 ;
        RECT 4.192 6.368 4.224 6.4 ;
  LAYER M1 ;
        RECT 4.256 3.912 4.288 6.42 ;
  LAYER M3 ;
        RECT 4.256 3.932 4.288 3.964 ;
  LAYER M1 ;
        RECT 4.32 3.912 4.352 6.42 ;
  LAYER M3 ;
        RECT 4.32 6.368 4.352 6.4 ;
  LAYER M1 ;
        RECT 4.384 3.912 4.416 6.42 ;
  LAYER M3 ;
        RECT 4.384 3.932 4.416 3.964 ;
  LAYER M1 ;
        RECT 4.448 3.912 4.48 6.42 ;
  LAYER M3 ;
        RECT 4.448 6.368 4.48 6.4 ;
  LAYER M1 ;
        RECT 4.512 3.912 4.544 6.42 ;
  LAYER M3 ;
        RECT 4.512 3.932 4.544 3.964 ;
  LAYER M1 ;
        RECT 4.576 3.912 4.608 6.42 ;
  LAYER M3 ;
        RECT 4.576 6.368 4.608 6.4 ;
  LAYER M1 ;
        RECT 4.64 3.912 4.672 6.42 ;
  LAYER M3 ;
        RECT 4.64 3.932 4.672 3.964 ;
  LAYER M1 ;
        RECT 4.704 3.912 4.736 6.42 ;
  LAYER M3 ;
        RECT 4.704 6.368 4.736 6.4 ;
  LAYER M1 ;
        RECT 4.768 3.912 4.8 6.42 ;
  LAYER M3 ;
        RECT 4.768 3.932 4.8 3.964 ;
  LAYER M1 ;
        RECT 4.832 3.912 4.864 6.42 ;
  LAYER M3 ;
        RECT 4.832 6.368 4.864 6.4 ;
  LAYER M1 ;
        RECT 4.896 3.912 4.928 6.42 ;
  LAYER M3 ;
        RECT 4.896 3.932 4.928 3.964 ;
  LAYER M1 ;
        RECT 4.96 3.912 4.992 6.42 ;
  LAYER M3 ;
        RECT 4.96 6.368 4.992 6.4 ;
  LAYER M1 ;
        RECT 5.024 3.912 5.056 6.42 ;
  LAYER M3 ;
        RECT 5.024 3.932 5.056 3.964 ;
  LAYER M1 ;
        RECT 5.088 3.912 5.12 6.42 ;
  LAYER M3 ;
        RECT 5.088 6.368 5.12 6.4 ;
  LAYER M1 ;
        RECT 5.152 3.912 5.184 6.42 ;
  LAYER M3 ;
        RECT 5.152 3.932 5.184 3.964 ;
  LAYER M1 ;
        RECT 5.216 3.912 5.248 6.42 ;
  LAYER M3 ;
        RECT 5.216 6.368 5.248 6.4 ;
  LAYER M1 ;
        RECT 5.28 3.912 5.312 6.42 ;
  LAYER M3 ;
        RECT 5.28 3.932 5.312 3.964 ;
  LAYER M1 ;
        RECT 5.344 3.912 5.376 6.42 ;
  LAYER M3 ;
        RECT 5.344 6.368 5.376 6.4 ;
  LAYER M1 ;
        RECT 5.408 3.912 5.44 6.42 ;
  LAYER M3 ;
        RECT 5.408 3.932 5.44 3.964 ;
  LAYER M1 ;
        RECT 5.472 3.912 5.504 6.42 ;
  LAYER M3 ;
        RECT 5.472 6.368 5.504 6.4 ;
  LAYER M1 ;
        RECT 5.536 3.912 5.568 6.42 ;
  LAYER M3 ;
        RECT 5.536 3.932 5.568 3.964 ;
  LAYER M1 ;
        RECT 5.6 3.912 5.632 6.42 ;
  LAYER M3 ;
        RECT 5.6 6.368 5.632 6.4 ;
  LAYER M1 ;
        RECT 5.664 3.912 5.696 6.42 ;
  LAYER M3 ;
        RECT 5.664 3.932 5.696 3.964 ;
  LAYER M1 ;
        RECT 5.728 3.912 5.76 6.42 ;
  LAYER M3 ;
        RECT 5.728 6.368 5.76 6.4 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 6.42 ;
  LAYER M3 ;
        RECT 3.424 3.996 3.456 4.028 ;
  LAYER M2 ;
        RECT 5.792 4.06 5.824 4.092 ;
  LAYER M2 ;
        RECT 3.424 4.124 3.456 4.156 ;
  LAYER M2 ;
        RECT 5.792 4.188 5.824 4.22 ;
  LAYER M2 ;
        RECT 3.424 4.252 3.456 4.284 ;
  LAYER M2 ;
        RECT 5.792 4.316 5.824 4.348 ;
  LAYER M2 ;
        RECT 3.424 4.38 3.456 4.412 ;
  LAYER M2 ;
        RECT 5.792 4.444 5.824 4.476 ;
  LAYER M2 ;
        RECT 3.424 4.508 3.456 4.54 ;
  LAYER M2 ;
        RECT 5.792 4.572 5.824 4.604 ;
  LAYER M2 ;
        RECT 3.424 4.636 3.456 4.668 ;
  LAYER M2 ;
        RECT 5.792 4.7 5.824 4.732 ;
  LAYER M2 ;
        RECT 3.424 4.764 3.456 4.796 ;
  LAYER M2 ;
        RECT 5.792 4.828 5.824 4.86 ;
  LAYER M2 ;
        RECT 3.424 4.892 3.456 4.924 ;
  LAYER M2 ;
        RECT 5.792 4.956 5.824 4.988 ;
  LAYER M2 ;
        RECT 3.424 5.02 3.456 5.052 ;
  LAYER M2 ;
        RECT 5.792 5.084 5.824 5.116 ;
  LAYER M2 ;
        RECT 3.424 5.148 3.456 5.18 ;
  LAYER M2 ;
        RECT 5.792 5.212 5.824 5.244 ;
  LAYER M2 ;
        RECT 3.424 5.276 3.456 5.308 ;
  LAYER M2 ;
        RECT 5.792 5.34 5.824 5.372 ;
  LAYER M2 ;
        RECT 3.424 5.404 3.456 5.436 ;
  LAYER M2 ;
        RECT 5.792 5.468 5.824 5.5 ;
  LAYER M2 ;
        RECT 3.424 5.532 3.456 5.564 ;
  LAYER M2 ;
        RECT 5.792 5.596 5.824 5.628 ;
  LAYER M2 ;
        RECT 3.424 5.66 3.456 5.692 ;
  LAYER M2 ;
        RECT 5.792 5.724 5.824 5.756 ;
  LAYER M2 ;
        RECT 3.424 5.788 3.456 5.82 ;
  LAYER M2 ;
        RECT 5.792 5.852 5.824 5.884 ;
  LAYER M2 ;
        RECT 3.424 5.916 3.456 5.948 ;
  LAYER M2 ;
        RECT 5.792 5.98 5.824 6.012 ;
  LAYER M2 ;
        RECT 3.424 6.044 3.456 6.076 ;
  LAYER M2 ;
        RECT 5.792 6.108 5.824 6.14 ;
  LAYER M2 ;
        RECT 3.424 6.172 3.456 6.204 ;
  LAYER M2 ;
        RECT 5.792 6.236 5.824 6.268 ;
  LAYER M2 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M1 ;
        RECT 3.424 7.02 3.456 9.528 ;
  LAYER M3 ;
        RECT 3.424 9.476 3.456 9.508 ;
  LAYER M1 ;
        RECT 3.488 7.02 3.52 9.528 ;
  LAYER M3 ;
        RECT 3.488 7.04 3.52 7.072 ;
  LAYER M1 ;
        RECT 3.552 7.02 3.584 9.528 ;
  LAYER M3 ;
        RECT 3.552 9.476 3.584 9.508 ;
  LAYER M1 ;
        RECT 3.616 7.02 3.648 9.528 ;
  LAYER M3 ;
        RECT 3.616 7.04 3.648 7.072 ;
  LAYER M1 ;
        RECT 3.68 7.02 3.712 9.528 ;
  LAYER M3 ;
        RECT 3.68 9.476 3.712 9.508 ;
  LAYER M1 ;
        RECT 3.744 7.02 3.776 9.528 ;
  LAYER M3 ;
        RECT 3.744 7.04 3.776 7.072 ;
  LAYER M1 ;
        RECT 3.808 7.02 3.84 9.528 ;
  LAYER M3 ;
        RECT 3.808 9.476 3.84 9.508 ;
  LAYER M1 ;
        RECT 3.872 7.02 3.904 9.528 ;
  LAYER M3 ;
        RECT 3.872 7.04 3.904 7.072 ;
  LAYER M1 ;
        RECT 3.936 7.02 3.968 9.528 ;
  LAYER M3 ;
        RECT 3.936 9.476 3.968 9.508 ;
  LAYER M1 ;
        RECT 4 7.02 4.032 9.528 ;
  LAYER M3 ;
        RECT 4 7.04 4.032 7.072 ;
  LAYER M1 ;
        RECT 4.064 7.02 4.096 9.528 ;
  LAYER M3 ;
        RECT 4.064 9.476 4.096 9.508 ;
  LAYER M1 ;
        RECT 4.128 7.02 4.16 9.528 ;
  LAYER M3 ;
        RECT 4.128 7.04 4.16 7.072 ;
  LAYER M1 ;
        RECT 4.192 7.02 4.224 9.528 ;
  LAYER M3 ;
        RECT 4.192 9.476 4.224 9.508 ;
  LAYER M1 ;
        RECT 4.256 7.02 4.288 9.528 ;
  LAYER M3 ;
        RECT 4.256 7.04 4.288 7.072 ;
  LAYER M1 ;
        RECT 4.32 7.02 4.352 9.528 ;
  LAYER M3 ;
        RECT 4.32 9.476 4.352 9.508 ;
  LAYER M1 ;
        RECT 4.384 7.02 4.416 9.528 ;
  LAYER M3 ;
        RECT 4.384 7.04 4.416 7.072 ;
  LAYER M1 ;
        RECT 4.448 7.02 4.48 9.528 ;
  LAYER M3 ;
        RECT 4.448 9.476 4.48 9.508 ;
  LAYER M1 ;
        RECT 4.512 7.02 4.544 9.528 ;
  LAYER M3 ;
        RECT 4.512 7.04 4.544 7.072 ;
  LAYER M1 ;
        RECT 4.576 7.02 4.608 9.528 ;
  LAYER M3 ;
        RECT 4.576 9.476 4.608 9.508 ;
  LAYER M1 ;
        RECT 4.64 7.02 4.672 9.528 ;
  LAYER M3 ;
        RECT 4.64 7.04 4.672 7.072 ;
  LAYER M1 ;
        RECT 4.704 7.02 4.736 9.528 ;
  LAYER M3 ;
        RECT 4.704 9.476 4.736 9.508 ;
  LAYER M1 ;
        RECT 4.768 7.02 4.8 9.528 ;
  LAYER M3 ;
        RECT 4.768 7.04 4.8 7.072 ;
  LAYER M1 ;
        RECT 4.832 7.02 4.864 9.528 ;
  LAYER M3 ;
        RECT 4.832 9.476 4.864 9.508 ;
  LAYER M1 ;
        RECT 4.896 7.02 4.928 9.528 ;
  LAYER M3 ;
        RECT 4.896 7.04 4.928 7.072 ;
  LAYER M1 ;
        RECT 4.96 7.02 4.992 9.528 ;
  LAYER M3 ;
        RECT 4.96 9.476 4.992 9.508 ;
  LAYER M1 ;
        RECT 5.024 7.02 5.056 9.528 ;
  LAYER M3 ;
        RECT 5.024 7.04 5.056 7.072 ;
  LAYER M1 ;
        RECT 5.088 7.02 5.12 9.528 ;
  LAYER M3 ;
        RECT 5.088 9.476 5.12 9.508 ;
  LAYER M1 ;
        RECT 5.152 7.02 5.184 9.528 ;
  LAYER M3 ;
        RECT 5.152 7.04 5.184 7.072 ;
  LAYER M1 ;
        RECT 5.216 7.02 5.248 9.528 ;
  LAYER M3 ;
        RECT 5.216 9.476 5.248 9.508 ;
  LAYER M1 ;
        RECT 5.28 7.02 5.312 9.528 ;
  LAYER M3 ;
        RECT 5.28 7.04 5.312 7.072 ;
  LAYER M1 ;
        RECT 5.344 7.02 5.376 9.528 ;
  LAYER M3 ;
        RECT 5.344 9.476 5.376 9.508 ;
  LAYER M1 ;
        RECT 5.408 7.02 5.44 9.528 ;
  LAYER M3 ;
        RECT 5.408 7.04 5.44 7.072 ;
  LAYER M1 ;
        RECT 5.472 7.02 5.504 9.528 ;
  LAYER M3 ;
        RECT 5.472 9.476 5.504 9.508 ;
  LAYER M1 ;
        RECT 5.536 7.02 5.568 9.528 ;
  LAYER M3 ;
        RECT 5.536 7.04 5.568 7.072 ;
  LAYER M1 ;
        RECT 5.6 7.02 5.632 9.528 ;
  LAYER M3 ;
        RECT 5.6 9.476 5.632 9.508 ;
  LAYER M1 ;
        RECT 5.664 7.02 5.696 9.528 ;
  LAYER M3 ;
        RECT 5.664 7.04 5.696 7.072 ;
  LAYER M1 ;
        RECT 5.728 7.02 5.76 9.528 ;
  LAYER M3 ;
        RECT 5.728 9.476 5.76 9.508 ;
  LAYER M1 ;
        RECT 5.792 7.02 5.824 9.528 ;
  LAYER M3 ;
        RECT 3.424 7.104 3.456 7.136 ;
  LAYER M2 ;
        RECT 5.792 7.168 5.824 7.2 ;
  LAYER M2 ;
        RECT 3.424 7.232 3.456 7.264 ;
  LAYER M2 ;
        RECT 5.792 7.296 5.824 7.328 ;
  LAYER M2 ;
        RECT 3.424 7.36 3.456 7.392 ;
  LAYER M2 ;
        RECT 5.792 7.424 5.824 7.456 ;
  LAYER M2 ;
        RECT 3.424 7.488 3.456 7.52 ;
  LAYER M2 ;
        RECT 5.792 7.552 5.824 7.584 ;
  LAYER M2 ;
        RECT 3.424 7.616 3.456 7.648 ;
  LAYER M2 ;
        RECT 5.792 7.68 5.824 7.712 ;
  LAYER M2 ;
        RECT 3.424 7.744 3.456 7.776 ;
  LAYER M2 ;
        RECT 5.792 7.808 5.824 7.84 ;
  LAYER M2 ;
        RECT 3.424 7.872 3.456 7.904 ;
  LAYER M2 ;
        RECT 5.792 7.936 5.824 7.968 ;
  LAYER M2 ;
        RECT 3.424 8 3.456 8.032 ;
  LAYER M2 ;
        RECT 5.792 8.064 5.824 8.096 ;
  LAYER M2 ;
        RECT 3.424 8.128 3.456 8.16 ;
  LAYER M2 ;
        RECT 5.792 8.192 5.824 8.224 ;
  LAYER M2 ;
        RECT 3.424 8.256 3.456 8.288 ;
  LAYER M2 ;
        RECT 5.792 8.32 5.824 8.352 ;
  LAYER M2 ;
        RECT 3.424 8.384 3.456 8.416 ;
  LAYER M2 ;
        RECT 5.792 8.448 5.824 8.48 ;
  LAYER M2 ;
        RECT 3.424 8.512 3.456 8.544 ;
  LAYER M2 ;
        RECT 5.792 8.576 5.824 8.608 ;
  LAYER M2 ;
        RECT 3.424 8.64 3.456 8.672 ;
  LAYER M2 ;
        RECT 5.792 8.704 5.824 8.736 ;
  LAYER M2 ;
        RECT 3.424 8.768 3.456 8.8 ;
  LAYER M2 ;
        RECT 5.792 8.832 5.824 8.864 ;
  LAYER M2 ;
        RECT 3.424 8.896 3.456 8.928 ;
  LAYER M2 ;
        RECT 5.792 8.96 5.824 8.992 ;
  LAYER M2 ;
        RECT 3.424 9.024 3.456 9.056 ;
  LAYER M2 ;
        RECT 5.792 9.088 5.824 9.12 ;
  LAYER M2 ;
        RECT 3.424 9.152 3.456 9.184 ;
  LAYER M2 ;
        RECT 5.792 9.216 5.824 9.248 ;
  LAYER M2 ;
        RECT 3.424 9.28 3.456 9.312 ;
  LAYER M2 ;
        RECT 5.792 9.344 5.824 9.376 ;
  LAYER M2 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M1 ;
        RECT 3.424 10.128 3.456 12.636 ;
  LAYER M3 ;
        RECT 3.424 12.584 3.456 12.616 ;
  LAYER M1 ;
        RECT 3.488 10.128 3.52 12.636 ;
  LAYER M3 ;
        RECT 3.488 10.148 3.52 10.18 ;
  LAYER M1 ;
        RECT 3.552 10.128 3.584 12.636 ;
  LAYER M3 ;
        RECT 3.552 12.584 3.584 12.616 ;
  LAYER M1 ;
        RECT 3.616 10.128 3.648 12.636 ;
  LAYER M3 ;
        RECT 3.616 10.148 3.648 10.18 ;
  LAYER M1 ;
        RECT 3.68 10.128 3.712 12.636 ;
  LAYER M3 ;
        RECT 3.68 12.584 3.712 12.616 ;
  LAYER M1 ;
        RECT 3.744 10.128 3.776 12.636 ;
  LAYER M3 ;
        RECT 3.744 10.148 3.776 10.18 ;
  LAYER M1 ;
        RECT 3.808 10.128 3.84 12.636 ;
  LAYER M3 ;
        RECT 3.808 12.584 3.84 12.616 ;
  LAYER M1 ;
        RECT 3.872 10.128 3.904 12.636 ;
  LAYER M3 ;
        RECT 3.872 10.148 3.904 10.18 ;
  LAYER M1 ;
        RECT 3.936 10.128 3.968 12.636 ;
  LAYER M3 ;
        RECT 3.936 12.584 3.968 12.616 ;
  LAYER M1 ;
        RECT 4 10.128 4.032 12.636 ;
  LAYER M3 ;
        RECT 4 10.148 4.032 10.18 ;
  LAYER M1 ;
        RECT 4.064 10.128 4.096 12.636 ;
  LAYER M3 ;
        RECT 4.064 12.584 4.096 12.616 ;
  LAYER M1 ;
        RECT 4.128 10.128 4.16 12.636 ;
  LAYER M3 ;
        RECT 4.128 10.148 4.16 10.18 ;
  LAYER M1 ;
        RECT 4.192 10.128 4.224 12.636 ;
  LAYER M3 ;
        RECT 4.192 12.584 4.224 12.616 ;
  LAYER M1 ;
        RECT 4.256 10.128 4.288 12.636 ;
  LAYER M3 ;
        RECT 4.256 10.148 4.288 10.18 ;
  LAYER M1 ;
        RECT 4.32 10.128 4.352 12.636 ;
  LAYER M3 ;
        RECT 4.32 12.584 4.352 12.616 ;
  LAYER M1 ;
        RECT 4.384 10.128 4.416 12.636 ;
  LAYER M3 ;
        RECT 4.384 10.148 4.416 10.18 ;
  LAYER M1 ;
        RECT 4.448 10.128 4.48 12.636 ;
  LAYER M3 ;
        RECT 4.448 12.584 4.48 12.616 ;
  LAYER M1 ;
        RECT 4.512 10.128 4.544 12.636 ;
  LAYER M3 ;
        RECT 4.512 10.148 4.544 10.18 ;
  LAYER M1 ;
        RECT 4.576 10.128 4.608 12.636 ;
  LAYER M3 ;
        RECT 4.576 12.584 4.608 12.616 ;
  LAYER M1 ;
        RECT 4.64 10.128 4.672 12.636 ;
  LAYER M3 ;
        RECT 4.64 10.148 4.672 10.18 ;
  LAYER M1 ;
        RECT 4.704 10.128 4.736 12.636 ;
  LAYER M3 ;
        RECT 4.704 12.584 4.736 12.616 ;
  LAYER M1 ;
        RECT 4.768 10.128 4.8 12.636 ;
  LAYER M3 ;
        RECT 4.768 10.148 4.8 10.18 ;
  LAYER M1 ;
        RECT 4.832 10.128 4.864 12.636 ;
  LAYER M3 ;
        RECT 4.832 12.584 4.864 12.616 ;
  LAYER M1 ;
        RECT 4.896 10.128 4.928 12.636 ;
  LAYER M3 ;
        RECT 4.896 10.148 4.928 10.18 ;
  LAYER M1 ;
        RECT 4.96 10.128 4.992 12.636 ;
  LAYER M3 ;
        RECT 4.96 12.584 4.992 12.616 ;
  LAYER M1 ;
        RECT 5.024 10.128 5.056 12.636 ;
  LAYER M3 ;
        RECT 5.024 10.148 5.056 10.18 ;
  LAYER M1 ;
        RECT 5.088 10.128 5.12 12.636 ;
  LAYER M3 ;
        RECT 5.088 12.584 5.12 12.616 ;
  LAYER M1 ;
        RECT 5.152 10.128 5.184 12.636 ;
  LAYER M3 ;
        RECT 5.152 10.148 5.184 10.18 ;
  LAYER M1 ;
        RECT 5.216 10.128 5.248 12.636 ;
  LAYER M3 ;
        RECT 5.216 12.584 5.248 12.616 ;
  LAYER M1 ;
        RECT 5.28 10.128 5.312 12.636 ;
  LAYER M3 ;
        RECT 5.28 10.148 5.312 10.18 ;
  LAYER M1 ;
        RECT 5.344 10.128 5.376 12.636 ;
  LAYER M3 ;
        RECT 5.344 12.584 5.376 12.616 ;
  LAYER M1 ;
        RECT 5.408 10.128 5.44 12.636 ;
  LAYER M3 ;
        RECT 5.408 10.148 5.44 10.18 ;
  LAYER M1 ;
        RECT 5.472 10.128 5.504 12.636 ;
  LAYER M3 ;
        RECT 5.472 12.584 5.504 12.616 ;
  LAYER M1 ;
        RECT 5.536 10.128 5.568 12.636 ;
  LAYER M3 ;
        RECT 5.536 10.148 5.568 10.18 ;
  LAYER M1 ;
        RECT 5.6 10.128 5.632 12.636 ;
  LAYER M3 ;
        RECT 5.6 12.584 5.632 12.616 ;
  LAYER M1 ;
        RECT 5.664 10.128 5.696 12.636 ;
  LAYER M3 ;
        RECT 5.664 10.148 5.696 10.18 ;
  LAYER M1 ;
        RECT 5.728 10.128 5.76 12.636 ;
  LAYER M3 ;
        RECT 5.728 12.584 5.76 12.616 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 12.636 ;
  LAYER M3 ;
        RECT 3.424 10.212 3.456 10.244 ;
  LAYER M2 ;
        RECT 5.792 10.276 5.824 10.308 ;
  LAYER M2 ;
        RECT 3.424 10.34 3.456 10.372 ;
  LAYER M2 ;
        RECT 5.792 10.404 5.824 10.436 ;
  LAYER M2 ;
        RECT 3.424 10.468 3.456 10.5 ;
  LAYER M2 ;
        RECT 5.792 10.532 5.824 10.564 ;
  LAYER M2 ;
        RECT 3.424 10.596 3.456 10.628 ;
  LAYER M2 ;
        RECT 5.792 10.66 5.824 10.692 ;
  LAYER M2 ;
        RECT 3.424 10.724 3.456 10.756 ;
  LAYER M2 ;
        RECT 5.792 10.788 5.824 10.82 ;
  LAYER M2 ;
        RECT 3.424 10.852 3.456 10.884 ;
  LAYER M2 ;
        RECT 5.792 10.916 5.824 10.948 ;
  LAYER M2 ;
        RECT 3.424 10.98 3.456 11.012 ;
  LAYER M2 ;
        RECT 5.792 11.044 5.824 11.076 ;
  LAYER M2 ;
        RECT 3.424 11.108 3.456 11.14 ;
  LAYER M2 ;
        RECT 5.792 11.172 5.824 11.204 ;
  LAYER M2 ;
        RECT 3.424 11.236 3.456 11.268 ;
  LAYER M2 ;
        RECT 5.792 11.3 5.824 11.332 ;
  LAYER M2 ;
        RECT 3.424 11.364 3.456 11.396 ;
  LAYER M2 ;
        RECT 5.792 11.428 5.824 11.46 ;
  LAYER M2 ;
        RECT 3.424 11.492 3.456 11.524 ;
  LAYER M2 ;
        RECT 5.792 11.556 5.824 11.588 ;
  LAYER M2 ;
        RECT 3.424 11.62 3.456 11.652 ;
  LAYER M2 ;
        RECT 5.792 11.684 5.824 11.716 ;
  LAYER M2 ;
        RECT 3.424 11.748 3.456 11.78 ;
  LAYER M2 ;
        RECT 5.792 11.812 5.824 11.844 ;
  LAYER M2 ;
        RECT 3.424 11.876 3.456 11.908 ;
  LAYER M2 ;
        RECT 5.792 11.94 5.824 11.972 ;
  LAYER M2 ;
        RECT 3.424 12.004 3.456 12.036 ;
  LAYER M2 ;
        RECT 5.792 12.068 5.824 12.1 ;
  LAYER M2 ;
        RECT 3.424 12.132 3.456 12.164 ;
  LAYER M2 ;
        RECT 5.792 12.196 5.824 12.228 ;
  LAYER M2 ;
        RECT 3.424 12.26 3.456 12.292 ;
  LAYER M2 ;
        RECT 5.792 12.324 5.824 12.356 ;
  LAYER M2 ;
        RECT 3.424 12.388 3.456 12.42 ;
  LAYER M2 ;
        RECT 5.792 12.452 5.824 12.484 ;
  LAYER M2 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M1 ;
        RECT 3.424 13.236 3.456 15.744 ;
  LAYER M3 ;
        RECT 3.424 15.692 3.456 15.724 ;
  LAYER M1 ;
        RECT 3.488 13.236 3.52 15.744 ;
  LAYER M3 ;
        RECT 3.488 13.256 3.52 13.288 ;
  LAYER M1 ;
        RECT 3.552 13.236 3.584 15.744 ;
  LAYER M3 ;
        RECT 3.552 15.692 3.584 15.724 ;
  LAYER M1 ;
        RECT 3.616 13.236 3.648 15.744 ;
  LAYER M3 ;
        RECT 3.616 13.256 3.648 13.288 ;
  LAYER M1 ;
        RECT 3.68 13.236 3.712 15.744 ;
  LAYER M3 ;
        RECT 3.68 15.692 3.712 15.724 ;
  LAYER M1 ;
        RECT 3.744 13.236 3.776 15.744 ;
  LAYER M3 ;
        RECT 3.744 13.256 3.776 13.288 ;
  LAYER M1 ;
        RECT 3.808 13.236 3.84 15.744 ;
  LAYER M3 ;
        RECT 3.808 15.692 3.84 15.724 ;
  LAYER M1 ;
        RECT 3.872 13.236 3.904 15.744 ;
  LAYER M3 ;
        RECT 3.872 13.256 3.904 13.288 ;
  LAYER M1 ;
        RECT 3.936 13.236 3.968 15.744 ;
  LAYER M3 ;
        RECT 3.936 15.692 3.968 15.724 ;
  LAYER M1 ;
        RECT 4 13.236 4.032 15.744 ;
  LAYER M3 ;
        RECT 4 13.256 4.032 13.288 ;
  LAYER M1 ;
        RECT 4.064 13.236 4.096 15.744 ;
  LAYER M3 ;
        RECT 4.064 15.692 4.096 15.724 ;
  LAYER M1 ;
        RECT 4.128 13.236 4.16 15.744 ;
  LAYER M3 ;
        RECT 4.128 13.256 4.16 13.288 ;
  LAYER M1 ;
        RECT 4.192 13.236 4.224 15.744 ;
  LAYER M3 ;
        RECT 4.192 15.692 4.224 15.724 ;
  LAYER M1 ;
        RECT 4.256 13.236 4.288 15.744 ;
  LAYER M3 ;
        RECT 4.256 13.256 4.288 13.288 ;
  LAYER M1 ;
        RECT 4.32 13.236 4.352 15.744 ;
  LAYER M3 ;
        RECT 4.32 15.692 4.352 15.724 ;
  LAYER M1 ;
        RECT 4.384 13.236 4.416 15.744 ;
  LAYER M3 ;
        RECT 4.384 13.256 4.416 13.288 ;
  LAYER M1 ;
        RECT 4.448 13.236 4.48 15.744 ;
  LAYER M3 ;
        RECT 4.448 15.692 4.48 15.724 ;
  LAYER M1 ;
        RECT 4.512 13.236 4.544 15.744 ;
  LAYER M3 ;
        RECT 4.512 13.256 4.544 13.288 ;
  LAYER M1 ;
        RECT 4.576 13.236 4.608 15.744 ;
  LAYER M3 ;
        RECT 4.576 15.692 4.608 15.724 ;
  LAYER M1 ;
        RECT 4.64 13.236 4.672 15.744 ;
  LAYER M3 ;
        RECT 4.64 13.256 4.672 13.288 ;
  LAYER M1 ;
        RECT 4.704 13.236 4.736 15.744 ;
  LAYER M3 ;
        RECT 4.704 15.692 4.736 15.724 ;
  LAYER M1 ;
        RECT 4.768 13.236 4.8 15.744 ;
  LAYER M3 ;
        RECT 4.768 13.256 4.8 13.288 ;
  LAYER M1 ;
        RECT 4.832 13.236 4.864 15.744 ;
  LAYER M3 ;
        RECT 4.832 15.692 4.864 15.724 ;
  LAYER M1 ;
        RECT 4.896 13.236 4.928 15.744 ;
  LAYER M3 ;
        RECT 4.896 13.256 4.928 13.288 ;
  LAYER M1 ;
        RECT 4.96 13.236 4.992 15.744 ;
  LAYER M3 ;
        RECT 4.96 15.692 4.992 15.724 ;
  LAYER M1 ;
        RECT 5.024 13.236 5.056 15.744 ;
  LAYER M3 ;
        RECT 5.024 13.256 5.056 13.288 ;
  LAYER M1 ;
        RECT 5.088 13.236 5.12 15.744 ;
  LAYER M3 ;
        RECT 5.088 15.692 5.12 15.724 ;
  LAYER M1 ;
        RECT 5.152 13.236 5.184 15.744 ;
  LAYER M3 ;
        RECT 5.152 13.256 5.184 13.288 ;
  LAYER M1 ;
        RECT 5.216 13.236 5.248 15.744 ;
  LAYER M3 ;
        RECT 5.216 15.692 5.248 15.724 ;
  LAYER M1 ;
        RECT 5.28 13.236 5.312 15.744 ;
  LAYER M3 ;
        RECT 5.28 13.256 5.312 13.288 ;
  LAYER M1 ;
        RECT 5.344 13.236 5.376 15.744 ;
  LAYER M3 ;
        RECT 5.344 15.692 5.376 15.724 ;
  LAYER M1 ;
        RECT 5.408 13.236 5.44 15.744 ;
  LAYER M3 ;
        RECT 5.408 13.256 5.44 13.288 ;
  LAYER M1 ;
        RECT 5.472 13.236 5.504 15.744 ;
  LAYER M3 ;
        RECT 5.472 15.692 5.504 15.724 ;
  LAYER M1 ;
        RECT 5.536 13.236 5.568 15.744 ;
  LAYER M3 ;
        RECT 5.536 13.256 5.568 13.288 ;
  LAYER M1 ;
        RECT 5.6 13.236 5.632 15.744 ;
  LAYER M3 ;
        RECT 5.6 15.692 5.632 15.724 ;
  LAYER M1 ;
        RECT 5.664 13.236 5.696 15.744 ;
  LAYER M3 ;
        RECT 5.664 13.256 5.696 13.288 ;
  LAYER M1 ;
        RECT 5.728 13.236 5.76 15.744 ;
  LAYER M3 ;
        RECT 5.728 15.692 5.76 15.724 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 15.744 ;
  LAYER M3 ;
        RECT 3.424 13.32 3.456 13.352 ;
  LAYER M2 ;
        RECT 5.792 13.384 5.824 13.416 ;
  LAYER M2 ;
        RECT 3.424 13.448 3.456 13.48 ;
  LAYER M2 ;
        RECT 5.792 13.512 5.824 13.544 ;
  LAYER M2 ;
        RECT 3.424 13.576 3.456 13.608 ;
  LAYER M2 ;
        RECT 5.792 13.64 5.824 13.672 ;
  LAYER M2 ;
        RECT 3.424 13.704 3.456 13.736 ;
  LAYER M2 ;
        RECT 5.792 13.768 5.824 13.8 ;
  LAYER M2 ;
        RECT 3.424 13.832 3.456 13.864 ;
  LAYER M2 ;
        RECT 5.792 13.896 5.824 13.928 ;
  LAYER M2 ;
        RECT 3.424 13.96 3.456 13.992 ;
  LAYER M2 ;
        RECT 5.792 14.024 5.824 14.056 ;
  LAYER M2 ;
        RECT 3.424 14.088 3.456 14.12 ;
  LAYER M2 ;
        RECT 5.792 14.152 5.824 14.184 ;
  LAYER M2 ;
        RECT 3.424 14.216 3.456 14.248 ;
  LAYER M2 ;
        RECT 5.792 14.28 5.824 14.312 ;
  LAYER M2 ;
        RECT 3.424 14.344 3.456 14.376 ;
  LAYER M2 ;
        RECT 5.792 14.408 5.824 14.44 ;
  LAYER M2 ;
        RECT 3.424 14.472 3.456 14.504 ;
  LAYER M2 ;
        RECT 5.792 14.536 5.824 14.568 ;
  LAYER M2 ;
        RECT 3.424 14.6 3.456 14.632 ;
  LAYER M2 ;
        RECT 5.792 14.664 5.824 14.696 ;
  LAYER M2 ;
        RECT 3.424 14.728 3.456 14.76 ;
  LAYER M2 ;
        RECT 5.792 14.792 5.824 14.824 ;
  LAYER M2 ;
        RECT 3.424 14.856 3.456 14.888 ;
  LAYER M2 ;
        RECT 5.792 14.92 5.824 14.952 ;
  LAYER M2 ;
        RECT 3.424 14.984 3.456 15.016 ;
  LAYER M2 ;
        RECT 5.792 15.048 5.824 15.08 ;
  LAYER M2 ;
        RECT 3.424 15.112 3.456 15.144 ;
  LAYER M2 ;
        RECT 5.792 15.176 5.824 15.208 ;
  LAYER M2 ;
        RECT 3.424 15.24 3.456 15.272 ;
  LAYER M2 ;
        RECT 5.792 15.304 5.824 15.336 ;
  LAYER M2 ;
        RECT 3.424 15.368 3.456 15.4 ;
  LAYER M2 ;
        RECT 5.792 15.432 5.824 15.464 ;
  LAYER M2 ;
        RECT 3.424 15.496 3.456 15.528 ;
  LAYER M2 ;
        RECT 5.792 15.56 5.824 15.592 ;
  LAYER M2 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M1 ;
        RECT 3.424 16.344 3.456 18.852 ;
  LAYER M3 ;
        RECT 3.424 18.8 3.456 18.832 ;
  LAYER M1 ;
        RECT 3.488 16.344 3.52 18.852 ;
  LAYER M3 ;
        RECT 3.488 16.364 3.52 16.396 ;
  LAYER M1 ;
        RECT 3.552 16.344 3.584 18.852 ;
  LAYER M3 ;
        RECT 3.552 18.8 3.584 18.832 ;
  LAYER M1 ;
        RECT 3.616 16.344 3.648 18.852 ;
  LAYER M3 ;
        RECT 3.616 16.364 3.648 16.396 ;
  LAYER M1 ;
        RECT 3.68 16.344 3.712 18.852 ;
  LAYER M3 ;
        RECT 3.68 18.8 3.712 18.832 ;
  LAYER M1 ;
        RECT 3.744 16.344 3.776 18.852 ;
  LAYER M3 ;
        RECT 3.744 16.364 3.776 16.396 ;
  LAYER M1 ;
        RECT 3.808 16.344 3.84 18.852 ;
  LAYER M3 ;
        RECT 3.808 18.8 3.84 18.832 ;
  LAYER M1 ;
        RECT 3.872 16.344 3.904 18.852 ;
  LAYER M3 ;
        RECT 3.872 16.364 3.904 16.396 ;
  LAYER M1 ;
        RECT 3.936 16.344 3.968 18.852 ;
  LAYER M3 ;
        RECT 3.936 18.8 3.968 18.832 ;
  LAYER M1 ;
        RECT 4 16.344 4.032 18.852 ;
  LAYER M3 ;
        RECT 4 16.364 4.032 16.396 ;
  LAYER M1 ;
        RECT 4.064 16.344 4.096 18.852 ;
  LAYER M3 ;
        RECT 4.064 18.8 4.096 18.832 ;
  LAYER M1 ;
        RECT 4.128 16.344 4.16 18.852 ;
  LAYER M3 ;
        RECT 4.128 16.364 4.16 16.396 ;
  LAYER M1 ;
        RECT 4.192 16.344 4.224 18.852 ;
  LAYER M3 ;
        RECT 4.192 18.8 4.224 18.832 ;
  LAYER M1 ;
        RECT 4.256 16.344 4.288 18.852 ;
  LAYER M3 ;
        RECT 4.256 16.364 4.288 16.396 ;
  LAYER M1 ;
        RECT 4.32 16.344 4.352 18.852 ;
  LAYER M3 ;
        RECT 4.32 18.8 4.352 18.832 ;
  LAYER M1 ;
        RECT 4.384 16.344 4.416 18.852 ;
  LAYER M3 ;
        RECT 4.384 16.364 4.416 16.396 ;
  LAYER M1 ;
        RECT 4.448 16.344 4.48 18.852 ;
  LAYER M3 ;
        RECT 4.448 18.8 4.48 18.832 ;
  LAYER M1 ;
        RECT 4.512 16.344 4.544 18.852 ;
  LAYER M3 ;
        RECT 4.512 16.364 4.544 16.396 ;
  LAYER M1 ;
        RECT 4.576 16.344 4.608 18.852 ;
  LAYER M3 ;
        RECT 4.576 18.8 4.608 18.832 ;
  LAYER M1 ;
        RECT 4.64 16.344 4.672 18.852 ;
  LAYER M3 ;
        RECT 4.64 16.364 4.672 16.396 ;
  LAYER M1 ;
        RECT 4.704 16.344 4.736 18.852 ;
  LAYER M3 ;
        RECT 4.704 18.8 4.736 18.832 ;
  LAYER M1 ;
        RECT 4.768 16.344 4.8 18.852 ;
  LAYER M3 ;
        RECT 4.768 16.364 4.8 16.396 ;
  LAYER M1 ;
        RECT 4.832 16.344 4.864 18.852 ;
  LAYER M3 ;
        RECT 4.832 18.8 4.864 18.832 ;
  LAYER M1 ;
        RECT 4.896 16.344 4.928 18.852 ;
  LAYER M3 ;
        RECT 4.896 16.364 4.928 16.396 ;
  LAYER M1 ;
        RECT 4.96 16.344 4.992 18.852 ;
  LAYER M3 ;
        RECT 4.96 18.8 4.992 18.832 ;
  LAYER M1 ;
        RECT 5.024 16.344 5.056 18.852 ;
  LAYER M3 ;
        RECT 5.024 16.364 5.056 16.396 ;
  LAYER M1 ;
        RECT 5.088 16.344 5.12 18.852 ;
  LAYER M3 ;
        RECT 5.088 18.8 5.12 18.832 ;
  LAYER M1 ;
        RECT 5.152 16.344 5.184 18.852 ;
  LAYER M3 ;
        RECT 5.152 16.364 5.184 16.396 ;
  LAYER M1 ;
        RECT 5.216 16.344 5.248 18.852 ;
  LAYER M3 ;
        RECT 5.216 18.8 5.248 18.832 ;
  LAYER M1 ;
        RECT 5.28 16.344 5.312 18.852 ;
  LAYER M3 ;
        RECT 5.28 16.364 5.312 16.396 ;
  LAYER M1 ;
        RECT 5.344 16.344 5.376 18.852 ;
  LAYER M3 ;
        RECT 5.344 18.8 5.376 18.832 ;
  LAYER M1 ;
        RECT 5.408 16.344 5.44 18.852 ;
  LAYER M3 ;
        RECT 5.408 16.364 5.44 16.396 ;
  LAYER M1 ;
        RECT 5.472 16.344 5.504 18.852 ;
  LAYER M3 ;
        RECT 5.472 18.8 5.504 18.832 ;
  LAYER M1 ;
        RECT 5.536 16.344 5.568 18.852 ;
  LAYER M3 ;
        RECT 5.536 16.364 5.568 16.396 ;
  LAYER M1 ;
        RECT 5.6 16.344 5.632 18.852 ;
  LAYER M3 ;
        RECT 5.6 18.8 5.632 18.832 ;
  LAYER M1 ;
        RECT 5.664 16.344 5.696 18.852 ;
  LAYER M3 ;
        RECT 5.664 16.364 5.696 16.396 ;
  LAYER M1 ;
        RECT 5.728 16.344 5.76 18.852 ;
  LAYER M3 ;
        RECT 5.728 18.8 5.76 18.832 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 18.852 ;
  LAYER M3 ;
        RECT 3.424 16.428 3.456 16.46 ;
  LAYER M2 ;
        RECT 5.792 16.492 5.824 16.524 ;
  LAYER M2 ;
        RECT 3.424 16.556 3.456 16.588 ;
  LAYER M2 ;
        RECT 5.792 16.62 5.824 16.652 ;
  LAYER M2 ;
        RECT 3.424 16.684 3.456 16.716 ;
  LAYER M2 ;
        RECT 5.792 16.748 5.824 16.78 ;
  LAYER M2 ;
        RECT 3.424 16.812 3.456 16.844 ;
  LAYER M2 ;
        RECT 5.792 16.876 5.824 16.908 ;
  LAYER M2 ;
        RECT 3.424 16.94 3.456 16.972 ;
  LAYER M2 ;
        RECT 5.792 17.004 5.824 17.036 ;
  LAYER M2 ;
        RECT 3.424 17.068 3.456 17.1 ;
  LAYER M2 ;
        RECT 5.792 17.132 5.824 17.164 ;
  LAYER M2 ;
        RECT 3.424 17.196 3.456 17.228 ;
  LAYER M2 ;
        RECT 5.792 17.26 5.824 17.292 ;
  LAYER M2 ;
        RECT 3.424 17.324 3.456 17.356 ;
  LAYER M2 ;
        RECT 5.792 17.388 5.824 17.42 ;
  LAYER M2 ;
        RECT 3.424 17.452 3.456 17.484 ;
  LAYER M2 ;
        RECT 5.792 17.516 5.824 17.548 ;
  LAYER M2 ;
        RECT 3.424 17.58 3.456 17.612 ;
  LAYER M2 ;
        RECT 5.792 17.644 5.824 17.676 ;
  LAYER M2 ;
        RECT 3.424 17.708 3.456 17.74 ;
  LAYER M2 ;
        RECT 5.792 17.772 5.824 17.804 ;
  LAYER M2 ;
        RECT 3.424 17.836 3.456 17.868 ;
  LAYER M2 ;
        RECT 5.792 17.9 5.824 17.932 ;
  LAYER M2 ;
        RECT 3.424 17.964 3.456 17.996 ;
  LAYER M2 ;
        RECT 5.792 18.028 5.824 18.06 ;
  LAYER M2 ;
        RECT 3.424 18.092 3.456 18.124 ;
  LAYER M2 ;
        RECT 5.792 18.156 5.824 18.188 ;
  LAYER M2 ;
        RECT 3.424 18.22 3.456 18.252 ;
  LAYER M2 ;
        RECT 5.792 18.284 5.824 18.316 ;
  LAYER M2 ;
        RECT 3.424 18.348 3.456 18.38 ;
  LAYER M2 ;
        RECT 5.792 18.412 5.824 18.444 ;
  LAYER M2 ;
        RECT 3.424 18.476 3.456 18.508 ;
  LAYER M2 ;
        RECT 5.792 18.54 5.824 18.572 ;
  LAYER M2 ;
        RECT 3.424 18.604 3.456 18.636 ;
  LAYER M2 ;
        RECT 5.792 18.668 5.824 18.7 ;
  LAYER M2 ;
        RECT 3.376 16.296 5.872 18.9 ;
  LAYER M1 ;
        RECT 3.424 19.452 3.456 21.96 ;
  LAYER M3 ;
        RECT 3.424 21.908 3.456 21.94 ;
  LAYER M1 ;
        RECT 3.488 19.452 3.52 21.96 ;
  LAYER M3 ;
        RECT 3.488 19.472 3.52 19.504 ;
  LAYER M1 ;
        RECT 3.552 19.452 3.584 21.96 ;
  LAYER M3 ;
        RECT 3.552 21.908 3.584 21.94 ;
  LAYER M1 ;
        RECT 3.616 19.452 3.648 21.96 ;
  LAYER M3 ;
        RECT 3.616 19.472 3.648 19.504 ;
  LAYER M1 ;
        RECT 3.68 19.452 3.712 21.96 ;
  LAYER M3 ;
        RECT 3.68 21.908 3.712 21.94 ;
  LAYER M1 ;
        RECT 3.744 19.452 3.776 21.96 ;
  LAYER M3 ;
        RECT 3.744 19.472 3.776 19.504 ;
  LAYER M1 ;
        RECT 3.808 19.452 3.84 21.96 ;
  LAYER M3 ;
        RECT 3.808 21.908 3.84 21.94 ;
  LAYER M1 ;
        RECT 3.872 19.452 3.904 21.96 ;
  LAYER M3 ;
        RECT 3.872 19.472 3.904 19.504 ;
  LAYER M1 ;
        RECT 3.936 19.452 3.968 21.96 ;
  LAYER M3 ;
        RECT 3.936 21.908 3.968 21.94 ;
  LAYER M1 ;
        RECT 4 19.452 4.032 21.96 ;
  LAYER M3 ;
        RECT 4 19.472 4.032 19.504 ;
  LAYER M1 ;
        RECT 4.064 19.452 4.096 21.96 ;
  LAYER M3 ;
        RECT 4.064 21.908 4.096 21.94 ;
  LAYER M1 ;
        RECT 4.128 19.452 4.16 21.96 ;
  LAYER M3 ;
        RECT 4.128 19.472 4.16 19.504 ;
  LAYER M1 ;
        RECT 4.192 19.452 4.224 21.96 ;
  LAYER M3 ;
        RECT 4.192 21.908 4.224 21.94 ;
  LAYER M1 ;
        RECT 4.256 19.452 4.288 21.96 ;
  LAYER M3 ;
        RECT 4.256 19.472 4.288 19.504 ;
  LAYER M1 ;
        RECT 4.32 19.452 4.352 21.96 ;
  LAYER M3 ;
        RECT 4.32 21.908 4.352 21.94 ;
  LAYER M1 ;
        RECT 4.384 19.452 4.416 21.96 ;
  LAYER M3 ;
        RECT 4.384 19.472 4.416 19.504 ;
  LAYER M1 ;
        RECT 4.448 19.452 4.48 21.96 ;
  LAYER M3 ;
        RECT 4.448 21.908 4.48 21.94 ;
  LAYER M1 ;
        RECT 4.512 19.452 4.544 21.96 ;
  LAYER M3 ;
        RECT 4.512 19.472 4.544 19.504 ;
  LAYER M1 ;
        RECT 4.576 19.452 4.608 21.96 ;
  LAYER M3 ;
        RECT 4.576 21.908 4.608 21.94 ;
  LAYER M1 ;
        RECT 4.64 19.452 4.672 21.96 ;
  LAYER M3 ;
        RECT 4.64 19.472 4.672 19.504 ;
  LAYER M1 ;
        RECT 4.704 19.452 4.736 21.96 ;
  LAYER M3 ;
        RECT 4.704 21.908 4.736 21.94 ;
  LAYER M1 ;
        RECT 4.768 19.452 4.8 21.96 ;
  LAYER M3 ;
        RECT 4.768 19.472 4.8 19.504 ;
  LAYER M1 ;
        RECT 4.832 19.452 4.864 21.96 ;
  LAYER M3 ;
        RECT 4.832 21.908 4.864 21.94 ;
  LAYER M1 ;
        RECT 4.896 19.452 4.928 21.96 ;
  LAYER M3 ;
        RECT 4.896 19.472 4.928 19.504 ;
  LAYER M1 ;
        RECT 4.96 19.452 4.992 21.96 ;
  LAYER M3 ;
        RECT 4.96 21.908 4.992 21.94 ;
  LAYER M1 ;
        RECT 5.024 19.452 5.056 21.96 ;
  LAYER M3 ;
        RECT 5.024 19.472 5.056 19.504 ;
  LAYER M1 ;
        RECT 5.088 19.452 5.12 21.96 ;
  LAYER M3 ;
        RECT 5.088 21.908 5.12 21.94 ;
  LAYER M1 ;
        RECT 5.152 19.452 5.184 21.96 ;
  LAYER M3 ;
        RECT 5.152 19.472 5.184 19.504 ;
  LAYER M1 ;
        RECT 5.216 19.452 5.248 21.96 ;
  LAYER M3 ;
        RECT 5.216 21.908 5.248 21.94 ;
  LAYER M1 ;
        RECT 5.28 19.452 5.312 21.96 ;
  LAYER M3 ;
        RECT 5.28 19.472 5.312 19.504 ;
  LAYER M1 ;
        RECT 5.344 19.452 5.376 21.96 ;
  LAYER M3 ;
        RECT 5.344 21.908 5.376 21.94 ;
  LAYER M1 ;
        RECT 5.408 19.452 5.44 21.96 ;
  LAYER M3 ;
        RECT 5.408 19.472 5.44 19.504 ;
  LAYER M1 ;
        RECT 5.472 19.452 5.504 21.96 ;
  LAYER M3 ;
        RECT 5.472 21.908 5.504 21.94 ;
  LAYER M1 ;
        RECT 5.536 19.452 5.568 21.96 ;
  LAYER M3 ;
        RECT 5.536 19.472 5.568 19.504 ;
  LAYER M1 ;
        RECT 5.6 19.452 5.632 21.96 ;
  LAYER M3 ;
        RECT 5.6 21.908 5.632 21.94 ;
  LAYER M1 ;
        RECT 5.664 19.452 5.696 21.96 ;
  LAYER M3 ;
        RECT 5.664 19.472 5.696 19.504 ;
  LAYER M1 ;
        RECT 5.728 19.452 5.76 21.96 ;
  LAYER M3 ;
        RECT 5.728 21.908 5.76 21.94 ;
  LAYER M1 ;
        RECT 5.792 19.452 5.824 21.96 ;
  LAYER M3 ;
        RECT 3.424 19.536 3.456 19.568 ;
  LAYER M2 ;
        RECT 5.792 19.6 5.824 19.632 ;
  LAYER M2 ;
        RECT 3.424 19.664 3.456 19.696 ;
  LAYER M2 ;
        RECT 5.792 19.728 5.824 19.76 ;
  LAYER M2 ;
        RECT 3.424 19.792 3.456 19.824 ;
  LAYER M2 ;
        RECT 5.792 19.856 5.824 19.888 ;
  LAYER M2 ;
        RECT 3.424 19.92 3.456 19.952 ;
  LAYER M2 ;
        RECT 5.792 19.984 5.824 20.016 ;
  LAYER M2 ;
        RECT 3.424 20.048 3.456 20.08 ;
  LAYER M2 ;
        RECT 5.792 20.112 5.824 20.144 ;
  LAYER M2 ;
        RECT 3.424 20.176 3.456 20.208 ;
  LAYER M2 ;
        RECT 5.792 20.24 5.824 20.272 ;
  LAYER M2 ;
        RECT 3.424 20.304 3.456 20.336 ;
  LAYER M2 ;
        RECT 5.792 20.368 5.824 20.4 ;
  LAYER M2 ;
        RECT 3.424 20.432 3.456 20.464 ;
  LAYER M2 ;
        RECT 5.792 20.496 5.824 20.528 ;
  LAYER M2 ;
        RECT 3.424 20.56 3.456 20.592 ;
  LAYER M2 ;
        RECT 5.792 20.624 5.824 20.656 ;
  LAYER M2 ;
        RECT 3.424 20.688 3.456 20.72 ;
  LAYER M2 ;
        RECT 5.792 20.752 5.824 20.784 ;
  LAYER M2 ;
        RECT 3.424 20.816 3.456 20.848 ;
  LAYER M2 ;
        RECT 5.792 20.88 5.824 20.912 ;
  LAYER M2 ;
        RECT 3.424 20.944 3.456 20.976 ;
  LAYER M2 ;
        RECT 5.792 21.008 5.824 21.04 ;
  LAYER M2 ;
        RECT 3.424 21.072 3.456 21.104 ;
  LAYER M2 ;
        RECT 5.792 21.136 5.824 21.168 ;
  LAYER M2 ;
        RECT 3.424 21.2 3.456 21.232 ;
  LAYER M2 ;
        RECT 5.792 21.264 5.824 21.296 ;
  LAYER M2 ;
        RECT 3.424 21.328 3.456 21.36 ;
  LAYER M2 ;
        RECT 5.792 21.392 5.824 21.424 ;
  LAYER M2 ;
        RECT 3.424 21.456 3.456 21.488 ;
  LAYER M2 ;
        RECT 5.792 21.52 5.824 21.552 ;
  LAYER M2 ;
        RECT 3.424 21.584 3.456 21.616 ;
  LAYER M2 ;
        RECT 5.792 21.648 5.824 21.68 ;
  LAYER M2 ;
        RECT 3.424 21.712 3.456 21.744 ;
  LAYER M2 ;
        RECT 5.792 21.776 5.824 21.808 ;
  LAYER M2 ;
        RECT 3.376 19.404 5.872 22.008 ;
  LAYER M1 ;
        RECT 3.424 22.56 3.456 25.068 ;
  LAYER M3 ;
        RECT 3.424 25.016 3.456 25.048 ;
  LAYER M1 ;
        RECT 3.488 22.56 3.52 25.068 ;
  LAYER M3 ;
        RECT 3.488 22.58 3.52 22.612 ;
  LAYER M1 ;
        RECT 3.552 22.56 3.584 25.068 ;
  LAYER M3 ;
        RECT 3.552 25.016 3.584 25.048 ;
  LAYER M1 ;
        RECT 3.616 22.56 3.648 25.068 ;
  LAYER M3 ;
        RECT 3.616 22.58 3.648 22.612 ;
  LAYER M1 ;
        RECT 3.68 22.56 3.712 25.068 ;
  LAYER M3 ;
        RECT 3.68 25.016 3.712 25.048 ;
  LAYER M1 ;
        RECT 3.744 22.56 3.776 25.068 ;
  LAYER M3 ;
        RECT 3.744 22.58 3.776 22.612 ;
  LAYER M1 ;
        RECT 3.808 22.56 3.84 25.068 ;
  LAYER M3 ;
        RECT 3.808 25.016 3.84 25.048 ;
  LAYER M1 ;
        RECT 3.872 22.56 3.904 25.068 ;
  LAYER M3 ;
        RECT 3.872 22.58 3.904 22.612 ;
  LAYER M1 ;
        RECT 3.936 22.56 3.968 25.068 ;
  LAYER M3 ;
        RECT 3.936 25.016 3.968 25.048 ;
  LAYER M1 ;
        RECT 4 22.56 4.032 25.068 ;
  LAYER M3 ;
        RECT 4 22.58 4.032 22.612 ;
  LAYER M1 ;
        RECT 4.064 22.56 4.096 25.068 ;
  LAYER M3 ;
        RECT 4.064 25.016 4.096 25.048 ;
  LAYER M1 ;
        RECT 4.128 22.56 4.16 25.068 ;
  LAYER M3 ;
        RECT 4.128 22.58 4.16 22.612 ;
  LAYER M1 ;
        RECT 4.192 22.56 4.224 25.068 ;
  LAYER M3 ;
        RECT 4.192 25.016 4.224 25.048 ;
  LAYER M1 ;
        RECT 4.256 22.56 4.288 25.068 ;
  LAYER M3 ;
        RECT 4.256 22.58 4.288 22.612 ;
  LAYER M1 ;
        RECT 4.32 22.56 4.352 25.068 ;
  LAYER M3 ;
        RECT 4.32 25.016 4.352 25.048 ;
  LAYER M1 ;
        RECT 4.384 22.56 4.416 25.068 ;
  LAYER M3 ;
        RECT 4.384 22.58 4.416 22.612 ;
  LAYER M1 ;
        RECT 4.448 22.56 4.48 25.068 ;
  LAYER M3 ;
        RECT 4.448 25.016 4.48 25.048 ;
  LAYER M1 ;
        RECT 4.512 22.56 4.544 25.068 ;
  LAYER M3 ;
        RECT 4.512 22.58 4.544 22.612 ;
  LAYER M1 ;
        RECT 4.576 22.56 4.608 25.068 ;
  LAYER M3 ;
        RECT 4.576 25.016 4.608 25.048 ;
  LAYER M1 ;
        RECT 4.64 22.56 4.672 25.068 ;
  LAYER M3 ;
        RECT 4.64 22.58 4.672 22.612 ;
  LAYER M1 ;
        RECT 4.704 22.56 4.736 25.068 ;
  LAYER M3 ;
        RECT 4.704 25.016 4.736 25.048 ;
  LAYER M1 ;
        RECT 4.768 22.56 4.8 25.068 ;
  LAYER M3 ;
        RECT 4.768 22.58 4.8 22.612 ;
  LAYER M1 ;
        RECT 4.832 22.56 4.864 25.068 ;
  LAYER M3 ;
        RECT 4.832 25.016 4.864 25.048 ;
  LAYER M1 ;
        RECT 4.896 22.56 4.928 25.068 ;
  LAYER M3 ;
        RECT 4.896 22.58 4.928 22.612 ;
  LAYER M1 ;
        RECT 4.96 22.56 4.992 25.068 ;
  LAYER M3 ;
        RECT 4.96 25.016 4.992 25.048 ;
  LAYER M1 ;
        RECT 5.024 22.56 5.056 25.068 ;
  LAYER M3 ;
        RECT 5.024 22.58 5.056 22.612 ;
  LAYER M1 ;
        RECT 5.088 22.56 5.12 25.068 ;
  LAYER M3 ;
        RECT 5.088 25.016 5.12 25.048 ;
  LAYER M1 ;
        RECT 5.152 22.56 5.184 25.068 ;
  LAYER M3 ;
        RECT 5.152 22.58 5.184 22.612 ;
  LAYER M1 ;
        RECT 5.216 22.56 5.248 25.068 ;
  LAYER M3 ;
        RECT 5.216 25.016 5.248 25.048 ;
  LAYER M1 ;
        RECT 5.28 22.56 5.312 25.068 ;
  LAYER M3 ;
        RECT 5.28 22.58 5.312 22.612 ;
  LAYER M1 ;
        RECT 5.344 22.56 5.376 25.068 ;
  LAYER M3 ;
        RECT 5.344 25.016 5.376 25.048 ;
  LAYER M1 ;
        RECT 5.408 22.56 5.44 25.068 ;
  LAYER M3 ;
        RECT 5.408 22.58 5.44 22.612 ;
  LAYER M1 ;
        RECT 5.472 22.56 5.504 25.068 ;
  LAYER M3 ;
        RECT 5.472 25.016 5.504 25.048 ;
  LAYER M1 ;
        RECT 5.536 22.56 5.568 25.068 ;
  LAYER M3 ;
        RECT 5.536 22.58 5.568 22.612 ;
  LAYER M1 ;
        RECT 5.6 22.56 5.632 25.068 ;
  LAYER M3 ;
        RECT 5.6 25.016 5.632 25.048 ;
  LAYER M1 ;
        RECT 5.664 22.56 5.696 25.068 ;
  LAYER M3 ;
        RECT 5.664 22.58 5.696 22.612 ;
  LAYER M1 ;
        RECT 5.728 22.56 5.76 25.068 ;
  LAYER M3 ;
        RECT 5.728 25.016 5.76 25.048 ;
  LAYER M1 ;
        RECT 5.792 22.56 5.824 25.068 ;
  LAYER M3 ;
        RECT 3.424 22.644 3.456 22.676 ;
  LAYER M2 ;
        RECT 5.792 22.708 5.824 22.74 ;
  LAYER M2 ;
        RECT 3.424 22.772 3.456 22.804 ;
  LAYER M2 ;
        RECT 5.792 22.836 5.824 22.868 ;
  LAYER M2 ;
        RECT 3.424 22.9 3.456 22.932 ;
  LAYER M2 ;
        RECT 5.792 22.964 5.824 22.996 ;
  LAYER M2 ;
        RECT 3.424 23.028 3.456 23.06 ;
  LAYER M2 ;
        RECT 5.792 23.092 5.824 23.124 ;
  LAYER M2 ;
        RECT 3.424 23.156 3.456 23.188 ;
  LAYER M2 ;
        RECT 5.792 23.22 5.824 23.252 ;
  LAYER M2 ;
        RECT 3.424 23.284 3.456 23.316 ;
  LAYER M2 ;
        RECT 5.792 23.348 5.824 23.38 ;
  LAYER M2 ;
        RECT 3.424 23.412 3.456 23.444 ;
  LAYER M2 ;
        RECT 5.792 23.476 5.824 23.508 ;
  LAYER M2 ;
        RECT 3.424 23.54 3.456 23.572 ;
  LAYER M2 ;
        RECT 5.792 23.604 5.824 23.636 ;
  LAYER M2 ;
        RECT 3.424 23.668 3.456 23.7 ;
  LAYER M2 ;
        RECT 5.792 23.732 5.824 23.764 ;
  LAYER M2 ;
        RECT 3.424 23.796 3.456 23.828 ;
  LAYER M2 ;
        RECT 5.792 23.86 5.824 23.892 ;
  LAYER M2 ;
        RECT 3.424 23.924 3.456 23.956 ;
  LAYER M2 ;
        RECT 5.792 23.988 5.824 24.02 ;
  LAYER M2 ;
        RECT 3.424 24.052 3.456 24.084 ;
  LAYER M2 ;
        RECT 5.792 24.116 5.824 24.148 ;
  LAYER M2 ;
        RECT 3.424 24.18 3.456 24.212 ;
  LAYER M2 ;
        RECT 5.792 24.244 5.824 24.276 ;
  LAYER M2 ;
        RECT 3.424 24.308 3.456 24.34 ;
  LAYER M2 ;
        RECT 5.792 24.372 5.824 24.404 ;
  LAYER M2 ;
        RECT 3.424 24.436 3.456 24.468 ;
  LAYER M2 ;
        RECT 5.792 24.5 5.824 24.532 ;
  LAYER M2 ;
        RECT 3.424 24.564 3.456 24.596 ;
  LAYER M2 ;
        RECT 5.792 24.628 5.824 24.66 ;
  LAYER M2 ;
        RECT 3.424 24.692 3.456 24.724 ;
  LAYER M2 ;
        RECT 5.792 24.756 5.824 24.788 ;
  LAYER M2 ;
        RECT 3.424 24.82 3.456 24.852 ;
  LAYER M2 ;
        RECT 5.792 24.884 5.824 24.916 ;
  LAYER M2 ;
        RECT 3.376 22.512 5.872 25.116 ;
  LAYER M1 ;
        RECT 6.4 0.804 6.432 3.312 ;
  LAYER M3 ;
        RECT 6.4 3.26 6.432 3.292 ;
  LAYER M1 ;
        RECT 6.464 0.804 6.496 3.312 ;
  LAYER M3 ;
        RECT 6.464 0.824 6.496 0.856 ;
  LAYER M1 ;
        RECT 6.528 0.804 6.56 3.312 ;
  LAYER M3 ;
        RECT 6.528 3.26 6.56 3.292 ;
  LAYER M1 ;
        RECT 6.592 0.804 6.624 3.312 ;
  LAYER M3 ;
        RECT 6.592 0.824 6.624 0.856 ;
  LAYER M1 ;
        RECT 6.656 0.804 6.688 3.312 ;
  LAYER M3 ;
        RECT 6.656 3.26 6.688 3.292 ;
  LAYER M1 ;
        RECT 6.72 0.804 6.752 3.312 ;
  LAYER M3 ;
        RECT 6.72 0.824 6.752 0.856 ;
  LAYER M1 ;
        RECT 6.784 0.804 6.816 3.312 ;
  LAYER M3 ;
        RECT 6.784 3.26 6.816 3.292 ;
  LAYER M1 ;
        RECT 6.848 0.804 6.88 3.312 ;
  LAYER M3 ;
        RECT 6.848 0.824 6.88 0.856 ;
  LAYER M1 ;
        RECT 6.912 0.804 6.944 3.312 ;
  LAYER M3 ;
        RECT 6.912 3.26 6.944 3.292 ;
  LAYER M1 ;
        RECT 6.976 0.804 7.008 3.312 ;
  LAYER M3 ;
        RECT 6.976 0.824 7.008 0.856 ;
  LAYER M1 ;
        RECT 7.04 0.804 7.072 3.312 ;
  LAYER M3 ;
        RECT 7.04 3.26 7.072 3.292 ;
  LAYER M1 ;
        RECT 7.104 0.804 7.136 3.312 ;
  LAYER M3 ;
        RECT 7.104 0.824 7.136 0.856 ;
  LAYER M1 ;
        RECT 7.168 0.804 7.2 3.312 ;
  LAYER M3 ;
        RECT 7.168 3.26 7.2 3.292 ;
  LAYER M1 ;
        RECT 7.232 0.804 7.264 3.312 ;
  LAYER M3 ;
        RECT 7.232 0.824 7.264 0.856 ;
  LAYER M1 ;
        RECT 7.296 0.804 7.328 3.312 ;
  LAYER M3 ;
        RECT 7.296 3.26 7.328 3.292 ;
  LAYER M1 ;
        RECT 7.36 0.804 7.392 3.312 ;
  LAYER M3 ;
        RECT 7.36 0.824 7.392 0.856 ;
  LAYER M1 ;
        RECT 7.424 0.804 7.456 3.312 ;
  LAYER M3 ;
        RECT 7.424 3.26 7.456 3.292 ;
  LAYER M1 ;
        RECT 7.488 0.804 7.52 3.312 ;
  LAYER M3 ;
        RECT 7.488 0.824 7.52 0.856 ;
  LAYER M1 ;
        RECT 7.552 0.804 7.584 3.312 ;
  LAYER M3 ;
        RECT 7.552 3.26 7.584 3.292 ;
  LAYER M1 ;
        RECT 7.616 0.804 7.648 3.312 ;
  LAYER M3 ;
        RECT 7.616 0.824 7.648 0.856 ;
  LAYER M1 ;
        RECT 7.68 0.804 7.712 3.312 ;
  LAYER M3 ;
        RECT 7.68 3.26 7.712 3.292 ;
  LAYER M1 ;
        RECT 7.744 0.804 7.776 3.312 ;
  LAYER M3 ;
        RECT 7.744 0.824 7.776 0.856 ;
  LAYER M1 ;
        RECT 7.808 0.804 7.84 3.312 ;
  LAYER M3 ;
        RECT 7.808 3.26 7.84 3.292 ;
  LAYER M1 ;
        RECT 7.872 0.804 7.904 3.312 ;
  LAYER M3 ;
        RECT 7.872 0.824 7.904 0.856 ;
  LAYER M1 ;
        RECT 7.936 0.804 7.968 3.312 ;
  LAYER M3 ;
        RECT 7.936 3.26 7.968 3.292 ;
  LAYER M1 ;
        RECT 8 0.804 8.032 3.312 ;
  LAYER M3 ;
        RECT 8 0.824 8.032 0.856 ;
  LAYER M1 ;
        RECT 8.064 0.804 8.096 3.312 ;
  LAYER M3 ;
        RECT 8.064 3.26 8.096 3.292 ;
  LAYER M1 ;
        RECT 8.128 0.804 8.16 3.312 ;
  LAYER M3 ;
        RECT 8.128 0.824 8.16 0.856 ;
  LAYER M1 ;
        RECT 8.192 0.804 8.224 3.312 ;
  LAYER M3 ;
        RECT 8.192 3.26 8.224 3.292 ;
  LAYER M1 ;
        RECT 8.256 0.804 8.288 3.312 ;
  LAYER M3 ;
        RECT 8.256 0.824 8.288 0.856 ;
  LAYER M1 ;
        RECT 8.32 0.804 8.352 3.312 ;
  LAYER M3 ;
        RECT 8.32 3.26 8.352 3.292 ;
  LAYER M1 ;
        RECT 8.384 0.804 8.416 3.312 ;
  LAYER M3 ;
        RECT 8.384 0.824 8.416 0.856 ;
  LAYER M1 ;
        RECT 8.448 0.804 8.48 3.312 ;
  LAYER M3 ;
        RECT 8.448 3.26 8.48 3.292 ;
  LAYER M1 ;
        RECT 8.512 0.804 8.544 3.312 ;
  LAYER M3 ;
        RECT 8.512 0.824 8.544 0.856 ;
  LAYER M1 ;
        RECT 8.576 0.804 8.608 3.312 ;
  LAYER M3 ;
        RECT 8.576 3.26 8.608 3.292 ;
  LAYER M1 ;
        RECT 8.64 0.804 8.672 3.312 ;
  LAYER M3 ;
        RECT 8.64 0.824 8.672 0.856 ;
  LAYER M1 ;
        RECT 8.704 0.804 8.736 3.312 ;
  LAYER M3 ;
        RECT 8.704 3.26 8.736 3.292 ;
  LAYER M1 ;
        RECT 8.768 0.804 8.8 3.312 ;
  LAYER M3 ;
        RECT 6.4 0.888 6.432 0.92 ;
  LAYER M2 ;
        RECT 8.768 0.952 8.8 0.984 ;
  LAYER M2 ;
        RECT 6.4 1.016 6.432 1.048 ;
  LAYER M2 ;
        RECT 8.768 1.08 8.8 1.112 ;
  LAYER M2 ;
        RECT 6.4 1.144 6.432 1.176 ;
  LAYER M2 ;
        RECT 8.768 1.208 8.8 1.24 ;
  LAYER M2 ;
        RECT 6.4 1.272 6.432 1.304 ;
  LAYER M2 ;
        RECT 8.768 1.336 8.8 1.368 ;
  LAYER M2 ;
        RECT 6.4 1.4 6.432 1.432 ;
  LAYER M2 ;
        RECT 8.768 1.464 8.8 1.496 ;
  LAYER M2 ;
        RECT 6.4 1.528 6.432 1.56 ;
  LAYER M2 ;
        RECT 8.768 1.592 8.8 1.624 ;
  LAYER M2 ;
        RECT 6.4 1.656 6.432 1.688 ;
  LAYER M2 ;
        RECT 8.768 1.72 8.8 1.752 ;
  LAYER M2 ;
        RECT 6.4 1.784 6.432 1.816 ;
  LAYER M2 ;
        RECT 8.768 1.848 8.8 1.88 ;
  LAYER M2 ;
        RECT 6.4 1.912 6.432 1.944 ;
  LAYER M2 ;
        RECT 8.768 1.976 8.8 2.008 ;
  LAYER M2 ;
        RECT 6.4 2.04 6.432 2.072 ;
  LAYER M2 ;
        RECT 8.768 2.104 8.8 2.136 ;
  LAYER M2 ;
        RECT 6.4 2.168 6.432 2.2 ;
  LAYER M2 ;
        RECT 8.768 2.232 8.8 2.264 ;
  LAYER M2 ;
        RECT 6.4 2.296 6.432 2.328 ;
  LAYER M2 ;
        RECT 8.768 2.36 8.8 2.392 ;
  LAYER M2 ;
        RECT 6.4 2.424 6.432 2.456 ;
  LAYER M2 ;
        RECT 8.768 2.488 8.8 2.52 ;
  LAYER M2 ;
        RECT 6.4 2.552 6.432 2.584 ;
  LAYER M2 ;
        RECT 8.768 2.616 8.8 2.648 ;
  LAYER M2 ;
        RECT 6.4 2.68 6.432 2.712 ;
  LAYER M2 ;
        RECT 8.768 2.744 8.8 2.776 ;
  LAYER M2 ;
        RECT 6.4 2.808 6.432 2.84 ;
  LAYER M2 ;
        RECT 8.768 2.872 8.8 2.904 ;
  LAYER M2 ;
        RECT 6.4 2.936 6.432 2.968 ;
  LAYER M2 ;
        RECT 8.768 3 8.8 3.032 ;
  LAYER M2 ;
        RECT 6.4 3.064 6.432 3.096 ;
  LAYER M2 ;
        RECT 8.768 3.128 8.8 3.16 ;
  LAYER M2 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M1 ;
        RECT 6.4 3.912 6.432 6.42 ;
  LAYER M3 ;
        RECT 6.4 6.368 6.432 6.4 ;
  LAYER M1 ;
        RECT 6.464 3.912 6.496 6.42 ;
  LAYER M3 ;
        RECT 6.464 3.932 6.496 3.964 ;
  LAYER M1 ;
        RECT 6.528 3.912 6.56 6.42 ;
  LAYER M3 ;
        RECT 6.528 6.368 6.56 6.4 ;
  LAYER M1 ;
        RECT 6.592 3.912 6.624 6.42 ;
  LAYER M3 ;
        RECT 6.592 3.932 6.624 3.964 ;
  LAYER M1 ;
        RECT 6.656 3.912 6.688 6.42 ;
  LAYER M3 ;
        RECT 6.656 6.368 6.688 6.4 ;
  LAYER M1 ;
        RECT 6.72 3.912 6.752 6.42 ;
  LAYER M3 ;
        RECT 6.72 3.932 6.752 3.964 ;
  LAYER M1 ;
        RECT 6.784 3.912 6.816 6.42 ;
  LAYER M3 ;
        RECT 6.784 6.368 6.816 6.4 ;
  LAYER M1 ;
        RECT 6.848 3.912 6.88 6.42 ;
  LAYER M3 ;
        RECT 6.848 3.932 6.88 3.964 ;
  LAYER M1 ;
        RECT 6.912 3.912 6.944 6.42 ;
  LAYER M3 ;
        RECT 6.912 6.368 6.944 6.4 ;
  LAYER M1 ;
        RECT 6.976 3.912 7.008 6.42 ;
  LAYER M3 ;
        RECT 6.976 3.932 7.008 3.964 ;
  LAYER M1 ;
        RECT 7.04 3.912 7.072 6.42 ;
  LAYER M3 ;
        RECT 7.04 6.368 7.072 6.4 ;
  LAYER M1 ;
        RECT 7.104 3.912 7.136 6.42 ;
  LAYER M3 ;
        RECT 7.104 3.932 7.136 3.964 ;
  LAYER M1 ;
        RECT 7.168 3.912 7.2 6.42 ;
  LAYER M3 ;
        RECT 7.168 6.368 7.2 6.4 ;
  LAYER M1 ;
        RECT 7.232 3.912 7.264 6.42 ;
  LAYER M3 ;
        RECT 7.232 3.932 7.264 3.964 ;
  LAYER M1 ;
        RECT 7.296 3.912 7.328 6.42 ;
  LAYER M3 ;
        RECT 7.296 6.368 7.328 6.4 ;
  LAYER M1 ;
        RECT 7.36 3.912 7.392 6.42 ;
  LAYER M3 ;
        RECT 7.36 3.932 7.392 3.964 ;
  LAYER M1 ;
        RECT 7.424 3.912 7.456 6.42 ;
  LAYER M3 ;
        RECT 7.424 6.368 7.456 6.4 ;
  LAYER M1 ;
        RECT 7.488 3.912 7.52 6.42 ;
  LAYER M3 ;
        RECT 7.488 3.932 7.52 3.964 ;
  LAYER M1 ;
        RECT 7.552 3.912 7.584 6.42 ;
  LAYER M3 ;
        RECT 7.552 6.368 7.584 6.4 ;
  LAYER M1 ;
        RECT 7.616 3.912 7.648 6.42 ;
  LAYER M3 ;
        RECT 7.616 3.932 7.648 3.964 ;
  LAYER M1 ;
        RECT 7.68 3.912 7.712 6.42 ;
  LAYER M3 ;
        RECT 7.68 6.368 7.712 6.4 ;
  LAYER M1 ;
        RECT 7.744 3.912 7.776 6.42 ;
  LAYER M3 ;
        RECT 7.744 3.932 7.776 3.964 ;
  LAYER M1 ;
        RECT 7.808 3.912 7.84 6.42 ;
  LAYER M3 ;
        RECT 7.808 6.368 7.84 6.4 ;
  LAYER M1 ;
        RECT 7.872 3.912 7.904 6.42 ;
  LAYER M3 ;
        RECT 7.872 3.932 7.904 3.964 ;
  LAYER M1 ;
        RECT 7.936 3.912 7.968 6.42 ;
  LAYER M3 ;
        RECT 7.936 6.368 7.968 6.4 ;
  LAYER M1 ;
        RECT 8 3.912 8.032 6.42 ;
  LAYER M3 ;
        RECT 8 3.932 8.032 3.964 ;
  LAYER M1 ;
        RECT 8.064 3.912 8.096 6.42 ;
  LAYER M3 ;
        RECT 8.064 6.368 8.096 6.4 ;
  LAYER M1 ;
        RECT 8.128 3.912 8.16 6.42 ;
  LAYER M3 ;
        RECT 8.128 3.932 8.16 3.964 ;
  LAYER M1 ;
        RECT 8.192 3.912 8.224 6.42 ;
  LAYER M3 ;
        RECT 8.192 6.368 8.224 6.4 ;
  LAYER M1 ;
        RECT 8.256 3.912 8.288 6.42 ;
  LAYER M3 ;
        RECT 8.256 3.932 8.288 3.964 ;
  LAYER M1 ;
        RECT 8.32 3.912 8.352 6.42 ;
  LAYER M3 ;
        RECT 8.32 6.368 8.352 6.4 ;
  LAYER M1 ;
        RECT 8.384 3.912 8.416 6.42 ;
  LAYER M3 ;
        RECT 8.384 3.932 8.416 3.964 ;
  LAYER M1 ;
        RECT 8.448 3.912 8.48 6.42 ;
  LAYER M3 ;
        RECT 8.448 6.368 8.48 6.4 ;
  LAYER M1 ;
        RECT 8.512 3.912 8.544 6.42 ;
  LAYER M3 ;
        RECT 8.512 3.932 8.544 3.964 ;
  LAYER M1 ;
        RECT 8.576 3.912 8.608 6.42 ;
  LAYER M3 ;
        RECT 8.576 6.368 8.608 6.4 ;
  LAYER M1 ;
        RECT 8.64 3.912 8.672 6.42 ;
  LAYER M3 ;
        RECT 8.64 3.932 8.672 3.964 ;
  LAYER M1 ;
        RECT 8.704 3.912 8.736 6.42 ;
  LAYER M3 ;
        RECT 8.704 6.368 8.736 6.4 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 6.42 ;
  LAYER M3 ;
        RECT 6.4 3.996 6.432 4.028 ;
  LAYER M2 ;
        RECT 8.768 4.06 8.8 4.092 ;
  LAYER M2 ;
        RECT 6.4 4.124 6.432 4.156 ;
  LAYER M2 ;
        RECT 8.768 4.188 8.8 4.22 ;
  LAYER M2 ;
        RECT 6.4 4.252 6.432 4.284 ;
  LAYER M2 ;
        RECT 8.768 4.316 8.8 4.348 ;
  LAYER M2 ;
        RECT 6.4 4.38 6.432 4.412 ;
  LAYER M2 ;
        RECT 8.768 4.444 8.8 4.476 ;
  LAYER M2 ;
        RECT 6.4 4.508 6.432 4.54 ;
  LAYER M2 ;
        RECT 8.768 4.572 8.8 4.604 ;
  LAYER M2 ;
        RECT 6.4 4.636 6.432 4.668 ;
  LAYER M2 ;
        RECT 8.768 4.7 8.8 4.732 ;
  LAYER M2 ;
        RECT 6.4 4.764 6.432 4.796 ;
  LAYER M2 ;
        RECT 8.768 4.828 8.8 4.86 ;
  LAYER M2 ;
        RECT 6.4 4.892 6.432 4.924 ;
  LAYER M2 ;
        RECT 8.768 4.956 8.8 4.988 ;
  LAYER M2 ;
        RECT 6.4 5.02 6.432 5.052 ;
  LAYER M2 ;
        RECT 8.768 5.084 8.8 5.116 ;
  LAYER M2 ;
        RECT 6.4 5.148 6.432 5.18 ;
  LAYER M2 ;
        RECT 8.768 5.212 8.8 5.244 ;
  LAYER M2 ;
        RECT 6.4 5.276 6.432 5.308 ;
  LAYER M2 ;
        RECT 8.768 5.34 8.8 5.372 ;
  LAYER M2 ;
        RECT 6.4 5.404 6.432 5.436 ;
  LAYER M2 ;
        RECT 8.768 5.468 8.8 5.5 ;
  LAYER M2 ;
        RECT 6.4 5.532 6.432 5.564 ;
  LAYER M2 ;
        RECT 8.768 5.596 8.8 5.628 ;
  LAYER M2 ;
        RECT 6.4 5.66 6.432 5.692 ;
  LAYER M2 ;
        RECT 8.768 5.724 8.8 5.756 ;
  LAYER M2 ;
        RECT 6.4 5.788 6.432 5.82 ;
  LAYER M2 ;
        RECT 8.768 5.852 8.8 5.884 ;
  LAYER M2 ;
        RECT 6.4 5.916 6.432 5.948 ;
  LAYER M2 ;
        RECT 8.768 5.98 8.8 6.012 ;
  LAYER M2 ;
        RECT 6.4 6.044 6.432 6.076 ;
  LAYER M2 ;
        RECT 8.768 6.108 8.8 6.14 ;
  LAYER M2 ;
        RECT 6.4 6.172 6.432 6.204 ;
  LAYER M2 ;
        RECT 8.768 6.236 8.8 6.268 ;
  LAYER M2 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M1 ;
        RECT 6.4 7.02 6.432 9.528 ;
  LAYER M3 ;
        RECT 6.4 9.476 6.432 9.508 ;
  LAYER M1 ;
        RECT 6.464 7.02 6.496 9.528 ;
  LAYER M3 ;
        RECT 6.464 7.04 6.496 7.072 ;
  LAYER M1 ;
        RECT 6.528 7.02 6.56 9.528 ;
  LAYER M3 ;
        RECT 6.528 9.476 6.56 9.508 ;
  LAYER M1 ;
        RECT 6.592 7.02 6.624 9.528 ;
  LAYER M3 ;
        RECT 6.592 7.04 6.624 7.072 ;
  LAYER M1 ;
        RECT 6.656 7.02 6.688 9.528 ;
  LAYER M3 ;
        RECT 6.656 9.476 6.688 9.508 ;
  LAYER M1 ;
        RECT 6.72 7.02 6.752 9.528 ;
  LAYER M3 ;
        RECT 6.72 7.04 6.752 7.072 ;
  LAYER M1 ;
        RECT 6.784 7.02 6.816 9.528 ;
  LAYER M3 ;
        RECT 6.784 9.476 6.816 9.508 ;
  LAYER M1 ;
        RECT 6.848 7.02 6.88 9.528 ;
  LAYER M3 ;
        RECT 6.848 7.04 6.88 7.072 ;
  LAYER M1 ;
        RECT 6.912 7.02 6.944 9.528 ;
  LAYER M3 ;
        RECT 6.912 9.476 6.944 9.508 ;
  LAYER M1 ;
        RECT 6.976 7.02 7.008 9.528 ;
  LAYER M3 ;
        RECT 6.976 7.04 7.008 7.072 ;
  LAYER M1 ;
        RECT 7.04 7.02 7.072 9.528 ;
  LAYER M3 ;
        RECT 7.04 9.476 7.072 9.508 ;
  LAYER M1 ;
        RECT 7.104 7.02 7.136 9.528 ;
  LAYER M3 ;
        RECT 7.104 7.04 7.136 7.072 ;
  LAYER M1 ;
        RECT 7.168 7.02 7.2 9.528 ;
  LAYER M3 ;
        RECT 7.168 9.476 7.2 9.508 ;
  LAYER M1 ;
        RECT 7.232 7.02 7.264 9.528 ;
  LAYER M3 ;
        RECT 7.232 7.04 7.264 7.072 ;
  LAYER M1 ;
        RECT 7.296 7.02 7.328 9.528 ;
  LAYER M3 ;
        RECT 7.296 9.476 7.328 9.508 ;
  LAYER M1 ;
        RECT 7.36 7.02 7.392 9.528 ;
  LAYER M3 ;
        RECT 7.36 7.04 7.392 7.072 ;
  LAYER M1 ;
        RECT 7.424 7.02 7.456 9.528 ;
  LAYER M3 ;
        RECT 7.424 9.476 7.456 9.508 ;
  LAYER M1 ;
        RECT 7.488 7.02 7.52 9.528 ;
  LAYER M3 ;
        RECT 7.488 7.04 7.52 7.072 ;
  LAYER M1 ;
        RECT 7.552 7.02 7.584 9.528 ;
  LAYER M3 ;
        RECT 7.552 9.476 7.584 9.508 ;
  LAYER M1 ;
        RECT 7.616 7.02 7.648 9.528 ;
  LAYER M3 ;
        RECT 7.616 7.04 7.648 7.072 ;
  LAYER M1 ;
        RECT 7.68 7.02 7.712 9.528 ;
  LAYER M3 ;
        RECT 7.68 9.476 7.712 9.508 ;
  LAYER M1 ;
        RECT 7.744 7.02 7.776 9.528 ;
  LAYER M3 ;
        RECT 7.744 7.04 7.776 7.072 ;
  LAYER M1 ;
        RECT 7.808 7.02 7.84 9.528 ;
  LAYER M3 ;
        RECT 7.808 9.476 7.84 9.508 ;
  LAYER M1 ;
        RECT 7.872 7.02 7.904 9.528 ;
  LAYER M3 ;
        RECT 7.872 7.04 7.904 7.072 ;
  LAYER M1 ;
        RECT 7.936 7.02 7.968 9.528 ;
  LAYER M3 ;
        RECT 7.936 9.476 7.968 9.508 ;
  LAYER M1 ;
        RECT 8 7.02 8.032 9.528 ;
  LAYER M3 ;
        RECT 8 7.04 8.032 7.072 ;
  LAYER M1 ;
        RECT 8.064 7.02 8.096 9.528 ;
  LAYER M3 ;
        RECT 8.064 9.476 8.096 9.508 ;
  LAYER M1 ;
        RECT 8.128 7.02 8.16 9.528 ;
  LAYER M3 ;
        RECT 8.128 7.04 8.16 7.072 ;
  LAYER M1 ;
        RECT 8.192 7.02 8.224 9.528 ;
  LAYER M3 ;
        RECT 8.192 9.476 8.224 9.508 ;
  LAYER M1 ;
        RECT 8.256 7.02 8.288 9.528 ;
  LAYER M3 ;
        RECT 8.256 7.04 8.288 7.072 ;
  LAYER M1 ;
        RECT 8.32 7.02 8.352 9.528 ;
  LAYER M3 ;
        RECT 8.32 9.476 8.352 9.508 ;
  LAYER M1 ;
        RECT 8.384 7.02 8.416 9.528 ;
  LAYER M3 ;
        RECT 8.384 7.04 8.416 7.072 ;
  LAYER M1 ;
        RECT 8.448 7.02 8.48 9.528 ;
  LAYER M3 ;
        RECT 8.448 9.476 8.48 9.508 ;
  LAYER M1 ;
        RECT 8.512 7.02 8.544 9.528 ;
  LAYER M3 ;
        RECT 8.512 7.04 8.544 7.072 ;
  LAYER M1 ;
        RECT 8.576 7.02 8.608 9.528 ;
  LAYER M3 ;
        RECT 8.576 9.476 8.608 9.508 ;
  LAYER M1 ;
        RECT 8.64 7.02 8.672 9.528 ;
  LAYER M3 ;
        RECT 8.64 7.04 8.672 7.072 ;
  LAYER M1 ;
        RECT 8.704 7.02 8.736 9.528 ;
  LAYER M3 ;
        RECT 8.704 9.476 8.736 9.508 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 9.528 ;
  LAYER M3 ;
        RECT 6.4 7.104 6.432 7.136 ;
  LAYER M2 ;
        RECT 8.768 7.168 8.8 7.2 ;
  LAYER M2 ;
        RECT 6.4 7.232 6.432 7.264 ;
  LAYER M2 ;
        RECT 8.768 7.296 8.8 7.328 ;
  LAYER M2 ;
        RECT 6.4 7.36 6.432 7.392 ;
  LAYER M2 ;
        RECT 8.768 7.424 8.8 7.456 ;
  LAYER M2 ;
        RECT 6.4 7.488 6.432 7.52 ;
  LAYER M2 ;
        RECT 8.768 7.552 8.8 7.584 ;
  LAYER M2 ;
        RECT 6.4 7.616 6.432 7.648 ;
  LAYER M2 ;
        RECT 8.768 7.68 8.8 7.712 ;
  LAYER M2 ;
        RECT 6.4 7.744 6.432 7.776 ;
  LAYER M2 ;
        RECT 8.768 7.808 8.8 7.84 ;
  LAYER M2 ;
        RECT 6.4 7.872 6.432 7.904 ;
  LAYER M2 ;
        RECT 8.768 7.936 8.8 7.968 ;
  LAYER M2 ;
        RECT 6.4 8 6.432 8.032 ;
  LAYER M2 ;
        RECT 8.768 8.064 8.8 8.096 ;
  LAYER M2 ;
        RECT 6.4 8.128 6.432 8.16 ;
  LAYER M2 ;
        RECT 8.768 8.192 8.8 8.224 ;
  LAYER M2 ;
        RECT 6.4 8.256 6.432 8.288 ;
  LAYER M2 ;
        RECT 8.768 8.32 8.8 8.352 ;
  LAYER M2 ;
        RECT 6.4 8.384 6.432 8.416 ;
  LAYER M2 ;
        RECT 8.768 8.448 8.8 8.48 ;
  LAYER M2 ;
        RECT 6.4 8.512 6.432 8.544 ;
  LAYER M2 ;
        RECT 8.768 8.576 8.8 8.608 ;
  LAYER M2 ;
        RECT 6.4 8.64 6.432 8.672 ;
  LAYER M2 ;
        RECT 8.768 8.704 8.8 8.736 ;
  LAYER M2 ;
        RECT 6.4 8.768 6.432 8.8 ;
  LAYER M2 ;
        RECT 8.768 8.832 8.8 8.864 ;
  LAYER M2 ;
        RECT 6.4 8.896 6.432 8.928 ;
  LAYER M2 ;
        RECT 8.768 8.96 8.8 8.992 ;
  LAYER M2 ;
        RECT 6.4 9.024 6.432 9.056 ;
  LAYER M2 ;
        RECT 8.768 9.088 8.8 9.12 ;
  LAYER M2 ;
        RECT 6.4 9.152 6.432 9.184 ;
  LAYER M2 ;
        RECT 8.768 9.216 8.8 9.248 ;
  LAYER M2 ;
        RECT 6.4 9.28 6.432 9.312 ;
  LAYER M2 ;
        RECT 8.768 9.344 8.8 9.376 ;
  LAYER M2 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M1 ;
        RECT 6.4 10.128 6.432 12.636 ;
  LAYER M3 ;
        RECT 6.4 12.584 6.432 12.616 ;
  LAYER M1 ;
        RECT 6.464 10.128 6.496 12.636 ;
  LAYER M3 ;
        RECT 6.464 10.148 6.496 10.18 ;
  LAYER M1 ;
        RECT 6.528 10.128 6.56 12.636 ;
  LAYER M3 ;
        RECT 6.528 12.584 6.56 12.616 ;
  LAYER M1 ;
        RECT 6.592 10.128 6.624 12.636 ;
  LAYER M3 ;
        RECT 6.592 10.148 6.624 10.18 ;
  LAYER M1 ;
        RECT 6.656 10.128 6.688 12.636 ;
  LAYER M3 ;
        RECT 6.656 12.584 6.688 12.616 ;
  LAYER M1 ;
        RECT 6.72 10.128 6.752 12.636 ;
  LAYER M3 ;
        RECT 6.72 10.148 6.752 10.18 ;
  LAYER M1 ;
        RECT 6.784 10.128 6.816 12.636 ;
  LAYER M3 ;
        RECT 6.784 12.584 6.816 12.616 ;
  LAYER M1 ;
        RECT 6.848 10.128 6.88 12.636 ;
  LAYER M3 ;
        RECT 6.848 10.148 6.88 10.18 ;
  LAYER M1 ;
        RECT 6.912 10.128 6.944 12.636 ;
  LAYER M3 ;
        RECT 6.912 12.584 6.944 12.616 ;
  LAYER M1 ;
        RECT 6.976 10.128 7.008 12.636 ;
  LAYER M3 ;
        RECT 6.976 10.148 7.008 10.18 ;
  LAYER M1 ;
        RECT 7.04 10.128 7.072 12.636 ;
  LAYER M3 ;
        RECT 7.04 12.584 7.072 12.616 ;
  LAYER M1 ;
        RECT 7.104 10.128 7.136 12.636 ;
  LAYER M3 ;
        RECT 7.104 10.148 7.136 10.18 ;
  LAYER M1 ;
        RECT 7.168 10.128 7.2 12.636 ;
  LAYER M3 ;
        RECT 7.168 12.584 7.2 12.616 ;
  LAYER M1 ;
        RECT 7.232 10.128 7.264 12.636 ;
  LAYER M3 ;
        RECT 7.232 10.148 7.264 10.18 ;
  LAYER M1 ;
        RECT 7.296 10.128 7.328 12.636 ;
  LAYER M3 ;
        RECT 7.296 12.584 7.328 12.616 ;
  LAYER M1 ;
        RECT 7.36 10.128 7.392 12.636 ;
  LAYER M3 ;
        RECT 7.36 10.148 7.392 10.18 ;
  LAYER M1 ;
        RECT 7.424 10.128 7.456 12.636 ;
  LAYER M3 ;
        RECT 7.424 12.584 7.456 12.616 ;
  LAYER M1 ;
        RECT 7.488 10.128 7.52 12.636 ;
  LAYER M3 ;
        RECT 7.488 10.148 7.52 10.18 ;
  LAYER M1 ;
        RECT 7.552 10.128 7.584 12.636 ;
  LAYER M3 ;
        RECT 7.552 12.584 7.584 12.616 ;
  LAYER M1 ;
        RECT 7.616 10.128 7.648 12.636 ;
  LAYER M3 ;
        RECT 7.616 10.148 7.648 10.18 ;
  LAYER M1 ;
        RECT 7.68 10.128 7.712 12.636 ;
  LAYER M3 ;
        RECT 7.68 12.584 7.712 12.616 ;
  LAYER M1 ;
        RECT 7.744 10.128 7.776 12.636 ;
  LAYER M3 ;
        RECT 7.744 10.148 7.776 10.18 ;
  LAYER M1 ;
        RECT 7.808 10.128 7.84 12.636 ;
  LAYER M3 ;
        RECT 7.808 12.584 7.84 12.616 ;
  LAYER M1 ;
        RECT 7.872 10.128 7.904 12.636 ;
  LAYER M3 ;
        RECT 7.872 10.148 7.904 10.18 ;
  LAYER M1 ;
        RECT 7.936 10.128 7.968 12.636 ;
  LAYER M3 ;
        RECT 7.936 12.584 7.968 12.616 ;
  LAYER M1 ;
        RECT 8 10.128 8.032 12.636 ;
  LAYER M3 ;
        RECT 8 10.148 8.032 10.18 ;
  LAYER M1 ;
        RECT 8.064 10.128 8.096 12.636 ;
  LAYER M3 ;
        RECT 8.064 12.584 8.096 12.616 ;
  LAYER M1 ;
        RECT 8.128 10.128 8.16 12.636 ;
  LAYER M3 ;
        RECT 8.128 10.148 8.16 10.18 ;
  LAYER M1 ;
        RECT 8.192 10.128 8.224 12.636 ;
  LAYER M3 ;
        RECT 8.192 12.584 8.224 12.616 ;
  LAYER M1 ;
        RECT 8.256 10.128 8.288 12.636 ;
  LAYER M3 ;
        RECT 8.256 10.148 8.288 10.18 ;
  LAYER M1 ;
        RECT 8.32 10.128 8.352 12.636 ;
  LAYER M3 ;
        RECT 8.32 12.584 8.352 12.616 ;
  LAYER M1 ;
        RECT 8.384 10.128 8.416 12.636 ;
  LAYER M3 ;
        RECT 8.384 10.148 8.416 10.18 ;
  LAYER M1 ;
        RECT 8.448 10.128 8.48 12.636 ;
  LAYER M3 ;
        RECT 8.448 12.584 8.48 12.616 ;
  LAYER M1 ;
        RECT 8.512 10.128 8.544 12.636 ;
  LAYER M3 ;
        RECT 8.512 10.148 8.544 10.18 ;
  LAYER M1 ;
        RECT 8.576 10.128 8.608 12.636 ;
  LAYER M3 ;
        RECT 8.576 12.584 8.608 12.616 ;
  LAYER M1 ;
        RECT 8.64 10.128 8.672 12.636 ;
  LAYER M3 ;
        RECT 8.64 10.148 8.672 10.18 ;
  LAYER M1 ;
        RECT 8.704 10.128 8.736 12.636 ;
  LAYER M3 ;
        RECT 8.704 12.584 8.736 12.616 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 12.636 ;
  LAYER M3 ;
        RECT 6.4 10.212 6.432 10.244 ;
  LAYER M2 ;
        RECT 8.768 10.276 8.8 10.308 ;
  LAYER M2 ;
        RECT 6.4 10.34 6.432 10.372 ;
  LAYER M2 ;
        RECT 8.768 10.404 8.8 10.436 ;
  LAYER M2 ;
        RECT 6.4 10.468 6.432 10.5 ;
  LAYER M2 ;
        RECT 8.768 10.532 8.8 10.564 ;
  LAYER M2 ;
        RECT 6.4 10.596 6.432 10.628 ;
  LAYER M2 ;
        RECT 8.768 10.66 8.8 10.692 ;
  LAYER M2 ;
        RECT 6.4 10.724 6.432 10.756 ;
  LAYER M2 ;
        RECT 8.768 10.788 8.8 10.82 ;
  LAYER M2 ;
        RECT 6.4 10.852 6.432 10.884 ;
  LAYER M2 ;
        RECT 8.768 10.916 8.8 10.948 ;
  LAYER M2 ;
        RECT 6.4 10.98 6.432 11.012 ;
  LAYER M2 ;
        RECT 8.768 11.044 8.8 11.076 ;
  LAYER M2 ;
        RECT 6.4 11.108 6.432 11.14 ;
  LAYER M2 ;
        RECT 8.768 11.172 8.8 11.204 ;
  LAYER M2 ;
        RECT 6.4 11.236 6.432 11.268 ;
  LAYER M2 ;
        RECT 8.768 11.3 8.8 11.332 ;
  LAYER M2 ;
        RECT 6.4 11.364 6.432 11.396 ;
  LAYER M2 ;
        RECT 8.768 11.428 8.8 11.46 ;
  LAYER M2 ;
        RECT 6.4 11.492 6.432 11.524 ;
  LAYER M2 ;
        RECT 8.768 11.556 8.8 11.588 ;
  LAYER M2 ;
        RECT 6.4 11.62 6.432 11.652 ;
  LAYER M2 ;
        RECT 8.768 11.684 8.8 11.716 ;
  LAYER M2 ;
        RECT 6.4 11.748 6.432 11.78 ;
  LAYER M2 ;
        RECT 8.768 11.812 8.8 11.844 ;
  LAYER M2 ;
        RECT 6.4 11.876 6.432 11.908 ;
  LAYER M2 ;
        RECT 8.768 11.94 8.8 11.972 ;
  LAYER M2 ;
        RECT 6.4 12.004 6.432 12.036 ;
  LAYER M2 ;
        RECT 8.768 12.068 8.8 12.1 ;
  LAYER M2 ;
        RECT 6.4 12.132 6.432 12.164 ;
  LAYER M2 ;
        RECT 8.768 12.196 8.8 12.228 ;
  LAYER M2 ;
        RECT 6.4 12.26 6.432 12.292 ;
  LAYER M2 ;
        RECT 8.768 12.324 8.8 12.356 ;
  LAYER M2 ;
        RECT 6.4 12.388 6.432 12.42 ;
  LAYER M2 ;
        RECT 8.768 12.452 8.8 12.484 ;
  LAYER M2 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M1 ;
        RECT 6.4 13.236 6.432 15.744 ;
  LAYER M3 ;
        RECT 6.4 15.692 6.432 15.724 ;
  LAYER M1 ;
        RECT 6.464 13.236 6.496 15.744 ;
  LAYER M3 ;
        RECT 6.464 13.256 6.496 13.288 ;
  LAYER M1 ;
        RECT 6.528 13.236 6.56 15.744 ;
  LAYER M3 ;
        RECT 6.528 15.692 6.56 15.724 ;
  LAYER M1 ;
        RECT 6.592 13.236 6.624 15.744 ;
  LAYER M3 ;
        RECT 6.592 13.256 6.624 13.288 ;
  LAYER M1 ;
        RECT 6.656 13.236 6.688 15.744 ;
  LAYER M3 ;
        RECT 6.656 15.692 6.688 15.724 ;
  LAYER M1 ;
        RECT 6.72 13.236 6.752 15.744 ;
  LAYER M3 ;
        RECT 6.72 13.256 6.752 13.288 ;
  LAYER M1 ;
        RECT 6.784 13.236 6.816 15.744 ;
  LAYER M3 ;
        RECT 6.784 15.692 6.816 15.724 ;
  LAYER M1 ;
        RECT 6.848 13.236 6.88 15.744 ;
  LAYER M3 ;
        RECT 6.848 13.256 6.88 13.288 ;
  LAYER M1 ;
        RECT 6.912 13.236 6.944 15.744 ;
  LAYER M3 ;
        RECT 6.912 15.692 6.944 15.724 ;
  LAYER M1 ;
        RECT 6.976 13.236 7.008 15.744 ;
  LAYER M3 ;
        RECT 6.976 13.256 7.008 13.288 ;
  LAYER M1 ;
        RECT 7.04 13.236 7.072 15.744 ;
  LAYER M3 ;
        RECT 7.04 15.692 7.072 15.724 ;
  LAYER M1 ;
        RECT 7.104 13.236 7.136 15.744 ;
  LAYER M3 ;
        RECT 7.104 13.256 7.136 13.288 ;
  LAYER M1 ;
        RECT 7.168 13.236 7.2 15.744 ;
  LAYER M3 ;
        RECT 7.168 15.692 7.2 15.724 ;
  LAYER M1 ;
        RECT 7.232 13.236 7.264 15.744 ;
  LAYER M3 ;
        RECT 7.232 13.256 7.264 13.288 ;
  LAYER M1 ;
        RECT 7.296 13.236 7.328 15.744 ;
  LAYER M3 ;
        RECT 7.296 15.692 7.328 15.724 ;
  LAYER M1 ;
        RECT 7.36 13.236 7.392 15.744 ;
  LAYER M3 ;
        RECT 7.36 13.256 7.392 13.288 ;
  LAYER M1 ;
        RECT 7.424 13.236 7.456 15.744 ;
  LAYER M3 ;
        RECT 7.424 15.692 7.456 15.724 ;
  LAYER M1 ;
        RECT 7.488 13.236 7.52 15.744 ;
  LAYER M3 ;
        RECT 7.488 13.256 7.52 13.288 ;
  LAYER M1 ;
        RECT 7.552 13.236 7.584 15.744 ;
  LAYER M3 ;
        RECT 7.552 15.692 7.584 15.724 ;
  LAYER M1 ;
        RECT 7.616 13.236 7.648 15.744 ;
  LAYER M3 ;
        RECT 7.616 13.256 7.648 13.288 ;
  LAYER M1 ;
        RECT 7.68 13.236 7.712 15.744 ;
  LAYER M3 ;
        RECT 7.68 15.692 7.712 15.724 ;
  LAYER M1 ;
        RECT 7.744 13.236 7.776 15.744 ;
  LAYER M3 ;
        RECT 7.744 13.256 7.776 13.288 ;
  LAYER M1 ;
        RECT 7.808 13.236 7.84 15.744 ;
  LAYER M3 ;
        RECT 7.808 15.692 7.84 15.724 ;
  LAYER M1 ;
        RECT 7.872 13.236 7.904 15.744 ;
  LAYER M3 ;
        RECT 7.872 13.256 7.904 13.288 ;
  LAYER M1 ;
        RECT 7.936 13.236 7.968 15.744 ;
  LAYER M3 ;
        RECT 7.936 15.692 7.968 15.724 ;
  LAYER M1 ;
        RECT 8 13.236 8.032 15.744 ;
  LAYER M3 ;
        RECT 8 13.256 8.032 13.288 ;
  LAYER M1 ;
        RECT 8.064 13.236 8.096 15.744 ;
  LAYER M3 ;
        RECT 8.064 15.692 8.096 15.724 ;
  LAYER M1 ;
        RECT 8.128 13.236 8.16 15.744 ;
  LAYER M3 ;
        RECT 8.128 13.256 8.16 13.288 ;
  LAYER M1 ;
        RECT 8.192 13.236 8.224 15.744 ;
  LAYER M3 ;
        RECT 8.192 15.692 8.224 15.724 ;
  LAYER M1 ;
        RECT 8.256 13.236 8.288 15.744 ;
  LAYER M3 ;
        RECT 8.256 13.256 8.288 13.288 ;
  LAYER M1 ;
        RECT 8.32 13.236 8.352 15.744 ;
  LAYER M3 ;
        RECT 8.32 15.692 8.352 15.724 ;
  LAYER M1 ;
        RECT 8.384 13.236 8.416 15.744 ;
  LAYER M3 ;
        RECT 8.384 13.256 8.416 13.288 ;
  LAYER M1 ;
        RECT 8.448 13.236 8.48 15.744 ;
  LAYER M3 ;
        RECT 8.448 15.692 8.48 15.724 ;
  LAYER M1 ;
        RECT 8.512 13.236 8.544 15.744 ;
  LAYER M3 ;
        RECT 8.512 13.256 8.544 13.288 ;
  LAYER M1 ;
        RECT 8.576 13.236 8.608 15.744 ;
  LAYER M3 ;
        RECT 8.576 15.692 8.608 15.724 ;
  LAYER M1 ;
        RECT 8.64 13.236 8.672 15.744 ;
  LAYER M3 ;
        RECT 8.64 13.256 8.672 13.288 ;
  LAYER M1 ;
        RECT 8.704 13.236 8.736 15.744 ;
  LAYER M3 ;
        RECT 8.704 15.692 8.736 15.724 ;
  LAYER M1 ;
        RECT 8.768 13.236 8.8 15.744 ;
  LAYER M3 ;
        RECT 6.4 13.32 6.432 13.352 ;
  LAYER M2 ;
        RECT 8.768 13.384 8.8 13.416 ;
  LAYER M2 ;
        RECT 6.4 13.448 6.432 13.48 ;
  LAYER M2 ;
        RECT 8.768 13.512 8.8 13.544 ;
  LAYER M2 ;
        RECT 6.4 13.576 6.432 13.608 ;
  LAYER M2 ;
        RECT 8.768 13.64 8.8 13.672 ;
  LAYER M2 ;
        RECT 6.4 13.704 6.432 13.736 ;
  LAYER M2 ;
        RECT 8.768 13.768 8.8 13.8 ;
  LAYER M2 ;
        RECT 6.4 13.832 6.432 13.864 ;
  LAYER M2 ;
        RECT 8.768 13.896 8.8 13.928 ;
  LAYER M2 ;
        RECT 6.4 13.96 6.432 13.992 ;
  LAYER M2 ;
        RECT 8.768 14.024 8.8 14.056 ;
  LAYER M2 ;
        RECT 6.4 14.088 6.432 14.12 ;
  LAYER M2 ;
        RECT 8.768 14.152 8.8 14.184 ;
  LAYER M2 ;
        RECT 6.4 14.216 6.432 14.248 ;
  LAYER M2 ;
        RECT 8.768 14.28 8.8 14.312 ;
  LAYER M2 ;
        RECT 6.4 14.344 6.432 14.376 ;
  LAYER M2 ;
        RECT 8.768 14.408 8.8 14.44 ;
  LAYER M2 ;
        RECT 6.4 14.472 6.432 14.504 ;
  LAYER M2 ;
        RECT 8.768 14.536 8.8 14.568 ;
  LAYER M2 ;
        RECT 6.4 14.6 6.432 14.632 ;
  LAYER M2 ;
        RECT 8.768 14.664 8.8 14.696 ;
  LAYER M2 ;
        RECT 6.4 14.728 6.432 14.76 ;
  LAYER M2 ;
        RECT 8.768 14.792 8.8 14.824 ;
  LAYER M2 ;
        RECT 6.4 14.856 6.432 14.888 ;
  LAYER M2 ;
        RECT 8.768 14.92 8.8 14.952 ;
  LAYER M2 ;
        RECT 6.4 14.984 6.432 15.016 ;
  LAYER M2 ;
        RECT 8.768 15.048 8.8 15.08 ;
  LAYER M2 ;
        RECT 6.4 15.112 6.432 15.144 ;
  LAYER M2 ;
        RECT 8.768 15.176 8.8 15.208 ;
  LAYER M2 ;
        RECT 6.4 15.24 6.432 15.272 ;
  LAYER M2 ;
        RECT 8.768 15.304 8.8 15.336 ;
  LAYER M2 ;
        RECT 6.4 15.368 6.432 15.4 ;
  LAYER M2 ;
        RECT 8.768 15.432 8.8 15.464 ;
  LAYER M2 ;
        RECT 6.4 15.496 6.432 15.528 ;
  LAYER M2 ;
        RECT 8.768 15.56 8.8 15.592 ;
  LAYER M2 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M1 ;
        RECT 6.4 16.344 6.432 18.852 ;
  LAYER M3 ;
        RECT 6.4 18.8 6.432 18.832 ;
  LAYER M1 ;
        RECT 6.464 16.344 6.496 18.852 ;
  LAYER M3 ;
        RECT 6.464 16.364 6.496 16.396 ;
  LAYER M1 ;
        RECT 6.528 16.344 6.56 18.852 ;
  LAYER M3 ;
        RECT 6.528 18.8 6.56 18.832 ;
  LAYER M1 ;
        RECT 6.592 16.344 6.624 18.852 ;
  LAYER M3 ;
        RECT 6.592 16.364 6.624 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 18.852 ;
  LAYER M3 ;
        RECT 6.656 18.8 6.688 18.832 ;
  LAYER M1 ;
        RECT 6.72 16.344 6.752 18.852 ;
  LAYER M3 ;
        RECT 6.72 16.364 6.752 16.396 ;
  LAYER M1 ;
        RECT 6.784 16.344 6.816 18.852 ;
  LAYER M3 ;
        RECT 6.784 18.8 6.816 18.832 ;
  LAYER M1 ;
        RECT 6.848 16.344 6.88 18.852 ;
  LAYER M3 ;
        RECT 6.848 16.364 6.88 16.396 ;
  LAYER M1 ;
        RECT 6.912 16.344 6.944 18.852 ;
  LAYER M3 ;
        RECT 6.912 18.8 6.944 18.832 ;
  LAYER M1 ;
        RECT 6.976 16.344 7.008 18.852 ;
  LAYER M3 ;
        RECT 6.976 16.364 7.008 16.396 ;
  LAYER M1 ;
        RECT 7.04 16.344 7.072 18.852 ;
  LAYER M3 ;
        RECT 7.04 18.8 7.072 18.832 ;
  LAYER M1 ;
        RECT 7.104 16.344 7.136 18.852 ;
  LAYER M3 ;
        RECT 7.104 16.364 7.136 16.396 ;
  LAYER M1 ;
        RECT 7.168 16.344 7.2 18.852 ;
  LAYER M3 ;
        RECT 7.168 18.8 7.2 18.832 ;
  LAYER M1 ;
        RECT 7.232 16.344 7.264 18.852 ;
  LAYER M3 ;
        RECT 7.232 16.364 7.264 16.396 ;
  LAYER M1 ;
        RECT 7.296 16.344 7.328 18.852 ;
  LAYER M3 ;
        RECT 7.296 18.8 7.328 18.832 ;
  LAYER M1 ;
        RECT 7.36 16.344 7.392 18.852 ;
  LAYER M3 ;
        RECT 7.36 16.364 7.392 16.396 ;
  LAYER M1 ;
        RECT 7.424 16.344 7.456 18.852 ;
  LAYER M3 ;
        RECT 7.424 18.8 7.456 18.832 ;
  LAYER M1 ;
        RECT 7.488 16.344 7.52 18.852 ;
  LAYER M3 ;
        RECT 7.488 16.364 7.52 16.396 ;
  LAYER M1 ;
        RECT 7.552 16.344 7.584 18.852 ;
  LAYER M3 ;
        RECT 7.552 18.8 7.584 18.832 ;
  LAYER M1 ;
        RECT 7.616 16.344 7.648 18.852 ;
  LAYER M3 ;
        RECT 7.616 16.364 7.648 16.396 ;
  LAYER M1 ;
        RECT 7.68 16.344 7.712 18.852 ;
  LAYER M3 ;
        RECT 7.68 18.8 7.712 18.832 ;
  LAYER M1 ;
        RECT 7.744 16.344 7.776 18.852 ;
  LAYER M3 ;
        RECT 7.744 16.364 7.776 16.396 ;
  LAYER M1 ;
        RECT 7.808 16.344 7.84 18.852 ;
  LAYER M3 ;
        RECT 7.808 18.8 7.84 18.832 ;
  LAYER M1 ;
        RECT 7.872 16.344 7.904 18.852 ;
  LAYER M3 ;
        RECT 7.872 16.364 7.904 16.396 ;
  LAYER M1 ;
        RECT 7.936 16.344 7.968 18.852 ;
  LAYER M3 ;
        RECT 7.936 18.8 7.968 18.832 ;
  LAYER M1 ;
        RECT 8 16.344 8.032 18.852 ;
  LAYER M3 ;
        RECT 8 16.364 8.032 16.396 ;
  LAYER M1 ;
        RECT 8.064 16.344 8.096 18.852 ;
  LAYER M3 ;
        RECT 8.064 18.8 8.096 18.832 ;
  LAYER M1 ;
        RECT 8.128 16.344 8.16 18.852 ;
  LAYER M3 ;
        RECT 8.128 16.364 8.16 16.396 ;
  LAYER M1 ;
        RECT 8.192 16.344 8.224 18.852 ;
  LAYER M3 ;
        RECT 8.192 18.8 8.224 18.832 ;
  LAYER M1 ;
        RECT 8.256 16.344 8.288 18.852 ;
  LAYER M3 ;
        RECT 8.256 16.364 8.288 16.396 ;
  LAYER M1 ;
        RECT 8.32 16.344 8.352 18.852 ;
  LAYER M3 ;
        RECT 8.32 18.8 8.352 18.832 ;
  LAYER M1 ;
        RECT 8.384 16.344 8.416 18.852 ;
  LAYER M3 ;
        RECT 8.384 16.364 8.416 16.396 ;
  LAYER M1 ;
        RECT 8.448 16.344 8.48 18.852 ;
  LAYER M3 ;
        RECT 8.448 18.8 8.48 18.832 ;
  LAYER M1 ;
        RECT 8.512 16.344 8.544 18.852 ;
  LAYER M3 ;
        RECT 8.512 16.364 8.544 16.396 ;
  LAYER M1 ;
        RECT 8.576 16.344 8.608 18.852 ;
  LAYER M3 ;
        RECT 8.576 18.8 8.608 18.832 ;
  LAYER M1 ;
        RECT 8.64 16.344 8.672 18.852 ;
  LAYER M3 ;
        RECT 8.64 16.364 8.672 16.396 ;
  LAYER M1 ;
        RECT 8.704 16.344 8.736 18.852 ;
  LAYER M3 ;
        RECT 8.704 18.8 8.736 18.832 ;
  LAYER M1 ;
        RECT 8.768 16.344 8.8 18.852 ;
  LAYER M3 ;
        RECT 6.4 16.428 6.432 16.46 ;
  LAYER M2 ;
        RECT 8.768 16.492 8.8 16.524 ;
  LAYER M2 ;
        RECT 6.4 16.556 6.432 16.588 ;
  LAYER M2 ;
        RECT 8.768 16.62 8.8 16.652 ;
  LAYER M2 ;
        RECT 6.4 16.684 6.432 16.716 ;
  LAYER M2 ;
        RECT 8.768 16.748 8.8 16.78 ;
  LAYER M2 ;
        RECT 6.4 16.812 6.432 16.844 ;
  LAYER M2 ;
        RECT 8.768 16.876 8.8 16.908 ;
  LAYER M2 ;
        RECT 6.4 16.94 6.432 16.972 ;
  LAYER M2 ;
        RECT 8.768 17.004 8.8 17.036 ;
  LAYER M2 ;
        RECT 6.4 17.068 6.432 17.1 ;
  LAYER M2 ;
        RECT 8.768 17.132 8.8 17.164 ;
  LAYER M2 ;
        RECT 6.4 17.196 6.432 17.228 ;
  LAYER M2 ;
        RECT 8.768 17.26 8.8 17.292 ;
  LAYER M2 ;
        RECT 6.4 17.324 6.432 17.356 ;
  LAYER M2 ;
        RECT 8.768 17.388 8.8 17.42 ;
  LAYER M2 ;
        RECT 6.4 17.452 6.432 17.484 ;
  LAYER M2 ;
        RECT 8.768 17.516 8.8 17.548 ;
  LAYER M2 ;
        RECT 6.4 17.58 6.432 17.612 ;
  LAYER M2 ;
        RECT 8.768 17.644 8.8 17.676 ;
  LAYER M2 ;
        RECT 6.4 17.708 6.432 17.74 ;
  LAYER M2 ;
        RECT 8.768 17.772 8.8 17.804 ;
  LAYER M2 ;
        RECT 6.4 17.836 6.432 17.868 ;
  LAYER M2 ;
        RECT 8.768 17.9 8.8 17.932 ;
  LAYER M2 ;
        RECT 6.4 17.964 6.432 17.996 ;
  LAYER M2 ;
        RECT 8.768 18.028 8.8 18.06 ;
  LAYER M2 ;
        RECT 6.4 18.092 6.432 18.124 ;
  LAYER M2 ;
        RECT 8.768 18.156 8.8 18.188 ;
  LAYER M2 ;
        RECT 6.4 18.22 6.432 18.252 ;
  LAYER M2 ;
        RECT 8.768 18.284 8.8 18.316 ;
  LAYER M2 ;
        RECT 6.4 18.348 6.432 18.38 ;
  LAYER M2 ;
        RECT 8.768 18.412 8.8 18.444 ;
  LAYER M2 ;
        RECT 6.4 18.476 6.432 18.508 ;
  LAYER M2 ;
        RECT 8.768 18.54 8.8 18.572 ;
  LAYER M2 ;
        RECT 6.4 18.604 6.432 18.636 ;
  LAYER M2 ;
        RECT 8.768 18.668 8.8 18.7 ;
  LAYER M2 ;
        RECT 6.352 16.296 8.848 18.9 ;
  LAYER M1 ;
        RECT 6.4 19.452 6.432 21.96 ;
  LAYER M3 ;
        RECT 6.4 21.908 6.432 21.94 ;
  LAYER M1 ;
        RECT 6.464 19.452 6.496 21.96 ;
  LAYER M3 ;
        RECT 6.464 19.472 6.496 19.504 ;
  LAYER M1 ;
        RECT 6.528 19.452 6.56 21.96 ;
  LAYER M3 ;
        RECT 6.528 21.908 6.56 21.94 ;
  LAYER M1 ;
        RECT 6.592 19.452 6.624 21.96 ;
  LAYER M3 ;
        RECT 6.592 19.472 6.624 19.504 ;
  LAYER M1 ;
        RECT 6.656 19.452 6.688 21.96 ;
  LAYER M3 ;
        RECT 6.656 21.908 6.688 21.94 ;
  LAYER M1 ;
        RECT 6.72 19.452 6.752 21.96 ;
  LAYER M3 ;
        RECT 6.72 19.472 6.752 19.504 ;
  LAYER M1 ;
        RECT 6.784 19.452 6.816 21.96 ;
  LAYER M3 ;
        RECT 6.784 21.908 6.816 21.94 ;
  LAYER M1 ;
        RECT 6.848 19.452 6.88 21.96 ;
  LAYER M3 ;
        RECT 6.848 19.472 6.88 19.504 ;
  LAYER M1 ;
        RECT 6.912 19.452 6.944 21.96 ;
  LAYER M3 ;
        RECT 6.912 21.908 6.944 21.94 ;
  LAYER M1 ;
        RECT 6.976 19.452 7.008 21.96 ;
  LAYER M3 ;
        RECT 6.976 19.472 7.008 19.504 ;
  LAYER M1 ;
        RECT 7.04 19.452 7.072 21.96 ;
  LAYER M3 ;
        RECT 7.04 21.908 7.072 21.94 ;
  LAYER M1 ;
        RECT 7.104 19.452 7.136 21.96 ;
  LAYER M3 ;
        RECT 7.104 19.472 7.136 19.504 ;
  LAYER M1 ;
        RECT 7.168 19.452 7.2 21.96 ;
  LAYER M3 ;
        RECT 7.168 21.908 7.2 21.94 ;
  LAYER M1 ;
        RECT 7.232 19.452 7.264 21.96 ;
  LAYER M3 ;
        RECT 7.232 19.472 7.264 19.504 ;
  LAYER M1 ;
        RECT 7.296 19.452 7.328 21.96 ;
  LAYER M3 ;
        RECT 7.296 21.908 7.328 21.94 ;
  LAYER M1 ;
        RECT 7.36 19.452 7.392 21.96 ;
  LAYER M3 ;
        RECT 7.36 19.472 7.392 19.504 ;
  LAYER M1 ;
        RECT 7.424 19.452 7.456 21.96 ;
  LAYER M3 ;
        RECT 7.424 21.908 7.456 21.94 ;
  LAYER M1 ;
        RECT 7.488 19.452 7.52 21.96 ;
  LAYER M3 ;
        RECT 7.488 19.472 7.52 19.504 ;
  LAYER M1 ;
        RECT 7.552 19.452 7.584 21.96 ;
  LAYER M3 ;
        RECT 7.552 21.908 7.584 21.94 ;
  LAYER M1 ;
        RECT 7.616 19.452 7.648 21.96 ;
  LAYER M3 ;
        RECT 7.616 19.472 7.648 19.504 ;
  LAYER M1 ;
        RECT 7.68 19.452 7.712 21.96 ;
  LAYER M3 ;
        RECT 7.68 21.908 7.712 21.94 ;
  LAYER M1 ;
        RECT 7.744 19.452 7.776 21.96 ;
  LAYER M3 ;
        RECT 7.744 19.472 7.776 19.504 ;
  LAYER M1 ;
        RECT 7.808 19.452 7.84 21.96 ;
  LAYER M3 ;
        RECT 7.808 21.908 7.84 21.94 ;
  LAYER M1 ;
        RECT 7.872 19.452 7.904 21.96 ;
  LAYER M3 ;
        RECT 7.872 19.472 7.904 19.504 ;
  LAYER M1 ;
        RECT 7.936 19.452 7.968 21.96 ;
  LAYER M3 ;
        RECT 7.936 21.908 7.968 21.94 ;
  LAYER M1 ;
        RECT 8 19.452 8.032 21.96 ;
  LAYER M3 ;
        RECT 8 19.472 8.032 19.504 ;
  LAYER M1 ;
        RECT 8.064 19.452 8.096 21.96 ;
  LAYER M3 ;
        RECT 8.064 21.908 8.096 21.94 ;
  LAYER M1 ;
        RECT 8.128 19.452 8.16 21.96 ;
  LAYER M3 ;
        RECT 8.128 19.472 8.16 19.504 ;
  LAYER M1 ;
        RECT 8.192 19.452 8.224 21.96 ;
  LAYER M3 ;
        RECT 8.192 21.908 8.224 21.94 ;
  LAYER M1 ;
        RECT 8.256 19.452 8.288 21.96 ;
  LAYER M3 ;
        RECT 8.256 19.472 8.288 19.504 ;
  LAYER M1 ;
        RECT 8.32 19.452 8.352 21.96 ;
  LAYER M3 ;
        RECT 8.32 21.908 8.352 21.94 ;
  LAYER M1 ;
        RECT 8.384 19.452 8.416 21.96 ;
  LAYER M3 ;
        RECT 8.384 19.472 8.416 19.504 ;
  LAYER M1 ;
        RECT 8.448 19.452 8.48 21.96 ;
  LAYER M3 ;
        RECT 8.448 21.908 8.48 21.94 ;
  LAYER M1 ;
        RECT 8.512 19.452 8.544 21.96 ;
  LAYER M3 ;
        RECT 8.512 19.472 8.544 19.504 ;
  LAYER M1 ;
        RECT 8.576 19.452 8.608 21.96 ;
  LAYER M3 ;
        RECT 8.576 21.908 8.608 21.94 ;
  LAYER M1 ;
        RECT 8.64 19.452 8.672 21.96 ;
  LAYER M3 ;
        RECT 8.64 19.472 8.672 19.504 ;
  LAYER M1 ;
        RECT 8.704 19.452 8.736 21.96 ;
  LAYER M3 ;
        RECT 8.704 21.908 8.736 21.94 ;
  LAYER M1 ;
        RECT 8.768 19.452 8.8 21.96 ;
  LAYER M3 ;
        RECT 6.4 19.536 6.432 19.568 ;
  LAYER M2 ;
        RECT 8.768 19.6 8.8 19.632 ;
  LAYER M2 ;
        RECT 6.4 19.664 6.432 19.696 ;
  LAYER M2 ;
        RECT 8.768 19.728 8.8 19.76 ;
  LAYER M2 ;
        RECT 6.4 19.792 6.432 19.824 ;
  LAYER M2 ;
        RECT 8.768 19.856 8.8 19.888 ;
  LAYER M2 ;
        RECT 6.4 19.92 6.432 19.952 ;
  LAYER M2 ;
        RECT 8.768 19.984 8.8 20.016 ;
  LAYER M2 ;
        RECT 6.4 20.048 6.432 20.08 ;
  LAYER M2 ;
        RECT 8.768 20.112 8.8 20.144 ;
  LAYER M2 ;
        RECT 6.4 20.176 6.432 20.208 ;
  LAYER M2 ;
        RECT 8.768 20.24 8.8 20.272 ;
  LAYER M2 ;
        RECT 6.4 20.304 6.432 20.336 ;
  LAYER M2 ;
        RECT 8.768 20.368 8.8 20.4 ;
  LAYER M2 ;
        RECT 6.4 20.432 6.432 20.464 ;
  LAYER M2 ;
        RECT 8.768 20.496 8.8 20.528 ;
  LAYER M2 ;
        RECT 6.4 20.56 6.432 20.592 ;
  LAYER M2 ;
        RECT 8.768 20.624 8.8 20.656 ;
  LAYER M2 ;
        RECT 6.4 20.688 6.432 20.72 ;
  LAYER M2 ;
        RECT 8.768 20.752 8.8 20.784 ;
  LAYER M2 ;
        RECT 6.4 20.816 6.432 20.848 ;
  LAYER M2 ;
        RECT 8.768 20.88 8.8 20.912 ;
  LAYER M2 ;
        RECT 6.4 20.944 6.432 20.976 ;
  LAYER M2 ;
        RECT 8.768 21.008 8.8 21.04 ;
  LAYER M2 ;
        RECT 6.4 21.072 6.432 21.104 ;
  LAYER M2 ;
        RECT 8.768 21.136 8.8 21.168 ;
  LAYER M2 ;
        RECT 6.4 21.2 6.432 21.232 ;
  LAYER M2 ;
        RECT 8.768 21.264 8.8 21.296 ;
  LAYER M2 ;
        RECT 6.4 21.328 6.432 21.36 ;
  LAYER M2 ;
        RECT 8.768 21.392 8.8 21.424 ;
  LAYER M2 ;
        RECT 6.4 21.456 6.432 21.488 ;
  LAYER M2 ;
        RECT 8.768 21.52 8.8 21.552 ;
  LAYER M2 ;
        RECT 6.4 21.584 6.432 21.616 ;
  LAYER M2 ;
        RECT 8.768 21.648 8.8 21.68 ;
  LAYER M2 ;
        RECT 6.4 21.712 6.432 21.744 ;
  LAYER M2 ;
        RECT 8.768 21.776 8.8 21.808 ;
  LAYER M2 ;
        RECT 6.352 19.404 8.848 22.008 ;
  LAYER M1 ;
        RECT 6.4 22.56 6.432 25.068 ;
  LAYER M3 ;
        RECT 6.4 25.016 6.432 25.048 ;
  LAYER M1 ;
        RECT 6.464 22.56 6.496 25.068 ;
  LAYER M3 ;
        RECT 6.464 22.58 6.496 22.612 ;
  LAYER M1 ;
        RECT 6.528 22.56 6.56 25.068 ;
  LAYER M3 ;
        RECT 6.528 25.016 6.56 25.048 ;
  LAYER M1 ;
        RECT 6.592 22.56 6.624 25.068 ;
  LAYER M3 ;
        RECT 6.592 22.58 6.624 22.612 ;
  LAYER M1 ;
        RECT 6.656 22.56 6.688 25.068 ;
  LAYER M3 ;
        RECT 6.656 25.016 6.688 25.048 ;
  LAYER M1 ;
        RECT 6.72 22.56 6.752 25.068 ;
  LAYER M3 ;
        RECT 6.72 22.58 6.752 22.612 ;
  LAYER M1 ;
        RECT 6.784 22.56 6.816 25.068 ;
  LAYER M3 ;
        RECT 6.784 25.016 6.816 25.048 ;
  LAYER M1 ;
        RECT 6.848 22.56 6.88 25.068 ;
  LAYER M3 ;
        RECT 6.848 22.58 6.88 22.612 ;
  LAYER M1 ;
        RECT 6.912 22.56 6.944 25.068 ;
  LAYER M3 ;
        RECT 6.912 25.016 6.944 25.048 ;
  LAYER M1 ;
        RECT 6.976 22.56 7.008 25.068 ;
  LAYER M3 ;
        RECT 6.976 22.58 7.008 22.612 ;
  LAYER M1 ;
        RECT 7.04 22.56 7.072 25.068 ;
  LAYER M3 ;
        RECT 7.04 25.016 7.072 25.048 ;
  LAYER M1 ;
        RECT 7.104 22.56 7.136 25.068 ;
  LAYER M3 ;
        RECT 7.104 22.58 7.136 22.612 ;
  LAYER M1 ;
        RECT 7.168 22.56 7.2 25.068 ;
  LAYER M3 ;
        RECT 7.168 25.016 7.2 25.048 ;
  LAYER M1 ;
        RECT 7.232 22.56 7.264 25.068 ;
  LAYER M3 ;
        RECT 7.232 22.58 7.264 22.612 ;
  LAYER M1 ;
        RECT 7.296 22.56 7.328 25.068 ;
  LAYER M3 ;
        RECT 7.296 25.016 7.328 25.048 ;
  LAYER M1 ;
        RECT 7.36 22.56 7.392 25.068 ;
  LAYER M3 ;
        RECT 7.36 22.58 7.392 22.612 ;
  LAYER M1 ;
        RECT 7.424 22.56 7.456 25.068 ;
  LAYER M3 ;
        RECT 7.424 25.016 7.456 25.048 ;
  LAYER M1 ;
        RECT 7.488 22.56 7.52 25.068 ;
  LAYER M3 ;
        RECT 7.488 22.58 7.52 22.612 ;
  LAYER M1 ;
        RECT 7.552 22.56 7.584 25.068 ;
  LAYER M3 ;
        RECT 7.552 25.016 7.584 25.048 ;
  LAYER M1 ;
        RECT 7.616 22.56 7.648 25.068 ;
  LAYER M3 ;
        RECT 7.616 22.58 7.648 22.612 ;
  LAYER M1 ;
        RECT 7.68 22.56 7.712 25.068 ;
  LAYER M3 ;
        RECT 7.68 25.016 7.712 25.048 ;
  LAYER M1 ;
        RECT 7.744 22.56 7.776 25.068 ;
  LAYER M3 ;
        RECT 7.744 22.58 7.776 22.612 ;
  LAYER M1 ;
        RECT 7.808 22.56 7.84 25.068 ;
  LAYER M3 ;
        RECT 7.808 25.016 7.84 25.048 ;
  LAYER M1 ;
        RECT 7.872 22.56 7.904 25.068 ;
  LAYER M3 ;
        RECT 7.872 22.58 7.904 22.612 ;
  LAYER M1 ;
        RECT 7.936 22.56 7.968 25.068 ;
  LAYER M3 ;
        RECT 7.936 25.016 7.968 25.048 ;
  LAYER M1 ;
        RECT 8 22.56 8.032 25.068 ;
  LAYER M3 ;
        RECT 8 22.58 8.032 22.612 ;
  LAYER M1 ;
        RECT 8.064 22.56 8.096 25.068 ;
  LAYER M3 ;
        RECT 8.064 25.016 8.096 25.048 ;
  LAYER M1 ;
        RECT 8.128 22.56 8.16 25.068 ;
  LAYER M3 ;
        RECT 8.128 22.58 8.16 22.612 ;
  LAYER M1 ;
        RECT 8.192 22.56 8.224 25.068 ;
  LAYER M3 ;
        RECT 8.192 25.016 8.224 25.048 ;
  LAYER M1 ;
        RECT 8.256 22.56 8.288 25.068 ;
  LAYER M3 ;
        RECT 8.256 22.58 8.288 22.612 ;
  LAYER M1 ;
        RECT 8.32 22.56 8.352 25.068 ;
  LAYER M3 ;
        RECT 8.32 25.016 8.352 25.048 ;
  LAYER M1 ;
        RECT 8.384 22.56 8.416 25.068 ;
  LAYER M3 ;
        RECT 8.384 22.58 8.416 22.612 ;
  LAYER M1 ;
        RECT 8.448 22.56 8.48 25.068 ;
  LAYER M3 ;
        RECT 8.448 25.016 8.48 25.048 ;
  LAYER M1 ;
        RECT 8.512 22.56 8.544 25.068 ;
  LAYER M3 ;
        RECT 8.512 22.58 8.544 22.612 ;
  LAYER M1 ;
        RECT 8.576 22.56 8.608 25.068 ;
  LAYER M3 ;
        RECT 8.576 25.016 8.608 25.048 ;
  LAYER M1 ;
        RECT 8.64 22.56 8.672 25.068 ;
  LAYER M3 ;
        RECT 8.64 22.58 8.672 22.612 ;
  LAYER M1 ;
        RECT 8.704 22.56 8.736 25.068 ;
  LAYER M3 ;
        RECT 8.704 25.016 8.736 25.048 ;
  LAYER M1 ;
        RECT 8.768 22.56 8.8 25.068 ;
  LAYER M3 ;
        RECT 6.4 22.644 6.432 22.676 ;
  LAYER M2 ;
        RECT 8.768 22.708 8.8 22.74 ;
  LAYER M2 ;
        RECT 6.4 22.772 6.432 22.804 ;
  LAYER M2 ;
        RECT 8.768 22.836 8.8 22.868 ;
  LAYER M2 ;
        RECT 6.4 22.9 6.432 22.932 ;
  LAYER M2 ;
        RECT 8.768 22.964 8.8 22.996 ;
  LAYER M2 ;
        RECT 6.4 23.028 6.432 23.06 ;
  LAYER M2 ;
        RECT 8.768 23.092 8.8 23.124 ;
  LAYER M2 ;
        RECT 6.4 23.156 6.432 23.188 ;
  LAYER M2 ;
        RECT 8.768 23.22 8.8 23.252 ;
  LAYER M2 ;
        RECT 6.4 23.284 6.432 23.316 ;
  LAYER M2 ;
        RECT 8.768 23.348 8.8 23.38 ;
  LAYER M2 ;
        RECT 6.4 23.412 6.432 23.444 ;
  LAYER M2 ;
        RECT 8.768 23.476 8.8 23.508 ;
  LAYER M2 ;
        RECT 6.4 23.54 6.432 23.572 ;
  LAYER M2 ;
        RECT 8.768 23.604 8.8 23.636 ;
  LAYER M2 ;
        RECT 6.4 23.668 6.432 23.7 ;
  LAYER M2 ;
        RECT 8.768 23.732 8.8 23.764 ;
  LAYER M2 ;
        RECT 6.4 23.796 6.432 23.828 ;
  LAYER M2 ;
        RECT 8.768 23.86 8.8 23.892 ;
  LAYER M2 ;
        RECT 6.4 23.924 6.432 23.956 ;
  LAYER M2 ;
        RECT 8.768 23.988 8.8 24.02 ;
  LAYER M2 ;
        RECT 6.4 24.052 6.432 24.084 ;
  LAYER M2 ;
        RECT 8.768 24.116 8.8 24.148 ;
  LAYER M2 ;
        RECT 6.4 24.18 6.432 24.212 ;
  LAYER M2 ;
        RECT 8.768 24.244 8.8 24.276 ;
  LAYER M2 ;
        RECT 6.4 24.308 6.432 24.34 ;
  LAYER M2 ;
        RECT 8.768 24.372 8.8 24.404 ;
  LAYER M2 ;
        RECT 6.4 24.436 6.432 24.468 ;
  LAYER M2 ;
        RECT 8.768 24.5 8.8 24.532 ;
  LAYER M2 ;
        RECT 6.4 24.564 6.432 24.596 ;
  LAYER M2 ;
        RECT 8.768 24.628 8.8 24.66 ;
  LAYER M2 ;
        RECT 6.4 24.692 6.432 24.724 ;
  LAYER M2 ;
        RECT 8.768 24.756 8.8 24.788 ;
  LAYER M2 ;
        RECT 6.4 24.82 6.432 24.852 ;
  LAYER M2 ;
        RECT 8.768 24.884 8.8 24.916 ;
  LAYER M2 ;
        RECT 6.352 22.512 8.848 25.116 ;
  END 
END Cap_60fF
