module testcase_EA_placer ( 0, 1 ); 
input 0, 1;

CMC_PMOS_S_n12_X1_Y1 m1 ( .G(0) );
CMC_PMOS_S_n12_X1_Y1 m2 ( .G(2) );
CMC_PMOS_S_n12_X1_Y1 m3 ( .G(2) );
CMC_PMOS_S_n12_X1_Y1 m4 ( .G(3) );
CMC_PMOS_S_n12_X1_Y1 m5 ( .G(3) );
CMC_PMOS_S_n12_X1_Y1 m6 ( .G(3) );
CMC_PMOS_S_n12_X1_Y1 m7 ( .G(3) );
CMC_PMOS_S_n12_X1_Y1 m8 ( .G(4) );
CMC_PMOS_S_n12_X1_Y1 m9 ( .G(4) );
CMC_PMOS_S_n12_X1_Y1 m10 ( .G(4) );
CMC_PMOS_S_n12_X1_Y1 m11 ( .G(4) );
CMC_PMOS_S_n12_X1_Y1 m12 ( .G(5) );
CMC_PMOS_S_n12_X1_Y1 m13 ( .G(5) );
CMC_PMOS_S_n12_X1_Y1 m14 ( .G(1) );

endmodule
