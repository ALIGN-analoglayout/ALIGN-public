.subckt common_source vin vop vccx vssx
mp0 vop vop vccx vccx p w=720e-9 nf=4 m=4
mn0 vop vin vssx vssx n w=720e-9 nf=4 m=4
.ends common_source
