MACRO switched_capacitor_filter
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_filter 0 0 ;
  SIZE 47.52 BY 39.48 ;
  PIN id
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.664 -0.016 23.696 0.016 ;
      LAYER M2 ;
        RECT 23.324 0.32 24.116 0.352 ;
      LAYER M2 ;
        RECT 23.664 0.32 23.696 0.352 ;
      LAYER M3 ;
        RECT 23.66 0 23.7 0.336 ;
      LAYER M2 ;
        RECT 23.664 -0.016 23.696 0.016 ;
    END
  END id
  PIN voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.824 39.464 15.856 39.496 ;
      LAYER M2 ;
        RECT 22.844 4.436 24.676 4.468 ;
      LAYER M2 ;
        RECT 22.684 3.008 25.316 3.04 ;
      LAYER M2 ;
        RECT 22.864 4.436 22.896 4.468 ;
      LAYER M3 ;
        RECT 22.86 3.024 22.9 4.452 ;
      LAYER M2 ;
        RECT 22.864 3.008 22.896 3.04 ;
      LAYER M2 ;
        RECT 7.964 0.824 8.036 0.856 ;
      LAYER M1 ;
        RECT 12.128 14.832 12.16 14.904 ;
      LAYER M2 ;
        RECT 12.108 14.852 12.18 14.884 ;
      LAYER M1 ;
        RECT 3.136 14.832 3.168 14.904 ;
      LAYER M2 ;
        RECT 3.116 14.852 3.188 14.884 ;
      LAYER M2 ;
        RECT 3.152 14.852 12.144 14.884 ;
      LAYER M2 ;
        RECT 7.984 0.824 8.016 0.856 ;
      LAYER M3 ;
        RECT 7.98 0.84 8.02 1.68 ;
      LAYER M4 ;
        RECT 8 1.66 8.16 1.7 ;
      LAYER M5 ;
        RECT 8.128 1.68 8.192 14.868 ;
      LAYER M4 ;
        RECT 8.14 14.848 8.18 14.888 ;
      LAYER M3 ;
        RECT 8.14 14.848 8.18 14.888 ;
      LAYER M2 ;
        RECT 8.144 14.852 8.176 14.884 ;
      LAYER M1 ;
        RECT 22.176 39.024 22.208 39.096 ;
      LAYER M2 ;
        RECT 22.156 39.044 22.228 39.076 ;
      LAYER M1 ;
        RECT 25.152 39.024 25.184 39.096 ;
      LAYER M2 ;
        RECT 25.132 39.044 25.204 39.076 ;
      LAYER M2 ;
        RECT 22.192 39.044 25.168 39.076 ;
      LAYER M2 ;
        RECT 22.704 3.008 22.736 3.04 ;
      LAYER M3 ;
        RECT 22.7 1.68 22.74 3.024 ;
      LAYER M4 ;
        RECT 8.16 1.66 22.72 1.7 ;
      LAYER M2 ;
        RECT 12.144 14.852 12.176 14.884 ;
      LAYER M3 ;
        RECT 12.14 14.868 12.18 16.8 ;
      LAYER M4 ;
        RECT 12.16 16.78 16.48 16.82 ;
      LAYER M3 ;
        RECT 16.46 16.8 16.5 36.96 ;
      LAYER M4 ;
        RECT 16.48 36.94 22.16 36.98 ;
      LAYER M3 ;
        RECT 22.14 36.96 22.18 39.06 ;
      LAYER M2 ;
        RECT 22.144 39.044 22.176 39.076 ;
      LAYER M3 ;
        RECT 16.46 36.96 16.5 39.48 ;
      LAYER M4 ;
        RECT 15.84 39.46 16.48 39.5 ;
      LAYER M3 ;
        RECT 15.82 39.46 15.86 39.5 ;
      LAYER M2 ;
        RECT 15.824 39.464 15.856 39.496 ;
    END
  END voutn
  PIN voutp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.664 39.464 31.696 39.496 ;
      LAYER M2 ;
        RECT 23.484 4.268 24.036 4.3 ;
      LAYER M2 ;
        RECT 22.044 3.176 24.676 3.208 ;
      LAYER M2 ;
        RECT 23.584 4.268 23.616 4.3 ;
      LAYER M3 ;
        RECT 23.58 3.192 23.62 4.284 ;
      LAYER M2 ;
        RECT 23.584 3.176 23.616 3.208 ;
      LAYER M2 ;
        RECT 39.484 0.824 39.556 0.856 ;
      LAYER M1 ;
        RECT 35.36 14.832 35.392 14.904 ;
      LAYER M2 ;
        RECT 35.34 14.852 35.412 14.884 ;
      LAYER M1 ;
        RECT 44.352 14.832 44.384 14.904 ;
      LAYER M2 ;
        RECT 44.332 14.852 44.404 14.884 ;
      LAYER M2 ;
        RECT 35.376 14.852 44.368 14.884 ;
      LAYER M2 ;
        RECT 39.504 0.824 39.536 0.856 ;
      LAYER M3 ;
        RECT 39.5 0.84 39.54 1.68 ;
      LAYER M4 ;
        RECT 39.36 1.66 39.52 1.7 ;
      LAYER M5 ;
        RECT 39.328 1.68 39.392 14.868 ;
      LAYER M4 ;
        RECT 39.34 14.848 39.38 14.888 ;
      LAYER M3 ;
        RECT 39.34 14.848 39.38 14.888 ;
      LAYER M2 ;
        RECT 39.344 14.852 39.376 14.884 ;
      LAYER M1 ;
        RECT 19.2 39.192 19.232 39.264 ;
      LAYER M2 ;
        RECT 19.18 39.212 19.252 39.244 ;
      LAYER M1 ;
        RECT 28.128 39.192 28.16 39.264 ;
      LAYER M2 ;
        RECT 28.108 39.212 28.18 39.244 ;
      LAYER M2 ;
        RECT 19.216 39.212 28.144 39.244 ;
      LAYER M2 ;
        RECT 24.624 3.176 24.656 3.208 ;
      LAYER M3 ;
        RECT 24.62 1.596 24.66 3.192 ;
      LAYER M4 ;
        RECT 24.64 1.576 39.312 1.616 ;
      LAYER M5 ;
        RECT 39.28 1.596 39.344 1.68 ;
      LAYER M5 ;
        RECT 39.28 1.68 39.344 1.744 ;
      LAYER M5 ;
        RECT 39.312 1.68 39.36 1.744 ;
      LAYER M2 ;
        RECT 35.344 14.852 35.376 14.884 ;
      LAYER M3 ;
        RECT 35.34 14.868 35.38 16.8 ;
      LAYER M4 ;
        RECT 32.112 16.78 35.36 16.82 ;
      LAYER M5 ;
        RECT 32.08 16.8 32.144 36.72 ;
      LAYER M6 ;
        RECT 30.384 36.688 32.112 36.752 ;
      LAYER M5 ;
        RECT 30.352 36.72 30.416 39.228 ;
      LAYER M4 ;
        RECT 28.16 39.208 30.384 39.248 ;
      LAYER M3 ;
        RECT 28.14 39.208 28.18 39.248 ;
      LAYER M2 ;
        RECT 28.144 39.212 28.176 39.244 ;
      LAYER M4 ;
        RECT 30.32 39.208 31.68 39.248 ;
      LAYER M3 ;
        RECT 31.66 39.228 31.7 39.48 ;
      LAYER M2 ;
        RECT 31.664 39.464 31.696 39.496 ;
    END
  END voutp
  PIN vss
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.824 -0.016 23.856 0.016 ;
      LAYER M2 ;
        RECT 21.564 0.236 26.116 0.268 ;
      LAYER M1 ;
        RECT 22.4 19.872 22.432 19.944 ;
      LAYER M2 ;
        RECT 22.38 19.892 22.452 19.924 ;
      LAYER M1 ;
        RECT 25.312 19.872 25.344 19.944 ;
      LAYER M2 ;
        RECT 25.292 19.892 25.364 19.924 ;
      LAYER M2 ;
        RECT 22.416 19.892 25.328 19.924 ;
      LAYER M1 ;
        RECT 19.36 19.704 19.392 19.776 ;
      LAYER M2 ;
        RECT 19.34 19.724 19.412 19.756 ;
      LAYER M1 ;
        RECT 28.352 19.704 28.384 19.776 ;
      LAYER M2 ;
        RECT 28.332 19.724 28.404 19.756 ;
      LAYER M2 ;
        RECT 19.376 19.724 28.368 19.756 ;
      LAYER M2 ;
        RECT 23.824 0.236 23.856 0.268 ;
      LAYER M3 ;
        RECT 23.82 0 23.86 0.252 ;
      LAYER M2 ;
        RECT 23.824 -0.016 23.856 0.016 ;
      LAYER M2 ;
        RECT 25.024 0.236 25.056 0.268 ;
      LAYER M3 ;
        RECT 25.02 0.252 25.06 19.908 ;
      LAYER M2 ;
        RECT 25.024 19.892 25.056 19.924 ;
      LAYER M3 ;
        RECT 25.02 19.72 25.06 19.76 ;
      LAYER M2 ;
        RECT 25.024 19.724 25.056 19.756 ;
    END
  END vss
  PIN vinn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.744 -0.016 15.776 0.016 ;
      LAYER M2 ;
        RECT 15.724 0.236 15.796 0.268 ;
      LAYER M1 ;
        RECT 28.288 5.844 28.32 5.916 ;
      LAYER M2 ;
        RECT 28.268 5.864 28.34 5.896 ;
      LAYER M1 ;
        RECT 19.36 5.844 19.392 5.916 ;
      LAYER M2 ;
        RECT 19.34 5.864 19.412 5.896 ;
      LAYER M2 ;
        RECT 19.376 5.864 28.304 5.896 ;
      LAYER M2 ;
        RECT 15.744 0.236 15.776 0.268 ;
      LAYER M3 ;
        RECT 15.74 0 15.78 0.252 ;
      LAYER M2 ;
        RECT 15.744 -0.016 15.776 0.016 ;
      LAYER M3 ;
        RECT 15.74 0.252 15.78 5.88 ;
      LAYER M4 ;
        RECT 15.76 5.86 19.36 5.9 ;
      LAYER M3 ;
        RECT 19.34 5.86 19.38 5.9 ;
      LAYER M2 ;
        RECT 19.344 5.864 19.376 5.896 ;
    END
  END vinn
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.904 -0.016 15.936 0.016 ;
      LAYER M2 ;
        RECT 5.244 0.236 5.316 0.268 ;
      LAYER M2 ;
        RECT 5.964 0.74 6.036 0.772 ;
      LAYER M2 ;
        RECT 7.324 0.74 7.396 0.772 ;
      LAYER M2 ;
        RECT 5.264 0.236 5.296 0.268 ;
      LAYER M3 ;
        RECT 5.26 0.252 5.3 0.756 ;
      LAYER M4 ;
        RECT 5.28 0.736 6 0.776 ;
      LAYER M3 ;
        RECT 5.98 0.736 6.02 0.776 ;
      LAYER M2 ;
        RECT 5.984 0.74 6.016 0.772 ;
      LAYER M4 ;
        RECT 6 0.736 7.36 0.776 ;
      LAYER M3 ;
        RECT 7.34 0.736 7.38 0.776 ;
      LAYER M2 ;
        RECT 7.344 0.74 7.376 0.772 ;
      LAYER M2 ;
        RECT 42.204 0.236 42.276 0.268 ;
      LAYER M2 ;
        RECT 41.484 0.74 41.556 0.772 ;
      LAYER M2 ;
        RECT 40.124 0.74 40.196 0.772 ;
      LAYER M2 ;
        RECT 42.224 0.236 42.256 0.268 ;
      LAYER M3 ;
        RECT 42.22 0.252 42.26 0.756 ;
      LAYER M4 ;
        RECT 41.52 0.736 42.24 0.776 ;
      LAYER M3 ;
        RECT 41.5 0.736 41.54 0.776 ;
      LAYER M2 ;
        RECT 41.504 0.74 41.536 0.772 ;
      LAYER M4 ;
        RECT 40.16 0.736 41.52 0.776 ;
      LAYER M3 ;
        RECT 40.14 0.736 40.18 0.776 ;
      LAYER M2 ;
        RECT 40.144 0.74 40.176 0.772 ;
      LAYER M4 ;
        RECT 7.26 0.736 7.3 0.776 ;
      LAYER M3 ;
        RECT 7.26 0.756 7.3 1.68 ;
      LAYER M2 ;
        RECT 7.28 1.664 15.92 1.696 ;
      LAYER M3 ;
        RECT 15.9 0 15.94 1.68 ;
      LAYER M2 ;
        RECT 15.904 -0.016 15.936 0.016 ;
      LAYER M3 ;
        RECT 15.9 1.68 15.94 1.764 ;
      LAYER M2 ;
        RECT 15.92 1.748 22.64 1.78 ;
      LAYER M3 ;
        RECT 22.62 1.744 22.66 1.784 ;
      LAYER M4 ;
        RECT 22.64 1.744 40.176 1.784 ;
      LAYER M5 ;
        RECT 40.144 0.756 40.208 1.764 ;
      LAYER M4 ;
        RECT 40.156 0.736 40.196 0.776 ;
    END
  END agnd
  PIN vinp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.744 -0.016 31.776 0.016 ;
      LAYER M2 ;
        RECT 31.724 0.236 31.796 0.268 ;
      LAYER M1 ;
        RECT 25.312 6.012 25.344 6.084 ;
      LAYER M2 ;
        RECT 25.292 6.032 25.364 6.064 ;
      LAYER M1 ;
        RECT 22.336 6.012 22.368 6.084 ;
      LAYER M2 ;
        RECT 22.316 6.032 22.388 6.064 ;
      LAYER M2 ;
        RECT 22.352 6.032 25.328 6.064 ;
      LAYER M2 ;
        RECT 31.744 0.236 31.776 0.268 ;
      LAYER M3 ;
        RECT 31.74 0.252 31.78 3.276 ;
      LAYER M2 ;
        RECT 26.88 3.26 31.76 3.292 ;
      LAYER M3 ;
        RECT 26.86 3.276 26.9 6.048 ;
      LAYER M4 ;
        RECT 25.36 6.028 26.88 6.068 ;
      LAYER M3 ;
        RECT 25.34 6.028 25.38 6.068 ;
      LAYER M2 ;
        RECT 25.344 6.032 25.376 6.064 ;
      LAYER M3 ;
        RECT 31.74 0 31.78 0.252 ;
      LAYER M2 ;
        RECT 31.744 -0.016 31.776 0.016 ;
    END
  END vinp
  OBS 
  LAYER M2 ;
        RECT 22.124 3.26 25.396 3.292 ;
  LAYER M2 ;
        RECT 21.484 0.488 26.036 0.52 ;
  LAYER M2 ;
        RECT 23.404 5.024 24.116 5.056 ;
  LAYER M2 ;
        RECT 22.764 4.184 24.756 4.216 ;
  LAYER M2 ;
        RECT 23.484 4.772 24.196 4.804 ;
  LAYER M3 ;
        RECT 23.5 1.56 23.54 2.472 ;
  LAYER M2 ;
        RECT 40.844 0.824 40.916 0.856 ;
  LAYER M1 ;
        RECT 35.2 31.212 35.232 31.284 ;
  LAYER M2 ;
        RECT 35.18 31.232 35.252 31.264 ;
  LAYER M1 ;
        RECT 44.128 31.212 44.16 31.284 ;
  LAYER M2 ;
        RECT 44.108 31.232 44.18 31.264 ;
  LAYER M2 ;
        RECT 35.216 31.232 44.144 31.264 ;
  LAYER M2 ;
        RECT 40.864 0.824 40.896 0.856 ;
  LAYER M3 ;
        RECT 40.86 0.84 40.9 1.68 ;
  LAYER M2 ;
        RECT 40.88 1.664 41.04 1.696 ;
  LAYER M3 ;
        RECT 41.02 1.68 41.06 31.248 ;
  LAYER M2 ;
        RECT 41.024 31.232 41.056 31.264 ;
  LAYER M1 ;
        RECT 28.128 19.116 28.16 19.188 ;
  LAYER M2 ;
        RECT 28.108 19.136 28.18 19.168 ;
  LAYER M1 ;
        RECT 19.136 19.116 19.168 19.188 ;
  LAYER M2 ;
        RECT 19.116 19.136 19.188 19.168 ;
  LAYER M2 ;
        RECT 19.152 19.136 28.144 19.168 ;
  LAYER M3 ;
        RECT 23.5 2.416 23.54 2.456 ;
  LAYER M4 ;
        RECT 23.52 2.416 25.2 2.456 ;
  LAYER M3 ;
        RECT 25.18 2.436 25.22 18.564 ;
  LAYER M2 ;
        RECT 25.2 18.548 41.04 18.58 ;
  LAYER M3 ;
        RECT 41.02 18.544 41.06 18.584 ;
  LAYER M3 ;
        RECT 25.18 18.564 25.22 19.152 ;
  LAYER M2 ;
        RECT 25.184 19.136 25.216 19.168 ;
  LAYER M3 ;
        RECT 23.82 1.476 23.86 2.388 ;
  LAYER M2 ;
        RECT 6.604 0.824 6.676 0.856 ;
  LAYER M1 ;
        RECT 12.288 31.212 12.32 31.284 ;
  LAYER M2 ;
        RECT 12.268 31.232 12.34 31.264 ;
  LAYER M1 ;
        RECT 3.36 31.212 3.392 31.284 ;
  LAYER M2 ;
        RECT 3.34 31.232 3.412 31.264 ;
  LAYER M2 ;
        RECT 3.376 31.232 12.304 31.264 ;
  LAYER M2 ;
        RECT 6.624 0.824 6.656 0.856 ;
  LAYER M3 ;
        RECT 6.62 0.84 6.66 1.68 ;
  LAYER M2 ;
        RECT 6.48 1.664 6.64 1.696 ;
  LAYER M3 ;
        RECT 6.46 1.68 6.5 31.248 ;
  LAYER M2 ;
        RECT 6.464 31.232 6.496 31.264 ;
  LAYER M1 ;
        RECT 25.088 18.948 25.12 19.02 ;
  LAYER M2 ;
        RECT 25.068 18.968 25.14 19 ;
  LAYER M1 ;
        RECT 22.176 18.948 22.208 19.02 ;
  LAYER M2 ;
        RECT 22.156 18.968 22.228 19 ;
  LAYER M2 ;
        RECT 22.192 18.968 25.104 19 ;
  LAYER M3 ;
        RECT 23.82 2.332 23.86 2.372 ;
  LAYER M4 ;
        RECT 22.08 2.332 23.84 2.372 ;
  LAYER M3 ;
        RECT 22.06 2.352 22.1 18.564 ;
  LAYER M2 ;
        RECT 6.48 18.548 22.08 18.58 ;
  LAYER M3 ;
        RECT 6.46 18.544 6.5 18.584 ;
  LAYER M3 ;
        RECT 22.06 18.564 22.1 18.984 ;
  LAYER M4 ;
        RECT 22.08 18.964 22.16 19.004 ;
  LAYER M3 ;
        RECT 22.14 18.964 22.18 19.004 ;
  LAYER M2 ;
        RECT 22.144 18.968 22.176 19 ;
  LAYER M2 ;
        RECT 15.644 0.404 15.716 0.436 ;
  LAYER M2 ;
        RECT 6.684 0.656 6.756 0.688 ;
  LAYER M2 ;
        RECT 8.044 0.656 8.116 0.688 ;
  LAYER M2 ;
        RECT 15.664 0.404 15.696 0.436 ;
  LAYER M3 ;
        RECT 15.66 0.42 15.7 0.588 ;
  LAYER M2 ;
        RECT 8.08 0.572 15.68 0.604 ;
  LAYER M3 ;
        RECT 8.06 0.588 8.1 0.672 ;
  LAYER M2 ;
        RECT 8.064 0.656 8.096 0.688 ;
  LAYER M3 ;
        RECT 8.06 0.652 8.1 0.692 ;
  LAYER M4 ;
        RECT 6.72 0.652 8.08 0.692 ;
  LAYER M3 ;
        RECT 6.7 0.652 6.74 0.692 ;
  LAYER M2 ;
        RECT 6.704 0.656 6.736 0.688 ;
  LAYER M2 ;
        RECT 31.804 0.404 31.876 0.436 ;
  LAYER M2 ;
        RECT 40.764 0.656 40.836 0.688 ;
  LAYER M2 ;
        RECT 39.404 0.656 39.476 0.688 ;
  LAYER M2 ;
        RECT 31.824 0.404 31.856 0.436 ;
  LAYER M3 ;
        RECT 31.82 0.42 31.86 0.588 ;
  LAYER M2 ;
        RECT 31.84 0.572 39.44 0.604 ;
  LAYER M3 ;
        RECT 39.42 0.588 39.46 0.672 ;
  LAYER M2 ;
        RECT 39.424 0.656 39.456 0.688 ;
  LAYER M3 ;
        RECT 39.42 0.652 39.46 0.692 ;
  LAYER M4 ;
        RECT 39.44 0.652 40.8 0.692 ;
  LAYER M3 ;
        RECT 40.78 0.652 40.82 0.692 ;
  LAYER M2 ;
        RECT 40.784 0.656 40.816 0.688 ;
  LAYER M2 ;
        RECT 15.184 0.572 15.216 0.604 ;
  LAYER M3 ;
        RECT 15.18 0.568 15.22 0.608 ;
  LAYER M4 ;
        RECT 15.12 0.568 15.2 0.608 ;
  LAYER M5 ;
        RECT 15.088 0.588 15.152 6.72 ;
  LAYER M4 ;
        RECT 15.12 6.7 30.24 6.74 ;
  LAYER M5 ;
        RECT 30.208 5.124 30.272 6.72 ;
  LAYER M4 ;
        RECT 30.24 5.104 31.84 5.144 ;
  LAYER M3 ;
        RECT 31.82 3.36 31.86 5.124 ;
  LAYER M2 ;
        RECT 31.84 3.344 32 3.376 ;
  LAYER M3 ;
        RECT 31.98 0.588 32.02 3.36 ;
  LAYER M2 ;
        RECT 31.984 0.572 32.016 0.604 ;
  LAYER M2 ;
        RECT 5.324 0.404 5.396 0.436 ;
  LAYER M2 ;
        RECT 6.044 0.572 6.116 0.604 ;
  LAYER M2 ;
        RECT 7.404 0.572 7.476 0.604 ;
  LAYER M2 ;
        RECT 5.344 0.404 5.376 0.436 ;
  LAYER M3 ;
        RECT 5.34 0.42 5.38 0.588 ;
  LAYER M4 ;
        RECT 5.36 0.568 6.08 0.608 ;
  LAYER M3 ;
        RECT 6.06 0.568 6.1 0.608 ;
  LAYER M2 ;
        RECT 6.064 0.572 6.096 0.604 ;
  LAYER M4 ;
        RECT 6.08 0.568 7.44 0.608 ;
  LAYER M3 ;
        RECT 7.42 0.568 7.46 0.608 ;
  LAYER M2 ;
        RECT 7.424 0.572 7.456 0.604 ;
  LAYER M2 ;
        RECT 42.124 0.404 42.196 0.436 ;
  LAYER M2 ;
        RECT 41.404 0.572 41.476 0.604 ;
  LAYER M2 ;
        RECT 40.044 0.572 40.116 0.604 ;
  LAYER M2 ;
        RECT 42.144 0.404 42.176 0.436 ;
  LAYER M3 ;
        RECT 42.14 0.42 42.18 0.588 ;
  LAYER M4 ;
        RECT 41.44 0.568 42.16 0.608 ;
  LAYER M3 ;
        RECT 41.42 0.568 41.46 0.608 ;
  LAYER M2 ;
        RECT 41.424 0.572 41.456 0.604 ;
  LAYER M4 ;
        RECT 40.08 0.568 41.44 0.608 ;
  LAYER M3 ;
        RECT 40.06 0.568 40.1 0.608 ;
  LAYER M2 ;
        RECT 40.064 0.572 40.096 0.604 ;
  LAYER M4 ;
        RECT 7.44 0.568 8.352 0.608 ;
  LAYER M5 ;
        RECT 8.32 0.588 8.384 3.36 ;
  LAYER M4 ;
        RECT 8.352 3.34 38.592 3.38 ;
  LAYER M5 ;
        RECT 38.56 0.84 38.624 3.36 ;
  LAYER M4 ;
        RECT 38.592 0.82 40.24 0.86 ;
  LAYER M3 ;
        RECT 40.22 0.588 40.26 0.84 ;
  LAYER M4 ;
        RECT 40.22 0.568 40.26 0.608 ;
  LAYER M2 ;
        RECT 23.964 4.856 24.036 4.888 ;
  LAYER M2 ;
        RECT 23.324 4.352 24.196 4.384 ;
  LAYER M2 ;
        RECT 23.984 4.856 24.016 4.888 ;
  LAYER M3 ;
        RECT 23.98 4.368 24.02 4.872 ;
  LAYER M2 ;
        RECT 23.984 4.352 24.016 4.384 ;
  LAYER M2 ;
        RECT 23.324 4.94 23.396 4.972 ;
  LAYER M2 ;
        RECT 22.684 4.52 24.836 4.552 ;
  LAYER M2 ;
        RECT 23.344 4.94 23.376 4.972 ;
  LAYER M3 ;
        RECT 23.34 4.536 23.38 4.956 ;
  LAYER M2 ;
        RECT 23.344 4.52 23.376 4.552 ;
  LAYER M3 ;
        RECT 23.58 1.728 23.62 2.64 ;
  LAYER M2 ;
        RECT 22.204 3.092 24.836 3.124 ;
  LAYER M3 ;
        RECT 23.58 2.584 23.62 2.624 ;
  LAYER M4 ;
        RECT 23.52 2.584 23.6 2.624 ;
  LAYER M3 ;
        RECT 23.5 2.604 23.54 3.108 ;
  LAYER M2 ;
        RECT 23.504 3.092 23.536 3.124 ;
  LAYER M3 ;
        RECT 23.66 1.812 23.7 2.724 ;
  LAYER M2 ;
        RECT 21.404 0.404 25.956 0.436 ;
  LAYER M3 ;
        RECT 23.66 1.828 23.7 1.868 ;
  LAYER M4 ;
        RECT 23.44 1.828 23.68 1.868 ;
  LAYER M3 ;
        RECT 23.42 0.42 23.46 1.848 ;
  LAYER M2 ;
        RECT 23.424 0.404 23.456 0.436 ;
  LAYER M3 ;
        RECT 23.74 1.644 23.78 2.556 ;
  LAYER M2 ;
        RECT 22.844 2.924 25.476 2.956 ;
  LAYER M3 ;
        RECT 23.74 2.5 23.78 2.54 ;
  LAYER M4 ;
        RECT 23.76 2.5 23.84 2.54 ;
  LAYER M3 ;
        RECT 23.82 2.52 23.86 2.94 ;
  LAYER M2 ;
        RECT 23.824 2.924 23.856 2.956 ;
  LAYER M1 ;
        RECT 24.064 4.752 24.096 5.412 ;
  LAYER M1 ;
        RECT 23.424 4.752 23.456 5.412 ;
  LAYER M1 ;
        RECT 24.144 4.752 24.176 5.412 ;
  LAYER M1 ;
        RECT 23.504 4.752 23.536 5.412 ;
  LAYER M1 ;
        RECT 23.984 4.752 24.016 5.412 ;
  LAYER M1 ;
        RECT 23.344 5.192 23.376 5.224 ;
  LAYER M1 ;
        RECT 22.144 2.064 22.176 2.724 ;
  LAYER M1 ;
        RECT 22.144 1.224 22.176 1.884 ;
  LAYER M1 ;
        RECT 23.424 2.064 23.456 2.724 ;
  LAYER M1 ;
        RECT 23.424 1.224 23.456 1.884 ;
  LAYER M1 ;
        RECT 24.704 2.064 24.736 2.724 ;
  LAYER M1 ;
        RECT 24.704 1.224 24.736 1.884 ;
  LAYER M1 ;
        RECT 22.784 2.064 22.816 2.724 ;
  LAYER M1 ;
        RECT 22.784 1.224 22.816 1.884 ;
  LAYER M1 ;
        RECT 24.064 2.064 24.096 2.724 ;
  LAYER M1 ;
        RECT 24.064 1.224 24.096 1.884 ;
  LAYER M1 ;
        RECT 25.344 2.064 25.376 2.724 ;
  LAYER M1 ;
        RECT 25.344 1.224 25.376 1.884 ;
  LAYER M1 ;
        RECT 22.064 2.064 22.096 2.724 ;
  LAYER M1 ;
        RECT 22.064 1.224 22.096 1.884 ;
  LAYER M1 ;
        RECT 23.344 2.064 23.376 2.724 ;
  LAYER M1 ;
        RECT 23.344 1.224 23.376 1.884 ;
  LAYER M1 ;
        RECT 24.624 2.064 24.656 2.724 ;
  LAYER M1 ;
        RECT 24.624 1.224 24.656 1.884 ;
  LAYER M1 ;
        RECT 22.704 2.064 22.736 2.724 ;
  LAYER M1 ;
        RECT 22.704 1.224 22.736 1.884 ;
  LAYER M1 ;
        RECT 23.984 2.064 24.016 2.724 ;
  LAYER M1 ;
        RECT 23.984 1.224 24.016 1.884 ;
  LAYER M1 ;
        RECT 25.264 2.064 25.296 2.724 ;
  LAYER M1 ;
        RECT 25.264 1.224 25.296 1.884 ;
  LAYER M1 ;
        RECT 22.224 2.064 22.256 2.724 ;
  LAYER M1 ;
        RECT 22.224 1.224 22.256 1.884 ;
  LAYER M1 ;
        RECT 23.504 2.064 23.536 2.724 ;
  LAYER M1 ;
        RECT 23.504 1.224 23.536 1.884 ;
  LAYER M1 ;
        RECT 24.784 2.064 24.816 2.724 ;
  LAYER M1 ;
        RECT 24.784 1.224 24.816 1.884 ;
  LAYER M1 ;
        RECT 22.864 2.064 22.896 2.724 ;
  LAYER M1 ;
        RECT 22.864 1.224 22.896 1.884 ;
  LAYER M1 ;
        RECT 24.144 2.064 24.176 2.724 ;
  LAYER M1 ;
        RECT 24.144 1.224 24.176 1.884 ;
  LAYER M1 ;
        RECT 25.424 2.064 25.456 2.724 ;
  LAYER M1 ;
        RECT 25.424 1.224 25.456 1.884 ;
  LAYER M2 ;
        RECT 22.044 2.672 25.316 2.704 ;
  LAYER M2 ;
        RECT 22.204 2.588 24.836 2.62 ;
  LAYER M2 ;
        RECT 22.844 2.504 25.476 2.536 ;
  LAYER M2 ;
        RECT 22.124 2.42 24.756 2.452 ;
  LAYER M2 ;
        RECT 22.764 2.336 25.396 2.368 ;
  LAYER M2 ;
        RECT 22.044 1.832 25.316 1.864 ;
  LAYER M2 ;
        RECT 22.844 1.748 25.476 1.78 ;
  LAYER M2 ;
        RECT 22.204 1.664 24.836 1.696 ;
  LAYER M2 ;
        RECT 22.764 1.58 25.396 1.612 ;
  LAYER M2 ;
        RECT 25.424 1.412 25.456 1.444 ;
  LAYER M1 ;
        RECT 24.064 0.216 24.096 0.876 ;
  LAYER M1 ;
        RECT 23.424 0.216 23.456 0.876 ;
  LAYER M1 ;
        RECT 25.984 0.216 26.016 0.876 ;
  LAYER M1 ;
        RECT 25.344 0.216 25.376 0.876 ;
  LAYER M1 ;
        RECT 24.704 0.216 24.736 0.876 ;
  LAYER M1 ;
        RECT 22.784 0.216 22.816 0.876 ;
  LAYER M1 ;
        RECT 22.144 0.216 22.176 0.876 ;
  LAYER M1 ;
        RECT 21.504 0.216 21.536 0.876 ;
  LAYER M1 ;
        RECT 24.144 0.216 24.176 0.876 ;
  LAYER M1 ;
        RECT 23.504 0.216 23.536 0.876 ;
  LAYER M1 ;
        RECT 26.064 0.216 26.096 0.876 ;
  LAYER M1 ;
        RECT 25.424 0.216 25.456 0.876 ;
  LAYER M1 ;
        RECT 24.784 0.216 24.816 0.876 ;
  LAYER M1 ;
        RECT 22.864 0.216 22.896 0.876 ;
  LAYER M1 ;
        RECT 22.224 0.216 22.256 0.876 ;
  LAYER M1 ;
        RECT 21.584 0.216 21.616 0.876 ;
  LAYER M1 ;
        RECT 23.984 0.216 24.016 0.876 ;
  LAYER M1 ;
        RECT 23.344 0.216 23.376 0.876 ;
  LAYER M1 ;
        RECT 25.904 0.216 25.936 0.876 ;
  LAYER M1 ;
        RECT 25.264 0.216 25.296 0.876 ;
  LAYER M1 ;
        RECT 24.624 0.216 24.656 0.876 ;
  LAYER M1 ;
        RECT 22.704 0.216 22.736 0.876 ;
  LAYER M1 ;
        RECT 22.064 0.216 22.096 0.876 ;
  LAYER M1 ;
        RECT 21.424 0.656 21.456 0.688 ;
  LAYER M1 ;
        RECT 22.784 3.912 22.816 4.572 ;
  LAYER M1 ;
        RECT 24.704 3.912 24.736 4.572 ;
  LAYER M1 ;
        RECT 23.424 3.912 23.456 4.572 ;
  LAYER M1 ;
        RECT 24.064 3.912 24.096 4.572 ;
  LAYER M1 ;
        RECT 22.704 3.912 22.736 4.572 ;
  LAYER M1 ;
        RECT 24.784 3.912 24.816 4.572 ;
  LAYER M1 ;
        RECT 23.344 3.912 23.376 4.572 ;
  LAYER M1 ;
        RECT 24.144 3.912 24.176 4.572 ;
  LAYER M1 ;
        RECT 22.864 3.912 22.896 4.572 ;
  LAYER M1 ;
        RECT 24.624 3.912 24.656 4.572 ;
  LAYER M1 ;
        RECT 23.504 3.912 23.536 4.572 ;
  LAYER M1 ;
        RECT 23.984 4.1 24.016 4.132 ;
  LAYER M1 ;
        RECT 25.344 2.904 25.376 3.564 ;
  LAYER M1 ;
        RECT 24.064 2.904 24.096 3.564 ;
  LAYER M1 ;
        RECT 22.784 2.904 22.816 3.564 ;
  LAYER M1 ;
        RECT 24.704 2.904 24.736 3.564 ;
  LAYER M1 ;
        RECT 23.424 2.904 23.456 3.564 ;
  LAYER M1 ;
        RECT 22.144 2.904 22.176 3.564 ;
  LAYER M1 ;
        RECT 25.424 2.904 25.456 3.564 ;
  LAYER M1 ;
        RECT 24.144 2.904 24.176 3.564 ;
  LAYER M1 ;
        RECT 22.864 2.904 22.896 3.564 ;
  LAYER M1 ;
        RECT 24.784 2.904 24.816 3.564 ;
  LAYER M1 ;
        RECT 23.504 2.904 23.536 3.564 ;
  LAYER M1 ;
        RECT 22.224 2.904 22.256 3.564 ;
  LAYER M1 ;
        RECT 25.264 2.904 25.296 3.564 ;
  LAYER M1 ;
        RECT 23.984 2.904 24.016 3.564 ;
  LAYER M1 ;
        RECT 22.704 2.904 22.736 3.564 ;
  LAYER M1 ;
        RECT 24.624 2.904 24.656 3.564 ;
  LAYER M1 ;
        RECT 23.344 2.904 23.376 3.564 ;
  LAYER M1 ;
        RECT 22.064 3.344 22.096 3.376 ;
  LAYER M1 ;
        RECT 6.48 14.244 6.512 14.316 ;
  LAYER M2 ;
        RECT 6.46 14.264 6.532 14.296 ;
  LAYER M1 ;
        RECT 9.392 14.244 9.424 14.316 ;
  LAYER M2 ;
        RECT 9.372 14.264 9.444 14.296 ;
  LAYER M2 ;
        RECT 6.496 14.264 9.408 14.296 ;
  LAYER M2 ;
        RECT 6.124 0.908 6.836 0.94 ;
  LAYER M1 ;
        RECT 9.312 31.044 9.344 31.116 ;
  LAYER M2 ;
        RECT 9.292 31.064 9.364 31.096 ;
  LAYER M1 ;
        RECT 6.336 31.044 6.368 31.116 ;
  LAYER M2 ;
        RECT 6.316 31.064 6.388 31.096 ;
  LAYER M2 ;
        RECT 6.352 31.064 9.328 31.096 ;
  LAYER M2 ;
        RECT 6.544 14.264 6.576 14.296 ;
  LAYER M3 ;
        RECT 6.54 0.924 6.58 14.28 ;
  LAYER M2 ;
        RECT 6.544 0.908 6.576 0.94 ;
  LAYER M2 ;
        RECT 9.344 14.264 9.376 14.296 ;
  LAYER M3 ;
        RECT 9.34 14.28 9.38 31.08 ;
  LAYER M2 ;
        RECT 9.344 31.064 9.376 31.096 ;
  LAYER M1 ;
        RECT 6.256 1.308 6.288 1.38 ;
  LAYER M2 ;
        RECT 6.236 1.328 6.308 1.36 ;
  LAYER M1 ;
        RECT 9.232 1.308 9.264 1.38 ;
  LAYER M2 ;
        RECT 9.212 1.328 9.284 1.36 ;
  LAYER M2 ;
        RECT 6.272 1.328 9.248 1.36 ;
  LAYER M2 ;
        RECT 5.404 0.32 5.476 0.352 ;
  LAYER M2 ;
        RECT 15.564 0.32 15.636 0.352 ;
  LAYER M2 ;
        RECT 6.224 1.328 6.256 1.36 ;
  LAYER M3 ;
        RECT 6.22 0.336 6.26 1.344 ;
  LAYER M4 ;
        RECT 5.44 0.316 6.24 0.356 ;
  LAYER M3 ;
        RECT 5.42 0.316 5.46 0.356 ;
  LAYER M2 ;
        RECT 5.424 0.32 5.456 0.352 ;
  LAYER M2 ;
        RECT 9.264 1.328 9.296 1.36 ;
  LAYER M3 ;
        RECT 9.26 0.336 9.3 1.344 ;
  LAYER M4 ;
        RECT 9.28 0.316 15.6 0.356 ;
  LAYER M3 ;
        RECT 15.58 0.316 15.62 0.356 ;
  LAYER M2 ;
        RECT 15.584 0.32 15.616 0.352 ;
  LAYER M2 ;
        RECT 7.484 0.908 8.196 0.94 ;
  LAYER M1 ;
        RECT 9.088 15 9.12 15.072 ;
  LAYER M2 ;
        RECT 9.068 15.02 9.14 15.052 ;
  LAYER M1 ;
        RECT 6.176 15 6.208 15.072 ;
  LAYER M2 ;
        RECT 6.156 15.02 6.228 15.052 ;
  LAYER M2 ;
        RECT 6.192 15.02 9.104 15.052 ;
  LAYER M2 ;
        RECT 7.504 0.908 7.536 0.94 ;
  LAYER M3 ;
        RECT 7.5 0.924 7.54 1.68 ;
  LAYER M4 ;
        RECT 7.44 1.66 7.52 1.7 ;
  LAYER M5 ;
        RECT 7.408 1.68 7.472 15.036 ;
  LAYER M4 ;
        RECT 7.42 15.016 7.46 15.056 ;
  LAYER M3 ;
        RECT 7.42 15.016 7.46 15.056 ;
  LAYER M2 ;
        RECT 7.424 15.02 7.456 15.052 ;
  LAYER M1 ;
        RECT 9.008 5.004 9.04 5.076 ;
  LAYER M2 ;
        RECT 8.988 5.024 9.06 5.056 ;
  LAYER M2 ;
        RECT 6.272 5.024 9.024 5.056 ;
  LAYER M1 ;
        RECT 6.256 5.004 6.288 5.076 ;
  LAYER M2 ;
        RECT 6.236 5.024 6.308 5.056 ;
  LAYER M1 ;
        RECT 9.008 8.112 9.04 8.184 ;
  LAYER M2 ;
        RECT 8.988 8.132 9.06 8.164 ;
  LAYER M2 ;
        RECT 6.272 8.132 9.024 8.164 ;
  LAYER M1 ;
        RECT 6.256 8.112 6.288 8.184 ;
  LAYER M2 ;
        RECT 6.236 8.132 6.308 8.164 ;
  LAYER M1 ;
        RECT 6.032 5.004 6.064 5.076 ;
  LAYER M2 ;
        RECT 6.012 5.024 6.084 5.056 ;
  LAYER M1 ;
        RECT 6.032 4.872 6.064 5.04 ;
  LAYER M1 ;
        RECT 6.032 4.836 6.064 4.908 ;
  LAYER M2 ;
        RECT 6.012 4.856 6.084 4.888 ;
  LAYER M2 ;
        RECT 6.048 4.856 6.272 4.888 ;
  LAYER M1 ;
        RECT 6.256 4.836 6.288 4.908 ;
  LAYER M2 ;
        RECT 6.236 4.856 6.308 4.888 ;
  LAYER M1 ;
        RECT 6.032 8.112 6.064 8.184 ;
  LAYER M2 ;
        RECT 6.012 8.132 6.084 8.164 ;
  LAYER M1 ;
        RECT 6.032 7.98 6.064 8.148 ;
  LAYER M1 ;
        RECT 6.032 7.944 6.064 8.016 ;
  LAYER M2 ;
        RECT 6.012 7.964 6.084 7.996 ;
  LAYER M2 ;
        RECT 6.048 7.964 6.272 7.996 ;
  LAYER M1 ;
        RECT 6.256 7.944 6.288 8.016 ;
  LAYER M2 ;
        RECT 6.236 7.964 6.308 7.996 ;
  LAYER M1 ;
        RECT 6.256 1.308 6.288 1.38 ;
  LAYER M2 ;
        RECT 6.236 1.328 6.308 1.36 ;
  LAYER M1 ;
        RECT 6.256 1.344 6.288 1.596 ;
  LAYER M1 ;
        RECT 6.256 1.596 6.288 8.148 ;
  LAYER M1 ;
        RECT 11.984 8.112 12.016 8.184 ;
  LAYER M2 ;
        RECT 11.964 8.132 12.036 8.164 ;
  LAYER M2 ;
        RECT 9.248 8.132 12 8.164 ;
  LAYER M1 ;
        RECT 9.232 8.112 9.264 8.184 ;
  LAYER M2 ;
        RECT 9.212 8.132 9.284 8.164 ;
  LAYER M1 ;
        RECT 11.984 5.004 12.016 5.076 ;
  LAYER M2 ;
        RECT 11.964 5.024 12.036 5.056 ;
  LAYER M2 ;
        RECT 9.248 5.024 12 5.056 ;
  LAYER M1 ;
        RECT 9.232 5.004 9.264 5.076 ;
  LAYER M2 ;
        RECT 9.212 5.024 9.284 5.056 ;
  LAYER M1 ;
        RECT 9.232 1.308 9.264 1.38 ;
  LAYER M2 ;
        RECT 9.212 1.328 9.284 1.36 ;
  LAYER M1 ;
        RECT 9.232 1.344 9.264 1.596 ;
  LAYER M1 ;
        RECT 9.232 1.596 9.264 8.148 ;
  LAYER M2 ;
        RECT 6.272 1.328 9.248 1.36 ;
  LAYER M1 ;
        RECT 3.056 1.896 3.088 1.968 ;
  LAYER M2 ;
        RECT 3.036 1.916 3.108 1.948 ;
  LAYER M1 ;
        RECT 3.056 1.764 3.088 1.932 ;
  LAYER M1 ;
        RECT 3.056 1.728 3.088 1.8 ;
  LAYER M2 ;
        RECT 3.036 1.748 3.108 1.78 ;
  LAYER M2 ;
        RECT 3.072 1.748 3.296 1.78 ;
  LAYER M1 ;
        RECT 3.28 1.728 3.312 1.8 ;
  LAYER M2 ;
        RECT 3.26 1.748 3.332 1.78 ;
  LAYER M1 ;
        RECT 3.056 5.004 3.088 5.076 ;
  LAYER M2 ;
        RECT 3.036 5.024 3.108 5.056 ;
  LAYER M1 ;
        RECT 3.056 4.872 3.088 5.04 ;
  LAYER M1 ;
        RECT 3.056 4.836 3.088 4.908 ;
  LAYER M2 ;
        RECT 3.036 4.856 3.108 4.888 ;
  LAYER M2 ;
        RECT 3.072 4.856 3.296 4.888 ;
  LAYER M1 ;
        RECT 3.28 4.836 3.312 4.908 ;
  LAYER M2 ;
        RECT 3.26 4.856 3.332 4.888 ;
  LAYER M1 ;
        RECT 3.056 8.112 3.088 8.184 ;
  LAYER M2 ;
        RECT 3.036 8.132 3.108 8.164 ;
  LAYER M1 ;
        RECT 3.056 7.98 3.088 8.148 ;
  LAYER M1 ;
        RECT 3.056 7.944 3.088 8.016 ;
  LAYER M2 ;
        RECT 3.036 7.964 3.108 7.996 ;
  LAYER M2 ;
        RECT 3.072 7.964 3.296 7.996 ;
  LAYER M1 ;
        RECT 3.28 7.944 3.312 8.016 ;
  LAYER M2 ;
        RECT 3.26 7.964 3.332 7.996 ;
  LAYER M1 ;
        RECT 3.056 11.22 3.088 11.292 ;
  LAYER M2 ;
        RECT 3.036 11.24 3.108 11.272 ;
  LAYER M1 ;
        RECT 3.056 11.088 3.088 11.256 ;
  LAYER M1 ;
        RECT 3.056 11.052 3.088 11.124 ;
  LAYER M2 ;
        RECT 3.036 11.072 3.108 11.104 ;
  LAYER M2 ;
        RECT 3.072 11.072 3.296 11.104 ;
  LAYER M1 ;
        RECT 3.28 11.052 3.312 11.124 ;
  LAYER M2 ;
        RECT 3.26 11.072 3.332 11.104 ;
  LAYER M1 ;
        RECT 6.032 1.896 6.064 1.968 ;
  LAYER M2 ;
        RECT 6.012 1.916 6.084 1.948 ;
  LAYER M2 ;
        RECT 3.296 1.916 6.048 1.948 ;
  LAYER M1 ;
        RECT 3.28 1.896 3.312 1.968 ;
  LAYER M2 ;
        RECT 3.26 1.916 3.332 1.948 ;
  LAYER M1 ;
        RECT 6.032 11.22 6.064 11.292 ;
  LAYER M2 ;
        RECT 6.012 11.24 6.084 11.272 ;
  LAYER M2 ;
        RECT 3.296 11.24 6.048 11.272 ;
  LAYER M1 ;
        RECT 3.28 11.22 3.312 11.292 ;
  LAYER M2 ;
        RECT 3.26 11.24 3.332 11.272 ;
  LAYER M1 ;
        RECT 3.28 1.14 3.312 1.212 ;
  LAYER M2 ;
        RECT 3.26 1.16 3.332 1.192 ;
  LAYER M1 ;
        RECT 3.28 1.176 3.312 1.596 ;
  LAYER M1 ;
        RECT 3.28 1.596 3.312 11.256 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 1.968 ;
  LAYER M2 ;
        RECT 11.964 1.916 12.036 1.948 ;
  LAYER M1 ;
        RECT 11.984 1.764 12.016 1.932 ;
  LAYER M1 ;
        RECT 11.984 1.728 12.016 1.8 ;
  LAYER M2 ;
        RECT 11.964 1.748 12.036 1.78 ;
  LAYER M2 ;
        RECT 12 1.748 12.224 1.78 ;
  LAYER M1 ;
        RECT 12.208 1.728 12.24 1.8 ;
  LAYER M2 ;
        RECT 12.188 1.748 12.26 1.78 ;
  LAYER M1 ;
        RECT 11.984 11.22 12.016 11.292 ;
  LAYER M2 ;
        RECT 11.964 11.24 12.036 11.272 ;
  LAYER M1 ;
        RECT 11.984 11.088 12.016 11.256 ;
  LAYER M1 ;
        RECT 11.984 11.052 12.016 11.124 ;
  LAYER M2 ;
        RECT 11.964 11.072 12.036 11.104 ;
  LAYER M2 ;
        RECT 12 11.072 12.224 11.104 ;
  LAYER M1 ;
        RECT 12.208 11.052 12.24 11.124 ;
  LAYER M2 ;
        RECT 12.188 11.072 12.26 11.104 ;
  LAYER M1 ;
        RECT 14.96 1.896 14.992 1.968 ;
  LAYER M2 ;
        RECT 14.94 1.916 15.012 1.948 ;
  LAYER M2 ;
        RECT 12.224 1.916 14.976 1.948 ;
  LAYER M1 ;
        RECT 12.208 1.896 12.24 1.968 ;
  LAYER M2 ;
        RECT 12.188 1.916 12.26 1.948 ;
  LAYER M1 ;
        RECT 14.96 5.004 14.992 5.076 ;
  LAYER M2 ;
        RECT 14.94 5.024 15.012 5.056 ;
  LAYER M2 ;
        RECT 12.224 5.024 14.976 5.056 ;
  LAYER M1 ;
        RECT 12.208 5.004 12.24 5.076 ;
  LAYER M2 ;
        RECT 12.188 5.024 12.26 5.056 ;
  LAYER M1 ;
        RECT 14.96 8.112 14.992 8.184 ;
  LAYER M2 ;
        RECT 14.94 8.132 15.012 8.164 ;
  LAYER M2 ;
        RECT 12.224 8.132 14.976 8.164 ;
  LAYER M1 ;
        RECT 12.208 8.112 12.24 8.184 ;
  LAYER M2 ;
        RECT 12.188 8.132 12.26 8.164 ;
  LAYER M1 ;
        RECT 14.96 11.22 14.992 11.292 ;
  LAYER M2 ;
        RECT 14.94 11.24 15.012 11.272 ;
  LAYER M2 ;
        RECT 12.224 11.24 14.976 11.272 ;
  LAYER M1 ;
        RECT 12.208 11.22 12.24 11.292 ;
  LAYER M2 ;
        RECT 12.188 11.24 12.26 11.272 ;
  LAYER M1 ;
        RECT 12.208 1.14 12.24 1.212 ;
  LAYER M2 ;
        RECT 12.188 1.16 12.26 1.192 ;
  LAYER M1 ;
        RECT 12.208 1.176 12.24 1.596 ;
  LAYER M1 ;
        RECT 12.208 1.596 12.24 11.256 ;
  LAYER M2 ;
        RECT 3.296 1.16 12.224 1.192 ;
  LAYER M1 ;
        RECT 9.008 11.22 9.04 11.292 ;
  LAYER M2 ;
        RECT 8.988 11.24 9.06 11.272 ;
  LAYER M2 ;
        RECT 6.048 11.24 9.024 11.272 ;
  LAYER M1 ;
        RECT 6.032 11.22 6.064 11.292 ;
  LAYER M2 ;
        RECT 6.012 11.24 6.084 11.272 ;
  LAYER M1 ;
        RECT 9.008 1.896 9.04 1.968 ;
  LAYER M2 ;
        RECT 8.988 1.916 9.06 1.948 ;
  LAYER M2 ;
        RECT 9.024 1.916 12 1.948 ;
  LAYER M1 ;
        RECT 11.984 1.896 12.016 1.968 ;
  LAYER M2 ;
        RECT 11.964 1.916 12.036 1.948 ;
  LAYER M1 ;
        RECT 6.64 7.44 6.672 7.512 ;
  LAYER M2 ;
        RECT 6.62 7.46 6.692 7.492 ;
  LAYER M2 ;
        RECT 6.432 7.46 6.656 7.492 ;
  LAYER M1 ;
        RECT 6.416 7.44 6.448 7.512 ;
  LAYER M2 ;
        RECT 6.396 7.46 6.468 7.492 ;
  LAYER M1 ;
        RECT 6.64 10.548 6.672 10.62 ;
  LAYER M2 ;
        RECT 6.62 10.568 6.692 10.6 ;
  LAYER M2 ;
        RECT 6.432 10.568 6.656 10.6 ;
  LAYER M1 ;
        RECT 6.416 10.548 6.448 10.62 ;
  LAYER M2 ;
        RECT 6.396 10.568 6.468 10.6 ;
  LAYER M1 ;
        RECT 3.664 7.44 3.696 7.512 ;
  LAYER M2 ;
        RECT 3.644 7.46 3.716 7.492 ;
  LAYER M1 ;
        RECT 3.68 7.46 6.432 7.492 ;
  LAYER M1 ;
        RECT 6.416 7.44 6.448 7.512 ;
  LAYER M2 ;
        RECT 6.396 7.46 6.468 7.492 ;
  LAYER M2 ;
        RECT 6.432 7.46 6.496 7.492 ;
  LAYER M1 ;
        RECT 6.48 7.44 6.512 7.512 ;
  LAYER M2 ;
        RECT 6.46 7.46 6.532 7.492 ;
  LAYER M1 ;
        RECT 3.664 10.548 3.696 10.62 ;
  LAYER M2 ;
        RECT 3.644 10.568 3.716 10.6 ;
  LAYER M1 ;
        RECT 3.68 10.568 6.432 10.6 ;
  LAYER M1 ;
        RECT 6.416 10.548 6.448 10.62 ;
  LAYER M2 ;
        RECT 6.396 10.568 6.468 10.6 ;
  LAYER M2 ;
        RECT 6.432 10.568 6.496 10.6 ;
  LAYER M1 ;
        RECT 6.48 10.548 6.512 10.62 ;
  LAYER M2 ;
        RECT 6.46 10.568 6.532 10.6 ;
  LAYER M1 ;
        RECT 6.48 14.244 6.512 14.316 ;
  LAYER M2 ;
        RECT 6.46 14.264 6.532 14.296 ;
  LAYER M1 ;
        RECT 6.48 14.028 6.512 14.28 ;
  LAYER M1 ;
        RECT 6.48 7.476 6.512 14.028 ;
  LAYER M1 ;
        RECT 9.616 10.548 9.648 10.62 ;
  LAYER M2 ;
        RECT 9.596 10.568 9.668 10.6 ;
  LAYER M2 ;
        RECT 9.408 10.568 9.632 10.6 ;
  LAYER M1 ;
        RECT 9.392 10.548 9.424 10.62 ;
  LAYER M2 ;
        RECT 9.372 10.568 9.444 10.6 ;
  LAYER M1 ;
        RECT 9.616 7.44 9.648 7.512 ;
  LAYER M2 ;
        RECT 9.596 7.46 9.668 7.492 ;
  LAYER M2 ;
        RECT 9.408 7.46 9.632 7.492 ;
  LAYER M1 ;
        RECT 9.392 7.44 9.424 7.512 ;
  LAYER M2 ;
        RECT 9.372 7.46 9.444 7.492 ;
  LAYER M1 ;
        RECT 9.392 14.244 9.424 14.316 ;
  LAYER M2 ;
        RECT 9.372 14.264 9.444 14.296 ;
  LAYER M1 ;
        RECT 9.392 14.028 9.424 14.28 ;
  LAYER M1 ;
        RECT 9.392 7.476 9.424 14.028 ;
  LAYER M2 ;
        RECT 6.496 14.264 9.408 14.296 ;
  LAYER M1 ;
        RECT 0.688 4.332 0.72 4.404 ;
  LAYER M2 ;
        RECT 0.668 4.352 0.74 4.384 ;
  LAYER M2 ;
        RECT 0.32 4.352 0.704 4.384 ;
  LAYER M1 ;
        RECT 0.304 4.332 0.336 4.404 ;
  LAYER M2 ;
        RECT 0.284 4.352 0.356 4.384 ;
  LAYER M1 ;
        RECT 0.688 7.44 0.72 7.512 ;
  LAYER M2 ;
        RECT 0.668 7.46 0.74 7.492 ;
  LAYER M2 ;
        RECT 0.32 7.46 0.704 7.492 ;
  LAYER M1 ;
        RECT 0.304 7.44 0.336 7.512 ;
  LAYER M2 ;
        RECT 0.284 7.46 0.356 7.492 ;
  LAYER M1 ;
        RECT 0.688 10.548 0.72 10.62 ;
  LAYER M2 ;
        RECT 0.668 10.568 0.74 10.6 ;
  LAYER M2 ;
        RECT 0.32 10.568 0.704 10.6 ;
  LAYER M1 ;
        RECT 0.304 10.548 0.336 10.62 ;
  LAYER M2 ;
        RECT 0.284 10.568 0.356 10.6 ;
  LAYER M1 ;
        RECT 0.688 13.656 0.72 13.728 ;
  LAYER M2 ;
        RECT 0.668 13.676 0.74 13.708 ;
  LAYER M2 ;
        RECT 0.32 13.676 0.704 13.708 ;
  LAYER M1 ;
        RECT 0.304 13.656 0.336 13.728 ;
  LAYER M2 ;
        RECT 0.284 13.676 0.356 13.708 ;
  LAYER M1 ;
        RECT 0.304 14.412 0.336 14.484 ;
  LAYER M2 ;
        RECT 0.284 14.432 0.356 14.464 ;
  LAYER M1 ;
        RECT 0.304 14.028 0.336 14.448 ;
  LAYER M1 ;
        RECT 0.304 4.368 0.336 14.028 ;
  LAYER M1 ;
        RECT 12.592 4.332 12.624 4.404 ;
  LAYER M2 ;
        RECT 12.572 4.352 12.644 4.384 ;
  LAYER M1 ;
        RECT 12.608 4.352 15.2 4.384 ;
  LAYER M1 ;
        RECT 15.184 4.332 15.216 4.404 ;
  LAYER M2 ;
        RECT 15.164 4.352 15.236 4.384 ;
  LAYER M2 ;
        RECT 15.2 4.352 15.264 4.384 ;
  LAYER M1 ;
        RECT 15.248 4.332 15.28 4.404 ;
  LAYER M2 ;
        RECT 15.228 4.352 15.3 4.384 ;
  LAYER M1 ;
        RECT 12.592 7.44 12.624 7.512 ;
  LAYER M2 ;
        RECT 12.572 7.46 12.644 7.492 ;
  LAYER M1 ;
        RECT 12.608 7.46 15.2 7.492 ;
  LAYER M1 ;
        RECT 15.184 7.44 15.216 7.512 ;
  LAYER M2 ;
        RECT 15.164 7.46 15.236 7.492 ;
  LAYER M2 ;
        RECT 15.2 7.46 15.264 7.492 ;
  LAYER M1 ;
        RECT 15.248 7.44 15.28 7.512 ;
  LAYER M2 ;
        RECT 15.228 7.46 15.3 7.492 ;
  LAYER M1 ;
        RECT 12.592 10.548 12.624 10.62 ;
  LAYER M2 ;
        RECT 12.572 10.568 12.644 10.6 ;
  LAYER M1 ;
        RECT 12.608 10.568 15.2 10.6 ;
  LAYER M1 ;
        RECT 15.184 10.548 15.216 10.62 ;
  LAYER M2 ;
        RECT 15.164 10.568 15.236 10.6 ;
  LAYER M2 ;
        RECT 15.2 10.568 15.264 10.6 ;
  LAYER M1 ;
        RECT 15.248 10.548 15.28 10.62 ;
  LAYER M2 ;
        RECT 15.228 10.568 15.3 10.6 ;
  LAYER M1 ;
        RECT 12.592 13.656 12.624 13.728 ;
  LAYER M2 ;
        RECT 12.572 13.676 12.644 13.708 ;
  LAYER M1 ;
        RECT 12.608 13.676 15.2 13.708 ;
  LAYER M1 ;
        RECT 15.184 13.656 15.216 13.728 ;
  LAYER M2 ;
        RECT 15.164 13.676 15.236 13.708 ;
  LAYER M2 ;
        RECT 15.2 13.676 15.264 13.708 ;
  LAYER M1 ;
        RECT 15.248 13.656 15.28 13.728 ;
  LAYER M2 ;
        RECT 15.228 13.676 15.3 13.708 ;
  LAYER M1 ;
        RECT 15.248 14.412 15.28 14.484 ;
  LAYER M2 ;
        RECT 15.228 14.432 15.3 14.464 ;
  LAYER M1 ;
        RECT 15.248 14.028 15.28 14.448 ;
  LAYER M1 ;
        RECT 15.248 4.536 15.28 14.028 ;
  LAYER M2 ;
        RECT 0.32 14.432 15.264 14.464 ;
  LAYER M1 ;
        RECT 3.664 4.332 3.696 4.404 ;
  LAYER M2 ;
        RECT 3.644 4.352 3.716 4.384 ;
  LAYER M2 ;
        RECT 0.704 4.352 3.68 4.384 ;
  LAYER M1 ;
        RECT 0.688 4.332 0.72 4.404 ;
  LAYER M2 ;
        RECT 0.668 4.352 0.74 4.384 ;
  LAYER M1 ;
        RECT 3.664 13.656 3.696 13.728 ;
  LAYER M2 ;
        RECT 3.644 13.676 3.716 13.708 ;
  LAYER M2 ;
        RECT 0.704 13.676 3.68 13.708 ;
  LAYER M1 ;
        RECT 0.688 13.656 0.72 13.728 ;
  LAYER M2 ;
        RECT 0.668 13.676 0.74 13.708 ;
  LAYER M1 ;
        RECT 6.64 13.656 6.672 13.728 ;
  LAYER M2 ;
        RECT 6.62 13.676 6.692 13.708 ;
  LAYER M2 ;
        RECT 3.68 13.676 6.656 13.708 ;
  LAYER M1 ;
        RECT 3.664 13.656 3.696 13.728 ;
  LAYER M2 ;
        RECT 3.644 13.676 3.716 13.708 ;
  LAYER M1 ;
        RECT 9.616 13.656 9.648 13.728 ;
  LAYER M2 ;
        RECT 9.596 13.676 9.668 13.708 ;
  LAYER M2 ;
        RECT 6.656 13.676 9.632 13.708 ;
  LAYER M1 ;
        RECT 6.64 13.656 6.672 13.728 ;
  LAYER M2 ;
        RECT 6.62 13.676 6.692 13.708 ;
  LAYER M1 ;
        RECT 9.616 4.332 9.648 4.404 ;
  LAYER M2 ;
        RECT 9.596 4.352 9.668 4.384 ;
  LAYER M2 ;
        RECT 9.632 4.352 12.608 4.384 ;
  LAYER M1 ;
        RECT 12.592 4.332 12.624 4.404 ;
  LAYER M2 ;
        RECT 12.572 4.352 12.644 4.384 ;
  LAYER M1 ;
        RECT 6.64 4.332 6.672 4.404 ;
  LAYER M2 ;
        RECT 6.62 4.352 6.692 4.384 ;
  LAYER M2 ;
        RECT 6.656 4.352 9.632 4.384 ;
  LAYER M1 ;
        RECT 9.616 4.332 9.648 4.404 ;
  LAYER M2 ;
        RECT 9.596 4.352 9.668 4.384 ;
  LAYER M1 ;
        RECT 0.64 1.848 3.136 4.452 ;
  LAYER M3 ;
        RECT 0.64 1.848 3.136 4.452 ;
  LAYER M2 ;
        RECT 0.64 1.848 3.136 4.452 ;
  LAYER M1 ;
        RECT 0.64 4.956 3.136 7.56 ;
  LAYER M3 ;
        RECT 0.64 4.956 3.136 7.56 ;
  LAYER M2 ;
        RECT 0.64 4.956 3.136 7.56 ;
  LAYER M1 ;
        RECT 0.64 8.064 3.136 10.668 ;
  LAYER M3 ;
        RECT 0.64 8.064 3.136 10.668 ;
  LAYER M2 ;
        RECT 0.64 8.064 3.136 10.668 ;
  LAYER M1 ;
        RECT 0.64 11.172 3.136 13.776 ;
  LAYER M3 ;
        RECT 0.64 11.172 3.136 13.776 ;
  LAYER M2 ;
        RECT 0.64 11.172 3.136 13.776 ;
  LAYER M1 ;
        RECT 3.616 1.848 6.112 4.452 ;
  LAYER M3 ;
        RECT 3.616 1.848 6.112 4.452 ;
  LAYER M2 ;
        RECT 3.616 1.848 6.112 4.452 ;
  LAYER M1 ;
        RECT 3.616 4.956 6.112 7.56 ;
  LAYER M3 ;
        RECT 3.616 4.956 6.112 7.56 ;
  LAYER M2 ;
        RECT 3.616 4.956 6.112 7.56 ;
  LAYER M1 ;
        RECT 3.616 8.064 6.112 10.668 ;
  LAYER M3 ;
        RECT 3.616 8.064 6.112 10.668 ;
  LAYER M2 ;
        RECT 3.616 8.064 6.112 10.668 ;
  LAYER M1 ;
        RECT 3.616 11.172 6.112 13.776 ;
  LAYER M3 ;
        RECT 3.616 11.172 6.112 13.776 ;
  LAYER M2 ;
        RECT 3.616 11.172 6.112 13.776 ;
  LAYER M1 ;
        RECT 6.592 1.848 9.088 4.452 ;
  LAYER M3 ;
        RECT 6.592 1.848 9.088 4.452 ;
  LAYER M2 ;
        RECT 6.592 1.848 9.088 4.452 ;
  LAYER M1 ;
        RECT 6.592 4.956 9.088 7.56 ;
  LAYER M3 ;
        RECT 6.592 4.956 9.088 7.56 ;
  LAYER M2 ;
        RECT 6.592 4.956 9.088 7.56 ;
  LAYER M1 ;
        RECT 6.592 8.064 9.088 10.668 ;
  LAYER M3 ;
        RECT 6.592 8.064 9.088 10.668 ;
  LAYER M2 ;
        RECT 6.592 8.064 9.088 10.668 ;
  LAYER M1 ;
        RECT 6.592 11.172 9.088 13.776 ;
  LAYER M3 ;
        RECT 6.592 11.172 9.088 13.776 ;
  LAYER M2 ;
        RECT 6.592 11.172 9.088 13.776 ;
  LAYER M1 ;
        RECT 9.568 1.848 12.064 4.452 ;
  LAYER M3 ;
        RECT 9.568 1.848 12.064 4.452 ;
  LAYER M2 ;
        RECT 9.568 1.848 12.064 4.452 ;
  LAYER M1 ;
        RECT 9.568 4.956 12.064 7.56 ;
  LAYER M3 ;
        RECT 9.568 4.956 12.064 7.56 ;
  LAYER M2 ;
        RECT 9.568 4.956 12.064 7.56 ;
  LAYER M1 ;
        RECT 9.568 8.064 12.064 10.668 ;
  LAYER M3 ;
        RECT 9.568 8.064 12.064 10.668 ;
  LAYER M2 ;
        RECT 9.568 8.064 12.064 10.668 ;
  LAYER M1 ;
        RECT 9.568 11.172 12.064 13.776 ;
  LAYER M3 ;
        RECT 9.568 11.172 12.064 13.776 ;
  LAYER M2 ;
        RECT 9.568 11.172 12.064 13.776 ;
  LAYER M1 ;
        RECT 12.544 1.848 15.04 4.452 ;
  LAYER M3 ;
        RECT 12.544 1.848 15.04 4.452 ;
  LAYER M2 ;
        RECT 12.544 1.848 15.04 4.452 ;
  LAYER M1 ;
        RECT 12.544 4.956 15.04 7.56 ;
  LAYER M3 ;
        RECT 12.544 4.956 15.04 7.56 ;
  LAYER M2 ;
        RECT 12.544 4.956 15.04 7.56 ;
  LAYER M1 ;
        RECT 12.544 8.064 15.04 10.668 ;
  LAYER M3 ;
        RECT 12.544 8.064 15.04 10.668 ;
  LAYER M2 ;
        RECT 12.544 8.064 15.04 10.668 ;
  LAYER M1 ;
        RECT 12.544 11.172 15.04 13.776 ;
  LAYER M3 ;
        RECT 12.544 11.172 15.04 13.776 ;
  LAYER M2 ;
        RECT 12.544 11.172 15.04 13.776 ;
  LAYER M1 ;
        RECT 5.344 0.216 5.376 0.876 ;
  LAYER M1 ;
        RECT 5.264 0.216 5.296 0.876 ;
  LAYER M1 ;
        RECT 5.424 0.656 5.456 0.688 ;
  LAYER M1 ;
        RECT 15.664 0.216 15.696 0.876 ;
  LAYER M1 ;
        RECT 15.744 0.216 15.776 0.876 ;
  LAYER M1 ;
        RECT 15.584 0.656 15.616 0.688 ;
  LAYER M1 ;
        RECT 6.704 0.3 6.736 0.96 ;
  LAYER M1 ;
        RECT 6.064 0.3 6.096 0.96 ;
  LAYER M1 ;
        RECT 6.784 0.3 6.816 0.96 ;
  LAYER M1 ;
        RECT 6.144 0.3 6.176 0.96 ;
  LAYER M1 ;
        RECT 6.624 0.3 6.656 0.96 ;
  LAYER M1 ;
        RECT 5.984 0.488 6.016 0.52 ;
  LAYER M1 ;
        RECT 8.064 0.3 8.096 0.96 ;
  LAYER M1 ;
        RECT 7.424 0.3 7.456 0.96 ;
  LAYER M1 ;
        RECT 8.144 0.3 8.176 0.96 ;
  LAYER M1 ;
        RECT 7.504 0.3 7.536 0.96 ;
  LAYER M1 ;
        RECT 7.984 0.3 8.016 0.96 ;
  LAYER M1 ;
        RECT 7.344 0.488 7.376 0.52 ;
  LAYER M1 ;
        RECT 6.56 24.24 6.592 24.312 ;
  LAYER M2 ;
        RECT 6.54 24.26 6.612 24.292 ;
  LAYER M2 ;
        RECT 6.576 24.26 9.328 24.292 ;
  LAYER M1 ;
        RECT 9.312 24.24 9.344 24.312 ;
  LAYER M2 ;
        RECT 9.292 24.26 9.364 24.292 ;
  LAYER M1 ;
        RECT 9.536 21.132 9.568 21.204 ;
  LAYER M2 ;
        RECT 9.516 21.152 9.588 21.184 ;
  LAYER M1 ;
        RECT 9.536 21.168 9.568 21.336 ;
  LAYER M1 ;
        RECT 9.536 21.3 9.568 21.372 ;
  LAYER M2 ;
        RECT 9.516 21.32 9.588 21.352 ;
  LAYER M2 ;
        RECT 9.328 21.32 9.552 21.352 ;
  LAYER M1 ;
        RECT 9.312 21.3 9.344 21.372 ;
  LAYER M2 ;
        RECT 9.292 21.32 9.364 21.352 ;
  LAYER M1 ;
        RECT 9.312 31.044 9.344 31.116 ;
  LAYER M2 ;
        RECT 9.292 31.064 9.364 31.096 ;
  LAYER M1 ;
        RECT 9.312 30.828 9.344 31.08 ;
  LAYER M1 ;
        RECT 9.312 21.336 9.344 30.828 ;
  LAYER M1 ;
        RECT 3.584 27.348 3.616 27.42 ;
  LAYER M2 ;
        RECT 3.564 27.368 3.636 27.4 ;
  LAYER M2 ;
        RECT 3.6 27.368 6.352 27.4 ;
  LAYER M1 ;
        RECT 6.336 27.348 6.368 27.42 ;
  LAYER M2 ;
        RECT 6.316 27.368 6.388 27.4 ;
  LAYER M1 ;
        RECT 6.336 31.044 6.368 31.116 ;
  LAYER M2 ;
        RECT 6.316 31.064 6.388 31.096 ;
  LAYER M1 ;
        RECT 6.336 30.828 6.368 31.08 ;
  LAYER M1 ;
        RECT 6.336 27.384 6.368 30.828 ;
  LAYER M2 ;
        RECT 6.352 31.064 9.328 31.096 ;
  LAYER M1 ;
        RECT 9.536 24.24 9.568 24.312 ;
  LAYER M2 ;
        RECT 9.516 24.26 9.588 24.292 ;
  LAYER M2 ;
        RECT 9.552 24.26 12.304 24.292 ;
  LAYER M1 ;
        RECT 12.288 24.24 12.32 24.312 ;
  LAYER M2 ;
        RECT 12.268 24.26 12.34 24.292 ;
  LAYER M1 ;
        RECT 9.536 27.348 9.568 27.42 ;
  LAYER M2 ;
        RECT 9.516 27.368 9.588 27.4 ;
  LAYER M2 ;
        RECT 9.552 27.368 12.304 27.4 ;
  LAYER M1 ;
        RECT 12.288 27.348 12.32 27.42 ;
  LAYER M2 ;
        RECT 12.268 27.368 12.34 27.4 ;
  LAYER M1 ;
        RECT 12.288 31.212 12.32 31.284 ;
  LAYER M2 ;
        RECT 12.268 31.232 12.34 31.264 ;
  LAYER M1 ;
        RECT 12.288 30.828 12.32 31.248 ;
  LAYER M1 ;
        RECT 12.288 24.276 12.32 30.828 ;
  LAYER M1 ;
        RECT 3.584 24.24 3.616 24.312 ;
  LAYER M2 ;
        RECT 3.564 24.26 3.636 24.292 ;
  LAYER M1 ;
        RECT 3.584 24.276 3.616 24.444 ;
  LAYER M1 ;
        RECT 3.584 24.408 3.616 24.48 ;
  LAYER M2 ;
        RECT 3.564 24.428 3.636 24.46 ;
  LAYER M2 ;
        RECT 3.376 24.428 3.6 24.46 ;
  LAYER M1 ;
        RECT 3.36 24.408 3.392 24.48 ;
  LAYER M2 ;
        RECT 3.34 24.428 3.412 24.46 ;
  LAYER M1 ;
        RECT 3.584 21.132 3.616 21.204 ;
  LAYER M2 ;
        RECT 3.564 21.152 3.636 21.184 ;
  LAYER M1 ;
        RECT 3.584 21.168 3.616 21.336 ;
  LAYER M1 ;
        RECT 3.584 21.3 3.616 21.372 ;
  LAYER M2 ;
        RECT 3.564 21.32 3.636 21.352 ;
  LAYER M2 ;
        RECT 3.376 21.32 3.6 21.352 ;
  LAYER M1 ;
        RECT 3.36 21.3 3.392 21.372 ;
  LAYER M2 ;
        RECT 3.34 21.32 3.412 21.352 ;
  LAYER M1 ;
        RECT 3.36 31.212 3.392 31.284 ;
  LAYER M2 ;
        RECT 3.34 31.232 3.412 31.264 ;
  LAYER M1 ;
        RECT 3.36 30.828 3.392 31.248 ;
  LAYER M1 ;
        RECT 3.36 21.336 3.392 30.828 ;
  LAYER M2 ;
        RECT 3.376 31.232 12.304 31.264 ;
  LAYER M1 ;
        RECT 6.56 27.348 6.592 27.42 ;
  LAYER M2 ;
        RECT 6.54 27.368 6.612 27.4 ;
  LAYER M2 ;
        RECT 6.576 27.368 9.552 27.4 ;
  LAYER M1 ;
        RECT 9.536 27.348 9.568 27.42 ;
  LAYER M2 ;
        RECT 9.516 27.368 9.588 27.4 ;
  LAYER M1 ;
        RECT 6.56 21.132 6.592 21.204 ;
  LAYER M2 ;
        RECT 6.54 21.152 6.612 21.184 ;
  LAYER M2 ;
        RECT 3.6 21.152 6.576 21.184 ;
  LAYER M1 ;
        RECT 3.584 21.132 3.616 21.204 ;
  LAYER M2 ;
        RECT 3.564 21.152 3.636 21.184 ;
  LAYER M1 ;
        RECT 12.512 30.456 12.544 30.528 ;
  LAYER M2 ;
        RECT 12.492 30.476 12.564 30.508 ;
  LAYER M2 ;
        RECT 12.528 30.476 15.28 30.508 ;
  LAYER M1 ;
        RECT 15.264 30.456 15.296 30.528 ;
  LAYER M2 ;
        RECT 15.244 30.476 15.316 30.508 ;
  LAYER M1 ;
        RECT 12.512 27.348 12.544 27.42 ;
  LAYER M2 ;
        RECT 12.492 27.368 12.564 27.4 ;
  LAYER M2 ;
        RECT 12.528 27.368 15.28 27.4 ;
  LAYER M1 ;
        RECT 15.264 27.348 15.296 27.42 ;
  LAYER M2 ;
        RECT 15.244 27.368 15.316 27.4 ;
  LAYER M1 ;
        RECT 12.512 24.24 12.544 24.312 ;
  LAYER M2 ;
        RECT 12.492 24.26 12.564 24.292 ;
  LAYER M2 ;
        RECT 12.528 24.26 15.28 24.292 ;
  LAYER M1 ;
        RECT 15.264 24.24 15.296 24.312 ;
  LAYER M2 ;
        RECT 15.244 24.26 15.316 24.292 ;
  LAYER M1 ;
        RECT 12.512 21.132 12.544 21.204 ;
  LAYER M2 ;
        RECT 12.492 21.152 12.564 21.184 ;
  LAYER M2 ;
        RECT 12.528 21.152 15.28 21.184 ;
  LAYER M1 ;
        RECT 15.264 21.132 15.296 21.204 ;
  LAYER M2 ;
        RECT 15.244 21.152 15.316 21.184 ;
  LAYER M1 ;
        RECT 12.512 18.024 12.544 18.096 ;
  LAYER M2 ;
        RECT 12.492 18.044 12.564 18.076 ;
  LAYER M2 ;
        RECT 12.528 18.044 15.28 18.076 ;
  LAYER M1 ;
        RECT 15.264 18.024 15.296 18.096 ;
  LAYER M2 ;
        RECT 15.244 18.044 15.316 18.076 ;
  LAYER M1 ;
        RECT 15.264 31.38 15.296 31.452 ;
  LAYER M2 ;
        RECT 15.244 31.4 15.316 31.432 ;
  LAYER M1 ;
        RECT 15.264 30.828 15.296 31.416 ;
  LAYER M1 ;
        RECT 15.264 18.06 15.296 30.828 ;
  LAYER M1 ;
        RECT 0.608 30.456 0.64 30.528 ;
  LAYER M2 ;
        RECT 0.588 30.476 0.66 30.508 ;
  LAYER M1 ;
        RECT 0.608 30.492 0.64 30.66 ;
  LAYER M1 ;
        RECT 0.608 30.624 0.64 30.696 ;
  LAYER M2 ;
        RECT 0.588 30.644 0.66 30.676 ;
  LAYER M2 ;
        RECT 0.4 30.644 0.624 30.676 ;
  LAYER M1 ;
        RECT 0.384 30.624 0.416 30.696 ;
  LAYER M2 ;
        RECT 0.364 30.644 0.436 30.676 ;
  LAYER M1 ;
        RECT 0.608 27.348 0.64 27.42 ;
  LAYER M2 ;
        RECT 0.588 27.368 0.66 27.4 ;
  LAYER M1 ;
        RECT 0.608 27.384 0.64 27.552 ;
  LAYER M1 ;
        RECT 0.608 27.516 0.64 27.588 ;
  LAYER M2 ;
        RECT 0.588 27.536 0.66 27.568 ;
  LAYER M2 ;
        RECT 0.4 27.536 0.624 27.568 ;
  LAYER M1 ;
        RECT 0.384 27.516 0.416 27.588 ;
  LAYER M2 ;
        RECT 0.364 27.536 0.436 27.568 ;
  LAYER M1 ;
        RECT 0.608 24.24 0.64 24.312 ;
  LAYER M2 ;
        RECT 0.588 24.26 0.66 24.292 ;
  LAYER M1 ;
        RECT 0.608 24.276 0.64 24.444 ;
  LAYER M1 ;
        RECT 0.608 24.408 0.64 24.48 ;
  LAYER M2 ;
        RECT 0.588 24.428 0.66 24.46 ;
  LAYER M2 ;
        RECT 0.4 24.428 0.624 24.46 ;
  LAYER M1 ;
        RECT 0.384 24.408 0.416 24.48 ;
  LAYER M2 ;
        RECT 0.364 24.428 0.436 24.46 ;
  LAYER M1 ;
        RECT 0.608 21.132 0.64 21.204 ;
  LAYER M2 ;
        RECT 0.588 21.152 0.66 21.184 ;
  LAYER M1 ;
        RECT 0.608 21.168 0.64 21.336 ;
  LAYER M1 ;
        RECT 0.608 21.3 0.64 21.372 ;
  LAYER M2 ;
        RECT 0.588 21.32 0.66 21.352 ;
  LAYER M2 ;
        RECT 0.4 21.32 0.624 21.352 ;
  LAYER M1 ;
        RECT 0.384 21.3 0.416 21.372 ;
  LAYER M2 ;
        RECT 0.364 21.32 0.436 21.352 ;
  LAYER M1 ;
        RECT 0.608 18.024 0.64 18.096 ;
  LAYER M2 ;
        RECT 0.588 18.044 0.66 18.076 ;
  LAYER M1 ;
        RECT 0.608 18.06 0.64 18.228 ;
  LAYER M1 ;
        RECT 0.608 18.192 0.64 18.264 ;
  LAYER M2 ;
        RECT 0.588 18.212 0.66 18.244 ;
  LAYER M2 ;
        RECT 0.4 18.212 0.624 18.244 ;
  LAYER M1 ;
        RECT 0.384 18.192 0.416 18.264 ;
  LAYER M2 ;
        RECT 0.364 18.212 0.436 18.244 ;
  LAYER M1 ;
        RECT 0.384 31.38 0.416 31.452 ;
  LAYER M2 ;
        RECT 0.364 31.4 0.436 31.432 ;
  LAYER M1 ;
        RECT 0.384 30.828 0.416 31.416 ;
  LAYER M1 ;
        RECT 0.384 18.228 0.416 30.828 ;
  LAYER M2 ;
        RECT 0.4 31.4 15.28 31.432 ;
  LAYER M1 ;
        RECT 9.536 30.456 9.568 30.528 ;
  LAYER M2 ;
        RECT 9.516 30.476 9.588 30.508 ;
  LAYER M2 ;
        RECT 9.552 30.476 12.528 30.508 ;
  LAYER M1 ;
        RECT 12.512 30.456 12.544 30.528 ;
  LAYER M2 ;
        RECT 12.492 30.476 12.564 30.508 ;
  LAYER M1 ;
        RECT 9.536 18.024 9.568 18.096 ;
  LAYER M2 ;
        RECT 9.516 18.044 9.588 18.076 ;
  LAYER M2 ;
        RECT 9.552 18.044 12.528 18.076 ;
  LAYER M1 ;
        RECT 12.512 18.024 12.544 18.096 ;
  LAYER M2 ;
        RECT 12.492 18.044 12.564 18.076 ;
  LAYER M1 ;
        RECT 6.56 18.024 6.592 18.096 ;
  LAYER M2 ;
        RECT 6.54 18.044 6.612 18.076 ;
  LAYER M2 ;
        RECT 6.576 18.044 9.552 18.076 ;
  LAYER M1 ;
        RECT 9.536 18.024 9.568 18.096 ;
  LAYER M2 ;
        RECT 9.516 18.044 9.588 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M2 ;
        RECT 3.6 18.044 6.576 18.076 ;
  LAYER M1 ;
        RECT 6.56 18.024 6.592 18.096 ;
  LAYER M2 ;
        RECT 6.54 18.044 6.612 18.076 ;
  LAYER M1 ;
        RECT 3.584 30.456 3.616 30.528 ;
  LAYER M2 ;
        RECT 3.564 30.476 3.636 30.508 ;
  LAYER M2 ;
        RECT 0.624 30.476 3.6 30.508 ;
  LAYER M1 ;
        RECT 0.608 30.456 0.64 30.528 ;
  LAYER M2 ;
        RECT 0.588 30.476 0.66 30.508 ;
  LAYER M1 ;
        RECT 6.56 30.456 6.592 30.528 ;
  LAYER M2 ;
        RECT 6.54 30.476 6.612 30.508 ;
  LAYER M2 ;
        RECT 3.6 30.476 6.576 30.508 ;
  LAYER M1 ;
        RECT 3.584 30.456 3.616 30.528 ;
  LAYER M2 ;
        RECT 3.564 30.476 3.636 30.508 ;
  LAYER M1 ;
        RECT 8.928 21.804 8.96 21.876 ;
  LAYER M2 ;
        RECT 8.908 21.824 8.98 21.856 ;
  LAYER M2 ;
        RECT 8.944 21.824 9.168 21.856 ;
  LAYER M1 ;
        RECT 9.152 21.804 9.184 21.876 ;
  LAYER M2 ;
        RECT 9.132 21.824 9.204 21.856 ;
  LAYER M1 ;
        RECT 11.904 18.696 11.936 18.768 ;
  LAYER M2 ;
        RECT 11.884 18.716 11.956 18.748 ;
  LAYER M1 ;
        RECT 9.168 18.716 11.92 18.748 ;
  LAYER M1 ;
        RECT 9.152 18.696 9.184 18.768 ;
  LAYER M2 ;
        RECT 9.132 18.716 9.204 18.748 ;
  LAYER M2 ;
        RECT 9.104 18.716 9.168 18.748 ;
  LAYER M1 ;
        RECT 9.088 18.696 9.12 18.768 ;
  LAYER M2 ;
        RECT 9.068 18.716 9.14 18.748 ;
  LAYER M1 ;
        RECT 9.088 15 9.12 15.072 ;
  LAYER M2 ;
        RECT 9.068 15.02 9.14 15.052 ;
  LAYER M1 ;
        RECT 9.088 15.036 9.12 15.288 ;
  LAYER M1 ;
        RECT 9.088 15.288 9.12 21.84 ;
  LAYER M1 ;
        RECT 5.952 24.912 5.984 24.984 ;
  LAYER M2 ;
        RECT 5.932 24.932 6.004 24.964 ;
  LAYER M2 ;
        RECT 5.968 24.932 6.192 24.964 ;
  LAYER M1 ;
        RECT 6.176 24.912 6.208 24.984 ;
  LAYER M2 ;
        RECT 6.156 24.932 6.228 24.964 ;
  LAYER M1 ;
        RECT 6.176 15 6.208 15.072 ;
  LAYER M2 ;
        RECT 6.156 15.02 6.228 15.052 ;
  LAYER M1 ;
        RECT 6.176 15.036 6.208 15.288 ;
  LAYER M1 ;
        RECT 6.176 15.288 6.208 24.948 ;
  LAYER M2 ;
        RECT 6.192 15.02 9.104 15.052 ;
  LAYER M1 ;
        RECT 11.904 21.804 11.936 21.876 ;
  LAYER M2 ;
        RECT 11.884 21.824 11.956 21.856 ;
  LAYER M2 ;
        RECT 11.92 21.824 12.144 21.856 ;
  LAYER M1 ;
        RECT 12.128 21.804 12.16 21.876 ;
  LAYER M2 ;
        RECT 12.108 21.824 12.18 21.856 ;
  LAYER M1 ;
        RECT 11.904 24.912 11.936 24.984 ;
  LAYER M2 ;
        RECT 11.884 24.932 11.956 24.964 ;
  LAYER M2 ;
        RECT 11.92 24.932 12.144 24.964 ;
  LAYER M1 ;
        RECT 12.128 24.912 12.16 24.984 ;
  LAYER M2 ;
        RECT 12.108 24.932 12.18 24.964 ;
  LAYER M1 ;
        RECT 12.128 14.832 12.16 14.904 ;
  LAYER M2 ;
        RECT 12.108 14.852 12.18 14.884 ;
  LAYER M1 ;
        RECT 12.128 14.868 12.16 15.288 ;
  LAYER M1 ;
        RECT 12.128 15.288 12.16 24.948 ;
  LAYER M1 ;
        RECT 5.952 21.804 5.984 21.876 ;
  LAYER M2 ;
        RECT 5.932 21.824 6.004 21.856 ;
  LAYER M1 ;
        RECT 3.216 21.824 5.968 21.856 ;
  LAYER M1 ;
        RECT 3.2 21.804 3.232 21.876 ;
  LAYER M2 ;
        RECT 3.18 21.824 3.252 21.856 ;
  LAYER M2 ;
        RECT 3.152 21.824 3.216 21.856 ;
  LAYER M1 ;
        RECT 3.136 21.804 3.168 21.876 ;
  LAYER M2 ;
        RECT 3.116 21.824 3.188 21.856 ;
  LAYER M1 ;
        RECT 5.952 18.696 5.984 18.768 ;
  LAYER M2 ;
        RECT 5.932 18.716 6.004 18.748 ;
  LAYER M1 ;
        RECT 3.216 18.716 5.968 18.748 ;
  LAYER M1 ;
        RECT 3.2 18.696 3.232 18.768 ;
  LAYER M2 ;
        RECT 3.18 18.716 3.252 18.748 ;
  LAYER M2 ;
        RECT 3.152 18.716 3.216 18.748 ;
  LAYER M1 ;
        RECT 3.136 18.696 3.168 18.768 ;
  LAYER M2 ;
        RECT 3.116 18.716 3.188 18.748 ;
  LAYER M1 ;
        RECT 3.136 14.832 3.168 14.904 ;
  LAYER M2 ;
        RECT 3.116 14.852 3.188 14.884 ;
  LAYER M1 ;
        RECT 3.136 14.868 3.168 15.288 ;
  LAYER M1 ;
        RECT 3.136 15.288 3.168 21.672 ;
  LAYER M2 ;
        RECT 3.152 14.852 12.144 14.884 ;
  LAYER M1 ;
        RECT 8.928 24.912 8.96 24.984 ;
  LAYER M2 ;
        RECT 8.908 24.932 8.98 24.964 ;
  LAYER M2 ;
        RECT 8.944 24.932 11.92 24.964 ;
  LAYER M1 ;
        RECT 11.904 24.912 11.936 24.984 ;
  LAYER M2 ;
        RECT 11.884 24.932 11.956 24.964 ;
  LAYER M1 ;
        RECT 8.928 18.696 8.96 18.768 ;
  LAYER M2 ;
        RECT 8.908 18.716 8.98 18.748 ;
  LAYER M2 ;
        RECT 5.968 18.716 8.944 18.748 ;
  LAYER M1 ;
        RECT 5.952 18.696 5.984 18.768 ;
  LAYER M2 ;
        RECT 5.932 18.716 6.004 18.748 ;
  LAYER M1 ;
        RECT 14.88 28.02 14.912 28.092 ;
  LAYER M2 ;
        RECT 14.86 28.04 14.932 28.072 ;
  LAYER M2 ;
        RECT 14.896 28.04 15.12 28.072 ;
  LAYER M1 ;
        RECT 15.104 28.02 15.136 28.092 ;
  LAYER M2 ;
        RECT 15.084 28.04 15.156 28.072 ;
  LAYER M1 ;
        RECT 14.88 24.912 14.912 24.984 ;
  LAYER M2 ;
        RECT 14.86 24.932 14.932 24.964 ;
  LAYER M2 ;
        RECT 14.896 24.932 15.12 24.964 ;
  LAYER M1 ;
        RECT 15.104 24.912 15.136 24.984 ;
  LAYER M2 ;
        RECT 15.084 24.932 15.156 24.964 ;
  LAYER M1 ;
        RECT 14.88 21.804 14.912 21.876 ;
  LAYER M2 ;
        RECT 14.86 21.824 14.932 21.856 ;
  LAYER M2 ;
        RECT 14.896 21.824 15.12 21.856 ;
  LAYER M1 ;
        RECT 15.104 21.804 15.136 21.876 ;
  LAYER M2 ;
        RECT 15.084 21.824 15.156 21.856 ;
  LAYER M1 ;
        RECT 14.88 18.696 14.912 18.768 ;
  LAYER M2 ;
        RECT 14.86 18.716 14.932 18.748 ;
  LAYER M2 ;
        RECT 14.896 18.716 15.12 18.748 ;
  LAYER M1 ;
        RECT 15.104 18.696 15.136 18.768 ;
  LAYER M2 ;
        RECT 15.084 18.716 15.156 18.748 ;
  LAYER M1 ;
        RECT 14.88 15.588 14.912 15.66 ;
  LAYER M2 ;
        RECT 14.86 15.608 14.932 15.64 ;
  LAYER M2 ;
        RECT 14.896 15.608 15.12 15.64 ;
  LAYER M1 ;
        RECT 15.104 15.588 15.136 15.66 ;
  LAYER M2 ;
        RECT 15.084 15.608 15.156 15.64 ;
  LAYER M1 ;
        RECT 15.104 14.664 15.136 14.736 ;
  LAYER M2 ;
        RECT 15.084 14.684 15.156 14.716 ;
  LAYER M1 ;
        RECT 15.104 14.7 15.136 15.288 ;
  LAYER M1 ;
        RECT 15.104 15.288 15.136 28.056 ;
  LAYER M1 ;
        RECT 2.976 28.02 3.008 28.092 ;
  LAYER M2 ;
        RECT 2.956 28.04 3.028 28.072 ;
  LAYER M1 ;
        RECT 0.24 28.04 2.992 28.072 ;
  LAYER M1 ;
        RECT 0.224 28.02 0.256 28.092 ;
  LAYER M2 ;
        RECT 0.204 28.04 0.276 28.072 ;
  LAYER M2 ;
        RECT 0.176 28.04 0.24 28.072 ;
  LAYER M1 ;
        RECT 0.16 28.02 0.192 28.092 ;
  LAYER M2 ;
        RECT 0.14 28.04 0.212 28.072 ;
  LAYER M1 ;
        RECT 2.976 24.912 3.008 24.984 ;
  LAYER M2 ;
        RECT 2.956 24.932 3.028 24.964 ;
  LAYER M1 ;
        RECT 0.24 24.932 2.992 24.964 ;
  LAYER M1 ;
        RECT 0.224 24.912 0.256 24.984 ;
  LAYER M2 ;
        RECT 0.204 24.932 0.276 24.964 ;
  LAYER M2 ;
        RECT 0.176 24.932 0.24 24.964 ;
  LAYER M1 ;
        RECT 0.16 24.912 0.192 24.984 ;
  LAYER M2 ;
        RECT 0.14 24.932 0.212 24.964 ;
  LAYER M1 ;
        RECT 2.976 21.804 3.008 21.876 ;
  LAYER M2 ;
        RECT 2.956 21.824 3.028 21.856 ;
  LAYER M1 ;
        RECT 0.24 21.824 2.992 21.856 ;
  LAYER M1 ;
        RECT 0.224 21.804 0.256 21.876 ;
  LAYER M2 ;
        RECT 0.204 21.824 0.276 21.856 ;
  LAYER M2 ;
        RECT 0.176 21.824 0.24 21.856 ;
  LAYER M1 ;
        RECT 0.16 21.804 0.192 21.876 ;
  LAYER M2 ;
        RECT 0.14 21.824 0.212 21.856 ;
  LAYER M1 ;
        RECT 2.976 18.696 3.008 18.768 ;
  LAYER M2 ;
        RECT 2.956 18.716 3.028 18.748 ;
  LAYER M1 ;
        RECT 0.24 18.716 2.992 18.748 ;
  LAYER M1 ;
        RECT 0.224 18.696 0.256 18.768 ;
  LAYER M2 ;
        RECT 0.204 18.716 0.276 18.748 ;
  LAYER M2 ;
        RECT 0.176 18.716 0.24 18.748 ;
  LAYER M1 ;
        RECT 0.16 18.696 0.192 18.768 ;
  LAYER M2 ;
        RECT 0.14 18.716 0.212 18.748 ;
  LAYER M1 ;
        RECT 2.976 15.588 3.008 15.66 ;
  LAYER M2 ;
        RECT 2.956 15.608 3.028 15.64 ;
  LAYER M1 ;
        RECT 0.24 15.608 2.992 15.64 ;
  LAYER M1 ;
        RECT 0.224 15.588 0.256 15.66 ;
  LAYER M2 ;
        RECT 0.204 15.608 0.276 15.64 ;
  LAYER M2 ;
        RECT 0.176 15.608 0.24 15.64 ;
  LAYER M1 ;
        RECT 0.16 15.588 0.192 15.66 ;
  LAYER M2 ;
        RECT 0.14 15.608 0.212 15.64 ;
  LAYER M1 ;
        RECT 0.16 14.664 0.192 14.736 ;
  LAYER M2 ;
        RECT 0.14 14.684 0.212 14.716 ;
  LAYER M1 ;
        RECT 0.16 14.7 0.192 15.288 ;
  LAYER M1 ;
        RECT 0.16 15.288 0.192 27.888 ;
  LAYER M2 ;
        RECT 0.176 14.684 15.12 14.716 ;
  LAYER M1 ;
        RECT 11.904 28.02 11.936 28.092 ;
  LAYER M2 ;
        RECT 11.884 28.04 11.956 28.072 ;
  LAYER M2 ;
        RECT 11.92 28.04 14.896 28.072 ;
  LAYER M1 ;
        RECT 14.88 28.02 14.912 28.092 ;
  LAYER M2 ;
        RECT 14.86 28.04 14.932 28.072 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 15.66 ;
  LAYER M2 ;
        RECT 11.884 15.608 11.956 15.64 ;
  LAYER M2 ;
        RECT 11.92 15.608 14.896 15.64 ;
  LAYER M1 ;
        RECT 14.88 15.588 14.912 15.66 ;
  LAYER M2 ;
        RECT 14.86 15.608 14.932 15.64 ;
  LAYER M1 ;
        RECT 8.928 15.588 8.96 15.66 ;
  LAYER M2 ;
        RECT 8.908 15.608 8.98 15.64 ;
  LAYER M2 ;
        RECT 8.944 15.608 11.92 15.64 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 15.66 ;
  LAYER M2 ;
        RECT 11.884 15.608 11.956 15.64 ;
  LAYER M1 ;
        RECT 5.952 15.588 5.984 15.66 ;
  LAYER M2 ;
        RECT 5.932 15.608 6.004 15.64 ;
  LAYER M2 ;
        RECT 5.968 15.608 8.944 15.64 ;
  LAYER M1 ;
        RECT 8.928 15.588 8.96 15.66 ;
  LAYER M2 ;
        RECT 8.908 15.608 8.98 15.64 ;
  LAYER M1 ;
        RECT 5.952 28.02 5.984 28.092 ;
  LAYER M2 ;
        RECT 5.932 28.04 6.004 28.072 ;
  LAYER M2 ;
        RECT 2.992 28.04 5.968 28.072 ;
  LAYER M1 ;
        RECT 2.976 28.02 3.008 28.092 ;
  LAYER M2 ;
        RECT 2.956 28.04 3.028 28.072 ;
  LAYER M1 ;
        RECT 8.928 28.02 8.96 28.092 ;
  LAYER M2 ;
        RECT 8.908 28.04 8.98 28.072 ;
  LAYER M2 ;
        RECT 5.968 28.04 8.944 28.072 ;
  LAYER M1 ;
        RECT 5.952 28.02 5.984 28.092 ;
  LAYER M2 ;
        RECT 5.932 28.04 6.004 28.072 ;
  LAYER M1 ;
        RECT 12.464 27.972 14.96 30.576 ;
  LAYER M3 ;
        RECT 12.464 27.972 14.96 30.576 ;
  LAYER M2 ;
        RECT 12.464 27.972 14.96 30.576 ;
  LAYER M1 ;
        RECT 12.464 24.864 14.96 27.468 ;
  LAYER M3 ;
        RECT 12.464 24.864 14.96 27.468 ;
  LAYER M2 ;
        RECT 12.464 24.864 14.96 27.468 ;
  LAYER M1 ;
        RECT 12.464 21.756 14.96 24.36 ;
  LAYER M3 ;
        RECT 12.464 21.756 14.96 24.36 ;
  LAYER M2 ;
        RECT 12.464 21.756 14.96 24.36 ;
  LAYER M1 ;
        RECT 12.464 18.648 14.96 21.252 ;
  LAYER M3 ;
        RECT 12.464 18.648 14.96 21.252 ;
  LAYER M2 ;
        RECT 12.464 18.648 14.96 21.252 ;
  LAYER M1 ;
        RECT 12.464 15.54 14.96 18.144 ;
  LAYER M3 ;
        RECT 12.464 15.54 14.96 18.144 ;
  LAYER M2 ;
        RECT 12.464 15.54 14.96 18.144 ;
  LAYER M1 ;
        RECT 9.488 27.972 11.984 30.576 ;
  LAYER M3 ;
        RECT 9.488 27.972 11.984 30.576 ;
  LAYER M2 ;
        RECT 9.488 27.972 11.984 30.576 ;
  LAYER M1 ;
        RECT 9.488 24.864 11.984 27.468 ;
  LAYER M3 ;
        RECT 9.488 24.864 11.984 27.468 ;
  LAYER M2 ;
        RECT 9.488 24.864 11.984 27.468 ;
  LAYER M1 ;
        RECT 9.488 21.756 11.984 24.36 ;
  LAYER M3 ;
        RECT 9.488 21.756 11.984 24.36 ;
  LAYER M2 ;
        RECT 9.488 21.756 11.984 24.36 ;
  LAYER M1 ;
        RECT 9.488 18.648 11.984 21.252 ;
  LAYER M3 ;
        RECT 9.488 18.648 11.984 21.252 ;
  LAYER M2 ;
        RECT 9.488 18.648 11.984 21.252 ;
  LAYER M1 ;
        RECT 9.488 15.54 11.984 18.144 ;
  LAYER M3 ;
        RECT 9.488 15.54 11.984 18.144 ;
  LAYER M2 ;
        RECT 9.488 15.54 11.984 18.144 ;
  LAYER M1 ;
        RECT 6.512 27.972 9.008 30.576 ;
  LAYER M3 ;
        RECT 6.512 27.972 9.008 30.576 ;
  LAYER M2 ;
        RECT 6.512 27.972 9.008 30.576 ;
  LAYER M1 ;
        RECT 6.512 24.864 9.008 27.468 ;
  LAYER M3 ;
        RECT 6.512 24.864 9.008 27.468 ;
  LAYER M2 ;
        RECT 6.512 24.864 9.008 27.468 ;
  LAYER M1 ;
        RECT 6.512 21.756 9.008 24.36 ;
  LAYER M3 ;
        RECT 6.512 21.756 9.008 24.36 ;
  LAYER M2 ;
        RECT 6.512 21.756 9.008 24.36 ;
  LAYER M1 ;
        RECT 6.512 18.648 9.008 21.252 ;
  LAYER M3 ;
        RECT 6.512 18.648 9.008 21.252 ;
  LAYER M2 ;
        RECT 6.512 18.648 9.008 21.252 ;
  LAYER M1 ;
        RECT 6.512 15.54 9.008 18.144 ;
  LAYER M3 ;
        RECT 6.512 15.54 9.008 18.144 ;
  LAYER M2 ;
        RECT 6.512 15.54 9.008 18.144 ;
  LAYER M1 ;
        RECT 3.536 27.972 6.032 30.576 ;
  LAYER M3 ;
        RECT 3.536 27.972 6.032 30.576 ;
  LAYER M2 ;
        RECT 3.536 27.972 6.032 30.576 ;
  LAYER M1 ;
        RECT 3.536 24.864 6.032 27.468 ;
  LAYER M3 ;
        RECT 3.536 24.864 6.032 27.468 ;
  LAYER M2 ;
        RECT 3.536 24.864 6.032 27.468 ;
  LAYER M1 ;
        RECT 3.536 21.756 6.032 24.36 ;
  LAYER M3 ;
        RECT 3.536 21.756 6.032 24.36 ;
  LAYER M2 ;
        RECT 3.536 21.756 6.032 24.36 ;
  LAYER M1 ;
        RECT 3.536 18.648 6.032 21.252 ;
  LAYER M3 ;
        RECT 3.536 18.648 6.032 21.252 ;
  LAYER M2 ;
        RECT 3.536 18.648 6.032 21.252 ;
  LAYER M1 ;
        RECT 3.536 15.54 6.032 18.144 ;
  LAYER M3 ;
        RECT 3.536 15.54 6.032 18.144 ;
  LAYER M2 ;
        RECT 3.536 15.54 6.032 18.144 ;
  LAYER M1 ;
        RECT 0.56 27.972 3.056 30.576 ;
  LAYER M3 ;
        RECT 0.56 27.972 3.056 30.576 ;
  LAYER M2 ;
        RECT 0.56 27.972 3.056 30.576 ;
  LAYER M1 ;
        RECT 0.56 24.864 3.056 27.468 ;
  LAYER M3 ;
        RECT 0.56 24.864 3.056 27.468 ;
  LAYER M2 ;
        RECT 0.56 24.864 3.056 27.468 ;
  LAYER M1 ;
        RECT 0.56 21.756 3.056 24.36 ;
  LAYER M3 ;
        RECT 0.56 21.756 3.056 24.36 ;
  LAYER M2 ;
        RECT 0.56 21.756 3.056 24.36 ;
  LAYER M1 ;
        RECT 0.56 18.648 3.056 21.252 ;
  LAYER M3 ;
        RECT 0.56 18.648 3.056 21.252 ;
  LAYER M2 ;
        RECT 0.56 18.648 3.056 21.252 ;
  LAYER M1 ;
        RECT 0.56 15.54 3.056 18.144 ;
  LAYER M3 ;
        RECT 0.56 15.54 3.056 18.144 ;
  LAYER M2 ;
        RECT 0.56 15.54 3.056 18.144 ;
  LAYER M1 ;
        RECT 41.008 14.244 41.04 14.316 ;
  LAYER M2 ;
        RECT 40.988 14.264 41.06 14.296 ;
  LAYER M1 ;
        RECT 38.096 14.244 38.128 14.316 ;
  LAYER M2 ;
        RECT 38.076 14.264 38.148 14.296 ;
  LAYER M2 ;
        RECT 38.112 14.264 41.024 14.296 ;
  LAYER M2 ;
        RECT 40.684 0.908 41.396 0.94 ;
  LAYER M1 ;
        RECT 38.176 31.044 38.208 31.116 ;
  LAYER M2 ;
        RECT 38.156 31.064 38.228 31.096 ;
  LAYER M1 ;
        RECT 41.152 31.044 41.184 31.116 ;
  LAYER M2 ;
        RECT 41.132 31.064 41.204 31.096 ;
  LAYER M2 ;
        RECT 38.192 31.064 41.168 31.096 ;
  LAYER M2 ;
        RECT 40.944 14.264 40.976 14.296 ;
  LAYER M3 ;
        RECT 40.94 0.924 40.98 14.28 ;
  LAYER M2 ;
        RECT 40.944 0.908 40.976 0.94 ;
  LAYER M2 ;
        RECT 38.144 14.264 38.176 14.296 ;
  LAYER M3 ;
        RECT 38.14 14.28 38.18 31.08 ;
  LAYER M2 ;
        RECT 38.144 31.064 38.176 31.096 ;
  LAYER M1 ;
        RECT 41.232 1.308 41.264 1.38 ;
  LAYER M2 ;
        RECT 41.212 1.328 41.284 1.36 ;
  LAYER M1 ;
        RECT 38.256 1.308 38.288 1.38 ;
  LAYER M2 ;
        RECT 38.236 1.328 38.308 1.36 ;
  LAYER M2 ;
        RECT 38.272 1.328 41.248 1.36 ;
  LAYER M2 ;
        RECT 42.044 0.32 42.116 0.352 ;
  LAYER M2 ;
        RECT 31.884 0.32 31.956 0.352 ;
  LAYER M2 ;
        RECT 41.264 1.328 41.296 1.36 ;
  LAYER M3 ;
        RECT 41.26 0.336 41.3 1.344 ;
  LAYER M4 ;
        RECT 41.28 0.316 42.08 0.356 ;
  LAYER M3 ;
        RECT 42.06 0.316 42.1 0.356 ;
  LAYER M2 ;
        RECT 42.064 0.32 42.096 0.352 ;
  LAYER M2 ;
        RECT 38.224 1.328 38.256 1.36 ;
  LAYER M3 ;
        RECT 38.22 0.336 38.26 1.344 ;
  LAYER M4 ;
        RECT 31.92 0.316 38.24 0.356 ;
  LAYER M3 ;
        RECT 31.9 0.316 31.94 0.356 ;
  LAYER M2 ;
        RECT 31.904 0.32 31.936 0.352 ;
  LAYER M2 ;
        RECT 39.324 0.908 40.036 0.94 ;
  LAYER M1 ;
        RECT 38.4 15 38.432 15.072 ;
  LAYER M2 ;
        RECT 38.38 15.02 38.452 15.052 ;
  LAYER M1 ;
        RECT 41.312 15 41.344 15.072 ;
  LAYER M2 ;
        RECT 41.292 15.02 41.364 15.052 ;
  LAYER M2 ;
        RECT 38.416 15.02 41.328 15.052 ;
  LAYER M2 ;
        RECT 39.984 0.908 40.016 0.94 ;
  LAYER M3 ;
        RECT 39.98 0.924 40.02 1.68 ;
  LAYER M4 ;
        RECT 40 1.66 40.08 1.7 ;
  LAYER M5 ;
        RECT 40.048 1.68 40.112 15.036 ;
  LAYER M4 ;
        RECT 40.06 15.016 40.1 15.056 ;
  LAYER M3 ;
        RECT 40.06 15.016 40.1 15.056 ;
  LAYER M2 ;
        RECT 40.064 15.02 40.096 15.052 ;
  LAYER M1 ;
        RECT 38.48 5.004 38.512 5.076 ;
  LAYER M2 ;
        RECT 38.46 5.024 38.532 5.056 ;
  LAYER M2 ;
        RECT 38.496 5.024 41.248 5.056 ;
  LAYER M1 ;
        RECT 41.232 5.004 41.264 5.076 ;
  LAYER M2 ;
        RECT 41.212 5.024 41.284 5.056 ;
  LAYER M1 ;
        RECT 38.48 8.112 38.512 8.184 ;
  LAYER M2 ;
        RECT 38.46 8.132 38.532 8.164 ;
  LAYER M2 ;
        RECT 38.496 8.132 41.248 8.164 ;
  LAYER M1 ;
        RECT 41.232 8.112 41.264 8.184 ;
  LAYER M2 ;
        RECT 41.212 8.132 41.284 8.164 ;
  LAYER M1 ;
        RECT 41.456 5.004 41.488 5.076 ;
  LAYER M2 ;
        RECT 41.436 5.024 41.508 5.056 ;
  LAYER M1 ;
        RECT 41.456 4.872 41.488 5.04 ;
  LAYER M1 ;
        RECT 41.456 4.836 41.488 4.908 ;
  LAYER M2 ;
        RECT 41.436 4.856 41.508 4.888 ;
  LAYER M2 ;
        RECT 41.248 4.856 41.472 4.888 ;
  LAYER M1 ;
        RECT 41.232 4.836 41.264 4.908 ;
  LAYER M2 ;
        RECT 41.212 4.856 41.284 4.888 ;
  LAYER M1 ;
        RECT 41.456 8.112 41.488 8.184 ;
  LAYER M2 ;
        RECT 41.436 8.132 41.508 8.164 ;
  LAYER M1 ;
        RECT 41.456 7.98 41.488 8.148 ;
  LAYER M1 ;
        RECT 41.456 7.944 41.488 8.016 ;
  LAYER M2 ;
        RECT 41.436 7.964 41.508 7.996 ;
  LAYER M2 ;
        RECT 41.248 7.964 41.472 7.996 ;
  LAYER M1 ;
        RECT 41.232 7.944 41.264 8.016 ;
  LAYER M2 ;
        RECT 41.212 7.964 41.284 7.996 ;
  LAYER M1 ;
        RECT 41.232 1.308 41.264 1.38 ;
  LAYER M2 ;
        RECT 41.212 1.328 41.284 1.36 ;
  LAYER M1 ;
        RECT 41.232 1.344 41.264 1.596 ;
  LAYER M1 ;
        RECT 41.232 1.596 41.264 8.148 ;
  LAYER M1 ;
        RECT 35.504 8.112 35.536 8.184 ;
  LAYER M2 ;
        RECT 35.484 8.132 35.556 8.164 ;
  LAYER M2 ;
        RECT 35.52 8.132 38.272 8.164 ;
  LAYER M1 ;
        RECT 38.256 8.112 38.288 8.184 ;
  LAYER M2 ;
        RECT 38.236 8.132 38.308 8.164 ;
  LAYER M1 ;
        RECT 35.504 5.004 35.536 5.076 ;
  LAYER M2 ;
        RECT 35.484 5.024 35.556 5.056 ;
  LAYER M2 ;
        RECT 35.52 5.024 38.272 5.056 ;
  LAYER M1 ;
        RECT 38.256 5.004 38.288 5.076 ;
  LAYER M2 ;
        RECT 38.236 5.024 38.308 5.056 ;
  LAYER M1 ;
        RECT 38.256 1.308 38.288 1.38 ;
  LAYER M2 ;
        RECT 38.236 1.328 38.308 1.36 ;
  LAYER M1 ;
        RECT 38.256 1.344 38.288 1.596 ;
  LAYER M1 ;
        RECT 38.256 1.596 38.288 8.148 ;
  LAYER M2 ;
        RECT 38.272 1.328 41.248 1.36 ;
  LAYER M1 ;
        RECT 44.432 1.896 44.464 1.968 ;
  LAYER M2 ;
        RECT 44.412 1.916 44.484 1.948 ;
  LAYER M1 ;
        RECT 44.432 1.764 44.464 1.932 ;
  LAYER M1 ;
        RECT 44.432 1.728 44.464 1.8 ;
  LAYER M2 ;
        RECT 44.412 1.748 44.484 1.78 ;
  LAYER M2 ;
        RECT 44.224 1.748 44.448 1.78 ;
  LAYER M1 ;
        RECT 44.208 1.728 44.24 1.8 ;
  LAYER M2 ;
        RECT 44.188 1.748 44.26 1.78 ;
  LAYER M1 ;
        RECT 44.432 5.004 44.464 5.076 ;
  LAYER M2 ;
        RECT 44.412 5.024 44.484 5.056 ;
  LAYER M1 ;
        RECT 44.432 4.872 44.464 5.04 ;
  LAYER M1 ;
        RECT 44.432 4.836 44.464 4.908 ;
  LAYER M2 ;
        RECT 44.412 4.856 44.484 4.888 ;
  LAYER M2 ;
        RECT 44.224 4.856 44.448 4.888 ;
  LAYER M1 ;
        RECT 44.208 4.836 44.24 4.908 ;
  LAYER M2 ;
        RECT 44.188 4.856 44.26 4.888 ;
  LAYER M1 ;
        RECT 44.432 8.112 44.464 8.184 ;
  LAYER M2 ;
        RECT 44.412 8.132 44.484 8.164 ;
  LAYER M1 ;
        RECT 44.432 7.98 44.464 8.148 ;
  LAYER M1 ;
        RECT 44.432 7.944 44.464 8.016 ;
  LAYER M2 ;
        RECT 44.412 7.964 44.484 7.996 ;
  LAYER M2 ;
        RECT 44.224 7.964 44.448 7.996 ;
  LAYER M1 ;
        RECT 44.208 7.944 44.24 8.016 ;
  LAYER M2 ;
        RECT 44.188 7.964 44.26 7.996 ;
  LAYER M1 ;
        RECT 44.432 11.22 44.464 11.292 ;
  LAYER M2 ;
        RECT 44.412 11.24 44.484 11.272 ;
  LAYER M1 ;
        RECT 44.432 11.088 44.464 11.256 ;
  LAYER M1 ;
        RECT 44.432 11.052 44.464 11.124 ;
  LAYER M2 ;
        RECT 44.412 11.072 44.484 11.104 ;
  LAYER M2 ;
        RECT 44.224 11.072 44.448 11.104 ;
  LAYER M1 ;
        RECT 44.208 11.052 44.24 11.124 ;
  LAYER M2 ;
        RECT 44.188 11.072 44.26 11.104 ;
  LAYER M1 ;
        RECT 41.456 1.896 41.488 1.968 ;
  LAYER M2 ;
        RECT 41.436 1.916 41.508 1.948 ;
  LAYER M2 ;
        RECT 41.472 1.916 44.224 1.948 ;
  LAYER M1 ;
        RECT 44.208 1.896 44.24 1.968 ;
  LAYER M2 ;
        RECT 44.188 1.916 44.26 1.948 ;
  LAYER M1 ;
        RECT 41.456 11.22 41.488 11.292 ;
  LAYER M2 ;
        RECT 41.436 11.24 41.508 11.272 ;
  LAYER M2 ;
        RECT 41.472 11.24 44.224 11.272 ;
  LAYER M1 ;
        RECT 44.208 11.22 44.24 11.292 ;
  LAYER M2 ;
        RECT 44.188 11.24 44.26 11.272 ;
  LAYER M1 ;
        RECT 44.208 1.14 44.24 1.212 ;
  LAYER M2 ;
        RECT 44.188 1.16 44.26 1.192 ;
  LAYER M1 ;
        RECT 44.208 1.176 44.24 1.596 ;
  LAYER M1 ;
        RECT 44.208 1.596 44.24 11.256 ;
  LAYER M1 ;
        RECT 35.504 1.896 35.536 1.968 ;
  LAYER M2 ;
        RECT 35.484 1.916 35.556 1.948 ;
  LAYER M1 ;
        RECT 35.504 1.764 35.536 1.932 ;
  LAYER M1 ;
        RECT 35.504 1.728 35.536 1.8 ;
  LAYER M2 ;
        RECT 35.484 1.748 35.556 1.78 ;
  LAYER M2 ;
        RECT 35.296 1.748 35.52 1.78 ;
  LAYER M1 ;
        RECT 35.28 1.728 35.312 1.8 ;
  LAYER M2 ;
        RECT 35.26 1.748 35.332 1.78 ;
  LAYER M1 ;
        RECT 35.504 11.22 35.536 11.292 ;
  LAYER M2 ;
        RECT 35.484 11.24 35.556 11.272 ;
  LAYER M1 ;
        RECT 35.504 11.088 35.536 11.256 ;
  LAYER M1 ;
        RECT 35.504 11.052 35.536 11.124 ;
  LAYER M2 ;
        RECT 35.484 11.072 35.556 11.104 ;
  LAYER M2 ;
        RECT 35.296 11.072 35.52 11.104 ;
  LAYER M1 ;
        RECT 35.28 11.052 35.312 11.124 ;
  LAYER M2 ;
        RECT 35.26 11.072 35.332 11.104 ;
  LAYER M1 ;
        RECT 32.528 1.896 32.56 1.968 ;
  LAYER M2 ;
        RECT 32.508 1.916 32.58 1.948 ;
  LAYER M2 ;
        RECT 32.544 1.916 35.296 1.948 ;
  LAYER M1 ;
        RECT 35.28 1.896 35.312 1.968 ;
  LAYER M2 ;
        RECT 35.26 1.916 35.332 1.948 ;
  LAYER M1 ;
        RECT 32.528 5.004 32.56 5.076 ;
  LAYER M2 ;
        RECT 32.508 5.024 32.58 5.056 ;
  LAYER M2 ;
        RECT 32.544 5.024 35.296 5.056 ;
  LAYER M1 ;
        RECT 35.28 5.004 35.312 5.076 ;
  LAYER M2 ;
        RECT 35.26 5.024 35.332 5.056 ;
  LAYER M1 ;
        RECT 32.528 8.112 32.56 8.184 ;
  LAYER M2 ;
        RECT 32.508 8.132 32.58 8.164 ;
  LAYER M2 ;
        RECT 32.544 8.132 35.296 8.164 ;
  LAYER M1 ;
        RECT 35.28 8.112 35.312 8.184 ;
  LAYER M2 ;
        RECT 35.26 8.132 35.332 8.164 ;
  LAYER M1 ;
        RECT 32.528 11.22 32.56 11.292 ;
  LAYER M2 ;
        RECT 32.508 11.24 32.58 11.272 ;
  LAYER M2 ;
        RECT 32.544 11.24 35.296 11.272 ;
  LAYER M1 ;
        RECT 35.28 11.22 35.312 11.292 ;
  LAYER M2 ;
        RECT 35.26 11.24 35.332 11.272 ;
  LAYER M1 ;
        RECT 35.28 1.14 35.312 1.212 ;
  LAYER M2 ;
        RECT 35.26 1.16 35.332 1.192 ;
  LAYER M1 ;
        RECT 35.28 1.176 35.312 1.596 ;
  LAYER M1 ;
        RECT 35.28 1.596 35.312 11.256 ;
  LAYER M2 ;
        RECT 35.296 1.16 44.224 1.192 ;
  LAYER M1 ;
        RECT 38.48 11.22 38.512 11.292 ;
  LAYER M2 ;
        RECT 38.46 11.24 38.532 11.272 ;
  LAYER M2 ;
        RECT 38.496 11.24 41.472 11.272 ;
  LAYER M1 ;
        RECT 41.456 11.22 41.488 11.292 ;
  LAYER M2 ;
        RECT 41.436 11.24 41.508 11.272 ;
  LAYER M1 ;
        RECT 38.48 1.896 38.512 1.968 ;
  LAYER M2 ;
        RECT 38.46 1.916 38.532 1.948 ;
  LAYER M2 ;
        RECT 35.52 1.916 38.496 1.948 ;
  LAYER M1 ;
        RECT 35.504 1.896 35.536 1.968 ;
  LAYER M2 ;
        RECT 35.484 1.916 35.556 1.948 ;
  LAYER M1 ;
        RECT 40.848 7.44 40.88 7.512 ;
  LAYER M2 ;
        RECT 40.828 7.46 40.9 7.492 ;
  LAYER M2 ;
        RECT 40.864 7.46 41.088 7.492 ;
  LAYER M1 ;
        RECT 41.072 7.44 41.104 7.512 ;
  LAYER M2 ;
        RECT 41.052 7.46 41.124 7.492 ;
  LAYER M1 ;
        RECT 40.848 10.548 40.88 10.62 ;
  LAYER M2 ;
        RECT 40.828 10.568 40.9 10.6 ;
  LAYER M2 ;
        RECT 40.864 10.568 41.088 10.6 ;
  LAYER M1 ;
        RECT 41.072 10.548 41.104 10.62 ;
  LAYER M2 ;
        RECT 41.052 10.568 41.124 10.6 ;
  LAYER M1 ;
        RECT 43.824 7.44 43.856 7.512 ;
  LAYER M2 ;
        RECT 43.804 7.46 43.876 7.492 ;
  LAYER M1 ;
        RECT 41.088 7.46 43.84 7.492 ;
  LAYER M1 ;
        RECT 41.072 7.44 41.104 7.512 ;
  LAYER M2 ;
        RECT 41.052 7.46 41.124 7.492 ;
  LAYER M2 ;
        RECT 41.024 7.46 41.088 7.492 ;
  LAYER M1 ;
        RECT 41.008 7.44 41.04 7.512 ;
  LAYER M2 ;
        RECT 40.988 7.46 41.06 7.492 ;
  LAYER M1 ;
        RECT 43.824 10.548 43.856 10.62 ;
  LAYER M2 ;
        RECT 43.804 10.568 43.876 10.6 ;
  LAYER M1 ;
        RECT 41.088 10.568 43.84 10.6 ;
  LAYER M1 ;
        RECT 41.072 10.548 41.104 10.62 ;
  LAYER M2 ;
        RECT 41.052 10.568 41.124 10.6 ;
  LAYER M2 ;
        RECT 41.024 10.568 41.088 10.6 ;
  LAYER M1 ;
        RECT 41.008 10.548 41.04 10.62 ;
  LAYER M2 ;
        RECT 40.988 10.568 41.06 10.6 ;
  LAYER M1 ;
        RECT 41.008 14.244 41.04 14.316 ;
  LAYER M2 ;
        RECT 40.988 14.264 41.06 14.296 ;
  LAYER M1 ;
        RECT 41.008 14.028 41.04 14.28 ;
  LAYER M1 ;
        RECT 41.008 7.476 41.04 14.028 ;
  LAYER M1 ;
        RECT 37.872 10.548 37.904 10.62 ;
  LAYER M2 ;
        RECT 37.852 10.568 37.924 10.6 ;
  LAYER M2 ;
        RECT 37.888 10.568 38.112 10.6 ;
  LAYER M1 ;
        RECT 38.096 10.548 38.128 10.62 ;
  LAYER M2 ;
        RECT 38.076 10.568 38.148 10.6 ;
  LAYER M1 ;
        RECT 37.872 7.44 37.904 7.512 ;
  LAYER M2 ;
        RECT 37.852 7.46 37.924 7.492 ;
  LAYER M2 ;
        RECT 37.888 7.46 38.112 7.492 ;
  LAYER M1 ;
        RECT 38.096 7.44 38.128 7.512 ;
  LAYER M2 ;
        RECT 38.076 7.46 38.148 7.492 ;
  LAYER M1 ;
        RECT 38.096 14.244 38.128 14.316 ;
  LAYER M2 ;
        RECT 38.076 14.264 38.148 14.296 ;
  LAYER M1 ;
        RECT 38.096 14.028 38.128 14.28 ;
  LAYER M1 ;
        RECT 38.096 7.476 38.128 14.028 ;
  LAYER M2 ;
        RECT 38.112 14.264 41.024 14.296 ;
  LAYER M1 ;
        RECT 46.8 4.332 46.832 4.404 ;
  LAYER M2 ;
        RECT 46.78 4.352 46.852 4.384 ;
  LAYER M2 ;
        RECT 46.816 4.352 47.2 4.384 ;
  LAYER M1 ;
        RECT 47.184 4.332 47.216 4.404 ;
  LAYER M2 ;
        RECT 47.164 4.352 47.236 4.384 ;
  LAYER M1 ;
        RECT 46.8 7.44 46.832 7.512 ;
  LAYER M2 ;
        RECT 46.78 7.46 46.852 7.492 ;
  LAYER M2 ;
        RECT 46.816 7.46 47.2 7.492 ;
  LAYER M1 ;
        RECT 47.184 7.44 47.216 7.512 ;
  LAYER M2 ;
        RECT 47.164 7.46 47.236 7.492 ;
  LAYER M1 ;
        RECT 46.8 10.548 46.832 10.62 ;
  LAYER M2 ;
        RECT 46.78 10.568 46.852 10.6 ;
  LAYER M2 ;
        RECT 46.816 10.568 47.2 10.6 ;
  LAYER M1 ;
        RECT 47.184 10.548 47.216 10.62 ;
  LAYER M2 ;
        RECT 47.164 10.568 47.236 10.6 ;
  LAYER M1 ;
        RECT 46.8 13.656 46.832 13.728 ;
  LAYER M2 ;
        RECT 46.78 13.676 46.852 13.708 ;
  LAYER M2 ;
        RECT 46.816 13.676 47.2 13.708 ;
  LAYER M1 ;
        RECT 47.184 13.656 47.216 13.728 ;
  LAYER M2 ;
        RECT 47.164 13.676 47.236 13.708 ;
  LAYER M1 ;
        RECT 47.184 14.412 47.216 14.484 ;
  LAYER M2 ;
        RECT 47.164 14.432 47.236 14.464 ;
  LAYER M1 ;
        RECT 47.184 14.028 47.216 14.448 ;
  LAYER M1 ;
        RECT 47.184 4.368 47.216 14.028 ;
  LAYER M1 ;
        RECT 34.896 4.332 34.928 4.404 ;
  LAYER M2 ;
        RECT 34.876 4.352 34.948 4.384 ;
  LAYER M1 ;
        RECT 32.32 4.352 34.912 4.384 ;
  LAYER M1 ;
        RECT 32.304 4.332 32.336 4.404 ;
  LAYER M2 ;
        RECT 32.284 4.352 32.356 4.384 ;
  LAYER M2 ;
        RECT 32.256 4.352 32.32 4.384 ;
  LAYER M1 ;
        RECT 32.24 4.332 32.272 4.404 ;
  LAYER M2 ;
        RECT 32.22 4.352 32.292 4.384 ;
  LAYER M1 ;
        RECT 34.896 7.44 34.928 7.512 ;
  LAYER M2 ;
        RECT 34.876 7.46 34.948 7.492 ;
  LAYER M1 ;
        RECT 32.32 7.46 34.912 7.492 ;
  LAYER M1 ;
        RECT 32.304 7.44 32.336 7.512 ;
  LAYER M2 ;
        RECT 32.284 7.46 32.356 7.492 ;
  LAYER M2 ;
        RECT 32.256 7.46 32.32 7.492 ;
  LAYER M1 ;
        RECT 32.24 7.44 32.272 7.512 ;
  LAYER M2 ;
        RECT 32.22 7.46 32.292 7.492 ;
  LAYER M1 ;
        RECT 34.896 10.548 34.928 10.62 ;
  LAYER M2 ;
        RECT 34.876 10.568 34.948 10.6 ;
  LAYER M1 ;
        RECT 32.32 10.568 34.912 10.6 ;
  LAYER M1 ;
        RECT 32.304 10.548 32.336 10.62 ;
  LAYER M2 ;
        RECT 32.284 10.568 32.356 10.6 ;
  LAYER M2 ;
        RECT 32.256 10.568 32.32 10.6 ;
  LAYER M1 ;
        RECT 32.24 10.548 32.272 10.62 ;
  LAYER M2 ;
        RECT 32.22 10.568 32.292 10.6 ;
  LAYER M1 ;
        RECT 34.896 13.656 34.928 13.728 ;
  LAYER M2 ;
        RECT 34.876 13.676 34.948 13.708 ;
  LAYER M1 ;
        RECT 32.32 13.676 34.912 13.708 ;
  LAYER M1 ;
        RECT 32.304 13.656 32.336 13.728 ;
  LAYER M2 ;
        RECT 32.284 13.676 32.356 13.708 ;
  LAYER M2 ;
        RECT 32.256 13.676 32.32 13.708 ;
  LAYER M1 ;
        RECT 32.24 13.656 32.272 13.728 ;
  LAYER M2 ;
        RECT 32.22 13.676 32.292 13.708 ;
  LAYER M1 ;
        RECT 32.24 14.412 32.272 14.484 ;
  LAYER M2 ;
        RECT 32.22 14.432 32.292 14.464 ;
  LAYER M1 ;
        RECT 32.24 14.028 32.272 14.448 ;
  LAYER M1 ;
        RECT 32.24 4.536 32.272 14.028 ;
  LAYER M2 ;
        RECT 32.256 14.432 47.2 14.464 ;
  LAYER M1 ;
        RECT 43.824 4.332 43.856 4.404 ;
  LAYER M2 ;
        RECT 43.804 4.352 43.876 4.384 ;
  LAYER M2 ;
        RECT 43.84 4.352 46.816 4.384 ;
  LAYER M1 ;
        RECT 46.8 4.332 46.832 4.404 ;
  LAYER M2 ;
        RECT 46.78 4.352 46.852 4.384 ;
  LAYER M1 ;
        RECT 43.824 13.656 43.856 13.728 ;
  LAYER M2 ;
        RECT 43.804 13.676 43.876 13.708 ;
  LAYER M2 ;
        RECT 43.84 13.676 46.816 13.708 ;
  LAYER M1 ;
        RECT 46.8 13.656 46.832 13.728 ;
  LAYER M2 ;
        RECT 46.78 13.676 46.852 13.708 ;
  LAYER M1 ;
        RECT 40.848 13.656 40.88 13.728 ;
  LAYER M2 ;
        RECT 40.828 13.676 40.9 13.708 ;
  LAYER M2 ;
        RECT 40.864 13.676 43.84 13.708 ;
  LAYER M1 ;
        RECT 43.824 13.656 43.856 13.728 ;
  LAYER M2 ;
        RECT 43.804 13.676 43.876 13.708 ;
  LAYER M1 ;
        RECT 37.872 13.656 37.904 13.728 ;
  LAYER M2 ;
        RECT 37.852 13.676 37.924 13.708 ;
  LAYER M2 ;
        RECT 37.888 13.676 40.864 13.708 ;
  LAYER M1 ;
        RECT 40.848 13.656 40.88 13.728 ;
  LAYER M2 ;
        RECT 40.828 13.676 40.9 13.708 ;
  LAYER M1 ;
        RECT 37.872 4.332 37.904 4.404 ;
  LAYER M2 ;
        RECT 37.852 4.352 37.924 4.384 ;
  LAYER M2 ;
        RECT 34.912 4.352 37.888 4.384 ;
  LAYER M1 ;
        RECT 34.896 4.332 34.928 4.404 ;
  LAYER M2 ;
        RECT 34.876 4.352 34.948 4.384 ;
  LAYER M1 ;
        RECT 40.848 4.332 40.88 4.404 ;
  LAYER M2 ;
        RECT 40.828 4.352 40.9 4.384 ;
  LAYER M2 ;
        RECT 37.888 4.352 40.864 4.384 ;
  LAYER M1 ;
        RECT 37.872 4.332 37.904 4.404 ;
  LAYER M2 ;
        RECT 37.852 4.352 37.924 4.384 ;
  LAYER M1 ;
        RECT 44.384 1.848 46.88 4.452 ;
  LAYER M3 ;
        RECT 44.384 1.848 46.88 4.452 ;
  LAYER M2 ;
        RECT 44.384 1.848 46.88 4.452 ;
  LAYER M1 ;
        RECT 44.384 4.956 46.88 7.56 ;
  LAYER M3 ;
        RECT 44.384 4.956 46.88 7.56 ;
  LAYER M2 ;
        RECT 44.384 4.956 46.88 7.56 ;
  LAYER M1 ;
        RECT 44.384 8.064 46.88 10.668 ;
  LAYER M3 ;
        RECT 44.384 8.064 46.88 10.668 ;
  LAYER M2 ;
        RECT 44.384 8.064 46.88 10.668 ;
  LAYER M1 ;
        RECT 44.384 11.172 46.88 13.776 ;
  LAYER M3 ;
        RECT 44.384 11.172 46.88 13.776 ;
  LAYER M2 ;
        RECT 44.384 11.172 46.88 13.776 ;
  LAYER M1 ;
        RECT 41.408 1.848 43.904 4.452 ;
  LAYER M3 ;
        RECT 41.408 1.848 43.904 4.452 ;
  LAYER M2 ;
        RECT 41.408 1.848 43.904 4.452 ;
  LAYER M1 ;
        RECT 41.408 4.956 43.904 7.56 ;
  LAYER M3 ;
        RECT 41.408 4.956 43.904 7.56 ;
  LAYER M2 ;
        RECT 41.408 4.956 43.904 7.56 ;
  LAYER M1 ;
        RECT 41.408 8.064 43.904 10.668 ;
  LAYER M3 ;
        RECT 41.408 8.064 43.904 10.668 ;
  LAYER M2 ;
        RECT 41.408 8.064 43.904 10.668 ;
  LAYER M1 ;
        RECT 41.408 11.172 43.904 13.776 ;
  LAYER M3 ;
        RECT 41.408 11.172 43.904 13.776 ;
  LAYER M2 ;
        RECT 41.408 11.172 43.904 13.776 ;
  LAYER M1 ;
        RECT 38.432 1.848 40.928 4.452 ;
  LAYER M3 ;
        RECT 38.432 1.848 40.928 4.452 ;
  LAYER M2 ;
        RECT 38.432 1.848 40.928 4.452 ;
  LAYER M1 ;
        RECT 38.432 4.956 40.928 7.56 ;
  LAYER M3 ;
        RECT 38.432 4.956 40.928 7.56 ;
  LAYER M2 ;
        RECT 38.432 4.956 40.928 7.56 ;
  LAYER M1 ;
        RECT 38.432 8.064 40.928 10.668 ;
  LAYER M3 ;
        RECT 38.432 8.064 40.928 10.668 ;
  LAYER M2 ;
        RECT 38.432 8.064 40.928 10.668 ;
  LAYER M1 ;
        RECT 38.432 11.172 40.928 13.776 ;
  LAYER M3 ;
        RECT 38.432 11.172 40.928 13.776 ;
  LAYER M2 ;
        RECT 38.432 11.172 40.928 13.776 ;
  LAYER M1 ;
        RECT 35.456 1.848 37.952 4.452 ;
  LAYER M3 ;
        RECT 35.456 1.848 37.952 4.452 ;
  LAYER M2 ;
        RECT 35.456 1.848 37.952 4.452 ;
  LAYER M1 ;
        RECT 35.456 4.956 37.952 7.56 ;
  LAYER M3 ;
        RECT 35.456 4.956 37.952 7.56 ;
  LAYER M2 ;
        RECT 35.456 4.956 37.952 7.56 ;
  LAYER M1 ;
        RECT 35.456 8.064 37.952 10.668 ;
  LAYER M3 ;
        RECT 35.456 8.064 37.952 10.668 ;
  LAYER M2 ;
        RECT 35.456 8.064 37.952 10.668 ;
  LAYER M1 ;
        RECT 35.456 11.172 37.952 13.776 ;
  LAYER M3 ;
        RECT 35.456 11.172 37.952 13.776 ;
  LAYER M2 ;
        RECT 35.456 11.172 37.952 13.776 ;
  LAYER M1 ;
        RECT 32.48 1.848 34.976 4.452 ;
  LAYER M3 ;
        RECT 32.48 1.848 34.976 4.452 ;
  LAYER M2 ;
        RECT 32.48 1.848 34.976 4.452 ;
  LAYER M1 ;
        RECT 32.48 4.956 34.976 7.56 ;
  LAYER M3 ;
        RECT 32.48 4.956 34.976 7.56 ;
  LAYER M2 ;
        RECT 32.48 4.956 34.976 7.56 ;
  LAYER M1 ;
        RECT 32.48 8.064 34.976 10.668 ;
  LAYER M3 ;
        RECT 32.48 8.064 34.976 10.668 ;
  LAYER M2 ;
        RECT 32.48 8.064 34.976 10.668 ;
  LAYER M1 ;
        RECT 32.48 11.172 34.976 13.776 ;
  LAYER M3 ;
        RECT 32.48 11.172 34.976 13.776 ;
  LAYER M2 ;
        RECT 32.48 11.172 34.976 13.776 ;
  LAYER M1 ;
        RECT 42.144 0.216 42.176 0.876 ;
  LAYER M1 ;
        RECT 42.224 0.216 42.256 0.876 ;
  LAYER M1 ;
        RECT 42.064 0.656 42.096 0.688 ;
  LAYER M1 ;
        RECT 31.824 0.216 31.856 0.876 ;
  LAYER M1 ;
        RECT 31.744 0.216 31.776 0.876 ;
  LAYER M1 ;
        RECT 31.904 0.656 31.936 0.688 ;
  LAYER M1 ;
        RECT 40.784 0.3 40.816 0.96 ;
  LAYER M1 ;
        RECT 41.424 0.3 41.456 0.96 ;
  LAYER M1 ;
        RECT 40.704 0.3 40.736 0.96 ;
  LAYER M1 ;
        RECT 41.344 0.3 41.376 0.96 ;
  LAYER M1 ;
        RECT 40.864 0.3 40.896 0.96 ;
  LAYER M1 ;
        RECT 41.504 0.488 41.536 0.52 ;
  LAYER M1 ;
        RECT 39.424 0.3 39.456 0.96 ;
  LAYER M1 ;
        RECT 40.064 0.3 40.096 0.96 ;
  LAYER M1 ;
        RECT 39.344 0.3 39.376 0.96 ;
  LAYER M1 ;
        RECT 39.984 0.3 40.016 0.96 ;
  LAYER M1 ;
        RECT 39.504 0.3 39.536 0.96 ;
  LAYER M1 ;
        RECT 40.144 0.488 40.176 0.52 ;
  LAYER M1 ;
        RECT 40.928 24.24 40.96 24.312 ;
  LAYER M2 ;
        RECT 40.908 24.26 40.98 24.292 ;
  LAYER M2 ;
        RECT 38.192 24.26 40.944 24.292 ;
  LAYER M1 ;
        RECT 38.176 24.24 38.208 24.312 ;
  LAYER M2 ;
        RECT 38.156 24.26 38.228 24.292 ;
  LAYER M1 ;
        RECT 37.952 21.132 37.984 21.204 ;
  LAYER M2 ;
        RECT 37.932 21.152 38.004 21.184 ;
  LAYER M1 ;
        RECT 37.952 21.168 37.984 21.336 ;
  LAYER M1 ;
        RECT 37.952 21.3 37.984 21.372 ;
  LAYER M2 ;
        RECT 37.932 21.32 38.004 21.352 ;
  LAYER M2 ;
        RECT 37.968 21.32 38.192 21.352 ;
  LAYER M1 ;
        RECT 38.176 21.3 38.208 21.372 ;
  LAYER M2 ;
        RECT 38.156 21.32 38.228 21.352 ;
  LAYER M1 ;
        RECT 38.176 31.044 38.208 31.116 ;
  LAYER M2 ;
        RECT 38.156 31.064 38.228 31.096 ;
  LAYER M1 ;
        RECT 38.176 30.828 38.208 31.08 ;
  LAYER M1 ;
        RECT 38.176 21.336 38.208 30.828 ;
  LAYER M1 ;
        RECT 43.904 27.348 43.936 27.42 ;
  LAYER M2 ;
        RECT 43.884 27.368 43.956 27.4 ;
  LAYER M2 ;
        RECT 41.168 27.368 43.92 27.4 ;
  LAYER M1 ;
        RECT 41.152 27.348 41.184 27.42 ;
  LAYER M2 ;
        RECT 41.132 27.368 41.204 27.4 ;
  LAYER M1 ;
        RECT 41.152 31.044 41.184 31.116 ;
  LAYER M2 ;
        RECT 41.132 31.064 41.204 31.096 ;
  LAYER M1 ;
        RECT 41.152 30.828 41.184 31.08 ;
  LAYER M1 ;
        RECT 41.152 27.384 41.184 30.828 ;
  LAYER M2 ;
        RECT 38.192 31.064 41.168 31.096 ;
  LAYER M1 ;
        RECT 37.952 24.24 37.984 24.312 ;
  LAYER M2 ;
        RECT 37.932 24.26 38.004 24.292 ;
  LAYER M2 ;
        RECT 35.216 24.26 37.968 24.292 ;
  LAYER M1 ;
        RECT 35.2 24.24 35.232 24.312 ;
  LAYER M2 ;
        RECT 35.18 24.26 35.252 24.292 ;
  LAYER M1 ;
        RECT 37.952 27.348 37.984 27.42 ;
  LAYER M2 ;
        RECT 37.932 27.368 38.004 27.4 ;
  LAYER M2 ;
        RECT 35.216 27.368 37.968 27.4 ;
  LAYER M1 ;
        RECT 35.2 27.348 35.232 27.42 ;
  LAYER M2 ;
        RECT 35.18 27.368 35.252 27.4 ;
  LAYER M1 ;
        RECT 35.2 31.212 35.232 31.284 ;
  LAYER M2 ;
        RECT 35.18 31.232 35.252 31.264 ;
  LAYER M1 ;
        RECT 35.2 30.828 35.232 31.248 ;
  LAYER M1 ;
        RECT 35.2 24.276 35.232 30.828 ;
  LAYER M1 ;
        RECT 43.904 24.24 43.936 24.312 ;
  LAYER M2 ;
        RECT 43.884 24.26 43.956 24.292 ;
  LAYER M1 ;
        RECT 43.904 24.276 43.936 24.444 ;
  LAYER M1 ;
        RECT 43.904 24.408 43.936 24.48 ;
  LAYER M2 ;
        RECT 43.884 24.428 43.956 24.46 ;
  LAYER M2 ;
        RECT 43.92 24.428 44.144 24.46 ;
  LAYER M1 ;
        RECT 44.128 24.408 44.16 24.48 ;
  LAYER M2 ;
        RECT 44.108 24.428 44.18 24.46 ;
  LAYER M1 ;
        RECT 43.904 21.132 43.936 21.204 ;
  LAYER M2 ;
        RECT 43.884 21.152 43.956 21.184 ;
  LAYER M1 ;
        RECT 43.904 21.168 43.936 21.336 ;
  LAYER M1 ;
        RECT 43.904 21.3 43.936 21.372 ;
  LAYER M2 ;
        RECT 43.884 21.32 43.956 21.352 ;
  LAYER M2 ;
        RECT 43.92 21.32 44.144 21.352 ;
  LAYER M1 ;
        RECT 44.128 21.3 44.16 21.372 ;
  LAYER M2 ;
        RECT 44.108 21.32 44.18 21.352 ;
  LAYER M1 ;
        RECT 44.128 31.212 44.16 31.284 ;
  LAYER M2 ;
        RECT 44.108 31.232 44.18 31.264 ;
  LAYER M1 ;
        RECT 44.128 30.828 44.16 31.248 ;
  LAYER M1 ;
        RECT 44.128 21.336 44.16 30.828 ;
  LAYER M2 ;
        RECT 35.216 31.232 44.144 31.264 ;
  LAYER M1 ;
        RECT 40.928 27.348 40.96 27.42 ;
  LAYER M2 ;
        RECT 40.908 27.368 40.98 27.4 ;
  LAYER M2 ;
        RECT 37.968 27.368 40.944 27.4 ;
  LAYER M1 ;
        RECT 37.952 27.348 37.984 27.42 ;
  LAYER M2 ;
        RECT 37.932 27.368 38.004 27.4 ;
  LAYER M1 ;
        RECT 40.928 21.132 40.96 21.204 ;
  LAYER M2 ;
        RECT 40.908 21.152 40.98 21.184 ;
  LAYER M2 ;
        RECT 40.944 21.152 43.92 21.184 ;
  LAYER M1 ;
        RECT 43.904 21.132 43.936 21.204 ;
  LAYER M2 ;
        RECT 43.884 21.152 43.956 21.184 ;
  LAYER M1 ;
        RECT 34.976 30.456 35.008 30.528 ;
  LAYER M2 ;
        RECT 34.956 30.476 35.028 30.508 ;
  LAYER M2 ;
        RECT 32.24 30.476 34.992 30.508 ;
  LAYER M1 ;
        RECT 32.224 30.456 32.256 30.528 ;
  LAYER M2 ;
        RECT 32.204 30.476 32.276 30.508 ;
  LAYER M1 ;
        RECT 34.976 27.348 35.008 27.42 ;
  LAYER M2 ;
        RECT 34.956 27.368 35.028 27.4 ;
  LAYER M2 ;
        RECT 32.24 27.368 34.992 27.4 ;
  LAYER M1 ;
        RECT 32.224 27.348 32.256 27.42 ;
  LAYER M2 ;
        RECT 32.204 27.368 32.276 27.4 ;
  LAYER M1 ;
        RECT 34.976 24.24 35.008 24.312 ;
  LAYER M2 ;
        RECT 34.956 24.26 35.028 24.292 ;
  LAYER M2 ;
        RECT 32.24 24.26 34.992 24.292 ;
  LAYER M1 ;
        RECT 32.224 24.24 32.256 24.312 ;
  LAYER M2 ;
        RECT 32.204 24.26 32.276 24.292 ;
  LAYER M1 ;
        RECT 34.976 21.132 35.008 21.204 ;
  LAYER M2 ;
        RECT 34.956 21.152 35.028 21.184 ;
  LAYER M2 ;
        RECT 32.24 21.152 34.992 21.184 ;
  LAYER M1 ;
        RECT 32.224 21.132 32.256 21.204 ;
  LAYER M2 ;
        RECT 32.204 21.152 32.276 21.184 ;
  LAYER M1 ;
        RECT 34.976 18.024 35.008 18.096 ;
  LAYER M2 ;
        RECT 34.956 18.044 35.028 18.076 ;
  LAYER M2 ;
        RECT 32.24 18.044 34.992 18.076 ;
  LAYER M1 ;
        RECT 32.224 18.024 32.256 18.096 ;
  LAYER M2 ;
        RECT 32.204 18.044 32.276 18.076 ;
  LAYER M1 ;
        RECT 32.224 31.38 32.256 31.452 ;
  LAYER M2 ;
        RECT 32.204 31.4 32.276 31.432 ;
  LAYER M1 ;
        RECT 32.224 30.828 32.256 31.416 ;
  LAYER M1 ;
        RECT 32.224 18.06 32.256 30.828 ;
  LAYER M1 ;
        RECT 46.88 30.456 46.912 30.528 ;
  LAYER M2 ;
        RECT 46.86 30.476 46.932 30.508 ;
  LAYER M1 ;
        RECT 46.88 30.492 46.912 30.66 ;
  LAYER M1 ;
        RECT 46.88 30.624 46.912 30.696 ;
  LAYER M2 ;
        RECT 46.86 30.644 46.932 30.676 ;
  LAYER M2 ;
        RECT 46.896 30.644 47.12 30.676 ;
  LAYER M1 ;
        RECT 47.104 30.624 47.136 30.696 ;
  LAYER M2 ;
        RECT 47.084 30.644 47.156 30.676 ;
  LAYER M1 ;
        RECT 46.88 27.348 46.912 27.42 ;
  LAYER M2 ;
        RECT 46.86 27.368 46.932 27.4 ;
  LAYER M1 ;
        RECT 46.88 27.384 46.912 27.552 ;
  LAYER M1 ;
        RECT 46.88 27.516 46.912 27.588 ;
  LAYER M2 ;
        RECT 46.86 27.536 46.932 27.568 ;
  LAYER M2 ;
        RECT 46.896 27.536 47.12 27.568 ;
  LAYER M1 ;
        RECT 47.104 27.516 47.136 27.588 ;
  LAYER M2 ;
        RECT 47.084 27.536 47.156 27.568 ;
  LAYER M1 ;
        RECT 46.88 24.24 46.912 24.312 ;
  LAYER M2 ;
        RECT 46.86 24.26 46.932 24.292 ;
  LAYER M1 ;
        RECT 46.88 24.276 46.912 24.444 ;
  LAYER M1 ;
        RECT 46.88 24.408 46.912 24.48 ;
  LAYER M2 ;
        RECT 46.86 24.428 46.932 24.46 ;
  LAYER M2 ;
        RECT 46.896 24.428 47.12 24.46 ;
  LAYER M1 ;
        RECT 47.104 24.408 47.136 24.48 ;
  LAYER M2 ;
        RECT 47.084 24.428 47.156 24.46 ;
  LAYER M1 ;
        RECT 46.88 21.132 46.912 21.204 ;
  LAYER M2 ;
        RECT 46.86 21.152 46.932 21.184 ;
  LAYER M1 ;
        RECT 46.88 21.168 46.912 21.336 ;
  LAYER M1 ;
        RECT 46.88 21.3 46.912 21.372 ;
  LAYER M2 ;
        RECT 46.86 21.32 46.932 21.352 ;
  LAYER M2 ;
        RECT 46.896 21.32 47.12 21.352 ;
  LAYER M1 ;
        RECT 47.104 21.3 47.136 21.372 ;
  LAYER M2 ;
        RECT 47.084 21.32 47.156 21.352 ;
  LAYER M1 ;
        RECT 46.88 18.024 46.912 18.096 ;
  LAYER M2 ;
        RECT 46.86 18.044 46.932 18.076 ;
  LAYER M1 ;
        RECT 46.88 18.06 46.912 18.228 ;
  LAYER M1 ;
        RECT 46.88 18.192 46.912 18.264 ;
  LAYER M2 ;
        RECT 46.86 18.212 46.932 18.244 ;
  LAYER M2 ;
        RECT 46.896 18.212 47.12 18.244 ;
  LAYER M1 ;
        RECT 47.104 18.192 47.136 18.264 ;
  LAYER M2 ;
        RECT 47.084 18.212 47.156 18.244 ;
  LAYER M1 ;
        RECT 47.104 31.38 47.136 31.452 ;
  LAYER M2 ;
        RECT 47.084 31.4 47.156 31.432 ;
  LAYER M1 ;
        RECT 47.104 30.828 47.136 31.416 ;
  LAYER M1 ;
        RECT 47.104 18.228 47.136 30.828 ;
  LAYER M2 ;
        RECT 32.24 31.4 47.12 31.432 ;
  LAYER M1 ;
        RECT 37.952 30.456 37.984 30.528 ;
  LAYER M2 ;
        RECT 37.932 30.476 38.004 30.508 ;
  LAYER M2 ;
        RECT 34.992 30.476 37.968 30.508 ;
  LAYER M1 ;
        RECT 34.976 30.456 35.008 30.528 ;
  LAYER M2 ;
        RECT 34.956 30.476 35.028 30.508 ;
  LAYER M1 ;
        RECT 37.952 18.024 37.984 18.096 ;
  LAYER M2 ;
        RECT 37.932 18.044 38.004 18.076 ;
  LAYER M2 ;
        RECT 34.992 18.044 37.968 18.076 ;
  LAYER M1 ;
        RECT 34.976 18.024 35.008 18.096 ;
  LAYER M2 ;
        RECT 34.956 18.044 35.028 18.076 ;
  LAYER M1 ;
        RECT 40.928 18.024 40.96 18.096 ;
  LAYER M2 ;
        RECT 40.908 18.044 40.98 18.076 ;
  LAYER M2 ;
        RECT 37.968 18.044 40.944 18.076 ;
  LAYER M1 ;
        RECT 37.952 18.024 37.984 18.096 ;
  LAYER M2 ;
        RECT 37.932 18.044 38.004 18.076 ;
  LAYER M1 ;
        RECT 43.904 18.024 43.936 18.096 ;
  LAYER M2 ;
        RECT 43.884 18.044 43.956 18.076 ;
  LAYER M2 ;
        RECT 40.944 18.044 43.92 18.076 ;
  LAYER M1 ;
        RECT 40.928 18.024 40.96 18.096 ;
  LAYER M2 ;
        RECT 40.908 18.044 40.98 18.076 ;
  LAYER M1 ;
        RECT 43.904 30.456 43.936 30.528 ;
  LAYER M2 ;
        RECT 43.884 30.476 43.956 30.508 ;
  LAYER M2 ;
        RECT 43.92 30.476 46.896 30.508 ;
  LAYER M1 ;
        RECT 46.88 30.456 46.912 30.528 ;
  LAYER M2 ;
        RECT 46.86 30.476 46.932 30.508 ;
  LAYER M1 ;
        RECT 40.928 30.456 40.96 30.528 ;
  LAYER M2 ;
        RECT 40.908 30.476 40.98 30.508 ;
  LAYER M2 ;
        RECT 40.944 30.476 43.92 30.508 ;
  LAYER M1 ;
        RECT 43.904 30.456 43.936 30.528 ;
  LAYER M2 ;
        RECT 43.884 30.476 43.956 30.508 ;
  LAYER M1 ;
        RECT 38.56 21.804 38.592 21.876 ;
  LAYER M2 ;
        RECT 38.54 21.824 38.612 21.856 ;
  LAYER M2 ;
        RECT 38.352 21.824 38.576 21.856 ;
  LAYER M1 ;
        RECT 38.336 21.804 38.368 21.876 ;
  LAYER M2 ;
        RECT 38.316 21.824 38.388 21.856 ;
  LAYER M1 ;
        RECT 35.584 18.696 35.616 18.768 ;
  LAYER M2 ;
        RECT 35.564 18.716 35.636 18.748 ;
  LAYER M1 ;
        RECT 35.6 18.716 38.352 18.748 ;
  LAYER M1 ;
        RECT 38.336 18.696 38.368 18.768 ;
  LAYER M2 ;
        RECT 38.316 18.716 38.388 18.748 ;
  LAYER M2 ;
        RECT 38.352 18.716 38.416 18.748 ;
  LAYER M1 ;
        RECT 38.4 18.696 38.432 18.768 ;
  LAYER M2 ;
        RECT 38.38 18.716 38.452 18.748 ;
  LAYER M1 ;
        RECT 38.4 15 38.432 15.072 ;
  LAYER M2 ;
        RECT 38.38 15.02 38.452 15.052 ;
  LAYER M1 ;
        RECT 38.4 15.036 38.432 15.288 ;
  LAYER M1 ;
        RECT 38.4 15.288 38.432 21.84 ;
  LAYER M1 ;
        RECT 41.536 24.912 41.568 24.984 ;
  LAYER M2 ;
        RECT 41.516 24.932 41.588 24.964 ;
  LAYER M2 ;
        RECT 41.328 24.932 41.552 24.964 ;
  LAYER M1 ;
        RECT 41.312 24.912 41.344 24.984 ;
  LAYER M2 ;
        RECT 41.292 24.932 41.364 24.964 ;
  LAYER M1 ;
        RECT 41.312 15 41.344 15.072 ;
  LAYER M2 ;
        RECT 41.292 15.02 41.364 15.052 ;
  LAYER M1 ;
        RECT 41.312 15.036 41.344 15.288 ;
  LAYER M1 ;
        RECT 41.312 15.288 41.344 24.948 ;
  LAYER M2 ;
        RECT 38.416 15.02 41.328 15.052 ;
  LAYER M1 ;
        RECT 35.584 21.804 35.616 21.876 ;
  LAYER M2 ;
        RECT 35.564 21.824 35.636 21.856 ;
  LAYER M2 ;
        RECT 35.376 21.824 35.6 21.856 ;
  LAYER M1 ;
        RECT 35.36 21.804 35.392 21.876 ;
  LAYER M2 ;
        RECT 35.34 21.824 35.412 21.856 ;
  LAYER M1 ;
        RECT 35.584 24.912 35.616 24.984 ;
  LAYER M2 ;
        RECT 35.564 24.932 35.636 24.964 ;
  LAYER M2 ;
        RECT 35.376 24.932 35.6 24.964 ;
  LAYER M1 ;
        RECT 35.36 24.912 35.392 24.984 ;
  LAYER M2 ;
        RECT 35.34 24.932 35.412 24.964 ;
  LAYER M1 ;
        RECT 35.36 14.832 35.392 14.904 ;
  LAYER M2 ;
        RECT 35.34 14.852 35.412 14.884 ;
  LAYER M1 ;
        RECT 35.36 14.868 35.392 15.288 ;
  LAYER M1 ;
        RECT 35.36 15.288 35.392 24.948 ;
  LAYER M1 ;
        RECT 41.536 21.804 41.568 21.876 ;
  LAYER M2 ;
        RECT 41.516 21.824 41.588 21.856 ;
  LAYER M1 ;
        RECT 41.552 21.824 44.304 21.856 ;
  LAYER M1 ;
        RECT 44.288 21.804 44.32 21.876 ;
  LAYER M2 ;
        RECT 44.268 21.824 44.34 21.856 ;
  LAYER M2 ;
        RECT 44.304 21.824 44.368 21.856 ;
  LAYER M1 ;
        RECT 44.352 21.804 44.384 21.876 ;
  LAYER M2 ;
        RECT 44.332 21.824 44.404 21.856 ;
  LAYER M1 ;
        RECT 41.536 18.696 41.568 18.768 ;
  LAYER M2 ;
        RECT 41.516 18.716 41.588 18.748 ;
  LAYER M1 ;
        RECT 41.552 18.716 44.304 18.748 ;
  LAYER M1 ;
        RECT 44.288 18.696 44.32 18.768 ;
  LAYER M2 ;
        RECT 44.268 18.716 44.34 18.748 ;
  LAYER M2 ;
        RECT 44.304 18.716 44.368 18.748 ;
  LAYER M1 ;
        RECT 44.352 18.696 44.384 18.768 ;
  LAYER M2 ;
        RECT 44.332 18.716 44.404 18.748 ;
  LAYER M1 ;
        RECT 44.352 14.832 44.384 14.904 ;
  LAYER M2 ;
        RECT 44.332 14.852 44.404 14.884 ;
  LAYER M1 ;
        RECT 44.352 14.868 44.384 15.288 ;
  LAYER M1 ;
        RECT 44.352 15.288 44.384 21.672 ;
  LAYER M2 ;
        RECT 35.376 14.852 44.368 14.884 ;
  LAYER M1 ;
        RECT 38.56 24.912 38.592 24.984 ;
  LAYER M2 ;
        RECT 38.54 24.932 38.612 24.964 ;
  LAYER M2 ;
        RECT 35.6 24.932 38.576 24.964 ;
  LAYER M1 ;
        RECT 35.584 24.912 35.616 24.984 ;
  LAYER M2 ;
        RECT 35.564 24.932 35.636 24.964 ;
  LAYER M1 ;
        RECT 38.56 18.696 38.592 18.768 ;
  LAYER M2 ;
        RECT 38.54 18.716 38.612 18.748 ;
  LAYER M2 ;
        RECT 38.576 18.716 41.552 18.748 ;
  LAYER M1 ;
        RECT 41.536 18.696 41.568 18.768 ;
  LAYER M2 ;
        RECT 41.516 18.716 41.588 18.748 ;
  LAYER M1 ;
        RECT 32.608 28.02 32.64 28.092 ;
  LAYER M2 ;
        RECT 32.588 28.04 32.66 28.072 ;
  LAYER M2 ;
        RECT 32.4 28.04 32.624 28.072 ;
  LAYER M1 ;
        RECT 32.384 28.02 32.416 28.092 ;
  LAYER M2 ;
        RECT 32.364 28.04 32.436 28.072 ;
  LAYER M1 ;
        RECT 32.608 24.912 32.64 24.984 ;
  LAYER M2 ;
        RECT 32.588 24.932 32.66 24.964 ;
  LAYER M2 ;
        RECT 32.4 24.932 32.624 24.964 ;
  LAYER M1 ;
        RECT 32.384 24.912 32.416 24.984 ;
  LAYER M2 ;
        RECT 32.364 24.932 32.436 24.964 ;
  LAYER M1 ;
        RECT 32.608 21.804 32.64 21.876 ;
  LAYER M2 ;
        RECT 32.588 21.824 32.66 21.856 ;
  LAYER M2 ;
        RECT 32.4 21.824 32.624 21.856 ;
  LAYER M1 ;
        RECT 32.384 21.804 32.416 21.876 ;
  LAYER M2 ;
        RECT 32.364 21.824 32.436 21.856 ;
  LAYER M1 ;
        RECT 32.608 18.696 32.64 18.768 ;
  LAYER M2 ;
        RECT 32.588 18.716 32.66 18.748 ;
  LAYER M2 ;
        RECT 32.4 18.716 32.624 18.748 ;
  LAYER M1 ;
        RECT 32.384 18.696 32.416 18.768 ;
  LAYER M2 ;
        RECT 32.364 18.716 32.436 18.748 ;
  LAYER M1 ;
        RECT 32.608 15.588 32.64 15.66 ;
  LAYER M2 ;
        RECT 32.588 15.608 32.66 15.64 ;
  LAYER M2 ;
        RECT 32.4 15.608 32.624 15.64 ;
  LAYER M1 ;
        RECT 32.384 15.588 32.416 15.66 ;
  LAYER M2 ;
        RECT 32.364 15.608 32.436 15.64 ;
  LAYER M1 ;
        RECT 32.384 14.664 32.416 14.736 ;
  LAYER M2 ;
        RECT 32.364 14.684 32.436 14.716 ;
  LAYER M1 ;
        RECT 32.384 14.7 32.416 15.288 ;
  LAYER M1 ;
        RECT 32.384 15.288 32.416 28.056 ;
  LAYER M1 ;
        RECT 44.512 28.02 44.544 28.092 ;
  LAYER M2 ;
        RECT 44.492 28.04 44.564 28.072 ;
  LAYER M1 ;
        RECT 44.528 28.04 47.28 28.072 ;
  LAYER M1 ;
        RECT 47.264 28.02 47.296 28.092 ;
  LAYER M2 ;
        RECT 47.244 28.04 47.316 28.072 ;
  LAYER M2 ;
        RECT 47.28 28.04 47.344 28.072 ;
  LAYER M1 ;
        RECT 47.328 28.02 47.36 28.092 ;
  LAYER M2 ;
        RECT 47.308 28.04 47.38 28.072 ;
  LAYER M1 ;
        RECT 44.512 24.912 44.544 24.984 ;
  LAYER M2 ;
        RECT 44.492 24.932 44.564 24.964 ;
  LAYER M1 ;
        RECT 44.528 24.932 47.28 24.964 ;
  LAYER M1 ;
        RECT 47.264 24.912 47.296 24.984 ;
  LAYER M2 ;
        RECT 47.244 24.932 47.316 24.964 ;
  LAYER M2 ;
        RECT 47.28 24.932 47.344 24.964 ;
  LAYER M1 ;
        RECT 47.328 24.912 47.36 24.984 ;
  LAYER M2 ;
        RECT 47.308 24.932 47.38 24.964 ;
  LAYER M1 ;
        RECT 44.512 21.804 44.544 21.876 ;
  LAYER M2 ;
        RECT 44.492 21.824 44.564 21.856 ;
  LAYER M1 ;
        RECT 44.528 21.824 47.28 21.856 ;
  LAYER M1 ;
        RECT 47.264 21.804 47.296 21.876 ;
  LAYER M2 ;
        RECT 47.244 21.824 47.316 21.856 ;
  LAYER M2 ;
        RECT 47.28 21.824 47.344 21.856 ;
  LAYER M1 ;
        RECT 47.328 21.804 47.36 21.876 ;
  LAYER M2 ;
        RECT 47.308 21.824 47.38 21.856 ;
  LAYER M1 ;
        RECT 44.512 18.696 44.544 18.768 ;
  LAYER M2 ;
        RECT 44.492 18.716 44.564 18.748 ;
  LAYER M1 ;
        RECT 44.528 18.716 47.28 18.748 ;
  LAYER M1 ;
        RECT 47.264 18.696 47.296 18.768 ;
  LAYER M2 ;
        RECT 47.244 18.716 47.316 18.748 ;
  LAYER M2 ;
        RECT 47.28 18.716 47.344 18.748 ;
  LAYER M1 ;
        RECT 47.328 18.696 47.36 18.768 ;
  LAYER M2 ;
        RECT 47.308 18.716 47.38 18.748 ;
  LAYER M1 ;
        RECT 44.512 15.588 44.544 15.66 ;
  LAYER M2 ;
        RECT 44.492 15.608 44.564 15.64 ;
  LAYER M1 ;
        RECT 44.528 15.608 47.28 15.64 ;
  LAYER M1 ;
        RECT 47.264 15.588 47.296 15.66 ;
  LAYER M2 ;
        RECT 47.244 15.608 47.316 15.64 ;
  LAYER M2 ;
        RECT 47.28 15.608 47.344 15.64 ;
  LAYER M1 ;
        RECT 47.328 15.588 47.36 15.66 ;
  LAYER M2 ;
        RECT 47.308 15.608 47.38 15.64 ;
  LAYER M1 ;
        RECT 47.328 14.664 47.36 14.736 ;
  LAYER M2 ;
        RECT 47.308 14.684 47.38 14.716 ;
  LAYER M1 ;
        RECT 47.328 14.7 47.36 15.288 ;
  LAYER M1 ;
        RECT 47.328 15.288 47.36 27.888 ;
  LAYER M2 ;
        RECT 32.4 14.684 47.344 14.716 ;
  LAYER M1 ;
        RECT 35.584 28.02 35.616 28.092 ;
  LAYER M2 ;
        RECT 35.564 28.04 35.636 28.072 ;
  LAYER M2 ;
        RECT 32.624 28.04 35.6 28.072 ;
  LAYER M1 ;
        RECT 32.608 28.02 32.64 28.092 ;
  LAYER M2 ;
        RECT 32.588 28.04 32.66 28.072 ;
  LAYER M1 ;
        RECT 35.584 15.588 35.616 15.66 ;
  LAYER M2 ;
        RECT 35.564 15.608 35.636 15.64 ;
  LAYER M2 ;
        RECT 32.624 15.608 35.6 15.64 ;
  LAYER M1 ;
        RECT 32.608 15.588 32.64 15.66 ;
  LAYER M2 ;
        RECT 32.588 15.608 32.66 15.64 ;
  LAYER M1 ;
        RECT 38.56 15.588 38.592 15.66 ;
  LAYER M2 ;
        RECT 38.54 15.608 38.612 15.64 ;
  LAYER M2 ;
        RECT 35.6 15.608 38.576 15.64 ;
  LAYER M1 ;
        RECT 35.584 15.588 35.616 15.66 ;
  LAYER M2 ;
        RECT 35.564 15.608 35.636 15.64 ;
  LAYER M1 ;
        RECT 41.536 15.588 41.568 15.66 ;
  LAYER M2 ;
        RECT 41.516 15.608 41.588 15.64 ;
  LAYER M2 ;
        RECT 38.576 15.608 41.552 15.64 ;
  LAYER M1 ;
        RECT 38.56 15.588 38.592 15.66 ;
  LAYER M2 ;
        RECT 38.54 15.608 38.612 15.64 ;
  LAYER M1 ;
        RECT 41.536 28.02 41.568 28.092 ;
  LAYER M2 ;
        RECT 41.516 28.04 41.588 28.072 ;
  LAYER M2 ;
        RECT 41.552 28.04 44.528 28.072 ;
  LAYER M1 ;
        RECT 44.512 28.02 44.544 28.092 ;
  LAYER M2 ;
        RECT 44.492 28.04 44.564 28.072 ;
  LAYER M1 ;
        RECT 38.56 28.02 38.592 28.092 ;
  LAYER M2 ;
        RECT 38.54 28.04 38.612 28.072 ;
  LAYER M2 ;
        RECT 38.576 28.04 41.552 28.072 ;
  LAYER M1 ;
        RECT 41.536 28.02 41.568 28.092 ;
  LAYER M2 ;
        RECT 41.516 28.04 41.588 28.072 ;
  LAYER M1 ;
        RECT 32.56 27.972 35.056 30.576 ;
  LAYER M3 ;
        RECT 32.56 27.972 35.056 30.576 ;
  LAYER M2 ;
        RECT 32.56 27.972 35.056 30.576 ;
  LAYER M1 ;
        RECT 32.56 24.864 35.056 27.468 ;
  LAYER M3 ;
        RECT 32.56 24.864 35.056 27.468 ;
  LAYER M2 ;
        RECT 32.56 24.864 35.056 27.468 ;
  LAYER M1 ;
        RECT 32.56 21.756 35.056 24.36 ;
  LAYER M3 ;
        RECT 32.56 21.756 35.056 24.36 ;
  LAYER M2 ;
        RECT 32.56 21.756 35.056 24.36 ;
  LAYER M1 ;
        RECT 32.56 18.648 35.056 21.252 ;
  LAYER M3 ;
        RECT 32.56 18.648 35.056 21.252 ;
  LAYER M2 ;
        RECT 32.56 18.648 35.056 21.252 ;
  LAYER M1 ;
        RECT 32.56 15.54 35.056 18.144 ;
  LAYER M3 ;
        RECT 32.56 15.54 35.056 18.144 ;
  LAYER M2 ;
        RECT 32.56 15.54 35.056 18.144 ;
  LAYER M1 ;
        RECT 35.536 27.972 38.032 30.576 ;
  LAYER M3 ;
        RECT 35.536 27.972 38.032 30.576 ;
  LAYER M2 ;
        RECT 35.536 27.972 38.032 30.576 ;
  LAYER M1 ;
        RECT 35.536 24.864 38.032 27.468 ;
  LAYER M3 ;
        RECT 35.536 24.864 38.032 27.468 ;
  LAYER M2 ;
        RECT 35.536 24.864 38.032 27.468 ;
  LAYER M1 ;
        RECT 35.536 21.756 38.032 24.36 ;
  LAYER M3 ;
        RECT 35.536 21.756 38.032 24.36 ;
  LAYER M2 ;
        RECT 35.536 21.756 38.032 24.36 ;
  LAYER M1 ;
        RECT 35.536 18.648 38.032 21.252 ;
  LAYER M3 ;
        RECT 35.536 18.648 38.032 21.252 ;
  LAYER M2 ;
        RECT 35.536 18.648 38.032 21.252 ;
  LAYER M1 ;
        RECT 35.536 15.54 38.032 18.144 ;
  LAYER M3 ;
        RECT 35.536 15.54 38.032 18.144 ;
  LAYER M2 ;
        RECT 35.536 15.54 38.032 18.144 ;
  LAYER M1 ;
        RECT 38.512 27.972 41.008 30.576 ;
  LAYER M3 ;
        RECT 38.512 27.972 41.008 30.576 ;
  LAYER M2 ;
        RECT 38.512 27.972 41.008 30.576 ;
  LAYER M1 ;
        RECT 38.512 24.864 41.008 27.468 ;
  LAYER M3 ;
        RECT 38.512 24.864 41.008 27.468 ;
  LAYER M2 ;
        RECT 38.512 24.864 41.008 27.468 ;
  LAYER M1 ;
        RECT 38.512 21.756 41.008 24.36 ;
  LAYER M3 ;
        RECT 38.512 21.756 41.008 24.36 ;
  LAYER M2 ;
        RECT 38.512 21.756 41.008 24.36 ;
  LAYER M1 ;
        RECT 38.512 18.648 41.008 21.252 ;
  LAYER M3 ;
        RECT 38.512 18.648 41.008 21.252 ;
  LAYER M2 ;
        RECT 38.512 18.648 41.008 21.252 ;
  LAYER M1 ;
        RECT 38.512 15.54 41.008 18.144 ;
  LAYER M3 ;
        RECT 38.512 15.54 41.008 18.144 ;
  LAYER M2 ;
        RECT 38.512 15.54 41.008 18.144 ;
  LAYER M1 ;
        RECT 41.488 27.972 43.984 30.576 ;
  LAYER M3 ;
        RECT 41.488 27.972 43.984 30.576 ;
  LAYER M2 ;
        RECT 41.488 27.972 43.984 30.576 ;
  LAYER M1 ;
        RECT 41.488 24.864 43.984 27.468 ;
  LAYER M3 ;
        RECT 41.488 24.864 43.984 27.468 ;
  LAYER M2 ;
        RECT 41.488 24.864 43.984 27.468 ;
  LAYER M1 ;
        RECT 41.488 21.756 43.984 24.36 ;
  LAYER M3 ;
        RECT 41.488 21.756 43.984 24.36 ;
  LAYER M2 ;
        RECT 41.488 21.756 43.984 24.36 ;
  LAYER M1 ;
        RECT 41.488 18.648 43.984 21.252 ;
  LAYER M3 ;
        RECT 41.488 18.648 43.984 21.252 ;
  LAYER M2 ;
        RECT 41.488 18.648 43.984 21.252 ;
  LAYER M1 ;
        RECT 41.488 15.54 43.984 18.144 ;
  LAYER M3 ;
        RECT 41.488 15.54 43.984 18.144 ;
  LAYER M2 ;
        RECT 41.488 15.54 43.984 18.144 ;
  LAYER M1 ;
        RECT 44.464 27.972 46.96 30.576 ;
  LAYER M3 ;
        RECT 44.464 27.972 46.96 30.576 ;
  LAYER M2 ;
        RECT 44.464 27.972 46.96 30.576 ;
  LAYER M1 ;
        RECT 44.464 24.864 46.96 27.468 ;
  LAYER M3 ;
        RECT 44.464 24.864 46.96 27.468 ;
  LAYER M2 ;
        RECT 44.464 24.864 46.96 27.468 ;
  LAYER M1 ;
        RECT 44.464 21.756 46.96 24.36 ;
  LAYER M3 ;
        RECT 44.464 21.756 46.96 24.36 ;
  LAYER M2 ;
        RECT 44.464 21.756 46.96 24.36 ;
  LAYER M1 ;
        RECT 44.464 18.648 46.96 21.252 ;
  LAYER M3 ;
        RECT 44.464 18.648 46.96 21.252 ;
  LAYER M2 ;
        RECT 44.464 18.648 46.96 21.252 ;
  LAYER M1 ;
        RECT 44.464 15.54 46.96 18.144 ;
  LAYER M3 ;
        RECT 44.464 15.54 46.96 18.144 ;
  LAYER M2 ;
        RECT 44.464 15.54 46.96 18.144 ;
  LAYER M1 ;
        RECT 22.56 12.816 22.592 12.888 ;
  LAYER M2 ;
        RECT 22.54 12.836 22.612 12.868 ;
  LAYER M2 ;
        RECT 22.576 12.836 25.328 12.868 ;
  LAYER M1 ;
        RECT 25.312 12.816 25.344 12.888 ;
  LAYER M2 ;
        RECT 25.292 12.836 25.364 12.868 ;
  LAYER M1 ;
        RECT 25.536 9.708 25.568 9.78 ;
  LAYER M2 ;
        RECT 25.516 9.728 25.588 9.76 ;
  LAYER M1 ;
        RECT 25.536 9.576 25.568 9.744 ;
  LAYER M1 ;
        RECT 25.536 9.54 25.568 9.612 ;
  LAYER M2 ;
        RECT 25.516 9.56 25.588 9.592 ;
  LAYER M2 ;
        RECT 25.328 9.56 25.552 9.592 ;
  LAYER M1 ;
        RECT 25.312 9.54 25.344 9.612 ;
  LAYER M2 ;
        RECT 25.292 9.56 25.364 9.592 ;
  LAYER M1 ;
        RECT 25.312 6.012 25.344 6.084 ;
  LAYER M2 ;
        RECT 25.292 6.032 25.364 6.064 ;
  LAYER M1 ;
        RECT 25.312 6.048 25.344 6.3 ;
  LAYER M1 ;
        RECT 25.312 6.3 25.344 12.852 ;
  LAYER M1 ;
        RECT 19.584 12.816 19.616 12.888 ;
  LAYER M2 ;
        RECT 19.564 12.836 19.636 12.868 ;
  LAYER M2 ;
        RECT 19.6 12.836 22.352 12.868 ;
  LAYER M1 ;
        RECT 22.336 12.816 22.368 12.888 ;
  LAYER M2 ;
        RECT 22.316 12.836 22.388 12.868 ;
  LAYER M1 ;
        RECT 22.336 6.012 22.368 6.084 ;
  LAYER M2 ;
        RECT 22.316 6.032 22.388 6.064 ;
  LAYER M1 ;
        RECT 22.336 6.048 22.368 6.3 ;
  LAYER M1 ;
        RECT 22.336 6.3 22.368 12.852 ;
  LAYER M2 ;
        RECT 22.352 6.032 25.328 6.064 ;
  LAYER M1 ;
        RECT 25.536 12.816 25.568 12.888 ;
  LAYER M2 ;
        RECT 25.516 12.836 25.588 12.868 ;
  LAYER M2 ;
        RECT 25.552 12.836 28.304 12.868 ;
  LAYER M1 ;
        RECT 28.288 12.816 28.32 12.888 ;
  LAYER M2 ;
        RECT 28.268 12.836 28.34 12.868 ;
  LAYER M1 ;
        RECT 28.288 5.844 28.32 5.916 ;
  LAYER M2 ;
        RECT 28.268 5.864 28.34 5.896 ;
  LAYER M1 ;
        RECT 28.288 5.88 28.32 6.3 ;
  LAYER M1 ;
        RECT 28.288 6.3 28.32 12.852 ;
  LAYER M1 ;
        RECT 19.584 9.708 19.616 9.78 ;
  LAYER M2 ;
        RECT 19.564 9.728 19.636 9.76 ;
  LAYER M1 ;
        RECT 19.584 9.576 19.616 9.744 ;
  LAYER M1 ;
        RECT 19.584 9.54 19.616 9.612 ;
  LAYER M2 ;
        RECT 19.564 9.56 19.636 9.592 ;
  LAYER M2 ;
        RECT 19.376 9.56 19.6 9.592 ;
  LAYER M1 ;
        RECT 19.36 9.54 19.392 9.612 ;
  LAYER M2 ;
        RECT 19.34 9.56 19.412 9.592 ;
  LAYER M1 ;
        RECT 19.36 5.844 19.392 5.916 ;
  LAYER M2 ;
        RECT 19.34 5.864 19.412 5.896 ;
  LAYER M1 ;
        RECT 19.36 5.88 19.392 6.3 ;
  LAYER M1 ;
        RECT 19.36 6.3 19.392 9.576 ;
  LAYER M2 ;
        RECT 19.376 5.864 28.304 5.896 ;
  LAYER M1 ;
        RECT 22.56 9.708 22.592 9.78 ;
  LAYER M2 ;
        RECT 22.54 9.728 22.612 9.76 ;
  LAYER M2 ;
        RECT 19.6 9.728 22.576 9.76 ;
  LAYER M1 ;
        RECT 19.584 9.708 19.616 9.78 ;
  LAYER M2 ;
        RECT 19.564 9.728 19.636 9.76 ;
  LAYER M1 ;
        RECT 28.512 6.6 28.544 6.672 ;
  LAYER M2 ;
        RECT 28.492 6.62 28.564 6.652 ;
  LAYER M2 ;
        RECT 28.528 6.62 31.28 6.652 ;
  LAYER M1 ;
        RECT 31.264 6.6 31.296 6.672 ;
  LAYER M2 ;
        RECT 31.244 6.62 31.316 6.652 ;
  LAYER M1 ;
        RECT 28.512 9.708 28.544 9.78 ;
  LAYER M2 ;
        RECT 28.492 9.728 28.564 9.76 ;
  LAYER M2 ;
        RECT 28.528 9.728 31.28 9.76 ;
  LAYER M1 ;
        RECT 31.264 9.708 31.296 9.78 ;
  LAYER M2 ;
        RECT 31.244 9.728 31.316 9.76 ;
  LAYER M1 ;
        RECT 28.512 12.816 28.544 12.888 ;
  LAYER M2 ;
        RECT 28.492 12.836 28.564 12.868 ;
  LAYER M2 ;
        RECT 28.528 12.836 31.28 12.868 ;
  LAYER M1 ;
        RECT 31.264 12.816 31.296 12.888 ;
  LAYER M2 ;
        RECT 31.244 12.836 31.316 12.868 ;
  LAYER M1 ;
        RECT 28.512 15.924 28.544 15.996 ;
  LAYER M2 ;
        RECT 28.492 15.944 28.564 15.976 ;
  LAYER M2 ;
        RECT 28.528 15.944 31.28 15.976 ;
  LAYER M1 ;
        RECT 31.264 15.924 31.296 15.996 ;
  LAYER M2 ;
        RECT 31.244 15.944 31.316 15.976 ;
  LAYER M1 ;
        RECT 31.264 5.676 31.296 5.748 ;
  LAYER M2 ;
        RECT 31.244 5.696 31.316 5.728 ;
  LAYER M1 ;
        RECT 31.264 5.712 31.296 6.3 ;
  LAYER M1 ;
        RECT 31.264 6.3 31.296 15.96 ;
  LAYER M1 ;
        RECT 16.608 6.6 16.64 6.672 ;
  LAYER M2 ;
        RECT 16.588 6.62 16.66 6.652 ;
  LAYER M1 ;
        RECT 16.608 6.468 16.64 6.636 ;
  LAYER M1 ;
        RECT 16.608 6.432 16.64 6.504 ;
  LAYER M2 ;
        RECT 16.588 6.452 16.66 6.484 ;
  LAYER M2 ;
        RECT 16.4 6.452 16.624 6.484 ;
  LAYER M1 ;
        RECT 16.384 6.432 16.416 6.504 ;
  LAYER M2 ;
        RECT 16.364 6.452 16.436 6.484 ;
  LAYER M1 ;
        RECT 16.608 9.708 16.64 9.78 ;
  LAYER M2 ;
        RECT 16.588 9.728 16.66 9.76 ;
  LAYER M1 ;
        RECT 16.608 9.576 16.64 9.744 ;
  LAYER M1 ;
        RECT 16.608 9.54 16.64 9.612 ;
  LAYER M2 ;
        RECT 16.588 9.56 16.66 9.592 ;
  LAYER M2 ;
        RECT 16.4 9.56 16.624 9.592 ;
  LAYER M1 ;
        RECT 16.384 9.54 16.416 9.612 ;
  LAYER M2 ;
        RECT 16.364 9.56 16.436 9.592 ;
  LAYER M1 ;
        RECT 16.608 12.816 16.64 12.888 ;
  LAYER M2 ;
        RECT 16.588 12.836 16.66 12.868 ;
  LAYER M1 ;
        RECT 16.608 12.684 16.64 12.852 ;
  LAYER M1 ;
        RECT 16.608 12.648 16.64 12.72 ;
  LAYER M2 ;
        RECT 16.588 12.668 16.66 12.7 ;
  LAYER M2 ;
        RECT 16.4 12.668 16.624 12.7 ;
  LAYER M1 ;
        RECT 16.384 12.648 16.416 12.72 ;
  LAYER M2 ;
        RECT 16.364 12.668 16.436 12.7 ;
  LAYER M1 ;
        RECT 16.608 15.924 16.64 15.996 ;
  LAYER M2 ;
        RECT 16.588 15.944 16.66 15.976 ;
  LAYER M1 ;
        RECT 16.608 15.792 16.64 15.96 ;
  LAYER M1 ;
        RECT 16.608 15.756 16.64 15.828 ;
  LAYER M2 ;
        RECT 16.588 15.776 16.66 15.808 ;
  LAYER M2 ;
        RECT 16.4 15.776 16.624 15.808 ;
  LAYER M1 ;
        RECT 16.384 15.756 16.416 15.828 ;
  LAYER M2 ;
        RECT 16.364 15.776 16.436 15.808 ;
  LAYER M1 ;
        RECT 16.384 5.676 16.416 5.748 ;
  LAYER M2 ;
        RECT 16.364 5.696 16.436 5.728 ;
  LAYER M1 ;
        RECT 16.384 5.712 16.416 6.3 ;
  LAYER M1 ;
        RECT 16.384 6.3 16.416 15.792 ;
  LAYER M2 ;
        RECT 16.4 5.696 31.28 5.728 ;
  LAYER M1 ;
        RECT 25.536 6.6 25.568 6.672 ;
  LAYER M2 ;
        RECT 25.516 6.62 25.588 6.652 ;
  LAYER M2 ;
        RECT 25.552 6.62 28.528 6.652 ;
  LAYER M1 ;
        RECT 28.512 6.6 28.544 6.672 ;
  LAYER M2 ;
        RECT 28.492 6.62 28.564 6.652 ;
  LAYER M1 ;
        RECT 25.536 15.924 25.568 15.996 ;
  LAYER M2 ;
        RECT 25.516 15.944 25.588 15.976 ;
  LAYER M2 ;
        RECT 25.552 15.944 28.528 15.976 ;
  LAYER M1 ;
        RECT 28.512 15.924 28.544 15.996 ;
  LAYER M2 ;
        RECT 28.492 15.944 28.564 15.976 ;
  LAYER M1 ;
        RECT 22.56 15.924 22.592 15.996 ;
  LAYER M2 ;
        RECT 22.54 15.944 22.612 15.976 ;
  LAYER M2 ;
        RECT 22.576 15.944 25.552 15.976 ;
  LAYER M1 ;
        RECT 25.536 15.924 25.568 15.996 ;
  LAYER M2 ;
        RECT 25.516 15.944 25.588 15.976 ;
  LAYER M1 ;
        RECT 19.584 15.924 19.616 15.996 ;
  LAYER M2 ;
        RECT 19.564 15.944 19.636 15.976 ;
  LAYER M2 ;
        RECT 19.6 15.944 22.576 15.976 ;
  LAYER M1 ;
        RECT 22.56 15.924 22.592 15.996 ;
  LAYER M2 ;
        RECT 22.54 15.944 22.612 15.976 ;
  LAYER M1 ;
        RECT 19.584 6.6 19.616 6.672 ;
  LAYER M2 ;
        RECT 19.564 6.62 19.636 6.652 ;
  LAYER M2 ;
        RECT 16.624 6.62 19.6 6.652 ;
  LAYER M1 ;
        RECT 16.608 6.6 16.64 6.672 ;
  LAYER M2 ;
        RECT 16.588 6.62 16.66 6.652 ;
  LAYER M1 ;
        RECT 22.56 6.6 22.592 6.672 ;
  LAYER M2 ;
        RECT 22.54 6.62 22.612 6.652 ;
  LAYER M2 ;
        RECT 19.6 6.62 22.576 6.652 ;
  LAYER M1 ;
        RECT 19.584 6.6 19.616 6.672 ;
  LAYER M2 ;
        RECT 19.564 6.62 19.636 6.652 ;
  LAYER M1 ;
        RECT 24.928 15.252 24.96 15.324 ;
  LAYER M2 ;
        RECT 24.908 15.272 24.98 15.304 ;
  LAYER M2 ;
        RECT 24.944 15.272 25.168 15.304 ;
  LAYER M1 ;
        RECT 25.152 15.252 25.184 15.324 ;
  LAYER M2 ;
        RECT 25.132 15.272 25.204 15.304 ;
  LAYER M1 ;
        RECT 27.904 12.144 27.936 12.216 ;
  LAYER M2 ;
        RECT 27.884 12.164 27.956 12.196 ;
  LAYER M1 ;
        RECT 25.168 12.164 27.92 12.196 ;
  LAYER M1 ;
        RECT 25.152 12.144 25.184 12.216 ;
  LAYER M2 ;
        RECT 25.132 12.164 25.204 12.196 ;
  LAYER M2 ;
        RECT 25.104 12.164 25.168 12.196 ;
  LAYER M1 ;
        RECT 25.088 12.144 25.12 12.216 ;
  LAYER M2 ;
        RECT 25.068 12.164 25.14 12.196 ;
  LAYER M1 ;
        RECT 25.088 18.948 25.12 19.02 ;
  LAYER M2 ;
        RECT 25.068 18.968 25.14 19 ;
  LAYER M1 ;
        RECT 25.088 18.732 25.12 18.984 ;
  LAYER M1 ;
        RECT 25.088 12.348 25.12 18.732 ;
  LAYER M1 ;
        RECT 21.952 15.252 21.984 15.324 ;
  LAYER M2 ;
        RECT 21.932 15.272 22.004 15.304 ;
  LAYER M2 ;
        RECT 21.968 15.272 22.192 15.304 ;
  LAYER M1 ;
        RECT 22.176 15.252 22.208 15.324 ;
  LAYER M2 ;
        RECT 22.156 15.272 22.228 15.304 ;
  LAYER M1 ;
        RECT 22.176 18.948 22.208 19.02 ;
  LAYER M2 ;
        RECT 22.156 18.968 22.228 19 ;
  LAYER M1 ;
        RECT 22.176 18.732 22.208 18.984 ;
  LAYER M1 ;
        RECT 22.176 15.288 22.208 18.732 ;
  LAYER M2 ;
        RECT 22.192 18.968 25.104 19 ;
  LAYER M1 ;
        RECT 27.904 15.252 27.936 15.324 ;
  LAYER M2 ;
        RECT 27.884 15.272 27.956 15.304 ;
  LAYER M2 ;
        RECT 27.92 15.272 28.144 15.304 ;
  LAYER M1 ;
        RECT 28.128 15.252 28.16 15.324 ;
  LAYER M2 ;
        RECT 28.108 15.272 28.18 15.304 ;
  LAYER M1 ;
        RECT 28.128 19.116 28.16 19.188 ;
  LAYER M2 ;
        RECT 28.108 19.136 28.18 19.168 ;
  LAYER M1 ;
        RECT 28.128 18.732 28.16 19.152 ;
  LAYER M1 ;
        RECT 28.128 15.288 28.16 18.732 ;
  LAYER M1 ;
        RECT 21.952 12.144 21.984 12.216 ;
  LAYER M2 ;
        RECT 21.932 12.164 22.004 12.196 ;
  LAYER M1 ;
        RECT 19.216 12.164 21.968 12.196 ;
  LAYER M1 ;
        RECT 19.2 12.144 19.232 12.216 ;
  LAYER M2 ;
        RECT 19.18 12.164 19.252 12.196 ;
  LAYER M2 ;
        RECT 19.152 12.164 19.216 12.196 ;
  LAYER M1 ;
        RECT 19.136 12.144 19.168 12.216 ;
  LAYER M2 ;
        RECT 19.116 12.164 19.188 12.196 ;
  LAYER M1 ;
        RECT 19.136 19.116 19.168 19.188 ;
  LAYER M2 ;
        RECT 19.116 19.136 19.188 19.168 ;
  LAYER M1 ;
        RECT 19.136 18.732 19.168 19.152 ;
  LAYER M1 ;
        RECT 19.136 12.348 19.168 18.732 ;
  LAYER M2 ;
        RECT 19.152 19.136 28.144 19.168 ;
  LAYER M1 ;
        RECT 24.928 12.144 24.96 12.216 ;
  LAYER M2 ;
        RECT 24.908 12.164 24.98 12.196 ;
  LAYER M2 ;
        RECT 21.968 12.164 24.944 12.196 ;
  LAYER M1 ;
        RECT 21.952 12.144 21.984 12.216 ;
  LAYER M2 ;
        RECT 21.932 12.164 22.004 12.196 ;
  LAYER M1 ;
        RECT 30.88 9.036 30.912 9.108 ;
  LAYER M2 ;
        RECT 30.86 9.056 30.932 9.088 ;
  LAYER M2 ;
        RECT 30.896 9.056 31.12 9.088 ;
  LAYER M1 ;
        RECT 31.104 9.036 31.136 9.108 ;
  LAYER M2 ;
        RECT 31.084 9.056 31.156 9.088 ;
  LAYER M1 ;
        RECT 30.88 12.144 30.912 12.216 ;
  LAYER M2 ;
        RECT 30.86 12.164 30.932 12.196 ;
  LAYER M2 ;
        RECT 30.896 12.164 31.12 12.196 ;
  LAYER M1 ;
        RECT 31.104 12.144 31.136 12.216 ;
  LAYER M2 ;
        RECT 31.084 12.164 31.156 12.196 ;
  LAYER M1 ;
        RECT 30.88 15.252 30.912 15.324 ;
  LAYER M2 ;
        RECT 30.86 15.272 30.932 15.304 ;
  LAYER M2 ;
        RECT 30.896 15.272 31.12 15.304 ;
  LAYER M1 ;
        RECT 31.104 15.252 31.136 15.324 ;
  LAYER M2 ;
        RECT 31.084 15.272 31.156 15.304 ;
  LAYER M1 ;
        RECT 30.88 18.36 30.912 18.432 ;
  LAYER M2 ;
        RECT 30.86 18.38 30.932 18.412 ;
  LAYER M2 ;
        RECT 30.896 18.38 31.12 18.412 ;
  LAYER M1 ;
        RECT 31.104 18.36 31.136 18.432 ;
  LAYER M2 ;
        RECT 31.084 18.38 31.156 18.412 ;
  LAYER M1 ;
        RECT 31.104 19.284 31.136 19.356 ;
  LAYER M2 ;
        RECT 31.084 19.304 31.156 19.336 ;
  LAYER M1 ;
        RECT 31.104 18.732 31.136 19.32 ;
  LAYER M1 ;
        RECT 31.104 9.072 31.136 18.732 ;
  LAYER M1 ;
        RECT 18.976 9.036 19.008 9.108 ;
  LAYER M2 ;
        RECT 18.956 9.056 19.028 9.088 ;
  LAYER M1 ;
        RECT 16.24 9.056 18.992 9.088 ;
  LAYER M1 ;
        RECT 16.224 9.036 16.256 9.108 ;
  LAYER M2 ;
        RECT 16.204 9.056 16.276 9.088 ;
  LAYER M2 ;
        RECT 16.176 9.056 16.24 9.088 ;
  LAYER M1 ;
        RECT 16.16 9.036 16.192 9.108 ;
  LAYER M2 ;
        RECT 16.14 9.056 16.212 9.088 ;
  LAYER M1 ;
        RECT 18.976 12.144 19.008 12.216 ;
  LAYER M2 ;
        RECT 18.956 12.164 19.028 12.196 ;
  LAYER M1 ;
        RECT 16.24 12.164 18.992 12.196 ;
  LAYER M1 ;
        RECT 16.224 12.144 16.256 12.216 ;
  LAYER M2 ;
        RECT 16.204 12.164 16.276 12.196 ;
  LAYER M2 ;
        RECT 16.176 12.164 16.24 12.196 ;
  LAYER M1 ;
        RECT 16.16 12.144 16.192 12.216 ;
  LAYER M2 ;
        RECT 16.14 12.164 16.212 12.196 ;
  LAYER M1 ;
        RECT 18.976 15.252 19.008 15.324 ;
  LAYER M2 ;
        RECT 18.956 15.272 19.028 15.304 ;
  LAYER M1 ;
        RECT 16.24 15.272 18.992 15.304 ;
  LAYER M1 ;
        RECT 16.224 15.252 16.256 15.324 ;
  LAYER M2 ;
        RECT 16.204 15.272 16.276 15.304 ;
  LAYER M2 ;
        RECT 16.176 15.272 16.24 15.304 ;
  LAYER M1 ;
        RECT 16.16 15.252 16.192 15.324 ;
  LAYER M2 ;
        RECT 16.14 15.272 16.212 15.304 ;
  LAYER M1 ;
        RECT 18.976 18.36 19.008 18.432 ;
  LAYER M2 ;
        RECT 18.956 18.38 19.028 18.412 ;
  LAYER M1 ;
        RECT 16.24 18.38 18.992 18.412 ;
  LAYER M1 ;
        RECT 16.224 18.36 16.256 18.432 ;
  LAYER M2 ;
        RECT 16.204 18.38 16.276 18.412 ;
  LAYER M2 ;
        RECT 16.176 18.38 16.24 18.412 ;
  LAYER M1 ;
        RECT 16.16 18.36 16.192 18.432 ;
  LAYER M2 ;
        RECT 16.14 18.38 16.212 18.412 ;
  LAYER M1 ;
        RECT 16.16 19.284 16.192 19.356 ;
  LAYER M2 ;
        RECT 16.14 19.304 16.212 19.336 ;
  LAYER M1 ;
        RECT 16.16 18.732 16.192 19.32 ;
  LAYER M1 ;
        RECT 16.16 9.24 16.192 18.732 ;
  LAYER M2 ;
        RECT 16.176 19.304 31.12 19.336 ;
  LAYER M1 ;
        RECT 27.904 9.036 27.936 9.108 ;
  LAYER M2 ;
        RECT 27.884 9.056 27.956 9.088 ;
  LAYER M2 ;
        RECT 27.92 9.056 30.896 9.088 ;
  LAYER M1 ;
        RECT 30.88 9.036 30.912 9.108 ;
  LAYER M2 ;
        RECT 30.86 9.056 30.932 9.088 ;
  LAYER M1 ;
        RECT 27.904 18.36 27.936 18.432 ;
  LAYER M2 ;
        RECT 27.884 18.38 27.956 18.412 ;
  LAYER M2 ;
        RECT 27.92 18.38 30.896 18.412 ;
  LAYER M1 ;
        RECT 30.88 18.36 30.912 18.432 ;
  LAYER M2 ;
        RECT 30.86 18.38 30.932 18.412 ;
  LAYER M1 ;
        RECT 24.928 18.36 24.96 18.432 ;
  LAYER M2 ;
        RECT 24.908 18.38 24.98 18.412 ;
  LAYER M2 ;
        RECT 24.944 18.38 27.92 18.412 ;
  LAYER M1 ;
        RECT 27.904 18.36 27.936 18.432 ;
  LAYER M2 ;
        RECT 27.884 18.38 27.956 18.412 ;
  LAYER M1 ;
        RECT 21.952 18.36 21.984 18.432 ;
  LAYER M2 ;
        RECT 21.932 18.38 22.004 18.412 ;
  LAYER M2 ;
        RECT 21.968 18.38 24.944 18.412 ;
  LAYER M1 ;
        RECT 24.928 18.36 24.96 18.432 ;
  LAYER M2 ;
        RECT 24.908 18.38 24.98 18.412 ;
  LAYER M1 ;
        RECT 21.952 9.036 21.984 9.108 ;
  LAYER M2 ;
        RECT 21.932 9.056 22.004 9.088 ;
  LAYER M2 ;
        RECT 18.992 9.056 21.968 9.088 ;
  LAYER M1 ;
        RECT 18.976 9.036 19.008 9.108 ;
  LAYER M2 ;
        RECT 18.956 9.056 19.028 9.088 ;
  LAYER M1 ;
        RECT 24.928 9.036 24.96 9.108 ;
  LAYER M2 ;
        RECT 24.908 9.056 24.98 9.088 ;
  LAYER M2 ;
        RECT 21.968 9.056 24.944 9.088 ;
  LAYER M1 ;
        RECT 21.952 9.036 21.984 9.108 ;
  LAYER M2 ;
        RECT 21.932 9.056 22.004 9.088 ;
  LAYER M1 ;
        RECT 28.464 6.552 30.96 9.156 ;
  LAYER M3 ;
        RECT 28.464 6.552 30.96 9.156 ;
  LAYER M2 ;
        RECT 28.464 6.552 30.96 9.156 ;
  LAYER M1 ;
        RECT 28.464 9.66 30.96 12.264 ;
  LAYER M3 ;
        RECT 28.464 9.66 30.96 12.264 ;
  LAYER M2 ;
        RECT 28.464 9.66 30.96 12.264 ;
  LAYER M1 ;
        RECT 28.464 12.768 30.96 15.372 ;
  LAYER M3 ;
        RECT 28.464 12.768 30.96 15.372 ;
  LAYER M2 ;
        RECT 28.464 12.768 30.96 15.372 ;
  LAYER M1 ;
        RECT 28.464 15.876 30.96 18.48 ;
  LAYER M3 ;
        RECT 28.464 15.876 30.96 18.48 ;
  LAYER M2 ;
        RECT 28.464 15.876 30.96 18.48 ;
  LAYER M1 ;
        RECT 25.488 6.552 27.984 9.156 ;
  LAYER M3 ;
        RECT 25.488 6.552 27.984 9.156 ;
  LAYER M2 ;
        RECT 25.488 6.552 27.984 9.156 ;
  LAYER M1 ;
        RECT 25.488 9.66 27.984 12.264 ;
  LAYER M3 ;
        RECT 25.488 9.66 27.984 12.264 ;
  LAYER M2 ;
        RECT 25.488 9.66 27.984 12.264 ;
  LAYER M1 ;
        RECT 25.488 12.768 27.984 15.372 ;
  LAYER M3 ;
        RECT 25.488 12.768 27.984 15.372 ;
  LAYER M2 ;
        RECT 25.488 12.768 27.984 15.372 ;
  LAYER M1 ;
        RECT 25.488 15.876 27.984 18.48 ;
  LAYER M3 ;
        RECT 25.488 15.876 27.984 18.48 ;
  LAYER M2 ;
        RECT 25.488 15.876 27.984 18.48 ;
  LAYER M1 ;
        RECT 22.512 6.552 25.008 9.156 ;
  LAYER M3 ;
        RECT 22.512 6.552 25.008 9.156 ;
  LAYER M2 ;
        RECT 22.512 6.552 25.008 9.156 ;
  LAYER M1 ;
        RECT 22.512 9.66 25.008 12.264 ;
  LAYER M3 ;
        RECT 22.512 9.66 25.008 12.264 ;
  LAYER M2 ;
        RECT 22.512 9.66 25.008 12.264 ;
  LAYER M1 ;
        RECT 22.512 12.768 25.008 15.372 ;
  LAYER M3 ;
        RECT 22.512 12.768 25.008 15.372 ;
  LAYER M2 ;
        RECT 22.512 12.768 25.008 15.372 ;
  LAYER M1 ;
        RECT 22.512 15.876 25.008 18.48 ;
  LAYER M3 ;
        RECT 22.512 15.876 25.008 18.48 ;
  LAYER M2 ;
        RECT 22.512 15.876 25.008 18.48 ;
  LAYER M1 ;
        RECT 19.536 6.552 22.032 9.156 ;
  LAYER M3 ;
        RECT 19.536 6.552 22.032 9.156 ;
  LAYER M2 ;
        RECT 19.536 6.552 22.032 9.156 ;
  LAYER M1 ;
        RECT 19.536 9.66 22.032 12.264 ;
  LAYER M3 ;
        RECT 19.536 9.66 22.032 12.264 ;
  LAYER M2 ;
        RECT 19.536 9.66 22.032 12.264 ;
  LAYER M1 ;
        RECT 19.536 12.768 22.032 15.372 ;
  LAYER M3 ;
        RECT 19.536 12.768 22.032 15.372 ;
  LAYER M2 ;
        RECT 19.536 12.768 22.032 15.372 ;
  LAYER M1 ;
        RECT 19.536 15.876 22.032 18.48 ;
  LAYER M3 ;
        RECT 19.536 15.876 22.032 18.48 ;
  LAYER M2 ;
        RECT 19.536 15.876 22.032 18.48 ;
  LAYER M1 ;
        RECT 16.56 6.552 19.056 9.156 ;
  LAYER M3 ;
        RECT 16.56 6.552 19.056 9.156 ;
  LAYER M2 ;
        RECT 16.56 6.552 19.056 9.156 ;
  LAYER M1 ;
        RECT 16.56 9.66 19.056 12.264 ;
  LAYER M3 ;
        RECT 16.56 9.66 19.056 12.264 ;
  LAYER M2 ;
        RECT 16.56 9.66 19.056 12.264 ;
  LAYER M1 ;
        RECT 16.56 12.768 19.056 15.372 ;
  LAYER M3 ;
        RECT 16.56 12.768 19.056 15.372 ;
  LAYER M2 ;
        RECT 16.56 12.768 19.056 15.372 ;
  LAYER M1 ;
        RECT 16.56 15.876 19.056 18.48 ;
  LAYER M3 ;
        RECT 16.56 15.876 19.056 18.48 ;
  LAYER M2 ;
        RECT 16.56 15.876 19.056 18.48 ;
  LAYER M1 ;
        RECT 24.928 32.22 24.96 32.292 ;
  LAYER M2 ;
        RECT 24.908 32.24 24.98 32.272 ;
  LAYER M2 ;
        RECT 22.192 32.24 24.944 32.272 ;
  LAYER M1 ;
        RECT 22.176 32.22 22.208 32.292 ;
  LAYER M2 ;
        RECT 22.156 32.24 22.228 32.272 ;
  LAYER M1 ;
        RECT 24.928 29.112 24.96 29.184 ;
  LAYER M2 ;
        RECT 24.908 29.132 24.98 29.164 ;
  LAYER M2 ;
        RECT 22.192 29.132 24.944 29.164 ;
  LAYER M1 ;
        RECT 22.176 29.112 22.208 29.184 ;
  LAYER M2 ;
        RECT 22.156 29.132 22.228 29.164 ;
  LAYER M1 ;
        RECT 21.952 32.22 21.984 32.292 ;
  LAYER M2 ;
        RECT 21.932 32.24 22.004 32.272 ;
  LAYER M1 ;
        RECT 21.952 32.256 21.984 32.424 ;
  LAYER M1 ;
        RECT 21.952 32.388 21.984 32.46 ;
  LAYER M2 ;
        RECT 21.932 32.408 22.004 32.44 ;
  LAYER M2 ;
        RECT 21.968 32.408 22.192 32.44 ;
  LAYER M1 ;
        RECT 22.176 32.388 22.208 32.46 ;
  LAYER M2 ;
        RECT 22.156 32.408 22.228 32.44 ;
  LAYER M1 ;
        RECT 21.952 29.112 21.984 29.184 ;
  LAYER M2 ;
        RECT 21.932 29.132 22.004 29.164 ;
  LAYER M1 ;
        RECT 21.952 29.148 21.984 29.316 ;
  LAYER M1 ;
        RECT 21.952 29.28 21.984 29.352 ;
  LAYER M2 ;
        RECT 21.932 29.3 22.004 29.332 ;
  LAYER M2 ;
        RECT 21.968 29.3 22.192 29.332 ;
  LAYER M1 ;
        RECT 22.176 29.28 22.208 29.352 ;
  LAYER M2 ;
        RECT 22.156 29.3 22.228 29.332 ;
  LAYER M1 ;
        RECT 22.176 39.024 22.208 39.096 ;
  LAYER M2 ;
        RECT 22.156 39.044 22.228 39.076 ;
  LAYER M1 ;
        RECT 22.176 38.808 22.208 39.06 ;
  LAYER M1 ;
        RECT 22.176 29.148 22.208 38.808 ;
  LAYER M1 ;
        RECT 27.904 29.112 27.936 29.184 ;
  LAYER M2 ;
        RECT 27.884 29.132 27.956 29.164 ;
  LAYER M2 ;
        RECT 25.168 29.132 27.92 29.164 ;
  LAYER M1 ;
        RECT 25.152 29.112 25.184 29.184 ;
  LAYER M2 ;
        RECT 25.132 29.132 25.204 29.164 ;
  LAYER M1 ;
        RECT 27.904 32.22 27.936 32.292 ;
  LAYER M2 ;
        RECT 27.884 32.24 27.956 32.272 ;
  LAYER M2 ;
        RECT 25.168 32.24 27.92 32.272 ;
  LAYER M1 ;
        RECT 25.152 32.22 25.184 32.292 ;
  LAYER M2 ;
        RECT 25.132 32.24 25.204 32.272 ;
  LAYER M1 ;
        RECT 25.152 39.024 25.184 39.096 ;
  LAYER M2 ;
        RECT 25.132 39.044 25.204 39.076 ;
  LAYER M1 ;
        RECT 25.152 38.808 25.184 39.06 ;
  LAYER M1 ;
        RECT 25.152 29.148 25.184 38.808 ;
  LAYER M2 ;
        RECT 22.192 39.044 25.168 39.076 ;
  LAYER M1 ;
        RECT 21.952 26.004 21.984 26.076 ;
  LAYER M2 ;
        RECT 21.932 26.024 22.004 26.056 ;
  LAYER M2 ;
        RECT 19.216 26.024 21.968 26.056 ;
  LAYER M1 ;
        RECT 19.2 26.004 19.232 26.076 ;
  LAYER M2 ;
        RECT 19.18 26.024 19.252 26.056 ;
  LAYER M1 ;
        RECT 21.952 35.328 21.984 35.4 ;
  LAYER M2 ;
        RECT 21.932 35.348 22.004 35.38 ;
  LAYER M2 ;
        RECT 19.216 35.348 21.968 35.38 ;
  LAYER M1 ;
        RECT 19.2 35.328 19.232 35.4 ;
  LAYER M2 ;
        RECT 19.18 35.348 19.252 35.38 ;
  LAYER M1 ;
        RECT 19.2 39.192 19.232 39.264 ;
  LAYER M2 ;
        RECT 19.18 39.212 19.252 39.244 ;
  LAYER M1 ;
        RECT 19.2 38.808 19.232 39.228 ;
  LAYER M1 ;
        RECT 19.2 26.04 19.232 38.808 ;
  LAYER M1 ;
        RECT 27.904 35.328 27.936 35.4 ;
  LAYER M2 ;
        RECT 27.884 35.348 27.956 35.38 ;
  LAYER M1 ;
        RECT 27.904 35.364 27.936 35.532 ;
  LAYER M1 ;
        RECT 27.904 35.496 27.936 35.568 ;
  LAYER M2 ;
        RECT 27.884 35.516 27.956 35.548 ;
  LAYER M2 ;
        RECT 27.92 35.516 28.144 35.548 ;
  LAYER M1 ;
        RECT 28.128 35.496 28.16 35.568 ;
  LAYER M2 ;
        RECT 28.108 35.516 28.18 35.548 ;
  LAYER M1 ;
        RECT 27.904 26.004 27.936 26.076 ;
  LAYER M2 ;
        RECT 27.884 26.024 27.956 26.056 ;
  LAYER M1 ;
        RECT 27.904 26.04 27.936 26.208 ;
  LAYER M1 ;
        RECT 27.904 26.172 27.936 26.244 ;
  LAYER M2 ;
        RECT 27.884 26.192 27.956 26.224 ;
  LAYER M2 ;
        RECT 27.92 26.192 28.144 26.224 ;
  LAYER M1 ;
        RECT 28.128 26.172 28.16 26.244 ;
  LAYER M2 ;
        RECT 28.108 26.192 28.18 26.224 ;
  LAYER M1 ;
        RECT 28.128 39.192 28.16 39.264 ;
  LAYER M2 ;
        RECT 28.108 39.212 28.18 39.244 ;
  LAYER M1 ;
        RECT 28.128 38.808 28.16 39.228 ;
  LAYER M1 ;
        RECT 28.128 26.208 28.16 38.808 ;
  LAYER M2 ;
        RECT 19.216 39.212 28.144 39.244 ;
  LAYER M1 ;
        RECT 24.928 35.328 24.96 35.4 ;
  LAYER M2 ;
        RECT 24.908 35.348 24.98 35.38 ;
  LAYER M2 ;
        RECT 24.944 35.348 27.92 35.38 ;
  LAYER M1 ;
        RECT 27.904 35.328 27.936 35.4 ;
  LAYER M2 ;
        RECT 27.884 35.348 27.956 35.38 ;
  LAYER M1 ;
        RECT 24.928 26.004 24.96 26.076 ;
  LAYER M2 ;
        RECT 24.908 26.024 24.98 26.056 ;
  LAYER M2 ;
        RECT 21.968 26.024 24.944 26.056 ;
  LAYER M1 ;
        RECT 21.952 26.004 21.984 26.076 ;
  LAYER M2 ;
        RECT 21.932 26.024 22.004 26.056 ;
  LAYER M1 ;
        RECT 18.976 38.436 19.008 38.508 ;
  LAYER M2 ;
        RECT 18.956 38.456 19.028 38.488 ;
  LAYER M2 ;
        RECT 16.24 38.456 18.992 38.488 ;
  LAYER M1 ;
        RECT 16.224 38.436 16.256 38.508 ;
  LAYER M2 ;
        RECT 16.204 38.456 16.276 38.488 ;
  LAYER M1 ;
        RECT 18.976 35.328 19.008 35.4 ;
  LAYER M2 ;
        RECT 18.956 35.348 19.028 35.38 ;
  LAYER M2 ;
        RECT 16.24 35.348 18.992 35.38 ;
  LAYER M1 ;
        RECT 16.224 35.328 16.256 35.4 ;
  LAYER M2 ;
        RECT 16.204 35.348 16.276 35.38 ;
  LAYER M1 ;
        RECT 18.976 32.22 19.008 32.292 ;
  LAYER M2 ;
        RECT 18.956 32.24 19.028 32.272 ;
  LAYER M2 ;
        RECT 16.24 32.24 18.992 32.272 ;
  LAYER M1 ;
        RECT 16.224 32.22 16.256 32.292 ;
  LAYER M2 ;
        RECT 16.204 32.24 16.276 32.272 ;
  LAYER M1 ;
        RECT 18.976 29.112 19.008 29.184 ;
  LAYER M2 ;
        RECT 18.956 29.132 19.028 29.164 ;
  LAYER M2 ;
        RECT 16.24 29.132 18.992 29.164 ;
  LAYER M1 ;
        RECT 16.224 29.112 16.256 29.184 ;
  LAYER M2 ;
        RECT 16.204 29.132 16.276 29.164 ;
  LAYER M1 ;
        RECT 18.976 26.004 19.008 26.076 ;
  LAYER M2 ;
        RECT 18.956 26.024 19.028 26.056 ;
  LAYER M2 ;
        RECT 16.24 26.024 18.992 26.056 ;
  LAYER M1 ;
        RECT 16.224 26.004 16.256 26.076 ;
  LAYER M2 ;
        RECT 16.204 26.024 16.276 26.056 ;
  LAYER M1 ;
        RECT 18.976 22.896 19.008 22.968 ;
  LAYER M2 ;
        RECT 18.956 22.916 19.028 22.948 ;
  LAYER M2 ;
        RECT 16.24 22.916 18.992 22.948 ;
  LAYER M1 ;
        RECT 16.224 22.896 16.256 22.968 ;
  LAYER M2 ;
        RECT 16.204 22.916 16.276 22.948 ;
  LAYER M1 ;
        RECT 16.224 39.36 16.256 39.432 ;
  LAYER M2 ;
        RECT 16.204 39.38 16.276 39.412 ;
  LAYER M1 ;
        RECT 16.224 38.808 16.256 39.396 ;
  LAYER M1 ;
        RECT 16.224 22.932 16.256 38.808 ;
  LAYER M1 ;
        RECT 30.88 38.436 30.912 38.508 ;
  LAYER M2 ;
        RECT 30.86 38.456 30.932 38.488 ;
  LAYER M1 ;
        RECT 30.88 38.472 30.912 38.64 ;
  LAYER M1 ;
        RECT 30.88 38.604 30.912 38.676 ;
  LAYER M2 ;
        RECT 30.86 38.624 30.932 38.656 ;
  LAYER M2 ;
        RECT 30.896 38.624 31.12 38.656 ;
  LAYER M1 ;
        RECT 31.104 38.604 31.136 38.676 ;
  LAYER M2 ;
        RECT 31.084 38.624 31.156 38.656 ;
  LAYER M1 ;
        RECT 30.88 35.328 30.912 35.4 ;
  LAYER M2 ;
        RECT 30.86 35.348 30.932 35.38 ;
  LAYER M1 ;
        RECT 30.88 35.364 30.912 35.532 ;
  LAYER M1 ;
        RECT 30.88 35.496 30.912 35.568 ;
  LAYER M2 ;
        RECT 30.86 35.516 30.932 35.548 ;
  LAYER M2 ;
        RECT 30.896 35.516 31.12 35.548 ;
  LAYER M1 ;
        RECT 31.104 35.496 31.136 35.568 ;
  LAYER M2 ;
        RECT 31.084 35.516 31.156 35.548 ;
  LAYER M1 ;
        RECT 30.88 32.22 30.912 32.292 ;
  LAYER M2 ;
        RECT 30.86 32.24 30.932 32.272 ;
  LAYER M1 ;
        RECT 30.88 32.256 30.912 32.424 ;
  LAYER M1 ;
        RECT 30.88 32.388 30.912 32.46 ;
  LAYER M2 ;
        RECT 30.86 32.408 30.932 32.44 ;
  LAYER M2 ;
        RECT 30.896 32.408 31.12 32.44 ;
  LAYER M1 ;
        RECT 31.104 32.388 31.136 32.46 ;
  LAYER M2 ;
        RECT 31.084 32.408 31.156 32.44 ;
  LAYER M1 ;
        RECT 30.88 29.112 30.912 29.184 ;
  LAYER M2 ;
        RECT 30.86 29.132 30.932 29.164 ;
  LAYER M1 ;
        RECT 30.88 29.148 30.912 29.316 ;
  LAYER M1 ;
        RECT 30.88 29.28 30.912 29.352 ;
  LAYER M2 ;
        RECT 30.86 29.3 30.932 29.332 ;
  LAYER M2 ;
        RECT 30.896 29.3 31.12 29.332 ;
  LAYER M1 ;
        RECT 31.104 29.28 31.136 29.352 ;
  LAYER M2 ;
        RECT 31.084 29.3 31.156 29.332 ;
  LAYER M1 ;
        RECT 30.88 26.004 30.912 26.076 ;
  LAYER M2 ;
        RECT 30.86 26.024 30.932 26.056 ;
  LAYER M1 ;
        RECT 30.88 26.04 30.912 26.208 ;
  LAYER M1 ;
        RECT 30.88 26.172 30.912 26.244 ;
  LAYER M2 ;
        RECT 30.86 26.192 30.932 26.224 ;
  LAYER M2 ;
        RECT 30.896 26.192 31.12 26.224 ;
  LAYER M1 ;
        RECT 31.104 26.172 31.136 26.244 ;
  LAYER M2 ;
        RECT 31.084 26.192 31.156 26.224 ;
  LAYER M1 ;
        RECT 30.88 22.896 30.912 22.968 ;
  LAYER M2 ;
        RECT 30.86 22.916 30.932 22.948 ;
  LAYER M1 ;
        RECT 30.88 22.932 30.912 23.1 ;
  LAYER M1 ;
        RECT 30.88 23.064 30.912 23.136 ;
  LAYER M2 ;
        RECT 30.86 23.084 30.932 23.116 ;
  LAYER M2 ;
        RECT 30.896 23.084 31.12 23.116 ;
  LAYER M1 ;
        RECT 31.104 23.064 31.136 23.136 ;
  LAYER M2 ;
        RECT 31.084 23.084 31.156 23.116 ;
  LAYER M1 ;
        RECT 31.104 39.36 31.136 39.432 ;
  LAYER M2 ;
        RECT 31.084 39.38 31.156 39.412 ;
  LAYER M1 ;
        RECT 31.104 38.808 31.136 39.396 ;
  LAYER M1 ;
        RECT 31.104 23.1 31.136 38.808 ;
  LAYER M2 ;
        RECT 16.24 39.38 31.12 39.412 ;
  LAYER M1 ;
        RECT 21.952 38.436 21.984 38.508 ;
  LAYER M2 ;
        RECT 21.932 38.456 22.004 38.488 ;
  LAYER M2 ;
        RECT 18.992 38.456 21.968 38.488 ;
  LAYER M1 ;
        RECT 18.976 38.436 19.008 38.508 ;
  LAYER M2 ;
        RECT 18.956 38.456 19.028 38.488 ;
  LAYER M1 ;
        RECT 21.952 22.896 21.984 22.968 ;
  LAYER M2 ;
        RECT 21.932 22.916 22.004 22.948 ;
  LAYER M2 ;
        RECT 18.992 22.916 21.968 22.948 ;
  LAYER M1 ;
        RECT 18.976 22.896 19.008 22.968 ;
  LAYER M2 ;
        RECT 18.956 22.916 19.028 22.948 ;
  LAYER M1 ;
        RECT 24.928 22.896 24.96 22.968 ;
  LAYER M2 ;
        RECT 24.908 22.916 24.98 22.948 ;
  LAYER M2 ;
        RECT 21.968 22.916 24.944 22.948 ;
  LAYER M1 ;
        RECT 21.952 22.896 21.984 22.968 ;
  LAYER M2 ;
        RECT 21.932 22.916 22.004 22.948 ;
  LAYER M1 ;
        RECT 27.904 22.896 27.936 22.968 ;
  LAYER M2 ;
        RECT 27.884 22.916 27.956 22.948 ;
  LAYER M2 ;
        RECT 24.944 22.916 27.92 22.948 ;
  LAYER M1 ;
        RECT 24.928 22.896 24.96 22.968 ;
  LAYER M2 ;
        RECT 24.908 22.916 24.98 22.948 ;
  LAYER M1 ;
        RECT 27.904 38.436 27.936 38.508 ;
  LAYER M2 ;
        RECT 27.884 38.456 27.956 38.488 ;
  LAYER M2 ;
        RECT 27.92 38.456 30.896 38.488 ;
  LAYER M1 ;
        RECT 30.88 38.436 30.912 38.508 ;
  LAYER M2 ;
        RECT 30.86 38.456 30.932 38.488 ;
  LAYER M1 ;
        RECT 24.928 38.436 24.96 38.508 ;
  LAYER M2 ;
        RECT 24.908 38.456 24.98 38.488 ;
  LAYER M2 ;
        RECT 24.944 38.456 27.92 38.488 ;
  LAYER M1 ;
        RECT 27.904 38.436 27.936 38.508 ;
  LAYER M2 ;
        RECT 27.884 38.456 27.956 38.488 ;
  LAYER M1 ;
        RECT 22.56 29.784 22.592 29.856 ;
  LAYER M2 ;
        RECT 22.54 29.804 22.612 29.836 ;
  LAYER M2 ;
        RECT 22.352 29.804 22.576 29.836 ;
  LAYER M1 ;
        RECT 22.336 29.784 22.368 29.856 ;
  LAYER M2 ;
        RECT 22.316 29.804 22.388 29.836 ;
  LAYER M1 ;
        RECT 22.56 26.676 22.592 26.748 ;
  LAYER M2 ;
        RECT 22.54 26.696 22.612 26.728 ;
  LAYER M2 ;
        RECT 22.352 26.696 22.576 26.728 ;
  LAYER M1 ;
        RECT 22.336 26.676 22.368 26.748 ;
  LAYER M2 ;
        RECT 22.316 26.696 22.388 26.728 ;
  LAYER M1 ;
        RECT 19.584 29.784 19.616 29.856 ;
  LAYER M2 ;
        RECT 19.564 29.804 19.636 29.836 ;
  LAYER M1 ;
        RECT 19.6 29.804 22.352 29.836 ;
  LAYER M1 ;
        RECT 22.336 29.784 22.368 29.856 ;
  LAYER M2 ;
        RECT 22.316 29.804 22.388 29.836 ;
  LAYER M2 ;
        RECT 22.352 29.804 22.416 29.836 ;
  LAYER M1 ;
        RECT 22.4 29.784 22.432 29.856 ;
  LAYER M2 ;
        RECT 22.38 29.804 22.452 29.836 ;
  LAYER M1 ;
        RECT 19.584 26.676 19.616 26.748 ;
  LAYER M2 ;
        RECT 19.564 26.696 19.636 26.728 ;
  LAYER M1 ;
        RECT 19.6 26.696 22.352 26.728 ;
  LAYER M1 ;
        RECT 22.336 26.676 22.368 26.748 ;
  LAYER M2 ;
        RECT 22.316 26.696 22.388 26.728 ;
  LAYER M2 ;
        RECT 22.352 26.696 22.416 26.728 ;
  LAYER M1 ;
        RECT 22.4 26.676 22.432 26.748 ;
  LAYER M2 ;
        RECT 22.38 26.696 22.452 26.728 ;
  LAYER M1 ;
        RECT 22.4 19.872 22.432 19.944 ;
  LAYER M2 ;
        RECT 22.38 19.892 22.452 19.924 ;
  LAYER M1 ;
        RECT 22.4 19.908 22.432 20.16 ;
  LAYER M1 ;
        RECT 22.4 20.16 22.432 29.82 ;
  LAYER M1 ;
        RECT 25.536 26.676 25.568 26.748 ;
  LAYER M2 ;
        RECT 25.516 26.696 25.588 26.728 ;
  LAYER M2 ;
        RECT 25.328 26.696 25.552 26.728 ;
  LAYER M1 ;
        RECT 25.312 26.676 25.344 26.748 ;
  LAYER M2 ;
        RECT 25.292 26.696 25.364 26.728 ;
  LAYER M1 ;
        RECT 25.536 29.784 25.568 29.856 ;
  LAYER M2 ;
        RECT 25.516 29.804 25.588 29.836 ;
  LAYER M2 ;
        RECT 25.328 29.804 25.552 29.836 ;
  LAYER M1 ;
        RECT 25.312 29.784 25.344 29.856 ;
  LAYER M2 ;
        RECT 25.292 29.804 25.364 29.836 ;
  LAYER M1 ;
        RECT 25.312 19.872 25.344 19.944 ;
  LAYER M2 ;
        RECT 25.292 19.892 25.364 19.924 ;
  LAYER M1 ;
        RECT 25.312 19.908 25.344 20.16 ;
  LAYER M1 ;
        RECT 25.312 20.16 25.344 29.82 ;
  LAYER M2 ;
        RECT 22.416 19.892 25.328 19.924 ;
  LAYER M1 ;
        RECT 19.584 23.568 19.616 23.64 ;
  LAYER M2 ;
        RECT 19.564 23.588 19.636 23.62 ;
  LAYER M2 ;
        RECT 19.376 23.588 19.6 23.62 ;
  LAYER M1 ;
        RECT 19.36 23.568 19.392 23.64 ;
  LAYER M2 ;
        RECT 19.34 23.588 19.412 23.62 ;
  LAYER M1 ;
        RECT 19.584 32.892 19.616 32.964 ;
  LAYER M2 ;
        RECT 19.564 32.912 19.636 32.944 ;
  LAYER M2 ;
        RECT 19.376 32.912 19.6 32.944 ;
  LAYER M1 ;
        RECT 19.36 32.892 19.392 32.964 ;
  LAYER M2 ;
        RECT 19.34 32.912 19.412 32.944 ;
  LAYER M1 ;
        RECT 19.36 19.704 19.392 19.776 ;
  LAYER M2 ;
        RECT 19.34 19.724 19.412 19.756 ;
  LAYER M1 ;
        RECT 19.36 19.74 19.392 20.16 ;
  LAYER M1 ;
        RECT 19.36 20.16 19.392 32.928 ;
  LAYER M1 ;
        RECT 25.536 32.892 25.568 32.964 ;
  LAYER M2 ;
        RECT 25.516 32.912 25.588 32.944 ;
  LAYER M1 ;
        RECT 25.552 32.912 28.304 32.944 ;
  LAYER M1 ;
        RECT 28.288 32.892 28.32 32.964 ;
  LAYER M2 ;
        RECT 28.268 32.912 28.34 32.944 ;
  LAYER M2 ;
        RECT 28.304 32.912 28.368 32.944 ;
  LAYER M1 ;
        RECT 28.352 32.892 28.384 32.964 ;
  LAYER M2 ;
        RECT 28.332 32.912 28.404 32.944 ;
  LAYER M1 ;
        RECT 25.536 23.568 25.568 23.64 ;
  LAYER M2 ;
        RECT 25.516 23.588 25.588 23.62 ;
  LAYER M1 ;
        RECT 25.552 23.588 28.304 23.62 ;
  LAYER M1 ;
        RECT 28.288 23.568 28.32 23.64 ;
  LAYER M2 ;
        RECT 28.268 23.588 28.34 23.62 ;
  LAYER M2 ;
        RECT 28.304 23.588 28.368 23.62 ;
  LAYER M1 ;
        RECT 28.352 23.568 28.384 23.64 ;
  LAYER M2 ;
        RECT 28.332 23.588 28.404 23.62 ;
  LAYER M1 ;
        RECT 28.352 19.704 28.384 19.776 ;
  LAYER M2 ;
        RECT 28.332 19.724 28.404 19.756 ;
  LAYER M1 ;
        RECT 28.352 19.74 28.384 20.16 ;
  LAYER M1 ;
        RECT 28.352 20.16 28.384 32.76 ;
  LAYER M2 ;
        RECT 19.376 19.724 28.368 19.756 ;
  LAYER M1 ;
        RECT 22.56 32.892 22.592 32.964 ;
  LAYER M2 ;
        RECT 22.54 32.912 22.612 32.944 ;
  LAYER M2 ;
        RECT 22.576 32.912 25.552 32.944 ;
  LAYER M1 ;
        RECT 25.536 32.892 25.568 32.964 ;
  LAYER M2 ;
        RECT 25.516 32.912 25.588 32.944 ;
  LAYER M1 ;
        RECT 22.56 23.568 22.592 23.64 ;
  LAYER M2 ;
        RECT 22.54 23.588 22.612 23.62 ;
  LAYER M2 ;
        RECT 19.6 23.588 22.576 23.62 ;
  LAYER M1 ;
        RECT 19.584 23.568 19.616 23.64 ;
  LAYER M2 ;
        RECT 19.564 23.588 19.636 23.62 ;
  LAYER M1 ;
        RECT 16.608 36 16.64 36.072 ;
  LAYER M2 ;
        RECT 16.588 36.02 16.66 36.052 ;
  LAYER M2 ;
        RECT 16.4 36.02 16.624 36.052 ;
  LAYER M1 ;
        RECT 16.384 36 16.416 36.072 ;
  LAYER M2 ;
        RECT 16.364 36.02 16.436 36.052 ;
  LAYER M1 ;
        RECT 16.608 32.892 16.64 32.964 ;
  LAYER M2 ;
        RECT 16.588 32.912 16.66 32.944 ;
  LAYER M2 ;
        RECT 16.4 32.912 16.624 32.944 ;
  LAYER M1 ;
        RECT 16.384 32.892 16.416 32.964 ;
  LAYER M2 ;
        RECT 16.364 32.912 16.436 32.944 ;
  LAYER M1 ;
        RECT 16.608 29.784 16.64 29.856 ;
  LAYER M2 ;
        RECT 16.588 29.804 16.66 29.836 ;
  LAYER M2 ;
        RECT 16.4 29.804 16.624 29.836 ;
  LAYER M1 ;
        RECT 16.384 29.784 16.416 29.856 ;
  LAYER M2 ;
        RECT 16.364 29.804 16.436 29.836 ;
  LAYER M1 ;
        RECT 16.608 26.676 16.64 26.748 ;
  LAYER M2 ;
        RECT 16.588 26.696 16.66 26.728 ;
  LAYER M2 ;
        RECT 16.4 26.696 16.624 26.728 ;
  LAYER M1 ;
        RECT 16.384 26.676 16.416 26.748 ;
  LAYER M2 ;
        RECT 16.364 26.696 16.436 26.728 ;
  LAYER M1 ;
        RECT 16.608 23.568 16.64 23.64 ;
  LAYER M2 ;
        RECT 16.588 23.588 16.66 23.62 ;
  LAYER M2 ;
        RECT 16.4 23.588 16.624 23.62 ;
  LAYER M1 ;
        RECT 16.384 23.568 16.416 23.64 ;
  LAYER M2 ;
        RECT 16.364 23.588 16.436 23.62 ;
  LAYER M1 ;
        RECT 16.608 20.46 16.64 20.532 ;
  LAYER M2 ;
        RECT 16.588 20.48 16.66 20.512 ;
  LAYER M2 ;
        RECT 16.4 20.48 16.624 20.512 ;
  LAYER M1 ;
        RECT 16.384 20.46 16.416 20.532 ;
  LAYER M2 ;
        RECT 16.364 20.48 16.436 20.512 ;
  LAYER M1 ;
        RECT 16.384 19.536 16.416 19.608 ;
  LAYER M2 ;
        RECT 16.364 19.556 16.436 19.588 ;
  LAYER M1 ;
        RECT 16.384 19.572 16.416 20.16 ;
  LAYER M1 ;
        RECT 16.384 20.16 16.416 36.036 ;
  LAYER M1 ;
        RECT 28.512 36 28.544 36.072 ;
  LAYER M2 ;
        RECT 28.492 36.02 28.564 36.052 ;
  LAYER M1 ;
        RECT 28.528 36.02 31.28 36.052 ;
  LAYER M1 ;
        RECT 31.264 36 31.296 36.072 ;
  LAYER M2 ;
        RECT 31.244 36.02 31.316 36.052 ;
  LAYER M2 ;
        RECT 31.28 36.02 31.344 36.052 ;
  LAYER M1 ;
        RECT 31.328 36 31.36 36.072 ;
  LAYER M2 ;
        RECT 31.308 36.02 31.38 36.052 ;
  LAYER M1 ;
        RECT 28.512 32.892 28.544 32.964 ;
  LAYER M2 ;
        RECT 28.492 32.912 28.564 32.944 ;
  LAYER M1 ;
        RECT 28.528 32.912 31.28 32.944 ;
  LAYER M1 ;
        RECT 31.264 32.892 31.296 32.964 ;
  LAYER M2 ;
        RECT 31.244 32.912 31.316 32.944 ;
  LAYER M2 ;
        RECT 31.28 32.912 31.344 32.944 ;
  LAYER M1 ;
        RECT 31.328 32.892 31.36 32.964 ;
  LAYER M2 ;
        RECT 31.308 32.912 31.38 32.944 ;
  LAYER M1 ;
        RECT 28.512 29.784 28.544 29.856 ;
  LAYER M2 ;
        RECT 28.492 29.804 28.564 29.836 ;
  LAYER M1 ;
        RECT 28.528 29.804 31.28 29.836 ;
  LAYER M1 ;
        RECT 31.264 29.784 31.296 29.856 ;
  LAYER M2 ;
        RECT 31.244 29.804 31.316 29.836 ;
  LAYER M2 ;
        RECT 31.28 29.804 31.344 29.836 ;
  LAYER M1 ;
        RECT 31.328 29.784 31.36 29.856 ;
  LAYER M2 ;
        RECT 31.308 29.804 31.38 29.836 ;
  LAYER M1 ;
        RECT 28.512 26.676 28.544 26.748 ;
  LAYER M2 ;
        RECT 28.492 26.696 28.564 26.728 ;
  LAYER M1 ;
        RECT 28.528 26.696 31.28 26.728 ;
  LAYER M1 ;
        RECT 31.264 26.676 31.296 26.748 ;
  LAYER M2 ;
        RECT 31.244 26.696 31.316 26.728 ;
  LAYER M2 ;
        RECT 31.28 26.696 31.344 26.728 ;
  LAYER M1 ;
        RECT 31.328 26.676 31.36 26.748 ;
  LAYER M2 ;
        RECT 31.308 26.696 31.38 26.728 ;
  LAYER M1 ;
        RECT 28.512 23.568 28.544 23.64 ;
  LAYER M2 ;
        RECT 28.492 23.588 28.564 23.62 ;
  LAYER M1 ;
        RECT 28.528 23.588 31.28 23.62 ;
  LAYER M1 ;
        RECT 31.264 23.568 31.296 23.64 ;
  LAYER M2 ;
        RECT 31.244 23.588 31.316 23.62 ;
  LAYER M2 ;
        RECT 31.28 23.588 31.344 23.62 ;
  LAYER M1 ;
        RECT 31.328 23.568 31.36 23.64 ;
  LAYER M2 ;
        RECT 31.308 23.588 31.38 23.62 ;
  LAYER M1 ;
        RECT 28.512 20.46 28.544 20.532 ;
  LAYER M2 ;
        RECT 28.492 20.48 28.564 20.512 ;
  LAYER M1 ;
        RECT 28.528 20.48 31.28 20.512 ;
  LAYER M1 ;
        RECT 31.264 20.46 31.296 20.532 ;
  LAYER M2 ;
        RECT 31.244 20.48 31.316 20.512 ;
  LAYER M2 ;
        RECT 31.28 20.48 31.344 20.512 ;
  LAYER M1 ;
        RECT 31.328 20.46 31.36 20.532 ;
  LAYER M2 ;
        RECT 31.308 20.48 31.38 20.512 ;
  LAYER M1 ;
        RECT 31.328 19.536 31.36 19.608 ;
  LAYER M2 ;
        RECT 31.308 19.556 31.38 19.588 ;
  LAYER M1 ;
        RECT 31.328 19.572 31.36 20.16 ;
  LAYER M1 ;
        RECT 31.328 20.16 31.36 35.868 ;
  LAYER M2 ;
        RECT 16.4 19.556 31.344 19.588 ;
  LAYER M1 ;
        RECT 19.584 36 19.616 36.072 ;
  LAYER M2 ;
        RECT 19.564 36.02 19.636 36.052 ;
  LAYER M2 ;
        RECT 16.624 36.02 19.6 36.052 ;
  LAYER M1 ;
        RECT 16.608 36 16.64 36.072 ;
  LAYER M2 ;
        RECT 16.588 36.02 16.66 36.052 ;
  LAYER M1 ;
        RECT 19.584 20.46 19.616 20.532 ;
  LAYER M2 ;
        RECT 19.564 20.48 19.636 20.512 ;
  LAYER M2 ;
        RECT 16.624 20.48 19.6 20.512 ;
  LAYER M1 ;
        RECT 16.608 20.46 16.64 20.532 ;
  LAYER M2 ;
        RECT 16.588 20.48 16.66 20.512 ;
  LAYER M1 ;
        RECT 22.56 20.46 22.592 20.532 ;
  LAYER M2 ;
        RECT 22.54 20.48 22.612 20.512 ;
  LAYER M2 ;
        RECT 19.6 20.48 22.576 20.512 ;
  LAYER M1 ;
        RECT 19.584 20.46 19.616 20.532 ;
  LAYER M2 ;
        RECT 19.564 20.48 19.636 20.512 ;
  LAYER M1 ;
        RECT 25.536 20.46 25.568 20.532 ;
  LAYER M2 ;
        RECT 25.516 20.48 25.588 20.512 ;
  LAYER M2 ;
        RECT 22.576 20.48 25.552 20.512 ;
  LAYER M1 ;
        RECT 22.56 20.46 22.592 20.532 ;
  LAYER M2 ;
        RECT 22.54 20.48 22.612 20.512 ;
  LAYER M1 ;
        RECT 25.536 36 25.568 36.072 ;
  LAYER M2 ;
        RECT 25.516 36.02 25.588 36.052 ;
  LAYER M2 ;
        RECT 25.552 36.02 28.528 36.052 ;
  LAYER M1 ;
        RECT 28.512 36 28.544 36.072 ;
  LAYER M2 ;
        RECT 28.492 36.02 28.564 36.052 ;
  LAYER M1 ;
        RECT 22.56 36 22.592 36.072 ;
  LAYER M2 ;
        RECT 22.54 36.02 22.612 36.052 ;
  LAYER M2 ;
        RECT 22.576 36.02 25.552 36.052 ;
  LAYER M1 ;
        RECT 25.536 36 25.568 36.072 ;
  LAYER M2 ;
        RECT 25.516 36.02 25.588 36.052 ;
  LAYER M1 ;
        RECT 16.56 35.952 19.056 38.556 ;
  LAYER M3 ;
        RECT 16.56 35.952 19.056 38.556 ;
  LAYER M2 ;
        RECT 16.56 35.952 19.056 38.556 ;
  LAYER M1 ;
        RECT 16.56 32.844 19.056 35.448 ;
  LAYER M3 ;
        RECT 16.56 32.844 19.056 35.448 ;
  LAYER M2 ;
        RECT 16.56 32.844 19.056 35.448 ;
  LAYER M1 ;
        RECT 16.56 29.736 19.056 32.34 ;
  LAYER M3 ;
        RECT 16.56 29.736 19.056 32.34 ;
  LAYER M2 ;
        RECT 16.56 29.736 19.056 32.34 ;
  LAYER M1 ;
        RECT 16.56 26.628 19.056 29.232 ;
  LAYER M3 ;
        RECT 16.56 26.628 19.056 29.232 ;
  LAYER M2 ;
        RECT 16.56 26.628 19.056 29.232 ;
  LAYER M1 ;
        RECT 16.56 23.52 19.056 26.124 ;
  LAYER M3 ;
        RECT 16.56 23.52 19.056 26.124 ;
  LAYER M2 ;
        RECT 16.56 23.52 19.056 26.124 ;
  LAYER M1 ;
        RECT 16.56 20.412 19.056 23.016 ;
  LAYER M3 ;
        RECT 16.56 20.412 19.056 23.016 ;
  LAYER M2 ;
        RECT 16.56 20.412 19.056 23.016 ;
  LAYER M1 ;
        RECT 19.536 35.952 22.032 38.556 ;
  LAYER M3 ;
        RECT 19.536 35.952 22.032 38.556 ;
  LAYER M2 ;
        RECT 19.536 35.952 22.032 38.556 ;
  LAYER M1 ;
        RECT 19.536 32.844 22.032 35.448 ;
  LAYER M3 ;
        RECT 19.536 32.844 22.032 35.448 ;
  LAYER M2 ;
        RECT 19.536 32.844 22.032 35.448 ;
  LAYER M1 ;
        RECT 19.536 29.736 22.032 32.34 ;
  LAYER M3 ;
        RECT 19.536 29.736 22.032 32.34 ;
  LAYER M2 ;
        RECT 19.536 29.736 22.032 32.34 ;
  LAYER M1 ;
        RECT 19.536 26.628 22.032 29.232 ;
  LAYER M3 ;
        RECT 19.536 26.628 22.032 29.232 ;
  LAYER M2 ;
        RECT 19.536 26.628 22.032 29.232 ;
  LAYER M1 ;
        RECT 19.536 23.52 22.032 26.124 ;
  LAYER M3 ;
        RECT 19.536 23.52 22.032 26.124 ;
  LAYER M2 ;
        RECT 19.536 23.52 22.032 26.124 ;
  LAYER M1 ;
        RECT 19.536 20.412 22.032 23.016 ;
  LAYER M3 ;
        RECT 19.536 20.412 22.032 23.016 ;
  LAYER M2 ;
        RECT 19.536 20.412 22.032 23.016 ;
  LAYER M1 ;
        RECT 22.512 35.952 25.008 38.556 ;
  LAYER M3 ;
        RECT 22.512 35.952 25.008 38.556 ;
  LAYER M2 ;
        RECT 22.512 35.952 25.008 38.556 ;
  LAYER M1 ;
        RECT 22.512 32.844 25.008 35.448 ;
  LAYER M3 ;
        RECT 22.512 32.844 25.008 35.448 ;
  LAYER M2 ;
        RECT 22.512 32.844 25.008 35.448 ;
  LAYER M1 ;
        RECT 22.512 29.736 25.008 32.34 ;
  LAYER M3 ;
        RECT 22.512 29.736 25.008 32.34 ;
  LAYER M2 ;
        RECT 22.512 29.736 25.008 32.34 ;
  LAYER M1 ;
        RECT 22.512 26.628 25.008 29.232 ;
  LAYER M3 ;
        RECT 22.512 26.628 25.008 29.232 ;
  LAYER M2 ;
        RECT 22.512 26.628 25.008 29.232 ;
  LAYER M1 ;
        RECT 22.512 23.52 25.008 26.124 ;
  LAYER M3 ;
        RECT 22.512 23.52 25.008 26.124 ;
  LAYER M2 ;
        RECT 22.512 23.52 25.008 26.124 ;
  LAYER M1 ;
        RECT 22.512 20.412 25.008 23.016 ;
  LAYER M3 ;
        RECT 22.512 20.412 25.008 23.016 ;
  LAYER M2 ;
        RECT 22.512 20.412 25.008 23.016 ;
  LAYER M1 ;
        RECT 25.488 35.952 27.984 38.556 ;
  LAYER M3 ;
        RECT 25.488 35.952 27.984 38.556 ;
  LAYER M2 ;
        RECT 25.488 35.952 27.984 38.556 ;
  LAYER M1 ;
        RECT 25.488 32.844 27.984 35.448 ;
  LAYER M3 ;
        RECT 25.488 32.844 27.984 35.448 ;
  LAYER M2 ;
        RECT 25.488 32.844 27.984 35.448 ;
  LAYER M1 ;
        RECT 25.488 29.736 27.984 32.34 ;
  LAYER M3 ;
        RECT 25.488 29.736 27.984 32.34 ;
  LAYER M2 ;
        RECT 25.488 29.736 27.984 32.34 ;
  LAYER M1 ;
        RECT 25.488 26.628 27.984 29.232 ;
  LAYER M3 ;
        RECT 25.488 26.628 27.984 29.232 ;
  LAYER M2 ;
        RECT 25.488 26.628 27.984 29.232 ;
  LAYER M1 ;
        RECT 25.488 23.52 27.984 26.124 ;
  LAYER M3 ;
        RECT 25.488 23.52 27.984 26.124 ;
  LAYER M2 ;
        RECT 25.488 23.52 27.984 26.124 ;
  LAYER M1 ;
        RECT 25.488 20.412 27.984 23.016 ;
  LAYER M3 ;
        RECT 25.488 20.412 27.984 23.016 ;
  LAYER M2 ;
        RECT 25.488 20.412 27.984 23.016 ;
  LAYER M1 ;
        RECT 28.464 35.952 30.96 38.556 ;
  LAYER M3 ;
        RECT 28.464 35.952 30.96 38.556 ;
  LAYER M2 ;
        RECT 28.464 35.952 30.96 38.556 ;
  LAYER M1 ;
        RECT 28.464 32.844 30.96 35.448 ;
  LAYER M3 ;
        RECT 28.464 32.844 30.96 35.448 ;
  LAYER M2 ;
        RECT 28.464 32.844 30.96 35.448 ;
  LAYER M1 ;
        RECT 28.464 29.736 30.96 32.34 ;
  LAYER M3 ;
        RECT 28.464 29.736 30.96 32.34 ;
  LAYER M2 ;
        RECT 28.464 29.736 30.96 32.34 ;
  LAYER M1 ;
        RECT 28.464 26.628 30.96 29.232 ;
  LAYER M3 ;
        RECT 28.464 26.628 30.96 29.232 ;
  LAYER M2 ;
        RECT 28.464 26.628 30.96 29.232 ;
  LAYER M1 ;
        RECT 28.464 23.52 30.96 26.124 ;
  LAYER M3 ;
        RECT 28.464 23.52 30.96 26.124 ;
  LAYER M2 ;
        RECT 28.464 23.52 30.96 26.124 ;
  LAYER M1 ;
        RECT 28.464 20.412 30.96 23.016 ;
  LAYER M3 ;
        RECT 28.464 20.412 30.96 23.016 ;
  LAYER M2 ;
        RECT 28.464 20.412 30.96 23.016 ;
  END 
END switched_capacitor_filter
