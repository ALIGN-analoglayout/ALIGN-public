MACRO CMC_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 1.5560 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 2.2760 0.4360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.3200 1.0560 0.3520 ;
    LAYER V1 ;
      RECT 1.5040 0.3200 1.5360 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
  END
END CMC_NMOS_n12_X2_Y1
MACRO CMC_PMOS_S_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X1_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 0.4360 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 1.0760 0.2680 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 0.9960 0.3520 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.3200 0.9760 0.3520 ;
  END
END CMC_PMOS_S_n12_X1_Y1
MACRO CMC_PMOS_n12_X5_Y2
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X5_Y2 0 0 ;
  SIZE 6.4000 BY 1.6800 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 5.3960 0.1000 ;
      LAYER M2 ;
        RECT 0.8440 0.9080 6.0360 0.9400 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 6.0360 0.2680 ;
      LAYER M2 ;
        RECT 0.2040 1.0760 5.3960 1.1080 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 5.5560 0.1840 ;
      LAYER M2 ;
        RECT 1.0040 0.9920 6.1960 1.0240 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 6.1960 0.3520 ;
      LAYER M2 ;
        RECT 0.3640 1.1600 5.5560 1.1920 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 6.1160 0.4360 ;
      LAYER M2 ;
        RECT 0.2840 1.2440 6.1160 1.2760 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 4.1440 0.0480 4.1760 0.7080 ;
    LAYER M1 ;
      RECT 5.4240 0.0480 5.4560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 4.7840 0.0480 4.8160 0.7080 ;
    LAYER M1 ;
      RECT 6.0640 0.0480 6.0960 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 4.0640 0.0480 4.0960 0.7080 ;
    LAYER V0 ;
      RECT 4.0640 0.2360 4.0960 0.2680 ;
    LAYER V0 ;
      RECT 4.0640 0.3620 4.0960 0.3940 ;
    LAYER V0 ;
      RECT 4.0640 0.4880 4.0960 0.5200 ;
    LAYER M1 ;
      RECT 5.3440 0.0480 5.3760 0.7080 ;
    LAYER V0 ;
      RECT 5.3440 0.2360 5.3760 0.2680 ;
    LAYER V0 ;
      RECT 5.3440 0.3620 5.3760 0.3940 ;
    LAYER V0 ;
      RECT 5.3440 0.4880 5.3760 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER V0 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V0 ;
      RECT 3.4240 0.3620 3.4560 0.3940 ;
    LAYER V0 ;
      RECT 3.4240 0.4880 3.4560 0.5200 ;
    LAYER M1 ;
      RECT 4.7040 0.0480 4.7360 0.7080 ;
    LAYER V0 ;
      RECT 4.7040 0.2360 4.7360 0.2680 ;
    LAYER V0 ;
      RECT 4.7040 0.3620 4.7360 0.3940 ;
    LAYER V0 ;
      RECT 4.7040 0.4880 4.7360 0.5200 ;
    LAYER M1 ;
      RECT 5.9840 0.0480 6.0160 0.7080 ;
    LAYER V0 ;
      RECT 5.9840 0.2360 6.0160 0.2680 ;
    LAYER V0 ;
      RECT 5.9840 0.3620 6.0160 0.3940 ;
    LAYER V0 ;
      RECT 5.9840 0.4880 6.0160 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER M1 ;
      RECT 4.2240 0.0480 4.2560 0.7080 ;
    LAYER V0 ;
      RECT 4.2240 0.2360 4.2560 0.2680 ;
    LAYER V0 ;
      RECT 4.2240 0.3620 4.2560 0.3940 ;
    LAYER V0 ;
      RECT 4.2240 0.4880 4.2560 0.5200 ;
    LAYER M1 ;
      RECT 5.5040 0.0480 5.5360 0.7080 ;
    LAYER V0 ;
      RECT 5.5040 0.2360 5.5360 0.2680 ;
    LAYER V0 ;
      RECT 5.5040 0.3620 5.5360 0.3940 ;
    LAYER V0 ;
      RECT 5.5040 0.4880 5.5360 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER V0 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V0 ;
      RECT 3.5840 0.3620 3.6160 0.3940 ;
    LAYER V0 ;
      RECT 3.5840 0.4880 3.6160 0.5200 ;
    LAYER M1 ;
      RECT 4.8640 0.0480 4.8960 0.7080 ;
    LAYER V0 ;
      RECT 4.8640 0.2360 4.8960 0.2680 ;
    LAYER V0 ;
      RECT 4.8640 0.3620 4.8960 0.3940 ;
    LAYER V0 ;
      RECT 4.8640 0.4880 4.8960 0.5200 ;
    LAYER M1 ;
      RECT 6.1440 0.0480 6.1760 0.7080 ;
    LAYER V0 ;
      RECT 6.1440 0.2360 6.1760 0.2680 ;
    LAYER V0 ;
      RECT 6.1440 0.3620 6.1760 0.3940 ;
    LAYER V0 ;
      RECT 6.1440 0.4880 6.1760 0.5200 ;
    LAYER M3 ;
      RECT 3.0200 0.0480 3.0600 0.1200 ;
    LAYER V2 ;
      RECT 3.0200 0.0680 3.0600 0.1000 ;
    LAYER V2 ;
      RECT 3.0200 0.0680 3.0600 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 4.0640 0.0680 4.0960 0.1000 ;
    LAYER V1 ;
      RECT 5.3440 0.0680 5.3760 0.1000 ;
    LAYER M3 ;
      RECT 2.9400 0.1320 2.9800 0.2040 ;
    LAYER V2 ;
      RECT 2.9400 0.1520 2.9800 0.1840 ;
    LAYER V2 ;
      RECT 2.9400 0.1520 2.9800 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER V1 ;
      RECT 4.2240 0.1520 4.2560 0.1840 ;
    LAYER V1 ;
      RECT 5.5040 0.1520 5.5360 0.1840 ;
    LAYER M3 ;
      RECT 3.1800 0.2160 3.2200 0.2880 ;
    LAYER V2 ;
      RECT 3.1800 0.2360 3.2200 0.2680 ;
    LAYER V2 ;
      RECT 3.1800 0.2360 3.2200 0.2680 ;
    LAYER V1 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V1 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V1 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V1 ;
      RECT 4.7040 0.2360 4.7360 0.2680 ;
    LAYER V1 ;
      RECT 5.9840 0.2360 6.0160 0.2680 ;
    LAYER M3 ;
      RECT 3.2600 0.3000 3.3000 0.3720 ;
    LAYER V2 ;
      RECT 3.2600 0.3200 3.3000 0.3520 ;
    LAYER V2 ;
      RECT 3.2600 0.3200 3.3000 0.3520 ;
    LAYER V1 ;
      RECT 1.0240 0.3200 1.0560 0.3520 ;
    LAYER V1 ;
      RECT 2.3040 0.3200 2.3360 0.3520 ;
    LAYER V1 ;
      RECT 3.5840 0.3200 3.6160 0.3520 ;
    LAYER V1 ;
      RECT 4.8640 0.3200 4.8960 0.3520 ;
    LAYER V1 ;
      RECT 6.1440 0.3200 6.1760 0.3520 ;
    LAYER M3 ;
      RECT 3.1000 0.3840 3.1400 0.4560 ;
    LAYER V2 ;
      RECT 3.1000 0.4040 3.1400 0.4360 ;
    LAYER V2 ;
      RECT 3.1000 0.4040 3.1400 0.4360 ;
    LAYER V1 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER V1 ;
      RECT 2.8640 0.4040 2.8960 0.4360 ;
    LAYER V1 ;
      RECT 4.1440 0.4040 4.1760 0.4360 ;
    LAYER V1 ;
      RECT 5.4240 0.4040 5.4560 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 3.5040 0.4040 3.5360 0.4360 ;
    LAYER V1 ;
      RECT 4.7840 0.4040 4.8160 0.4360 ;
    LAYER V1 ;
      RECT 6.0640 0.4040 6.0960 0.4360 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 4.1440 0.8880 4.1760 1.5480 ;
    LAYER M1 ;
      RECT 5.4240 0.8880 5.4560 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 3.5040 0.8880 3.5360 1.5480 ;
    LAYER M1 ;
      RECT 4.7840 0.8880 4.8160 1.5480 ;
    LAYER M1 ;
      RECT 6.0640 0.8880 6.0960 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER V0 ;
      RECT 2.7840 1.0760 2.8160 1.1080 ;
    LAYER V0 ;
      RECT 2.7840 1.2020 2.8160 1.2340 ;
    LAYER V0 ;
      RECT 2.7840 1.3280 2.8160 1.3600 ;
    LAYER M1 ;
      RECT 4.0640 0.8880 4.0960 1.5480 ;
    LAYER V0 ;
      RECT 4.0640 1.0760 4.0960 1.1080 ;
    LAYER V0 ;
      RECT 4.0640 1.2020 4.0960 1.2340 ;
    LAYER V0 ;
      RECT 4.0640 1.3280 4.0960 1.3600 ;
    LAYER M1 ;
      RECT 5.3440 0.8880 5.3760 1.5480 ;
    LAYER V0 ;
      RECT 5.3440 1.0760 5.3760 1.1080 ;
    LAYER V0 ;
      RECT 5.3440 1.2020 5.3760 1.2340 ;
    LAYER V0 ;
      RECT 5.3440 1.3280 5.3760 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER V0 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER V0 ;
      RECT 2.1440 1.2020 2.1760 1.2340 ;
    LAYER V0 ;
      RECT 2.1440 1.3280 2.1760 1.3600 ;
    LAYER M1 ;
      RECT 3.4240 0.8880 3.4560 1.5480 ;
    LAYER V0 ;
      RECT 3.4240 1.0760 3.4560 1.1080 ;
    LAYER V0 ;
      RECT 3.4240 1.2020 3.4560 1.2340 ;
    LAYER V0 ;
      RECT 3.4240 1.3280 3.4560 1.3600 ;
    LAYER M1 ;
      RECT 4.7040 0.8880 4.7360 1.5480 ;
    LAYER V0 ;
      RECT 4.7040 1.0760 4.7360 1.1080 ;
    LAYER V0 ;
      RECT 4.7040 1.2020 4.7360 1.2340 ;
    LAYER V0 ;
      RECT 4.7040 1.3280 4.7360 1.3600 ;
    LAYER M1 ;
      RECT 5.9840 0.8880 6.0160 1.5480 ;
    LAYER V0 ;
      RECT 5.9840 1.0760 6.0160 1.1080 ;
    LAYER V0 ;
      RECT 5.9840 1.2020 6.0160 1.2340 ;
    LAYER V0 ;
      RECT 5.9840 1.3280 6.0160 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER V0 ;
      RECT 2.9440 1.0760 2.9760 1.1080 ;
    LAYER V0 ;
      RECT 2.9440 1.2020 2.9760 1.2340 ;
    LAYER V0 ;
      RECT 2.9440 1.3280 2.9760 1.3600 ;
    LAYER M1 ;
      RECT 4.2240 0.8880 4.2560 1.5480 ;
    LAYER V0 ;
      RECT 4.2240 1.0760 4.2560 1.1080 ;
    LAYER V0 ;
      RECT 4.2240 1.2020 4.2560 1.2340 ;
    LAYER V0 ;
      RECT 4.2240 1.3280 4.2560 1.3600 ;
    LAYER M1 ;
      RECT 5.5040 0.8880 5.5360 1.5480 ;
    LAYER V0 ;
      RECT 5.5040 1.0760 5.5360 1.1080 ;
    LAYER V0 ;
      RECT 5.5040 1.2020 5.5360 1.2340 ;
    LAYER V0 ;
      RECT 5.5040 1.3280 5.5360 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER V0 ;
      RECT 2.3040 1.0760 2.3360 1.1080 ;
    LAYER V0 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER V0 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER M1 ;
      RECT 3.5840 0.8880 3.6160 1.5480 ;
    LAYER V0 ;
      RECT 3.5840 1.0760 3.6160 1.1080 ;
    LAYER V0 ;
      RECT 3.5840 1.2020 3.6160 1.2340 ;
    LAYER V0 ;
      RECT 3.5840 1.3280 3.6160 1.3600 ;
    LAYER M1 ;
      RECT 4.8640 0.8880 4.8960 1.5480 ;
    LAYER V0 ;
      RECT 4.8640 1.0760 4.8960 1.1080 ;
    LAYER V0 ;
      RECT 4.8640 1.2020 4.8960 1.2340 ;
    LAYER V0 ;
      RECT 4.8640 1.3280 4.8960 1.3600 ;
    LAYER M1 ;
      RECT 6.1440 0.8880 6.1760 1.5480 ;
    LAYER V0 ;
      RECT 6.1440 1.0760 6.1760 1.1080 ;
    LAYER V0 ;
      RECT 6.1440 1.2020 6.1760 1.2340 ;
    LAYER V0 ;
      RECT 6.1440 1.3280 6.1760 1.3600 ;
    LAYER M3 ;
      RECT 3.0200 0.0480 3.0600 0.9600 ;
    LAYER V2 ;
      RECT 3.0200 0.0680 3.0600 0.1000 ;
    LAYER V2 ;
      RECT 3.0200 0.9080 3.0600 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 2.1440 0.9080 2.1760 0.9400 ;
    LAYER V1 ;
      RECT 3.4240 0.9080 3.4560 0.9400 ;
    LAYER V1 ;
      RECT 4.7040 0.9080 4.7360 0.9400 ;
    LAYER V1 ;
      RECT 5.9840 0.9080 6.0160 0.9400 ;
    LAYER M3 ;
      RECT 2.9400 0.1320 2.9800 1.0440 ;
    LAYER V2 ;
      RECT 2.9400 0.1520 2.9800 0.1840 ;
    LAYER V2 ;
      RECT 2.9400 0.9920 2.9800 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 2.3040 0.9920 2.3360 1.0240 ;
    LAYER V1 ;
      RECT 3.5840 0.9920 3.6160 1.0240 ;
    LAYER V1 ;
      RECT 4.8640 0.9920 4.8960 1.0240 ;
    LAYER V1 ;
      RECT 6.1440 0.9920 6.1760 1.0240 ;
    LAYER M3 ;
      RECT 3.1800 0.2160 3.2200 1.1280 ;
    LAYER V2 ;
      RECT 3.1800 0.2360 3.2200 0.2680 ;
    LAYER V2 ;
      RECT 3.1800 1.0760 3.2200 1.1080 ;
    LAYER V1 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V1 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V1 ;
      RECT 2.7840 1.0760 2.8160 1.1080 ;
    LAYER V1 ;
      RECT 4.0640 1.0760 4.0960 1.1080 ;
    LAYER V1 ;
      RECT 5.3440 1.0760 5.3760 1.1080 ;
    LAYER M3 ;
      RECT 3.2600 0.3000 3.3000 1.2120 ;
    LAYER V2 ;
      RECT 3.2600 0.3200 3.3000 0.3520 ;
    LAYER V2 ;
      RECT 3.2600 1.1600 3.3000 1.1920 ;
    LAYER V1 ;
      RECT 0.3840 1.1600 0.4160 1.1920 ;
    LAYER V1 ;
      RECT 1.6640 1.1600 1.6960 1.1920 ;
    LAYER V1 ;
      RECT 2.9440 1.1600 2.9760 1.1920 ;
    LAYER V1 ;
      RECT 4.2240 1.1600 4.2560 1.1920 ;
    LAYER V1 ;
      RECT 5.5040 1.1600 5.5360 1.1920 ;
    LAYER M3 ;
      RECT 3.1000 0.3840 3.1400 1.2960 ;
    LAYER V2 ;
      RECT 3.1000 0.4040 3.1400 0.4360 ;
    LAYER V2 ;
      RECT 3.1000 1.2440 3.1400 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V1 ;
      RECT 1.5840 1.2440 1.6160 1.2760 ;
    LAYER V1 ;
      RECT 2.8640 1.2440 2.8960 1.2760 ;
    LAYER V1 ;
      RECT 4.1440 1.2440 4.1760 1.2760 ;
    LAYER V1 ;
      RECT 5.4240 1.2440 5.4560 1.2760 ;
    LAYER V1 ;
      RECT 0.9440 1.2440 0.9760 1.2760 ;
    LAYER V1 ;
      RECT 2.2240 1.2440 2.2560 1.2760 ;
    LAYER V1 ;
      RECT 3.5040 1.2440 3.5360 1.2760 ;
    LAYER V1 ;
      RECT 4.7840 1.2440 4.8160 1.2760 ;
    LAYER V1 ;
      RECT 6.0640 1.2440 6.0960 1.2760 ;
  END
END CMC_PMOS_n12_X5_Y2
MACRO DCL_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.2760 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.4360 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
  END
END DCL_NMOS_n12_X1_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 1.0760 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DCL_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.2760 0.1000 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.4360 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
  END
END DCL_PMOS_n12_X1_Y1
MACRO DP_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 3.4760 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 3.6360 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 2.9160 0.3520 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4040 3.5560 0.4360 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER V0 ;
      RECT 3.4240 0.2360 3.4560 0.2680 ;
    LAYER V0 ;
      RECT 3.4240 0.3620 3.4560 0.3940 ;
    LAYER V0 ;
      RECT 3.4240 0.4880 3.4560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER V0 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V0 ;
      RECT 3.5840 0.3620 3.6160 0.3940 ;
    LAYER V0 ;
      RECT 3.5840 0.4880 3.6160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 3.4240 0.0680 3.4560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V1 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 1.5840 0.3200 1.6160 0.3520 ;
    LAYER V1 ;
      RECT 2.8640 0.3200 2.8960 0.3520 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 2.2240 0.4040 2.2560 0.4360 ;
    LAYER V1 ;
      RECT 3.5040 0.4040 3.5360 0.4360 ;
  END
END DP_NMOS_n12_X3_Y1
MACRO SCM_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 2.2760 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 1.5560 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 2.2240 0.1520 2.2560 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 1.5840 0.1520 1.6160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
  END
END SCM_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.9160 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.9960 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.0760 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
  END
END Switch_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y1 0 0 ;
  SIZE 1.9200 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.5560 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 1.6360 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 1.7160 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
  END
END Switch_NMOS_n12_X3_Y1
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 0.2760 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.3560 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 0.4360 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X5_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X5_Y1 0 0 ;
  SIZE 3.2000 BY 0.8400 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.8360 0.1000 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 2.9160 0.2680 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.3040 0.1520 2.3360 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
    LAYER V1 ;
      RECT 2.2240 0.2360 2.2560 0.2680 ;
    LAYER V1 ;
      RECT 2.8640 0.2360 2.8960 0.2680 ;
  END
END Switch_PMOS_n12_X5_Y1
MACRO Switch_PMOS_n12_X5_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X5_Y2 0 0 ;
  SIZE 3.2000 BY 1.6800 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.8360 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 2.8360 0.9400 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 2.9160 0.2680 ;
      LAYER M2 ;
        RECT 0.2840 1.0760 2.9160 1.1080 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
      LAYER M2 ;
        RECT 0.3640 0.9920 2.9960 1.0240 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER V0 ;
      RECT 2.7840 0.2360 2.8160 0.2680 ;
    LAYER V0 ;
      RECT 2.7840 0.3620 2.8160 0.3940 ;
    LAYER V0 ;
      RECT 2.7840 0.4880 2.8160 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER V0 ;
      RECT 2.9440 0.2360 2.9760 0.2680 ;
    LAYER V0 ;
      RECT 2.9440 0.3620 2.9760 0.3940 ;
    LAYER V0 ;
      RECT 2.9440 0.4880 2.9760 0.5200 ;
    LAYER M3 ;
      RECT 1.5000 0.0480 1.5400 0.1200 ;
    LAYER V2 ;
      RECT 1.5000 0.0680 1.5400 0.1000 ;
    LAYER V2 ;
      RECT 1.5000 0.0680 1.5400 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER M3 ;
      RECT 1.5800 0.1320 1.6200 0.2040 ;
    LAYER V2 ;
      RECT 1.5800 0.1520 1.6200 0.1840 ;
    LAYER V2 ;
      RECT 1.5800 0.1520 1.6200 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 2.3040 0.1520 2.3360 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER M3 ;
      RECT 1.4200 0.2160 1.4600 0.2880 ;
    LAYER V2 ;
      RECT 1.4200 0.2360 1.4600 0.2680 ;
    LAYER V2 ;
      RECT 1.4200 0.2360 1.4600 0.2680 ;
    LAYER V1 ;
      RECT 0.3040 0.2360 0.3360 0.2680 ;
    LAYER V1 ;
      RECT 0.9440 0.2360 0.9760 0.2680 ;
    LAYER V1 ;
      RECT 1.5840 0.2360 1.6160 0.2680 ;
    LAYER V1 ;
      RECT 2.2240 0.2360 2.2560 0.2680 ;
    LAYER V1 ;
      RECT 2.8640 0.2360 2.8960 0.2680 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER V0 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER V0 ;
      RECT 2.1440 1.2020 2.1760 1.2340 ;
    LAYER V0 ;
      RECT 2.1440 1.3280 2.1760 1.3600 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER V0 ;
      RECT 2.7840 1.0760 2.8160 1.1080 ;
    LAYER V0 ;
      RECT 2.7840 1.2020 2.8160 1.2340 ;
    LAYER V0 ;
      RECT 2.7840 1.3280 2.8160 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER V0 ;
      RECT 2.3040 1.0760 2.3360 1.1080 ;
    LAYER V0 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER V0 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER V0 ;
      RECT 2.9440 1.0760 2.9760 1.1080 ;
    LAYER V0 ;
      RECT 2.9440 1.2020 2.9760 1.2340 ;
    LAYER V0 ;
      RECT 2.9440 1.3280 2.9760 1.3600 ;
    LAYER M3 ;
      RECT 1.5000 0.0480 1.5400 0.9600 ;
    LAYER V2 ;
      RECT 1.5000 0.0680 1.5400 0.1000 ;
    LAYER V2 ;
      RECT 1.5000 0.9080 1.5400 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 1.5040 0.9080 1.5360 0.9400 ;
    LAYER V1 ;
      RECT 2.1440 0.9080 2.1760 0.9400 ;
    LAYER V1 ;
      RECT 2.7840 0.9080 2.8160 0.9400 ;
    LAYER M3 ;
      RECT 1.5800 0.1320 1.6200 1.0440 ;
    LAYER V2 ;
      RECT 1.5800 0.1520 1.6200 0.1840 ;
    LAYER V2 ;
      RECT 1.5800 0.9920 1.6200 1.0240 ;
    LAYER V1 ;
      RECT 0.3840 0.9920 0.4160 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.6640 0.9920 1.6960 1.0240 ;
    LAYER V1 ;
      RECT 2.3040 0.9920 2.3360 1.0240 ;
    LAYER V1 ;
      RECT 2.9440 0.9920 2.9760 1.0240 ;
    LAYER M3 ;
      RECT 1.4200 0.2160 1.4600 1.1280 ;
    LAYER V2 ;
      RECT 1.4200 0.2360 1.4600 0.2680 ;
    LAYER V2 ;
      RECT 1.4200 1.0760 1.4600 1.1080 ;
    LAYER V1 ;
      RECT 0.3040 1.0760 0.3360 1.1080 ;
    LAYER V1 ;
      RECT 0.9440 1.0760 0.9760 1.1080 ;
    LAYER V1 ;
      RECT 1.5840 1.0760 1.6160 1.1080 ;
    LAYER V1 ;
      RECT 2.2240 1.0760 2.2560 1.1080 ;
    LAYER V1 ;
      RECT 2.8640 1.0760 2.8960 1.1080 ;
  END
END Switch_PMOS_n12_X5_Y2
