.subckt TEST gnd ibias vdd vref vrefp
xm72 net0211 net0211 net0211 gnd nfet w=w0 l=l0
xm71 gnd gnd gnd gnd nfet w=w1 l=l0
xm70 net0176 net0176 net0176 gnd nfet w=w2 l=l1
xm69 net0211 net0211 net0211 gnd nfet w=w3 l=l1
xm54 net0144 net0144 net0144 gnd nfet w=w4 l=l1
xm51 net0111 net0111 net0111 gnd nfet w=w4 l=l1
xm50 net0111 net0111 net0111 gnd nfet w=w4 l=l1
xm48 net0129 net0129 net0129 gnd nfet w=w4 l=l1
xm43 net0109 net0109 net0109 gnd nfet w=w4 l=l1
xm68 net0160 net0160 net0160 gnd nfet w=w3 l=l1
xm62 net0147 net0147 net0147 gnd nfet w=w3 l=l2
xm65 net0149 net0149 net0149 gnd nfet w=w0 l=l0
xm58 net0103 net0103 net0103 gnd nfet w=w3 l=l2
xm55 net0103 net0103 net0103 gnd nfet w=w4 l=l1
xm57 net0111 net0111 net0111 gnd nfet w=w2 l=l1
xm59 net0144 net0144 net0144 gnd nfet w=w3 l=l2
xm61 net0149 net0149 net0149 gnd nfet w=w3 l=l2
xm25 net0147 vdd gnd gnd nfet w=w5 l=l0
xm24 net0148 vdd gnd gnd nfet w=w0 l=l0
xm23 net0149 vdd gnd gnd nfet w=w5 l=l0
xm22 net0144 net0103 net0147 gnd nfet w=w6 l=l2
xm1 net0103 net0103 net0149 gnd nfet w=w6 l=l2
xm20 net0111 ibias net0148 gnd nfet w=w3 l=l1
xm19 net0129 vfb net0111 gnd nfet w=w7 l=l1
xm18 net0103 vfb net0111 gnd nfet w=w7 l=l1
xm17 net0109 vref net0111 gnd nfet w=w7 l=l1
xm16 net0144 vref net0111 gnd nfet w=w7 l=l1
xm67 net0211 vdd gnd gnd nfet w=w5 l=l0
xm21 net0160 ibias net0211 gnd nfet w=w6 l=l1
xm63 gnd gnd gnd gnd nfet w=w1 l=l0
xm64 net0147 net0147 net0147 gnd nfet w=w0 l=l0
xm30 net0176 ibias net0207 gnd nfet w=w8 l=l1
xm14 net0140 net0140 net0140 gnd nfet w=w3 l=l1
xm8 net0140 ibias net016 gnd nfet w=w6 l=l1
xm7 ibias ibias net017 gnd nfet w=w6 l=l1
xm6 net017 vdd gnd gnd nfet w=w0 l=l0
xm3 net016 vdd gnd gnd nfet w=w5 l=l0
xm9 gnd gnd gnd gnd nfet w=w1 l=l0
xm10 net016 net016 net016 gnd nfet w=w0 l=l0
xm11 ibias ibias ibias gnd nfet w=w3 l=l1
xm66 net0207 vdd gnd gnd nfet w=w9 l=l0
xm13 net016 net016 net016 gnd nfet w=w3 l=l1
xm12 net017 net017 net017 gnd nfet w=w3 l=l1
xm35 vdd net0144 vdd vdd pfet_lvt w=w10 l=l3
xm2 vfb vfb vfb vdd pfet_lvt w=w11 l=l1
xm4 net0168 net0168 net0168 vdd pfet_lvt w=w12 l=l1
xm5 vrefp vrefp vrefp vdd pfet_lvt w=w13 l=l1
xm31 net0160 net0160 net0160 vdd pfet_lvt w=w14 l=l1
xm28 vrefp net0176 net0168 vdd pfet_lvt w=w15 l=l1
xm26 vfb vfb vfb vdd pfet_lvt w=w14 l=l1
xm0 net0156 net0156 net0156 vdd pfet_lvt w=w11 l=l1
xm34 vdd net0160 vdd vdd pfet_lvt w=w16 l=l4
xm29 net0176 net0160 vrefp vdd pfet_lvt w=w17 l=l1
xm15 vfb net0144 net0156 vdd pfet_lvt w=w18 l=l1
xm27 net0160 net0160 vfb vdd pfet_lvt w=w19 l=l1
xm79 net0122 net0122 net0122 vdd pfet w=w20 l=l1
xm75 vdd vdd vdd vdd pfet w=w21 l=l0
xm60 net0134 gnd vdd vdd pfet w=w22 l=l0
xm56 net0118 gnd vdd vdd pfet w=w10 l=l0
xm53 net0122 gnd vdd vdd pfet w=w10 l=l0
xm52 net0101 gnd vdd vdd pfet w=w22 l=l0
xm49 net093 gnd vdd vdd pfet w=w9 l=l0
xm47 net0144 net0140 net0133 vdd pfet w=w23 l=l1
xm46 net0103 net0140 net0102 vdd pfet w=w23 l=l1
xm45 net0140 net0140 net093 vdd pfet w=w24 l=l5
xm44 net0129 net0129 net0122 vdd pfet w=w4 l=l1
xm42 net0133 net0129 net0134 vdd pfet w=w25 l=l1
xm41 net0109 net0109 net0118 vdd pfet w=w4 l=l1
xm40 net0102 net0109 net0101 vdd pfet w=w25 l=l1
xm85 net0133 net0133 net0133 vdd pfet w=w23 l=l1
xm84 net0102 net0102 net0102 vdd pfet w=w23 l=l1
xm83 net0134 net0134 net0134 vdd pfet w=w26 l=l1
xm82 net0101 net0101 net0101 vdd pfet w=w26 l=l1
xm81 net0129 net0129 net0129 vdd pfet w=w20 l=l1
xm80 net0109 net0109 net0109 vdd pfet w=w20 l=l1
xm73 net0140 net0140 net0140 vdd pfet w=w27 l=l5
xm77 net0118 net0118 net0118 vdd pfet w=w9 l=l0
xm78 net0118 net0118 net0118 vdd pfet w=w20 l=l1
xm74 net093 net093 net093 vdd pfet w=w27 l=l5
xm89 net0156 net0156 net0156 vdd pfet w=w9 l=l0
xm88 vdd vdd vdd vdd pfet w=w28 l=l0
xm86 net0168 gnd vdd vdd pfet w=w22 l=l0
xm87 net0156 gnd vdd vdd pfet w=w10 l=l0
xm76 net0122 net0122 net0122 vdd pfet w=w9 l=l0
.ends TEST

