VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO CMC_NMOS_25_1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_25_1 0 0 ;
  SIZE 2.16 BY 0.466 ;
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.192 2.012 0.21 ;
    END
  END D2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.448 2.16 0.466 ;
    END
  END VDD
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.32 2.066 0.338 ;
    END
  END G
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.256 1.904 0.274 ;
    END
  END D1
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.064 2.12 0.082 ;
    END
  END S2
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.128 1.796 0.146 ;
    END
  END S1
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 2.16 0.018 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0 0 2.16 0.466 ;
  END
END CMC_NMOS_25_1

MACRO CMC_PMOS_10_1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_10_1 0 0 ;
  SIZE 0.864 BY 0.402 ;
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 0.608 0.146 ;
    END
  END D1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.864 0.402 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
    END
  END VSS
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 0.77 0.082 ;
    END
  END G
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.32 0.824 0.338 ;
    END
  END S2
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.192 0.716 0.21 ;
    END
  END D2
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 0.5 0.274 ;
    END
  END S1
  OBS
    LAYER M1 ;
      RECT 0 0 0.864 0.402 ;
  END
END CMC_PMOS_10_1


MACRO CMC_PMOS_15_1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_15_1 0 0 ;
  SIZE 1.296 BY 0.402 ;
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.256 0.932 0.274 ;
    END
  END S1
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 1.296 0.018 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 1.296 0.402 ;
    END
  END VDD
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.364 0.32 1.256 0.338 ;
    END
  END S2
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.064 1.202 0.082 ;
    END
  END G
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.192 1.148 0.21 ;
    END
  END D2
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 1.04 0.146 ;
    END
  END D1
  OBS
    LAYER M1 ;
      RECT 0 0 1.296 0.402 ;
  END
END CMC_PMOS_15_1

MACRO Cap_192f
  ORIGIN 0 0 ;
  FOREIGN Cap_192f 0 0 ;
  SIZE 24.184 BY 4.024 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 24.184 0.023 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.001 24.184 4.019 ;
    END
  END PLUS
END Cap_192f


MACRO Cap_32f
  ORIGIN 0 0 ;
  FOREIGN Cap_32f 0 0 ;
  SIZE 4.024 BY 4.024 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 4.024 0.023 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.001 4.024 4.019 ;
    END
  END PLUS
END Cap_32f

MACRO Cap_352f
  ORIGIN 0 0 ;
  FOREIGN Cap_352f 0 0 ;
  SIZE 13.384 BY 13.384 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 13.361 13.384 13.379 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 13.384 0.023 ;
    END
  END MINUS
END Cap_352f


MACRO Cap_96f
  ORIGIN 0 0 ;
  FOREIGN Cap_96f 0 0 ;
  SIZE 12.087 BY 4.024 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 4.001 12.087 4.019 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.005 12.088 0.023 ;
    END
  END MINUS
END Cap_96f

MACRO DP_NMOS_70_1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_70_1 0 0 ;
  SIZE 6.048 BY 0.402 ;
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 6.048 0.018 ;
    END
  END VSS
  PIN G1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.32 5.954 0.338 ;
    END
  END G1
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.256 5.792 0.274 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.256 0.192 5.9 0.21 ;
    END
  END D2
  PIN G2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.31 0.128 5.954 0.146 ;
    END
  END G2
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.064 6.008 0.082 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 6.048 0.402 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0 0 6.048 0.402 ;
  END
END DP_NMOS_70_1

MACRO SCM_NMOS_50
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_50 0 0 ;
  SIZE 2.592 BY 0.402 ;
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.228 0.192 1.364 0.21 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.336 0.192 1.364 0.21 ;
    END
  END D1
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 2.592 0.018 ;
    END
  END VSS
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.064 2.552 0.082 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 2.592 0.402 ;
    END
  END VDD
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.128 2.444 0.146 ;
    END
  END D2
  OBS
    LAYER M1 ;
      RECT 0 0 2.592 0.402 ;
  END
END SCM_NMOS_50

MACRO Switch_NMOS_10
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_10 0 0 ;
  SIZE 0.432 BY 0.466 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.064 0.392 0.082 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.384 0.284 0.402 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.128 0.338 0.146 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.448 0.432 0.466 ;
    END
  END VDD
END Switch_NMOS_10

MACRO Switch_PMOS_10
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_10 0 0 ;
  SIZE 0.432 BY 0.466 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.32 0.392 0.338 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.064 0.284 0.082 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.256 0.338 0.274 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.448 0.432 0.466 ;
    END
  END VDD
END Switch_PMOS_10

END LIBRARY
