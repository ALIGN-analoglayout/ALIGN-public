MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 9.92 BY 24.864 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.584 24.408 3.616 24.48 ;
      LAYER M2 ;
        RECT 3.564 24.428 3.636 24.46 ;
      LAYER M1 ;
        RECT 6.784 24.408 6.816 24.48 ;
      LAYER M2 ;
        RECT 6.764 24.428 6.836 24.46 ;
      LAYER M2 ;
        RECT 3.6 24.428 6.8 24.46 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.264 0.384 3.296 0.456 ;
      LAYER M2 ;
        RECT 3.244 0.404 3.316 0.436 ;
      LAYER M1 ;
        RECT 6.464 0.384 6.496 0.456 ;
      LAYER M2 ;
        RECT 6.444 0.404 6.516 0.436 ;
      LAYER M2 ;
        RECT 3.28 0.404 6.48 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.744 24.576 3.776 24.648 ;
      LAYER M2 ;
        RECT 3.724 24.596 3.796 24.628 ;
      LAYER M1 ;
        RECT 6.944 24.576 6.976 24.648 ;
      LAYER M2 ;
        RECT 6.924 24.596 6.996 24.628 ;
      LAYER M2 ;
        RECT 3.76 24.596 6.96 24.628 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.424 0.216 3.456 0.288 ;
      LAYER M2 ;
        RECT 3.404 0.236 3.476 0.268 ;
      LAYER M1 ;
        RECT 6.624 0.216 6.656 0.288 ;
      LAYER M2 ;
        RECT 6.604 0.236 6.676 0.268 ;
      LAYER M2 ;
        RECT 3.44 0.236 6.64 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 3.904 12.648 3.936 12.72 ;
  LAYER M2 ;
        RECT 3.884 12.668 3.956 12.7 ;
  LAYER M2 ;
        RECT 3.28 12.668 3.92 12.7 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 12.72 ;
  LAYER M2 ;
        RECT 3.244 12.668 3.316 12.7 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 6.84 ;
  LAYER M2 ;
        RECT 3.884 6.788 3.956 6.82 ;
  LAYER M2 ;
        RECT 3.28 6.788 3.92 6.82 ;
  LAYER M1 ;
        RECT 3.264 6.768 3.296 6.84 ;
  LAYER M2 ;
        RECT 3.244 6.788 3.316 6.82 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 15.66 ;
  LAYER M2 ;
        RECT 3.884 15.608 3.956 15.64 ;
  LAYER M2 ;
        RECT 3.28 15.608 3.92 15.64 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M1 ;
        RECT 3.264 0.384 3.296 0.456 ;
  LAYER M2 ;
        RECT 3.244 0.404 3.316 0.436 ;
  LAYER M1 ;
        RECT 3.264 0.42 3.296 0.588 ;
  LAYER M1 ;
        RECT 3.264 0.588 3.296 15.624 ;
  LAYER M1 ;
        RECT 3.904 12.648 3.936 12.72 ;
  LAYER M2 ;
        RECT 3.884 12.668 3.956 12.7 ;
  LAYER M1 ;
        RECT 3.904 12.516 3.936 12.684 ;
  LAYER M1 ;
        RECT 3.904 12.48 3.936 12.552 ;
  LAYER M2 ;
        RECT 3.884 12.5 3.956 12.532 ;
  LAYER M2 ;
        RECT 3.92 12.5 6.48 12.532 ;
  LAYER M1 ;
        RECT 6.464 12.48 6.496 12.552 ;
  LAYER M2 ;
        RECT 6.444 12.5 6.516 12.532 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 6.84 ;
  LAYER M2 ;
        RECT 3.884 6.788 3.956 6.82 ;
  LAYER M1 ;
        RECT 3.904 6.636 3.936 6.804 ;
  LAYER M1 ;
        RECT 3.904 6.6 3.936 6.672 ;
  LAYER M2 ;
        RECT 3.884 6.62 3.956 6.652 ;
  LAYER M2 ;
        RECT 3.92 6.62 6.48 6.652 ;
  LAYER M1 ;
        RECT 6.464 6.6 6.496 6.672 ;
  LAYER M2 ;
        RECT 6.444 6.62 6.516 6.652 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 15.66 ;
  LAYER M2 ;
        RECT 3.884 15.608 3.956 15.64 ;
  LAYER M1 ;
        RECT 3.904 15.456 3.936 15.624 ;
  LAYER M1 ;
        RECT 3.904 15.42 3.936 15.492 ;
  LAYER M2 ;
        RECT 3.884 15.44 3.956 15.472 ;
  LAYER M2 ;
        RECT 3.92 15.44 6.48 15.472 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 15.492 ;
  LAYER M2 ;
        RECT 6.444 15.44 6.516 15.472 ;
  LAYER M1 ;
        RECT 6.464 0.384 6.496 0.456 ;
  LAYER M2 ;
        RECT 6.444 0.404 6.516 0.436 ;
  LAYER M1 ;
        RECT 6.464 0.42 6.496 0.588 ;
  LAYER M1 ;
        RECT 6.464 0.588 6.496 15.456 ;
  LAYER M2 ;
        RECT 3.28 0.404 6.48 0.436 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 9.78 ;
  LAYER M2 ;
        RECT 3.884 9.728 3.956 9.76 ;
  LAYER M2 ;
        RECT 3.44 9.728 3.92 9.76 ;
  LAYER M1 ;
        RECT 3.424 9.708 3.456 9.78 ;
  LAYER M2 ;
        RECT 3.404 9.728 3.476 9.76 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 3.9 ;
  LAYER M2 ;
        RECT 3.884 3.848 3.956 3.88 ;
  LAYER M2 ;
        RECT 3.44 3.848 3.92 3.88 ;
  LAYER M1 ;
        RECT 3.424 3.828 3.456 3.9 ;
  LAYER M2 ;
        RECT 3.404 3.848 3.476 3.88 ;
  LAYER M1 ;
        RECT 3.904 18.528 3.936 18.6 ;
  LAYER M2 ;
        RECT 3.884 18.548 3.956 18.58 ;
  LAYER M2 ;
        RECT 3.44 18.548 3.92 18.58 ;
  LAYER M1 ;
        RECT 3.424 18.528 3.456 18.6 ;
  LAYER M2 ;
        RECT 3.404 18.548 3.476 18.58 ;
  LAYER M1 ;
        RECT 3.424 0.216 3.456 0.288 ;
  LAYER M2 ;
        RECT 3.404 0.236 3.476 0.268 ;
  LAYER M1 ;
        RECT 3.424 0.252 3.456 0.588 ;
  LAYER M1 ;
        RECT 3.424 0.588 3.456 18.564 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 9.78 ;
  LAYER M2 ;
        RECT 3.884 9.728 3.956 9.76 ;
  LAYER M1 ;
        RECT 3.904 9.576 3.936 9.744 ;
  LAYER M1 ;
        RECT 3.904 9.54 3.936 9.612 ;
  LAYER M2 ;
        RECT 3.884 9.56 3.956 9.592 ;
  LAYER M2 ;
        RECT 3.92 9.56 6.64 9.592 ;
  LAYER M1 ;
        RECT 6.624 9.54 6.656 9.612 ;
  LAYER M2 ;
        RECT 6.604 9.56 6.676 9.592 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 3.9 ;
  LAYER M2 ;
        RECT 3.884 3.848 3.956 3.88 ;
  LAYER M1 ;
        RECT 3.904 3.696 3.936 3.864 ;
  LAYER M1 ;
        RECT 3.904 3.66 3.936 3.732 ;
  LAYER M2 ;
        RECT 3.884 3.68 3.956 3.712 ;
  LAYER M2 ;
        RECT 3.92 3.68 6.64 3.712 ;
  LAYER M1 ;
        RECT 6.624 3.66 6.656 3.732 ;
  LAYER M2 ;
        RECT 6.604 3.68 6.676 3.712 ;
  LAYER M1 ;
        RECT 3.904 18.528 3.936 18.6 ;
  LAYER M2 ;
        RECT 3.884 18.548 3.956 18.58 ;
  LAYER M1 ;
        RECT 3.904 18.396 3.936 18.564 ;
  LAYER M1 ;
        RECT 3.904 18.36 3.936 18.432 ;
  LAYER M2 ;
        RECT 3.884 18.38 3.956 18.412 ;
  LAYER M2 ;
        RECT 3.92 18.38 6.64 18.412 ;
  LAYER M1 ;
        RECT 6.624 18.36 6.656 18.432 ;
  LAYER M2 ;
        RECT 6.604 18.38 6.676 18.412 ;
  LAYER M1 ;
        RECT 6.624 0.216 6.656 0.288 ;
  LAYER M2 ;
        RECT 6.604 0.236 6.676 0.268 ;
  LAYER M1 ;
        RECT 6.624 0.252 6.656 0.588 ;
  LAYER M1 ;
        RECT 6.624 0.588 6.656 18.396 ;
  LAYER M2 ;
        RECT 3.44 0.236 6.64 0.268 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 0.96 ;
  LAYER M2 ;
        RECT 0.684 0.908 0.756 0.94 ;
  LAYER M2 ;
        RECT 0.08 0.908 0.72 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 0.704 3.828 0.736 3.9 ;
  LAYER M2 ;
        RECT 0.684 3.848 0.756 3.88 ;
  LAYER M2 ;
        RECT 0.08 3.848 0.72 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 0.704 6.768 0.736 6.84 ;
  LAYER M2 ;
        RECT 0.684 6.788 0.756 6.82 ;
  LAYER M2 ;
        RECT 0.08 6.788 0.72 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.704 9.708 0.736 9.78 ;
  LAYER M2 ;
        RECT 0.684 9.728 0.756 9.76 ;
  LAYER M2 ;
        RECT 0.08 9.728 0.72 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.704 12.648 0.736 12.72 ;
  LAYER M2 ;
        RECT 0.684 12.668 0.756 12.7 ;
  LAYER M2 ;
        RECT 0.08 12.668 0.72 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.704 15.588 0.736 15.66 ;
  LAYER M2 ;
        RECT 0.684 15.608 0.756 15.64 ;
  LAYER M2 ;
        RECT 0.08 15.608 0.72 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.704 18.528 0.736 18.6 ;
  LAYER M2 ;
        RECT 0.684 18.548 0.756 18.58 ;
  LAYER M2 ;
        RECT 0.08 18.548 0.72 18.58 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M1 ;
        RECT 0.704 21.468 0.736 21.54 ;
  LAYER M2 ;
        RECT 0.684 21.488 0.756 21.52 ;
  LAYER M2 ;
        RECT 0.08 21.488 0.72 21.52 ;
  LAYER M1 ;
        RECT 0.064 21.468 0.096 21.54 ;
  LAYER M2 ;
        RECT 0.044 21.488 0.116 21.52 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.588 ;
  LAYER M1 ;
        RECT 0.064 0.588 0.096 21.504 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 0.96 ;
  LAYER M2 ;
        RECT 7.084 0.908 7.156 0.94 ;
  LAYER M1 ;
        RECT 7.104 0.756 7.136 0.924 ;
  LAYER M1 ;
        RECT 7.104 0.72 7.136 0.792 ;
  LAYER M2 ;
        RECT 7.084 0.74 7.156 0.772 ;
  LAYER M2 ;
        RECT 7.12 0.74 9.68 0.772 ;
  LAYER M1 ;
        RECT 9.664 0.72 9.696 0.792 ;
  LAYER M2 ;
        RECT 9.644 0.74 9.716 0.772 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 3.9 ;
  LAYER M2 ;
        RECT 7.084 3.848 7.156 3.88 ;
  LAYER M1 ;
        RECT 7.104 3.696 7.136 3.864 ;
  LAYER M1 ;
        RECT 7.104 3.66 7.136 3.732 ;
  LAYER M2 ;
        RECT 7.084 3.68 7.156 3.712 ;
  LAYER M2 ;
        RECT 7.12 3.68 9.68 3.712 ;
  LAYER M1 ;
        RECT 9.664 3.66 9.696 3.732 ;
  LAYER M2 ;
        RECT 9.644 3.68 9.716 3.712 ;
  LAYER M1 ;
        RECT 7.104 6.768 7.136 6.84 ;
  LAYER M2 ;
        RECT 7.084 6.788 7.156 6.82 ;
  LAYER M1 ;
        RECT 7.104 6.636 7.136 6.804 ;
  LAYER M1 ;
        RECT 7.104 6.6 7.136 6.672 ;
  LAYER M2 ;
        RECT 7.084 6.62 7.156 6.652 ;
  LAYER M2 ;
        RECT 7.12 6.62 9.68 6.652 ;
  LAYER M1 ;
        RECT 9.664 6.6 9.696 6.672 ;
  LAYER M2 ;
        RECT 9.644 6.62 9.716 6.652 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 9.78 ;
  LAYER M2 ;
        RECT 7.084 9.728 7.156 9.76 ;
  LAYER M1 ;
        RECT 7.104 9.576 7.136 9.744 ;
  LAYER M1 ;
        RECT 7.104 9.54 7.136 9.612 ;
  LAYER M2 ;
        RECT 7.084 9.56 7.156 9.592 ;
  LAYER M2 ;
        RECT 7.12 9.56 9.68 9.592 ;
  LAYER M1 ;
        RECT 9.664 9.54 9.696 9.612 ;
  LAYER M2 ;
        RECT 9.644 9.56 9.716 9.592 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 12.72 ;
  LAYER M2 ;
        RECT 7.084 12.668 7.156 12.7 ;
  LAYER M1 ;
        RECT 7.104 12.516 7.136 12.684 ;
  LAYER M1 ;
        RECT 7.104 12.48 7.136 12.552 ;
  LAYER M2 ;
        RECT 7.084 12.5 7.156 12.532 ;
  LAYER M2 ;
        RECT 7.12 12.5 9.68 12.532 ;
  LAYER M1 ;
        RECT 9.664 12.48 9.696 12.552 ;
  LAYER M2 ;
        RECT 9.644 12.5 9.716 12.532 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 15.66 ;
  LAYER M2 ;
        RECT 7.084 15.608 7.156 15.64 ;
  LAYER M1 ;
        RECT 7.104 15.456 7.136 15.624 ;
  LAYER M1 ;
        RECT 7.104 15.42 7.136 15.492 ;
  LAYER M2 ;
        RECT 7.084 15.44 7.156 15.472 ;
  LAYER M2 ;
        RECT 7.12 15.44 9.68 15.472 ;
  LAYER M1 ;
        RECT 9.664 15.42 9.696 15.492 ;
  LAYER M2 ;
        RECT 9.644 15.44 9.716 15.472 ;
  LAYER M1 ;
        RECT 7.104 18.528 7.136 18.6 ;
  LAYER M2 ;
        RECT 7.084 18.548 7.156 18.58 ;
  LAYER M1 ;
        RECT 7.104 18.396 7.136 18.564 ;
  LAYER M1 ;
        RECT 7.104 18.36 7.136 18.432 ;
  LAYER M2 ;
        RECT 7.084 18.38 7.156 18.412 ;
  LAYER M2 ;
        RECT 7.12 18.38 9.68 18.412 ;
  LAYER M1 ;
        RECT 9.664 18.36 9.696 18.432 ;
  LAYER M2 ;
        RECT 9.644 18.38 9.716 18.412 ;
  LAYER M1 ;
        RECT 7.104 21.468 7.136 21.54 ;
  LAYER M2 ;
        RECT 7.084 21.488 7.156 21.52 ;
  LAYER M1 ;
        RECT 7.104 21.336 7.136 21.504 ;
  LAYER M1 ;
        RECT 7.104 21.3 7.136 21.372 ;
  LAYER M2 ;
        RECT 7.084 21.32 7.156 21.352 ;
  LAYER M2 ;
        RECT 7.12 21.32 9.68 21.352 ;
  LAYER M1 ;
        RECT 9.664 21.3 9.696 21.372 ;
  LAYER M2 ;
        RECT 9.644 21.32 9.716 21.352 ;
  LAYER M1 ;
        RECT 9.664 0.048 9.696 0.12 ;
  LAYER M2 ;
        RECT 9.644 0.068 9.716 0.1 ;
  LAYER M1 ;
        RECT 9.664 0.084 9.696 0.588 ;
  LAYER M1 ;
        RECT 9.664 0.588 9.696 21.336 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.68 0.1 ;
  LAYER M1 ;
        RECT 3.904 0.888 3.936 0.96 ;
  LAYER M2 ;
        RECT 3.884 0.908 3.956 0.94 ;
  LAYER M2 ;
        RECT 0.72 0.908 3.92 0.94 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 0.96 ;
  LAYER M2 ;
        RECT 0.684 0.908 0.756 0.94 ;
  LAYER M1 ;
        RECT 3.904 21.468 3.936 21.54 ;
  LAYER M2 ;
        RECT 3.884 21.488 3.956 21.52 ;
  LAYER M2 ;
        RECT 0.72 21.488 3.92 21.52 ;
  LAYER M1 ;
        RECT 0.704 21.468 0.736 21.54 ;
  LAYER M2 ;
        RECT 0.684 21.488 0.756 21.52 ;
  LAYER M1 ;
        RECT 6.304 15.084 6.336 15.156 ;
  LAYER M2 ;
        RECT 6.284 15.104 6.356 15.136 ;
  LAYER M2 ;
        RECT 3.6 15.104 6.32 15.136 ;
  LAYER M1 ;
        RECT 3.584 15.084 3.616 15.156 ;
  LAYER M2 ;
        RECT 3.564 15.104 3.636 15.136 ;
  LAYER M1 ;
        RECT 6.304 9.204 6.336 9.276 ;
  LAYER M2 ;
        RECT 6.284 9.224 6.356 9.256 ;
  LAYER M2 ;
        RECT 3.6 9.224 6.32 9.256 ;
  LAYER M1 ;
        RECT 3.584 9.204 3.616 9.276 ;
  LAYER M2 ;
        RECT 3.564 9.224 3.636 9.256 ;
  LAYER M1 ;
        RECT 6.304 18.024 6.336 18.096 ;
  LAYER M2 ;
        RECT 6.284 18.044 6.356 18.076 ;
  LAYER M2 ;
        RECT 3.6 18.044 6.32 18.076 ;
  LAYER M1 ;
        RECT 3.584 18.024 3.616 18.096 ;
  LAYER M2 ;
        RECT 3.564 18.044 3.636 18.076 ;
  LAYER M1 ;
        RECT 3.584 24.408 3.616 24.48 ;
  LAYER M2 ;
        RECT 3.564 24.428 3.636 24.46 ;
  LAYER M1 ;
        RECT 3.584 24.276 3.616 24.444 ;
  LAYER M1 ;
        RECT 3.584 9.24 3.616 24.276 ;
  LAYER M1 ;
        RECT 6.304 15.084 6.336 15.156 ;
  LAYER M2 ;
        RECT 6.284 15.104 6.356 15.136 ;
  LAYER M1 ;
        RECT 6.304 15.12 6.336 15.288 ;
  LAYER M1 ;
        RECT 6.304 15.252 6.336 15.324 ;
  LAYER M2 ;
        RECT 6.284 15.272 6.356 15.304 ;
  LAYER M2 ;
        RECT 6.32 15.272 6.8 15.304 ;
  LAYER M1 ;
        RECT 6.784 15.252 6.816 15.324 ;
  LAYER M2 ;
        RECT 6.764 15.272 6.836 15.304 ;
  LAYER M1 ;
        RECT 6.304 9.204 6.336 9.276 ;
  LAYER M2 ;
        RECT 6.284 9.224 6.356 9.256 ;
  LAYER M1 ;
        RECT 6.304 9.24 6.336 9.408 ;
  LAYER M1 ;
        RECT 6.304 9.372 6.336 9.444 ;
  LAYER M2 ;
        RECT 6.284 9.392 6.356 9.424 ;
  LAYER M2 ;
        RECT 6.32 9.392 6.8 9.424 ;
  LAYER M1 ;
        RECT 6.784 9.372 6.816 9.444 ;
  LAYER M2 ;
        RECT 6.764 9.392 6.836 9.424 ;
  LAYER M1 ;
        RECT 6.304 18.024 6.336 18.096 ;
  LAYER M2 ;
        RECT 6.284 18.044 6.356 18.076 ;
  LAYER M1 ;
        RECT 6.304 18.06 6.336 18.228 ;
  LAYER M1 ;
        RECT 6.304 18.192 6.336 18.264 ;
  LAYER M2 ;
        RECT 6.284 18.212 6.356 18.244 ;
  LAYER M2 ;
        RECT 6.32 18.212 6.8 18.244 ;
  LAYER M1 ;
        RECT 6.784 18.192 6.816 18.264 ;
  LAYER M2 ;
        RECT 6.764 18.212 6.836 18.244 ;
  LAYER M1 ;
        RECT 6.784 24.408 6.816 24.48 ;
  LAYER M2 ;
        RECT 6.764 24.428 6.836 24.46 ;
  LAYER M1 ;
        RECT 6.784 24.276 6.816 24.444 ;
  LAYER M1 ;
        RECT 6.784 9.408 6.816 24.276 ;
  LAYER M2 ;
        RECT 3.6 24.428 6.8 24.46 ;
  LAYER M1 ;
        RECT 6.304 12.144 6.336 12.216 ;
  LAYER M2 ;
        RECT 6.284 12.164 6.356 12.196 ;
  LAYER M2 ;
        RECT 3.76 12.164 6.32 12.196 ;
  LAYER M1 ;
        RECT 3.744 12.144 3.776 12.216 ;
  LAYER M2 ;
        RECT 3.724 12.164 3.796 12.196 ;
  LAYER M1 ;
        RECT 6.304 6.264 6.336 6.336 ;
  LAYER M2 ;
        RECT 6.284 6.284 6.356 6.316 ;
  LAYER M2 ;
        RECT 3.76 6.284 6.32 6.316 ;
  LAYER M1 ;
        RECT 3.744 6.264 3.776 6.336 ;
  LAYER M2 ;
        RECT 3.724 6.284 3.796 6.316 ;
  LAYER M1 ;
        RECT 6.304 20.964 6.336 21.036 ;
  LAYER M2 ;
        RECT 6.284 20.984 6.356 21.016 ;
  LAYER M2 ;
        RECT 3.76 20.984 6.32 21.016 ;
  LAYER M1 ;
        RECT 3.744 20.964 3.776 21.036 ;
  LAYER M2 ;
        RECT 3.724 20.984 3.796 21.016 ;
  LAYER M1 ;
        RECT 3.744 24.576 3.776 24.648 ;
  LAYER M2 ;
        RECT 3.724 24.596 3.796 24.628 ;
  LAYER M1 ;
        RECT 3.744 24.276 3.776 24.612 ;
  LAYER M1 ;
        RECT 3.744 6.3 3.776 24.276 ;
  LAYER M1 ;
        RECT 6.304 12.144 6.336 12.216 ;
  LAYER M2 ;
        RECT 6.284 12.164 6.356 12.196 ;
  LAYER M1 ;
        RECT 6.304 12.18 6.336 12.348 ;
  LAYER M1 ;
        RECT 6.304 12.312 6.336 12.384 ;
  LAYER M2 ;
        RECT 6.284 12.332 6.356 12.364 ;
  LAYER M2 ;
        RECT 6.32 12.332 6.96 12.364 ;
  LAYER M1 ;
        RECT 6.944 12.312 6.976 12.384 ;
  LAYER M2 ;
        RECT 6.924 12.332 6.996 12.364 ;
  LAYER M1 ;
        RECT 6.304 6.264 6.336 6.336 ;
  LAYER M2 ;
        RECT 6.284 6.284 6.356 6.316 ;
  LAYER M1 ;
        RECT 6.304 6.3 6.336 6.468 ;
  LAYER M1 ;
        RECT 6.304 6.432 6.336 6.504 ;
  LAYER M2 ;
        RECT 6.284 6.452 6.356 6.484 ;
  LAYER M2 ;
        RECT 6.32 6.452 6.96 6.484 ;
  LAYER M1 ;
        RECT 6.944 6.432 6.976 6.504 ;
  LAYER M2 ;
        RECT 6.924 6.452 6.996 6.484 ;
  LAYER M1 ;
        RECT 6.304 20.964 6.336 21.036 ;
  LAYER M2 ;
        RECT 6.284 20.984 6.356 21.016 ;
  LAYER M1 ;
        RECT 6.304 21 6.336 21.168 ;
  LAYER M1 ;
        RECT 6.304 21.132 6.336 21.204 ;
  LAYER M2 ;
        RECT 6.284 21.152 6.356 21.184 ;
  LAYER M2 ;
        RECT 6.32 21.152 6.96 21.184 ;
  LAYER M1 ;
        RECT 6.944 21.132 6.976 21.204 ;
  LAYER M2 ;
        RECT 6.924 21.152 6.996 21.184 ;
  LAYER M1 ;
        RECT 6.944 24.576 6.976 24.648 ;
  LAYER M2 ;
        RECT 6.924 24.596 6.996 24.628 ;
  LAYER M1 ;
        RECT 6.944 24.276 6.976 24.612 ;
  LAYER M1 ;
        RECT 6.944 6.468 6.976 24.276 ;
  LAYER M2 ;
        RECT 3.76 24.596 6.96 24.628 ;
  LAYER M1 ;
        RECT 3.104 3.324 3.136 3.396 ;
  LAYER M2 ;
        RECT 3.084 3.344 3.156 3.376 ;
  LAYER M2 ;
        RECT 0.24 3.344 3.12 3.376 ;
  LAYER M1 ;
        RECT 0.224 3.324 0.256 3.396 ;
  LAYER M2 ;
        RECT 0.204 3.344 0.276 3.376 ;
  LAYER M1 ;
        RECT 3.104 6.264 3.136 6.336 ;
  LAYER M2 ;
        RECT 3.084 6.284 3.156 6.316 ;
  LAYER M2 ;
        RECT 0.24 6.284 3.12 6.316 ;
  LAYER M1 ;
        RECT 0.224 6.264 0.256 6.336 ;
  LAYER M2 ;
        RECT 0.204 6.284 0.276 6.316 ;
  LAYER M1 ;
        RECT 3.104 9.204 3.136 9.276 ;
  LAYER M2 ;
        RECT 3.084 9.224 3.156 9.256 ;
  LAYER M2 ;
        RECT 0.24 9.224 3.12 9.256 ;
  LAYER M1 ;
        RECT 0.224 9.204 0.256 9.276 ;
  LAYER M2 ;
        RECT 0.204 9.224 0.276 9.256 ;
  LAYER M1 ;
        RECT 3.104 12.144 3.136 12.216 ;
  LAYER M2 ;
        RECT 3.084 12.164 3.156 12.196 ;
  LAYER M2 ;
        RECT 0.24 12.164 3.12 12.196 ;
  LAYER M1 ;
        RECT 0.224 12.144 0.256 12.216 ;
  LAYER M2 ;
        RECT 0.204 12.164 0.276 12.196 ;
  LAYER M1 ;
        RECT 3.104 15.084 3.136 15.156 ;
  LAYER M2 ;
        RECT 3.084 15.104 3.156 15.136 ;
  LAYER M2 ;
        RECT 0.24 15.104 3.12 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.084 0.256 15.156 ;
  LAYER M2 ;
        RECT 0.204 15.104 0.276 15.136 ;
  LAYER M1 ;
        RECT 3.104 18.024 3.136 18.096 ;
  LAYER M2 ;
        RECT 3.084 18.044 3.156 18.076 ;
  LAYER M2 ;
        RECT 0.24 18.044 3.12 18.076 ;
  LAYER M1 ;
        RECT 0.224 18.024 0.256 18.096 ;
  LAYER M2 ;
        RECT 0.204 18.044 0.276 18.076 ;
  LAYER M1 ;
        RECT 3.104 20.964 3.136 21.036 ;
  LAYER M2 ;
        RECT 3.084 20.984 3.156 21.016 ;
  LAYER M2 ;
        RECT 0.24 20.984 3.12 21.016 ;
  LAYER M1 ;
        RECT 0.224 20.964 0.256 21.036 ;
  LAYER M2 ;
        RECT 0.204 20.984 0.276 21.016 ;
  LAYER M1 ;
        RECT 3.104 23.904 3.136 23.976 ;
  LAYER M2 ;
        RECT 3.084 23.924 3.156 23.956 ;
  LAYER M2 ;
        RECT 0.24 23.924 3.12 23.956 ;
  LAYER M1 ;
        RECT 0.224 23.904 0.256 23.976 ;
  LAYER M2 ;
        RECT 0.204 23.924 0.276 23.956 ;
  LAYER M1 ;
        RECT 0.224 24.744 0.256 24.816 ;
  LAYER M2 ;
        RECT 0.204 24.764 0.276 24.796 ;
  LAYER M1 ;
        RECT 0.224 24.276 0.256 24.78 ;
  LAYER M1 ;
        RECT 0.224 3.36 0.256 24.276 ;
  LAYER M1 ;
        RECT 9.504 3.324 9.536 3.396 ;
  LAYER M2 ;
        RECT 9.484 3.344 9.556 3.376 ;
  LAYER M1 ;
        RECT 9.504 3.36 9.536 3.528 ;
  LAYER M1 ;
        RECT 9.504 3.492 9.536 3.564 ;
  LAYER M2 ;
        RECT 9.484 3.512 9.556 3.544 ;
  LAYER M2 ;
        RECT 9.52 3.512 9.84 3.544 ;
  LAYER M1 ;
        RECT 9.824 3.492 9.856 3.564 ;
  LAYER M2 ;
        RECT 9.804 3.512 9.876 3.544 ;
  LAYER M1 ;
        RECT 9.504 6.264 9.536 6.336 ;
  LAYER M2 ;
        RECT 9.484 6.284 9.556 6.316 ;
  LAYER M1 ;
        RECT 9.504 6.3 9.536 6.468 ;
  LAYER M1 ;
        RECT 9.504 6.432 9.536 6.504 ;
  LAYER M2 ;
        RECT 9.484 6.452 9.556 6.484 ;
  LAYER M2 ;
        RECT 9.52 6.452 9.84 6.484 ;
  LAYER M1 ;
        RECT 9.824 6.432 9.856 6.504 ;
  LAYER M2 ;
        RECT 9.804 6.452 9.876 6.484 ;
  LAYER M1 ;
        RECT 9.504 9.204 9.536 9.276 ;
  LAYER M2 ;
        RECT 9.484 9.224 9.556 9.256 ;
  LAYER M1 ;
        RECT 9.504 9.24 9.536 9.408 ;
  LAYER M1 ;
        RECT 9.504 9.372 9.536 9.444 ;
  LAYER M2 ;
        RECT 9.484 9.392 9.556 9.424 ;
  LAYER M2 ;
        RECT 9.52 9.392 9.84 9.424 ;
  LAYER M1 ;
        RECT 9.824 9.372 9.856 9.444 ;
  LAYER M2 ;
        RECT 9.804 9.392 9.876 9.424 ;
  LAYER M1 ;
        RECT 9.504 12.144 9.536 12.216 ;
  LAYER M2 ;
        RECT 9.484 12.164 9.556 12.196 ;
  LAYER M1 ;
        RECT 9.504 12.18 9.536 12.348 ;
  LAYER M1 ;
        RECT 9.504 12.312 9.536 12.384 ;
  LAYER M2 ;
        RECT 9.484 12.332 9.556 12.364 ;
  LAYER M2 ;
        RECT 9.52 12.332 9.84 12.364 ;
  LAYER M1 ;
        RECT 9.824 12.312 9.856 12.384 ;
  LAYER M2 ;
        RECT 9.804 12.332 9.876 12.364 ;
  LAYER M1 ;
        RECT 9.504 15.084 9.536 15.156 ;
  LAYER M2 ;
        RECT 9.484 15.104 9.556 15.136 ;
  LAYER M1 ;
        RECT 9.504 15.12 9.536 15.288 ;
  LAYER M1 ;
        RECT 9.504 15.252 9.536 15.324 ;
  LAYER M2 ;
        RECT 9.484 15.272 9.556 15.304 ;
  LAYER M2 ;
        RECT 9.52 15.272 9.84 15.304 ;
  LAYER M1 ;
        RECT 9.824 15.252 9.856 15.324 ;
  LAYER M2 ;
        RECT 9.804 15.272 9.876 15.304 ;
  LAYER M1 ;
        RECT 9.504 18.024 9.536 18.096 ;
  LAYER M2 ;
        RECT 9.484 18.044 9.556 18.076 ;
  LAYER M1 ;
        RECT 9.504 18.06 9.536 18.228 ;
  LAYER M1 ;
        RECT 9.504 18.192 9.536 18.264 ;
  LAYER M2 ;
        RECT 9.484 18.212 9.556 18.244 ;
  LAYER M2 ;
        RECT 9.52 18.212 9.84 18.244 ;
  LAYER M1 ;
        RECT 9.824 18.192 9.856 18.264 ;
  LAYER M2 ;
        RECT 9.804 18.212 9.876 18.244 ;
  LAYER M1 ;
        RECT 9.504 20.964 9.536 21.036 ;
  LAYER M2 ;
        RECT 9.484 20.984 9.556 21.016 ;
  LAYER M1 ;
        RECT 9.504 21 9.536 21.168 ;
  LAYER M1 ;
        RECT 9.504 21.132 9.536 21.204 ;
  LAYER M2 ;
        RECT 9.484 21.152 9.556 21.184 ;
  LAYER M2 ;
        RECT 9.52 21.152 9.84 21.184 ;
  LAYER M1 ;
        RECT 9.824 21.132 9.856 21.204 ;
  LAYER M2 ;
        RECT 9.804 21.152 9.876 21.184 ;
  LAYER M1 ;
        RECT 9.504 23.904 9.536 23.976 ;
  LAYER M2 ;
        RECT 9.484 23.924 9.556 23.956 ;
  LAYER M1 ;
        RECT 9.504 23.94 9.536 24.108 ;
  LAYER M1 ;
        RECT 9.504 24.072 9.536 24.144 ;
  LAYER M2 ;
        RECT 9.484 24.092 9.556 24.124 ;
  LAYER M2 ;
        RECT 9.52 24.092 9.84 24.124 ;
  LAYER M1 ;
        RECT 9.824 24.072 9.856 24.144 ;
  LAYER M2 ;
        RECT 9.804 24.092 9.876 24.124 ;
  LAYER M1 ;
        RECT 9.824 24.744 9.856 24.816 ;
  LAYER M2 ;
        RECT 9.804 24.764 9.876 24.796 ;
  LAYER M1 ;
        RECT 9.824 24.276 9.856 24.78 ;
  LAYER M1 ;
        RECT 9.824 3.528 9.856 24.276 ;
  LAYER M2 ;
        RECT 0.24 24.764 9.84 24.796 ;
  LAYER M1 ;
        RECT 6.304 3.324 6.336 3.396 ;
  LAYER M2 ;
        RECT 6.284 3.344 6.356 3.376 ;
  LAYER M2 ;
        RECT 3.12 3.344 6.32 3.376 ;
  LAYER M1 ;
        RECT 3.104 3.324 3.136 3.396 ;
  LAYER M2 ;
        RECT 3.084 3.344 3.156 3.376 ;
  LAYER M1 ;
        RECT 6.304 23.904 6.336 23.976 ;
  LAYER M2 ;
        RECT 6.284 23.924 6.356 23.956 ;
  LAYER M2 ;
        RECT 3.12 23.924 6.32 23.956 ;
  LAYER M1 ;
        RECT 3.104 23.904 3.136 23.976 ;
  LAYER M2 ;
        RECT 3.084 23.924 3.156 23.956 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M1 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M1 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M1 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M1 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M1 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M1 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M1 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M1 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M1 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M1 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M1 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M1 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M1 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M1 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M1 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M1 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M1 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M1 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M1 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M1 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M1 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M1 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M1 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M1 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M1 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M1 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M1 ;
        RECT 2.432 0.888 2.464 3.396 ;
  LAYER M1 ;
        RECT 2.496 0.888 2.528 3.396 ;
  LAYER M1 ;
        RECT 2.56 0.888 2.592 3.396 ;
  LAYER M1 ;
        RECT 2.624 0.888 2.656 3.396 ;
  LAYER M1 ;
        RECT 2.688 0.888 2.72 3.396 ;
  LAYER M1 ;
        RECT 2.752 0.888 2.784 3.396 ;
  LAYER M1 ;
        RECT 2.816 0.888 2.848 3.396 ;
  LAYER M1 ;
        RECT 2.88 0.888 2.912 3.396 ;
  LAYER M1 ;
        RECT 2.944 0.888 2.976 3.396 ;
  LAYER M1 ;
        RECT 3.008 0.888 3.04 3.396 ;
  LAYER M2 ;
        RECT 0.684 0.972 3.156 1.004 ;
  LAYER M2 ;
        RECT 0.684 1.036 3.156 1.068 ;
  LAYER M2 ;
        RECT 0.684 1.1 3.156 1.132 ;
  LAYER M2 ;
        RECT 0.684 1.164 3.156 1.196 ;
  LAYER M2 ;
        RECT 0.684 1.228 3.156 1.26 ;
  LAYER M2 ;
        RECT 0.684 1.292 3.156 1.324 ;
  LAYER M2 ;
        RECT 0.684 1.356 3.156 1.388 ;
  LAYER M2 ;
        RECT 0.684 1.42 3.156 1.452 ;
  LAYER M2 ;
        RECT 0.684 1.484 3.156 1.516 ;
  LAYER M2 ;
        RECT 0.684 1.548 3.156 1.58 ;
  LAYER M2 ;
        RECT 0.684 1.612 3.156 1.644 ;
  LAYER M2 ;
        RECT 0.684 1.676 3.156 1.708 ;
  LAYER M2 ;
        RECT 0.684 1.74 3.156 1.772 ;
  LAYER M2 ;
        RECT 0.684 1.804 3.156 1.836 ;
  LAYER M2 ;
        RECT 0.684 1.868 3.156 1.9 ;
  LAYER M2 ;
        RECT 0.684 1.932 3.156 1.964 ;
  LAYER M2 ;
        RECT 0.684 1.996 3.156 2.028 ;
  LAYER M2 ;
        RECT 0.684 2.06 3.156 2.092 ;
  LAYER M2 ;
        RECT 0.684 2.124 3.156 2.156 ;
  LAYER M2 ;
        RECT 0.684 2.188 3.156 2.22 ;
  LAYER M2 ;
        RECT 0.684 2.252 3.156 2.284 ;
  LAYER M2 ;
        RECT 0.684 2.316 3.156 2.348 ;
  LAYER M2 ;
        RECT 0.684 2.38 3.156 2.412 ;
  LAYER M2 ;
        RECT 0.684 2.444 3.156 2.476 ;
  LAYER M2 ;
        RECT 0.684 2.508 3.156 2.54 ;
  LAYER M2 ;
        RECT 0.684 2.572 3.156 2.604 ;
  LAYER M2 ;
        RECT 0.684 2.636 3.156 2.668 ;
  LAYER M2 ;
        RECT 0.684 2.7 3.156 2.732 ;
  LAYER M2 ;
        RECT 0.684 2.764 3.156 2.796 ;
  LAYER M2 ;
        RECT 0.684 2.828 3.156 2.86 ;
  LAYER M2 ;
        RECT 0.684 2.892 3.156 2.924 ;
  LAYER M2 ;
        RECT 0.684 2.956 3.156 2.988 ;
  LAYER M2 ;
        RECT 0.684 3.02 3.156 3.052 ;
  LAYER M2 ;
        RECT 0.684 3.084 3.156 3.116 ;
  LAYER M2 ;
        RECT 0.684 3.148 3.156 3.18 ;
  LAYER M2 ;
        RECT 0.684 3.212 3.156 3.244 ;
  LAYER M3 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M3 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M3 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M3 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M3 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M3 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M3 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M3 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M3 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M3 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M3 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M3 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M3 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M3 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M3 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M3 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M3 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M3 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M3 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M3 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M3 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M3 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M3 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M3 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M3 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M3 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M3 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M3 ;
        RECT 2.432 0.888 2.464 3.396 ;
  LAYER M3 ;
        RECT 2.496 0.888 2.528 3.396 ;
  LAYER M3 ;
        RECT 2.56 0.888 2.592 3.396 ;
  LAYER M3 ;
        RECT 2.624 0.888 2.656 3.396 ;
  LAYER M3 ;
        RECT 2.688 0.888 2.72 3.396 ;
  LAYER M3 ;
        RECT 2.752 0.888 2.784 3.396 ;
  LAYER M3 ;
        RECT 2.816 0.888 2.848 3.396 ;
  LAYER M3 ;
        RECT 2.88 0.888 2.912 3.396 ;
  LAYER M3 ;
        RECT 2.944 0.888 2.976 3.396 ;
  LAYER M3 ;
        RECT 3.008 0.888 3.04 3.396 ;
  LAYER M3 ;
        RECT 3.104 0.888 3.136 3.396 ;
  LAYER M1 ;
        RECT 0.719 0.924 0.721 3.36 ;
  LAYER M1 ;
        RECT 0.799 0.924 0.801 3.36 ;
  LAYER M1 ;
        RECT 0.879 0.924 0.881 3.36 ;
  LAYER M1 ;
        RECT 0.959 0.924 0.961 3.36 ;
  LAYER M1 ;
        RECT 1.039 0.924 1.041 3.36 ;
  LAYER M1 ;
        RECT 1.119 0.924 1.121 3.36 ;
  LAYER M1 ;
        RECT 1.199 0.924 1.201 3.36 ;
  LAYER M1 ;
        RECT 1.279 0.924 1.281 3.36 ;
  LAYER M1 ;
        RECT 1.359 0.924 1.361 3.36 ;
  LAYER M1 ;
        RECT 1.439 0.924 1.441 3.36 ;
  LAYER M1 ;
        RECT 1.519 0.924 1.521 3.36 ;
  LAYER M1 ;
        RECT 1.599 0.924 1.601 3.36 ;
  LAYER M1 ;
        RECT 1.679 0.924 1.681 3.36 ;
  LAYER M1 ;
        RECT 1.759 0.924 1.761 3.36 ;
  LAYER M1 ;
        RECT 1.839 0.924 1.841 3.36 ;
  LAYER M1 ;
        RECT 1.919 0.924 1.921 3.36 ;
  LAYER M1 ;
        RECT 1.999 0.924 2.001 3.36 ;
  LAYER M1 ;
        RECT 2.079 0.924 2.081 3.36 ;
  LAYER M1 ;
        RECT 2.159 0.924 2.161 3.36 ;
  LAYER M1 ;
        RECT 2.239 0.924 2.241 3.36 ;
  LAYER M1 ;
        RECT 2.319 0.924 2.321 3.36 ;
  LAYER M1 ;
        RECT 2.399 0.924 2.401 3.36 ;
  LAYER M1 ;
        RECT 2.479 0.924 2.481 3.36 ;
  LAYER M1 ;
        RECT 2.559 0.924 2.561 3.36 ;
  LAYER M1 ;
        RECT 2.639 0.924 2.641 3.36 ;
  LAYER M1 ;
        RECT 2.719 0.924 2.721 3.36 ;
  LAYER M1 ;
        RECT 2.799 0.924 2.801 3.36 ;
  LAYER M1 ;
        RECT 2.879 0.924 2.881 3.36 ;
  LAYER M1 ;
        RECT 2.959 0.924 2.961 3.36 ;
  LAYER M1 ;
        RECT 3.039 0.924 3.041 3.36 ;
  LAYER M2 ;
        RECT 0.72 0.923 3.12 0.925 ;
  LAYER M2 ;
        RECT 0.72 1.007 3.12 1.009 ;
  LAYER M2 ;
        RECT 0.72 1.091 3.12 1.093 ;
  LAYER M2 ;
        RECT 0.72 1.175 3.12 1.177 ;
  LAYER M2 ;
        RECT 0.72 1.259 3.12 1.261 ;
  LAYER M2 ;
        RECT 0.72 1.343 3.12 1.345 ;
  LAYER M2 ;
        RECT 0.72 1.427 3.12 1.429 ;
  LAYER M2 ;
        RECT 0.72 1.511 3.12 1.513 ;
  LAYER M2 ;
        RECT 0.72 1.595 3.12 1.597 ;
  LAYER M2 ;
        RECT 0.72 1.679 3.12 1.681 ;
  LAYER M2 ;
        RECT 0.72 1.763 3.12 1.765 ;
  LAYER M2 ;
        RECT 0.72 1.847 3.12 1.849 ;
  LAYER M2 ;
        RECT 0.72 1.9305 3.12 1.9325 ;
  LAYER M2 ;
        RECT 0.72 2.015 3.12 2.017 ;
  LAYER M2 ;
        RECT 0.72 2.099 3.12 2.101 ;
  LAYER M2 ;
        RECT 0.72 2.183 3.12 2.185 ;
  LAYER M2 ;
        RECT 0.72 2.267 3.12 2.269 ;
  LAYER M2 ;
        RECT 0.72 2.351 3.12 2.353 ;
  LAYER M2 ;
        RECT 0.72 2.435 3.12 2.437 ;
  LAYER M2 ;
        RECT 0.72 2.519 3.12 2.521 ;
  LAYER M2 ;
        RECT 0.72 2.603 3.12 2.605 ;
  LAYER M2 ;
        RECT 0.72 2.687 3.12 2.689 ;
  LAYER M2 ;
        RECT 0.72 2.771 3.12 2.773 ;
  LAYER M2 ;
        RECT 0.72 2.855 3.12 2.857 ;
  LAYER M2 ;
        RECT 0.72 2.939 3.12 2.941 ;
  LAYER M2 ;
        RECT 0.72 3.023 3.12 3.025 ;
  LAYER M2 ;
        RECT 0.72 3.107 3.12 3.109 ;
  LAYER M2 ;
        RECT 0.72 3.191 3.12 3.193 ;
  LAYER M2 ;
        RECT 0.72 3.275 3.12 3.277 ;
  LAYER M1 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M1 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M1 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M1 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M1 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M1 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M1 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M1 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M1 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M1 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M1 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M1 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M1 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M1 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M1 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M1 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M1 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M1 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M1 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M1 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M1 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M1 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M1 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M1 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M1 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M1 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M1 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M1 ;
        RECT 2.432 3.828 2.464 6.336 ;
  LAYER M1 ;
        RECT 2.496 3.828 2.528 6.336 ;
  LAYER M1 ;
        RECT 2.56 3.828 2.592 6.336 ;
  LAYER M1 ;
        RECT 2.624 3.828 2.656 6.336 ;
  LAYER M1 ;
        RECT 2.688 3.828 2.72 6.336 ;
  LAYER M1 ;
        RECT 2.752 3.828 2.784 6.336 ;
  LAYER M1 ;
        RECT 2.816 3.828 2.848 6.336 ;
  LAYER M1 ;
        RECT 2.88 3.828 2.912 6.336 ;
  LAYER M1 ;
        RECT 2.944 3.828 2.976 6.336 ;
  LAYER M1 ;
        RECT 3.008 3.828 3.04 6.336 ;
  LAYER M2 ;
        RECT 0.684 3.912 3.156 3.944 ;
  LAYER M2 ;
        RECT 0.684 3.976 3.156 4.008 ;
  LAYER M2 ;
        RECT 0.684 4.04 3.156 4.072 ;
  LAYER M2 ;
        RECT 0.684 4.104 3.156 4.136 ;
  LAYER M2 ;
        RECT 0.684 4.168 3.156 4.2 ;
  LAYER M2 ;
        RECT 0.684 4.232 3.156 4.264 ;
  LAYER M2 ;
        RECT 0.684 4.296 3.156 4.328 ;
  LAYER M2 ;
        RECT 0.684 4.36 3.156 4.392 ;
  LAYER M2 ;
        RECT 0.684 4.424 3.156 4.456 ;
  LAYER M2 ;
        RECT 0.684 4.488 3.156 4.52 ;
  LAYER M2 ;
        RECT 0.684 4.552 3.156 4.584 ;
  LAYER M2 ;
        RECT 0.684 4.616 3.156 4.648 ;
  LAYER M2 ;
        RECT 0.684 4.68 3.156 4.712 ;
  LAYER M2 ;
        RECT 0.684 4.744 3.156 4.776 ;
  LAYER M2 ;
        RECT 0.684 4.808 3.156 4.84 ;
  LAYER M2 ;
        RECT 0.684 4.872 3.156 4.904 ;
  LAYER M2 ;
        RECT 0.684 4.936 3.156 4.968 ;
  LAYER M2 ;
        RECT 0.684 5 3.156 5.032 ;
  LAYER M2 ;
        RECT 0.684 5.064 3.156 5.096 ;
  LAYER M2 ;
        RECT 0.684 5.128 3.156 5.16 ;
  LAYER M2 ;
        RECT 0.684 5.192 3.156 5.224 ;
  LAYER M2 ;
        RECT 0.684 5.256 3.156 5.288 ;
  LAYER M2 ;
        RECT 0.684 5.32 3.156 5.352 ;
  LAYER M2 ;
        RECT 0.684 5.384 3.156 5.416 ;
  LAYER M2 ;
        RECT 0.684 5.448 3.156 5.48 ;
  LAYER M2 ;
        RECT 0.684 5.512 3.156 5.544 ;
  LAYER M2 ;
        RECT 0.684 5.576 3.156 5.608 ;
  LAYER M2 ;
        RECT 0.684 5.64 3.156 5.672 ;
  LAYER M2 ;
        RECT 0.684 5.704 3.156 5.736 ;
  LAYER M2 ;
        RECT 0.684 5.768 3.156 5.8 ;
  LAYER M2 ;
        RECT 0.684 5.832 3.156 5.864 ;
  LAYER M2 ;
        RECT 0.684 5.896 3.156 5.928 ;
  LAYER M2 ;
        RECT 0.684 5.96 3.156 5.992 ;
  LAYER M2 ;
        RECT 0.684 6.024 3.156 6.056 ;
  LAYER M2 ;
        RECT 0.684 6.088 3.156 6.12 ;
  LAYER M2 ;
        RECT 0.684 6.152 3.156 6.184 ;
  LAYER M3 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M3 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M3 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M3 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M3 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M3 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M3 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M3 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M3 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M3 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M3 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M3 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M3 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M3 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M3 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M3 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M3 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M3 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M3 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M3 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M3 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M3 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M3 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M3 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M3 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M3 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M3 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M3 ;
        RECT 2.432 3.828 2.464 6.336 ;
  LAYER M3 ;
        RECT 2.496 3.828 2.528 6.336 ;
  LAYER M3 ;
        RECT 2.56 3.828 2.592 6.336 ;
  LAYER M3 ;
        RECT 2.624 3.828 2.656 6.336 ;
  LAYER M3 ;
        RECT 2.688 3.828 2.72 6.336 ;
  LAYER M3 ;
        RECT 2.752 3.828 2.784 6.336 ;
  LAYER M3 ;
        RECT 2.816 3.828 2.848 6.336 ;
  LAYER M3 ;
        RECT 2.88 3.828 2.912 6.336 ;
  LAYER M3 ;
        RECT 2.944 3.828 2.976 6.336 ;
  LAYER M3 ;
        RECT 3.008 3.828 3.04 6.336 ;
  LAYER M3 ;
        RECT 3.104 3.828 3.136 6.336 ;
  LAYER M1 ;
        RECT 0.719 3.864 0.721 6.3 ;
  LAYER M1 ;
        RECT 0.799 3.864 0.801 6.3 ;
  LAYER M1 ;
        RECT 0.879 3.864 0.881 6.3 ;
  LAYER M1 ;
        RECT 0.959 3.864 0.961 6.3 ;
  LAYER M1 ;
        RECT 1.039 3.864 1.041 6.3 ;
  LAYER M1 ;
        RECT 1.119 3.864 1.121 6.3 ;
  LAYER M1 ;
        RECT 1.199 3.864 1.201 6.3 ;
  LAYER M1 ;
        RECT 1.279 3.864 1.281 6.3 ;
  LAYER M1 ;
        RECT 1.359 3.864 1.361 6.3 ;
  LAYER M1 ;
        RECT 1.439 3.864 1.441 6.3 ;
  LAYER M1 ;
        RECT 1.519 3.864 1.521 6.3 ;
  LAYER M1 ;
        RECT 1.599 3.864 1.601 6.3 ;
  LAYER M1 ;
        RECT 1.679 3.864 1.681 6.3 ;
  LAYER M1 ;
        RECT 1.759 3.864 1.761 6.3 ;
  LAYER M1 ;
        RECT 1.839 3.864 1.841 6.3 ;
  LAYER M1 ;
        RECT 1.919 3.864 1.921 6.3 ;
  LAYER M1 ;
        RECT 1.999 3.864 2.001 6.3 ;
  LAYER M1 ;
        RECT 2.079 3.864 2.081 6.3 ;
  LAYER M1 ;
        RECT 2.159 3.864 2.161 6.3 ;
  LAYER M1 ;
        RECT 2.239 3.864 2.241 6.3 ;
  LAYER M1 ;
        RECT 2.319 3.864 2.321 6.3 ;
  LAYER M1 ;
        RECT 2.399 3.864 2.401 6.3 ;
  LAYER M1 ;
        RECT 2.479 3.864 2.481 6.3 ;
  LAYER M1 ;
        RECT 2.559 3.864 2.561 6.3 ;
  LAYER M1 ;
        RECT 2.639 3.864 2.641 6.3 ;
  LAYER M1 ;
        RECT 2.719 3.864 2.721 6.3 ;
  LAYER M1 ;
        RECT 2.799 3.864 2.801 6.3 ;
  LAYER M1 ;
        RECT 2.879 3.864 2.881 6.3 ;
  LAYER M1 ;
        RECT 2.959 3.864 2.961 6.3 ;
  LAYER M1 ;
        RECT 3.039 3.864 3.041 6.3 ;
  LAYER M2 ;
        RECT 0.72 3.863 3.12 3.865 ;
  LAYER M2 ;
        RECT 0.72 3.947 3.12 3.949 ;
  LAYER M2 ;
        RECT 0.72 4.031 3.12 4.033 ;
  LAYER M2 ;
        RECT 0.72 4.115 3.12 4.117 ;
  LAYER M2 ;
        RECT 0.72 4.199 3.12 4.201 ;
  LAYER M2 ;
        RECT 0.72 4.283 3.12 4.285 ;
  LAYER M2 ;
        RECT 0.72 4.367 3.12 4.369 ;
  LAYER M2 ;
        RECT 0.72 4.451 3.12 4.453 ;
  LAYER M2 ;
        RECT 0.72 4.535 3.12 4.537 ;
  LAYER M2 ;
        RECT 0.72 4.619 3.12 4.621 ;
  LAYER M2 ;
        RECT 0.72 4.703 3.12 4.705 ;
  LAYER M2 ;
        RECT 0.72 4.787 3.12 4.789 ;
  LAYER M2 ;
        RECT 0.72 4.8705 3.12 4.8725 ;
  LAYER M2 ;
        RECT 0.72 4.955 3.12 4.957 ;
  LAYER M2 ;
        RECT 0.72 5.039 3.12 5.041 ;
  LAYER M2 ;
        RECT 0.72 5.123 3.12 5.125 ;
  LAYER M2 ;
        RECT 0.72 5.207 3.12 5.209 ;
  LAYER M2 ;
        RECT 0.72 5.291 3.12 5.293 ;
  LAYER M2 ;
        RECT 0.72 5.375 3.12 5.377 ;
  LAYER M2 ;
        RECT 0.72 5.459 3.12 5.461 ;
  LAYER M2 ;
        RECT 0.72 5.543 3.12 5.545 ;
  LAYER M2 ;
        RECT 0.72 5.627 3.12 5.629 ;
  LAYER M2 ;
        RECT 0.72 5.711 3.12 5.713 ;
  LAYER M2 ;
        RECT 0.72 5.795 3.12 5.797 ;
  LAYER M2 ;
        RECT 0.72 5.879 3.12 5.881 ;
  LAYER M2 ;
        RECT 0.72 5.963 3.12 5.965 ;
  LAYER M2 ;
        RECT 0.72 6.047 3.12 6.049 ;
  LAYER M2 ;
        RECT 0.72 6.131 3.12 6.133 ;
  LAYER M2 ;
        RECT 0.72 6.215 3.12 6.217 ;
  LAYER M1 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M1 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M1 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M1 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M1 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M1 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M1 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M1 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M1 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M1 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M1 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M1 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M1 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M1 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M1 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M1 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M1 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M1 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M1 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M1 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M1 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M1 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M1 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M1 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M1 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M1 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M1 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M1 ;
        RECT 2.432 6.768 2.464 9.276 ;
  LAYER M1 ;
        RECT 2.496 6.768 2.528 9.276 ;
  LAYER M1 ;
        RECT 2.56 6.768 2.592 9.276 ;
  LAYER M1 ;
        RECT 2.624 6.768 2.656 9.276 ;
  LAYER M1 ;
        RECT 2.688 6.768 2.72 9.276 ;
  LAYER M1 ;
        RECT 2.752 6.768 2.784 9.276 ;
  LAYER M1 ;
        RECT 2.816 6.768 2.848 9.276 ;
  LAYER M1 ;
        RECT 2.88 6.768 2.912 9.276 ;
  LAYER M1 ;
        RECT 2.944 6.768 2.976 9.276 ;
  LAYER M1 ;
        RECT 3.008 6.768 3.04 9.276 ;
  LAYER M2 ;
        RECT 0.684 6.852 3.156 6.884 ;
  LAYER M2 ;
        RECT 0.684 6.916 3.156 6.948 ;
  LAYER M2 ;
        RECT 0.684 6.98 3.156 7.012 ;
  LAYER M2 ;
        RECT 0.684 7.044 3.156 7.076 ;
  LAYER M2 ;
        RECT 0.684 7.108 3.156 7.14 ;
  LAYER M2 ;
        RECT 0.684 7.172 3.156 7.204 ;
  LAYER M2 ;
        RECT 0.684 7.236 3.156 7.268 ;
  LAYER M2 ;
        RECT 0.684 7.3 3.156 7.332 ;
  LAYER M2 ;
        RECT 0.684 7.364 3.156 7.396 ;
  LAYER M2 ;
        RECT 0.684 7.428 3.156 7.46 ;
  LAYER M2 ;
        RECT 0.684 7.492 3.156 7.524 ;
  LAYER M2 ;
        RECT 0.684 7.556 3.156 7.588 ;
  LAYER M2 ;
        RECT 0.684 7.62 3.156 7.652 ;
  LAYER M2 ;
        RECT 0.684 7.684 3.156 7.716 ;
  LAYER M2 ;
        RECT 0.684 7.748 3.156 7.78 ;
  LAYER M2 ;
        RECT 0.684 7.812 3.156 7.844 ;
  LAYER M2 ;
        RECT 0.684 7.876 3.156 7.908 ;
  LAYER M2 ;
        RECT 0.684 7.94 3.156 7.972 ;
  LAYER M2 ;
        RECT 0.684 8.004 3.156 8.036 ;
  LAYER M2 ;
        RECT 0.684 8.068 3.156 8.1 ;
  LAYER M2 ;
        RECT 0.684 8.132 3.156 8.164 ;
  LAYER M2 ;
        RECT 0.684 8.196 3.156 8.228 ;
  LAYER M2 ;
        RECT 0.684 8.26 3.156 8.292 ;
  LAYER M2 ;
        RECT 0.684 8.324 3.156 8.356 ;
  LAYER M2 ;
        RECT 0.684 8.388 3.156 8.42 ;
  LAYER M2 ;
        RECT 0.684 8.452 3.156 8.484 ;
  LAYER M2 ;
        RECT 0.684 8.516 3.156 8.548 ;
  LAYER M2 ;
        RECT 0.684 8.58 3.156 8.612 ;
  LAYER M2 ;
        RECT 0.684 8.644 3.156 8.676 ;
  LAYER M2 ;
        RECT 0.684 8.708 3.156 8.74 ;
  LAYER M2 ;
        RECT 0.684 8.772 3.156 8.804 ;
  LAYER M2 ;
        RECT 0.684 8.836 3.156 8.868 ;
  LAYER M2 ;
        RECT 0.684 8.9 3.156 8.932 ;
  LAYER M2 ;
        RECT 0.684 8.964 3.156 8.996 ;
  LAYER M2 ;
        RECT 0.684 9.028 3.156 9.06 ;
  LAYER M2 ;
        RECT 0.684 9.092 3.156 9.124 ;
  LAYER M3 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M3 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M3 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M3 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M3 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M3 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M3 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M3 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M3 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M3 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M3 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M3 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M3 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M3 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M3 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M3 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M3 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M3 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M3 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M3 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M3 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M3 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M3 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M3 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M3 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M3 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M3 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M3 ;
        RECT 2.432 6.768 2.464 9.276 ;
  LAYER M3 ;
        RECT 2.496 6.768 2.528 9.276 ;
  LAYER M3 ;
        RECT 2.56 6.768 2.592 9.276 ;
  LAYER M3 ;
        RECT 2.624 6.768 2.656 9.276 ;
  LAYER M3 ;
        RECT 2.688 6.768 2.72 9.276 ;
  LAYER M3 ;
        RECT 2.752 6.768 2.784 9.276 ;
  LAYER M3 ;
        RECT 2.816 6.768 2.848 9.276 ;
  LAYER M3 ;
        RECT 2.88 6.768 2.912 9.276 ;
  LAYER M3 ;
        RECT 2.944 6.768 2.976 9.276 ;
  LAYER M3 ;
        RECT 3.008 6.768 3.04 9.276 ;
  LAYER M3 ;
        RECT 3.104 6.768 3.136 9.276 ;
  LAYER M1 ;
        RECT 0.719 6.804 0.721 9.24 ;
  LAYER M1 ;
        RECT 0.799 6.804 0.801 9.24 ;
  LAYER M1 ;
        RECT 0.879 6.804 0.881 9.24 ;
  LAYER M1 ;
        RECT 0.959 6.804 0.961 9.24 ;
  LAYER M1 ;
        RECT 1.039 6.804 1.041 9.24 ;
  LAYER M1 ;
        RECT 1.119 6.804 1.121 9.24 ;
  LAYER M1 ;
        RECT 1.199 6.804 1.201 9.24 ;
  LAYER M1 ;
        RECT 1.279 6.804 1.281 9.24 ;
  LAYER M1 ;
        RECT 1.359 6.804 1.361 9.24 ;
  LAYER M1 ;
        RECT 1.439 6.804 1.441 9.24 ;
  LAYER M1 ;
        RECT 1.519 6.804 1.521 9.24 ;
  LAYER M1 ;
        RECT 1.599 6.804 1.601 9.24 ;
  LAYER M1 ;
        RECT 1.679 6.804 1.681 9.24 ;
  LAYER M1 ;
        RECT 1.759 6.804 1.761 9.24 ;
  LAYER M1 ;
        RECT 1.839 6.804 1.841 9.24 ;
  LAYER M1 ;
        RECT 1.919 6.804 1.921 9.24 ;
  LAYER M1 ;
        RECT 1.999 6.804 2.001 9.24 ;
  LAYER M1 ;
        RECT 2.079 6.804 2.081 9.24 ;
  LAYER M1 ;
        RECT 2.159 6.804 2.161 9.24 ;
  LAYER M1 ;
        RECT 2.239 6.804 2.241 9.24 ;
  LAYER M1 ;
        RECT 2.319 6.804 2.321 9.24 ;
  LAYER M1 ;
        RECT 2.399 6.804 2.401 9.24 ;
  LAYER M1 ;
        RECT 2.479 6.804 2.481 9.24 ;
  LAYER M1 ;
        RECT 2.559 6.804 2.561 9.24 ;
  LAYER M1 ;
        RECT 2.639 6.804 2.641 9.24 ;
  LAYER M1 ;
        RECT 2.719 6.804 2.721 9.24 ;
  LAYER M1 ;
        RECT 2.799 6.804 2.801 9.24 ;
  LAYER M1 ;
        RECT 2.879 6.804 2.881 9.24 ;
  LAYER M1 ;
        RECT 2.959 6.804 2.961 9.24 ;
  LAYER M1 ;
        RECT 3.039 6.804 3.041 9.24 ;
  LAYER M2 ;
        RECT 0.72 6.803 3.12 6.805 ;
  LAYER M2 ;
        RECT 0.72 6.887 3.12 6.889 ;
  LAYER M2 ;
        RECT 0.72 6.971 3.12 6.973 ;
  LAYER M2 ;
        RECT 0.72 7.055 3.12 7.057 ;
  LAYER M2 ;
        RECT 0.72 7.139 3.12 7.141 ;
  LAYER M2 ;
        RECT 0.72 7.223 3.12 7.225 ;
  LAYER M2 ;
        RECT 0.72 7.307 3.12 7.309 ;
  LAYER M2 ;
        RECT 0.72 7.391 3.12 7.393 ;
  LAYER M2 ;
        RECT 0.72 7.475 3.12 7.477 ;
  LAYER M2 ;
        RECT 0.72 7.559 3.12 7.561 ;
  LAYER M2 ;
        RECT 0.72 7.643 3.12 7.645 ;
  LAYER M2 ;
        RECT 0.72 7.727 3.12 7.729 ;
  LAYER M2 ;
        RECT 0.72 7.8105 3.12 7.8125 ;
  LAYER M2 ;
        RECT 0.72 7.895 3.12 7.897 ;
  LAYER M2 ;
        RECT 0.72 7.979 3.12 7.981 ;
  LAYER M2 ;
        RECT 0.72 8.063 3.12 8.065 ;
  LAYER M2 ;
        RECT 0.72 8.147 3.12 8.149 ;
  LAYER M2 ;
        RECT 0.72 8.231 3.12 8.233 ;
  LAYER M2 ;
        RECT 0.72 8.315 3.12 8.317 ;
  LAYER M2 ;
        RECT 0.72 8.399 3.12 8.401 ;
  LAYER M2 ;
        RECT 0.72 8.483 3.12 8.485 ;
  LAYER M2 ;
        RECT 0.72 8.567 3.12 8.569 ;
  LAYER M2 ;
        RECT 0.72 8.651 3.12 8.653 ;
  LAYER M2 ;
        RECT 0.72 8.735 3.12 8.737 ;
  LAYER M2 ;
        RECT 0.72 8.819 3.12 8.821 ;
  LAYER M2 ;
        RECT 0.72 8.903 3.12 8.905 ;
  LAYER M2 ;
        RECT 0.72 8.987 3.12 8.989 ;
  LAYER M2 ;
        RECT 0.72 9.071 3.12 9.073 ;
  LAYER M2 ;
        RECT 0.72 9.155 3.12 9.157 ;
  LAYER M1 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M1 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M1 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M1 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M1 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M1 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M1 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M1 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M1 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M1 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M1 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M1 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M1 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M1 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M1 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M1 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M1 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M1 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M1 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M1 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M1 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M1 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M1 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M1 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M1 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M1 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M1 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M1 ;
        RECT 2.432 9.708 2.464 12.216 ;
  LAYER M1 ;
        RECT 2.496 9.708 2.528 12.216 ;
  LAYER M1 ;
        RECT 2.56 9.708 2.592 12.216 ;
  LAYER M1 ;
        RECT 2.624 9.708 2.656 12.216 ;
  LAYER M1 ;
        RECT 2.688 9.708 2.72 12.216 ;
  LAYER M1 ;
        RECT 2.752 9.708 2.784 12.216 ;
  LAYER M1 ;
        RECT 2.816 9.708 2.848 12.216 ;
  LAYER M1 ;
        RECT 2.88 9.708 2.912 12.216 ;
  LAYER M1 ;
        RECT 2.944 9.708 2.976 12.216 ;
  LAYER M1 ;
        RECT 3.008 9.708 3.04 12.216 ;
  LAYER M2 ;
        RECT 0.684 9.792 3.156 9.824 ;
  LAYER M2 ;
        RECT 0.684 9.856 3.156 9.888 ;
  LAYER M2 ;
        RECT 0.684 9.92 3.156 9.952 ;
  LAYER M2 ;
        RECT 0.684 9.984 3.156 10.016 ;
  LAYER M2 ;
        RECT 0.684 10.048 3.156 10.08 ;
  LAYER M2 ;
        RECT 0.684 10.112 3.156 10.144 ;
  LAYER M2 ;
        RECT 0.684 10.176 3.156 10.208 ;
  LAYER M2 ;
        RECT 0.684 10.24 3.156 10.272 ;
  LAYER M2 ;
        RECT 0.684 10.304 3.156 10.336 ;
  LAYER M2 ;
        RECT 0.684 10.368 3.156 10.4 ;
  LAYER M2 ;
        RECT 0.684 10.432 3.156 10.464 ;
  LAYER M2 ;
        RECT 0.684 10.496 3.156 10.528 ;
  LAYER M2 ;
        RECT 0.684 10.56 3.156 10.592 ;
  LAYER M2 ;
        RECT 0.684 10.624 3.156 10.656 ;
  LAYER M2 ;
        RECT 0.684 10.688 3.156 10.72 ;
  LAYER M2 ;
        RECT 0.684 10.752 3.156 10.784 ;
  LAYER M2 ;
        RECT 0.684 10.816 3.156 10.848 ;
  LAYER M2 ;
        RECT 0.684 10.88 3.156 10.912 ;
  LAYER M2 ;
        RECT 0.684 10.944 3.156 10.976 ;
  LAYER M2 ;
        RECT 0.684 11.008 3.156 11.04 ;
  LAYER M2 ;
        RECT 0.684 11.072 3.156 11.104 ;
  LAYER M2 ;
        RECT 0.684 11.136 3.156 11.168 ;
  LAYER M2 ;
        RECT 0.684 11.2 3.156 11.232 ;
  LAYER M2 ;
        RECT 0.684 11.264 3.156 11.296 ;
  LAYER M2 ;
        RECT 0.684 11.328 3.156 11.36 ;
  LAYER M2 ;
        RECT 0.684 11.392 3.156 11.424 ;
  LAYER M2 ;
        RECT 0.684 11.456 3.156 11.488 ;
  LAYER M2 ;
        RECT 0.684 11.52 3.156 11.552 ;
  LAYER M2 ;
        RECT 0.684 11.584 3.156 11.616 ;
  LAYER M2 ;
        RECT 0.684 11.648 3.156 11.68 ;
  LAYER M2 ;
        RECT 0.684 11.712 3.156 11.744 ;
  LAYER M2 ;
        RECT 0.684 11.776 3.156 11.808 ;
  LAYER M2 ;
        RECT 0.684 11.84 3.156 11.872 ;
  LAYER M2 ;
        RECT 0.684 11.904 3.156 11.936 ;
  LAYER M2 ;
        RECT 0.684 11.968 3.156 12 ;
  LAYER M2 ;
        RECT 0.684 12.032 3.156 12.064 ;
  LAYER M3 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M3 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M3 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M3 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M3 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M3 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M3 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M3 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M3 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M3 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M3 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M3 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M3 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M3 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M3 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M3 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M3 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M3 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M3 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M3 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M3 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M3 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M3 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M3 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M3 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M3 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M3 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M3 ;
        RECT 2.432 9.708 2.464 12.216 ;
  LAYER M3 ;
        RECT 2.496 9.708 2.528 12.216 ;
  LAYER M3 ;
        RECT 2.56 9.708 2.592 12.216 ;
  LAYER M3 ;
        RECT 2.624 9.708 2.656 12.216 ;
  LAYER M3 ;
        RECT 2.688 9.708 2.72 12.216 ;
  LAYER M3 ;
        RECT 2.752 9.708 2.784 12.216 ;
  LAYER M3 ;
        RECT 2.816 9.708 2.848 12.216 ;
  LAYER M3 ;
        RECT 2.88 9.708 2.912 12.216 ;
  LAYER M3 ;
        RECT 2.944 9.708 2.976 12.216 ;
  LAYER M3 ;
        RECT 3.008 9.708 3.04 12.216 ;
  LAYER M3 ;
        RECT 3.104 9.708 3.136 12.216 ;
  LAYER M1 ;
        RECT 0.719 9.744 0.721 12.18 ;
  LAYER M1 ;
        RECT 0.799 9.744 0.801 12.18 ;
  LAYER M1 ;
        RECT 0.879 9.744 0.881 12.18 ;
  LAYER M1 ;
        RECT 0.959 9.744 0.961 12.18 ;
  LAYER M1 ;
        RECT 1.039 9.744 1.041 12.18 ;
  LAYER M1 ;
        RECT 1.119 9.744 1.121 12.18 ;
  LAYER M1 ;
        RECT 1.199 9.744 1.201 12.18 ;
  LAYER M1 ;
        RECT 1.279 9.744 1.281 12.18 ;
  LAYER M1 ;
        RECT 1.359 9.744 1.361 12.18 ;
  LAYER M1 ;
        RECT 1.439 9.744 1.441 12.18 ;
  LAYER M1 ;
        RECT 1.519 9.744 1.521 12.18 ;
  LAYER M1 ;
        RECT 1.599 9.744 1.601 12.18 ;
  LAYER M1 ;
        RECT 1.679 9.744 1.681 12.18 ;
  LAYER M1 ;
        RECT 1.759 9.744 1.761 12.18 ;
  LAYER M1 ;
        RECT 1.839 9.744 1.841 12.18 ;
  LAYER M1 ;
        RECT 1.919 9.744 1.921 12.18 ;
  LAYER M1 ;
        RECT 1.999 9.744 2.001 12.18 ;
  LAYER M1 ;
        RECT 2.079 9.744 2.081 12.18 ;
  LAYER M1 ;
        RECT 2.159 9.744 2.161 12.18 ;
  LAYER M1 ;
        RECT 2.239 9.744 2.241 12.18 ;
  LAYER M1 ;
        RECT 2.319 9.744 2.321 12.18 ;
  LAYER M1 ;
        RECT 2.399 9.744 2.401 12.18 ;
  LAYER M1 ;
        RECT 2.479 9.744 2.481 12.18 ;
  LAYER M1 ;
        RECT 2.559 9.744 2.561 12.18 ;
  LAYER M1 ;
        RECT 2.639 9.744 2.641 12.18 ;
  LAYER M1 ;
        RECT 2.719 9.744 2.721 12.18 ;
  LAYER M1 ;
        RECT 2.799 9.744 2.801 12.18 ;
  LAYER M1 ;
        RECT 2.879 9.744 2.881 12.18 ;
  LAYER M1 ;
        RECT 2.959 9.744 2.961 12.18 ;
  LAYER M1 ;
        RECT 3.039 9.744 3.041 12.18 ;
  LAYER M2 ;
        RECT 0.72 9.743 3.12 9.745 ;
  LAYER M2 ;
        RECT 0.72 9.827 3.12 9.829 ;
  LAYER M2 ;
        RECT 0.72 9.911 3.12 9.913 ;
  LAYER M2 ;
        RECT 0.72 9.995 3.12 9.997 ;
  LAYER M2 ;
        RECT 0.72 10.079 3.12 10.081 ;
  LAYER M2 ;
        RECT 0.72 10.163 3.12 10.165 ;
  LAYER M2 ;
        RECT 0.72 10.247 3.12 10.249 ;
  LAYER M2 ;
        RECT 0.72 10.331 3.12 10.333 ;
  LAYER M2 ;
        RECT 0.72 10.415 3.12 10.417 ;
  LAYER M2 ;
        RECT 0.72 10.499 3.12 10.501 ;
  LAYER M2 ;
        RECT 0.72 10.583 3.12 10.585 ;
  LAYER M2 ;
        RECT 0.72 10.667 3.12 10.669 ;
  LAYER M2 ;
        RECT 0.72 10.7505 3.12 10.7525 ;
  LAYER M2 ;
        RECT 0.72 10.835 3.12 10.837 ;
  LAYER M2 ;
        RECT 0.72 10.919 3.12 10.921 ;
  LAYER M2 ;
        RECT 0.72 11.003 3.12 11.005 ;
  LAYER M2 ;
        RECT 0.72 11.087 3.12 11.089 ;
  LAYER M2 ;
        RECT 0.72 11.171 3.12 11.173 ;
  LAYER M2 ;
        RECT 0.72 11.255 3.12 11.257 ;
  LAYER M2 ;
        RECT 0.72 11.339 3.12 11.341 ;
  LAYER M2 ;
        RECT 0.72 11.423 3.12 11.425 ;
  LAYER M2 ;
        RECT 0.72 11.507 3.12 11.509 ;
  LAYER M2 ;
        RECT 0.72 11.591 3.12 11.593 ;
  LAYER M2 ;
        RECT 0.72 11.675 3.12 11.677 ;
  LAYER M2 ;
        RECT 0.72 11.759 3.12 11.761 ;
  LAYER M2 ;
        RECT 0.72 11.843 3.12 11.845 ;
  LAYER M2 ;
        RECT 0.72 11.927 3.12 11.929 ;
  LAYER M2 ;
        RECT 0.72 12.011 3.12 12.013 ;
  LAYER M2 ;
        RECT 0.72 12.095 3.12 12.097 ;
  LAYER M1 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M1 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M1 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M1 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M1 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M1 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M1 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M1 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M1 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M1 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M1 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M1 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M1 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M1 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M1 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M1 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M1 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M1 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M1 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M1 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M1 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M1 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M1 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M1 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M1 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M1 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M1 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M1 ;
        RECT 2.432 12.648 2.464 15.156 ;
  LAYER M1 ;
        RECT 2.496 12.648 2.528 15.156 ;
  LAYER M1 ;
        RECT 2.56 12.648 2.592 15.156 ;
  LAYER M1 ;
        RECT 2.624 12.648 2.656 15.156 ;
  LAYER M1 ;
        RECT 2.688 12.648 2.72 15.156 ;
  LAYER M1 ;
        RECT 2.752 12.648 2.784 15.156 ;
  LAYER M1 ;
        RECT 2.816 12.648 2.848 15.156 ;
  LAYER M1 ;
        RECT 2.88 12.648 2.912 15.156 ;
  LAYER M1 ;
        RECT 2.944 12.648 2.976 15.156 ;
  LAYER M1 ;
        RECT 3.008 12.648 3.04 15.156 ;
  LAYER M2 ;
        RECT 0.684 12.732 3.156 12.764 ;
  LAYER M2 ;
        RECT 0.684 12.796 3.156 12.828 ;
  LAYER M2 ;
        RECT 0.684 12.86 3.156 12.892 ;
  LAYER M2 ;
        RECT 0.684 12.924 3.156 12.956 ;
  LAYER M2 ;
        RECT 0.684 12.988 3.156 13.02 ;
  LAYER M2 ;
        RECT 0.684 13.052 3.156 13.084 ;
  LAYER M2 ;
        RECT 0.684 13.116 3.156 13.148 ;
  LAYER M2 ;
        RECT 0.684 13.18 3.156 13.212 ;
  LAYER M2 ;
        RECT 0.684 13.244 3.156 13.276 ;
  LAYER M2 ;
        RECT 0.684 13.308 3.156 13.34 ;
  LAYER M2 ;
        RECT 0.684 13.372 3.156 13.404 ;
  LAYER M2 ;
        RECT 0.684 13.436 3.156 13.468 ;
  LAYER M2 ;
        RECT 0.684 13.5 3.156 13.532 ;
  LAYER M2 ;
        RECT 0.684 13.564 3.156 13.596 ;
  LAYER M2 ;
        RECT 0.684 13.628 3.156 13.66 ;
  LAYER M2 ;
        RECT 0.684 13.692 3.156 13.724 ;
  LAYER M2 ;
        RECT 0.684 13.756 3.156 13.788 ;
  LAYER M2 ;
        RECT 0.684 13.82 3.156 13.852 ;
  LAYER M2 ;
        RECT 0.684 13.884 3.156 13.916 ;
  LAYER M2 ;
        RECT 0.684 13.948 3.156 13.98 ;
  LAYER M2 ;
        RECT 0.684 14.012 3.156 14.044 ;
  LAYER M2 ;
        RECT 0.684 14.076 3.156 14.108 ;
  LAYER M2 ;
        RECT 0.684 14.14 3.156 14.172 ;
  LAYER M2 ;
        RECT 0.684 14.204 3.156 14.236 ;
  LAYER M2 ;
        RECT 0.684 14.268 3.156 14.3 ;
  LAYER M2 ;
        RECT 0.684 14.332 3.156 14.364 ;
  LAYER M2 ;
        RECT 0.684 14.396 3.156 14.428 ;
  LAYER M2 ;
        RECT 0.684 14.46 3.156 14.492 ;
  LAYER M2 ;
        RECT 0.684 14.524 3.156 14.556 ;
  LAYER M2 ;
        RECT 0.684 14.588 3.156 14.62 ;
  LAYER M2 ;
        RECT 0.684 14.652 3.156 14.684 ;
  LAYER M2 ;
        RECT 0.684 14.716 3.156 14.748 ;
  LAYER M2 ;
        RECT 0.684 14.78 3.156 14.812 ;
  LAYER M2 ;
        RECT 0.684 14.844 3.156 14.876 ;
  LAYER M2 ;
        RECT 0.684 14.908 3.156 14.94 ;
  LAYER M2 ;
        RECT 0.684 14.972 3.156 15.004 ;
  LAYER M3 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M3 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M3 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M3 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M3 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M3 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M3 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M3 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M3 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M3 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M3 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M3 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M3 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M3 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M3 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M3 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M3 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M3 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M3 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M3 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M3 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M3 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M3 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M3 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M3 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M3 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M3 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M3 ;
        RECT 2.432 12.648 2.464 15.156 ;
  LAYER M3 ;
        RECT 2.496 12.648 2.528 15.156 ;
  LAYER M3 ;
        RECT 2.56 12.648 2.592 15.156 ;
  LAYER M3 ;
        RECT 2.624 12.648 2.656 15.156 ;
  LAYER M3 ;
        RECT 2.688 12.648 2.72 15.156 ;
  LAYER M3 ;
        RECT 2.752 12.648 2.784 15.156 ;
  LAYER M3 ;
        RECT 2.816 12.648 2.848 15.156 ;
  LAYER M3 ;
        RECT 2.88 12.648 2.912 15.156 ;
  LAYER M3 ;
        RECT 2.944 12.648 2.976 15.156 ;
  LAYER M3 ;
        RECT 3.008 12.648 3.04 15.156 ;
  LAYER M3 ;
        RECT 3.104 12.648 3.136 15.156 ;
  LAYER M1 ;
        RECT 0.719 12.684 0.721 15.12 ;
  LAYER M1 ;
        RECT 0.799 12.684 0.801 15.12 ;
  LAYER M1 ;
        RECT 0.879 12.684 0.881 15.12 ;
  LAYER M1 ;
        RECT 0.959 12.684 0.961 15.12 ;
  LAYER M1 ;
        RECT 1.039 12.684 1.041 15.12 ;
  LAYER M1 ;
        RECT 1.119 12.684 1.121 15.12 ;
  LAYER M1 ;
        RECT 1.199 12.684 1.201 15.12 ;
  LAYER M1 ;
        RECT 1.279 12.684 1.281 15.12 ;
  LAYER M1 ;
        RECT 1.359 12.684 1.361 15.12 ;
  LAYER M1 ;
        RECT 1.439 12.684 1.441 15.12 ;
  LAYER M1 ;
        RECT 1.519 12.684 1.521 15.12 ;
  LAYER M1 ;
        RECT 1.599 12.684 1.601 15.12 ;
  LAYER M1 ;
        RECT 1.679 12.684 1.681 15.12 ;
  LAYER M1 ;
        RECT 1.759 12.684 1.761 15.12 ;
  LAYER M1 ;
        RECT 1.839 12.684 1.841 15.12 ;
  LAYER M1 ;
        RECT 1.919 12.684 1.921 15.12 ;
  LAYER M1 ;
        RECT 1.999 12.684 2.001 15.12 ;
  LAYER M1 ;
        RECT 2.079 12.684 2.081 15.12 ;
  LAYER M1 ;
        RECT 2.159 12.684 2.161 15.12 ;
  LAYER M1 ;
        RECT 2.239 12.684 2.241 15.12 ;
  LAYER M1 ;
        RECT 2.319 12.684 2.321 15.12 ;
  LAYER M1 ;
        RECT 2.399 12.684 2.401 15.12 ;
  LAYER M1 ;
        RECT 2.479 12.684 2.481 15.12 ;
  LAYER M1 ;
        RECT 2.559 12.684 2.561 15.12 ;
  LAYER M1 ;
        RECT 2.639 12.684 2.641 15.12 ;
  LAYER M1 ;
        RECT 2.719 12.684 2.721 15.12 ;
  LAYER M1 ;
        RECT 2.799 12.684 2.801 15.12 ;
  LAYER M1 ;
        RECT 2.879 12.684 2.881 15.12 ;
  LAYER M1 ;
        RECT 2.959 12.684 2.961 15.12 ;
  LAYER M1 ;
        RECT 3.039 12.684 3.041 15.12 ;
  LAYER M2 ;
        RECT 0.72 12.683 3.12 12.685 ;
  LAYER M2 ;
        RECT 0.72 12.767 3.12 12.769 ;
  LAYER M2 ;
        RECT 0.72 12.851 3.12 12.853 ;
  LAYER M2 ;
        RECT 0.72 12.935 3.12 12.937 ;
  LAYER M2 ;
        RECT 0.72 13.019 3.12 13.021 ;
  LAYER M2 ;
        RECT 0.72 13.103 3.12 13.105 ;
  LAYER M2 ;
        RECT 0.72 13.187 3.12 13.189 ;
  LAYER M2 ;
        RECT 0.72 13.271 3.12 13.273 ;
  LAYER M2 ;
        RECT 0.72 13.355 3.12 13.357 ;
  LAYER M2 ;
        RECT 0.72 13.439 3.12 13.441 ;
  LAYER M2 ;
        RECT 0.72 13.523 3.12 13.525 ;
  LAYER M2 ;
        RECT 0.72 13.607 3.12 13.609 ;
  LAYER M2 ;
        RECT 0.72 13.6905 3.12 13.6925 ;
  LAYER M2 ;
        RECT 0.72 13.775 3.12 13.777 ;
  LAYER M2 ;
        RECT 0.72 13.859 3.12 13.861 ;
  LAYER M2 ;
        RECT 0.72 13.943 3.12 13.945 ;
  LAYER M2 ;
        RECT 0.72 14.027 3.12 14.029 ;
  LAYER M2 ;
        RECT 0.72 14.111 3.12 14.113 ;
  LAYER M2 ;
        RECT 0.72 14.195 3.12 14.197 ;
  LAYER M2 ;
        RECT 0.72 14.279 3.12 14.281 ;
  LAYER M2 ;
        RECT 0.72 14.363 3.12 14.365 ;
  LAYER M2 ;
        RECT 0.72 14.447 3.12 14.449 ;
  LAYER M2 ;
        RECT 0.72 14.531 3.12 14.533 ;
  LAYER M2 ;
        RECT 0.72 14.615 3.12 14.617 ;
  LAYER M2 ;
        RECT 0.72 14.699 3.12 14.701 ;
  LAYER M2 ;
        RECT 0.72 14.783 3.12 14.785 ;
  LAYER M2 ;
        RECT 0.72 14.867 3.12 14.869 ;
  LAYER M2 ;
        RECT 0.72 14.951 3.12 14.953 ;
  LAYER M2 ;
        RECT 0.72 15.035 3.12 15.037 ;
  LAYER M1 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M1 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M1 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M1 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M1 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M1 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M1 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M1 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M1 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M1 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M1 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M1 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M1 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M1 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M1 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M1 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M1 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M1 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M1 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M1 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M1 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M1 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M1 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M1 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M1 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M1 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M1 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M1 ;
        RECT 2.432 15.588 2.464 18.096 ;
  LAYER M1 ;
        RECT 2.496 15.588 2.528 18.096 ;
  LAYER M1 ;
        RECT 2.56 15.588 2.592 18.096 ;
  LAYER M1 ;
        RECT 2.624 15.588 2.656 18.096 ;
  LAYER M1 ;
        RECT 2.688 15.588 2.72 18.096 ;
  LAYER M1 ;
        RECT 2.752 15.588 2.784 18.096 ;
  LAYER M1 ;
        RECT 2.816 15.588 2.848 18.096 ;
  LAYER M1 ;
        RECT 2.88 15.588 2.912 18.096 ;
  LAYER M1 ;
        RECT 2.944 15.588 2.976 18.096 ;
  LAYER M1 ;
        RECT 3.008 15.588 3.04 18.096 ;
  LAYER M2 ;
        RECT 0.684 15.672 3.156 15.704 ;
  LAYER M2 ;
        RECT 0.684 15.736 3.156 15.768 ;
  LAYER M2 ;
        RECT 0.684 15.8 3.156 15.832 ;
  LAYER M2 ;
        RECT 0.684 15.864 3.156 15.896 ;
  LAYER M2 ;
        RECT 0.684 15.928 3.156 15.96 ;
  LAYER M2 ;
        RECT 0.684 15.992 3.156 16.024 ;
  LAYER M2 ;
        RECT 0.684 16.056 3.156 16.088 ;
  LAYER M2 ;
        RECT 0.684 16.12 3.156 16.152 ;
  LAYER M2 ;
        RECT 0.684 16.184 3.156 16.216 ;
  LAYER M2 ;
        RECT 0.684 16.248 3.156 16.28 ;
  LAYER M2 ;
        RECT 0.684 16.312 3.156 16.344 ;
  LAYER M2 ;
        RECT 0.684 16.376 3.156 16.408 ;
  LAYER M2 ;
        RECT 0.684 16.44 3.156 16.472 ;
  LAYER M2 ;
        RECT 0.684 16.504 3.156 16.536 ;
  LAYER M2 ;
        RECT 0.684 16.568 3.156 16.6 ;
  LAYER M2 ;
        RECT 0.684 16.632 3.156 16.664 ;
  LAYER M2 ;
        RECT 0.684 16.696 3.156 16.728 ;
  LAYER M2 ;
        RECT 0.684 16.76 3.156 16.792 ;
  LAYER M2 ;
        RECT 0.684 16.824 3.156 16.856 ;
  LAYER M2 ;
        RECT 0.684 16.888 3.156 16.92 ;
  LAYER M2 ;
        RECT 0.684 16.952 3.156 16.984 ;
  LAYER M2 ;
        RECT 0.684 17.016 3.156 17.048 ;
  LAYER M2 ;
        RECT 0.684 17.08 3.156 17.112 ;
  LAYER M2 ;
        RECT 0.684 17.144 3.156 17.176 ;
  LAYER M2 ;
        RECT 0.684 17.208 3.156 17.24 ;
  LAYER M2 ;
        RECT 0.684 17.272 3.156 17.304 ;
  LAYER M2 ;
        RECT 0.684 17.336 3.156 17.368 ;
  LAYER M2 ;
        RECT 0.684 17.4 3.156 17.432 ;
  LAYER M2 ;
        RECT 0.684 17.464 3.156 17.496 ;
  LAYER M2 ;
        RECT 0.684 17.528 3.156 17.56 ;
  LAYER M2 ;
        RECT 0.684 17.592 3.156 17.624 ;
  LAYER M2 ;
        RECT 0.684 17.656 3.156 17.688 ;
  LAYER M2 ;
        RECT 0.684 17.72 3.156 17.752 ;
  LAYER M2 ;
        RECT 0.684 17.784 3.156 17.816 ;
  LAYER M2 ;
        RECT 0.684 17.848 3.156 17.88 ;
  LAYER M2 ;
        RECT 0.684 17.912 3.156 17.944 ;
  LAYER M3 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M3 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M3 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M3 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M3 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M3 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M3 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M3 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M3 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M3 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M3 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M3 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M3 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M3 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M3 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M3 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M3 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M3 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M3 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M3 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M3 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M3 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M3 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M3 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M3 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M3 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M3 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M3 ;
        RECT 2.432 15.588 2.464 18.096 ;
  LAYER M3 ;
        RECT 2.496 15.588 2.528 18.096 ;
  LAYER M3 ;
        RECT 2.56 15.588 2.592 18.096 ;
  LAYER M3 ;
        RECT 2.624 15.588 2.656 18.096 ;
  LAYER M3 ;
        RECT 2.688 15.588 2.72 18.096 ;
  LAYER M3 ;
        RECT 2.752 15.588 2.784 18.096 ;
  LAYER M3 ;
        RECT 2.816 15.588 2.848 18.096 ;
  LAYER M3 ;
        RECT 2.88 15.588 2.912 18.096 ;
  LAYER M3 ;
        RECT 2.944 15.588 2.976 18.096 ;
  LAYER M3 ;
        RECT 3.008 15.588 3.04 18.096 ;
  LAYER M3 ;
        RECT 3.104 15.588 3.136 18.096 ;
  LAYER M1 ;
        RECT 0.719 15.624 0.721 18.06 ;
  LAYER M1 ;
        RECT 0.799 15.624 0.801 18.06 ;
  LAYER M1 ;
        RECT 0.879 15.624 0.881 18.06 ;
  LAYER M1 ;
        RECT 0.959 15.624 0.961 18.06 ;
  LAYER M1 ;
        RECT 1.039 15.624 1.041 18.06 ;
  LAYER M1 ;
        RECT 1.119 15.624 1.121 18.06 ;
  LAYER M1 ;
        RECT 1.199 15.624 1.201 18.06 ;
  LAYER M1 ;
        RECT 1.279 15.624 1.281 18.06 ;
  LAYER M1 ;
        RECT 1.359 15.624 1.361 18.06 ;
  LAYER M1 ;
        RECT 1.439 15.624 1.441 18.06 ;
  LAYER M1 ;
        RECT 1.519 15.624 1.521 18.06 ;
  LAYER M1 ;
        RECT 1.599 15.624 1.601 18.06 ;
  LAYER M1 ;
        RECT 1.679 15.624 1.681 18.06 ;
  LAYER M1 ;
        RECT 1.759 15.624 1.761 18.06 ;
  LAYER M1 ;
        RECT 1.839 15.624 1.841 18.06 ;
  LAYER M1 ;
        RECT 1.919 15.624 1.921 18.06 ;
  LAYER M1 ;
        RECT 1.999 15.624 2.001 18.06 ;
  LAYER M1 ;
        RECT 2.079 15.624 2.081 18.06 ;
  LAYER M1 ;
        RECT 2.159 15.624 2.161 18.06 ;
  LAYER M1 ;
        RECT 2.239 15.624 2.241 18.06 ;
  LAYER M1 ;
        RECT 2.319 15.624 2.321 18.06 ;
  LAYER M1 ;
        RECT 2.399 15.624 2.401 18.06 ;
  LAYER M1 ;
        RECT 2.479 15.624 2.481 18.06 ;
  LAYER M1 ;
        RECT 2.559 15.624 2.561 18.06 ;
  LAYER M1 ;
        RECT 2.639 15.624 2.641 18.06 ;
  LAYER M1 ;
        RECT 2.719 15.624 2.721 18.06 ;
  LAYER M1 ;
        RECT 2.799 15.624 2.801 18.06 ;
  LAYER M1 ;
        RECT 2.879 15.624 2.881 18.06 ;
  LAYER M1 ;
        RECT 2.959 15.624 2.961 18.06 ;
  LAYER M1 ;
        RECT 3.039 15.624 3.041 18.06 ;
  LAYER M2 ;
        RECT 0.72 15.623 3.12 15.625 ;
  LAYER M2 ;
        RECT 0.72 15.707 3.12 15.709 ;
  LAYER M2 ;
        RECT 0.72 15.791 3.12 15.793 ;
  LAYER M2 ;
        RECT 0.72 15.875 3.12 15.877 ;
  LAYER M2 ;
        RECT 0.72 15.959 3.12 15.961 ;
  LAYER M2 ;
        RECT 0.72 16.043 3.12 16.045 ;
  LAYER M2 ;
        RECT 0.72 16.127 3.12 16.129 ;
  LAYER M2 ;
        RECT 0.72 16.211 3.12 16.213 ;
  LAYER M2 ;
        RECT 0.72 16.295 3.12 16.297 ;
  LAYER M2 ;
        RECT 0.72 16.379 3.12 16.381 ;
  LAYER M2 ;
        RECT 0.72 16.463 3.12 16.465 ;
  LAYER M2 ;
        RECT 0.72 16.547 3.12 16.549 ;
  LAYER M2 ;
        RECT 0.72 16.6305 3.12 16.6325 ;
  LAYER M2 ;
        RECT 0.72 16.715 3.12 16.717 ;
  LAYER M2 ;
        RECT 0.72 16.799 3.12 16.801 ;
  LAYER M2 ;
        RECT 0.72 16.883 3.12 16.885 ;
  LAYER M2 ;
        RECT 0.72 16.967 3.12 16.969 ;
  LAYER M2 ;
        RECT 0.72 17.051 3.12 17.053 ;
  LAYER M2 ;
        RECT 0.72 17.135 3.12 17.137 ;
  LAYER M2 ;
        RECT 0.72 17.219 3.12 17.221 ;
  LAYER M2 ;
        RECT 0.72 17.303 3.12 17.305 ;
  LAYER M2 ;
        RECT 0.72 17.387 3.12 17.389 ;
  LAYER M2 ;
        RECT 0.72 17.471 3.12 17.473 ;
  LAYER M2 ;
        RECT 0.72 17.555 3.12 17.557 ;
  LAYER M2 ;
        RECT 0.72 17.639 3.12 17.641 ;
  LAYER M2 ;
        RECT 0.72 17.723 3.12 17.725 ;
  LAYER M2 ;
        RECT 0.72 17.807 3.12 17.809 ;
  LAYER M2 ;
        RECT 0.72 17.891 3.12 17.893 ;
  LAYER M2 ;
        RECT 0.72 17.975 3.12 17.977 ;
  LAYER M1 ;
        RECT 0.704 18.528 0.736 21.036 ;
  LAYER M1 ;
        RECT 0.768 18.528 0.8 21.036 ;
  LAYER M1 ;
        RECT 0.832 18.528 0.864 21.036 ;
  LAYER M1 ;
        RECT 0.896 18.528 0.928 21.036 ;
  LAYER M1 ;
        RECT 0.96 18.528 0.992 21.036 ;
  LAYER M1 ;
        RECT 1.024 18.528 1.056 21.036 ;
  LAYER M1 ;
        RECT 1.088 18.528 1.12 21.036 ;
  LAYER M1 ;
        RECT 1.152 18.528 1.184 21.036 ;
  LAYER M1 ;
        RECT 1.216 18.528 1.248 21.036 ;
  LAYER M1 ;
        RECT 1.28 18.528 1.312 21.036 ;
  LAYER M1 ;
        RECT 1.344 18.528 1.376 21.036 ;
  LAYER M1 ;
        RECT 1.408 18.528 1.44 21.036 ;
  LAYER M1 ;
        RECT 1.472 18.528 1.504 21.036 ;
  LAYER M1 ;
        RECT 1.536 18.528 1.568 21.036 ;
  LAYER M1 ;
        RECT 1.6 18.528 1.632 21.036 ;
  LAYER M1 ;
        RECT 1.664 18.528 1.696 21.036 ;
  LAYER M1 ;
        RECT 1.728 18.528 1.76 21.036 ;
  LAYER M1 ;
        RECT 1.792 18.528 1.824 21.036 ;
  LAYER M1 ;
        RECT 1.856 18.528 1.888 21.036 ;
  LAYER M1 ;
        RECT 1.92 18.528 1.952 21.036 ;
  LAYER M1 ;
        RECT 1.984 18.528 2.016 21.036 ;
  LAYER M1 ;
        RECT 2.048 18.528 2.08 21.036 ;
  LAYER M1 ;
        RECT 2.112 18.528 2.144 21.036 ;
  LAYER M1 ;
        RECT 2.176 18.528 2.208 21.036 ;
  LAYER M1 ;
        RECT 2.24 18.528 2.272 21.036 ;
  LAYER M1 ;
        RECT 2.304 18.528 2.336 21.036 ;
  LAYER M1 ;
        RECT 2.368 18.528 2.4 21.036 ;
  LAYER M1 ;
        RECT 2.432 18.528 2.464 21.036 ;
  LAYER M1 ;
        RECT 2.496 18.528 2.528 21.036 ;
  LAYER M1 ;
        RECT 2.56 18.528 2.592 21.036 ;
  LAYER M1 ;
        RECT 2.624 18.528 2.656 21.036 ;
  LAYER M1 ;
        RECT 2.688 18.528 2.72 21.036 ;
  LAYER M1 ;
        RECT 2.752 18.528 2.784 21.036 ;
  LAYER M1 ;
        RECT 2.816 18.528 2.848 21.036 ;
  LAYER M1 ;
        RECT 2.88 18.528 2.912 21.036 ;
  LAYER M1 ;
        RECT 2.944 18.528 2.976 21.036 ;
  LAYER M1 ;
        RECT 3.008 18.528 3.04 21.036 ;
  LAYER M2 ;
        RECT 0.684 18.612 3.156 18.644 ;
  LAYER M2 ;
        RECT 0.684 18.676 3.156 18.708 ;
  LAYER M2 ;
        RECT 0.684 18.74 3.156 18.772 ;
  LAYER M2 ;
        RECT 0.684 18.804 3.156 18.836 ;
  LAYER M2 ;
        RECT 0.684 18.868 3.156 18.9 ;
  LAYER M2 ;
        RECT 0.684 18.932 3.156 18.964 ;
  LAYER M2 ;
        RECT 0.684 18.996 3.156 19.028 ;
  LAYER M2 ;
        RECT 0.684 19.06 3.156 19.092 ;
  LAYER M2 ;
        RECT 0.684 19.124 3.156 19.156 ;
  LAYER M2 ;
        RECT 0.684 19.188 3.156 19.22 ;
  LAYER M2 ;
        RECT 0.684 19.252 3.156 19.284 ;
  LAYER M2 ;
        RECT 0.684 19.316 3.156 19.348 ;
  LAYER M2 ;
        RECT 0.684 19.38 3.156 19.412 ;
  LAYER M2 ;
        RECT 0.684 19.444 3.156 19.476 ;
  LAYER M2 ;
        RECT 0.684 19.508 3.156 19.54 ;
  LAYER M2 ;
        RECT 0.684 19.572 3.156 19.604 ;
  LAYER M2 ;
        RECT 0.684 19.636 3.156 19.668 ;
  LAYER M2 ;
        RECT 0.684 19.7 3.156 19.732 ;
  LAYER M2 ;
        RECT 0.684 19.764 3.156 19.796 ;
  LAYER M2 ;
        RECT 0.684 19.828 3.156 19.86 ;
  LAYER M2 ;
        RECT 0.684 19.892 3.156 19.924 ;
  LAYER M2 ;
        RECT 0.684 19.956 3.156 19.988 ;
  LAYER M2 ;
        RECT 0.684 20.02 3.156 20.052 ;
  LAYER M2 ;
        RECT 0.684 20.084 3.156 20.116 ;
  LAYER M2 ;
        RECT 0.684 20.148 3.156 20.18 ;
  LAYER M2 ;
        RECT 0.684 20.212 3.156 20.244 ;
  LAYER M2 ;
        RECT 0.684 20.276 3.156 20.308 ;
  LAYER M2 ;
        RECT 0.684 20.34 3.156 20.372 ;
  LAYER M2 ;
        RECT 0.684 20.404 3.156 20.436 ;
  LAYER M2 ;
        RECT 0.684 20.468 3.156 20.5 ;
  LAYER M2 ;
        RECT 0.684 20.532 3.156 20.564 ;
  LAYER M2 ;
        RECT 0.684 20.596 3.156 20.628 ;
  LAYER M2 ;
        RECT 0.684 20.66 3.156 20.692 ;
  LAYER M2 ;
        RECT 0.684 20.724 3.156 20.756 ;
  LAYER M2 ;
        RECT 0.684 20.788 3.156 20.82 ;
  LAYER M2 ;
        RECT 0.684 20.852 3.156 20.884 ;
  LAYER M3 ;
        RECT 0.704 18.528 0.736 21.036 ;
  LAYER M3 ;
        RECT 0.768 18.528 0.8 21.036 ;
  LAYER M3 ;
        RECT 0.832 18.528 0.864 21.036 ;
  LAYER M3 ;
        RECT 0.896 18.528 0.928 21.036 ;
  LAYER M3 ;
        RECT 0.96 18.528 0.992 21.036 ;
  LAYER M3 ;
        RECT 1.024 18.528 1.056 21.036 ;
  LAYER M3 ;
        RECT 1.088 18.528 1.12 21.036 ;
  LAYER M3 ;
        RECT 1.152 18.528 1.184 21.036 ;
  LAYER M3 ;
        RECT 1.216 18.528 1.248 21.036 ;
  LAYER M3 ;
        RECT 1.28 18.528 1.312 21.036 ;
  LAYER M3 ;
        RECT 1.344 18.528 1.376 21.036 ;
  LAYER M3 ;
        RECT 1.408 18.528 1.44 21.036 ;
  LAYER M3 ;
        RECT 1.472 18.528 1.504 21.036 ;
  LAYER M3 ;
        RECT 1.536 18.528 1.568 21.036 ;
  LAYER M3 ;
        RECT 1.6 18.528 1.632 21.036 ;
  LAYER M3 ;
        RECT 1.664 18.528 1.696 21.036 ;
  LAYER M3 ;
        RECT 1.728 18.528 1.76 21.036 ;
  LAYER M3 ;
        RECT 1.792 18.528 1.824 21.036 ;
  LAYER M3 ;
        RECT 1.856 18.528 1.888 21.036 ;
  LAYER M3 ;
        RECT 1.92 18.528 1.952 21.036 ;
  LAYER M3 ;
        RECT 1.984 18.528 2.016 21.036 ;
  LAYER M3 ;
        RECT 2.048 18.528 2.08 21.036 ;
  LAYER M3 ;
        RECT 2.112 18.528 2.144 21.036 ;
  LAYER M3 ;
        RECT 2.176 18.528 2.208 21.036 ;
  LAYER M3 ;
        RECT 2.24 18.528 2.272 21.036 ;
  LAYER M3 ;
        RECT 2.304 18.528 2.336 21.036 ;
  LAYER M3 ;
        RECT 2.368 18.528 2.4 21.036 ;
  LAYER M3 ;
        RECT 2.432 18.528 2.464 21.036 ;
  LAYER M3 ;
        RECT 2.496 18.528 2.528 21.036 ;
  LAYER M3 ;
        RECT 2.56 18.528 2.592 21.036 ;
  LAYER M3 ;
        RECT 2.624 18.528 2.656 21.036 ;
  LAYER M3 ;
        RECT 2.688 18.528 2.72 21.036 ;
  LAYER M3 ;
        RECT 2.752 18.528 2.784 21.036 ;
  LAYER M3 ;
        RECT 2.816 18.528 2.848 21.036 ;
  LAYER M3 ;
        RECT 2.88 18.528 2.912 21.036 ;
  LAYER M3 ;
        RECT 2.944 18.528 2.976 21.036 ;
  LAYER M3 ;
        RECT 3.008 18.528 3.04 21.036 ;
  LAYER M3 ;
        RECT 3.104 18.528 3.136 21.036 ;
  LAYER M1 ;
        RECT 0.719 18.564 0.721 21 ;
  LAYER M1 ;
        RECT 0.799 18.564 0.801 21 ;
  LAYER M1 ;
        RECT 0.879 18.564 0.881 21 ;
  LAYER M1 ;
        RECT 0.959 18.564 0.961 21 ;
  LAYER M1 ;
        RECT 1.039 18.564 1.041 21 ;
  LAYER M1 ;
        RECT 1.119 18.564 1.121 21 ;
  LAYER M1 ;
        RECT 1.199 18.564 1.201 21 ;
  LAYER M1 ;
        RECT 1.279 18.564 1.281 21 ;
  LAYER M1 ;
        RECT 1.359 18.564 1.361 21 ;
  LAYER M1 ;
        RECT 1.439 18.564 1.441 21 ;
  LAYER M1 ;
        RECT 1.519 18.564 1.521 21 ;
  LAYER M1 ;
        RECT 1.599 18.564 1.601 21 ;
  LAYER M1 ;
        RECT 1.679 18.564 1.681 21 ;
  LAYER M1 ;
        RECT 1.759 18.564 1.761 21 ;
  LAYER M1 ;
        RECT 1.839 18.564 1.841 21 ;
  LAYER M1 ;
        RECT 1.919 18.564 1.921 21 ;
  LAYER M1 ;
        RECT 1.999 18.564 2.001 21 ;
  LAYER M1 ;
        RECT 2.079 18.564 2.081 21 ;
  LAYER M1 ;
        RECT 2.159 18.564 2.161 21 ;
  LAYER M1 ;
        RECT 2.239 18.564 2.241 21 ;
  LAYER M1 ;
        RECT 2.319 18.564 2.321 21 ;
  LAYER M1 ;
        RECT 2.399 18.564 2.401 21 ;
  LAYER M1 ;
        RECT 2.479 18.564 2.481 21 ;
  LAYER M1 ;
        RECT 2.559 18.564 2.561 21 ;
  LAYER M1 ;
        RECT 2.639 18.564 2.641 21 ;
  LAYER M1 ;
        RECT 2.719 18.564 2.721 21 ;
  LAYER M1 ;
        RECT 2.799 18.564 2.801 21 ;
  LAYER M1 ;
        RECT 2.879 18.564 2.881 21 ;
  LAYER M1 ;
        RECT 2.959 18.564 2.961 21 ;
  LAYER M1 ;
        RECT 3.039 18.564 3.041 21 ;
  LAYER M2 ;
        RECT 0.72 18.563 3.12 18.565 ;
  LAYER M2 ;
        RECT 0.72 18.647 3.12 18.649 ;
  LAYER M2 ;
        RECT 0.72 18.731 3.12 18.733 ;
  LAYER M2 ;
        RECT 0.72 18.815 3.12 18.817 ;
  LAYER M2 ;
        RECT 0.72 18.899 3.12 18.901 ;
  LAYER M2 ;
        RECT 0.72 18.983 3.12 18.985 ;
  LAYER M2 ;
        RECT 0.72 19.067 3.12 19.069 ;
  LAYER M2 ;
        RECT 0.72 19.151 3.12 19.153 ;
  LAYER M2 ;
        RECT 0.72 19.235 3.12 19.237 ;
  LAYER M2 ;
        RECT 0.72 19.319 3.12 19.321 ;
  LAYER M2 ;
        RECT 0.72 19.403 3.12 19.405 ;
  LAYER M2 ;
        RECT 0.72 19.487 3.12 19.489 ;
  LAYER M2 ;
        RECT 0.72 19.5705 3.12 19.5725 ;
  LAYER M2 ;
        RECT 0.72 19.655 3.12 19.657 ;
  LAYER M2 ;
        RECT 0.72 19.739 3.12 19.741 ;
  LAYER M2 ;
        RECT 0.72 19.823 3.12 19.825 ;
  LAYER M2 ;
        RECT 0.72 19.907 3.12 19.909 ;
  LAYER M2 ;
        RECT 0.72 19.991 3.12 19.993 ;
  LAYER M2 ;
        RECT 0.72 20.075 3.12 20.077 ;
  LAYER M2 ;
        RECT 0.72 20.159 3.12 20.161 ;
  LAYER M2 ;
        RECT 0.72 20.243 3.12 20.245 ;
  LAYER M2 ;
        RECT 0.72 20.327 3.12 20.329 ;
  LAYER M2 ;
        RECT 0.72 20.411 3.12 20.413 ;
  LAYER M2 ;
        RECT 0.72 20.495 3.12 20.497 ;
  LAYER M2 ;
        RECT 0.72 20.579 3.12 20.581 ;
  LAYER M2 ;
        RECT 0.72 20.663 3.12 20.665 ;
  LAYER M2 ;
        RECT 0.72 20.747 3.12 20.749 ;
  LAYER M2 ;
        RECT 0.72 20.831 3.12 20.833 ;
  LAYER M2 ;
        RECT 0.72 20.915 3.12 20.917 ;
  LAYER M1 ;
        RECT 0.704 21.468 0.736 23.976 ;
  LAYER M1 ;
        RECT 0.768 21.468 0.8 23.976 ;
  LAYER M1 ;
        RECT 0.832 21.468 0.864 23.976 ;
  LAYER M1 ;
        RECT 0.896 21.468 0.928 23.976 ;
  LAYER M1 ;
        RECT 0.96 21.468 0.992 23.976 ;
  LAYER M1 ;
        RECT 1.024 21.468 1.056 23.976 ;
  LAYER M1 ;
        RECT 1.088 21.468 1.12 23.976 ;
  LAYER M1 ;
        RECT 1.152 21.468 1.184 23.976 ;
  LAYER M1 ;
        RECT 1.216 21.468 1.248 23.976 ;
  LAYER M1 ;
        RECT 1.28 21.468 1.312 23.976 ;
  LAYER M1 ;
        RECT 1.344 21.468 1.376 23.976 ;
  LAYER M1 ;
        RECT 1.408 21.468 1.44 23.976 ;
  LAYER M1 ;
        RECT 1.472 21.468 1.504 23.976 ;
  LAYER M1 ;
        RECT 1.536 21.468 1.568 23.976 ;
  LAYER M1 ;
        RECT 1.6 21.468 1.632 23.976 ;
  LAYER M1 ;
        RECT 1.664 21.468 1.696 23.976 ;
  LAYER M1 ;
        RECT 1.728 21.468 1.76 23.976 ;
  LAYER M1 ;
        RECT 1.792 21.468 1.824 23.976 ;
  LAYER M1 ;
        RECT 1.856 21.468 1.888 23.976 ;
  LAYER M1 ;
        RECT 1.92 21.468 1.952 23.976 ;
  LAYER M1 ;
        RECT 1.984 21.468 2.016 23.976 ;
  LAYER M1 ;
        RECT 2.048 21.468 2.08 23.976 ;
  LAYER M1 ;
        RECT 2.112 21.468 2.144 23.976 ;
  LAYER M1 ;
        RECT 2.176 21.468 2.208 23.976 ;
  LAYER M1 ;
        RECT 2.24 21.468 2.272 23.976 ;
  LAYER M1 ;
        RECT 2.304 21.468 2.336 23.976 ;
  LAYER M1 ;
        RECT 2.368 21.468 2.4 23.976 ;
  LAYER M1 ;
        RECT 2.432 21.468 2.464 23.976 ;
  LAYER M1 ;
        RECT 2.496 21.468 2.528 23.976 ;
  LAYER M1 ;
        RECT 2.56 21.468 2.592 23.976 ;
  LAYER M1 ;
        RECT 2.624 21.468 2.656 23.976 ;
  LAYER M1 ;
        RECT 2.688 21.468 2.72 23.976 ;
  LAYER M1 ;
        RECT 2.752 21.468 2.784 23.976 ;
  LAYER M1 ;
        RECT 2.816 21.468 2.848 23.976 ;
  LAYER M1 ;
        RECT 2.88 21.468 2.912 23.976 ;
  LAYER M1 ;
        RECT 2.944 21.468 2.976 23.976 ;
  LAYER M1 ;
        RECT 3.008 21.468 3.04 23.976 ;
  LAYER M2 ;
        RECT 0.684 21.552 3.156 21.584 ;
  LAYER M2 ;
        RECT 0.684 21.616 3.156 21.648 ;
  LAYER M2 ;
        RECT 0.684 21.68 3.156 21.712 ;
  LAYER M2 ;
        RECT 0.684 21.744 3.156 21.776 ;
  LAYER M2 ;
        RECT 0.684 21.808 3.156 21.84 ;
  LAYER M2 ;
        RECT 0.684 21.872 3.156 21.904 ;
  LAYER M2 ;
        RECT 0.684 21.936 3.156 21.968 ;
  LAYER M2 ;
        RECT 0.684 22 3.156 22.032 ;
  LAYER M2 ;
        RECT 0.684 22.064 3.156 22.096 ;
  LAYER M2 ;
        RECT 0.684 22.128 3.156 22.16 ;
  LAYER M2 ;
        RECT 0.684 22.192 3.156 22.224 ;
  LAYER M2 ;
        RECT 0.684 22.256 3.156 22.288 ;
  LAYER M2 ;
        RECT 0.684 22.32 3.156 22.352 ;
  LAYER M2 ;
        RECT 0.684 22.384 3.156 22.416 ;
  LAYER M2 ;
        RECT 0.684 22.448 3.156 22.48 ;
  LAYER M2 ;
        RECT 0.684 22.512 3.156 22.544 ;
  LAYER M2 ;
        RECT 0.684 22.576 3.156 22.608 ;
  LAYER M2 ;
        RECT 0.684 22.64 3.156 22.672 ;
  LAYER M2 ;
        RECT 0.684 22.704 3.156 22.736 ;
  LAYER M2 ;
        RECT 0.684 22.768 3.156 22.8 ;
  LAYER M2 ;
        RECT 0.684 22.832 3.156 22.864 ;
  LAYER M2 ;
        RECT 0.684 22.896 3.156 22.928 ;
  LAYER M2 ;
        RECT 0.684 22.96 3.156 22.992 ;
  LAYER M2 ;
        RECT 0.684 23.024 3.156 23.056 ;
  LAYER M2 ;
        RECT 0.684 23.088 3.156 23.12 ;
  LAYER M2 ;
        RECT 0.684 23.152 3.156 23.184 ;
  LAYER M2 ;
        RECT 0.684 23.216 3.156 23.248 ;
  LAYER M2 ;
        RECT 0.684 23.28 3.156 23.312 ;
  LAYER M2 ;
        RECT 0.684 23.344 3.156 23.376 ;
  LAYER M2 ;
        RECT 0.684 23.408 3.156 23.44 ;
  LAYER M2 ;
        RECT 0.684 23.472 3.156 23.504 ;
  LAYER M2 ;
        RECT 0.684 23.536 3.156 23.568 ;
  LAYER M2 ;
        RECT 0.684 23.6 3.156 23.632 ;
  LAYER M2 ;
        RECT 0.684 23.664 3.156 23.696 ;
  LAYER M2 ;
        RECT 0.684 23.728 3.156 23.76 ;
  LAYER M2 ;
        RECT 0.684 23.792 3.156 23.824 ;
  LAYER M3 ;
        RECT 0.704 21.468 0.736 23.976 ;
  LAYER M3 ;
        RECT 0.768 21.468 0.8 23.976 ;
  LAYER M3 ;
        RECT 0.832 21.468 0.864 23.976 ;
  LAYER M3 ;
        RECT 0.896 21.468 0.928 23.976 ;
  LAYER M3 ;
        RECT 0.96 21.468 0.992 23.976 ;
  LAYER M3 ;
        RECT 1.024 21.468 1.056 23.976 ;
  LAYER M3 ;
        RECT 1.088 21.468 1.12 23.976 ;
  LAYER M3 ;
        RECT 1.152 21.468 1.184 23.976 ;
  LAYER M3 ;
        RECT 1.216 21.468 1.248 23.976 ;
  LAYER M3 ;
        RECT 1.28 21.468 1.312 23.976 ;
  LAYER M3 ;
        RECT 1.344 21.468 1.376 23.976 ;
  LAYER M3 ;
        RECT 1.408 21.468 1.44 23.976 ;
  LAYER M3 ;
        RECT 1.472 21.468 1.504 23.976 ;
  LAYER M3 ;
        RECT 1.536 21.468 1.568 23.976 ;
  LAYER M3 ;
        RECT 1.6 21.468 1.632 23.976 ;
  LAYER M3 ;
        RECT 1.664 21.468 1.696 23.976 ;
  LAYER M3 ;
        RECT 1.728 21.468 1.76 23.976 ;
  LAYER M3 ;
        RECT 1.792 21.468 1.824 23.976 ;
  LAYER M3 ;
        RECT 1.856 21.468 1.888 23.976 ;
  LAYER M3 ;
        RECT 1.92 21.468 1.952 23.976 ;
  LAYER M3 ;
        RECT 1.984 21.468 2.016 23.976 ;
  LAYER M3 ;
        RECT 2.048 21.468 2.08 23.976 ;
  LAYER M3 ;
        RECT 2.112 21.468 2.144 23.976 ;
  LAYER M3 ;
        RECT 2.176 21.468 2.208 23.976 ;
  LAYER M3 ;
        RECT 2.24 21.468 2.272 23.976 ;
  LAYER M3 ;
        RECT 2.304 21.468 2.336 23.976 ;
  LAYER M3 ;
        RECT 2.368 21.468 2.4 23.976 ;
  LAYER M3 ;
        RECT 2.432 21.468 2.464 23.976 ;
  LAYER M3 ;
        RECT 2.496 21.468 2.528 23.976 ;
  LAYER M3 ;
        RECT 2.56 21.468 2.592 23.976 ;
  LAYER M3 ;
        RECT 2.624 21.468 2.656 23.976 ;
  LAYER M3 ;
        RECT 2.688 21.468 2.72 23.976 ;
  LAYER M3 ;
        RECT 2.752 21.468 2.784 23.976 ;
  LAYER M3 ;
        RECT 2.816 21.468 2.848 23.976 ;
  LAYER M3 ;
        RECT 2.88 21.468 2.912 23.976 ;
  LAYER M3 ;
        RECT 2.944 21.468 2.976 23.976 ;
  LAYER M3 ;
        RECT 3.008 21.468 3.04 23.976 ;
  LAYER M3 ;
        RECT 3.104 21.468 3.136 23.976 ;
  LAYER M1 ;
        RECT 0.719 21.504 0.721 23.94 ;
  LAYER M1 ;
        RECT 0.799 21.504 0.801 23.94 ;
  LAYER M1 ;
        RECT 0.879 21.504 0.881 23.94 ;
  LAYER M1 ;
        RECT 0.959 21.504 0.961 23.94 ;
  LAYER M1 ;
        RECT 1.039 21.504 1.041 23.94 ;
  LAYER M1 ;
        RECT 1.119 21.504 1.121 23.94 ;
  LAYER M1 ;
        RECT 1.199 21.504 1.201 23.94 ;
  LAYER M1 ;
        RECT 1.279 21.504 1.281 23.94 ;
  LAYER M1 ;
        RECT 1.359 21.504 1.361 23.94 ;
  LAYER M1 ;
        RECT 1.439 21.504 1.441 23.94 ;
  LAYER M1 ;
        RECT 1.519 21.504 1.521 23.94 ;
  LAYER M1 ;
        RECT 1.599 21.504 1.601 23.94 ;
  LAYER M1 ;
        RECT 1.679 21.504 1.681 23.94 ;
  LAYER M1 ;
        RECT 1.759 21.504 1.761 23.94 ;
  LAYER M1 ;
        RECT 1.839 21.504 1.841 23.94 ;
  LAYER M1 ;
        RECT 1.919 21.504 1.921 23.94 ;
  LAYER M1 ;
        RECT 1.999 21.504 2.001 23.94 ;
  LAYER M1 ;
        RECT 2.079 21.504 2.081 23.94 ;
  LAYER M1 ;
        RECT 2.159 21.504 2.161 23.94 ;
  LAYER M1 ;
        RECT 2.239 21.504 2.241 23.94 ;
  LAYER M1 ;
        RECT 2.319 21.504 2.321 23.94 ;
  LAYER M1 ;
        RECT 2.399 21.504 2.401 23.94 ;
  LAYER M1 ;
        RECT 2.479 21.504 2.481 23.94 ;
  LAYER M1 ;
        RECT 2.559 21.504 2.561 23.94 ;
  LAYER M1 ;
        RECT 2.639 21.504 2.641 23.94 ;
  LAYER M1 ;
        RECT 2.719 21.504 2.721 23.94 ;
  LAYER M1 ;
        RECT 2.799 21.504 2.801 23.94 ;
  LAYER M1 ;
        RECT 2.879 21.504 2.881 23.94 ;
  LAYER M1 ;
        RECT 2.959 21.504 2.961 23.94 ;
  LAYER M1 ;
        RECT 3.039 21.504 3.041 23.94 ;
  LAYER M2 ;
        RECT 0.72 21.503 3.12 21.505 ;
  LAYER M2 ;
        RECT 0.72 21.587 3.12 21.589 ;
  LAYER M2 ;
        RECT 0.72 21.671 3.12 21.673 ;
  LAYER M2 ;
        RECT 0.72 21.755 3.12 21.757 ;
  LAYER M2 ;
        RECT 0.72 21.839 3.12 21.841 ;
  LAYER M2 ;
        RECT 0.72 21.923 3.12 21.925 ;
  LAYER M2 ;
        RECT 0.72 22.007 3.12 22.009 ;
  LAYER M2 ;
        RECT 0.72 22.091 3.12 22.093 ;
  LAYER M2 ;
        RECT 0.72 22.175 3.12 22.177 ;
  LAYER M2 ;
        RECT 0.72 22.259 3.12 22.261 ;
  LAYER M2 ;
        RECT 0.72 22.343 3.12 22.345 ;
  LAYER M2 ;
        RECT 0.72 22.427 3.12 22.429 ;
  LAYER M2 ;
        RECT 0.72 22.5105 3.12 22.5125 ;
  LAYER M2 ;
        RECT 0.72 22.595 3.12 22.597 ;
  LAYER M2 ;
        RECT 0.72 22.679 3.12 22.681 ;
  LAYER M2 ;
        RECT 0.72 22.763 3.12 22.765 ;
  LAYER M2 ;
        RECT 0.72 22.847 3.12 22.849 ;
  LAYER M2 ;
        RECT 0.72 22.931 3.12 22.933 ;
  LAYER M2 ;
        RECT 0.72 23.015 3.12 23.017 ;
  LAYER M2 ;
        RECT 0.72 23.099 3.12 23.101 ;
  LAYER M2 ;
        RECT 0.72 23.183 3.12 23.185 ;
  LAYER M2 ;
        RECT 0.72 23.267 3.12 23.269 ;
  LAYER M2 ;
        RECT 0.72 23.351 3.12 23.353 ;
  LAYER M2 ;
        RECT 0.72 23.435 3.12 23.437 ;
  LAYER M2 ;
        RECT 0.72 23.519 3.12 23.521 ;
  LAYER M2 ;
        RECT 0.72 23.603 3.12 23.605 ;
  LAYER M2 ;
        RECT 0.72 23.687 3.12 23.689 ;
  LAYER M2 ;
        RECT 0.72 23.771 3.12 23.773 ;
  LAYER M2 ;
        RECT 0.72 23.855 3.12 23.857 ;
  LAYER M1 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M1 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M1 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M1 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M1 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M1 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M1 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M1 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M1 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M1 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M1 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M1 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M1 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M1 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M1 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M1 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M1 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M1 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M1 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M1 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M1 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M1 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M1 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M1 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M1 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M1 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M1 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M1 ;
        RECT 5.632 0.888 5.664 3.396 ;
  LAYER M1 ;
        RECT 5.696 0.888 5.728 3.396 ;
  LAYER M1 ;
        RECT 5.76 0.888 5.792 3.396 ;
  LAYER M1 ;
        RECT 5.824 0.888 5.856 3.396 ;
  LAYER M1 ;
        RECT 5.888 0.888 5.92 3.396 ;
  LAYER M1 ;
        RECT 5.952 0.888 5.984 3.396 ;
  LAYER M1 ;
        RECT 6.016 0.888 6.048 3.396 ;
  LAYER M1 ;
        RECT 6.08 0.888 6.112 3.396 ;
  LAYER M1 ;
        RECT 6.144 0.888 6.176 3.396 ;
  LAYER M1 ;
        RECT 6.208 0.888 6.24 3.396 ;
  LAYER M2 ;
        RECT 3.884 0.972 6.356 1.004 ;
  LAYER M2 ;
        RECT 3.884 1.036 6.356 1.068 ;
  LAYER M2 ;
        RECT 3.884 1.1 6.356 1.132 ;
  LAYER M2 ;
        RECT 3.884 1.164 6.356 1.196 ;
  LAYER M2 ;
        RECT 3.884 1.228 6.356 1.26 ;
  LAYER M2 ;
        RECT 3.884 1.292 6.356 1.324 ;
  LAYER M2 ;
        RECT 3.884 1.356 6.356 1.388 ;
  LAYER M2 ;
        RECT 3.884 1.42 6.356 1.452 ;
  LAYER M2 ;
        RECT 3.884 1.484 6.356 1.516 ;
  LAYER M2 ;
        RECT 3.884 1.548 6.356 1.58 ;
  LAYER M2 ;
        RECT 3.884 1.612 6.356 1.644 ;
  LAYER M2 ;
        RECT 3.884 1.676 6.356 1.708 ;
  LAYER M2 ;
        RECT 3.884 1.74 6.356 1.772 ;
  LAYER M2 ;
        RECT 3.884 1.804 6.356 1.836 ;
  LAYER M2 ;
        RECT 3.884 1.868 6.356 1.9 ;
  LAYER M2 ;
        RECT 3.884 1.932 6.356 1.964 ;
  LAYER M2 ;
        RECT 3.884 1.996 6.356 2.028 ;
  LAYER M2 ;
        RECT 3.884 2.06 6.356 2.092 ;
  LAYER M2 ;
        RECT 3.884 2.124 6.356 2.156 ;
  LAYER M2 ;
        RECT 3.884 2.188 6.356 2.22 ;
  LAYER M2 ;
        RECT 3.884 2.252 6.356 2.284 ;
  LAYER M2 ;
        RECT 3.884 2.316 6.356 2.348 ;
  LAYER M2 ;
        RECT 3.884 2.38 6.356 2.412 ;
  LAYER M2 ;
        RECT 3.884 2.444 6.356 2.476 ;
  LAYER M2 ;
        RECT 3.884 2.508 6.356 2.54 ;
  LAYER M2 ;
        RECT 3.884 2.572 6.356 2.604 ;
  LAYER M2 ;
        RECT 3.884 2.636 6.356 2.668 ;
  LAYER M2 ;
        RECT 3.884 2.7 6.356 2.732 ;
  LAYER M2 ;
        RECT 3.884 2.764 6.356 2.796 ;
  LAYER M2 ;
        RECT 3.884 2.828 6.356 2.86 ;
  LAYER M2 ;
        RECT 3.884 2.892 6.356 2.924 ;
  LAYER M2 ;
        RECT 3.884 2.956 6.356 2.988 ;
  LAYER M2 ;
        RECT 3.884 3.02 6.356 3.052 ;
  LAYER M2 ;
        RECT 3.884 3.084 6.356 3.116 ;
  LAYER M2 ;
        RECT 3.884 3.148 6.356 3.18 ;
  LAYER M2 ;
        RECT 3.884 3.212 6.356 3.244 ;
  LAYER M3 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M3 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M3 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M3 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M3 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M3 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M3 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M3 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M3 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M3 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M3 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M3 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M3 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M3 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M3 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M3 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M3 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M3 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M3 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M3 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M3 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M3 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M3 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M3 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M3 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M3 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M3 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M3 ;
        RECT 5.632 0.888 5.664 3.396 ;
  LAYER M3 ;
        RECT 5.696 0.888 5.728 3.396 ;
  LAYER M3 ;
        RECT 5.76 0.888 5.792 3.396 ;
  LAYER M3 ;
        RECT 5.824 0.888 5.856 3.396 ;
  LAYER M3 ;
        RECT 5.888 0.888 5.92 3.396 ;
  LAYER M3 ;
        RECT 5.952 0.888 5.984 3.396 ;
  LAYER M3 ;
        RECT 6.016 0.888 6.048 3.396 ;
  LAYER M3 ;
        RECT 6.08 0.888 6.112 3.396 ;
  LAYER M3 ;
        RECT 6.144 0.888 6.176 3.396 ;
  LAYER M3 ;
        RECT 6.208 0.888 6.24 3.396 ;
  LAYER M3 ;
        RECT 6.304 0.888 6.336 3.396 ;
  LAYER M1 ;
        RECT 3.919 0.924 3.921 3.36 ;
  LAYER M1 ;
        RECT 3.999 0.924 4.001 3.36 ;
  LAYER M1 ;
        RECT 4.079 0.924 4.081 3.36 ;
  LAYER M1 ;
        RECT 4.159 0.924 4.161 3.36 ;
  LAYER M1 ;
        RECT 4.239 0.924 4.241 3.36 ;
  LAYER M1 ;
        RECT 4.319 0.924 4.321 3.36 ;
  LAYER M1 ;
        RECT 4.399 0.924 4.401 3.36 ;
  LAYER M1 ;
        RECT 4.479 0.924 4.481 3.36 ;
  LAYER M1 ;
        RECT 4.559 0.924 4.561 3.36 ;
  LAYER M1 ;
        RECT 4.639 0.924 4.641 3.36 ;
  LAYER M1 ;
        RECT 4.719 0.924 4.721 3.36 ;
  LAYER M1 ;
        RECT 4.799 0.924 4.801 3.36 ;
  LAYER M1 ;
        RECT 4.879 0.924 4.881 3.36 ;
  LAYER M1 ;
        RECT 4.959 0.924 4.961 3.36 ;
  LAYER M1 ;
        RECT 5.039 0.924 5.041 3.36 ;
  LAYER M1 ;
        RECT 5.119 0.924 5.121 3.36 ;
  LAYER M1 ;
        RECT 5.199 0.924 5.201 3.36 ;
  LAYER M1 ;
        RECT 5.279 0.924 5.281 3.36 ;
  LAYER M1 ;
        RECT 5.359 0.924 5.361 3.36 ;
  LAYER M1 ;
        RECT 5.439 0.924 5.441 3.36 ;
  LAYER M1 ;
        RECT 5.519 0.924 5.521 3.36 ;
  LAYER M1 ;
        RECT 5.599 0.924 5.601 3.36 ;
  LAYER M1 ;
        RECT 5.679 0.924 5.681 3.36 ;
  LAYER M1 ;
        RECT 5.759 0.924 5.761 3.36 ;
  LAYER M1 ;
        RECT 5.839 0.924 5.841 3.36 ;
  LAYER M1 ;
        RECT 5.919 0.924 5.921 3.36 ;
  LAYER M1 ;
        RECT 5.999 0.924 6.001 3.36 ;
  LAYER M1 ;
        RECT 6.079 0.924 6.081 3.36 ;
  LAYER M1 ;
        RECT 6.159 0.924 6.161 3.36 ;
  LAYER M1 ;
        RECT 6.239 0.924 6.241 3.36 ;
  LAYER M2 ;
        RECT 3.92 0.923 6.32 0.925 ;
  LAYER M2 ;
        RECT 3.92 1.007 6.32 1.009 ;
  LAYER M2 ;
        RECT 3.92 1.091 6.32 1.093 ;
  LAYER M2 ;
        RECT 3.92 1.175 6.32 1.177 ;
  LAYER M2 ;
        RECT 3.92 1.259 6.32 1.261 ;
  LAYER M2 ;
        RECT 3.92 1.343 6.32 1.345 ;
  LAYER M2 ;
        RECT 3.92 1.427 6.32 1.429 ;
  LAYER M2 ;
        RECT 3.92 1.511 6.32 1.513 ;
  LAYER M2 ;
        RECT 3.92 1.595 6.32 1.597 ;
  LAYER M2 ;
        RECT 3.92 1.679 6.32 1.681 ;
  LAYER M2 ;
        RECT 3.92 1.763 6.32 1.765 ;
  LAYER M2 ;
        RECT 3.92 1.847 6.32 1.849 ;
  LAYER M2 ;
        RECT 3.92 1.9305 6.32 1.9325 ;
  LAYER M2 ;
        RECT 3.92 2.015 6.32 2.017 ;
  LAYER M2 ;
        RECT 3.92 2.099 6.32 2.101 ;
  LAYER M2 ;
        RECT 3.92 2.183 6.32 2.185 ;
  LAYER M2 ;
        RECT 3.92 2.267 6.32 2.269 ;
  LAYER M2 ;
        RECT 3.92 2.351 6.32 2.353 ;
  LAYER M2 ;
        RECT 3.92 2.435 6.32 2.437 ;
  LAYER M2 ;
        RECT 3.92 2.519 6.32 2.521 ;
  LAYER M2 ;
        RECT 3.92 2.603 6.32 2.605 ;
  LAYER M2 ;
        RECT 3.92 2.687 6.32 2.689 ;
  LAYER M2 ;
        RECT 3.92 2.771 6.32 2.773 ;
  LAYER M2 ;
        RECT 3.92 2.855 6.32 2.857 ;
  LAYER M2 ;
        RECT 3.92 2.939 6.32 2.941 ;
  LAYER M2 ;
        RECT 3.92 3.023 6.32 3.025 ;
  LAYER M2 ;
        RECT 3.92 3.107 6.32 3.109 ;
  LAYER M2 ;
        RECT 3.92 3.191 6.32 3.193 ;
  LAYER M2 ;
        RECT 3.92 3.275 6.32 3.277 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M1 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M1 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M1 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M1 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M1 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M1 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M1 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M1 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M1 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M1 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M1 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M1 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M1 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M1 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M1 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M1 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M1 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M1 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M1 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M1 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M1 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M1 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M1 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M1 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M1 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M1 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M1 ;
        RECT 5.632 3.828 5.664 6.336 ;
  LAYER M1 ;
        RECT 5.696 3.828 5.728 6.336 ;
  LAYER M1 ;
        RECT 5.76 3.828 5.792 6.336 ;
  LAYER M1 ;
        RECT 5.824 3.828 5.856 6.336 ;
  LAYER M1 ;
        RECT 5.888 3.828 5.92 6.336 ;
  LAYER M1 ;
        RECT 5.952 3.828 5.984 6.336 ;
  LAYER M1 ;
        RECT 6.016 3.828 6.048 6.336 ;
  LAYER M1 ;
        RECT 6.08 3.828 6.112 6.336 ;
  LAYER M1 ;
        RECT 6.144 3.828 6.176 6.336 ;
  LAYER M1 ;
        RECT 6.208 3.828 6.24 6.336 ;
  LAYER M2 ;
        RECT 3.884 3.912 6.356 3.944 ;
  LAYER M2 ;
        RECT 3.884 3.976 6.356 4.008 ;
  LAYER M2 ;
        RECT 3.884 4.04 6.356 4.072 ;
  LAYER M2 ;
        RECT 3.884 4.104 6.356 4.136 ;
  LAYER M2 ;
        RECT 3.884 4.168 6.356 4.2 ;
  LAYER M2 ;
        RECT 3.884 4.232 6.356 4.264 ;
  LAYER M2 ;
        RECT 3.884 4.296 6.356 4.328 ;
  LAYER M2 ;
        RECT 3.884 4.36 6.356 4.392 ;
  LAYER M2 ;
        RECT 3.884 4.424 6.356 4.456 ;
  LAYER M2 ;
        RECT 3.884 4.488 6.356 4.52 ;
  LAYER M2 ;
        RECT 3.884 4.552 6.356 4.584 ;
  LAYER M2 ;
        RECT 3.884 4.616 6.356 4.648 ;
  LAYER M2 ;
        RECT 3.884 4.68 6.356 4.712 ;
  LAYER M2 ;
        RECT 3.884 4.744 6.356 4.776 ;
  LAYER M2 ;
        RECT 3.884 4.808 6.356 4.84 ;
  LAYER M2 ;
        RECT 3.884 4.872 6.356 4.904 ;
  LAYER M2 ;
        RECT 3.884 4.936 6.356 4.968 ;
  LAYER M2 ;
        RECT 3.884 5 6.356 5.032 ;
  LAYER M2 ;
        RECT 3.884 5.064 6.356 5.096 ;
  LAYER M2 ;
        RECT 3.884 5.128 6.356 5.16 ;
  LAYER M2 ;
        RECT 3.884 5.192 6.356 5.224 ;
  LAYER M2 ;
        RECT 3.884 5.256 6.356 5.288 ;
  LAYER M2 ;
        RECT 3.884 5.32 6.356 5.352 ;
  LAYER M2 ;
        RECT 3.884 5.384 6.356 5.416 ;
  LAYER M2 ;
        RECT 3.884 5.448 6.356 5.48 ;
  LAYER M2 ;
        RECT 3.884 5.512 6.356 5.544 ;
  LAYER M2 ;
        RECT 3.884 5.576 6.356 5.608 ;
  LAYER M2 ;
        RECT 3.884 5.64 6.356 5.672 ;
  LAYER M2 ;
        RECT 3.884 5.704 6.356 5.736 ;
  LAYER M2 ;
        RECT 3.884 5.768 6.356 5.8 ;
  LAYER M2 ;
        RECT 3.884 5.832 6.356 5.864 ;
  LAYER M2 ;
        RECT 3.884 5.896 6.356 5.928 ;
  LAYER M2 ;
        RECT 3.884 5.96 6.356 5.992 ;
  LAYER M2 ;
        RECT 3.884 6.024 6.356 6.056 ;
  LAYER M2 ;
        RECT 3.884 6.088 6.356 6.12 ;
  LAYER M2 ;
        RECT 3.884 6.152 6.356 6.184 ;
  LAYER M3 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M3 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M3 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M3 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M3 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M3 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M3 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M3 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M3 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M3 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M3 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M3 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M3 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M3 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M3 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M3 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M3 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M3 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M3 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M3 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M3 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M3 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M3 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M3 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M3 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M3 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M3 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M3 ;
        RECT 5.632 3.828 5.664 6.336 ;
  LAYER M3 ;
        RECT 5.696 3.828 5.728 6.336 ;
  LAYER M3 ;
        RECT 5.76 3.828 5.792 6.336 ;
  LAYER M3 ;
        RECT 5.824 3.828 5.856 6.336 ;
  LAYER M3 ;
        RECT 5.888 3.828 5.92 6.336 ;
  LAYER M3 ;
        RECT 5.952 3.828 5.984 6.336 ;
  LAYER M3 ;
        RECT 6.016 3.828 6.048 6.336 ;
  LAYER M3 ;
        RECT 6.08 3.828 6.112 6.336 ;
  LAYER M3 ;
        RECT 6.144 3.828 6.176 6.336 ;
  LAYER M3 ;
        RECT 6.208 3.828 6.24 6.336 ;
  LAYER M3 ;
        RECT 6.304 3.828 6.336 6.336 ;
  LAYER M1 ;
        RECT 3.919 3.864 3.921 6.3 ;
  LAYER M1 ;
        RECT 3.999 3.864 4.001 6.3 ;
  LAYER M1 ;
        RECT 4.079 3.864 4.081 6.3 ;
  LAYER M1 ;
        RECT 4.159 3.864 4.161 6.3 ;
  LAYER M1 ;
        RECT 4.239 3.864 4.241 6.3 ;
  LAYER M1 ;
        RECT 4.319 3.864 4.321 6.3 ;
  LAYER M1 ;
        RECT 4.399 3.864 4.401 6.3 ;
  LAYER M1 ;
        RECT 4.479 3.864 4.481 6.3 ;
  LAYER M1 ;
        RECT 4.559 3.864 4.561 6.3 ;
  LAYER M1 ;
        RECT 4.639 3.864 4.641 6.3 ;
  LAYER M1 ;
        RECT 4.719 3.864 4.721 6.3 ;
  LAYER M1 ;
        RECT 4.799 3.864 4.801 6.3 ;
  LAYER M1 ;
        RECT 4.879 3.864 4.881 6.3 ;
  LAYER M1 ;
        RECT 4.959 3.864 4.961 6.3 ;
  LAYER M1 ;
        RECT 5.039 3.864 5.041 6.3 ;
  LAYER M1 ;
        RECT 5.119 3.864 5.121 6.3 ;
  LAYER M1 ;
        RECT 5.199 3.864 5.201 6.3 ;
  LAYER M1 ;
        RECT 5.279 3.864 5.281 6.3 ;
  LAYER M1 ;
        RECT 5.359 3.864 5.361 6.3 ;
  LAYER M1 ;
        RECT 5.439 3.864 5.441 6.3 ;
  LAYER M1 ;
        RECT 5.519 3.864 5.521 6.3 ;
  LAYER M1 ;
        RECT 5.599 3.864 5.601 6.3 ;
  LAYER M1 ;
        RECT 5.679 3.864 5.681 6.3 ;
  LAYER M1 ;
        RECT 5.759 3.864 5.761 6.3 ;
  LAYER M1 ;
        RECT 5.839 3.864 5.841 6.3 ;
  LAYER M1 ;
        RECT 5.919 3.864 5.921 6.3 ;
  LAYER M1 ;
        RECT 5.999 3.864 6.001 6.3 ;
  LAYER M1 ;
        RECT 6.079 3.864 6.081 6.3 ;
  LAYER M1 ;
        RECT 6.159 3.864 6.161 6.3 ;
  LAYER M1 ;
        RECT 6.239 3.864 6.241 6.3 ;
  LAYER M2 ;
        RECT 3.92 3.863 6.32 3.865 ;
  LAYER M2 ;
        RECT 3.92 3.947 6.32 3.949 ;
  LAYER M2 ;
        RECT 3.92 4.031 6.32 4.033 ;
  LAYER M2 ;
        RECT 3.92 4.115 6.32 4.117 ;
  LAYER M2 ;
        RECT 3.92 4.199 6.32 4.201 ;
  LAYER M2 ;
        RECT 3.92 4.283 6.32 4.285 ;
  LAYER M2 ;
        RECT 3.92 4.367 6.32 4.369 ;
  LAYER M2 ;
        RECT 3.92 4.451 6.32 4.453 ;
  LAYER M2 ;
        RECT 3.92 4.535 6.32 4.537 ;
  LAYER M2 ;
        RECT 3.92 4.619 6.32 4.621 ;
  LAYER M2 ;
        RECT 3.92 4.703 6.32 4.705 ;
  LAYER M2 ;
        RECT 3.92 4.787 6.32 4.789 ;
  LAYER M2 ;
        RECT 3.92 4.8705 6.32 4.8725 ;
  LAYER M2 ;
        RECT 3.92 4.955 6.32 4.957 ;
  LAYER M2 ;
        RECT 3.92 5.039 6.32 5.041 ;
  LAYER M2 ;
        RECT 3.92 5.123 6.32 5.125 ;
  LAYER M2 ;
        RECT 3.92 5.207 6.32 5.209 ;
  LAYER M2 ;
        RECT 3.92 5.291 6.32 5.293 ;
  LAYER M2 ;
        RECT 3.92 5.375 6.32 5.377 ;
  LAYER M2 ;
        RECT 3.92 5.459 6.32 5.461 ;
  LAYER M2 ;
        RECT 3.92 5.543 6.32 5.545 ;
  LAYER M2 ;
        RECT 3.92 5.627 6.32 5.629 ;
  LAYER M2 ;
        RECT 3.92 5.711 6.32 5.713 ;
  LAYER M2 ;
        RECT 3.92 5.795 6.32 5.797 ;
  LAYER M2 ;
        RECT 3.92 5.879 6.32 5.881 ;
  LAYER M2 ;
        RECT 3.92 5.963 6.32 5.965 ;
  LAYER M2 ;
        RECT 3.92 6.047 6.32 6.049 ;
  LAYER M2 ;
        RECT 3.92 6.131 6.32 6.133 ;
  LAYER M2 ;
        RECT 3.92 6.215 6.32 6.217 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M1 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M1 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M1 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M1 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M1 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M1 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M1 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M1 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M1 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M1 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M1 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M1 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M1 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M1 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M1 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M1 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M1 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M1 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M1 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M1 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M1 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M1 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M1 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M1 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M1 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M1 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M1 ;
        RECT 5.632 6.768 5.664 9.276 ;
  LAYER M1 ;
        RECT 5.696 6.768 5.728 9.276 ;
  LAYER M1 ;
        RECT 5.76 6.768 5.792 9.276 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 9.276 ;
  LAYER M1 ;
        RECT 5.888 6.768 5.92 9.276 ;
  LAYER M1 ;
        RECT 5.952 6.768 5.984 9.276 ;
  LAYER M1 ;
        RECT 6.016 6.768 6.048 9.276 ;
  LAYER M1 ;
        RECT 6.08 6.768 6.112 9.276 ;
  LAYER M1 ;
        RECT 6.144 6.768 6.176 9.276 ;
  LAYER M1 ;
        RECT 6.208 6.768 6.24 9.276 ;
  LAYER M2 ;
        RECT 3.884 6.852 6.356 6.884 ;
  LAYER M2 ;
        RECT 3.884 6.916 6.356 6.948 ;
  LAYER M2 ;
        RECT 3.884 6.98 6.356 7.012 ;
  LAYER M2 ;
        RECT 3.884 7.044 6.356 7.076 ;
  LAYER M2 ;
        RECT 3.884 7.108 6.356 7.14 ;
  LAYER M2 ;
        RECT 3.884 7.172 6.356 7.204 ;
  LAYER M2 ;
        RECT 3.884 7.236 6.356 7.268 ;
  LAYER M2 ;
        RECT 3.884 7.3 6.356 7.332 ;
  LAYER M2 ;
        RECT 3.884 7.364 6.356 7.396 ;
  LAYER M2 ;
        RECT 3.884 7.428 6.356 7.46 ;
  LAYER M2 ;
        RECT 3.884 7.492 6.356 7.524 ;
  LAYER M2 ;
        RECT 3.884 7.556 6.356 7.588 ;
  LAYER M2 ;
        RECT 3.884 7.62 6.356 7.652 ;
  LAYER M2 ;
        RECT 3.884 7.684 6.356 7.716 ;
  LAYER M2 ;
        RECT 3.884 7.748 6.356 7.78 ;
  LAYER M2 ;
        RECT 3.884 7.812 6.356 7.844 ;
  LAYER M2 ;
        RECT 3.884 7.876 6.356 7.908 ;
  LAYER M2 ;
        RECT 3.884 7.94 6.356 7.972 ;
  LAYER M2 ;
        RECT 3.884 8.004 6.356 8.036 ;
  LAYER M2 ;
        RECT 3.884 8.068 6.356 8.1 ;
  LAYER M2 ;
        RECT 3.884 8.132 6.356 8.164 ;
  LAYER M2 ;
        RECT 3.884 8.196 6.356 8.228 ;
  LAYER M2 ;
        RECT 3.884 8.26 6.356 8.292 ;
  LAYER M2 ;
        RECT 3.884 8.324 6.356 8.356 ;
  LAYER M2 ;
        RECT 3.884 8.388 6.356 8.42 ;
  LAYER M2 ;
        RECT 3.884 8.452 6.356 8.484 ;
  LAYER M2 ;
        RECT 3.884 8.516 6.356 8.548 ;
  LAYER M2 ;
        RECT 3.884 8.58 6.356 8.612 ;
  LAYER M2 ;
        RECT 3.884 8.644 6.356 8.676 ;
  LAYER M2 ;
        RECT 3.884 8.708 6.356 8.74 ;
  LAYER M2 ;
        RECT 3.884 8.772 6.356 8.804 ;
  LAYER M2 ;
        RECT 3.884 8.836 6.356 8.868 ;
  LAYER M2 ;
        RECT 3.884 8.9 6.356 8.932 ;
  LAYER M2 ;
        RECT 3.884 8.964 6.356 8.996 ;
  LAYER M2 ;
        RECT 3.884 9.028 6.356 9.06 ;
  LAYER M2 ;
        RECT 3.884 9.092 6.356 9.124 ;
  LAYER M3 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M3 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M3 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M3 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M3 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M3 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M3 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M3 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M3 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M3 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M3 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M3 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M3 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M3 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M3 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M3 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M3 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M3 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M3 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M3 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M3 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M3 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M3 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M3 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M3 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M3 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M3 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M3 ;
        RECT 5.632 6.768 5.664 9.276 ;
  LAYER M3 ;
        RECT 5.696 6.768 5.728 9.276 ;
  LAYER M3 ;
        RECT 5.76 6.768 5.792 9.276 ;
  LAYER M3 ;
        RECT 5.824 6.768 5.856 9.276 ;
  LAYER M3 ;
        RECT 5.888 6.768 5.92 9.276 ;
  LAYER M3 ;
        RECT 5.952 6.768 5.984 9.276 ;
  LAYER M3 ;
        RECT 6.016 6.768 6.048 9.276 ;
  LAYER M3 ;
        RECT 6.08 6.768 6.112 9.276 ;
  LAYER M3 ;
        RECT 6.144 6.768 6.176 9.276 ;
  LAYER M3 ;
        RECT 6.208 6.768 6.24 9.276 ;
  LAYER M3 ;
        RECT 6.304 6.768 6.336 9.276 ;
  LAYER M1 ;
        RECT 3.919 6.804 3.921 9.24 ;
  LAYER M1 ;
        RECT 3.999 6.804 4.001 9.24 ;
  LAYER M1 ;
        RECT 4.079 6.804 4.081 9.24 ;
  LAYER M1 ;
        RECT 4.159 6.804 4.161 9.24 ;
  LAYER M1 ;
        RECT 4.239 6.804 4.241 9.24 ;
  LAYER M1 ;
        RECT 4.319 6.804 4.321 9.24 ;
  LAYER M1 ;
        RECT 4.399 6.804 4.401 9.24 ;
  LAYER M1 ;
        RECT 4.479 6.804 4.481 9.24 ;
  LAYER M1 ;
        RECT 4.559 6.804 4.561 9.24 ;
  LAYER M1 ;
        RECT 4.639 6.804 4.641 9.24 ;
  LAYER M1 ;
        RECT 4.719 6.804 4.721 9.24 ;
  LAYER M1 ;
        RECT 4.799 6.804 4.801 9.24 ;
  LAYER M1 ;
        RECT 4.879 6.804 4.881 9.24 ;
  LAYER M1 ;
        RECT 4.959 6.804 4.961 9.24 ;
  LAYER M1 ;
        RECT 5.039 6.804 5.041 9.24 ;
  LAYER M1 ;
        RECT 5.119 6.804 5.121 9.24 ;
  LAYER M1 ;
        RECT 5.199 6.804 5.201 9.24 ;
  LAYER M1 ;
        RECT 5.279 6.804 5.281 9.24 ;
  LAYER M1 ;
        RECT 5.359 6.804 5.361 9.24 ;
  LAYER M1 ;
        RECT 5.439 6.804 5.441 9.24 ;
  LAYER M1 ;
        RECT 5.519 6.804 5.521 9.24 ;
  LAYER M1 ;
        RECT 5.599 6.804 5.601 9.24 ;
  LAYER M1 ;
        RECT 5.679 6.804 5.681 9.24 ;
  LAYER M1 ;
        RECT 5.759 6.804 5.761 9.24 ;
  LAYER M1 ;
        RECT 5.839 6.804 5.841 9.24 ;
  LAYER M1 ;
        RECT 5.919 6.804 5.921 9.24 ;
  LAYER M1 ;
        RECT 5.999 6.804 6.001 9.24 ;
  LAYER M1 ;
        RECT 6.079 6.804 6.081 9.24 ;
  LAYER M1 ;
        RECT 6.159 6.804 6.161 9.24 ;
  LAYER M1 ;
        RECT 6.239 6.804 6.241 9.24 ;
  LAYER M2 ;
        RECT 3.92 6.803 6.32 6.805 ;
  LAYER M2 ;
        RECT 3.92 6.887 6.32 6.889 ;
  LAYER M2 ;
        RECT 3.92 6.971 6.32 6.973 ;
  LAYER M2 ;
        RECT 3.92 7.055 6.32 7.057 ;
  LAYER M2 ;
        RECT 3.92 7.139 6.32 7.141 ;
  LAYER M2 ;
        RECT 3.92 7.223 6.32 7.225 ;
  LAYER M2 ;
        RECT 3.92 7.307 6.32 7.309 ;
  LAYER M2 ;
        RECT 3.92 7.391 6.32 7.393 ;
  LAYER M2 ;
        RECT 3.92 7.475 6.32 7.477 ;
  LAYER M2 ;
        RECT 3.92 7.559 6.32 7.561 ;
  LAYER M2 ;
        RECT 3.92 7.643 6.32 7.645 ;
  LAYER M2 ;
        RECT 3.92 7.727 6.32 7.729 ;
  LAYER M2 ;
        RECT 3.92 7.8105 6.32 7.8125 ;
  LAYER M2 ;
        RECT 3.92 7.895 6.32 7.897 ;
  LAYER M2 ;
        RECT 3.92 7.979 6.32 7.981 ;
  LAYER M2 ;
        RECT 3.92 8.063 6.32 8.065 ;
  LAYER M2 ;
        RECT 3.92 8.147 6.32 8.149 ;
  LAYER M2 ;
        RECT 3.92 8.231 6.32 8.233 ;
  LAYER M2 ;
        RECT 3.92 8.315 6.32 8.317 ;
  LAYER M2 ;
        RECT 3.92 8.399 6.32 8.401 ;
  LAYER M2 ;
        RECT 3.92 8.483 6.32 8.485 ;
  LAYER M2 ;
        RECT 3.92 8.567 6.32 8.569 ;
  LAYER M2 ;
        RECT 3.92 8.651 6.32 8.653 ;
  LAYER M2 ;
        RECT 3.92 8.735 6.32 8.737 ;
  LAYER M2 ;
        RECT 3.92 8.819 6.32 8.821 ;
  LAYER M2 ;
        RECT 3.92 8.903 6.32 8.905 ;
  LAYER M2 ;
        RECT 3.92 8.987 6.32 8.989 ;
  LAYER M2 ;
        RECT 3.92 9.071 6.32 9.073 ;
  LAYER M2 ;
        RECT 3.92 9.155 6.32 9.157 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M1 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M1 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M1 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M1 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M1 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M1 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M1 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M1 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M1 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M1 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M1 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M1 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M1 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M1 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M1 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M1 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M1 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M1 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M1 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M1 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M1 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M1 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M1 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M1 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M1 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M1 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M1 ;
        RECT 5.632 9.708 5.664 12.216 ;
  LAYER M1 ;
        RECT 5.696 9.708 5.728 12.216 ;
  LAYER M1 ;
        RECT 5.76 9.708 5.792 12.216 ;
  LAYER M1 ;
        RECT 5.824 9.708 5.856 12.216 ;
  LAYER M1 ;
        RECT 5.888 9.708 5.92 12.216 ;
  LAYER M1 ;
        RECT 5.952 9.708 5.984 12.216 ;
  LAYER M1 ;
        RECT 6.016 9.708 6.048 12.216 ;
  LAYER M1 ;
        RECT 6.08 9.708 6.112 12.216 ;
  LAYER M1 ;
        RECT 6.144 9.708 6.176 12.216 ;
  LAYER M1 ;
        RECT 6.208 9.708 6.24 12.216 ;
  LAYER M2 ;
        RECT 3.884 9.792 6.356 9.824 ;
  LAYER M2 ;
        RECT 3.884 9.856 6.356 9.888 ;
  LAYER M2 ;
        RECT 3.884 9.92 6.356 9.952 ;
  LAYER M2 ;
        RECT 3.884 9.984 6.356 10.016 ;
  LAYER M2 ;
        RECT 3.884 10.048 6.356 10.08 ;
  LAYER M2 ;
        RECT 3.884 10.112 6.356 10.144 ;
  LAYER M2 ;
        RECT 3.884 10.176 6.356 10.208 ;
  LAYER M2 ;
        RECT 3.884 10.24 6.356 10.272 ;
  LAYER M2 ;
        RECT 3.884 10.304 6.356 10.336 ;
  LAYER M2 ;
        RECT 3.884 10.368 6.356 10.4 ;
  LAYER M2 ;
        RECT 3.884 10.432 6.356 10.464 ;
  LAYER M2 ;
        RECT 3.884 10.496 6.356 10.528 ;
  LAYER M2 ;
        RECT 3.884 10.56 6.356 10.592 ;
  LAYER M2 ;
        RECT 3.884 10.624 6.356 10.656 ;
  LAYER M2 ;
        RECT 3.884 10.688 6.356 10.72 ;
  LAYER M2 ;
        RECT 3.884 10.752 6.356 10.784 ;
  LAYER M2 ;
        RECT 3.884 10.816 6.356 10.848 ;
  LAYER M2 ;
        RECT 3.884 10.88 6.356 10.912 ;
  LAYER M2 ;
        RECT 3.884 10.944 6.356 10.976 ;
  LAYER M2 ;
        RECT 3.884 11.008 6.356 11.04 ;
  LAYER M2 ;
        RECT 3.884 11.072 6.356 11.104 ;
  LAYER M2 ;
        RECT 3.884 11.136 6.356 11.168 ;
  LAYER M2 ;
        RECT 3.884 11.2 6.356 11.232 ;
  LAYER M2 ;
        RECT 3.884 11.264 6.356 11.296 ;
  LAYER M2 ;
        RECT 3.884 11.328 6.356 11.36 ;
  LAYER M2 ;
        RECT 3.884 11.392 6.356 11.424 ;
  LAYER M2 ;
        RECT 3.884 11.456 6.356 11.488 ;
  LAYER M2 ;
        RECT 3.884 11.52 6.356 11.552 ;
  LAYER M2 ;
        RECT 3.884 11.584 6.356 11.616 ;
  LAYER M2 ;
        RECT 3.884 11.648 6.356 11.68 ;
  LAYER M2 ;
        RECT 3.884 11.712 6.356 11.744 ;
  LAYER M2 ;
        RECT 3.884 11.776 6.356 11.808 ;
  LAYER M2 ;
        RECT 3.884 11.84 6.356 11.872 ;
  LAYER M2 ;
        RECT 3.884 11.904 6.356 11.936 ;
  LAYER M2 ;
        RECT 3.884 11.968 6.356 12 ;
  LAYER M2 ;
        RECT 3.884 12.032 6.356 12.064 ;
  LAYER M3 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M3 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M3 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M3 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M3 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M3 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M3 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M3 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M3 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M3 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M3 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M3 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M3 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M3 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M3 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M3 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M3 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M3 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M3 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M3 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M3 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M3 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M3 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M3 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M3 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M3 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M3 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M3 ;
        RECT 5.632 9.708 5.664 12.216 ;
  LAYER M3 ;
        RECT 5.696 9.708 5.728 12.216 ;
  LAYER M3 ;
        RECT 5.76 9.708 5.792 12.216 ;
  LAYER M3 ;
        RECT 5.824 9.708 5.856 12.216 ;
  LAYER M3 ;
        RECT 5.888 9.708 5.92 12.216 ;
  LAYER M3 ;
        RECT 5.952 9.708 5.984 12.216 ;
  LAYER M3 ;
        RECT 6.016 9.708 6.048 12.216 ;
  LAYER M3 ;
        RECT 6.08 9.708 6.112 12.216 ;
  LAYER M3 ;
        RECT 6.144 9.708 6.176 12.216 ;
  LAYER M3 ;
        RECT 6.208 9.708 6.24 12.216 ;
  LAYER M3 ;
        RECT 6.304 9.708 6.336 12.216 ;
  LAYER M1 ;
        RECT 3.919 9.744 3.921 12.18 ;
  LAYER M1 ;
        RECT 3.999 9.744 4.001 12.18 ;
  LAYER M1 ;
        RECT 4.079 9.744 4.081 12.18 ;
  LAYER M1 ;
        RECT 4.159 9.744 4.161 12.18 ;
  LAYER M1 ;
        RECT 4.239 9.744 4.241 12.18 ;
  LAYER M1 ;
        RECT 4.319 9.744 4.321 12.18 ;
  LAYER M1 ;
        RECT 4.399 9.744 4.401 12.18 ;
  LAYER M1 ;
        RECT 4.479 9.744 4.481 12.18 ;
  LAYER M1 ;
        RECT 4.559 9.744 4.561 12.18 ;
  LAYER M1 ;
        RECT 4.639 9.744 4.641 12.18 ;
  LAYER M1 ;
        RECT 4.719 9.744 4.721 12.18 ;
  LAYER M1 ;
        RECT 4.799 9.744 4.801 12.18 ;
  LAYER M1 ;
        RECT 4.879 9.744 4.881 12.18 ;
  LAYER M1 ;
        RECT 4.959 9.744 4.961 12.18 ;
  LAYER M1 ;
        RECT 5.039 9.744 5.041 12.18 ;
  LAYER M1 ;
        RECT 5.119 9.744 5.121 12.18 ;
  LAYER M1 ;
        RECT 5.199 9.744 5.201 12.18 ;
  LAYER M1 ;
        RECT 5.279 9.744 5.281 12.18 ;
  LAYER M1 ;
        RECT 5.359 9.744 5.361 12.18 ;
  LAYER M1 ;
        RECT 5.439 9.744 5.441 12.18 ;
  LAYER M1 ;
        RECT 5.519 9.744 5.521 12.18 ;
  LAYER M1 ;
        RECT 5.599 9.744 5.601 12.18 ;
  LAYER M1 ;
        RECT 5.679 9.744 5.681 12.18 ;
  LAYER M1 ;
        RECT 5.759 9.744 5.761 12.18 ;
  LAYER M1 ;
        RECT 5.839 9.744 5.841 12.18 ;
  LAYER M1 ;
        RECT 5.919 9.744 5.921 12.18 ;
  LAYER M1 ;
        RECT 5.999 9.744 6.001 12.18 ;
  LAYER M1 ;
        RECT 6.079 9.744 6.081 12.18 ;
  LAYER M1 ;
        RECT 6.159 9.744 6.161 12.18 ;
  LAYER M1 ;
        RECT 6.239 9.744 6.241 12.18 ;
  LAYER M2 ;
        RECT 3.92 9.743 6.32 9.745 ;
  LAYER M2 ;
        RECT 3.92 9.827 6.32 9.829 ;
  LAYER M2 ;
        RECT 3.92 9.911 6.32 9.913 ;
  LAYER M2 ;
        RECT 3.92 9.995 6.32 9.997 ;
  LAYER M2 ;
        RECT 3.92 10.079 6.32 10.081 ;
  LAYER M2 ;
        RECT 3.92 10.163 6.32 10.165 ;
  LAYER M2 ;
        RECT 3.92 10.247 6.32 10.249 ;
  LAYER M2 ;
        RECT 3.92 10.331 6.32 10.333 ;
  LAYER M2 ;
        RECT 3.92 10.415 6.32 10.417 ;
  LAYER M2 ;
        RECT 3.92 10.499 6.32 10.501 ;
  LAYER M2 ;
        RECT 3.92 10.583 6.32 10.585 ;
  LAYER M2 ;
        RECT 3.92 10.667 6.32 10.669 ;
  LAYER M2 ;
        RECT 3.92 10.7505 6.32 10.7525 ;
  LAYER M2 ;
        RECT 3.92 10.835 6.32 10.837 ;
  LAYER M2 ;
        RECT 3.92 10.919 6.32 10.921 ;
  LAYER M2 ;
        RECT 3.92 11.003 6.32 11.005 ;
  LAYER M2 ;
        RECT 3.92 11.087 6.32 11.089 ;
  LAYER M2 ;
        RECT 3.92 11.171 6.32 11.173 ;
  LAYER M2 ;
        RECT 3.92 11.255 6.32 11.257 ;
  LAYER M2 ;
        RECT 3.92 11.339 6.32 11.341 ;
  LAYER M2 ;
        RECT 3.92 11.423 6.32 11.425 ;
  LAYER M2 ;
        RECT 3.92 11.507 6.32 11.509 ;
  LAYER M2 ;
        RECT 3.92 11.591 6.32 11.593 ;
  LAYER M2 ;
        RECT 3.92 11.675 6.32 11.677 ;
  LAYER M2 ;
        RECT 3.92 11.759 6.32 11.761 ;
  LAYER M2 ;
        RECT 3.92 11.843 6.32 11.845 ;
  LAYER M2 ;
        RECT 3.92 11.927 6.32 11.929 ;
  LAYER M2 ;
        RECT 3.92 12.011 6.32 12.013 ;
  LAYER M2 ;
        RECT 3.92 12.095 6.32 12.097 ;
  LAYER M1 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M1 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M1 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M1 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M1 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M1 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M1 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M1 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M1 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M1 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M1 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M1 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M1 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M1 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M1 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M1 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M1 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M1 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M1 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M1 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M1 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M1 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M1 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M1 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M1 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M1 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M1 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M1 ;
        RECT 5.632 12.648 5.664 15.156 ;
  LAYER M1 ;
        RECT 5.696 12.648 5.728 15.156 ;
  LAYER M1 ;
        RECT 5.76 12.648 5.792 15.156 ;
  LAYER M1 ;
        RECT 5.824 12.648 5.856 15.156 ;
  LAYER M1 ;
        RECT 5.888 12.648 5.92 15.156 ;
  LAYER M1 ;
        RECT 5.952 12.648 5.984 15.156 ;
  LAYER M1 ;
        RECT 6.016 12.648 6.048 15.156 ;
  LAYER M1 ;
        RECT 6.08 12.648 6.112 15.156 ;
  LAYER M1 ;
        RECT 6.144 12.648 6.176 15.156 ;
  LAYER M1 ;
        RECT 6.208 12.648 6.24 15.156 ;
  LAYER M2 ;
        RECT 3.884 12.732 6.356 12.764 ;
  LAYER M2 ;
        RECT 3.884 12.796 6.356 12.828 ;
  LAYER M2 ;
        RECT 3.884 12.86 6.356 12.892 ;
  LAYER M2 ;
        RECT 3.884 12.924 6.356 12.956 ;
  LAYER M2 ;
        RECT 3.884 12.988 6.356 13.02 ;
  LAYER M2 ;
        RECT 3.884 13.052 6.356 13.084 ;
  LAYER M2 ;
        RECT 3.884 13.116 6.356 13.148 ;
  LAYER M2 ;
        RECT 3.884 13.18 6.356 13.212 ;
  LAYER M2 ;
        RECT 3.884 13.244 6.356 13.276 ;
  LAYER M2 ;
        RECT 3.884 13.308 6.356 13.34 ;
  LAYER M2 ;
        RECT 3.884 13.372 6.356 13.404 ;
  LAYER M2 ;
        RECT 3.884 13.436 6.356 13.468 ;
  LAYER M2 ;
        RECT 3.884 13.5 6.356 13.532 ;
  LAYER M2 ;
        RECT 3.884 13.564 6.356 13.596 ;
  LAYER M2 ;
        RECT 3.884 13.628 6.356 13.66 ;
  LAYER M2 ;
        RECT 3.884 13.692 6.356 13.724 ;
  LAYER M2 ;
        RECT 3.884 13.756 6.356 13.788 ;
  LAYER M2 ;
        RECT 3.884 13.82 6.356 13.852 ;
  LAYER M2 ;
        RECT 3.884 13.884 6.356 13.916 ;
  LAYER M2 ;
        RECT 3.884 13.948 6.356 13.98 ;
  LAYER M2 ;
        RECT 3.884 14.012 6.356 14.044 ;
  LAYER M2 ;
        RECT 3.884 14.076 6.356 14.108 ;
  LAYER M2 ;
        RECT 3.884 14.14 6.356 14.172 ;
  LAYER M2 ;
        RECT 3.884 14.204 6.356 14.236 ;
  LAYER M2 ;
        RECT 3.884 14.268 6.356 14.3 ;
  LAYER M2 ;
        RECT 3.884 14.332 6.356 14.364 ;
  LAYER M2 ;
        RECT 3.884 14.396 6.356 14.428 ;
  LAYER M2 ;
        RECT 3.884 14.46 6.356 14.492 ;
  LAYER M2 ;
        RECT 3.884 14.524 6.356 14.556 ;
  LAYER M2 ;
        RECT 3.884 14.588 6.356 14.62 ;
  LAYER M2 ;
        RECT 3.884 14.652 6.356 14.684 ;
  LAYER M2 ;
        RECT 3.884 14.716 6.356 14.748 ;
  LAYER M2 ;
        RECT 3.884 14.78 6.356 14.812 ;
  LAYER M2 ;
        RECT 3.884 14.844 6.356 14.876 ;
  LAYER M2 ;
        RECT 3.884 14.908 6.356 14.94 ;
  LAYER M2 ;
        RECT 3.884 14.972 6.356 15.004 ;
  LAYER M3 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M3 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M3 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M3 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M3 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M3 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M3 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M3 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M3 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M3 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M3 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M3 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M3 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M3 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M3 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M3 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M3 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M3 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M3 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M3 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M3 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M3 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M3 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M3 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M3 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M3 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M3 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M3 ;
        RECT 5.632 12.648 5.664 15.156 ;
  LAYER M3 ;
        RECT 5.696 12.648 5.728 15.156 ;
  LAYER M3 ;
        RECT 5.76 12.648 5.792 15.156 ;
  LAYER M3 ;
        RECT 5.824 12.648 5.856 15.156 ;
  LAYER M3 ;
        RECT 5.888 12.648 5.92 15.156 ;
  LAYER M3 ;
        RECT 5.952 12.648 5.984 15.156 ;
  LAYER M3 ;
        RECT 6.016 12.648 6.048 15.156 ;
  LAYER M3 ;
        RECT 6.08 12.648 6.112 15.156 ;
  LAYER M3 ;
        RECT 6.144 12.648 6.176 15.156 ;
  LAYER M3 ;
        RECT 6.208 12.648 6.24 15.156 ;
  LAYER M3 ;
        RECT 6.304 12.648 6.336 15.156 ;
  LAYER M1 ;
        RECT 3.919 12.684 3.921 15.12 ;
  LAYER M1 ;
        RECT 3.999 12.684 4.001 15.12 ;
  LAYER M1 ;
        RECT 4.079 12.684 4.081 15.12 ;
  LAYER M1 ;
        RECT 4.159 12.684 4.161 15.12 ;
  LAYER M1 ;
        RECT 4.239 12.684 4.241 15.12 ;
  LAYER M1 ;
        RECT 4.319 12.684 4.321 15.12 ;
  LAYER M1 ;
        RECT 4.399 12.684 4.401 15.12 ;
  LAYER M1 ;
        RECT 4.479 12.684 4.481 15.12 ;
  LAYER M1 ;
        RECT 4.559 12.684 4.561 15.12 ;
  LAYER M1 ;
        RECT 4.639 12.684 4.641 15.12 ;
  LAYER M1 ;
        RECT 4.719 12.684 4.721 15.12 ;
  LAYER M1 ;
        RECT 4.799 12.684 4.801 15.12 ;
  LAYER M1 ;
        RECT 4.879 12.684 4.881 15.12 ;
  LAYER M1 ;
        RECT 4.959 12.684 4.961 15.12 ;
  LAYER M1 ;
        RECT 5.039 12.684 5.041 15.12 ;
  LAYER M1 ;
        RECT 5.119 12.684 5.121 15.12 ;
  LAYER M1 ;
        RECT 5.199 12.684 5.201 15.12 ;
  LAYER M1 ;
        RECT 5.279 12.684 5.281 15.12 ;
  LAYER M1 ;
        RECT 5.359 12.684 5.361 15.12 ;
  LAYER M1 ;
        RECT 5.439 12.684 5.441 15.12 ;
  LAYER M1 ;
        RECT 5.519 12.684 5.521 15.12 ;
  LAYER M1 ;
        RECT 5.599 12.684 5.601 15.12 ;
  LAYER M1 ;
        RECT 5.679 12.684 5.681 15.12 ;
  LAYER M1 ;
        RECT 5.759 12.684 5.761 15.12 ;
  LAYER M1 ;
        RECT 5.839 12.684 5.841 15.12 ;
  LAYER M1 ;
        RECT 5.919 12.684 5.921 15.12 ;
  LAYER M1 ;
        RECT 5.999 12.684 6.001 15.12 ;
  LAYER M1 ;
        RECT 6.079 12.684 6.081 15.12 ;
  LAYER M1 ;
        RECT 6.159 12.684 6.161 15.12 ;
  LAYER M1 ;
        RECT 6.239 12.684 6.241 15.12 ;
  LAYER M2 ;
        RECT 3.92 12.683 6.32 12.685 ;
  LAYER M2 ;
        RECT 3.92 12.767 6.32 12.769 ;
  LAYER M2 ;
        RECT 3.92 12.851 6.32 12.853 ;
  LAYER M2 ;
        RECT 3.92 12.935 6.32 12.937 ;
  LAYER M2 ;
        RECT 3.92 13.019 6.32 13.021 ;
  LAYER M2 ;
        RECT 3.92 13.103 6.32 13.105 ;
  LAYER M2 ;
        RECT 3.92 13.187 6.32 13.189 ;
  LAYER M2 ;
        RECT 3.92 13.271 6.32 13.273 ;
  LAYER M2 ;
        RECT 3.92 13.355 6.32 13.357 ;
  LAYER M2 ;
        RECT 3.92 13.439 6.32 13.441 ;
  LAYER M2 ;
        RECT 3.92 13.523 6.32 13.525 ;
  LAYER M2 ;
        RECT 3.92 13.607 6.32 13.609 ;
  LAYER M2 ;
        RECT 3.92 13.6905 6.32 13.6925 ;
  LAYER M2 ;
        RECT 3.92 13.775 6.32 13.777 ;
  LAYER M2 ;
        RECT 3.92 13.859 6.32 13.861 ;
  LAYER M2 ;
        RECT 3.92 13.943 6.32 13.945 ;
  LAYER M2 ;
        RECT 3.92 14.027 6.32 14.029 ;
  LAYER M2 ;
        RECT 3.92 14.111 6.32 14.113 ;
  LAYER M2 ;
        RECT 3.92 14.195 6.32 14.197 ;
  LAYER M2 ;
        RECT 3.92 14.279 6.32 14.281 ;
  LAYER M2 ;
        RECT 3.92 14.363 6.32 14.365 ;
  LAYER M2 ;
        RECT 3.92 14.447 6.32 14.449 ;
  LAYER M2 ;
        RECT 3.92 14.531 6.32 14.533 ;
  LAYER M2 ;
        RECT 3.92 14.615 6.32 14.617 ;
  LAYER M2 ;
        RECT 3.92 14.699 6.32 14.701 ;
  LAYER M2 ;
        RECT 3.92 14.783 6.32 14.785 ;
  LAYER M2 ;
        RECT 3.92 14.867 6.32 14.869 ;
  LAYER M2 ;
        RECT 3.92 14.951 6.32 14.953 ;
  LAYER M2 ;
        RECT 3.92 15.035 6.32 15.037 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M1 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M1 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M1 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M1 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M1 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M1 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M1 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M1 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M1 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M1 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M1 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M1 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M1 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M1 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M1 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M1 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M1 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M1 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M1 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M1 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M1 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M1 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M1 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M1 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M1 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M1 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M1 ;
        RECT 5.632 15.588 5.664 18.096 ;
  LAYER M1 ;
        RECT 5.696 15.588 5.728 18.096 ;
  LAYER M1 ;
        RECT 5.76 15.588 5.792 18.096 ;
  LAYER M1 ;
        RECT 5.824 15.588 5.856 18.096 ;
  LAYER M1 ;
        RECT 5.888 15.588 5.92 18.096 ;
  LAYER M1 ;
        RECT 5.952 15.588 5.984 18.096 ;
  LAYER M1 ;
        RECT 6.016 15.588 6.048 18.096 ;
  LAYER M1 ;
        RECT 6.08 15.588 6.112 18.096 ;
  LAYER M1 ;
        RECT 6.144 15.588 6.176 18.096 ;
  LAYER M1 ;
        RECT 6.208 15.588 6.24 18.096 ;
  LAYER M2 ;
        RECT 3.884 15.672 6.356 15.704 ;
  LAYER M2 ;
        RECT 3.884 15.736 6.356 15.768 ;
  LAYER M2 ;
        RECT 3.884 15.8 6.356 15.832 ;
  LAYER M2 ;
        RECT 3.884 15.864 6.356 15.896 ;
  LAYER M2 ;
        RECT 3.884 15.928 6.356 15.96 ;
  LAYER M2 ;
        RECT 3.884 15.992 6.356 16.024 ;
  LAYER M2 ;
        RECT 3.884 16.056 6.356 16.088 ;
  LAYER M2 ;
        RECT 3.884 16.12 6.356 16.152 ;
  LAYER M2 ;
        RECT 3.884 16.184 6.356 16.216 ;
  LAYER M2 ;
        RECT 3.884 16.248 6.356 16.28 ;
  LAYER M2 ;
        RECT 3.884 16.312 6.356 16.344 ;
  LAYER M2 ;
        RECT 3.884 16.376 6.356 16.408 ;
  LAYER M2 ;
        RECT 3.884 16.44 6.356 16.472 ;
  LAYER M2 ;
        RECT 3.884 16.504 6.356 16.536 ;
  LAYER M2 ;
        RECT 3.884 16.568 6.356 16.6 ;
  LAYER M2 ;
        RECT 3.884 16.632 6.356 16.664 ;
  LAYER M2 ;
        RECT 3.884 16.696 6.356 16.728 ;
  LAYER M2 ;
        RECT 3.884 16.76 6.356 16.792 ;
  LAYER M2 ;
        RECT 3.884 16.824 6.356 16.856 ;
  LAYER M2 ;
        RECT 3.884 16.888 6.356 16.92 ;
  LAYER M2 ;
        RECT 3.884 16.952 6.356 16.984 ;
  LAYER M2 ;
        RECT 3.884 17.016 6.356 17.048 ;
  LAYER M2 ;
        RECT 3.884 17.08 6.356 17.112 ;
  LAYER M2 ;
        RECT 3.884 17.144 6.356 17.176 ;
  LAYER M2 ;
        RECT 3.884 17.208 6.356 17.24 ;
  LAYER M2 ;
        RECT 3.884 17.272 6.356 17.304 ;
  LAYER M2 ;
        RECT 3.884 17.336 6.356 17.368 ;
  LAYER M2 ;
        RECT 3.884 17.4 6.356 17.432 ;
  LAYER M2 ;
        RECT 3.884 17.464 6.356 17.496 ;
  LAYER M2 ;
        RECT 3.884 17.528 6.356 17.56 ;
  LAYER M2 ;
        RECT 3.884 17.592 6.356 17.624 ;
  LAYER M2 ;
        RECT 3.884 17.656 6.356 17.688 ;
  LAYER M2 ;
        RECT 3.884 17.72 6.356 17.752 ;
  LAYER M2 ;
        RECT 3.884 17.784 6.356 17.816 ;
  LAYER M2 ;
        RECT 3.884 17.848 6.356 17.88 ;
  LAYER M2 ;
        RECT 3.884 17.912 6.356 17.944 ;
  LAYER M3 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M3 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M3 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M3 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M3 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M3 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M3 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M3 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M3 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M3 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M3 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M3 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M3 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M3 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M3 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M3 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M3 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M3 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M3 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M3 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M3 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M3 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M3 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M3 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M3 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M3 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M3 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M3 ;
        RECT 5.632 15.588 5.664 18.096 ;
  LAYER M3 ;
        RECT 5.696 15.588 5.728 18.096 ;
  LAYER M3 ;
        RECT 5.76 15.588 5.792 18.096 ;
  LAYER M3 ;
        RECT 5.824 15.588 5.856 18.096 ;
  LAYER M3 ;
        RECT 5.888 15.588 5.92 18.096 ;
  LAYER M3 ;
        RECT 5.952 15.588 5.984 18.096 ;
  LAYER M3 ;
        RECT 6.016 15.588 6.048 18.096 ;
  LAYER M3 ;
        RECT 6.08 15.588 6.112 18.096 ;
  LAYER M3 ;
        RECT 6.144 15.588 6.176 18.096 ;
  LAYER M3 ;
        RECT 6.208 15.588 6.24 18.096 ;
  LAYER M3 ;
        RECT 6.304 15.588 6.336 18.096 ;
  LAYER M1 ;
        RECT 3.919 15.624 3.921 18.06 ;
  LAYER M1 ;
        RECT 3.999 15.624 4.001 18.06 ;
  LAYER M1 ;
        RECT 4.079 15.624 4.081 18.06 ;
  LAYER M1 ;
        RECT 4.159 15.624 4.161 18.06 ;
  LAYER M1 ;
        RECT 4.239 15.624 4.241 18.06 ;
  LAYER M1 ;
        RECT 4.319 15.624 4.321 18.06 ;
  LAYER M1 ;
        RECT 4.399 15.624 4.401 18.06 ;
  LAYER M1 ;
        RECT 4.479 15.624 4.481 18.06 ;
  LAYER M1 ;
        RECT 4.559 15.624 4.561 18.06 ;
  LAYER M1 ;
        RECT 4.639 15.624 4.641 18.06 ;
  LAYER M1 ;
        RECT 4.719 15.624 4.721 18.06 ;
  LAYER M1 ;
        RECT 4.799 15.624 4.801 18.06 ;
  LAYER M1 ;
        RECT 4.879 15.624 4.881 18.06 ;
  LAYER M1 ;
        RECT 4.959 15.624 4.961 18.06 ;
  LAYER M1 ;
        RECT 5.039 15.624 5.041 18.06 ;
  LAYER M1 ;
        RECT 5.119 15.624 5.121 18.06 ;
  LAYER M1 ;
        RECT 5.199 15.624 5.201 18.06 ;
  LAYER M1 ;
        RECT 5.279 15.624 5.281 18.06 ;
  LAYER M1 ;
        RECT 5.359 15.624 5.361 18.06 ;
  LAYER M1 ;
        RECT 5.439 15.624 5.441 18.06 ;
  LAYER M1 ;
        RECT 5.519 15.624 5.521 18.06 ;
  LAYER M1 ;
        RECT 5.599 15.624 5.601 18.06 ;
  LAYER M1 ;
        RECT 5.679 15.624 5.681 18.06 ;
  LAYER M1 ;
        RECT 5.759 15.624 5.761 18.06 ;
  LAYER M1 ;
        RECT 5.839 15.624 5.841 18.06 ;
  LAYER M1 ;
        RECT 5.919 15.624 5.921 18.06 ;
  LAYER M1 ;
        RECT 5.999 15.624 6.001 18.06 ;
  LAYER M1 ;
        RECT 6.079 15.624 6.081 18.06 ;
  LAYER M1 ;
        RECT 6.159 15.624 6.161 18.06 ;
  LAYER M1 ;
        RECT 6.239 15.624 6.241 18.06 ;
  LAYER M2 ;
        RECT 3.92 15.623 6.32 15.625 ;
  LAYER M2 ;
        RECT 3.92 15.707 6.32 15.709 ;
  LAYER M2 ;
        RECT 3.92 15.791 6.32 15.793 ;
  LAYER M2 ;
        RECT 3.92 15.875 6.32 15.877 ;
  LAYER M2 ;
        RECT 3.92 15.959 6.32 15.961 ;
  LAYER M2 ;
        RECT 3.92 16.043 6.32 16.045 ;
  LAYER M2 ;
        RECT 3.92 16.127 6.32 16.129 ;
  LAYER M2 ;
        RECT 3.92 16.211 6.32 16.213 ;
  LAYER M2 ;
        RECT 3.92 16.295 6.32 16.297 ;
  LAYER M2 ;
        RECT 3.92 16.379 6.32 16.381 ;
  LAYER M2 ;
        RECT 3.92 16.463 6.32 16.465 ;
  LAYER M2 ;
        RECT 3.92 16.547 6.32 16.549 ;
  LAYER M2 ;
        RECT 3.92 16.6305 6.32 16.6325 ;
  LAYER M2 ;
        RECT 3.92 16.715 6.32 16.717 ;
  LAYER M2 ;
        RECT 3.92 16.799 6.32 16.801 ;
  LAYER M2 ;
        RECT 3.92 16.883 6.32 16.885 ;
  LAYER M2 ;
        RECT 3.92 16.967 6.32 16.969 ;
  LAYER M2 ;
        RECT 3.92 17.051 6.32 17.053 ;
  LAYER M2 ;
        RECT 3.92 17.135 6.32 17.137 ;
  LAYER M2 ;
        RECT 3.92 17.219 6.32 17.221 ;
  LAYER M2 ;
        RECT 3.92 17.303 6.32 17.305 ;
  LAYER M2 ;
        RECT 3.92 17.387 6.32 17.389 ;
  LAYER M2 ;
        RECT 3.92 17.471 6.32 17.473 ;
  LAYER M2 ;
        RECT 3.92 17.555 6.32 17.557 ;
  LAYER M2 ;
        RECT 3.92 17.639 6.32 17.641 ;
  LAYER M2 ;
        RECT 3.92 17.723 6.32 17.725 ;
  LAYER M2 ;
        RECT 3.92 17.807 6.32 17.809 ;
  LAYER M2 ;
        RECT 3.92 17.891 6.32 17.893 ;
  LAYER M2 ;
        RECT 3.92 17.975 6.32 17.977 ;
  LAYER M1 ;
        RECT 3.904 18.528 3.936 21.036 ;
  LAYER M1 ;
        RECT 3.968 18.528 4 21.036 ;
  LAYER M1 ;
        RECT 4.032 18.528 4.064 21.036 ;
  LAYER M1 ;
        RECT 4.096 18.528 4.128 21.036 ;
  LAYER M1 ;
        RECT 4.16 18.528 4.192 21.036 ;
  LAYER M1 ;
        RECT 4.224 18.528 4.256 21.036 ;
  LAYER M1 ;
        RECT 4.288 18.528 4.32 21.036 ;
  LAYER M1 ;
        RECT 4.352 18.528 4.384 21.036 ;
  LAYER M1 ;
        RECT 4.416 18.528 4.448 21.036 ;
  LAYER M1 ;
        RECT 4.48 18.528 4.512 21.036 ;
  LAYER M1 ;
        RECT 4.544 18.528 4.576 21.036 ;
  LAYER M1 ;
        RECT 4.608 18.528 4.64 21.036 ;
  LAYER M1 ;
        RECT 4.672 18.528 4.704 21.036 ;
  LAYER M1 ;
        RECT 4.736 18.528 4.768 21.036 ;
  LAYER M1 ;
        RECT 4.8 18.528 4.832 21.036 ;
  LAYER M1 ;
        RECT 4.864 18.528 4.896 21.036 ;
  LAYER M1 ;
        RECT 4.928 18.528 4.96 21.036 ;
  LAYER M1 ;
        RECT 4.992 18.528 5.024 21.036 ;
  LAYER M1 ;
        RECT 5.056 18.528 5.088 21.036 ;
  LAYER M1 ;
        RECT 5.12 18.528 5.152 21.036 ;
  LAYER M1 ;
        RECT 5.184 18.528 5.216 21.036 ;
  LAYER M1 ;
        RECT 5.248 18.528 5.28 21.036 ;
  LAYER M1 ;
        RECT 5.312 18.528 5.344 21.036 ;
  LAYER M1 ;
        RECT 5.376 18.528 5.408 21.036 ;
  LAYER M1 ;
        RECT 5.44 18.528 5.472 21.036 ;
  LAYER M1 ;
        RECT 5.504 18.528 5.536 21.036 ;
  LAYER M1 ;
        RECT 5.568 18.528 5.6 21.036 ;
  LAYER M1 ;
        RECT 5.632 18.528 5.664 21.036 ;
  LAYER M1 ;
        RECT 5.696 18.528 5.728 21.036 ;
  LAYER M1 ;
        RECT 5.76 18.528 5.792 21.036 ;
  LAYER M1 ;
        RECT 5.824 18.528 5.856 21.036 ;
  LAYER M1 ;
        RECT 5.888 18.528 5.92 21.036 ;
  LAYER M1 ;
        RECT 5.952 18.528 5.984 21.036 ;
  LAYER M1 ;
        RECT 6.016 18.528 6.048 21.036 ;
  LAYER M1 ;
        RECT 6.08 18.528 6.112 21.036 ;
  LAYER M1 ;
        RECT 6.144 18.528 6.176 21.036 ;
  LAYER M1 ;
        RECT 6.208 18.528 6.24 21.036 ;
  LAYER M2 ;
        RECT 3.884 18.612 6.356 18.644 ;
  LAYER M2 ;
        RECT 3.884 18.676 6.356 18.708 ;
  LAYER M2 ;
        RECT 3.884 18.74 6.356 18.772 ;
  LAYER M2 ;
        RECT 3.884 18.804 6.356 18.836 ;
  LAYER M2 ;
        RECT 3.884 18.868 6.356 18.9 ;
  LAYER M2 ;
        RECT 3.884 18.932 6.356 18.964 ;
  LAYER M2 ;
        RECT 3.884 18.996 6.356 19.028 ;
  LAYER M2 ;
        RECT 3.884 19.06 6.356 19.092 ;
  LAYER M2 ;
        RECT 3.884 19.124 6.356 19.156 ;
  LAYER M2 ;
        RECT 3.884 19.188 6.356 19.22 ;
  LAYER M2 ;
        RECT 3.884 19.252 6.356 19.284 ;
  LAYER M2 ;
        RECT 3.884 19.316 6.356 19.348 ;
  LAYER M2 ;
        RECT 3.884 19.38 6.356 19.412 ;
  LAYER M2 ;
        RECT 3.884 19.444 6.356 19.476 ;
  LAYER M2 ;
        RECT 3.884 19.508 6.356 19.54 ;
  LAYER M2 ;
        RECT 3.884 19.572 6.356 19.604 ;
  LAYER M2 ;
        RECT 3.884 19.636 6.356 19.668 ;
  LAYER M2 ;
        RECT 3.884 19.7 6.356 19.732 ;
  LAYER M2 ;
        RECT 3.884 19.764 6.356 19.796 ;
  LAYER M2 ;
        RECT 3.884 19.828 6.356 19.86 ;
  LAYER M2 ;
        RECT 3.884 19.892 6.356 19.924 ;
  LAYER M2 ;
        RECT 3.884 19.956 6.356 19.988 ;
  LAYER M2 ;
        RECT 3.884 20.02 6.356 20.052 ;
  LAYER M2 ;
        RECT 3.884 20.084 6.356 20.116 ;
  LAYER M2 ;
        RECT 3.884 20.148 6.356 20.18 ;
  LAYER M2 ;
        RECT 3.884 20.212 6.356 20.244 ;
  LAYER M2 ;
        RECT 3.884 20.276 6.356 20.308 ;
  LAYER M2 ;
        RECT 3.884 20.34 6.356 20.372 ;
  LAYER M2 ;
        RECT 3.884 20.404 6.356 20.436 ;
  LAYER M2 ;
        RECT 3.884 20.468 6.356 20.5 ;
  LAYER M2 ;
        RECT 3.884 20.532 6.356 20.564 ;
  LAYER M2 ;
        RECT 3.884 20.596 6.356 20.628 ;
  LAYER M2 ;
        RECT 3.884 20.66 6.356 20.692 ;
  LAYER M2 ;
        RECT 3.884 20.724 6.356 20.756 ;
  LAYER M2 ;
        RECT 3.884 20.788 6.356 20.82 ;
  LAYER M2 ;
        RECT 3.884 20.852 6.356 20.884 ;
  LAYER M3 ;
        RECT 3.904 18.528 3.936 21.036 ;
  LAYER M3 ;
        RECT 3.968 18.528 4 21.036 ;
  LAYER M3 ;
        RECT 4.032 18.528 4.064 21.036 ;
  LAYER M3 ;
        RECT 4.096 18.528 4.128 21.036 ;
  LAYER M3 ;
        RECT 4.16 18.528 4.192 21.036 ;
  LAYER M3 ;
        RECT 4.224 18.528 4.256 21.036 ;
  LAYER M3 ;
        RECT 4.288 18.528 4.32 21.036 ;
  LAYER M3 ;
        RECT 4.352 18.528 4.384 21.036 ;
  LAYER M3 ;
        RECT 4.416 18.528 4.448 21.036 ;
  LAYER M3 ;
        RECT 4.48 18.528 4.512 21.036 ;
  LAYER M3 ;
        RECT 4.544 18.528 4.576 21.036 ;
  LAYER M3 ;
        RECT 4.608 18.528 4.64 21.036 ;
  LAYER M3 ;
        RECT 4.672 18.528 4.704 21.036 ;
  LAYER M3 ;
        RECT 4.736 18.528 4.768 21.036 ;
  LAYER M3 ;
        RECT 4.8 18.528 4.832 21.036 ;
  LAYER M3 ;
        RECT 4.864 18.528 4.896 21.036 ;
  LAYER M3 ;
        RECT 4.928 18.528 4.96 21.036 ;
  LAYER M3 ;
        RECT 4.992 18.528 5.024 21.036 ;
  LAYER M3 ;
        RECT 5.056 18.528 5.088 21.036 ;
  LAYER M3 ;
        RECT 5.12 18.528 5.152 21.036 ;
  LAYER M3 ;
        RECT 5.184 18.528 5.216 21.036 ;
  LAYER M3 ;
        RECT 5.248 18.528 5.28 21.036 ;
  LAYER M3 ;
        RECT 5.312 18.528 5.344 21.036 ;
  LAYER M3 ;
        RECT 5.376 18.528 5.408 21.036 ;
  LAYER M3 ;
        RECT 5.44 18.528 5.472 21.036 ;
  LAYER M3 ;
        RECT 5.504 18.528 5.536 21.036 ;
  LAYER M3 ;
        RECT 5.568 18.528 5.6 21.036 ;
  LAYER M3 ;
        RECT 5.632 18.528 5.664 21.036 ;
  LAYER M3 ;
        RECT 5.696 18.528 5.728 21.036 ;
  LAYER M3 ;
        RECT 5.76 18.528 5.792 21.036 ;
  LAYER M3 ;
        RECT 5.824 18.528 5.856 21.036 ;
  LAYER M3 ;
        RECT 5.888 18.528 5.92 21.036 ;
  LAYER M3 ;
        RECT 5.952 18.528 5.984 21.036 ;
  LAYER M3 ;
        RECT 6.016 18.528 6.048 21.036 ;
  LAYER M3 ;
        RECT 6.08 18.528 6.112 21.036 ;
  LAYER M3 ;
        RECT 6.144 18.528 6.176 21.036 ;
  LAYER M3 ;
        RECT 6.208 18.528 6.24 21.036 ;
  LAYER M3 ;
        RECT 6.304 18.528 6.336 21.036 ;
  LAYER M1 ;
        RECT 3.919 18.564 3.921 21 ;
  LAYER M1 ;
        RECT 3.999 18.564 4.001 21 ;
  LAYER M1 ;
        RECT 4.079 18.564 4.081 21 ;
  LAYER M1 ;
        RECT 4.159 18.564 4.161 21 ;
  LAYER M1 ;
        RECT 4.239 18.564 4.241 21 ;
  LAYER M1 ;
        RECT 4.319 18.564 4.321 21 ;
  LAYER M1 ;
        RECT 4.399 18.564 4.401 21 ;
  LAYER M1 ;
        RECT 4.479 18.564 4.481 21 ;
  LAYER M1 ;
        RECT 4.559 18.564 4.561 21 ;
  LAYER M1 ;
        RECT 4.639 18.564 4.641 21 ;
  LAYER M1 ;
        RECT 4.719 18.564 4.721 21 ;
  LAYER M1 ;
        RECT 4.799 18.564 4.801 21 ;
  LAYER M1 ;
        RECT 4.879 18.564 4.881 21 ;
  LAYER M1 ;
        RECT 4.959 18.564 4.961 21 ;
  LAYER M1 ;
        RECT 5.039 18.564 5.041 21 ;
  LAYER M1 ;
        RECT 5.119 18.564 5.121 21 ;
  LAYER M1 ;
        RECT 5.199 18.564 5.201 21 ;
  LAYER M1 ;
        RECT 5.279 18.564 5.281 21 ;
  LAYER M1 ;
        RECT 5.359 18.564 5.361 21 ;
  LAYER M1 ;
        RECT 5.439 18.564 5.441 21 ;
  LAYER M1 ;
        RECT 5.519 18.564 5.521 21 ;
  LAYER M1 ;
        RECT 5.599 18.564 5.601 21 ;
  LAYER M1 ;
        RECT 5.679 18.564 5.681 21 ;
  LAYER M1 ;
        RECT 5.759 18.564 5.761 21 ;
  LAYER M1 ;
        RECT 5.839 18.564 5.841 21 ;
  LAYER M1 ;
        RECT 5.919 18.564 5.921 21 ;
  LAYER M1 ;
        RECT 5.999 18.564 6.001 21 ;
  LAYER M1 ;
        RECT 6.079 18.564 6.081 21 ;
  LAYER M1 ;
        RECT 6.159 18.564 6.161 21 ;
  LAYER M1 ;
        RECT 6.239 18.564 6.241 21 ;
  LAYER M2 ;
        RECT 3.92 18.563 6.32 18.565 ;
  LAYER M2 ;
        RECT 3.92 18.647 6.32 18.649 ;
  LAYER M2 ;
        RECT 3.92 18.731 6.32 18.733 ;
  LAYER M2 ;
        RECT 3.92 18.815 6.32 18.817 ;
  LAYER M2 ;
        RECT 3.92 18.899 6.32 18.901 ;
  LAYER M2 ;
        RECT 3.92 18.983 6.32 18.985 ;
  LAYER M2 ;
        RECT 3.92 19.067 6.32 19.069 ;
  LAYER M2 ;
        RECT 3.92 19.151 6.32 19.153 ;
  LAYER M2 ;
        RECT 3.92 19.235 6.32 19.237 ;
  LAYER M2 ;
        RECT 3.92 19.319 6.32 19.321 ;
  LAYER M2 ;
        RECT 3.92 19.403 6.32 19.405 ;
  LAYER M2 ;
        RECT 3.92 19.487 6.32 19.489 ;
  LAYER M2 ;
        RECT 3.92 19.5705 6.32 19.5725 ;
  LAYER M2 ;
        RECT 3.92 19.655 6.32 19.657 ;
  LAYER M2 ;
        RECT 3.92 19.739 6.32 19.741 ;
  LAYER M2 ;
        RECT 3.92 19.823 6.32 19.825 ;
  LAYER M2 ;
        RECT 3.92 19.907 6.32 19.909 ;
  LAYER M2 ;
        RECT 3.92 19.991 6.32 19.993 ;
  LAYER M2 ;
        RECT 3.92 20.075 6.32 20.077 ;
  LAYER M2 ;
        RECT 3.92 20.159 6.32 20.161 ;
  LAYER M2 ;
        RECT 3.92 20.243 6.32 20.245 ;
  LAYER M2 ;
        RECT 3.92 20.327 6.32 20.329 ;
  LAYER M2 ;
        RECT 3.92 20.411 6.32 20.413 ;
  LAYER M2 ;
        RECT 3.92 20.495 6.32 20.497 ;
  LAYER M2 ;
        RECT 3.92 20.579 6.32 20.581 ;
  LAYER M2 ;
        RECT 3.92 20.663 6.32 20.665 ;
  LAYER M2 ;
        RECT 3.92 20.747 6.32 20.749 ;
  LAYER M2 ;
        RECT 3.92 20.831 6.32 20.833 ;
  LAYER M2 ;
        RECT 3.92 20.915 6.32 20.917 ;
  LAYER M1 ;
        RECT 3.904 21.468 3.936 23.976 ;
  LAYER M1 ;
        RECT 3.968 21.468 4 23.976 ;
  LAYER M1 ;
        RECT 4.032 21.468 4.064 23.976 ;
  LAYER M1 ;
        RECT 4.096 21.468 4.128 23.976 ;
  LAYER M1 ;
        RECT 4.16 21.468 4.192 23.976 ;
  LAYER M1 ;
        RECT 4.224 21.468 4.256 23.976 ;
  LAYER M1 ;
        RECT 4.288 21.468 4.32 23.976 ;
  LAYER M1 ;
        RECT 4.352 21.468 4.384 23.976 ;
  LAYER M1 ;
        RECT 4.416 21.468 4.448 23.976 ;
  LAYER M1 ;
        RECT 4.48 21.468 4.512 23.976 ;
  LAYER M1 ;
        RECT 4.544 21.468 4.576 23.976 ;
  LAYER M1 ;
        RECT 4.608 21.468 4.64 23.976 ;
  LAYER M1 ;
        RECT 4.672 21.468 4.704 23.976 ;
  LAYER M1 ;
        RECT 4.736 21.468 4.768 23.976 ;
  LAYER M1 ;
        RECT 4.8 21.468 4.832 23.976 ;
  LAYER M1 ;
        RECT 4.864 21.468 4.896 23.976 ;
  LAYER M1 ;
        RECT 4.928 21.468 4.96 23.976 ;
  LAYER M1 ;
        RECT 4.992 21.468 5.024 23.976 ;
  LAYER M1 ;
        RECT 5.056 21.468 5.088 23.976 ;
  LAYER M1 ;
        RECT 5.12 21.468 5.152 23.976 ;
  LAYER M1 ;
        RECT 5.184 21.468 5.216 23.976 ;
  LAYER M1 ;
        RECT 5.248 21.468 5.28 23.976 ;
  LAYER M1 ;
        RECT 5.312 21.468 5.344 23.976 ;
  LAYER M1 ;
        RECT 5.376 21.468 5.408 23.976 ;
  LAYER M1 ;
        RECT 5.44 21.468 5.472 23.976 ;
  LAYER M1 ;
        RECT 5.504 21.468 5.536 23.976 ;
  LAYER M1 ;
        RECT 5.568 21.468 5.6 23.976 ;
  LAYER M1 ;
        RECT 5.632 21.468 5.664 23.976 ;
  LAYER M1 ;
        RECT 5.696 21.468 5.728 23.976 ;
  LAYER M1 ;
        RECT 5.76 21.468 5.792 23.976 ;
  LAYER M1 ;
        RECT 5.824 21.468 5.856 23.976 ;
  LAYER M1 ;
        RECT 5.888 21.468 5.92 23.976 ;
  LAYER M1 ;
        RECT 5.952 21.468 5.984 23.976 ;
  LAYER M1 ;
        RECT 6.016 21.468 6.048 23.976 ;
  LAYER M1 ;
        RECT 6.08 21.468 6.112 23.976 ;
  LAYER M1 ;
        RECT 6.144 21.468 6.176 23.976 ;
  LAYER M1 ;
        RECT 6.208 21.468 6.24 23.976 ;
  LAYER M2 ;
        RECT 3.884 21.552 6.356 21.584 ;
  LAYER M2 ;
        RECT 3.884 21.616 6.356 21.648 ;
  LAYER M2 ;
        RECT 3.884 21.68 6.356 21.712 ;
  LAYER M2 ;
        RECT 3.884 21.744 6.356 21.776 ;
  LAYER M2 ;
        RECT 3.884 21.808 6.356 21.84 ;
  LAYER M2 ;
        RECT 3.884 21.872 6.356 21.904 ;
  LAYER M2 ;
        RECT 3.884 21.936 6.356 21.968 ;
  LAYER M2 ;
        RECT 3.884 22 6.356 22.032 ;
  LAYER M2 ;
        RECT 3.884 22.064 6.356 22.096 ;
  LAYER M2 ;
        RECT 3.884 22.128 6.356 22.16 ;
  LAYER M2 ;
        RECT 3.884 22.192 6.356 22.224 ;
  LAYER M2 ;
        RECT 3.884 22.256 6.356 22.288 ;
  LAYER M2 ;
        RECT 3.884 22.32 6.356 22.352 ;
  LAYER M2 ;
        RECT 3.884 22.384 6.356 22.416 ;
  LAYER M2 ;
        RECT 3.884 22.448 6.356 22.48 ;
  LAYER M2 ;
        RECT 3.884 22.512 6.356 22.544 ;
  LAYER M2 ;
        RECT 3.884 22.576 6.356 22.608 ;
  LAYER M2 ;
        RECT 3.884 22.64 6.356 22.672 ;
  LAYER M2 ;
        RECT 3.884 22.704 6.356 22.736 ;
  LAYER M2 ;
        RECT 3.884 22.768 6.356 22.8 ;
  LAYER M2 ;
        RECT 3.884 22.832 6.356 22.864 ;
  LAYER M2 ;
        RECT 3.884 22.896 6.356 22.928 ;
  LAYER M2 ;
        RECT 3.884 22.96 6.356 22.992 ;
  LAYER M2 ;
        RECT 3.884 23.024 6.356 23.056 ;
  LAYER M2 ;
        RECT 3.884 23.088 6.356 23.12 ;
  LAYER M2 ;
        RECT 3.884 23.152 6.356 23.184 ;
  LAYER M2 ;
        RECT 3.884 23.216 6.356 23.248 ;
  LAYER M2 ;
        RECT 3.884 23.28 6.356 23.312 ;
  LAYER M2 ;
        RECT 3.884 23.344 6.356 23.376 ;
  LAYER M2 ;
        RECT 3.884 23.408 6.356 23.44 ;
  LAYER M2 ;
        RECT 3.884 23.472 6.356 23.504 ;
  LAYER M2 ;
        RECT 3.884 23.536 6.356 23.568 ;
  LAYER M2 ;
        RECT 3.884 23.6 6.356 23.632 ;
  LAYER M2 ;
        RECT 3.884 23.664 6.356 23.696 ;
  LAYER M2 ;
        RECT 3.884 23.728 6.356 23.76 ;
  LAYER M2 ;
        RECT 3.884 23.792 6.356 23.824 ;
  LAYER M3 ;
        RECT 3.904 21.468 3.936 23.976 ;
  LAYER M3 ;
        RECT 3.968 21.468 4 23.976 ;
  LAYER M3 ;
        RECT 4.032 21.468 4.064 23.976 ;
  LAYER M3 ;
        RECT 4.096 21.468 4.128 23.976 ;
  LAYER M3 ;
        RECT 4.16 21.468 4.192 23.976 ;
  LAYER M3 ;
        RECT 4.224 21.468 4.256 23.976 ;
  LAYER M3 ;
        RECT 4.288 21.468 4.32 23.976 ;
  LAYER M3 ;
        RECT 4.352 21.468 4.384 23.976 ;
  LAYER M3 ;
        RECT 4.416 21.468 4.448 23.976 ;
  LAYER M3 ;
        RECT 4.48 21.468 4.512 23.976 ;
  LAYER M3 ;
        RECT 4.544 21.468 4.576 23.976 ;
  LAYER M3 ;
        RECT 4.608 21.468 4.64 23.976 ;
  LAYER M3 ;
        RECT 4.672 21.468 4.704 23.976 ;
  LAYER M3 ;
        RECT 4.736 21.468 4.768 23.976 ;
  LAYER M3 ;
        RECT 4.8 21.468 4.832 23.976 ;
  LAYER M3 ;
        RECT 4.864 21.468 4.896 23.976 ;
  LAYER M3 ;
        RECT 4.928 21.468 4.96 23.976 ;
  LAYER M3 ;
        RECT 4.992 21.468 5.024 23.976 ;
  LAYER M3 ;
        RECT 5.056 21.468 5.088 23.976 ;
  LAYER M3 ;
        RECT 5.12 21.468 5.152 23.976 ;
  LAYER M3 ;
        RECT 5.184 21.468 5.216 23.976 ;
  LAYER M3 ;
        RECT 5.248 21.468 5.28 23.976 ;
  LAYER M3 ;
        RECT 5.312 21.468 5.344 23.976 ;
  LAYER M3 ;
        RECT 5.376 21.468 5.408 23.976 ;
  LAYER M3 ;
        RECT 5.44 21.468 5.472 23.976 ;
  LAYER M3 ;
        RECT 5.504 21.468 5.536 23.976 ;
  LAYER M3 ;
        RECT 5.568 21.468 5.6 23.976 ;
  LAYER M3 ;
        RECT 5.632 21.468 5.664 23.976 ;
  LAYER M3 ;
        RECT 5.696 21.468 5.728 23.976 ;
  LAYER M3 ;
        RECT 5.76 21.468 5.792 23.976 ;
  LAYER M3 ;
        RECT 5.824 21.468 5.856 23.976 ;
  LAYER M3 ;
        RECT 5.888 21.468 5.92 23.976 ;
  LAYER M3 ;
        RECT 5.952 21.468 5.984 23.976 ;
  LAYER M3 ;
        RECT 6.016 21.468 6.048 23.976 ;
  LAYER M3 ;
        RECT 6.08 21.468 6.112 23.976 ;
  LAYER M3 ;
        RECT 6.144 21.468 6.176 23.976 ;
  LAYER M3 ;
        RECT 6.208 21.468 6.24 23.976 ;
  LAYER M3 ;
        RECT 6.304 21.468 6.336 23.976 ;
  LAYER M1 ;
        RECT 3.919 21.504 3.921 23.94 ;
  LAYER M1 ;
        RECT 3.999 21.504 4.001 23.94 ;
  LAYER M1 ;
        RECT 4.079 21.504 4.081 23.94 ;
  LAYER M1 ;
        RECT 4.159 21.504 4.161 23.94 ;
  LAYER M1 ;
        RECT 4.239 21.504 4.241 23.94 ;
  LAYER M1 ;
        RECT 4.319 21.504 4.321 23.94 ;
  LAYER M1 ;
        RECT 4.399 21.504 4.401 23.94 ;
  LAYER M1 ;
        RECT 4.479 21.504 4.481 23.94 ;
  LAYER M1 ;
        RECT 4.559 21.504 4.561 23.94 ;
  LAYER M1 ;
        RECT 4.639 21.504 4.641 23.94 ;
  LAYER M1 ;
        RECT 4.719 21.504 4.721 23.94 ;
  LAYER M1 ;
        RECT 4.799 21.504 4.801 23.94 ;
  LAYER M1 ;
        RECT 4.879 21.504 4.881 23.94 ;
  LAYER M1 ;
        RECT 4.959 21.504 4.961 23.94 ;
  LAYER M1 ;
        RECT 5.039 21.504 5.041 23.94 ;
  LAYER M1 ;
        RECT 5.119 21.504 5.121 23.94 ;
  LAYER M1 ;
        RECT 5.199 21.504 5.201 23.94 ;
  LAYER M1 ;
        RECT 5.279 21.504 5.281 23.94 ;
  LAYER M1 ;
        RECT 5.359 21.504 5.361 23.94 ;
  LAYER M1 ;
        RECT 5.439 21.504 5.441 23.94 ;
  LAYER M1 ;
        RECT 5.519 21.504 5.521 23.94 ;
  LAYER M1 ;
        RECT 5.599 21.504 5.601 23.94 ;
  LAYER M1 ;
        RECT 5.679 21.504 5.681 23.94 ;
  LAYER M1 ;
        RECT 5.759 21.504 5.761 23.94 ;
  LAYER M1 ;
        RECT 5.839 21.504 5.841 23.94 ;
  LAYER M1 ;
        RECT 5.919 21.504 5.921 23.94 ;
  LAYER M1 ;
        RECT 5.999 21.504 6.001 23.94 ;
  LAYER M1 ;
        RECT 6.079 21.504 6.081 23.94 ;
  LAYER M1 ;
        RECT 6.159 21.504 6.161 23.94 ;
  LAYER M1 ;
        RECT 6.239 21.504 6.241 23.94 ;
  LAYER M2 ;
        RECT 3.92 21.503 6.32 21.505 ;
  LAYER M2 ;
        RECT 3.92 21.587 6.32 21.589 ;
  LAYER M2 ;
        RECT 3.92 21.671 6.32 21.673 ;
  LAYER M2 ;
        RECT 3.92 21.755 6.32 21.757 ;
  LAYER M2 ;
        RECT 3.92 21.839 6.32 21.841 ;
  LAYER M2 ;
        RECT 3.92 21.923 6.32 21.925 ;
  LAYER M2 ;
        RECT 3.92 22.007 6.32 22.009 ;
  LAYER M2 ;
        RECT 3.92 22.091 6.32 22.093 ;
  LAYER M2 ;
        RECT 3.92 22.175 6.32 22.177 ;
  LAYER M2 ;
        RECT 3.92 22.259 6.32 22.261 ;
  LAYER M2 ;
        RECT 3.92 22.343 6.32 22.345 ;
  LAYER M2 ;
        RECT 3.92 22.427 6.32 22.429 ;
  LAYER M2 ;
        RECT 3.92 22.5105 6.32 22.5125 ;
  LAYER M2 ;
        RECT 3.92 22.595 6.32 22.597 ;
  LAYER M2 ;
        RECT 3.92 22.679 6.32 22.681 ;
  LAYER M2 ;
        RECT 3.92 22.763 6.32 22.765 ;
  LAYER M2 ;
        RECT 3.92 22.847 6.32 22.849 ;
  LAYER M2 ;
        RECT 3.92 22.931 6.32 22.933 ;
  LAYER M2 ;
        RECT 3.92 23.015 6.32 23.017 ;
  LAYER M2 ;
        RECT 3.92 23.099 6.32 23.101 ;
  LAYER M2 ;
        RECT 3.92 23.183 6.32 23.185 ;
  LAYER M2 ;
        RECT 3.92 23.267 6.32 23.269 ;
  LAYER M2 ;
        RECT 3.92 23.351 6.32 23.353 ;
  LAYER M2 ;
        RECT 3.92 23.435 6.32 23.437 ;
  LAYER M2 ;
        RECT 3.92 23.519 6.32 23.521 ;
  LAYER M2 ;
        RECT 3.92 23.603 6.32 23.605 ;
  LAYER M2 ;
        RECT 3.92 23.687 6.32 23.689 ;
  LAYER M2 ;
        RECT 3.92 23.771 6.32 23.773 ;
  LAYER M2 ;
        RECT 3.92 23.855 6.32 23.857 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M1 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M1 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M1 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M1 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M1 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M1 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M1 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M1 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M1 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M1 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M1 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M1 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M1 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M1 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M1 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M1 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M1 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M1 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M1 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M1 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M1 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M1 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M1 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M1 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M1 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M1 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M1 ;
        RECT 8.832 0.888 8.864 3.396 ;
  LAYER M1 ;
        RECT 8.896 0.888 8.928 3.396 ;
  LAYER M1 ;
        RECT 8.96 0.888 8.992 3.396 ;
  LAYER M1 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M1 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M1 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M1 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M1 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M1 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M1 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M2 ;
        RECT 7.084 0.972 9.556 1.004 ;
  LAYER M2 ;
        RECT 7.084 1.036 9.556 1.068 ;
  LAYER M2 ;
        RECT 7.084 1.1 9.556 1.132 ;
  LAYER M2 ;
        RECT 7.084 1.164 9.556 1.196 ;
  LAYER M2 ;
        RECT 7.084 1.228 9.556 1.26 ;
  LAYER M2 ;
        RECT 7.084 1.292 9.556 1.324 ;
  LAYER M2 ;
        RECT 7.084 1.356 9.556 1.388 ;
  LAYER M2 ;
        RECT 7.084 1.42 9.556 1.452 ;
  LAYER M2 ;
        RECT 7.084 1.484 9.556 1.516 ;
  LAYER M2 ;
        RECT 7.084 1.548 9.556 1.58 ;
  LAYER M2 ;
        RECT 7.084 1.612 9.556 1.644 ;
  LAYER M2 ;
        RECT 7.084 1.676 9.556 1.708 ;
  LAYER M2 ;
        RECT 7.084 1.74 9.556 1.772 ;
  LAYER M2 ;
        RECT 7.084 1.804 9.556 1.836 ;
  LAYER M2 ;
        RECT 7.084 1.868 9.556 1.9 ;
  LAYER M2 ;
        RECT 7.084 1.932 9.556 1.964 ;
  LAYER M2 ;
        RECT 7.084 1.996 9.556 2.028 ;
  LAYER M2 ;
        RECT 7.084 2.06 9.556 2.092 ;
  LAYER M2 ;
        RECT 7.084 2.124 9.556 2.156 ;
  LAYER M2 ;
        RECT 7.084 2.188 9.556 2.22 ;
  LAYER M2 ;
        RECT 7.084 2.252 9.556 2.284 ;
  LAYER M2 ;
        RECT 7.084 2.316 9.556 2.348 ;
  LAYER M2 ;
        RECT 7.084 2.38 9.556 2.412 ;
  LAYER M2 ;
        RECT 7.084 2.444 9.556 2.476 ;
  LAYER M2 ;
        RECT 7.084 2.508 9.556 2.54 ;
  LAYER M2 ;
        RECT 7.084 2.572 9.556 2.604 ;
  LAYER M2 ;
        RECT 7.084 2.636 9.556 2.668 ;
  LAYER M2 ;
        RECT 7.084 2.7 9.556 2.732 ;
  LAYER M2 ;
        RECT 7.084 2.764 9.556 2.796 ;
  LAYER M2 ;
        RECT 7.084 2.828 9.556 2.86 ;
  LAYER M2 ;
        RECT 7.084 2.892 9.556 2.924 ;
  LAYER M2 ;
        RECT 7.084 2.956 9.556 2.988 ;
  LAYER M2 ;
        RECT 7.084 3.02 9.556 3.052 ;
  LAYER M2 ;
        RECT 7.084 3.084 9.556 3.116 ;
  LAYER M2 ;
        RECT 7.084 3.148 9.556 3.18 ;
  LAYER M2 ;
        RECT 7.084 3.212 9.556 3.244 ;
  LAYER M3 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M3 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M3 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M3 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M3 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M3 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M3 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M3 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M3 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M3 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M3 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M3 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M3 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M3 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M3 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M3 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M3 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M3 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M3 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M3 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M3 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M3 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M3 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M3 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M3 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M3 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M3 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M3 ;
        RECT 8.832 0.888 8.864 3.396 ;
  LAYER M3 ;
        RECT 8.896 0.888 8.928 3.396 ;
  LAYER M3 ;
        RECT 8.96 0.888 8.992 3.396 ;
  LAYER M3 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M3 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M3 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M3 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M3 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M3 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M3 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M3 ;
        RECT 9.504 0.888 9.536 3.396 ;
  LAYER M1 ;
        RECT 7.119 0.924 7.121 3.36 ;
  LAYER M1 ;
        RECT 7.199 0.924 7.201 3.36 ;
  LAYER M1 ;
        RECT 7.279 0.924 7.281 3.36 ;
  LAYER M1 ;
        RECT 7.359 0.924 7.361 3.36 ;
  LAYER M1 ;
        RECT 7.439 0.924 7.441 3.36 ;
  LAYER M1 ;
        RECT 7.519 0.924 7.521 3.36 ;
  LAYER M1 ;
        RECT 7.599 0.924 7.601 3.36 ;
  LAYER M1 ;
        RECT 7.679 0.924 7.681 3.36 ;
  LAYER M1 ;
        RECT 7.759 0.924 7.761 3.36 ;
  LAYER M1 ;
        RECT 7.839 0.924 7.841 3.36 ;
  LAYER M1 ;
        RECT 7.919 0.924 7.921 3.36 ;
  LAYER M1 ;
        RECT 7.999 0.924 8.001 3.36 ;
  LAYER M1 ;
        RECT 8.079 0.924 8.081 3.36 ;
  LAYER M1 ;
        RECT 8.159 0.924 8.161 3.36 ;
  LAYER M1 ;
        RECT 8.239 0.924 8.241 3.36 ;
  LAYER M1 ;
        RECT 8.319 0.924 8.321 3.36 ;
  LAYER M1 ;
        RECT 8.399 0.924 8.401 3.36 ;
  LAYER M1 ;
        RECT 8.479 0.924 8.481 3.36 ;
  LAYER M1 ;
        RECT 8.559 0.924 8.561 3.36 ;
  LAYER M1 ;
        RECT 8.639 0.924 8.641 3.36 ;
  LAYER M1 ;
        RECT 8.719 0.924 8.721 3.36 ;
  LAYER M1 ;
        RECT 8.799 0.924 8.801 3.36 ;
  LAYER M1 ;
        RECT 8.879 0.924 8.881 3.36 ;
  LAYER M1 ;
        RECT 8.959 0.924 8.961 3.36 ;
  LAYER M1 ;
        RECT 9.039 0.924 9.041 3.36 ;
  LAYER M1 ;
        RECT 9.119 0.924 9.121 3.36 ;
  LAYER M1 ;
        RECT 9.199 0.924 9.201 3.36 ;
  LAYER M1 ;
        RECT 9.279 0.924 9.281 3.36 ;
  LAYER M1 ;
        RECT 9.359 0.924 9.361 3.36 ;
  LAYER M1 ;
        RECT 9.439 0.924 9.441 3.36 ;
  LAYER M2 ;
        RECT 7.12 0.923 9.52 0.925 ;
  LAYER M2 ;
        RECT 7.12 1.007 9.52 1.009 ;
  LAYER M2 ;
        RECT 7.12 1.091 9.52 1.093 ;
  LAYER M2 ;
        RECT 7.12 1.175 9.52 1.177 ;
  LAYER M2 ;
        RECT 7.12 1.259 9.52 1.261 ;
  LAYER M2 ;
        RECT 7.12 1.343 9.52 1.345 ;
  LAYER M2 ;
        RECT 7.12 1.427 9.52 1.429 ;
  LAYER M2 ;
        RECT 7.12 1.511 9.52 1.513 ;
  LAYER M2 ;
        RECT 7.12 1.595 9.52 1.597 ;
  LAYER M2 ;
        RECT 7.12 1.679 9.52 1.681 ;
  LAYER M2 ;
        RECT 7.12 1.763 9.52 1.765 ;
  LAYER M2 ;
        RECT 7.12 1.847 9.52 1.849 ;
  LAYER M2 ;
        RECT 7.12 1.9305 9.52 1.9325 ;
  LAYER M2 ;
        RECT 7.12 2.015 9.52 2.017 ;
  LAYER M2 ;
        RECT 7.12 2.099 9.52 2.101 ;
  LAYER M2 ;
        RECT 7.12 2.183 9.52 2.185 ;
  LAYER M2 ;
        RECT 7.12 2.267 9.52 2.269 ;
  LAYER M2 ;
        RECT 7.12 2.351 9.52 2.353 ;
  LAYER M2 ;
        RECT 7.12 2.435 9.52 2.437 ;
  LAYER M2 ;
        RECT 7.12 2.519 9.52 2.521 ;
  LAYER M2 ;
        RECT 7.12 2.603 9.52 2.605 ;
  LAYER M2 ;
        RECT 7.12 2.687 9.52 2.689 ;
  LAYER M2 ;
        RECT 7.12 2.771 9.52 2.773 ;
  LAYER M2 ;
        RECT 7.12 2.855 9.52 2.857 ;
  LAYER M2 ;
        RECT 7.12 2.939 9.52 2.941 ;
  LAYER M2 ;
        RECT 7.12 3.023 9.52 3.025 ;
  LAYER M2 ;
        RECT 7.12 3.107 9.52 3.109 ;
  LAYER M2 ;
        RECT 7.12 3.191 9.52 3.193 ;
  LAYER M2 ;
        RECT 7.12 3.275 9.52 3.277 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M1 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M1 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M1 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M1 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M1 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M1 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M1 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M1 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M1 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M1 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M1 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M1 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M1 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M1 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M1 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M1 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M1 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M1 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M1 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M1 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M1 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M1 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M1 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M1 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M1 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M1 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M1 ;
        RECT 8.832 3.828 8.864 6.336 ;
  LAYER M1 ;
        RECT 8.896 3.828 8.928 6.336 ;
  LAYER M1 ;
        RECT 8.96 3.828 8.992 6.336 ;
  LAYER M1 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M1 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M1 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M1 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M1 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M1 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M1 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M2 ;
        RECT 7.084 3.912 9.556 3.944 ;
  LAYER M2 ;
        RECT 7.084 3.976 9.556 4.008 ;
  LAYER M2 ;
        RECT 7.084 4.04 9.556 4.072 ;
  LAYER M2 ;
        RECT 7.084 4.104 9.556 4.136 ;
  LAYER M2 ;
        RECT 7.084 4.168 9.556 4.2 ;
  LAYER M2 ;
        RECT 7.084 4.232 9.556 4.264 ;
  LAYER M2 ;
        RECT 7.084 4.296 9.556 4.328 ;
  LAYER M2 ;
        RECT 7.084 4.36 9.556 4.392 ;
  LAYER M2 ;
        RECT 7.084 4.424 9.556 4.456 ;
  LAYER M2 ;
        RECT 7.084 4.488 9.556 4.52 ;
  LAYER M2 ;
        RECT 7.084 4.552 9.556 4.584 ;
  LAYER M2 ;
        RECT 7.084 4.616 9.556 4.648 ;
  LAYER M2 ;
        RECT 7.084 4.68 9.556 4.712 ;
  LAYER M2 ;
        RECT 7.084 4.744 9.556 4.776 ;
  LAYER M2 ;
        RECT 7.084 4.808 9.556 4.84 ;
  LAYER M2 ;
        RECT 7.084 4.872 9.556 4.904 ;
  LAYER M2 ;
        RECT 7.084 4.936 9.556 4.968 ;
  LAYER M2 ;
        RECT 7.084 5 9.556 5.032 ;
  LAYER M2 ;
        RECT 7.084 5.064 9.556 5.096 ;
  LAYER M2 ;
        RECT 7.084 5.128 9.556 5.16 ;
  LAYER M2 ;
        RECT 7.084 5.192 9.556 5.224 ;
  LAYER M2 ;
        RECT 7.084 5.256 9.556 5.288 ;
  LAYER M2 ;
        RECT 7.084 5.32 9.556 5.352 ;
  LAYER M2 ;
        RECT 7.084 5.384 9.556 5.416 ;
  LAYER M2 ;
        RECT 7.084 5.448 9.556 5.48 ;
  LAYER M2 ;
        RECT 7.084 5.512 9.556 5.544 ;
  LAYER M2 ;
        RECT 7.084 5.576 9.556 5.608 ;
  LAYER M2 ;
        RECT 7.084 5.64 9.556 5.672 ;
  LAYER M2 ;
        RECT 7.084 5.704 9.556 5.736 ;
  LAYER M2 ;
        RECT 7.084 5.768 9.556 5.8 ;
  LAYER M2 ;
        RECT 7.084 5.832 9.556 5.864 ;
  LAYER M2 ;
        RECT 7.084 5.896 9.556 5.928 ;
  LAYER M2 ;
        RECT 7.084 5.96 9.556 5.992 ;
  LAYER M2 ;
        RECT 7.084 6.024 9.556 6.056 ;
  LAYER M2 ;
        RECT 7.084 6.088 9.556 6.12 ;
  LAYER M2 ;
        RECT 7.084 6.152 9.556 6.184 ;
  LAYER M3 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M3 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M3 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M3 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M3 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M3 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M3 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M3 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M3 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M3 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M3 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M3 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M3 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M3 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M3 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M3 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M3 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M3 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M3 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M3 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M3 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M3 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M3 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M3 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M3 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M3 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M3 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M3 ;
        RECT 8.832 3.828 8.864 6.336 ;
  LAYER M3 ;
        RECT 8.896 3.828 8.928 6.336 ;
  LAYER M3 ;
        RECT 8.96 3.828 8.992 6.336 ;
  LAYER M3 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M3 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M3 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M3 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M3 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M3 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M3 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M3 ;
        RECT 9.504 3.828 9.536 6.336 ;
  LAYER M1 ;
        RECT 7.119 3.864 7.121 6.3 ;
  LAYER M1 ;
        RECT 7.199 3.864 7.201 6.3 ;
  LAYER M1 ;
        RECT 7.279 3.864 7.281 6.3 ;
  LAYER M1 ;
        RECT 7.359 3.864 7.361 6.3 ;
  LAYER M1 ;
        RECT 7.439 3.864 7.441 6.3 ;
  LAYER M1 ;
        RECT 7.519 3.864 7.521 6.3 ;
  LAYER M1 ;
        RECT 7.599 3.864 7.601 6.3 ;
  LAYER M1 ;
        RECT 7.679 3.864 7.681 6.3 ;
  LAYER M1 ;
        RECT 7.759 3.864 7.761 6.3 ;
  LAYER M1 ;
        RECT 7.839 3.864 7.841 6.3 ;
  LAYER M1 ;
        RECT 7.919 3.864 7.921 6.3 ;
  LAYER M1 ;
        RECT 7.999 3.864 8.001 6.3 ;
  LAYER M1 ;
        RECT 8.079 3.864 8.081 6.3 ;
  LAYER M1 ;
        RECT 8.159 3.864 8.161 6.3 ;
  LAYER M1 ;
        RECT 8.239 3.864 8.241 6.3 ;
  LAYER M1 ;
        RECT 8.319 3.864 8.321 6.3 ;
  LAYER M1 ;
        RECT 8.399 3.864 8.401 6.3 ;
  LAYER M1 ;
        RECT 8.479 3.864 8.481 6.3 ;
  LAYER M1 ;
        RECT 8.559 3.864 8.561 6.3 ;
  LAYER M1 ;
        RECT 8.639 3.864 8.641 6.3 ;
  LAYER M1 ;
        RECT 8.719 3.864 8.721 6.3 ;
  LAYER M1 ;
        RECT 8.799 3.864 8.801 6.3 ;
  LAYER M1 ;
        RECT 8.879 3.864 8.881 6.3 ;
  LAYER M1 ;
        RECT 8.959 3.864 8.961 6.3 ;
  LAYER M1 ;
        RECT 9.039 3.864 9.041 6.3 ;
  LAYER M1 ;
        RECT 9.119 3.864 9.121 6.3 ;
  LAYER M1 ;
        RECT 9.199 3.864 9.201 6.3 ;
  LAYER M1 ;
        RECT 9.279 3.864 9.281 6.3 ;
  LAYER M1 ;
        RECT 9.359 3.864 9.361 6.3 ;
  LAYER M1 ;
        RECT 9.439 3.864 9.441 6.3 ;
  LAYER M2 ;
        RECT 7.12 3.863 9.52 3.865 ;
  LAYER M2 ;
        RECT 7.12 3.947 9.52 3.949 ;
  LAYER M2 ;
        RECT 7.12 4.031 9.52 4.033 ;
  LAYER M2 ;
        RECT 7.12 4.115 9.52 4.117 ;
  LAYER M2 ;
        RECT 7.12 4.199 9.52 4.201 ;
  LAYER M2 ;
        RECT 7.12 4.283 9.52 4.285 ;
  LAYER M2 ;
        RECT 7.12 4.367 9.52 4.369 ;
  LAYER M2 ;
        RECT 7.12 4.451 9.52 4.453 ;
  LAYER M2 ;
        RECT 7.12 4.535 9.52 4.537 ;
  LAYER M2 ;
        RECT 7.12 4.619 9.52 4.621 ;
  LAYER M2 ;
        RECT 7.12 4.703 9.52 4.705 ;
  LAYER M2 ;
        RECT 7.12 4.787 9.52 4.789 ;
  LAYER M2 ;
        RECT 7.12 4.8705 9.52 4.8725 ;
  LAYER M2 ;
        RECT 7.12 4.955 9.52 4.957 ;
  LAYER M2 ;
        RECT 7.12 5.039 9.52 5.041 ;
  LAYER M2 ;
        RECT 7.12 5.123 9.52 5.125 ;
  LAYER M2 ;
        RECT 7.12 5.207 9.52 5.209 ;
  LAYER M2 ;
        RECT 7.12 5.291 9.52 5.293 ;
  LAYER M2 ;
        RECT 7.12 5.375 9.52 5.377 ;
  LAYER M2 ;
        RECT 7.12 5.459 9.52 5.461 ;
  LAYER M2 ;
        RECT 7.12 5.543 9.52 5.545 ;
  LAYER M2 ;
        RECT 7.12 5.627 9.52 5.629 ;
  LAYER M2 ;
        RECT 7.12 5.711 9.52 5.713 ;
  LAYER M2 ;
        RECT 7.12 5.795 9.52 5.797 ;
  LAYER M2 ;
        RECT 7.12 5.879 9.52 5.881 ;
  LAYER M2 ;
        RECT 7.12 5.963 9.52 5.965 ;
  LAYER M2 ;
        RECT 7.12 6.047 9.52 6.049 ;
  LAYER M2 ;
        RECT 7.12 6.131 9.52 6.133 ;
  LAYER M2 ;
        RECT 7.12 6.215 9.52 6.217 ;
  LAYER M1 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M1 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M1 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M1 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M1 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M1 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M1 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M1 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M1 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M1 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M1 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M1 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M1 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M1 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M1 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M1 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M1 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M1 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M1 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M1 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M1 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M1 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M1 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M1 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M1 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M1 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M1 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M1 ;
        RECT 8.832 6.768 8.864 9.276 ;
  LAYER M1 ;
        RECT 8.896 6.768 8.928 9.276 ;
  LAYER M1 ;
        RECT 8.96 6.768 8.992 9.276 ;
  LAYER M1 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M1 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M1 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M1 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M1 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M1 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M1 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M2 ;
        RECT 7.084 6.852 9.556 6.884 ;
  LAYER M2 ;
        RECT 7.084 6.916 9.556 6.948 ;
  LAYER M2 ;
        RECT 7.084 6.98 9.556 7.012 ;
  LAYER M2 ;
        RECT 7.084 7.044 9.556 7.076 ;
  LAYER M2 ;
        RECT 7.084 7.108 9.556 7.14 ;
  LAYER M2 ;
        RECT 7.084 7.172 9.556 7.204 ;
  LAYER M2 ;
        RECT 7.084 7.236 9.556 7.268 ;
  LAYER M2 ;
        RECT 7.084 7.3 9.556 7.332 ;
  LAYER M2 ;
        RECT 7.084 7.364 9.556 7.396 ;
  LAYER M2 ;
        RECT 7.084 7.428 9.556 7.46 ;
  LAYER M2 ;
        RECT 7.084 7.492 9.556 7.524 ;
  LAYER M2 ;
        RECT 7.084 7.556 9.556 7.588 ;
  LAYER M2 ;
        RECT 7.084 7.62 9.556 7.652 ;
  LAYER M2 ;
        RECT 7.084 7.684 9.556 7.716 ;
  LAYER M2 ;
        RECT 7.084 7.748 9.556 7.78 ;
  LAYER M2 ;
        RECT 7.084 7.812 9.556 7.844 ;
  LAYER M2 ;
        RECT 7.084 7.876 9.556 7.908 ;
  LAYER M2 ;
        RECT 7.084 7.94 9.556 7.972 ;
  LAYER M2 ;
        RECT 7.084 8.004 9.556 8.036 ;
  LAYER M2 ;
        RECT 7.084 8.068 9.556 8.1 ;
  LAYER M2 ;
        RECT 7.084 8.132 9.556 8.164 ;
  LAYER M2 ;
        RECT 7.084 8.196 9.556 8.228 ;
  LAYER M2 ;
        RECT 7.084 8.26 9.556 8.292 ;
  LAYER M2 ;
        RECT 7.084 8.324 9.556 8.356 ;
  LAYER M2 ;
        RECT 7.084 8.388 9.556 8.42 ;
  LAYER M2 ;
        RECT 7.084 8.452 9.556 8.484 ;
  LAYER M2 ;
        RECT 7.084 8.516 9.556 8.548 ;
  LAYER M2 ;
        RECT 7.084 8.58 9.556 8.612 ;
  LAYER M2 ;
        RECT 7.084 8.644 9.556 8.676 ;
  LAYER M2 ;
        RECT 7.084 8.708 9.556 8.74 ;
  LAYER M2 ;
        RECT 7.084 8.772 9.556 8.804 ;
  LAYER M2 ;
        RECT 7.084 8.836 9.556 8.868 ;
  LAYER M2 ;
        RECT 7.084 8.9 9.556 8.932 ;
  LAYER M2 ;
        RECT 7.084 8.964 9.556 8.996 ;
  LAYER M2 ;
        RECT 7.084 9.028 9.556 9.06 ;
  LAYER M2 ;
        RECT 7.084 9.092 9.556 9.124 ;
  LAYER M3 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M3 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M3 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M3 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M3 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M3 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M3 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M3 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M3 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M3 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M3 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M3 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M3 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M3 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M3 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M3 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M3 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M3 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M3 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M3 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M3 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M3 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M3 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M3 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M3 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M3 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M3 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M3 ;
        RECT 8.832 6.768 8.864 9.276 ;
  LAYER M3 ;
        RECT 8.896 6.768 8.928 9.276 ;
  LAYER M3 ;
        RECT 8.96 6.768 8.992 9.276 ;
  LAYER M3 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M3 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M3 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M3 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M3 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M3 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M3 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M3 ;
        RECT 9.504 6.768 9.536 9.276 ;
  LAYER M1 ;
        RECT 7.119 6.804 7.121 9.24 ;
  LAYER M1 ;
        RECT 7.199 6.804 7.201 9.24 ;
  LAYER M1 ;
        RECT 7.279 6.804 7.281 9.24 ;
  LAYER M1 ;
        RECT 7.359 6.804 7.361 9.24 ;
  LAYER M1 ;
        RECT 7.439 6.804 7.441 9.24 ;
  LAYER M1 ;
        RECT 7.519 6.804 7.521 9.24 ;
  LAYER M1 ;
        RECT 7.599 6.804 7.601 9.24 ;
  LAYER M1 ;
        RECT 7.679 6.804 7.681 9.24 ;
  LAYER M1 ;
        RECT 7.759 6.804 7.761 9.24 ;
  LAYER M1 ;
        RECT 7.839 6.804 7.841 9.24 ;
  LAYER M1 ;
        RECT 7.919 6.804 7.921 9.24 ;
  LAYER M1 ;
        RECT 7.999 6.804 8.001 9.24 ;
  LAYER M1 ;
        RECT 8.079 6.804 8.081 9.24 ;
  LAYER M1 ;
        RECT 8.159 6.804 8.161 9.24 ;
  LAYER M1 ;
        RECT 8.239 6.804 8.241 9.24 ;
  LAYER M1 ;
        RECT 8.319 6.804 8.321 9.24 ;
  LAYER M1 ;
        RECT 8.399 6.804 8.401 9.24 ;
  LAYER M1 ;
        RECT 8.479 6.804 8.481 9.24 ;
  LAYER M1 ;
        RECT 8.559 6.804 8.561 9.24 ;
  LAYER M1 ;
        RECT 8.639 6.804 8.641 9.24 ;
  LAYER M1 ;
        RECT 8.719 6.804 8.721 9.24 ;
  LAYER M1 ;
        RECT 8.799 6.804 8.801 9.24 ;
  LAYER M1 ;
        RECT 8.879 6.804 8.881 9.24 ;
  LAYER M1 ;
        RECT 8.959 6.804 8.961 9.24 ;
  LAYER M1 ;
        RECT 9.039 6.804 9.041 9.24 ;
  LAYER M1 ;
        RECT 9.119 6.804 9.121 9.24 ;
  LAYER M1 ;
        RECT 9.199 6.804 9.201 9.24 ;
  LAYER M1 ;
        RECT 9.279 6.804 9.281 9.24 ;
  LAYER M1 ;
        RECT 9.359 6.804 9.361 9.24 ;
  LAYER M1 ;
        RECT 9.439 6.804 9.441 9.24 ;
  LAYER M2 ;
        RECT 7.12 6.803 9.52 6.805 ;
  LAYER M2 ;
        RECT 7.12 6.887 9.52 6.889 ;
  LAYER M2 ;
        RECT 7.12 6.971 9.52 6.973 ;
  LAYER M2 ;
        RECT 7.12 7.055 9.52 7.057 ;
  LAYER M2 ;
        RECT 7.12 7.139 9.52 7.141 ;
  LAYER M2 ;
        RECT 7.12 7.223 9.52 7.225 ;
  LAYER M2 ;
        RECT 7.12 7.307 9.52 7.309 ;
  LAYER M2 ;
        RECT 7.12 7.391 9.52 7.393 ;
  LAYER M2 ;
        RECT 7.12 7.475 9.52 7.477 ;
  LAYER M2 ;
        RECT 7.12 7.559 9.52 7.561 ;
  LAYER M2 ;
        RECT 7.12 7.643 9.52 7.645 ;
  LAYER M2 ;
        RECT 7.12 7.727 9.52 7.729 ;
  LAYER M2 ;
        RECT 7.12 7.8105 9.52 7.8125 ;
  LAYER M2 ;
        RECT 7.12 7.895 9.52 7.897 ;
  LAYER M2 ;
        RECT 7.12 7.979 9.52 7.981 ;
  LAYER M2 ;
        RECT 7.12 8.063 9.52 8.065 ;
  LAYER M2 ;
        RECT 7.12 8.147 9.52 8.149 ;
  LAYER M2 ;
        RECT 7.12 8.231 9.52 8.233 ;
  LAYER M2 ;
        RECT 7.12 8.315 9.52 8.317 ;
  LAYER M2 ;
        RECT 7.12 8.399 9.52 8.401 ;
  LAYER M2 ;
        RECT 7.12 8.483 9.52 8.485 ;
  LAYER M2 ;
        RECT 7.12 8.567 9.52 8.569 ;
  LAYER M2 ;
        RECT 7.12 8.651 9.52 8.653 ;
  LAYER M2 ;
        RECT 7.12 8.735 9.52 8.737 ;
  LAYER M2 ;
        RECT 7.12 8.819 9.52 8.821 ;
  LAYER M2 ;
        RECT 7.12 8.903 9.52 8.905 ;
  LAYER M2 ;
        RECT 7.12 8.987 9.52 8.989 ;
  LAYER M2 ;
        RECT 7.12 9.071 9.52 9.073 ;
  LAYER M2 ;
        RECT 7.12 9.155 9.52 9.157 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M1 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M1 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M1 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M1 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M1 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M1 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M1 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M1 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M1 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M1 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M1 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M1 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M1 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M1 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M1 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M1 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M1 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M1 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M1 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M1 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M1 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M1 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M1 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M1 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M1 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M1 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M1 ;
        RECT 8.832 9.708 8.864 12.216 ;
  LAYER M1 ;
        RECT 8.896 9.708 8.928 12.216 ;
  LAYER M1 ;
        RECT 8.96 9.708 8.992 12.216 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M1 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M1 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M1 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M1 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M1 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M1 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M2 ;
        RECT 7.084 9.792 9.556 9.824 ;
  LAYER M2 ;
        RECT 7.084 9.856 9.556 9.888 ;
  LAYER M2 ;
        RECT 7.084 9.92 9.556 9.952 ;
  LAYER M2 ;
        RECT 7.084 9.984 9.556 10.016 ;
  LAYER M2 ;
        RECT 7.084 10.048 9.556 10.08 ;
  LAYER M2 ;
        RECT 7.084 10.112 9.556 10.144 ;
  LAYER M2 ;
        RECT 7.084 10.176 9.556 10.208 ;
  LAYER M2 ;
        RECT 7.084 10.24 9.556 10.272 ;
  LAYER M2 ;
        RECT 7.084 10.304 9.556 10.336 ;
  LAYER M2 ;
        RECT 7.084 10.368 9.556 10.4 ;
  LAYER M2 ;
        RECT 7.084 10.432 9.556 10.464 ;
  LAYER M2 ;
        RECT 7.084 10.496 9.556 10.528 ;
  LAYER M2 ;
        RECT 7.084 10.56 9.556 10.592 ;
  LAYER M2 ;
        RECT 7.084 10.624 9.556 10.656 ;
  LAYER M2 ;
        RECT 7.084 10.688 9.556 10.72 ;
  LAYER M2 ;
        RECT 7.084 10.752 9.556 10.784 ;
  LAYER M2 ;
        RECT 7.084 10.816 9.556 10.848 ;
  LAYER M2 ;
        RECT 7.084 10.88 9.556 10.912 ;
  LAYER M2 ;
        RECT 7.084 10.944 9.556 10.976 ;
  LAYER M2 ;
        RECT 7.084 11.008 9.556 11.04 ;
  LAYER M2 ;
        RECT 7.084 11.072 9.556 11.104 ;
  LAYER M2 ;
        RECT 7.084 11.136 9.556 11.168 ;
  LAYER M2 ;
        RECT 7.084 11.2 9.556 11.232 ;
  LAYER M2 ;
        RECT 7.084 11.264 9.556 11.296 ;
  LAYER M2 ;
        RECT 7.084 11.328 9.556 11.36 ;
  LAYER M2 ;
        RECT 7.084 11.392 9.556 11.424 ;
  LAYER M2 ;
        RECT 7.084 11.456 9.556 11.488 ;
  LAYER M2 ;
        RECT 7.084 11.52 9.556 11.552 ;
  LAYER M2 ;
        RECT 7.084 11.584 9.556 11.616 ;
  LAYER M2 ;
        RECT 7.084 11.648 9.556 11.68 ;
  LAYER M2 ;
        RECT 7.084 11.712 9.556 11.744 ;
  LAYER M2 ;
        RECT 7.084 11.776 9.556 11.808 ;
  LAYER M2 ;
        RECT 7.084 11.84 9.556 11.872 ;
  LAYER M2 ;
        RECT 7.084 11.904 9.556 11.936 ;
  LAYER M2 ;
        RECT 7.084 11.968 9.556 12 ;
  LAYER M2 ;
        RECT 7.084 12.032 9.556 12.064 ;
  LAYER M3 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M3 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M3 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M3 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M3 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M3 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M3 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M3 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M3 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M3 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M3 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M3 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M3 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M3 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M3 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M3 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M3 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M3 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M3 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M3 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M3 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M3 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M3 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M3 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M3 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M3 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M3 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M3 ;
        RECT 8.832 9.708 8.864 12.216 ;
  LAYER M3 ;
        RECT 8.896 9.708 8.928 12.216 ;
  LAYER M3 ;
        RECT 8.96 9.708 8.992 12.216 ;
  LAYER M3 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M3 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M3 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M3 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M3 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M3 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M3 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M3 ;
        RECT 9.504 9.708 9.536 12.216 ;
  LAYER M1 ;
        RECT 7.119 9.744 7.121 12.18 ;
  LAYER M1 ;
        RECT 7.199 9.744 7.201 12.18 ;
  LAYER M1 ;
        RECT 7.279 9.744 7.281 12.18 ;
  LAYER M1 ;
        RECT 7.359 9.744 7.361 12.18 ;
  LAYER M1 ;
        RECT 7.439 9.744 7.441 12.18 ;
  LAYER M1 ;
        RECT 7.519 9.744 7.521 12.18 ;
  LAYER M1 ;
        RECT 7.599 9.744 7.601 12.18 ;
  LAYER M1 ;
        RECT 7.679 9.744 7.681 12.18 ;
  LAYER M1 ;
        RECT 7.759 9.744 7.761 12.18 ;
  LAYER M1 ;
        RECT 7.839 9.744 7.841 12.18 ;
  LAYER M1 ;
        RECT 7.919 9.744 7.921 12.18 ;
  LAYER M1 ;
        RECT 7.999 9.744 8.001 12.18 ;
  LAYER M1 ;
        RECT 8.079 9.744 8.081 12.18 ;
  LAYER M1 ;
        RECT 8.159 9.744 8.161 12.18 ;
  LAYER M1 ;
        RECT 8.239 9.744 8.241 12.18 ;
  LAYER M1 ;
        RECT 8.319 9.744 8.321 12.18 ;
  LAYER M1 ;
        RECT 8.399 9.744 8.401 12.18 ;
  LAYER M1 ;
        RECT 8.479 9.744 8.481 12.18 ;
  LAYER M1 ;
        RECT 8.559 9.744 8.561 12.18 ;
  LAYER M1 ;
        RECT 8.639 9.744 8.641 12.18 ;
  LAYER M1 ;
        RECT 8.719 9.744 8.721 12.18 ;
  LAYER M1 ;
        RECT 8.799 9.744 8.801 12.18 ;
  LAYER M1 ;
        RECT 8.879 9.744 8.881 12.18 ;
  LAYER M1 ;
        RECT 8.959 9.744 8.961 12.18 ;
  LAYER M1 ;
        RECT 9.039 9.744 9.041 12.18 ;
  LAYER M1 ;
        RECT 9.119 9.744 9.121 12.18 ;
  LAYER M1 ;
        RECT 9.199 9.744 9.201 12.18 ;
  LAYER M1 ;
        RECT 9.279 9.744 9.281 12.18 ;
  LAYER M1 ;
        RECT 9.359 9.744 9.361 12.18 ;
  LAYER M1 ;
        RECT 9.439 9.744 9.441 12.18 ;
  LAYER M2 ;
        RECT 7.12 9.743 9.52 9.745 ;
  LAYER M2 ;
        RECT 7.12 9.827 9.52 9.829 ;
  LAYER M2 ;
        RECT 7.12 9.911 9.52 9.913 ;
  LAYER M2 ;
        RECT 7.12 9.995 9.52 9.997 ;
  LAYER M2 ;
        RECT 7.12 10.079 9.52 10.081 ;
  LAYER M2 ;
        RECT 7.12 10.163 9.52 10.165 ;
  LAYER M2 ;
        RECT 7.12 10.247 9.52 10.249 ;
  LAYER M2 ;
        RECT 7.12 10.331 9.52 10.333 ;
  LAYER M2 ;
        RECT 7.12 10.415 9.52 10.417 ;
  LAYER M2 ;
        RECT 7.12 10.499 9.52 10.501 ;
  LAYER M2 ;
        RECT 7.12 10.583 9.52 10.585 ;
  LAYER M2 ;
        RECT 7.12 10.667 9.52 10.669 ;
  LAYER M2 ;
        RECT 7.12 10.7505 9.52 10.7525 ;
  LAYER M2 ;
        RECT 7.12 10.835 9.52 10.837 ;
  LAYER M2 ;
        RECT 7.12 10.919 9.52 10.921 ;
  LAYER M2 ;
        RECT 7.12 11.003 9.52 11.005 ;
  LAYER M2 ;
        RECT 7.12 11.087 9.52 11.089 ;
  LAYER M2 ;
        RECT 7.12 11.171 9.52 11.173 ;
  LAYER M2 ;
        RECT 7.12 11.255 9.52 11.257 ;
  LAYER M2 ;
        RECT 7.12 11.339 9.52 11.341 ;
  LAYER M2 ;
        RECT 7.12 11.423 9.52 11.425 ;
  LAYER M2 ;
        RECT 7.12 11.507 9.52 11.509 ;
  LAYER M2 ;
        RECT 7.12 11.591 9.52 11.593 ;
  LAYER M2 ;
        RECT 7.12 11.675 9.52 11.677 ;
  LAYER M2 ;
        RECT 7.12 11.759 9.52 11.761 ;
  LAYER M2 ;
        RECT 7.12 11.843 9.52 11.845 ;
  LAYER M2 ;
        RECT 7.12 11.927 9.52 11.929 ;
  LAYER M2 ;
        RECT 7.12 12.011 9.52 12.013 ;
  LAYER M2 ;
        RECT 7.12 12.095 9.52 12.097 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M1 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M1 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M1 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M1 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M1 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M1 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M1 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M1 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M1 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M1 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M1 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M1 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M1 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M1 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M1 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M1 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M1 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M1 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M1 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M1 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M1 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M1 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M1 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M1 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M1 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M1 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M1 ;
        RECT 8.832 12.648 8.864 15.156 ;
  LAYER M1 ;
        RECT 8.896 12.648 8.928 15.156 ;
  LAYER M1 ;
        RECT 8.96 12.648 8.992 15.156 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M1 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M1 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M1 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M1 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M1 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M1 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M2 ;
        RECT 7.084 12.732 9.556 12.764 ;
  LAYER M2 ;
        RECT 7.084 12.796 9.556 12.828 ;
  LAYER M2 ;
        RECT 7.084 12.86 9.556 12.892 ;
  LAYER M2 ;
        RECT 7.084 12.924 9.556 12.956 ;
  LAYER M2 ;
        RECT 7.084 12.988 9.556 13.02 ;
  LAYER M2 ;
        RECT 7.084 13.052 9.556 13.084 ;
  LAYER M2 ;
        RECT 7.084 13.116 9.556 13.148 ;
  LAYER M2 ;
        RECT 7.084 13.18 9.556 13.212 ;
  LAYER M2 ;
        RECT 7.084 13.244 9.556 13.276 ;
  LAYER M2 ;
        RECT 7.084 13.308 9.556 13.34 ;
  LAYER M2 ;
        RECT 7.084 13.372 9.556 13.404 ;
  LAYER M2 ;
        RECT 7.084 13.436 9.556 13.468 ;
  LAYER M2 ;
        RECT 7.084 13.5 9.556 13.532 ;
  LAYER M2 ;
        RECT 7.084 13.564 9.556 13.596 ;
  LAYER M2 ;
        RECT 7.084 13.628 9.556 13.66 ;
  LAYER M2 ;
        RECT 7.084 13.692 9.556 13.724 ;
  LAYER M2 ;
        RECT 7.084 13.756 9.556 13.788 ;
  LAYER M2 ;
        RECT 7.084 13.82 9.556 13.852 ;
  LAYER M2 ;
        RECT 7.084 13.884 9.556 13.916 ;
  LAYER M2 ;
        RECT 7.084 13.948 9.556 13.98 ;
  LAYER M2 ;
        RECT 7.084 14.012 9.556 14.044 ;
  LAYER M2 ;
        RECT 7.084 14.076 9.556 14.108 ;
  LAYER M2 ;
        RECT 7.084 14.14 9.556 14.172 ;
  LAYER M2 ;
        RECT 7.084 14.204 9.556 14.236 ;
  LAYER M2 ;
        RECT 7.084 14.268 9.556 14.3 ;
  LAYER M2 ;
        RECT 7.084 14.332 9.556 14.364 ;
  LAYER M2 ;
        RECT 7.084 14.396 9.556 14.428 ;
  LAYER M2 ;
        RECT 7.084 14.46 9.556 14.492 ;
  LAYER M2 ;
        RECT 7.084 14.524 9.556 14.556 ;
  LAYER M2 ;
        RECT 7.084 14.588 9.556 14.62 ;
  LAYER M2 ;
        RECT 7.084 14.652 9.556 14.684 ;
  LAYER M2 ;
        RECT 7.084 14.716 9.556 14.748 ;
  LAYER M2 ;
        RECT 7.084 14.78 9.556 14.812 ;
  LAYER M2 ;
        RECT 7.084 14.844 9.556 14.876 ;
  LAYER M2 ;
        RECT 7.084 14.908 9.556 14.94 ;
  LAYER M2 ;
        RECT 7.084 14.972 9.556 15.004 ;
  LAYER M3 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M3 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M3 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M3 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M3 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M3 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M3 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M3 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M3 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M3 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M3 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M3 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M3 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M3 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M3 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M3 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M3 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M3 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M3 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M3 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M3 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M3 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M3 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M3 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M3 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M3 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M3 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M3 ;
        RECT 8.832 12.648 8.864 15.156 ;
  LAYER M3 ;
        RECT 8.896 12.648 8.928 15.156 ;
  LAYER M3 ;
        RECT 8.96 12.648 8.992 15.156 ;
  LAYER M3 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M3 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M3 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M3 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M3 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M3 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M3 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M3 ;
        RECT 9.504 12.648 9.536 15.156 ;
  LAYER M1 ;
        RECT 7.119 12.684 7.121 15.12 ;
  LAYER M1 ;
        RECT 7.199 12.684 7.201 15.12 ;
  LAYER M1 ;
        RECT 7.279 12.684 7.281 15.12 ;
  LAYER M1 ;
        RECT 7.359 12.684 7.361 15.12 ;
  LAYER M1 ;
        RECT 7.439 12.684 7.441 15.12 ;
  LAYER M1 ;
        RECT 7.519 12.684 7.521 15.12 ;
  LAYER M1 ;
        RECT 7.599 12.684 7.601 15.12 ;
  LAYER M1 ;
        RECT 7.679 12.684 7.681 15.12 ;
  LAYER M1 ;
        RECT 7.759 12.684 7.761 15.12 ;
  LAYER M1 ;
        RECT 7.839 12.684 7.841 15.12 ;
  LAYER M1 ;
        RECT 7.919 12.684 7.921 15.12 ;
  LAYER M1 ;
        RECT 7.999 12.684 8.001 15.12 ;
  LAYER M1 ;
        RECT 8.079 12.684 8.081 15.12 ;
  LAYER M1 ;
        RECT 8.159 12.684 8.161 15.12 ;
  LAYER M1 ;
        RECT 8.239 12.684 8.241 15.12 ;
  LAYER M1 ;
        RECT 8.319 12.684 8.321 15.12 ;
  LAYER M1 ;
        RECT 8.399 12.684 8.401 15.12 ;
  LAYER M1 ;
        RECT 8.479 12.684 8.481 15.12 ;
  LAYER M1 ;
        RECT 8.559 12.684 8.561 15.12 ;
  LAYER M1 ;
        RECT 8.639 12.684 8.641 15.12 ;
  LAYER M1 ;
        RECT 8.719 12.684 8.721 15.12 ;
  LAYER M1 ;
        RECT 8.799 12.684 8.801 15.12 ;
  LAYER M1 ;
        RECT 8.879 12.684 8.881 15.12 ;
  LAYER M1 ;
        RECT 8.959 12.684 8.961 15.12 ;
  LAYER M1 ;
        RECT 9.039 12.684 9.041 15.12 ;
  LAYER M1 ;
        RECT 9.119 12.684 9.121 15.12 ;
  LAYER M1 ;
        RECT 9.199 12.684 9.201 15.12 ;
  LAYER M1 ;
        RECT 9.279 12.684 9.281 15.12 ;
  LAYER M1 ;
        RECT 9.359 12.684 9.361 15.12 ;
  LAYER M1 ;
        RECT 9.439 12.684 9.441 15.12 ;
  LAYER M2 ;
        RECT 7.12 12.683 9.52 12.685 ;
  LAYER M2 ;
        RECT 7.12 12.767 9.52 12.769 ;
  LAYER M2 ;
        RECT 7.12 12.851 9.52 12.853 ;
  LAYER M2 ;
        RECT 7.12 12.935 9.52 12.937 ;
  LAYER M2 ;
        RECT 7.12 13.019 9.52 13.021 ;
  LAYER M2 ;
        RECT 7.12 13.103 9.52 13.105 ;
  LAYER M2 ;
        RECT 7.12 13.187 9.52 13.189 ;
  LAYER M2 ;
        RECT 7.12 13.271 9.52 13.273 ;
  LAYER M2 ;
        RECT 7.12 13.355 9.52 13.357 ;
  LAYER M2 ;
        RECT 7.12 13.439 9.52 13.441 ;
  LAYER M2 ;
        RECT 7.12 13.523 9.52 13.525 ;
  LAYER M2 ;
        RECT 7.12 13.607 9.52 13.609 ;
  LAYER M2 ;
        RECT 7.12 13.6905 9.52 13.6925 ;
  LAYER M2 ;
        RECT 7.12 13.775 9.52 13.777 ;
  LAYER M2 ;
        RECT 7.12 13.859 9.52 13.861 ;
  LAYER M2 ;
        RECT 7.12 13.943 9.52 13.945 ;
  LAYER M2 ;
        RECT 7.12 14.027 9.52 14.029 ;
  LAYER M2 ;
        RECT 7.12 14.111 9.52 14.113 ;
  LAYER M2 ;
        RECT 7.12 14.195 9.52 14.197 ;
  LAYER M2 ;
        RECT 7.12 14.279 9.52 14.281 ;
  LAYER M2 ;
        RECT 7.12 14.363 9.52 14.365 ;
  LAYER M2 ;
        RECT 7.12 14.447 9.52 14.449 ;
  LAYER M2 ;
        RECT 7.12 14.531 9.52 14.533 ;
  LAYER M2 ;
        RECT 7.12 14.615 9.52 14.617 ;
  LAYER M2 ;
        RECT 7.12 14.699 9.52 14.701 ;
  LAYER M2 ;
        RECT 7.12 14.783 9.52 14.785 ;
  LAYER M2 ;
        RECT 7.12 14.867 9.52 14.869 ;
  LAYER M2 ;
        RECT 7.12 14.951 9.52 14.953 ;
  LAYER M2 ;
        RECT 7.12 15.035 9.52 15.037 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M1 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M1 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M1 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M1 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M1 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M1 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M1 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M1 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M1 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M1 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M1 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M1 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M1 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M1 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M1 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M1 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M1 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M1 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M1 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M1 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M1 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M1 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M1 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M1 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M1 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M1 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M1 ;
        RECT 8.832 15.588 8.864 18.096 ;
  LAYER M1 ;
        RECT 8.896 15.588 8.928 18.096 ;
  LAYER M1 ;
        RECT 8.96 15.588 8.992 18.096 ;
  LAYER M1 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M1 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M1 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M1 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M1 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M1 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M1 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M2 ;
        RECT 7.084 15.672 9.556 15.704 ;
  LAYER M2 ;
        RECT 7.084 15.736 9.556 15.768 ;
  LAYER M2 ;
        RECT 7.084 15.8 9.556 15.832 ;
  LAYER M2 ;
        RECT 7.084 15.864 9.556 15.896 ;
  LAYER M2 ;
        RECT 7.084 15.928 9.556 15.96 ;
  LAYER M2 ;
        RECT 7.084 15.992 9.556 16.024 ;
  LAYER M2 ;
        RECT 7.084 16.056 9.556 16.088 ;
  LAYER M2 ;
        RECT 7.084 16.12 9.556 16.152 ;
  LAYER M2 ;
        RECT 7.084 16.184 9.556 16.216 ;
  LAYER M2 ;
        RECT 7.084 16.248 9.556 16.28 ;
  LAYER M2 ;
        RECT 7.084 16.312 9.556 16.344 ;
  LAYER M2 ;
        RECT 7.084 16.376 9.556 16.408 ;
  LAYER M2 ;
        RECT 7.084 16.44 9.556 16.472 ;
  LAYER M2 ;
        RECT 7.084 16.504 9.556 16.536 ;
  LAYER M2 ;
        RECT 7.084 16.568 9.556 16.6 ;
  LAYER M2 ;
        RECT 7.084 16.632 9.556 16.664 ;
  LAYER M2 ;
        RECT 7.084 16.696 9.556 16.728 ;
  LAYER M2 ;
        RECT 7.084 16.76 9.556 16.792 ;
  LAYER M2 ;
        RECT 7.084 16.824 9.556 16.856 ;
  LAYER M2 ;
        RECT 7.084 16.888 9.556 16.92 ;
  LAYER M2 ;
        RECT 7.084 16.952 9.556 16.984 ;
  LAYER M2 ;
        RECT 7.084 17.016 9.556 17.048 ;
  LAYER M2 ;
        RECT 7.084 17.08 9.556 17.112 ;
  LAYER M2 ;
        RECT 7.084 17.144 9.556 17.176 ;
  LAYER M2 ;
        RECT 7.084 17.208 9.556 17.24 ;
  LAYER M2 ;
        RECT 7.084 17.272 9.556 17.304 ;
  LAYER M2 ;
        RECT 7.084 17.336 9.556 17.368 ;
  LAYER M2 ;
        RECT 7.084 17.4 9.556 17.432 ;
  LAYER M2 ;
        RECT 7.084 17.464 9.556 17.496 ;
  LAYER M2 ;
        RECT 7.084 17.528 9.556 17.56 ;
  LAYER M2 ;
        RECT 7.084 17.592 9.556 17.624 ;
  LAYER M2 ;
        RECT 7.084 17.656 9.556 17.688 ;
  LAYER M2 ;
        RECT 7.084 17.72 9.556 17.752 ;
  LAYER M2 ;
        RECT 7.084 17.784 9.556 17.816 ;
  LAYER M2 ;
        RECT 7.084 17.848 9.556 17.88 ;
  LAYER M2 ;
        RECT 7.084 17.912 9.556 17.944 ;
  LAYER M3 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M3 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M3 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M3 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M3 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M3 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M3 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M3 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M3 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M3 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M3 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M3 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M3 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M3 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M3 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M3 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M3 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M3 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M3 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M3 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M3 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M3 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M3 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M3 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M3 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M3 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M3 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M3 ;
        RECT 8.832 15.588 8.864 18.096 ;
  LAYER M3 ;
        RECT 8.896 15.588 8.928 18.096 ;
  LAYER M3 ;
        RECT 8.96 15.588 8.992 18.096 ;
  LAYER M3 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M3 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M3 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M3 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M3 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M3 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M3 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M3 ;
        RECT 9.504 15.588 9.536 18.096 ;
  LAYER M1 ;
        RECT 7.119 15.624 7.121 18.06 ;
  LAYER M1 ;
        RECT 7.199 15.624 7.201 18.06 ;
  LAYER M1 ;
        RECT 7.279 15.624 7.281 18.06 ;
  LAYER M1 ;
        RECT 7.359 15.624 7.361 18.06 ;
  LAYER M1 ;
        RECT 7.439 15.624 7.441 18.06 ;
  LAYER M1 ;
        RECT 7.519 15.624 7.521 18.06 ;
  LAYER M1 ;
        RECT 7.599 15.624 7.601 18.06 ;
  LAYER M1 ;
        RECT 7.679 15.624 7.681 18.06 ;
  LAYER M1 ;
        RECT 7.759 15.624 7.761 18.06 ;
  LAYER M1 ;
        RECT 7.839 15.624 7.841 18.06 ;
  LAYER M1 ;
        RECT 7.919 15.624 7.921 18.06 ;
  LAYER M1 ;
        RECT 7.999 15.624 8.001 18.06 ;
  LAYER M1 ;
        RECT 8.079 15.624 8.081 18.06 ;
  LAYER M1 ;
        RECT 8.159 15.624 8.161 18.06 ;
  LAYER M1 ;
        RECT 8.239 15.624 8.241 18.06 ;
  LAYER M1 ;
        RECT 8.319 15.624 8.321 18.06 ;
  LAYER M1 ;
        RECT 8.399 15.624 8.401 18.06 ;
  LAYER M1 ;
        RECT 8.479 15.624 8.481 18.06 ;
  LAYER M1 ;
        RECT 8.559 15.624 8.561 18.06 ;
  LAYER M1 ;
        RECT 8.639 15.624 8.641 18.06 ;
  LAYER M1 ;
        RECT 8.719 15.624 8.721 18.06 ;
  LAYER M1 ;
        RECT 8.799 15.624 8.801 18.06 ;
  LAYER M1 ;
        RECT 8.879 15.624 8.881 18.06 ;
  LAYER M1 ;
        RECT 8.959 15.624 8.961 18.06 ;
  LAYER M1 ;
        RECT 9.039 15.624 9.041 18.06 ;
  LAYER M1 ;
        RECT 9.119 15.624 9.121 18.06 ;
  LAYER M1 ;
        RECT 9.199 15.624 9.201 18.06 ;
  LAYER M1 ;
        RECT 9.279 15.624 9.281 18.06 ;
  LAYER M1 ;
        RECT 9.359 15.624 9.361 18.06 ;
  LAYER M1 ;
        RECT 9.439 15.624 9.441 18.06 ;
  LAYER M2 ;
        RECT 7.12 15.623 9.52 15.625 ;
  LAYER M2 ;
        RECT 7.12 15.707 9.52 15.709 ;
  LAYER M2 ;
        RECT 7.12 15.791 9.52 15.793 ;
  LAYER M2 ;
        RECT 7.12 15.875 9.52 15.877 ;
  LAYER M2 ;
        RECT 7.12 15.959 9.52 15.961 ;
  LAYER M2 ;
        RECT 7.12 16.043 9.52 16.045 ;
  LAYER M2 ;
        RECT 7.12 16.127 9.52 16.129 ;
  LAYER M2 ;
        RECT 7.12 16.211 9.52 16.213 ;
  LAYER M2 ;
        RECT 7.12 16.295 9.52 16.297 ;
  LAYER M2 ;
        RECT 7.12 16.379 9.52 16.381 ;
  LAYER M2 ;
        RECT 7.12 16.463 9.52 16.465 ;
  LAYER M2 ;
        RECT 7.12 16.547 9.52 16.549 ;
  LAYER M2 ;
        RECT 7.12 16.6305 9.52 16.6325 ;
  LAYER M2 ;
        RECT 7.12 16.715 9.52 16.717 ;
  LAYER M2 ;
        RECT 7.12 16.799 9.52 16.801 ;
  LAYER M2 ;
        RECT 7.12 16.883 9.52 16.885 ;
  LAYER M2 ;
        RECT 7.12 16.967 9.52 16.969 ;
  LAYER M2 ;
        RECT 7.12 17.051 9.52 17.053 ;
  LAYER M2 ;
        RECT 7.12 17.135 9.52 17.137 ;
  LAYER M2 ;
        RECT 7.12 17.219 9.52 17.221 ;
  LAYER M2 ;
        RECT 7.12 17.303 9.52 17.305 ;
  LAYER M2 ;
        RECT 7.12 17.387 9.52 17.389 ;
  LAYER M2 ;
        RECT 7.12 17.471 9.52 17.473 ;
  LAYER M2 ;
        RECT 7.12 17.555 9.52 17.557 ;
  LAYER M2 ;
        RECT 7.12 17.639 9.52 17.641 ;
  LAYER M2 ;
        RECT 7.12 17.723 9.52 17.725 ;
  LAYER M2 ;
        RECT 7.12 17.807 9.52 17.809 ;
  LAYER M2 ;
        RECT 7.12 17.891 9.52 17.893 ;
  LAYER M2 ;
        RECT 7.12 17.975 9.52 17.977 ;
  LAYER M1 ;
        RECT 7.104 18.528 7.136 21.036 ;
  LAYER M1 ;
        RECT 7.168 18.528 7.2 21.036 ;
  LAYER M1 ;
        RECT 7.232 18.528 7.264 21.036 ;
  LAYER M1 ;
        RECT 7.296 18.528 7.328 21.036 ;
  LAYER M1 ;
        RECT 7.36 18.528 7.392 21.036 ;
  LAYER M1 ;
        RECT 7.424 18.528 7.456 21.036 ;
  LAYER M1 ;
        RECT 7.488 18.528 7.52 21.036 ;
  LAYER M1 ;
        RECT 7.552 18.528 7.584 21.036 ;
  LAYER M1 ;
        RECT 7.616 18.528 7.648 21.036 ;
  LAYER M1 ;
        RECT 7.68 18.528 7.712 21.036 ;
  LAYER M1 ;
        RECT 7.744 18.528 7.776 21.036 ;
  LAYER M1 ;
        RECT 7.808 18.528 7.84 21.036 ;
  LAYER M1 ;
        RECT 7.872 18.528 7.904 21.036 ;
  LAYER M1 ;
        RECT 7.936 18.528 7.968 21.036 ;
  LAYER M1 ;
        RECT 8 18.528 8.032 21.036 ;
  LAYER M1 ;
        RECT 8.064 18.528 8.096 21.036 ;
  LAYER M1 ;
        RECT 8.128 18.528 8.16 21.036 ;
  LAYER M1 ;
        RECT 8.192 18.528 8.224 21.036 ;
  LAYER M1 ;
        RECT 8.256 18.528 8.288 21.036 ;
  LAYER M1 ;
        RECT 8.32 18.528 8.352 21.036 ;
  LAYER M1 ;
        RECT 8.384 18.528 8.416 21.036 ;
  LAYER M1 ;
        RECT 8.448 18.528 8.48 21.036 ;
  LAYER M1 ;
        RECT 8.512 18.528 8.544 21.036 ;
  LAYER M1 ;
        RECT 8.576 18.528 8.608 21.036 ;
  LAYER M1 ;
        RECT 8.64 18.528 8.672 21.036 ;
  LAYER M1 ;
        RECT 8.704 18.528 8.736 21.036 ;
  LAYER M1 ;
        RECT 8.768 18.528 8.8 21.036 ;
  LAYER M1 ;
        RECT 8.832 18.528 8.864 21.036 ;
  LAYER M1 ;
        RECT 8.896 18.528 8.928 21.036 ;
  LAYER M1 ;
        RECT 8.96 18.528 8.992 21.036 ;
  LAYER M1 ;
        RECT 9.024 18.528 9.056 21.036 ;
  LAYER M1 ;
        RECT 9.088 18.528 9.12 21.036 ;
  LAYER M1 ;
        RECT 9.152 18.528 9.184 21.036 ;
  LAYER M1 ;
        RECT 9.216 18.528 9.248 21.036 ;
  LAYER M1 ;
        RECT 9.28 18.528 9.312 21.036 ;
  LAYER M1 ;
        RECT 9.344 18.528 9.376 21.036 ;
  LAYER M1 ;
        RECT 9.408 18.528 9.44 21.036 ;
  LAYER M2 ;
        RECT 7.084 18.612 9.556 18.644 ;
  LAYER M2 ;
        RECT 7.084 18.676 9.556 18.708 ;
  LAYER M2 ;
        RECT 7.084 18.74 9.556 18.772 ;
  LAYER M2 ;
        RECT 7.084 18.804 9.556 18.836 ;
  LAYER M2 ;
        RECT 7.084 18.868 9.556 18.9 ;
  LAYER M2 ;
        RECT 7.084 18.932 9.556 18.964 ;
  LAYER M2 ;
        RECT 7.084 18.996 9.556 19.028 ;
  LAYER M2 ;
        RECT 7.084 19.06 9.556 19.092 ;
  LAYER M2 ;
        RECT 7.084 19.124 9.556 19.156 ;
  LAYER M2 ;
        RECT 7.084 19.188 9.556 19.22 ;
  LAYER M2 ;
        RECT 7.084 19.252 9.556 19.284 ;
  LAYER M2 ;
        RECT 7.084 19.316 9.556 19.348 ;
  LAYER M2 ;
        RECT 7.084 19.38 9.556 19.412 ;
  LAYER M2 ;
        RECT 7.084 19.444 9.556 19.476 ;
  LAYER M2 ;
        RECT 7.084 19.508 9.556 19.54 ;
  LAYER M2 ;
        RECT 7.084 19.572 9.556 19.604 ;
  LAYER M2 ;
        RECT 7.084 19.636 9.556 19.668 ;
  LAYER M2 ;
        RECT 7.084 19.7 9.556 19.732 ;
  LAYER M2 ;
        RECT 7.084 19.764 9.556 19.796 ;
  LAYER M2 ;
        RECT 7.084 19.828 9.556 19.86 ;
  LAYER M2 ;
        RECT 7.084 19.892 9.556 19.924 ;
  LAYER M2 ;
        RECT 7.084 19.956 9.556 19.988 ;
  LAYER M2 ;
        RECT 7.084 20.02 9.556 20.052 ;
  LAYER M2 ;
        RECT 7.084 20.084 9.556 20.116 ;
  LAYER M2 ;
        RECT 7.084 20.148 9.556 20.18 ;
  LAYER M2 ;
        RECT 7.084 20.212 9.556 20.244 ;
  LAYER M2 ;
        RECT 7.084 20.276 9.556 20.308 ;
  LAYER M2 ;
        RECT 7.084 20.34 9.556 20.372 ;
  LAYER M2 ;
        RECT 7.084 20.404 9.556 20.436 ;
  LAYER M2 ;
        RECT 7.084 20.468 9.556 20.5 ;
  LAYER M2 ;
        RECT 7.084 20.532 9.556 20.564 ;
  LAYER M2 ;
        RECT 7.084 20.596 9.556 20.628 ;
  LAYER M2 ;
        RECT 7.084 20.66 9.556 20.692 ;
  LAYER M2 ;
        RECT 7.084 20.724 9.556 20.756 ;
  LAYER M2 ;
        RECT 7.084 20.788 9.556 20.82 ;
  LAYER M2 ;
        RECT 7.084 20.852 9.556 20.884 ;
  LAYER M3 ;
        RECT 7.104 18.528 7.136 21.036 ;
  LAYER M3 ;
        RECT 7.168 18.528 7.2 21.036 ;
  LAYER M3 ;
        RECT 7.232 18.528 7.264 21.036 ;
  LAYER M3 ;
        RECT 7.296 18.528 7.328 21.036 ;
  LAYER M3 ;
        RECT 7.36 18.528 7.392 21.036 ;
  LAYER M3 ;
        RECT 7.424 18.528 7.456 21.036 ;
  LAYER M3 ;
        RECT 7.488 18.528 7.52 21.036 ;
  LAYER M3 ;
        RECT 7.552 18.528 7.584 21.036 ;
  LAYER M3 ;
        RECT 7.616 18.528 7.648 21.036 ;
  LAYER M3 ;
        RECT 7.68 18.528 7.712 21.036 ;
  LAYER M3 ;
        RECT 7.744 18.528 7.776 21.036 ;
  LAYER M3 ;
        RECT 7.808 18.528 7.84 21.036 ;
  LAYER M3 ;
        RECT 7.872 18.528 7.904 21.036 ;
  LAYER M3 ;
        RECT 7.936 18.528 7.968 21.036 ;
  LAYER M3 ;
        RECT 8 18.528 8.032 21.036 ;
  LAYER M3 ;
        RECT 8.064 18.528 8.096 21.036 ;
  LAYER M3 ;
        RECT 8.128 18.528 8.16 21.036 ;
  LAYER M3 ;
        RECT 8.192 18.528 8.224 21.036 ;
  LAYER M3 ;
        RECT 8.256 18.528 8.288 21.036 ;
  LAYER M3 ;
        RECT 8.32 18.528 8.352 21.036 ;
  LAYER M3 ;
        RECT 8.384 18.528 8.416 21.036 ;
  LAYER M3 ;
        RECT 8.448 18.528 8.48 21.036 ;
  LAYER M3 ;
        RECT 8.512 18.528 8.544 21.036 ;
  LAYER M3 ;
        RECT 8.576 18.528 8.608 21.036 ;
  LAYER M3 ;
        RECT 8.64 18.528 8.672 21.036 ;
  LAYER M3 ;
        RECT 8.704 18.528 8.736 21.036 ;
  LAYER M3 ;
        RECT 8.768 18.528 8.8 21.036 ;
  LAYER M3 ;
        RECT 8.832 18.528 8.864 21.036 ;
  LAYER M3 ;
        RECT 8.896 18.528 8.928 21.036 ;
  LAYER M3 ;
        RECT 8.96 18.528 8.992 21.036 ;
  LAYER M3 ;
        RECT 9.024 18.528 9.056 21.036 ;
  LAYER M3 ;
        RECT 9.088 18.528 9.12 21.036 ;
  LAYER M3 ;
        RECT 9.152 18.528 9.184 21.036 ;
  LAYER M3 ;
        RECT 9.216 18.528 9.248 21.036 ;
  LAYER M3 ;
        RECT 9.28 18.528 9.312 21.036 ;
  LAYER M3 ;
        RECT 9.344 18.528 9.376 21.036 ;
  LAYER M3 ;
        RECT 9.408 18.528 9.44 21.036 ;
  LAYER M3 ;
        RECT 9.504 18.528 9.536 21.036 ;
  LAYER M1 ;
        RECT 7.119 18.564 7.121 21 ;
  LAYER M1 ;
        RECT 7.199 18.564 7.201 21 ;
  LAYER M1 ;
        RECT 7.279 18.564 7.281 21 ;
  LAYER M1 ;
        RECT 7.359 18.564 7.361 21 ;
  LAYER M1 ;
        RECT 7.439 18.564 7.441 21 ;
  LAYER M1 ;
        RECT 7.519 18.564 7.521 21 ;
  LAYER M1 ;
        RECT 7.599 18.564 7.601 21 ;
  LAYER M1 ;
        RECT 7.679 18.564 7.681 21 ;
  LAYER M1 ;
        RECT 7.759 18.564 7.761 21 ;
  LAYER M1 ;
        RECT 7.839 18.564 7.841 21 ;
  LAYER M1 ;
        RECT 7.919 18.564 7.921 21 ;
  LAYER M1 ;
        RECT 7.999 18.564 8.001 21 ;
  LAYER M1 ;
        RECT 8.079 18.564 8.081 21 ;
  LAYER M1 ;
        RECT 8.159 18.564 8.161 21 ;
  LAYER M1 ;
        RECT 8.239 18.564 8.241 21 ;
  LAYER M1 ;
        RECT 8.319 18.564 8.321 21 ;
  LAYER M1 ;
        RECT 8.399 18.564 8.401 21 ;
  LAYER M1 ;
        RECT 8.479 18.564 8.481 21 ;
  LAYER M1 ;
        RECT 8.559 18.564 8.561 21 ;
  LAYER M1 ;
        RECT 8.639 18.564 8.641 21 ;
  LAYER M1 ;
        RECT 8.719 18.564 8.721 21 ;
  LAYER M1 ;
        RECT 8.799 18.564 8.801 21 ;
  LAYER M1 ;
        RECT 8.879 18.564 8.881 21 ;
  LAYER M1 ;
        RECT 8.959 18.564 8.961 21 ;
  LAYER M1 ;
        RECT 9.039 18.564 9.041 21 ;
  LAYER M1 ;
        RECT 9.119 18.564 9.121 21 ;
  LAYER M1 ;
        RECT 9.199 18.564 9.201 21 ;
  LAYER M1 ;
        RECT 9.279 18.564 9.281 21 ;
  LAYER M1 ;
        RECT 9.359 18.564 9.361 21 ;
  LAYER M1 ;
        RECT 9.439 18.564 9.441 21 ;
  LAYER M2 ;
        RECT 7.12 18.563 9.52 18.565 ;
  LAYER M2 ;
        RECT 7.12 18.647 9.52 18.649 ;
  LAYER M2 ;
        RECT 7.12 18.731 9.52 18.733 ;
  LAYER M2 ;
        RECT 7.12 18.815 9.52 18.817 ;
  LAYER M2 ;
        RECT 7.12 18.899 9.52 18.901 ;
  LAYER M2 ;
        RECT 7.12 18.983 9.52 18.985 ;
  LAYER M2 ;
        RECT 7.12 19.067 9.52 19.069 ;
  LAYER M2 ;
        RECT 7.12 19.151 9.52 19.153 ;
  LAYER M2 ;
        RECT 7.12 19.235 9.52 19.237 ;
  LAYER M2 ;
        RECT 7.12 19.319 9.52 19.321 ;
  LAYER M2 ;
        RECT 7.12 19.403 9.52 19.405 ;
  LAYER M2 ;
        RECT 7.12 19.487 9.52 19.489 ;
  LAYER M2 ;
        RECT 7.12 19.5705 9.52 19.5725 ;
  LAYER M2 ;
        RECT 7.12 19.655 9.52 19.657 ;
  LAYER M2 ;
        RECT 7.12 19.739 9.52 19.741 ;
  LAYER M2 ;
        RECT 7.12 19.823 9.52 19.825 ;
  LAYER M2 ;
        RECT 7.12 19.907 9.52 19.909 ;
  LAYER M2 ;
        RECT 7.12 19.991 9.52 19.993 ;
  LAYER M2 ;
        RECT 7.12 20.075 9.52 20.077 ;
  LAYER M2 ;
        RECT 7.12 20.159 9.52 20.161 ;
  LAYER M2 ;
        RECT 7.12 20.243 9.52 20.245 ;
  LAYER M2 ;
        RECT 7.12 20.327 9.52 20.329 ;
  LAYER M2 ;
        RECT 7.12 20.411 9.52 20.413 ;
  LAYER M2 ;
        RECT 7.12 20.495 9.52 20.497 ;
  LAYER M2 ;
        RECT 7.12 20.579 9.52 20.581 ;
  LAYER M2 ;
        RECT 7.12 20.663 9.52 20.665 ;
  LAYER M2 ;
        RECT 7.12 20.747 9.52 20.749 ;
  LAYER M2 ;
        RECT 7.12 20.831 9.52 20.833 ;
  LAYER M2 ;
        RECT 7.12 20.915 9.52 20.917 ;
  LAYER M1 ;
        RECT 7.104 21.468 7.136 23.976 ;
  LAYER M1 ;
        RECT 7.168 21.468 7.2 23.976 ;
  LAYER M1 ;
        RECT 7.232 21.468 7.264 23.976 ;
  LAYER M1 ;
        RECT 7.296 21.468 7.328 23.976 ;
  LAYER M1 ;
        RECT 7.36 21.468 7.392 23.976 ;
  LAYER M1 ;
        RECT 7.424 21.468 7.456 23.976 ;
  LAYER M1 ;
        RECT 7.488 21.468 7.52 23.976 ;
  LAYER M1 ;
        RECT 7.552 21.468 7.584 23.976 ;
  LAYER M1 ;
        RECT 7.616 21.468 7.648 23.976 ;
  LAYER M1 ;
        RECT 7.68 21.468 7.712 23.976 ;
  LAYER M1 ;
        RECT 7.744 21.468 7.776 23.976 ;
  LAYER M1 ;
        RECT 7.808 21.468 7.84 23.976 ;
  LAYER M1 ;
        RECT 7.872 21.468 7.904 23.976 ;
  LAYER M1 ;
        RECT 7.936 21.468 7.968 23.976 ;
  LAYER M1 ;
        RECT 8 21.468 8.032 23.976 ;
  LAYER M1 ;
        RECT 8.064 21.468 8.096 23.976 ;
  LAYER M1 ;
        RECT 8.128 21.468 8.16 23.976 ;
  LAYER M1 ;
        RECT 8.192 21.468 8.224 23.976 ;
  LAYER M1 ;
        RECT 8.256 21.468 8.288 23.976 ;
  LAYER M1 ;
        RECT 8.32 21.468 8.352 23.976 ;
  LAYER M1 ;
        RECT 8.384 21.468 8.416 23.976 ;
  LAYER M1 ;
        RECT 8.448 21.468 8.48 23.976 ;
  LAYER M1 ;
        RECT 8.512 21.468 8.544 23.976 ;
  LAYER M1 ;
        RECT 8.576 21.468 8.608 23.976 ;
  LAYER M1 ;
        RECT 8.64 21.468 8.672 23.976 ;
  LAYER M1 ;
        RECT 8.704 21.468 8.736 23.976 ;
  LAYER M1 ;
        RECT 8.768 21.468 8.8 23.976 ;
  LAYER M1 ;
        RECT 8.832 21.468 8.864 23.976 ;
  LAYER M1 ;
        RECT 8.896 21.468 8.928 23.976 ;
  LAYER M1 ;
        RECT 8.96 21.468 8.992 23.976 ;
  LAYER M1 ;
        RECT 9.024 21.468 9.056 23.976 ;
  LAYER M1 ;
        RECT 9.088 21.468 9.12 23.976 ;
  LAYER M1 ;
        RECT 9.152 21.468 9.184 23.976 ;
  LAYER M1 ;
        RECT 9.216 21.468 9.248 23.976 ;
  LAYER M1 ;
        RECT 9.28 21.468 9.312 23.976 ;
  LAYER M1 ;
        RECT 9.344 21.468 9.376 23.976 ;
  LAYER M1 ;
        RECT 9.408 21.468 9.44 23.976 ;
  LAYER M2 ;
        RECT 7.084 21.552 9.556 21.584 ;
  LAYER M2 ;
        RECT 7.084 21.616 9.556 21.648 ;
  LAYER M2 ;
        RECT 7.084 21.68 9.556 21.712 ;
  LAYER M2 ;
        RECT 7.084 21.744 9.556 21.776 ;
  LAYER M2 ;
        RECT 7.084 21.808 9.556 21.84 ;
  LAYER M2 ;
        RECT 7.084 21.872 9.556 21.904 ;
  LAYER M2 ;
        RECT 7.084 21.936 9.556 21.968 ;
  LAYER M2 ;
        RECT 7.084 22 9.556 22.032 ;
  LAYER M2 ;
        RECT 7.084 22.064 9.556 22.096 ;
  LAYER M2 ;
        RECT 7.084 22.128 9.556 22.16 ;
  LAYER M2 ;
        RECT 7.084 22.192 9.556 22.224 ;
  LAYER M2 ;
        RECT 7.084 22.256 9.556 22.288 ;
  LAYER M2 ;
        RECT 7.084 22.32 9.556 22.352 ;
  LAYER M2 ;
        RECT 7.084 22.384 9.556 22.416 ;
  LAYER M2 ;
        RECT 7.084 22.448 9.556 22.48 ;
  LAYER M2 ;
        RECT 7.084 22.512 9.556 22.544 ;
  LAYER M2 ;
        RECT 7.084 22.576 9.556 22.608 ;
  LAYER M2 ;
        RECT 7.084 22.64 9.556 22.672 ;
  LAYER M2 ;
        RECT 7.084 22.704 9.556 22.736 ;
  LAYER M2 ;
        RECT 7.084 22.768 9.556 22.8 ;
  LAYER M2 ;
        RECT 7.084 22.832 9.556 22.864 ;
  LAYER M2 ;
        RECT 7.084 22.896 9.556 22.928 ;
  LAYER M2 ;
        RECT 7.084 22.96 9.556 22.992 ;
  LAYER M2 ;
        RECT 7.084 23.024 9.556 23.056 ;
  LAYER M2 ;
        RECT 7.084 23.088 9.556 23.12 ;
  LAYER M2 ;
        RECT 7.084 23.152 9.556 23.184 ;
  LAYER M2 ;
        RECT 7.084 23.216 9.556 23.248 ;
  LAYER M2 ;
        RECT 7.084 23.28 9.556 23.312 ;
  LAYER M2 ;
        RECT 7.084 23.344 9.556 23.376 ;
  LAYER M2 ;
        RECT 7.084 23.408 9.556 23.44 ;
  LAYER M2 ;
        RECT 7.084 23.472 9.556 23.504 ;
  LAYER M2 ;
        RECT 7.084 23.536 9.556 23.568 ;
  LAYER M2 ;
        RECT 7.084 23.6 9.556 23.632 ;
  LAYER M2 ;
        RECT 7.084 23.664 9.556 23.696 ;
  LAYER M2 ;
        RECT 7.084 23.728 9.556 23.76 ;
  LAYER M2 ;
        RECT 7.084 23.792 9.556 23.824 ;
  LAYER M3 ;
        RECT 7.104 21.468 7.136 23.976 ;
  LAYER M3 ;
        RECT 7.168 21.468 7.2 23.976 ;
  LAYER M3 ;
        RECT 7.232 21.468 7.264 23.976 ;
  LAYER M3 ;
        RECT 7.296 21.468 7.328 23.976 ;
  LAYER M3 ;
        RECT 7.36 21.468 7.392 23.976 ;
  LAYER M3 ;
        RECT 7.424 21.468 7.456 23.976 ;
  LAYER M3 ;
        RECT 7.488 21.468 7.52 23.976 ;
  LAYER M3 ;
        RECT 7.552 21.468 7.584 23.976 ;
  LAYER M3 ;
        RECT 7.616 21.468 7.648 23.976 ;
  LAYER M3 ;
        RECT 7.68 21.468 7.712 23.976 ;
  LAYER M3 ;
        RECT 7.744 21.468 7.776 23.976 ;
  LAYER M3 ;
        RECT 7.808 21.468 7.84 23.976 ;
  LAYER M3 ;
        RECT 7.872 21.468 7.904 23.976 ;
  LAYER M3 ;
        RECT 7.936 21.468 7.968 23.976 ;
  LAYER M3 ;
        RECT 8 21.468 8.032 23.976 ;
  LAYER M3 ;
        RECT 8.064 21.468 8.096 23.976 ;
  LAYER M3 ;
        RECT 8.128 21.468 8.16 23.976 ;
  LAYER M3 ;
        RECT 8.192 21.468 8.224 23.976 ;
  LAYER M3 ;
        RECT 8.256 21.468 8.288 23.976 ;
  LAYER M3 ;
        RECT 8.32 21.468 8.352 23.976 ;
  LAYER M3 ;
        RECT 8.384 21.468 8.416 23.976 ;
  LAYER M3 ;
        RECT 8.448 21.468 8.48 23.976 ;
  LAYER M3 ;
        RECT 8.512 21.468 8.544 23.976 ;
  LAYER M3 ;
        RECT 8.576 21.468 8.608 23.976 ;
  LAYER M3 ;
        RECT 8.64 21.468 8.672 23.976 ;
  LAYER M3 ;
        RECT 8.704 21.468 8.736 23.976 ;
  LAYER M3 ;
        RECT 8.768 21.468 8.8 23.976 ;
  LAYER M3 ;
        RECT 8.832 21.468 8.864 23.976 ;
  LAYER M3 ;
        RECT 8.896 21.468 8.928 23.976 ;
  LAYER M3 ;
        RECT 8.96 21.468 8.992 23.976 ;
  LAYER M3 ;
        RECT 9.024 21.468 9.056 23.976 ;
  LAYER M3 ;
        RECT 9.088 21.468 9.12 23.976 ;
  LAYER M3 ;
        RECT 9.152 21.468 9.184 23.976 ;
  LAYER M3 ;
        RECT 9.216 21.468 9.248 23.976 ;
  LAYER M3 ;
        RECT 9.28 21.468 9.312 23.976 ;
  LAYER M3 ;
        RECT 9.344 21.468 9.376 23.976 ;
  LAYER M3 ;
        RECT 9.408 21.468 9.44 23.976 ;
  LAYER M3 ;
        RECT 9.504 21.468 9.536 23.976 ;
  LAYER M1 ;
        RECT 7.119 21.504 7.121 23.94 ;
  LAYER M1 ;
        RECT 7.199 21.504 7.201 23.94 ;
  LAYER M1 ;
        RECT 7.279 21.504 7.281 23.94 ;
  LAYER M1 ;
        RECT 7.359 21.504 7.361 23.94 ;
  LAYER M1 ;
        RECT 7.439 21.504 7.441 23.94 ;
  LAYER M1 ;
        RECT 7.519 21.504 7.521 23.94 ;
  LAYER M1 ;
        RECT 7.599 21.504 7.601 23.94 ;
  LAYER M1 ;
        RECT 7.679 21.504 7.681 23.94 ;
  LAYER M1 ;
        RECT 7.759 21.504 7.761 23.94 ;
  LAYER M1 ;
        RECT 7.839 21.504 7.841 23.94 ;
  LAYER M1 ;
        RECT 7.919 21.504 7.921 23.94 ;
  LAYER M1 ;
        RECT 7.999 21.504 8.001 23.94 ;
  LAYER M1 ;
        RECT 8.079 21.504 8.081 23.94 ;
  LAYER M1 ;
        RECT 8.159 21.504 8.161 23.94 ;
  LAYER M1 ;
        RECT 8.239 21.504 8.241 23.94 ;
  LAYER M1 ;
        RECT 8.319 21.504 8.321 23.94 ;
  LAYER M1 ;
        RECT 8.399 21.504 8.401 23.94 ;
  LAYER M1 ;
        RECT 8.479 21.504 8.481 23.94 ;
  LAYER M1 ;
        RECT 8.559 21.504 8.561 23.94 ;
  LAYER M1 ;
        RECT 8.639 21.504 8.641 23.94 ;
  LAYER M1 ;
        RECT 8.719 21.504 8.721 23.94 ;
  LAYER M1 ;
        RECT 8.799 21.504 8.801 23.94 ;
  LAYER M1 ;
        RECT 8.879 21.504 8.881 23.94 ;
  LAYER M1 ;
        RECT 8.959 21.504 8.961 23.94 ;
  LAYER M1 ;
        RECT 9.039 21.504 9.041 23.94 ;
  LAYER M1 ;
        RECT 9.119 21.504 9.121 23.94 ;
  LAYER M1 ;
        RECT 9.199 21.504 9.201 23.94 ;
  LAYER M1 ;
        RECT 9.279 21.504 9.281 23.94 ;
  LAYER M1 ;
        RECT 9.359 21.504 9.361 23.94 ;
  LAYER M1 ;
        RECT 9.439 21.504 9.441 23.94 ;
  LAYER M2 ;
        RECT 7.12 21.503 9.52 21.505 ;
  LAYER M2 ;
        RECT 7.12 21.587 9.52 21.589 ;
  LAYER M2 ;
        RECT 7.12 21.671 9.52 21.673 ;
  LAYER M2 ;
        RECT 7.12 21.755 9.52 21.757 ;
  LAYER M2 ;
        RECT 7.12 21.839 9.52 21.841 ;
  LAYER M2 ;
        RECT 7.12 21.923 9.52 21.925 ;
  LAYER M2 ;
        RECT 7.12 22.007 9.52 22.009 ;
  LAYER M2 ;
        RECT 7.12 22.091 9.52 22.093 ;
  LAYER M2 ;
        RECT 7.12 22.175 9.52 22.177 ;
  LAYER M2 ;
        RECT 7.12 22.259 9.52 22.261 ;
  LAYER M2 ;
        RECT 7.12 22.343 9.52 22.345 ;
  LAYER M2 ;
        RECT 7.12 22.427 9.52 22.429 ;
  LAYER M2 ;
        RECT 7.12 22.5105 9.52 22.5125 ;
  LAYER M2 ;
        RECT 7.12 22.595 9.52 22.597 ;
  LAYER M2 ;
        RECT 7.12 22.679 9.52 22.681 ;
  LAYER M2 ;
        RECT 7.12 22.763 9.52 22.765 ;
  LAYER M2 ;
        RECT 7.12 22.847 9.52 22.849 ;
  LAYER M2 ;
        RECT 7.12 22.931 9.52 22.933 ;
  LAYER M2 ;
        RECT 7.12 23.015 9.52 23.017 ;
  LAYER M2 ;
        RECT 7.12 23.099 9.52 23.101 ;
  LAYER M2 ;
        RECT 7.12 23.183 9.52 23.185 ;
  LAYER M2 ;
        RECT 7.12 23.267 9.52 23.269 ;
  LAYER M2 ;
        RECT 7.12 23.351 9.52 23.353 ;
  LAYER M2 ;
        RECT 7.12 23.435 9.52 23.437 ;
  LAYER M2 ;
        RECT 7.12 23.519 9.52 23.521 ;
  LAYER M2 ;
        RECT 7.12 23.603 9.52 23.605 ;
  LAYER M2 ;
        RECT 7.12 23.687 9.52 23.689 ;
  LAYER M2 ;
        RECT 7.12 23.771 9.52 23.773 ;
  LAYER M2 ;
        RECT 7.12 23.855 9.52 23.857 ;
  END 
END Cap_30fF_Cap_30fF
