MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 17.04 BY 19.992 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.844 19.536 6.876 19.608 ;
      LAYER M2 ;
        RECT 6.824 19.556 6.896 19.588 ;
      LAYER M1 ;
        RECT 10.46 19.536 10.492 19.608 ;
      LAYER M2 ;
        RECT 10.44 19.556 10.512 19.588 ;
      LAYER M2 ;
        RECT 6.86 19.556 10.476 19.588 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.236 0.384 6.268 0.456 ;
      LAYER M2 ;
        RECT 6.216 0.404 6.288 0.436 ;
      LAYER M1 ;
        RECT 9.852 0.384 9.884 0.456 ;
      LAYER M2 ;
        RECT 9.832 0.404 9.904 0.436 ;
      LAYER M2 ;
        RECT 6.252 0.404 9.868 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 7.004 19.704 7.036 19.776 ;
      LAYER M2 ;
        RECT 6.984 19.724 7.056 19.756 ;
      LAYER M1 ;
        RECT 10.62 19.704 10.652 19.776 ;
      LAYER M2 ;
        RECT 10.6 19.724 10.672 19.756 ;
      LAYER M2 ;
        RECT 7.02 19.724 10.636 19.756 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.396 0.216 6.428 0.288 ;
      LAYER M2 ;
        RECT 6.376 0.236 6.448 0.268 ;
      LAYER M1 ;
        RECT 10.012 0.216 10.044 0.288 ;
      LAYER M2 ;
        RECT 9.992 0.236 10.064 0.268 ;
      LAYER M2 ;
        RECT 6.412 0.236 10.028 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 9.692 7.188 9.724 7.26 ;
  LAYER M2 ;
        RECT 9.672 7.208 9.744 7.24 ;
  LAYER M2 ;
        RECT 6.252 7.208 9.708 7.24 ;
  LAYER M1 ;
        RECT 6.236 7.188 6.268 7.26 ;
  LAYER M2 ;
        RECT 6.216 7.208 6.288 7.24 ;
  LAYER M1 ;
        RECT 6.076 13.404 6.108 13.476 ;
  LAYER M2 ;
        RECT 6.056 13.424 6.128 13.456 ;
  LAYER M1 ;
        RECT 6.076 13.272 6.108 13.44 ;
  LAYER M1 ;
        RECT 6.076 13.236 6.108 13.308 ;
  LAYER M2 ;
        RECT 6.056 13.256 6.128 13.288 ;
  LAYER M2 ;
        RECT 6.092 13.256 6.252 13.288 ;
  LAYER M1 ;
        RECT 6.236 13.236 6.268 13.308 ;
  LAYER M2 ;
        RECT 6.216 13.256 6.288 13.288 ;
  LAYER M1 ;
        RECT 6.236 0.384 6.268 0.456 ;
  LAYER M2 ;
        RECT 6.216 0.404 6.288 0.436 ;
  LAYER M1 ;
        RECT 6.236 0.42 6.268 0.672 ;
  LAYER M1 ;
        RECT 6.236 0.672 6.268 13.272 ;
  LAYER M1 ;
        RECT 13.308 4.08 13.34 4.152 ;
  LAYER M2 ;
        RECT 13.288 4.1 13.36 4.132 ;
  LAYER M2 ;
        RECT 9.868 4.1 13.324 4.132 ;
  LAYER M1 ;
        RECT 9.852 4.08 9.884 4.152 ;
  LAYER M2 ;
        RECT 9.832 4.1 9.904 4.132 ;
  LAYER M1 ;
        RECT 9.852 0.384 9.884 0.456 ;
  LAYER M2 ;
        RECT 9.832 0.404 9.904 0.436 ;
  LAYER M1 ;
        RECT 9.852 0.42 9.884 0.672 ;
  LAYER M1 ;
        RECT 9.852 0.672 9.884 4.116 ;
  LAYER M2 ;
        RECT 6.252 0.404 9.868 0.436 ;
  LAYER M1 ;
        RECT 6.076 7.188 6.108 7.26 ;
  LAYER M2 ;
        RECT 6.056 7.208 6.128 7.24 ;
  LAYER M1 ;
        RECT 6.076 7.056 6.108 7.224 ;
  LAYER M1 ;
        RECT 6.076 7.02 6.108 7.092 ;
  LAYER M2 ;
        RECT 6.056 7.04 6.128 7.072 ;
  LAYER M2 ;
        RECT 6.092 7.04 6.412 7.072 ;
  LAYER M1 ;
        RECT 6.396 7.02 6.428 7.092 ;
  LAYER M2 ;
        RECT 6.376 7.04 6.448 7.072 ;
  LAYER M1 ;
        RECT 6.076 10.296 6.108 10.368 ;
  LAYER M2 ;
        RECT 6.056 10.316 6.128 10.348 ;
  LAYER M1 ;
        RECT 6.076 10.164 6.108 10.332 ;
  LAYER M1 ;
        RECT 6.076 10.128 6.108 10.2 ;
  LAYER M2 ;
        RECT 6.056 10.148 6.128 10.18 ;
  LAYER M2 ;
        RECT 6.092 10.148 6.412 10.18 ;
  LAYER M1 ;
        RECT 6.396 10.128 6.428 10.2 ;
  LAYER M2 ;
        RECT 6.376 10.148 6.448 10.18 ;
  LAYER M1 ;
        RECT 9.692 4.08 9.724 4.152 ;
  LAYER M2 ;
        RECT 9.672 4.1 9.744 4.132 ;
  LAYER M2 ;
        RECT 6.412 4.1 9.708 4.132 ;
  LAYER M1 ;
        RECT 6.396 4.08 6.428 4.152 ;
  LAYER M2 ;
        RECT 6.376 4.1 6.448 4.132 ;
  LAYER M1 ;
        RECT 9.692 13.404 9.724 13.476 ;
  LAYER M2 ;
        RECT 9.672 13.424 9.744 13.456 ;
  LAYER M2 ;
        RECT 6.412 13.424 9.708 13.456 ;
  LAYER M1 ;
        RECT 6.396 13.404 6.428 13.476 ;
  LAYER M2 ;
        RECT 6.376 13.424 6.448 13.456 ;
  LAYER M1 ;
        RECT 6.396 0.216 6.428 0.288 ;
  LAYER M2 ;
        RECT 6.376 0.236 6.448 0.268 ;
  LAYER M1 ;
        RECT 6.396 0.252 6.428 0.672 ;
  LAYER M1 ;
        RECT 6.396 0.672 6.428 13.44 ;
  LAYER M1 ;
        RECT 13.308 10.296 13.34 10.368 ;
  LAYER M2 ;
        RECT 13.288 10.316 13.36 10.348 ;
  LAYER M2 ;
        RECT 10.028 10.316 13.324 10.348 ;
  LAYER M1 ;
        RECT 10.012 10.296 10.044 10.368 ;
  LAYER M2 ;
        RECT 9.992 10.316 10.064 10.348 ;
  LAYER M1 ;
        RECT 13.308 7.188 13.34 7.26 ;
  LAYER M2 ;
        RECT 13.288 7.208 13.36 7.24 ;
  LAYER M2 ;
        RECT 10.028 7.208 13.324 7.24 ;
  LAYER M1 ;
        RECT 10.012 7.188 10.044 7.26 ;
  LAYER M2 ;
        RECT 9.992 7.208 10.064 7.24 ;
  LAYER M1 ;
        RECT 10.012 0.216 10.044 0.288 ;
  LAYER M2 ;
        RECT 9.992 0.236 10.064 0.268 ;
  LAYER M1 ;
        RECT 10.012 0.252 10.044 0.672 ;
  LAYER M1 ;
        RECT 10.012 0.672 10.044 10.332 ;
  LAYER M2 ;
        RECT 6.412 0.236 10.028 0.268 ;
  LAYER M1 ;
        RECT 6.076 0.972 6.108 1.044 ;
  LAYER M2 ;
        RECT 6.056 0.992 6.128 1.024 ;
  LAYER M1 ;
        RECT 6.076 0.84 6.108 1.008 ;
  LAYER M1 ;
        RECT 6.076 0.804 6.108 0.876 ;
  LAYER M2 ;
        RECT 6.056 0.824 6.128 0.856 ;
  LAYER M2 ;
        RECT 6.092 0.824 6.572 0.856 ;
  LAYER M1 ;
        RECT 6.556 0.804 6.588 0.876 ;
  LAYER M2 ;
        RECT 6.536 0.824 6.608 0.856 ;
  LAYER M1 ;
        RECT 6.076 4.08 6.108 4.152 ;
  LAYER M2 ;
        RECT 6.056 4.1 6.128 4.132 ;
  LAYER M1 ;
        RECT 6.076 3.948 6.108 4.116 ;
  LAYER M1 ;
        RECT 6.076 3.912 6.108 3.984 ;
  LAYER M2 ;
        RECT 6.056 3.932 6.128 3.964 ;
  LAYER M2 ;
        RECT 6.092 3.932 6.572 3.964 ;
  LAYER M1 ;
        RECT 6.556 3.912 6.588 3.984 ;
  LAYER M2 ;
        RECT 6.536 3.932 6.608 3.964 ;
  LAYER M1 ;
        RECT 6.076 16.512 6.108 16.584 ;
  LAYER M2 ;
        RECT 6.056 16.532 6.128 16.564 ;
  LAYER M1 ;
        RECT 6.076 16.38 6.108 16.548 ;
  LAYER M1 ;
        RECT 6.076 16.344 6.108 16.416 ;
  LAYER M2 ;
        RECT 6.056 16.364 6.128 16.396 ;
  LAYER M2 ;
        RECT 6.092 16.364 6.572 16.396 ;
  LAYER M1 ;
        RECT 6.556 16.344 6.588 16.416 ;
  LAYER M2 ;
        RECT 6.536 16.364 6.608 16.396 ;
  LAYER M1 ;
        RECT 9.692 0.972 9.724 1.044 ;
  LAYER M2 ;
        RECT 9.672 0.992 9.744 1.024 ;
  LAYER M2 ;
        RECT 6.572 0.992 9.708 1.024 ;
  LAYER M1 ;
        RECT 6.556 0.972 6.588 1.044 ;
  LAYER M2 ;
        RECT 6.536 0.992 6.608 1.024 ;
  LAYER M1 ;
        RECT 9.692 10.296 9.724 10.368 ;
  LAYER M2 ;
        RECT 9.672 10.316 9.744 10.348 ;
  LAYER M2 ;
        RECT 6.572 10.316 9.708 10.348 ;
  LAYER M1 ;
        RECT 6.556 10.296 6.588 10.368 ;
  LAYER M2 ;
        RECT 6.536 10.316 6.608 10.348 ;
  LAYER M1 ;
        RECT 9.692 16.512 9.724 16.584 ;
  LAYER M2 ;
        RECT 9.672 16.532 9.744 16.564 ;
  LAYER M2 ;
        RECT 6.572 16.532 9.708 16.564 ;
  LAYER M1 ;
        RECT 6.556 16.512 6.588 16.584 ;
  LAYER M2 ;
        RECT 6.536 16.532 6.608 16.564 ;
  LAYER M1 ;
        RECT 6.556 0.048 6.588 0.12 ;
  LAYER M2 ;
        RECT 6.536 0.068 6.608 0.1 ;
  LAYER M1 ;
        RECT 6.556 0.084 6.588 0.672 ;
  LAYER M1 ;
        RECT 6.556 0.672 6.588 16.548 ;
  LAYER M1 ;
        RECT 13.308 0.972 13.34 1.044 ;
  LAYER M2 ;
        RECT 13.288 0.992 13.36 1.024 ;
  LAYER M2 ;
        RECT 10.188 0.992 13.324 1.024 ;
  LAYER M1 ;
        RECT 10.172 0.972 10.204 1.044 ;
  LAYER M2 ;
        RECT 10.152 0.992 10.224 1.024 ;
  LAYER M1 ;
        RECT 13.308 13.404 13.34 13.476 ;
  LAYER M2 ;
        RECT 13.288 13.424 13.36 13.456 ;
  LAYER M2 ;
        RECT 10.188 13.424 13.324 13.456 ;
  LAYER M1 ;
        RECT 10.172 13.404 10.204 13.476 ;
  LAYER M2 ;
        RECT 10.152 13.424 10.224 13.456 ;
  LAYER M1 ;
        RECT 13.308 16.512 13.34 16.584 ;
  LAYER M2 ;
        RECT 13.288 16.532 13.36 16.564 ;
  LAYER M2 ;
        RECT 10.188 16.532 13.324 16.564 ;
  LAYER M1 ;
        RECT 10.172 16.512 10.204 16.584 ;
  LAYER M2 ;
        RECT 10.152 16.532 10.224 16.564 ;
  LAYER M1 ;
        RECT 10.172 0.048 10.204 0.12 ;
  LAYER M2 ;
        RECT 10.152 0.068 10.224 0.1 ;
  LAYER M1 ;
        RECT 10.172 0.084 10.204 0.672 ;
  LAYER M1 ;
        RECT 10.172 0.672 10.204 16.548 ;
  LAYER M2 ;
        RECT 6.572 0.068 10.188 0.1 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M2 ;
        RECT 2.476 16.532 6.092 16.564 ;
  LAYER M1 ;
        RECT 6.076 16.512 6.108 16.584 ;
  LAYER M2 ;
        RECT 6.056 16.532 6.128 16.564 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 13.44 2.492 16.548 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 10.332 2.492 13.44 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 7.224 2.492 10.332 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 2.46 4.116 2.492 7.224 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 1.044 ;
  LAYER M2 ;
        RECT 2.44 0.992 2.512 1.024 ;
  LAYER M1 ;
        RECT 2.46 1.008 2.492 4.116 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 16.924 16.512 16.956 16.584 ;
  LAYER M2 ;
        RECT 16.904 16.532 16.976 16.564 ;
  LAYER M2 ;
        RECT 13.324 16.532 16.94 16.564 ;
  LAYER M1 ;
        RECT 13.308 16.512 13.34 16.584 ;
  LAYER M2 ;
        RECT 13.288 16.532 13.36 16.564 ;
  LAYER M1 ;
        RECT 16.924 13.404 16.956 13.476 ;
  LAYER M2 ;
        RECT 16.904 13.424 16.976 13.456 ;
  LAYER M2 ;
        RECT 13.324 13.424 16.94 13.456 ;
  LAYER M1 ;
        RECT 13.308 13.404 13.34 13.476 ;
  LAYER M2 ;
        RECT 13.288 13.424 13.36 13.456 ;
  LAYER M1 ;
        RECT 16.924 10.296 16.956 10.368 ;
  LAYER M2 ;
        RECT 16.904 10.316 16.976 10.348 ;
  LAYER M1 ;
        RECT 16.924 10.332 16.956 13.44 ;
  LAYER M1 ;
        RECT 16.924 13.404 16.956 13.476 ;
  LAYER M2 ;
        RECT 16.904 13.424 16.976 13.456 ;
  LAYER M1 ;
        RECT 16.924 7.188 16.956 7.26 ;
  LAYER M2 ;
        RECT 16.904 7.208 16.976 7.24 ;
  LAYER M1 ;
        RECT 16.924 7.224 16.956 10.332 ;
  LAYER M1 ;
        RECT 16.924 10.296 16.956 10.368 ;
  LAYER M2 ;
        RECT 16.904 10.316 16.976 10.348 ;
  LAYER M1 ;
        RECT 16.924 4.08 16.956 4.152 ;
  LAYER M2 ;
        RECT 16.904 4.1 16.976 4.132 ;
  LAYER M1 ;
        RECT 16.924 4.116 16.956 7.224 ;
  LAYER M1 ;
        RECT 16.924 7.188 16.956 7.26 ;
  LAYER M2 ;
        RECT 16.904 7.208 16.976 7.24 ;
  LAYER M1 ;
        RECT 16.924 0.972 16.956 1.044 ;
  LAYER M2 ;
        RECT 16.904 0.992 16.976 1.024 ;
  LAYER M1 ;
        RECT 16.924 1.008 16.956 4.116 ;
  LAYER M1 ;
        RECT 16.924 4.08 16.956 4.152 ;
  LAYER M2 ;
        RECT 16.904 4.1 16.976 4.132 ;
  LAYER M1 ;
        RECT 7.324 9.624 7.356 9.696 ;
  LAYER M2 ;
        RECT 7.304 9.644 7.376 9.676 ;
  LAYER M2 ;
        RECT 6.86 9.644 7.34 9.676 ;
  LAYER M1 ;
        RECT 6.844 9.624 6.876 9.696 ;
  LAYER M2 ;
        RECT 6.824 9.644 6.896 9.676 ;
  LAYER M1 ;
        RECT 3.708 15.84 3.74 15.912 ;
  LAYER M2 ;
        RECT 3.688 15.86 3.76 15.892 ;
  LAYER M1 ;
        RECT 3.708 15.876 3.74 16.044 ;
  LAYER M1 ;
        RECT 3.708 16.008 3.74 16.08 ;
  LAYER M2 ;
        RECT 3.688 16.028 3.76 16.06 ;
  LAYER M2 ;
        RECT 3.724 16.028 6.86 16.06 ;
  LAYER M1 ;
        RECT 6.844 16.008 6.876 16.08 ;
  LAYER M2 ;
        RECT 6.824 16.028 6.896 16.06 ;
  LAYER M1 ;
        RECT 6.844 19.536 6.876 19.608 ;
  LAYER M2 ;
        RECT 6.824 19.556 6.896 19.588 ;
  LAYER M1 ;
        RECT 6.844 19.32 6.876 19.572 ;
  LAYER M1 ;
        RECT 6.844 9.66 6.876 19.32 ;
  LAYER M1 ;
        RECT 10.94 6.516 10.972 6.588 ;
  LAYER M2 ;
        RECT 10.92 6.536 10.992 6.568 ;
  LAYER M2 ;
        RECT 10.476 6.536 10.956 6.568 ;
  LAYER M1 ;
        RECT 10.46 6.516 10.492 6.588 ;
  LAYER M2 ;
        RECT 10.44 6.536 10.512 6.568 ;
  LAYER M1 ;
        RECT 10.46 19.536 10.492 19.608 ;
  LAYER M2 ;
        RECT 10.44 19.556 10.512 19.588 ;
  LAYER M1 ;
        RECT 10.46 19.32 10.492 19.572 ;
  LAYER M1 ;
        RECT 10.46 6.552 10.492 19.32 ;
  LAYER M2 ;
        RECT 6.86 19.556 10.476 19.588 ;
  LAYER M1 ;
        RECT 3.708 9.624 3.74 9.696 ;
  LAYER M2 ;
        RECT 3.688 9.644 3.76 9.676 ;
  LAYER M1 ;
        RECT 3.708 9.66 3.74 9.828 ;
  LAYER M1 ;
        RECT 3.708 9.792 3.74 9.864 ;
  LAYER M2 ;
        RECT 3.688 9.812 3.76 9.844 ;
  LAYER M2 ;
        RECT 3.724 9.812 7.02 9.844 ;
  LAYER M1 ;
        RECT 7.004 9.792 7.036 9.864 ;
  LAYER M2 ;
        RECT 6.984 9.812 7.056 9.844 ;
  LAYER M1 ;
        RECT 3.708 12.732 3.74 12.804 ;
  LAYER M2 ;
        RECT 3.688 12.752 3.76 12.784 ;
  LAYER M1 ;
        RECT 3.708 12.768 3.74 12.936 ;
  LAYER M1 ;
        RECT 3.708 12.9 3.74 12.972 ;
  LAYER M2 ;
        RECT 3.688 12.92 3.76 12.952 ;
  LAYER M2 ;
        RECT 3.724 12.92 7.02 12.952 ;
  LAYER M1 ;
        RECT 7.004 12.9 7.036 12.972 ;
  LAYER M2 ;
        RECT 6.984 12.92 7.056 12.952 ;
  LAYER M1 ;
        RECT 7.324 6.516 7.356 6.588 ;
  LAYER M2 ;
        RECT 7.304 6.536 7.376 6.568 ;
  LAYER M2 ;
        RECT 7.02 6.536 7.34 6.568 ;
  LAYER M1 ;
        RECT 7.004 6.516 7.036 6.588 ;
  LAYER M2 ;
        RECT 6.984 6.536 7.056 6.568 ;
  LAYER M1 ;
        RECT 7.324 15.84 7.356 15.912 ;
  LAYER M2 ;
        RECT 7.304 15.86 7.376 15.892 ;
  LAYER M2 ;
        RECT 7.02 15.86 7.34 15.892 ;
  LAYER M1 ;
        RECT 7.004 15.84 7.036 15.912 ;
  LAYER M2 ;
        RECT 6.984 15.86 7.056 15.892 ;
  LAYER M1 ;
        RECT 7.004 19.704 7.036 19.776 ;
  LAYER M2 ;
        RECT 6.984 19.724 7.056 19.756 ;
  LAYER M1 ;
        RECT 7.004 19.32 7.036 19.74 ;
  LAYER M1 ;
        RECT 7.004 6.552 7.036 19.32 ;
  LAYER M1 ;
        RECT 10.94 12.732 10.972 12.804 ;
  LAYER M2 ;
        RECT 10.92 12.752 10.992 12.784 ;
  LAYER M2 ;
        RECT 10.636 12.752 10.956 12.784 ;
  LAYER M1 ;
        RECT 10.62 12.732 10.652 12.804 ;
  LAYER M2 ;
        RECT 10.6 12.752 10.672 12.784 ;
  LAYER M1 ;
        RECT 10.94 9.624 10.972 9.696 ;
  LAYER M2 ;
        RECT 10.92 9.644 10.992 9.676 ;
  LAYER M2 ;
        RECT 10.636 9.644 10.956 9.676 ;
  LAYER M1 ;
        RECT 10.62 9.624 10.652 9.696 ;
  LAYER M2 ;
        RECT 10.6 9.644 10.672 9.676 ;
  LAYER M1 ;
        RECT 10.62 19.704 10.652 19.776 ;
  LAYER M2 ;
        RECT 10.6 19.724 10.672 19.756 ;
  LAYER M1 ;
        RECT 10.62 19.32 10.652 19.74 ;
  LAYER M1 ;
        RECT 10.62 9.66 10.652 19.32 ;
  LAYER M2 ;
        RECT 7.02 19.724 10.636 19.756 ;
  LAYER M1 ;
        RECT 3.708 3.408 3.74 3.48 ;
  LAYER M2 ;
        RECT 3.688 3.428 3.76 3.46 ;
  LAYER M1 ;
        RECT 3.708 3.444 3.74 3.612 ;
  LAYER M1 ;
        RECT 3.708 3.576 3.74 3.648 ;
  LAYER M2 ;
        RECT 3.688 3.596 3.76 3.628 ;
  LAYER M2 ;
        RECT 3.724 3.596 7.18 3.628 ;
  LAYER M1 ;
        RECT 7.164 3.576 7.196 3.648 ;
  LAYER M2 ;
        RECT 7.144 3.596 7.216 3.628 ;
  LAYER M1 ;
        RECT 3.708 6.516 3.74 6.588 ;
  LAYER M2 ;
        RECT 3.688 6.536 3.76 6.568 ;
  LAYER M1 ;
        RECT 3.708 6.552 3.74 6.72 ;
  LAYER M1 ;
        RECT 3.708 6.684 3.74 6.756 ;
  LAYER M2 ;
        RECT 3.688 6.704 3.76 6.736 ;
  LAYER M2 ;
        RECT 3.724 6.704 7.18 6.736 ;
  LAYER M1 ;
        RECT 7.164 6.684 7.196 6.756 ;
  LAYER M2 ;
        RECT 7.144 6.704 7.216 6.736 ;
  LAYER M1 ;
        RECT 3.708 18.948 3.74 19.02 ;
  LAYER M2 ;
        RECT 3.688 18.968 3.76 19 ;
  LAYER M1 ;
        RECT 3.708 18.984 3.74 19.152 ;
  LAYER M1 ;
        RECT 3.708 19.116 3.74 19.188 ;
  LAYER M2 ;
        RECT 3.688 19.136 3.76 19.168 ;
  LAYER M2 ;
        RECT 3.724 19.136 7.18 19.168 ;
  LAYER M1 ;
        RECT 7.164 19.116 7.196 19.188 ;
  LAYER M2 ;
        RECT 7.144 19.136 7.216 19.168 ;
  LAYER M1 ;
        RECT 7.324 3.408 7.356 3.48 ;
  LAYER M2 ;
        RECT 7.304 3.428 7.376 3.46 ;
  LAYER M2 ;
        RECT 7.18 3.428 7.34 3.46 ;
  LAYER M1 ;
        RECT 7.164 3.408 7.196 3.48 ;
  LAYER M2 ;
        RECT 7.144 3.428 7.216 3.46 ;
  LAYER M1 ;
        RECT 7.324 12.732 7.356 12.804 ;
  LAYER M2 ;
        RECT 7.304 12.752 7.376 12.784 ;
  LAYER M2 ;
        RECT 7.18 12.752 7.34 12.784 ;
  LAYER M1 ;
        RECT 7.164 12.732 7.196 12.804 ;
  LAYER M2 ;
        RECT 7.144 12.752 7.216 12.784 ;
  LAYER M1 ;
        RECT 7.324 18.948 7.356 19.02 ;
  LAYER M2 ;
        RECT 7.304 18.968 7.376 19 ;
  LAYER M2 ;
        RECT 7.18 18.968 7.34 19 ;
  LAYER M1 ;
        RECT 7.164 18.948 7.196 19.02 ;
  LAYER M2 ;
        RECT 7.144 18.968 7.216 19 ;
  LAYER M1 ;
        RECT 7.164 19.872 7.196 19.944 ;
  LAYER M2 ;
        RECT 7.144 19.892 7.216 19.924 ;
  LAYER M1 ;
        RECT 7.164 19.32 7.196 19.908 ;
  LAYER M1 ;
        RECT 7.164 3.444 7.196 19.32 ;
  LAYER M1 ;
        RECT 10.94 3.408 10.972 3.48 ;
  LAYER M2 ;
        RECT 10.92 3.428 10.992 3.46 ;
  LAYER M2 ;
        RECT 10.796 3.428 10.956 3.46 ;
  LAYER M1 ;
        RECT 10.78 3.408 10.812 3.48 ;
  LAYER M2 ;
        RECT 10.76 3.428 10.832 3.46 ;
  LAYER M1 ;
        RECT 10.94 15.84 10.972 15.912 ;
  LAYER M2 ;
        RECT 10.92 15.86 10.992 15.892 ;
  LAYER M2 ;
        RECT 10.796 15.86 10.956 15.892 ;
  LAYER M1 ;
        RECT 10.78 15.84 10.812 15.912 ;
  LAYER M2 ;
        RECT 10.76 15.86 10.832 15.892 ;
  LAYER M1 ;
        RECT 10.94 18.948 10.972 19.02 ;
  LAYER M2 ;
        RECT 10.92 18.968 10.992 19 ;
  LAYER M2 ;
        RECT 10.796 18.968 10.956 19 ;
  LAYER M1 ;
        RECT 10.78 18.948 10.812 19.02 ;
  LAYER M2 ;
        RECT 10.76 18.968 10.832 19 ;
  LAYER M1 ;
        RECT 10.78 19.872 10.812 19.944 ;
  LAYER M2 ;
        RECT 10.76 19.892 10.832 19.924 ;
  LAYER M1 ;
        RECT 10.78 19.32 10.812 19.908 ;
  LAYER M1 ;
        RECT 10.78 3.444 10.812 19.32 ;
  LAYER M2 ;
        RECT 7.18 19.892 10.796 19.924 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M2 ;
        RECT 0.108 18.968 3.724 19 ;
  LAYER M1 ;
        RECT 3.708 18.948 3.74 19.02 ;
  LAYER M2 ;
        RECT 3.688 18.968 3.76 19 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 15.876 0.124 18.984 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 12.768 0.124 15.876 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 9.66 0.124 12.768 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 0.092 6.552 0.124 9.66 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 3.408 0.124 3.48 ;
  LAYER M2 ;
        RECT 0.072 3.428 0.144 3.46 ;
  LAYER M1 ;
        RECT 0.092 3.444 0.124 6.552 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 14.556 18.948 14.588 19.02 ;
  LAYER M2 ;
        RECT 14.536 18.968 14.608 19 ;
  LAYER M2 ;
        RECT 10.956 18.968 14.572 19 ;
  LAYER M1 ;
        RECT 10.94 18.948 10.972 19.02 ;
  LAYER M2 ;
        RECT 10.92 18.968 10.992 19 ;
  LAYER M1 ;
        RECT 14.556 15.84 14.588 15.912 ;
  LAYER M2 ;
        RECT 14.536 15.86 14.608 15.892 ;
  LAYER M2 ;
        RECT 10.956 15.86 14.572 15.892 ;
  LAYER M1 ;
        RECT 10.94 15.84 10.972 15.912 ;
  LAYER M2 ;
        RECT 10.92 15.86 10.992 15.892 ;
  LAYER M1 ;
        RECT 14.556 12.732 14.588 12.804 ;
  LAYER M2 ;
        RECT 14.536 12.752 14.608 12.784 ;
  LAYER M1 ;
        RECT 14.556 12.768 14.588 15.876 ;
  LAYER M1 ;
        RECT 14.556 15.84 14.588 15.912 ;
  LAYER M2 ;
        RECT 14.536 15.86 14.608 15.892 ;
  LAYER M1 ;
        RECT 14.556 9.624 14.588 9.696 ;
  LAYER M2 ;
        RECT 14.536 9.644 14.608 9.676 ;
  LAYER M1 ;
        RECT 14.556 9.66 14.588 12.768 ;
  LAYER M1 ;
        RECT 14.556 12.732 14.588 12.804 ;
  LAYER M2 ;
        RECT 14.536 12.752 14.608 12.784 ;
  LAYER M1 ;
        RECT 14.556 6.516 14.588 6.588 ;
  LAYER M2 ;
        RECT 14.536 6.536 14.608 6.568 ;
  LAYER M1 ;
        RECT 14.556 6.552 14.588 9.66 ;
  LAYER M1 ;
        RECT 14.556 9.624 14.588 9.696 ;
  LAYER M2 ;
        RECT 14.536 9.644 14.608 9.676 ;
  LAYER M1 ;
        RECT 14.556 3.408 14.588 3.48 ;
  LAYER M2 ;
        RECT 14.536 3.428 14.608 3.46 ;
  LAYER M1 ;
        RECT 14.556 3.444 14.588 6.552 ;
  LAYER M1 ;
        RECT 14.556 6.516 14.588 6.588 ;
  LAYER M2 ;
        RECT 14.536 6.536 14.608 6.568 ;
  LAYER M1 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M3 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M2 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M1 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M3 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M2 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M1 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M3 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M2 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M1 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M3 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M2 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M1 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M3 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M2 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M1 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M3 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M2 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M1 ;
        RECT 3.66 0.924 6.156 3.528 ;
  LAYER M3 ;
        RECT 3.66 0.924 6.156 3.528 ;
  LAYER M2 ;
        RECT 3.66 0.924 6.156 3.528 ;
  LAYER M1 ;
        RECT 3.66 4.032 6.156 6.636 ;
  LAYER M3 ;
        RECT 3.66 4.032 6.156 6.636 ;
  LAYER M2 ;
        RECT 3.66 4.032 6.156 6.636 ;
  LAYER M1 ;
        RECT 3.66 7.14 6.156 9.744 ;
  LAYER M3 ;
        RECT 3.66 7.14 6.156 9.744 ;
  LAYER M2 ;
        RECT 3.66 7.14 6.156 9.744 ;
  LAYER M1 ;
        RECT 3.66 10.248 6.156 12.852 ;
  LAYER M3 ;
        RECT 3.66 10.248 6.156 12.852 ;
  LAYER M2 ;
        RECT 3.66 10.248 6.156 12.852 ;
  LAYER M1 ;
        RECT 3.66 13.356 6.156 15.96 ;
  LAYER M3 ;
        RECT 3.66 13.356 6.156 15.96 ;
  LAYER M2 ;
        RECT 3.66 13.356 6.156 15.96 ;
  LAYER M1 ;
        RECT 3.66 16.464 6.156 19.068 ;
  LAYER M3 ;
        RECT 3.66 16.464 6.156 19.068 ;
  LAYER M2 ;
        RECT 3.66 16.464 6.156 19.068 ;
  LAYER M1 ;
        RECT 7.276 0.924 9.772 3.528 ;
  LAYER M3 ;
        RECT 7.276 0.924 9.772 3.528 ;
  LAYER M2 ;
        RECT 7.276 0.924 9.772 3.528 ;
  LAYER M1 ;
        RECT 7.276 4.032 9.772 6.636 ;
  LAYER M3 ;
        RECT 7.276 4.032 9.772 6.636 ;
  LAYER M2 ;
        RECT 7.276 4.032 9.772 6.636 ;
  LAYER M1 ;
        RECT 7.276 7.14 9.772 9.744 ;
  LAYER M3 ;
        RECT 7.276 7.14 9.772 9.744 ;
  LAYER M2 ;
        RECT 7.276 7.14 9.772 9.744 ;
  LAYER M1 ;
        RECT 7.276 10.248 9.772 12.852 ;
  LAYER M3 ;
        RECT 7.276 10.248 9.772 12.852 ;
  LAYER M2 ;
        RECT 7.276 10.248 9.772 12.852 ;
  LAYER M1 ;
        RECT 7.276 13.356 9.772 15.96 ;
  LAYER M3 ;
        RECT 7.276 13.356 9.772 15.96 ;
  LAYER M2 ;
        RECT 7.276 13.356 9.772 15.96 ;
  LAYER M1 ;
        RECT 7.276 16.464 9.772 19.068 ;
  LAYER M3 ;
        RECT 7.276 16.464 9.772 19.068 ;
  LAYER M2 ;
        RECT 7.276 16.464 9.772 19.068 ;
  LAYER M1 ;
        RECT 10.892 0.924 13.388 3.528 ;
  LAYER M3 ;
        RECT 10.892 0.924 13.388 3.528 ;
  LAYER M2 ;
        RECT 10.892 0.924 13.388 3.528 ;
  LAYER M1 ;
        RECT 10.892 4.032 13.388 6.636 ;
  LAYER M3 ;
        RECT 10.892 4.032 13.388 6.636 ;
  LAYER M2 ;
        RECT 10.892 4.032 13.388 6.636 ;
  LAYER M1 ;
        RECT 10.892 7.14 13.388 9.744 ;
  LAYER M3 ;
        RECT 10.892 7.14 13.388 9.744 ;
  LAYER M2 ;
        RECT 10.892 7.14 13.388 9.744 ;
  LAYER M1 ;
        RECT 10.892 10.248 13.388 12.852 ;
  LAYER M3 ;
        RECT 10.892 10.248 13.388 12.852 ;
  LAYER M2 ;
        RECT 10.892 10.248 13.388 12.852 ;
  LAYER M1 ;
        RECT 10.892 13.356 13.388 15.96 ;
  LAYER M3 ;
        RECT 10.892 13.356 13.388 15.96 ;
  LAYER M2 ;
        RECT 10.892 13.356 13.388 15.96 ;
  LAYER M1 ;
        RECT 10.892 16.464 13.388 19.068 ;
  LAYER M3 ;
        RECT 10.892 16.464 13.388 19.068 ;
  LAYER M2 ;
        RECT 10.892 16.464 13.388 19.068 ;
  LAYER M1 ;
        RECT 14.508 0.924 17.004 3.528 ;
  LAYER M3 ;
        RECT 14.508 0.924 17.004 3.528 ;
  LAYER M2 ;
        RECT 14.508 0.924 17.004 3.528 ;
  LAYER M1 ;
        RECT 14.508 4.032 17.004 6.636 ;
  LAYER M3 ;
        RECT 14.508 4.032 17.004 6.636 ;
  LAYER M2 ;
        RECT 14.508 4.032 17.004 6.636 ;
  LAYER M1 ;
        RECT 14.508 7.14 17.004 9.744 ;
  LAYER M3 ;
        RECT 14.508 7.14 17.004 9.744 ;
  LAYER M2 ;
        RECT 14.508 7.14 17.004 9.744 ;
  LAYER M1 ;
        RECT 14.508 10.248 17.004 12.852 ;
  LAYER M3 ;
        RECT 14.508 10.248 17.004 12.852 ;
  LAYER M2 ;
        RECT 14.508 10.248 17.004 12.852 ;
  LAYER M1 ;
        RECT 14.508 13.356 17.004 15.96 ;
  LAYER M3 ;
        RECT 14.508 13.356 17.004 15.96 ;
  LAYER M2 ;
        RECT 14.508 13.356 17.004 15.96 ;
  LAYER M1 ;
        RECT 14.508 16.464 17.004 19.068 ;
  LAYER M3 ;
        RECT 14.508 16.464 17.004 19.068 ;
  LAYER M2 ;
        RECT 14.508 16.464 17.004 19.068 ;
  END 
END Cap_30fF_Cap_60fF
