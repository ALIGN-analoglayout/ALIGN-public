MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 8.96 BY 24.528 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 24.24 3.136 24.312 ;
      LAYER M2 ;
        RECT 3.084 24.26 3.156 24.292 ;
      LAYER M1 ;
        RECT 5.984 24.24 6.016 24.312 ;
      LAYER M2 ;
        RECT 5.964 24.26 6.036 24.292 ;
      LAYER M2 ;
        RECT 3.12 24.26 6 24.292 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
      LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
      LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
      LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
      LAYER M2 ;
        RECT 2.96 0.236 5.84 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 3.264 9.54 3.296 9.612 ;
  LAYER M2 ;
        RECT 3.244 9.56 3.316 9.592 ;
  LAYER M2 ;
        RECT 2.96 9.56 3.28 9.592 ;
  LAYER M1 ;
        RECT 2.944 9.54 2.976 9.612 ;
  LAYER M2 ;
        RECT 2.924 9.56 2.996 9.592 ;
  LAYER M1 ;
        RECT 3.264 12.48 3.296 12.552 ;
  LAYER M2 ;
        RECT 3.244 12.5 3.316 12.532 ;
  LAYER M2 ;
        RECT 2.96 12.5 3.28 12.532 ;
  LAYER M1 ;
        RECT 2.944 12.48 2.976 12.552 ;
  LAYER M2 ;
        RECT 2.924 12.5 2.996 12.532 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 6.672 ;
  LAYER M2 ;
        RECT 3.244 6.62 3.316 6.652 ;
  LAYER M2 ;
        RECT 2.96 6.62 3.28 6.652 ;
  LAYER M1 ;
        RECT 2.944 6.6 2.976 6.672 ;
  LAYER M2 ;
        RECT 2.924 6.62 2.996 6.652 ;
  LAYER M1 ;
        RECT 3.264 15.42 3.296 15.492 ;
  LAYER M2 ;
        RECT 3.244 15.44 3.316 15.472 ;
  LAYER M2 ;
        RECT 2.96 15.44 3.28 15.472 ;
  LAYER M1 ;
        RECT 2.944 15.42 2.976 15.492 ;
  LAYER M2 ;
        RECT 2.924 15.44 2.996 15.472 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 3.732 ;
  LAYER M2 ;
        RECT 3.244 3.68 3.316 3.712 ;
  LAYER M2 ;
        RECT 2.96 3.68 3.28 3.712 ;
  LAYER M1 ;
        RECT 2.944 3.66 2.976 3.732 ;
  LAYER M2 ;
        RECT 2.924 3.68 2.996 3.712 ;
  LAYER M1 ;
        RECT 3.264 18.36 3.296 18.432 ;
  LAYER M2 ;
        RECT 3.244 18.38 3.316 18.412 ;
  LAYER M2 ;
        RECT 2.96 18.38 3.28 18.412 ;
  LAYER M1 ;
        RECT 2.944 18.36 2.976 18.432 ;
  LAYER M2 ;
        RECT 2.924 18.38 2.996 18.412 ;
  LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
  LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
  LAYER M1 ;
        RECT 2.944 0.252 2.976 0.42 ;
  LAYER M1 ;
        RECT 2.944 0.42 2.976 18.396 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 9.612 ;
  LAYER M2 ;
        RECT 3.244 9.56 3.316 9.592 ;
  LAYER M1 ;
        RECT 3.264 9.408 3.296 9.576 ;
  LAYER M1 ;
        RECT 3.264 9.372 3.296 9.444 ;
  LAYER M2 ;
        RECT 3.244 9.392 3.316 9.424 ;
  LAYER M2 ;
        RECT 3.28 9.392 5.84 9.424 ;
  LAYER M1 ;
        RECT 5.824 9.372 5.856 9.444 ;
  LAYER M2 ;
        RECT 5.804 9.392 5.876 9.424 ;
  LAYER M1 ;
        RECT 3.264 12.48 3.296 12.552 ;
  LAYER M2 ;
        RECT 3.244 12.5 3.316 12.532 ;
  LAYER M1 ;
        RECT 3.264 12.348 3.296 12.516 ;
  LAYER M1 ;
        RECT 3.264 12.312 3.296 12.384 ;
  LAYER M2 ;
        RECT 3.244 12.332 3.316 12.364 ;
  LAYER M2 ;
        RECT 3.28 12.332 5.84 12.364 ;
  LAYER M1 ;
        RECT 5.824 12.312 5.856 12.384 ;
  LAYER M2 ;
        RECT 5.804 12.332 5.876 12.364 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 6.672 ;
  LAYER M2 ;
        RECT 3.244 6.62 3.316 6.652 ;
  LAYER M1 ;
        RECT 3.264 6.468 3.296 6.636 ;
  LAYER M1 ;
        RECT 3.264 6.432 3.296 6.504 ;
  LAYER M2 ;
        RECT 3.244 6.452 3.316 6.484 ;
  LAYER M2 ;
        RECT 3.28 6.452 5.84 6.484 ;
  LAYER M1 ;
        RECT 5.824 6.432 5.856 6.504 ;
  LAYER M2 ;
        RECT 5.804 6.452 5.876 6.484 ;
  LAYER M1 ;
        RECT 3.264 15.42 3.296 15.492 ;
  LAYER M2 ;
        RECT 3.244 15.44 3.316 15.472 ;
  LAYER M1 ;
        RECT 3.264 15.288 3.296 15.456 ;
  LAYER M1 ;
        RECT 3.264 15.252 3.296 15.324 ;
  LAYER M2 ;
        RECT 3.244 15.272 3.316 15.304 ;
  LAYER M2 ;
        RECT 3.28 15.272 5.84 15.304 ;
  LAYER M1 ;
        RECT 5.824 15.252 5.856 15.324 ;
  LAYER M2 ;
        RECT 5.804 15.272 5.876 15.304 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 3.732 ;
  LAYER M2 ;
        RECT 3.244 3.68 3.316 3.712 ;
  LAYER M1 ;
        RECT 3.264 3.528 3.296 3.696 ;
  LAYER M1 ;
        RECT 3.264 3.492 3.296 3.564 ;
  LAYER M2 ;
        RECT 3.244 3.512 3.316 3.544 ;
  LAYER M2 ;
        RECT 3.28 3.512 5.84 3.544 ;
  LAYER M1 ;
        RECT 5.824 3.492 5.856 3.564 ;
  LAYER M2 ;
        RECT 5.804 3.512 5.876 3.544 ;
  LAYER M1 ;
        RECT 3.264 18.36 3.296 18.432 ;
  LAYER M2 ;
        RECT 3.244 18.38 3.316 18.412 ;
  LAYER M1 ;
        RECT 3.264 18.228 3.296 18.396 ;
  LAYER M1 ;
        RECT 3.264 18.192 3.296 18.264 ;
  LAYER M2 ;
        RECT 3.244 18.212 3.316 18.244 ;
  LAYER M2 ;
        RECT 3.28 18.212 5.84 18.244 ;
  LAYER M1 ;
        RECT 5.824 18.192 5.856 18.264 ;
  LAYER M2 ;
        RECT 5.804 18.212 5.876 18.244 ;
  LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
  LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
  LAYER M1 ;
        RECT 5.824 0.252 5.856 0.42 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 18.228 ;
  LAYER M2 ;
        RECT 2.96 0.236 5.84 0.268 ;
  LAYER M1 ;
        RECT 0.384 0.72 0.416 0.792 ;
  LAYER M2 ;
        RECT 0.364 0.74 0.436 0.772 ;
  LAYER M2 ;
        RECT 0.08 0.74 0.4 0.772 ;
  LAYER M1 ;
        RECT 0.064 0.72 0.096 0.792 ;
  LAYER M2 ;
        RECT 0.044 0.74 0.116 0.772 ;
  LAYER M1 ;
        RECT 0.384 3.66 0.416 3.732 ;
  LAYER M2 ;
        RECT 0.364 3.68 0.436 3.712 ;
  LAYER M2 ;
        RECT 0.08 3.68 0.4 3.712 ;
  LAYER M1 ;
        RECT 0.064 3.66 0.096 3.732 ;
  LAYER M2 ;
        RECT 0.044 3.68 0.116 3.712 ;
  LAYER M1 ;
        RECT 0.384 6.6 0.416 6.672 ;
  LAYER M2 ;
        RECT 0.364 6.62 0.436 6.652 ;
  LAYER M2 ;
        RECT 0.08 6.62 0.4 6.652 ;
  LAYER M1 ;
        RECT 0.064 6.6 0.096 6.672 ;
  LAYER M2 ;
        RECT 0.044 6.62 0.116 6.652 ;
  LAYER M1 ;
        RECT 0.384 9.54 0.416 9.612 ;
  LAYER M2 ;
        RECT 0.364 9.56 0.436 9.592 ;
  LAYER M2 ;
        RECT 0.08 9.56 0.4 9.592 ;
  LAYER M1 ;
        RECT 0.064 9.54 0.096 9.612 ;
  LAYER M2 ;
        RECT 0.044 9.56 0.116 9.592 ;
  LAYER M1 ;
        RECT 0.384 12.48 0.416 12.552 ;
  LAYER M2 ;
        RECT 0.364 12.5 0.436 12.532 ;
  LAYER M2 ;
        RECT 0.08 12.5 0.4 12.532 ;
  LAYER M1 ;
        RECT 0.064 12.48 0.096 12.552 ;
  LAYER M2 ;
        RECT 0.044 12.5 0.116 12.532 ;
  LAYER M1 ;
        RECT 0.384 15.42 0.416 15.492 ;
  LAYER M2 ;
        RECT 0.364 15.44 0.436 15.472 ;
  LAYER M2 ;
        RECT 0.08 15.44 0.4 15.472 ;
  LAYER M1 ;
        RECT 0.064 15.42 0.096 15.492 ;
  LAYER M2 ;
        RECT 0.044 15.44 0.116 15.472 ;
  LAYER M1 ;
        RECT 0.384 18.36 0.416 18.432 ;
  LAYER M2 ;
        RECT 0.364 18.38 0.436 18.412 ;
  LAYER M2 ;
        RECT 0.08 18.38 0.4 18.412 ;
  LAYER M1 ;
        RECT 0.064 18.36 0.096 18.432 ;
  LAYER M2 ;
        RECT 0.044 18.38 0.116 18.412 ;
  LAYER M1 ;
        RECT 0.384 21.3 0.416 21.372 ;
  LAYER M2 ;
        RECT 0.364 21.32 0.436 21.352 ;
  LAYER M2 ;
        RECT 0.08 21.32 0.4 21.352 ;
  LAYER M1 ;
        RECT 0.064 21.3 0.096 21.372 ;
  LAYER M2 ;
        RECT 0.044 21.32 0.116 21.352 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.42 ;
  LAYER M1 ;
        RECT 0.064 0.42 0.096 21.336 ;
  LAYER M1 ;
        RECT 6.144 0.72 6.176 0.792 ;
  LAYER M2 ;
        RECT 6.124 0.74 6.196 0.772 ;
  LAYER M1 ;
        RECT 6.144 0.588 6.176 0.756 ;
  LAYER M1 ;
        RECT 6.144 0.552 6.176 0.624 ;
  LAYER M2 ;
        RECT 6.124 0.572 6.196 0.604 ;
  LAYER M2 ;
        RECT 6.16 0.572 8.72 0.604 ;
  LAYER M1 ;
        RECT 8.704 0.552 8.736 0.624 ;
  LAYER M2 ;
        RECT 8.684 0.572 8.756 0.604 ;
  LAYER M1 ;
        RECT 6.144 3.66 6.176 3.732 ;
  LAYER M2 ;
        RECT 6.124 3.68 6.196 3.712 ;
  LAYER M1 ;
        RECT 6.144 3.528 6.176 3.696 ;
  LAYER M1 ;
        RECT 6.144 3.492 6.176 3.564 ;
  LAYER M2 ;
        RECT 6.124 3.512 6.196 3.544 ;
  LAYER M2 ;
        RECT 6.16 3.512 8.72 3.544 ;
  LAYER M1 ;
        RECT 8.704 3.492 8.736 3.564 ;
  LAYER M2 ;
        RECT 8.684 3.512 8.756 3.544 ;
  LAYER M1 ;
        RECT 6.144 6.6 6.176 6.672 ;
  LAYER M2 ;
        RECT 6.124 6.62 6.196 6.652 ;
  LAYER M1 ;
        RECT 6.144 6.468 6.176 6.636 ;
  LAYER M1 ;
        RECT 6.144 6.432 6.176 6.504 ;
  LAYER M2 ;
        RECT 6.124 6.452 6.196 6.484 ;
  LAYER M2 ;
        RECT 6.16 6.452 8.72 6.484 ;
  LAYER M1 ;
        RECT 8.704 6.432 8.736 6.504 ;
  LAYER M2 ;
        RECT 8.684 6.452 8.756 6.484 ;
  LAYER M1 ;
        RECT 6.144 9.54 6.176 9.612 ;
  LAYER M2 ;
        RECT 6.124 9.56 6.196 9.592 ;
  LAYER M1 ;
        RECT 6.144 9.408 6.176 9.576 ;
  LAYER M1 ;
        RECT 6.144 9.372 6.176 9.444 ;
  LAYER M2 ;
        RECT 6.124 9.392 6.196 9.424 ;
  LAYER M2 ;
        RECT 6.16 9.392 8.72 9.424 ;
  LAYER M1 ;
        RECT 8.704 9.372 8.736 9.444 ;
  LAYER M2 ;
        RECT 8.684 9.392 8.756 9.424 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 12.552 ;
  LAYER M2 ;
        RECT 6.124 12.5 6.196 12.532 ;
  LAYER M1 ;
        RECT 6.144 12.348 6.176 12.516 ;
  LAYER M1 ;
        RECT 6.144 12.312 6.176 12.384 ;
  LAYER M2 ;
        RECT 6.124 12.332 6.196 12.364 ;
  LAYER M2 ;
        RECT 6.16 12.332 8.72 12.364 ;
  LAYER M1 ;
        RECT 8.704 12.312 8.736 12.384 ;
  LAYER M2 ;
        RECT 8.684 12.332 8.756 12.364 ;
  LAYER M1 ;
        RECT 6.144 15.42 6.176 15.492 ;
  LAYER M2 ;
        RECT 6.124 15.44 6.196 15.472 ;
  LAYER M1 ;
        RECT 6.144 15.288 6.176 15.456 ;
  LAYER M1 ;
        RECT 6.144 15.252 6.176 15.324 ;
  LAYER M2 ;
        RECT 6.124 15.272 6.196 15.304 ;
  LAYER M2 ;
        RECT 6.16 15.272 8.72 15.304 ;
  LAYER M1 ;
        RECT 8.704 15.252 8.736 15.324 ;
  LAYER M2 ;
        RECT 8.684 15.272 8.756 15.304 ;
  LAYER M1 ;
        RECT 6.144 18.36 6.176 18.432 ;
  LAYER M2 ;
        RECT 6.124 18.38 6.196 18.412 ;
  LAYER M1 ;
        RECT 6.144 18.228 6.176 18.396 ;
  LAYER M1 ;
        RECT 6.144 18.192 6.176 18.264 ;
  LAYER M2 ;
        RECT 6.124 18.212 6.196 18.244 ;
  LAYER M2 ;
        RECT 6.16 18.212 8.72 18.244 ;
  LAYER M1 ;
        RECT 8.704 18.192 8.736 18.264 ;
  LAYER M2 ;
        RECT 8.684 18.212 8.756 18.244 ;
  LAYER M1 ;
        RECT 6.144 21.3 6.176 21.372 ;
  LAYER M2 ;
        RECT 6.124 21.32 6.196 21.352 ;
  LAYER M1 ;
        RECT 6.144 21.168 6.176 21.336 ;
  LAYER M1 ;
        RECT 6.144 21.132 6.176 21.204 ;
  LAYER M2 ;
        RECT 6.124 21.152 6.196 21.184 ;
  LAYER M2 ;
        RECT 6.16 21.152 8.72 21.184 ;
  LAYER M1 ;
        RECT 8.704 21.132 8.736 21.204 ;
  LAYER M2 ;
        RECT 8.684 21.152 8.756 21.184 ;
  LAYER M1 ;
        RECT 8.704 0.048 8.736 0.12 ;
  LAYER M2 ;
        RECT 8.684 0.068 8.756 0.1 ;
  LAYER M1 ;
        RECT 8.704 0.084 8.736 0.42 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 21.168 ;
  LAYER M2 ;
        RECT 0.08 0.068 8.72 0.1 ;
  LAYER M1 ;
        RECT 3.264 0.72 3.296 0.792 ;
  LAYER M2 ;
        RECT 3.244 0.74 3.316 0.772 ;
  LAYER M2 ;
        RECT 0.4 0.74 3.28 0.772 ;
  LAYER M1 ;
        RECT 0.384 0.72 0.416 0.792 ;
  LAYER M2 ;
        RECT 0.364 0.74 0.436 0.772 ;
  LAYER M1 ;
        RECT 3.264 21.3 3.296 21.372 ;
  LAYER M2 ;
        RECT 3.244 21.32 3.316 21.352 ;
  LAYER M2 ;
        RECT 0.4 21.32 3.28 21.352 ;
  LAYER M1 ;
        RECT 0.384 21.3 0.416 21.372 ;
  LAYER M2 ;
        RECT 0.364 21.32 0.436 21.352 ;
  LAYER M1 ;
        RECT 5.664 11.976 5.696 12.048 ;
  LAYER M2 ;
        RECT 5.644 11.996 5.716 12.028 ;
  LAYER M2 ;
        RECT 3.12 11.996 5.68 12.028 ;
  LAYER M1 ;
        RECT 3.104 11.976 3.136 12.048 ;
  LAYER M2 ;
        RECT 3.084 11.996 3.156 12.028 ;
  LAYER M1 ;
        RECT 5.664 14.916 5.696 14.988 ;
  LAYER M2 ;
        RECT 5.644 14.936 5.716 14.968 ;
  LAYER M2 ;
        RECT 3.12 14.936 5.68 14.968 ;
  LAYER M1 ;
        RECT 3.104 14.916 3.136 14.988 ;
  LAYER M2 ;
        RECT 3.084 14.936 3.156 14.968 ;
  LAYER M1 ;
        RECT 5.664 9.036 5.696 9.108 ;
  LAYER M2 ;
        RECT 5.644 9.056 5.716 9.088 ;
  LAYER M2 ;
        RECT 3.12 9.056 5.68 9.088 ;
  LAYER M1 ;
        RECT 3.104 9.036 3.136 9.108 ;
  LAYER M2 ;
        RECT 3.084 9.056 3.156 9.088 ;
  LAYER M1 ;
        RECT 5.664 17.856 5.696 17.928 ;
  LAYER M2 ;
        RECT 5.644 17.876 5.716 17.908 ;
  LAYER M2 ;
        RECT 3.12 17.876 5.68 17.908 ;
  LAYER M1 ;
        RECT 3.104 17.856 3.136 17.928 ;
  LAYER M2 ;
        RECT 3.084 17.876 3.156 17.908 ;
  LAYER M1 ;
        RECT 5.664 6.096 5.696 6.168 ;
  LAYER M2 ;
        RECT 5.644 6.116 5.716 6.148 ;
  LAYER M2 ;
        RECT 3.12 6.116 5.68 6.148 ;
  LAYER M1 ;
        RECT 3.104 6.096 3.136 6.168 ;
  LAYER M2 ;
        RECT 3.084 6.116 3.156 6.148 ;
  LAYER M1 ;
        RECT 5.664 20.796 5.696 20.868 ;
  LAYER M2 ;
        RECT 5.644 20.816 5.716 20.848 ;
  LAYER M2 ;
        RECT 3.12 20.816 5.68 20.848 ;
  LAYER M1 ;
        RECT 3.104 20.796 3.136 20.868 ;
  LAYER M2 ;
        RECT 3.084 20.816 3.156 20.848 ;
  LAYER M1 ;
        RECT 3.104 24.24 3.136 24.312 ;
  LAYER M2 ;
        RECT 3.084 24.26 3.156 24.292 ;
  LAYER M1 ;
        RECT 3.104 24.108 3.136 24.276 ;
  LAYER M1 ;
        RECT 3.104 6.132 3.136 24.108 ;
  LAYER M1 ;
        RECT 5.664 11.976 5.696 12.048 ;
  LAYER M2 ;
        RECT 5.644 11.996 5.716 12.028 ;
  LAYER M1 ;
        RECT 5.664 12.012 5.696 12.18 ;
  LAYER M1 ;
        RECT 5.664 12.144 5.696 12.216 ;
  LAYER M2 ;
        RECT 5.644 12.164 5.716 12.196 ;
  LAYER M2 ;
        RECT 5.68 12.164 6 12.196 ;
  LAYER M1 ;
        RECT 5.984 12.144 6.016 12.216 ;
  LAYER M2 ;
        RECT 5.964 12.164 6.036 12.196 ;
  LAYER M1 ;
        RECT 5.664 14.916 5.696 14.988 ;
  LAYER M2 ;
        RECT 5.644 14.936 5.716 14.968 ;
  LAYER M1 ;
        RECT 5.664 14.952 5.696 15.12 ;
  LAYER M1 ;
        RECT 5.664 15.084 5.696 15.156 ;
  LAYER M2 ;
        RECT 5.644 15.104 5.716 15.136 ;
  LAYER M2 ;
        RECT 5.68 15.104 6 15.136 ;
  LAYER M1 ;
        RECT 5.984 15.084 6.016 15.156 ;
  LAYER M2 ;
        RECT 5.964 15.104 6.036 15.136 ;
  LAYER M1 ;
        RECT 5.664 9.036 5.696 9.108 ;
  LAYER M2 ;
        RECT 5.644 9.056 5.716 9.088 ;
  LAYER M1 ;
        RECT 5.664 9.072 5.696 9.24 ;
  LAYER M1 ;
        RECT 5.664 9.204 5.696 9.276 ;
  LAYER M2 ;
        RECT 5.644 9.224 5.716 9.256 ;
  LAYER M2 ;
        RECT 5.68 9.224 6 9.256 ;
  LAYER M1 ;
        RECT 5.984 9.204 6.016 9.276 ;
  LAYER M2 ;
        RECT 5.964 9.224 6.036 9.256 ;
  LAYER M1 ;
        RECT 5.664 17.856 5.696 17.928 ;
  LAYER M2 ;
        RECT 5.644 17.876 5.716 17.908 ;
  LAYER M1 ;
        RECT 5.664 17.892 5.696 18.06 ;
  LAYER M1 ;
        RECT 5.664 18.024 5.696 18.096 ;
  LAYER M2 ;
        RECT 5.644 18.044 5.716 18.076 ;
  LAYER M2 ;
        RECT 5.68 18.044 6 18.076 ;
  LAYER M1 ;
        RECT 5.984 18.024 6.016 18.096 ;
  LAYER M2 ;
        RECT 5.964 18.044 6.036 18.076 ;
  LAYER M1 ;
        RECT 5.664 6.096 5.696 6.168 ;
  LAYER M2 ;
        RECT 5.644 6.116 5.716 6.148 ;
  LAYER M1 ;
        RECT 5.664 6.132 5.696 6.3 ;
  LAYER M1 ;
        RECT 5.664 6.264 5.696 6.336 ;
  LAYER M2 ;
        RECT 5.644 6.284 5.716 6.316 ;
  LAYER M2 ;
        RECT 5.68 6.284 6 6.316 ;
  LAYER M1 ;
        RECT 5.984 6.264 6.016 6.336 ;
  LAYER M2 ;
        RECT 5.964 6.284 6.036 6.316 ;
  LAYER M1 ;
        RECT 5.664 20.796 5.696 20.868 ;
  LAYER M2 ;
        RECT 5.644 20.816 5.716 20.848 ;
  LAYER M1 ;
        RECT 5.664 20.832 5.696 21 ;
  LAYER M1 ;
        RECT 5.664 20.964 5.696 21.036 ;
  LAYER M2 ;
        RECT 5.644 20.984 5.716 21.016 ;
  LAYER M2 ;
        RECT 5.68 20.984 6 21.016 ;
  LAYER M1 ;
        RECT 5.984 20.964 6.016 21.036 ;
  LAYER M2 ;
        RECT 5.964 20.984 6.036 21.016 ;
  LAYER M1 ;
        RECT 5.984 24.24 6.016 24.312 ;
  LAYER M2 ;
        RECT 5.964 24.26 6.036 24.292 ;
  LAYER M1 ;
        RECT 5.984 24.108 6.016 24.276 ;
  LAYER M1 ;
        RECT 5.984 6.3 6.016 24.108 ;
  LAYER M2 ;
        RECT 3.12 24.26 6 24.292 ;
  LAYER M1 ;
        RECT 2.784 3.156 2.816 3.228 ;
  LAYER M2 ;
        RECT 2.764 3.176 2.836 3.208 ;
  LAYER M2 ;
        RECT 0.24 3.176 2.8 3.208 ;
  LAYER M1 ;
        RECT 0.224 3.156 0.256 3.228 ;
  LAYER M2 ;
        RECT 0.204 3.176 0.276 3.208 ;
  LAYER M1 ;
        RECT 2.784 6.096 2.816 6.168 ;
  LAYER M2 ;
        RECT 2.764 6.116 2.836 6.148 ;
  LAYER M2 ;
        RECT 0.24 6.116 2.8 6.148 ;
  LAYER M1 ;
        RECT 0.224 6.096 0.256 6.168 ;
  LAYER M2 ;
        RECT 0.204 6.116 0.276 6.148 ;
  LAYER M1 ;
        RECT 2.784 9.036 2.816 9.108 ;
  LAYER M2 ;
        RECT 2.764 9.056 2.836 9.088 ;
  LAYER M2 ;
        RECT 0.24 9.056 2.8 9.088 ;
  LAYER M1 ;
        RECT 0.224 9.036 0.256 9.108 ;
  LAYER M2 ;
        RECT 0.204 9.056 0.276 9.088 ;
  LAYER M1 ;
        RECT 2.784 11.976 2.816 12.048 ;
  LAYER M2 ;
        RECT 2.764 11.996 2.836 12.028 ;
  LAYER M2 ;
        RECT 0.24 11.996 2.8 12.028 ;
  LAYER M1 ;
        RECT 0.224 11.976 0.256 12.048 ;
  LAYER M2 ;
        RECT 0.204 11.996 0.276 12.028 ;
  LAYER M1 ;
        RECT 2.784 14.916 2.816 14.988 ;
  LAYER M2 ;
        RECT 2.764 14.936 2.836 14.968 ;
  LAYER M2 ;
        RECT 0.24 14.936 2.8 14.968 ;
  LAYER M1 ;
        RECT 0.224 14.916 0.256 14.988 ;
  LAYER M2 ;
        RECT 0.204 14.936 0.276 14.968 ;
  LAYER M1 ;
        RECT 2.784 17.856 2.816 17.928 ;
  LAYER M2 ;
        RECT 2.764 17.876 2.836 17.908 ;
  LAYER M2 ;
        RECT 0.24 17.876 2.8 17.908 ;
  LAYER M1 ;
        RECT 0.224 17.856 0.256 17.928 ;
  LAYER M2 ;
        RECT 0.204 17.876 0.276 17.908 ;
  LAYER M1 ;
        RECT 2.784 20.796 2.816 20.868 ;
  LAYER M2 ;
        RECT 2.764 20.816 2.836 20.848 ;
  LAYER M2 ;
        RECT 0.24 20.816 2.8 20.848 ;
  LAYER M1 ;
        RECT 0.224 20.796 0.256 20.868 ;
  LAYER M2 ;
        RECT 0.204 20.816 0.276 20.848 ;
  LAYER M1 ;
        RECT 2.784 23.736 2.816 23.808 ;
  LAYER M2 ;
        RECT 2.764 23.756 2.836 23.788 ;
  LAYER M2 ;
        RECT 0.24 23.756 2.8 23.788 ;
  LAYER M1 ;
        RECT 0.224 23.736 0.256 23.808 ;
  LAYER M2 ;
        RECT 0.204 23.756 0.276 23.788 ;
  LAYER M1 ;
        RECT 0.224 24.408 0.256 24.48 ;
  LAYER M2 ;
        RECT 0.204 24.428 0.276 24.46 ;
  LAYER M1 ;
        RECT 0.224 24.108 0.256 24.444 ;
  LAYER M1 ;
        RECT 0.224 3.192 0.256 24.108 ;
  LAYER M1 ;
        RECT 8.544 3.156 8.576 3.228 ;
  LAYER M2 ;
        RECT 8.524 3.176 8.596 3.208 ;
  LAYER M1 ;
        RECT 8.544 3.192 8.576 3.36 ;
  LAYER M1 ;
        RECT 8.544 3.324 8.576 3.396 ;
  LAYER M2 ;
        RECT 8.524 3.344 8.596 3.376 ;
  LAYER M2 ;
        RECT 8.56 3.344 8.88 3.376 ;
  LAYER M1 ;
        RECT 8.864 3.324 8.896 3.396 ;
  LAYER M2 ;
        RECT 8.844 3.344 8.916 3.376 ;
  LAYER M1 ;
        RECT 8.544 6.096 8.576 6.168 ;
  LAYER M2 ;
        RECT 8.524 6.116 8.596 6.148 ;
  LAYER M1 ;
        RECT 8.544 6.132 8.576 6.3 ;
  LAYER M1 ;
        RECT 8.544 6.264 8.576 6.336 ;
  LAYER M2 ;
        RECT 8.524 6.284 8.596 6.316 ;
  LAYER M2 ;
        RECT 8.56 6.284 8.88 6.316 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M1 ;
        RECT 8.544 9.036 8.576 9.108 ;
  LAYER M2 ;
        RECT 8.524 9.056 8.596 9.088 ;
  LAYER M1 ;
        RECT 8.544 9.072 8.576 9.24 ;
  LAYER M1 ;
        RECT 8.544 9.204 8.576 9.276 ;
  LAYER M2 ;
        RECT 8.524 9.224 8.596 9.256 ;
  LAYER M2 ;
        RECT 8.56 9.224 8.88 9.256 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M1 ;
        RECT 8.544 11.976 8.576 12.048 ;
  LAYER M2 ;
        RECT 8.524 11.996 8.596 12.028 ;
  LAYER M1 ;
        RECT 8.544 12.012 8.576 12.18 ;
  LAYER M1 ;
        RECT 8.544 12.144 8.576 12.216 ;
  LAYER M2 ;
        RECT 8.524 12.164 8.596 12.196 ;
  LAYER M2 ;
        RECT 8.56 12.164 8.88 12.196 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M1 ;
        RECT 8.544 14.916 8.576 14.988 ;
  LAYER M2 ;
        RECT 8.524 14.936 8.596 14.968 ;
  LAYER M1 ;
        RECT 8.544 14.952 8.576 15.12 ;
  LAYER M1 ;
        RECT 8.544 15.084 8.576 15.156 ;
  LAYER M2 ;
        RECT 8.524 15.104 8.596 15.136 ;
  LAYER M2 ;
        RECT 8.56 15.104 8.88 15.136 ;
  LAYER M1 ;
        RECT 8.864 15.084 8.896 15.156 ;
  LAYER M2 ;
        RECT 8.844 15.104 8.916 15.136 ;
  LAYER M1 ;
        RECT 8.544 17.856 8.576 17.928 ;
  LAYER M2 ;
        RECT 8.524 17.876 8.596 17.908 ;
  LAYER M1 ;
        RECT 8.544 17.892 8.576 18.06 ;
  LAYER M1 ;
        RECT 8.544 18.024 8.576 18.096 ;
  LAYER M2 ;
        RECT 8.524 18.044 8.596 18.076 ;
  LAYER M2 ;
        RECT 8.56 18.044 8.88 18.076 ;
  LAYER M1 ;
        RECT 8.864 18.024 8.896 18.096 ;
  LAYER M2 ;
        RECT 8.844 18.044 8.916 18.076 ;
  LAYER M1 ;
        RECT 8.544 20.796 8.576 20.868 ;
  LAYER M2 ;
        RECT 8.524 20.816 8.596 20.848 ;
  LAYER M1 ;
        RECT 8.544 20.832 8.576 21 ;
  LAYER M1 ;
        RECT 8.544 20.964 8.576 21.036 ;
  LAYER M2 ;
        RECT 8.524 20.984 8.596 21.016 ;
  LAYER M2 ;
        RECT 8.56 20.984 8.88 21.016 ;
  LAYER M1 ;
        RECT 8.864 20.964 8.896 21.036 ;
  LAYER M2 ;
        RECT 8.844 20.984 8.916 21.016 ;
  LAYER M1 ;
        RECT 8.544 23.736 8.576 23.808 ;
  LAYER M2 ;
        RECT 8.524 23.756 8.596 23.788 ;
  LAYER M1 ;
        RECT 8.544 23.772 8.576 23.94 ;
  LAYER M1 ;
        RECT 8.544 23.904 8.576 23.976 ;
  LAYER M2 ;
        RECT 8.524 23.924 8.596 23.956 ;
  LAYER M2 ;
        RECT 8.56 23.924 8.88 23.956 ;
  LAYER M1 ;
        RECT 8.864 23.904 8.896 23.976 ;
  LAYER M2 ;
        RECT 8.844 23.924 8.916 23.956 ;
  LAYER M1 ;
        RECT 8.864 24.408 8.896 24.48 ;
  LAYER M2 ;
        RECT 8.844 24.428 8.916 24.46 ;
  LAYER M1 ;
        RECT 8.864 24.108 8.896 24.444 ;
  LAYER M1 ;
        RECT 8.864 3.36 8.896 24.108 ;
  LAYER M2 ;
        RECT 0.24 24.428 8.88 24.46 ;
  LAYER M1 ;
        RECT 5.664 3.156 5.696 3.228 ;
  LAYER M2 ;
        RECT 5.644 3.176 5.716 3.208 ;
  LAYER M2 ;
        RECT 2.8 3.176 5.68 3.208 ;
  LAYER M1 ;
        RECT 2.784 3.156 2.816 3.228 ;
  LAYER M2 ;
        RECT 2.764 3.176 2.836 3.208 ;
  LAYER M1 ;
        RECT 5.664 23.736 5.696 23.808 ;
  LAYER M2 ;
        RECT 5.644 23.756 5.716 23.788 ;
  LAYER M2 ;
        RECT 2.8 23.756 5.68 23.788 ;
  LAYER M1 ;
        RECT 2.784 23.736 2.816 23.808 ;
  LAYER M2 ;
        RECT 2.764 23.756 2.836 23.788 ;
  LAYER M1 ;
        RECT 0.384 0.72 0.416 3.228 ;
  LAYER M1 ;
        RECT 0.448 0.72 0.48 3.228 ;
  LAYER M1 ;
        RECT 0.512 0.72 0.544 3.228 ;
  LAYER M1 ;
        RECT 0.576 0.72 0.608 3.228 ;
  LAYER M1 ;
        RECT 0.64 0.72 0.672 3.228 ;
  LAYER M1 ;
        RECT 0.704 0.72 0.736 3.228 ;
  LAYER M1 ;
        RECT 0.768 0.72 0.8 3.228 ;
  LAYER M1 ;
        RECT 0.832 0.72 0.864 3.228 ;
  LAYER M1 ;
        RECT 0.896 0.72 0.928 3.228 ;
  LAYER M1 ;
        RECT 0.96 0.72 0.992 3.228 ;
  LAYER M1 ;
        RECT 1.024 0.72 1.056 3.228 ;
  LAYER M1 ;
        RECT 1.088 0.72 1.12 3.228 ;
  LAYER M1 ;
        RECT 1.152 0.72 1.184 3.228 ;
  LAYER M1 ;
        RECT 1.216 0.72 1.248 3.228 ;
  LAYER M1 ;
        RECT 1.28 0.72 1.312 3.228 ;
  LAYER M1 ;
        RECT 1.344 0.72 1.376 3.228 ;
  LAYER M1 ;
        RECT 1.408 0.72 1.44 3.228 ;
  LAYER M1 ;
        RECT 1.472 0.72 1.504 3.228 ;
  LAYER M1 ;
        RECT 1.536 0.72 1.568 3.228 ;
  LAYER M1 ;
        RECT 1.6 0.72 1.632 3.228 ;
  LAYER M1 ;
        RECT 1.664 0.72 1.696 3.228 ;
  LAYER M1 ;
        RECT 1.728 0.72 1.76 3.228 ;
  LAYER M1 ;
        RECT 1.792 0.72 1.824 3.228 ;
  LAYER M1 ;
        RECT 1.856 0.72 1.888 3.228 ;
  LAYER M1 ;
        RECT 1.92 0.72 1.952 3.228 ;
  LAYER M1 ;
        RECT 1.984 0.72 2.016 3.228 ;
  LAYER M1 ;
        RECT 2.048 0.72 2.08 3.228 ;
  LAYER M1 ;
        RECT 2.112 0.72 2.144 3.228 ;
  LAYER M1 ;
        RECT 2.176 0.72 2.208 3.228 ;
  LAYER M1 ;
        RECT 2.24 0.72 2.272 3.228 ;
  LAYER M1 ;
        RECT 2.304 0.72 2.336 3.228 ;
  LAYER M1 ;
        RECT 2.368 0.72 2.4 3.228 ;
  LAYER M1 ;
        RECT 2.432 0.72 2.464 3.228 ;
  LAYER M1 ;
        RECT 2.496 0.72 2.528 3.228 ;
  LAYER M1 ;
        RECT 2.56 0.72 2.592 3.228 ;
  LAYER M1 ;
        RECT 2.624 0.72 2.656 3.228 ;
  LAYER M1 ;
        RECT 2.688 0.72 2.72 3.228 ;
  LAYER M2 ;
        RECT 0.364 0.804 2.836 0.836 ;
  LAYER M2 ;
        RECT 0.364 0.868 2.836 0.9 ;
  LAYER M2 ;
        RECT 0.364 0.932 2.836 0.964 ;
  LAYER M2 ;
        RECT 0.364 0.996 2.836 1.028 ;
  LAYER M2 ;
        RECT 0.364 1.06 2.836 1.092 ;
  LAYER M2 ;
        RECT 0.364 1.124 2.836 1.156 ;
  LAYER M2 ;
        RECT 0.364 1.188 2.836 1.22 ;
  LAYER M2 ;
        RECT 0.364 1.252 2.836 1.284 ;
  LAYER M2 ;
        RECT 0.364 1.316 2.836 1.348 ;
  LAYER M2 ;
        RECT 0.364 1.38 2.836 1.412 ;
  LAYER M2 ;
        RECT 0.364 1.444 2.836 1.476 ;
  LAYER M2 ;
        RECT 0.364 1.508 2.836 1.54 ;
  LAYER M2 ;
        RECT 0.364 1.572 2.836 1.604 ;
  LAYER M2 ;
        RECT 0.364 1.636 2.836 1.668 ;
  LAYER M2 ;
        RECT 0.364 1.7 2.836 1.732 ;
  LAYER M2 ;
        RECT 0.364 1.764 2.836 1.796 ;
  LAYER M2 ;
        RECT 0.364 1.828 2.836 1.86 ;
  LAYER M2 ;
        RECT 0.364 1.892 2.836 1.924 ;
  LAYER M2 ;
        RECT 0.364 1.956 2.836 1.988 ;
  LAYER M2 ;
        RECT 0.364 2.02 2.836 2.052 ;
  LAYER M2 ;
        RECT 0.364 2.084 2.836 2.116 ;
  LAYER M2 ;
        RECT 0.364 2.148 2.836 2.18 ;
  LAYER M2 ;
        RECT 0.364 2.212 2.836 2.244 ;
  LAYER M2 ;
        RECT 0.364 2.276 2.836 2.308 ;
  LAYER M2 ;
        RECT 0.364 2.34 2.836 2.372 ;
  LAYER M2 ;
        RECT 0.364 2.404 2.836 2.436 ;
  LAYER M2 ;
        RECT 0.364 2.468 2.836 2.5 ;
  LAYER M2 ;
        RECT 0.364 2.532 2.836 2.564 ;
  LAYER M2 ;
        RECT 0.364 2.596 2.836 2.628 ;
  LAYER M2 ;
        RECT 0.364 2.66 2.836 2.692 ;
  LAYER M2 ;
        RECT 0.364 2.724 2.836 2.756 ;
  LAYER M2 ;
        RECT 0.364 2.788 2.836 2.82 ;
  LAYER M2 ;
        RECT 0.364 2.852 2.836 2.884 ;
  LAYER M2 ;
        RECT 0.364 2.916 2.836 2.948 ;
  LAYER M2 ;
        RECT 0.364 2.98 2.836 3.012 ;
  LAYER M2 ;
        RECT 0.364 3.044 2.836 3.076 ;
  LAYER M3 ;
        RECT 0.384 0.72 0.416 3.228 ;
  LAYER M3 ;
        RECT 0.448 0.72 0.48 3.228 ;
  LAYER M3 ;
        RECT 0.512 0.72 0.544 3.228 ;
  LAYER M3 ;
        RECT 0.576 0.72 0.608 3.228 ;
  LAYER M3 ;
        RECT 0.64 0.72 0.672 3.228 ;
  LAYER M3 ;
        RECT 0.704 0.72 0.736 3.228 ;
  LAYER M3 ;
        RECT 0.768 0.72 0.8 3.228 ;
  LAYER M3 ;
        RECT 0.832 0.72 0.864 3.228 ;
  LAYER M3 ;
        RECT 0.896 0.72 0.928 3.228 ;
  LAYER M3 ;
        RECT 0.96 0.72 0.992 3.228 ;
  LAYER M3 ;
        RECT 1.024 0.72 1.056 3.228 ;
  LAYER M3 ;
        RECT 1.088 0.72 1.12 3.228 ;
  LAYER M3 ;
        RECT 1.152 0.72 1.184 3.228 ;
  LAYER M3 ;
        RECT 1.216 0.72 1.248 3.228 ;
  LAYER M3 ;
        RECT 1.28 0.72 1.312 3.228 ;
  LAYER M3 ;
        RECT 1.344 0.72 1.376 3.228 ;
  LAYER M3 ;
        RECT 1.408 0.72 1.44 3.228 ;
  LAYER M3 ;
        RECT 1.472 0.72 1.504 3.228 ;
  LAYER M3 ;
        RECT 1.536 0.72 1.568 3.228 ;
  LAYER M3 ;
        RECT 1.6 0.72 1.632 3.228 ;
  LAYER M3 ;
        RECT 1.664 0.72 1.696 3.228 ;
  LAYER M3 ;
        RECT 1.728 0.72 1.76 3.228 ;
  LAYER M3 ;
        RECT 1.792 0.72 1.824 3.228 ;
  LAYER M3 ;
        RECT 1.856 0.72 1.888 3.228 ;
  LAYER M3 ;
        RECT 1.92 0.72 1.952 3.228 ;
  LAYER M3 ;
        RECT 1.984 0.72 2.016 3.228 ;
  LAYER M3 ;
        RECT 2.048 0.72 2.08 3.228 ;
  LAYER M3 ;
        RECT 2.112 0.72 2.144 3.228 ;
  LAYER M3 ;
        RECT 2.176 0.72 2.208 3.228 ;
  LAYER M3 ;
        RECT 2.24 0.72 2.272 3.228 ;
  LAYER M3 ;
        RECT 2.304 0.72 2.336 3.228 ;
  LAYER M3 ;
        RECT 2.368 0.72 2.4 3.228 ;
  LAYER M3 ;
        RECT 2.432 0.72 2.464 3.228 ;
  LAYER M3 ;
        RECT 2.496 0.72 2.528 3.228 ;
  LAYER M3 ;
        RECT 2.56 0.72 2.592 3.228 ;
  LAYER M3 ;
        RECT 2.624 0.72 2.656 3.228 ;
  LAYER M3 ;
        RECT 2.688 0.72 2.72 3.228 ;
  LAYER M3 ;
        RECT 2.784 0.72 2.816 3.228 ;
  LAYER M1 ;
        RECT 0.399 0.756 0.401 3.192 ;
  LAYER M1 ;
        RECT 0.479 0.756 0.481 3.192 ;
  LAYER M1 ;
        RECT 0.559 0.756 0.561 3.192 ;
  LAYER M1 ;
        RECT 0.639 0.756 0.641 3.192 ;
  LAYER M1 ;
        RECT 0.719 0.756 0.721 3.192 ;
  LAYER M1 ;
        RECT 0.799 0.756 0.801 3.192 ;
  LAYER M1 ;
        RECT 0.879 0.756 0.881 3.192 ;
  LAYER M1 ;
        RECT 0.959 0.756 0.961 3.192 ;
  LAYER M1 ;
        RECT 1.039 0.756 1.041 3.192 ;
  LAYER M1 ;
        RECT 1.119 0.756 1.121 3.192 ;
  LAYER M1 ;
        RECT 1.199 0.756 1.201 3.192 ;
  LAYER M1 ;
        RECT 1.279 0.756 1.281 3.192 ;
  LAYER M1 ;
        RECT 1.359 0.756 1.361 3.192 ;
  LAYER M1 ;
        RECT 1.439 0.756 1.441 3.192 ;
  LAYER M1 ;
        RECT 1.519 0.756 1.521 3.192 ;
  LAYER M1 ;
        RECT 1.599 0.756 1.601 3.192 ;
  LAYER M1 ;
        RECT 1.679 0.756 1.681 3.192 ;
  LAYER M1 ;
        RECT 1.759 0.756 1.761 3.192 ;
  LAYER M1 ;
        RECT 1.839 0.756 1.841 3.192 ;
  LAYER M1 ;
        RECT 1.919 0.756 1.921 3.192 ;
  LAYER M1 ;
        RECT 1.999 0.756 2.001 3.192 ;
  LAYER M1 ;
        RECT 2.079 0.756 2.081 3.192 ;
  LAYER M1 ;
        RECT 2.159 0.756 2.161 3.192 ;
  LAYER M1 ;
        RECT 2.239 0.756 2.241 3.192 ;
  LAYER M1 ;
        RECT 2.319 0.756 2.321 3.192 ;
  LAYER M1 ;
        RECT 2.399 0.756 2.401 3.192 ;
  LAYER M1 ;
        RECT 2.479 0.756 2.481 3.192 ;
  LAYER M1 ;
        RECT 2.559 0.756 2.561 3.192 ;
  LAYER M1 ;
        RECT 2.639 0.756 2.641 3.192 ;
  LAYER M1 ;
        RECT 2.719 0.756 2.721 3.192 ;
  LAYER M2 ;
        RECT 0.4 0.755 2.8 0.757 ;
  LAYER M2 ;
        RECT 0.4 0.839 2.8 0.841 ;
  LAYER M2 ;
        RECT 0.4 0.923 2.8 0.925 ;
  LAYER M2 ;
        RECT 0.4 1.007 2.8 1.009 ;
  LAYER M2 ;
        RECT 0.4 1.091 2.8 1.093 ;
  LAYER M2 ;
        RECT 0.4 1.175 2.8 1.177 ;
  LAYER M2 ;
        RECT 0.4 1.259 2.8 1.261 ;
  LAYER M2 ;
        RECT 0.4 1.343 2.8 1.345 ;
  LAYER M2 ;
        RECT 0.4 1.427 2.8 1.429 ;
  LAYER M2 ;
        RECT 0.4 1.511 2.8 1.513 ;
  LAYER M2 ;
        RECT 0.4 1.595 2.8 1.597 ;
  LAYER M2 ;
        RECT 0.4 1.679 2.8 1.681 ;
  LAYER M2 ;
        RECT 0.4 1.7625 2.8 1.7645 ;
  LAYER M2 ;
        RECT 0.4 1.847 2.8 1.849 ;
  LAYER M2 ;
        RECT 0.4 1.931 2.8 1.933 ;
  LAYER M2 ;
        RECT 0.4 2.015 2.8 2.017 ;
  LAYER M2 ;
        RECT 0.4 2.099 2.8 2.101 ;
  LAYER M2 ;
        RECT 0.4 2.183 2.8 2.185 ;
  LAYER M2 ;
        RECT 0.4 2.267 2.8 2.269 ;
  LAYER M2 ;
        RECT 0.4 2.351 2.8 2.353 ;
  LAYER M2 ;
        RECT 0.4 2.435 2.8 2.437 ;
  LAYER M2 ;
        RECT 0.4 2.519 2.8 2.521 ;
  LAYER M2 ;
        RECT 0.4 2.603 2.8 2.605 ;
  LAYER M2 ;
        RECT 0.4 2.687 2.8 2.689 ;
  LAYER M2 ;
        RECT 0.4 2.771 2.8 2.773 ;
  LAYER M2 ;
        RECT 0.4 2.855 2.8 2.857 ;
  LAYER M2 ;
        RECT 0.4 2.939 2.8 2.941 ;
  LAYER M2 ;
        RECT 0.4 3.023 2.8 3.025 ;
  LAYER M2 ;
        RECT 0.4 3.107 2.8 3.109 ;
  LAYER M1 ;
        RECT 0.384 3.66 0.416 6.168 ;
  LAYER M1 ;
        RECT 0.448 3.66 0.48 6.168 ;
  LAYER M1 ;
        RECT 0.512 3.66 0.544 6.168 ;
  LAYER M1 ;
        RECT 0.576 3.66 0.608 6.168 ;
  LAYER M1 ;
        RECT 0.64 3.66 0.672 6.168 ;
  LAYER M1 ;
        RECT 0.704 3.66 0.736 6.168 ;
  LAYER M1 ;
        RECT 0.768 3.66 0.8 6.168 ;
  LAYER M1 ;
        RECT 0.832 3.66 0.864 6.168 ;
  LAYER M1 ;
        RECT 0.896 3.66 0.928 6.168 ;
  LAYER M1 ;
        RECT 0.96 3.66 0.992 6.168 ;
  LAYER M1 ;
        RECT 1.024 3.66 1.056 6.168 ;
  LAYER M1 ;
        RECT 1.088 3.66 1.12 6.168 ;
  LAYER M1 ;
        RECT 1.152 3.66 1.184 6.168 ;
  LAYER M1 ;
        RECT 1.216 3.66 1.248 6.168 ;
  LAYER M1 ;
        RECT 1.28 3.66 1.312 6.168 ;
  LAYER M1 ;
        RECT 1.344 3.66 1.376 6.168 ;
  LAYER M1 ;
        RECT 1.408 3.66 1.44 6.168 ;
  LAYER M1 ;
        RECT 1.472 3.66 1.504 6.168 ;
  LAYER M1 ;
        RECT 1.536 3.66 1.568 6.168 ;
  LAYER M1 ;
        RECT 1.6 3.66 1.632 6.168 ;
  LAYER M1 ;
        RECT 1.664 3.66 1.696 6.168 ;
  LAYER M1 ;
        RECT 1.728 3.66 1.76 6.168 ;
  LAYER M1 ;
        RECT 1.792 3.66 1.824 6.168 ;
  LAYER M1 ;
        RECT 1.856 3.66 1.888 6.168 ;
  LAYER M1 ;
        RECT 1.92 3.66 1.952 6.168 ;
  LAYER M1 ;
        RECT 1.984 3.66 2.016 6.168 ;
  LAYER M1 ;
        RECT 2.048 3.66 2.08 6.168 ;
  LAYER M1 ;
        RECT 2.112 3.66 2.144 6.168 ;
  LAYER M1 ;
        RECT 2.176 3.66 2.208 6.168 ;
  LAYER M1 ;
        RECT 2.24 3.66 2.272 6.168 ;
  LAYER M1 ;
        RECT 2.304 3.66 2.336 6.168 ;
  LAYER M1 ;
        RECT 2.368 3.66 2.4 6.168 ;
  LAYER M1 ;
        RECT 2.432 3.66 2.464 6.168 ;
  LAYER M1 ;
        RECT 2.496 3.66 2.528 6.168 ;
  LAYER M1 ;
        RECT 2.56 3.66 2.592 6.168 ;
  LAYER M1 ;
        RECT 2.624 3.66 2.656 6.168 ;
  LAYER M1 ;
        RECT 2.688 3.66 2.72 6.168 ;
  LAYER M2 ;
        RECT 0.364 3.744 2.836 3.776 ;
  LAYER M2 ;
        RECT 0.364 3.808 2.836 3.84 ;
  LAYER M2 ;
        RECT 0.364 3.872 2.836 3.904 ;
  LAYER M2 ;
        RECT 0.364 3.936 2.836 3.968 ;
  LAYER M2 ;
        RECT 0.364 4 2.836 4.032 ;
  LAYER M2 ;
        RECT 0.364 4.064 2.836 4.096 ;
  LAYER M2 ;
        RECT 0.364 4.128 2.836 4.16 ;
  LAYER M2 ;
        RECT 0.364 4.192 2.836 4.224 ;
  LAYER M2 ;
        RECT 0.364 4.256 2.836 4.288 ;
  LAYER M2 ;
        RECT 0.364 4.32 2.836 4.352 ;
  LAYER M2 ;
        RECT 0.364 4.384 2.836 4.416 ;
  LAYER M2 ;
        RECT 0.364 4.448 2.836 4.48 ;
  LAYER M2 ;
        RECT 0.364 4.512 2.836 4.544 ;
  LAYER M2 ;
        RECT 0.364 4.576 2.836 4.608 ;
  LAYER M2 ;
        RECT 0.364 4.64 2.836 4.672 ;
  LAYER M2 ;
        RECT 0.364 4.704 2.836 4.736 ;
  LAYER M2 ;
        RECT 0.364 4.768 2.836 4.8 ;
  LAYER M2 ;
        RECT 0.364 4.832 2.836 4.864 ;
  LAYER M2 ;
        RECT 0.364 4.896 2.836 4.928 ;
  LAYER M2 ;
        RECT 0.364 4.96 2.836 4.992 ;
  LAYER M2 ;
        RECT 0.364 5.024 2.836 5.056 ;
  LAYER M2 ;
        RECT 0.364 5.088 2.836 5.12 ;
  LAYER M2 ;
        RECT 0.364 5.152 2.836 5.184 ;
  LAYER M2 ;
        RECT 0.364 5.216 2.836 5.248 ;
  LAYER M2 ;
        RECT 0.364 5.28 2.836 5.312 ;
  LAYER M2 ;
        RECT 0.364 5.344 2.836 5.376 ;
  LAYER M2 ;
        RECT 0.364 5.408 2.836 5.44 ;
  LAYER M2 ;
        RECT 0.364 5.472 2.836 5.504 ;
  LAYER M2 ;
        RECT 0.364 5.536 2.836 5.568 ;
  LAYER M2 ;
        RECT 0.364 5.6 2.836 5.632 ;
  LAYER M2 ;
        RECT 0.364 5.664 2.836 5.696 ;
  LAYER M2 ;
        RECT 0.364 5.728 2.836 5.76 ;
  LAYER M2 ;
        RECT 0.364 5.792 2.836 5.824 ;
  LAYER M2 ;
        RECT 0.364 5.856 2.836 5.888 ;
  LAYER M2 ;
        RECT 0.364 5.92 2.836 5.952 ;
  LAYER M2 ;
        RECT 0.364 5.984 2.836 6.016 ;
  LAYER M3 ;
        RECT 0.384 3.66 0.416 6.168 ;
  LAYER M3 ;
        RECT 0.448 3.66 0.48 6.168 ;
  LAYER M3 ;
        RECT 0.512 3.66 0.544 6.168 ;
  LAYER M3 ;
        RECT 0.576 3.66 0.608 6.168 ;
  LAYER M3 ;
        RECT 0.64 3.66 0.672 6.168 ;
  LAYER M3 ;
        RECT 0.704 3.66 0.736 6.168 ;
  LAYER M3 ;
        RECT 0.768 3.66 0.8 6.168 ;
  LAYER M3 ;
        RECT 0.832 3.66 0.864 6.168 ;
  LAYER M3 ;
        RECT 0.896 3.66 0.928 6.168 ;
  LAYER M3 ;
        RECT 0.96 3.66 0.992 6.168 ;
  LAYER M3 ;
        RECT 1.024 3.66 1.056 6.168 ;
  LAYER M3 ;
        RECT 1.088 3.66 1.12 6.168 ;
  LAYER M3 ;
        RECT 1.152 3.66 1.184 6.168 ;
  LAYER M3 ;
        RECT 1.216 3.66 1.248 6.168 ;
  LAYER M3 ;
        RECT 1.28 3.66 1.312 6.168 ;
  LAYER M3 ;
        RECT 1.344 3.66 1.376 6.168 ;
  LAYER M3 ;
        RECT 1.408 3.66 1.44 6.168 ;
  LAYER M3 ;
        RECT 1.472 3.66 1.504 6.168 ;
  LAYER M3 ;
        RECT 1.536 3.66 1.568 6.168 ;
  LAYER M3 ;
        RECT 1.6 3.66 1.632 6.168 ;
  LAYER M3 ;
        RECT 1.664 3.66 1.696 6.168 ;
  LAYER M3 ;
        RECT 1.728 3.66 1.76 6.168 ;
  LAYER M3 ;
        RECT 1.792 3.66 1.824 6.168 ;
  LAYER M3 ;
        RECT 1.856 3.66 1.888 6.168 ;
  LAYER M3 ;
        RECT 1.92 3.66 1.952 6.168 ;
  LAYER M3 ;
        RECT 1.984 3.66 2.016 6.168 ;
  LAYER M3 ;
        RECT 2.048 3.66 2.08 6.168 ;
  LAYER M3 ;
        RECT 2.112 3.66 2.144 6.168 ;
  LAYER M3 ;
        RECT 2.176 3.66 2.208 6.168 ;
  LAYER M3 ;
        RECT 2.24 3.66 2.272 6.168 ;
  LAYER M3 ;
        RECT 2.304 3.66 2.336 6.168 ;
  LAYER M3 ;
        RECT 2.368 3.66 2.4 6.168 ;
  LAYER M3 ;
        RECT 2.432 3.66 2.464 6.168 ;
  LAYER M3 ;
        RECT 2.496 3.66 2.528 6.168 ;
  LAYER M3 ;
        RECT 2.56 3.66 2.592 6.168 ;
  LAYER M3 ;
        RECT 2.624 3.66 2.656 6.168 ;
  LAYER M3 ;
        RECT 2.688 3.66 2.72 6.168 ;
  LAYER M3 ;
        RECT 2.784 3.66 2.816 6.168 ;
  LAYER M1 ;
        RECT 0.399 3.696 0.401 6.132 ;
  LAYER M1 ;
        RECT 0.479 3.696 0.481 6.132 ;
  LAYER M1 ;
        RECT 0.559 3.696 0.561 6.132 ;
  LAYER M1 ;
        RECT 0.639 3.696 0.641 6.132 ;
  LAYER M1 ;
        RECT 0.719 3.696 0.721 6.132 ;
  LAYER M1 ;
        RECT 0.799 3.696 0.801 6.132 ;
  LAYER M1 ;
        RECT 0.879 3.696 0.881 6.132 ;
  LAYER M1 ;
        RECT 0.959 3.696 0.961 6.132 ;
  LAYER M1 ;
        RECT 1.039 3.696 1.041 6.132 ;
  LAYER M1 ;
        RECT 1.119 3.696 1.121 6.132 ;
  LAYER M1 ;
        RECT 1.199 3.696 1.201 6.132 ;
  LAYER M1 ;
        RECT 1.279 3.696 1.281 6.132 ;
  LAYER M1 ;
        RECT 1.359 3.696 1.361 6.132 ;
  LAYER M1 ;
        RECT 1.439 3.696 1.441 6.132 ;
  LAYER M1 ;
        RECT 1.519 3.696 1.521 6.132 ;
  LAYER M1 ;
        RECT 1.599 3.696 1.601 6.132 ;
  LAYER M1 ;
        RECT 1.679 3.696 1.681 6.132 ;
  LAYER M1 ;
        RECT 1.759 3.696 1.761 6.132 ;
  LAYER M1 ;
        RECT 1.839 3.696 1.841 6.132 ;
  LAYER M1 ;
        RECT 1.919 3.696 1.921 6.132 ;
  LAYER M1 ;
        RECT 1.999 3.696 2.001 6.132 ;
  LAYER M1 ;
        RECT 2.079 3.696 2.081 6.132 ;
  LAYER M1 ;
        RECT 2.159 3.696 2.161 6.132 ;
  LAYER M1 ;
        RECT 2.239 3.696 2.241 6.132 ;
  LAYER M1 ;
        RECT 2.319 3.696 2.321 6.132 ;
  LAYER M1 ;
        RECT 2.399 3.696 2.401 6.132 ;
  LAYER M1 ;
        RECT 2.479 3.696 2.481 6.132 ;
  LAYER M1 ;
        RECT 2.559 3.696 2.561 6.132 ;
  LAYER M1 ;
        RECT 2.639 3.696 2.641 6.132 ;
  LAYER M1 ;
        RECT 2.719 3.696 2.721 6.132 ;
  LAYER M2 ;
        RECT 0.4 3.695 2.8 3.697 ;
  LAYER M2 ;
        RECT 0.4 3.779 2.8 3.781 ;
  LAYER M2 ;
        RECT 0.4 3.863 2.8 3.865 ;
  LAYER M2 ;
        RECT 0.4 3.947 2.8 3.949 ;
  LAYER M2 ;
        RECT 0.4 4.031 2.8 4.033 ;
  LAYER M2 ;
        RECT 0.4 4.115 2.8 4.117 ;
  LAYER M2 ;
        RECT 0.4 4.199 2.8 4.201 ;
  LAYER M2 ;
        RECT 0.4 4.283 2.8 4.285 ;
  LAYER M2 ;
        RECT 0.4 4.367 2.8 4.369 ;
  LAYER M2 ;
        RECT 0.4 4.451 2.8 4.453 ;
  LAYER M2 ;
        RECT 0.4 4.535 2.8 4.537 ;
  LAYER M2 ;
        RECT 0.4 4.619 2.8 4.621 ;
  LAYER M2 ;
        RECT 0.4 4.7025 2.8 4.7045 ;
  LAYER M2 ;
        RECT 0.4 4.787 2.8 4.789 ;
  LAYER M2 ;
        RECT 0.4 4.871 2.8 4.873 ;
  LAYER M2 ;
        RECT 0.4 4.955 2.8 4.957 ;
  LAYER M2 ;
        RECT 0.4 5.039 2.8 5.041 ;
  LAYER M2 ;
        RECT 0.4 5.123 2.8 5.125 ;
  LAYER M2 ;
        RECT 0.4 5.207 2.8 5.209 ;
  LAYER M2 ;
        RECT 0.4 5.291 2.8 5.293 ;
  LAYER M2 ;
        RECT 0.4 5.375 2.8 5.377 ;
  LAYER M2 ;
        RECT 0.4 5.459 2.8 5.461 ;
  LAYER M2 ;
        RECT 0.4 5.543 2.8 5.545 ;
  LAYER M2 ;
        RECT 0.4 5.627 2.8 5.629 ;
  LAYER M2 ;
        RECT 0.4 5.711 2.8 5.713 ;
  LAYER M2 ;
        RECT 0.4 5.795 2.8 5.797 ;
  LAYER M2 ;
        RECT 0.4 5.879 2.8 5.881 ;
  LAYER M2 ;
        RECT 0.4 5.963 2.8 5.965 ;
  LAYER M2 ;
        RECT 0.4 6.047 2.8 6.049 ;
  LAYER M1 ;
        RECT 0.384 6.6 0.416 9.108 ;
  LAYER M1 ;
        RECT 0.448 6.6 0.48 9.108 ;
  LAYER M1 ;
        RECT 0.512 6.6 0.544 9.108 ;
  LAYER M1 ;
        RECT 0.576 6.6 0.608 9.108 ;
  LAYER M1 ;
        RECT 0.64 6.6 0.672 9.108 ;
  LAYER M1 ;
        RECT 0.704 6.6 0.736 9.108 ;
  LAYER M1 ;
        RECT 0.768 6.6 0.8 9.108 ;
  LAYER M1 ;
        RECT 0.832 6.6 0.864 9.108 ;
  LAYER M1 ;
        RECT 0.896 6.6 0.928 9.108 ;
  LAYER M1 ;
        RECT 0.96 6.6 0.992 9.108 ;
  LAYER M1 ;
        RECT 1.024 6.6 1.056 9.108 ;
  LAYER M1 ;
        RECT 1.088 6.6 1.12 9.108 ;
  LAYER M1 ;
        RECT 1.152 6.6 1.184 9.108 ;
  LAYER M1 ;
        RECT 1.216 6.6 1.248 9.108 ;
  LAYER M1 ;
        RECT 1.28 6.6 1.312 9.108 ;
  LAYER M1 ;
        RECT 1.344 6.6 1.376 9.108 ;
  LAYER M1 ;
        RECT 1.408 6.6 1.44 9.108 ;
  LAYER M1 ;
        RECT 1.472 6.6 1.504 9.108 ;
  LAYER M1 ;
        RECT 1.536 6.6 1.568 9.108 ;
  LAYER M1 ;
        RECT 1.6 6.6 1.632 9.108 ;
  LAYER M1 ;
        RECT 1.664 6.6 1.696 9.108 ;
  LAYER M1 ;
        RECT 1.728 6.6 1.76 9.108 ;
  LAYER M1 ;
        RECT 1.792 6.6 1.824 9.108 ;
  LAYER M1 ;
        RECT 1.856 6.6 1.888 9.108 ;
  LAYER M1 ;
        RECT 1.92 6.6 1.952 9.108 ;
  LAYER M1 ;
        RECT 1.984 6.6 2.016 9.108 ;
  LAYER M1 ;
        RECT 2.048 6.6 2.08 9.108 ;
  LAYER M1 ;
        RECT 2.112 6.6 2.144 9.108 ;
  LAYER M1 ;
        RECT 2.176 6.6 2.208 9.108 ;
  LAYER M1 ;
        RECT 2.24 6.6 2.272 9.108 ;
  LAYER M1 ;
        RECT 2.304 6.6 2.336 9.108 ;
  LAYER M1 ;
        RECT 2.368 6.6 2.4 9.108 ;
  LAYER M1 ;
        RECT 2.432 6.6 2.464 9.108 ;
  LAYER M1 ;
        RECT 2.496 6.6 2.528 9.108 ;
  LAYER M1 ;
        RECT 2.56 6.6 2.592 9.108 ;
  LAYER M1 ;
        RECT 2.624 6.6 2.656 9.108 ;
  LAYER M1 ;
        RECT 2.688 6.6 2.72 9.108 ;
  LAYER M2 ;
        RECT 0.364 6.684 2.836 6.716 ;
  LAYER M2 ;
        RECT 0.364 6.748 2.836 6.78 ;
  LAYER M2 ;
        RECT 0.364 6.812 2.836 6.844 ;
  LAYER M2 ;
        RECT 0.364 6.876 2.836 6.908 ;
  LAYER M2 ;
        RECT 0.364 6.94 2.836 6.972 ;
  LAYER M2 ;
        RECT 0.364 7.004 2.836 7.036 ;
  LAYER M2 ;
        RECT 0.364 7.068 2.836 7.1 ;
  LAYER M2 ;
        RECT 0.364 7.132 2.836 7.164 ;
  LAYER M2 ;
        RECT 0.364 7.196 2.836 7.228 ;
  LAYER M2 ;
        RECT 0.364 7.26 2.836 7.292 ;
  LAYER M2 ;
        RECT 0.364 7.324 2.836 7.356 ;
  LAYER M2 ;
        RECT 0.364 7.388 2.836 7.42 ;
  LAYER M2 ;
        RECT 0.364 7.452 2.836 7.484 ;
  LAYER M2 ;
        RECT 0.364 7.516 2.836 7.548 ;
  LAYER M2 ;
        RECT 0.364 7.58 2.836 7.612 ;
  LAYER M2 ;
        RECT 0.364 7.644 2.836 7.676 ;
  LAYER M2 ;
        RECT 0.364 7.708 2.836 7.74 ;
  LAYER M2 ;
        RECT 0.364 7.772 2.836 7.804 ;
  LAYER M2 ;
        RECT 0.364 7.836 2.836 7.868 ;
  LAYER M2 ;
        RECT 0.364 7.9 2.836 7.932 ;
  LAYER M2 ;
        RECT 0.364 7.964 2.836 7.996 ;
  LAYER M2 ;
        RECT 0.364 8.028 2.836 8.06 ;
  LAYER M2 ;
        RECT 0.364 8.092 2.836 8.124 ;
  LAYER M2 ;
        RECT 0.364 8.156 2.836 8.188 ;
  LAYER M2 ;
        RECT 0.364 8.22 2.836 8.252 ;
  LAYER M2 ;
        RECT 0.364 8.284 2.836 8.316 ;
  LAYER M2 ;
        RECT 0.364 8.348 2.836 8.38 ;
  LAYER M2 ;
        RECT 0.364 8.412 2.836 8.444 ;
  LAYER M2 ;
        RECT 0.364 8.476 2.836 8.508 ;
  LAYER M2 ;
        RECT 0.364 8.54 2.836 8.572 ;
  LAYER M2 ;
        RECT 0.364 8.604 2.836 8.636 ;
  LAYER M2 ;
        RECT 0.364 8.668 2.836 8.7 ;
  LAYER M2 ;
        RECT 0.364 8.732 2.836 8.764 ;
  LAYER M2 ;
        RECT 0.364 8.796 2.836 8.828 ;
  LAYER M2 ;
        RECT 0.364 8.86 2.836 8.892 ;
  LAYER M2 ;
        RECT 0.364 8.924 2.836 8.956 ;
  LAYER M3 ;
        RECT 0.384 6.6 0.416 9.108 ;
  LAYER M3 ;
        RECT 0.448 6.6 0.48 9.108 ;
  LAYER M3 ;
        RECT 0.512 6.6 0.544 9.108 ;
  LAYER M3 ;
        RECT 0.576 6.6 0.608 9.108 ;
  LAYER M3 ;
        RECT 0.64 6.6 0.672 9.108 ;
  LAYER M3 ;
        RECT 0.704 6.6 0.736 9.108 ;
  LAYER M3 ;
        RECT 0.768 6.6 0.8 9.108 ;
  LAYER M3 ;
        RECT 0.832 6.6 0.864 9.108 ;
  LAYER M3 ;
        RECT 0.896 6.6 0.928 9.108 ;
  LAYER M3 ;
        RECT 0.96 6.6 0.992 9.108 ;
  LAYER M3 ;
        RECT 1.024 6.6 1.056 9.108 ;
  LAYER M3 ;
        RECT 1.088 6.6 1.12 9.108 ;
  LAYER M3 ;
        RECT 1.152 6.6 1.184 9.108 ;
  LAYER M3 ;
        RECT 1.216 6.6 1.248 9.108 ;
  LAYER M3 ;
        RECT 1.28 6.6 1.312 9.108 ;
  LAYER M3 ;
        RECT 1.344 6.6 1.376 9.108 ;
  LAYER M3 ;
        RECT 1.408 6.6 1.44 9.108 ;
  LAYER M3 ;
        RECT 1.472 6.6 1.504 9.108 ;
  LAYER M3 ;
        RECT 1.536 6.6 1.568 9.108 ;
  LAYER M3 ;
        RECT 1.6 6.6 1.632 9.108 ;
  LAYER M3 ;
        RECT 1.664 6.6 1.696 9.108 ;
  LAYER M3 ;
        RECT 1.728 6.6 1.76 9.108 ;
  LAYER M3 ;
        RECT 1.792 6.6 1.824 9.108 ;
  LAYER M3 ;
        RECT 1.856 6.6 1.888 9.108 ;
  LAYER M3 ;
        RECT 1.92 6.6 1.952 9.108 ;
  LAYER M3 ;
        RECT 1.984 6.6 2.016 9.108 ;
  LAYER M3 ;
        RECT 2.048 6.6 2.08 9.108 ;
  LAYER M3 ;
        RECT 2.112 6.6 2.144 9.108 ;
  LAYER M3 ;
        RECT 2.176 6.6 2.208 9.108 ;
  LAYER M3 ;
        RECT 2.24 6.6 2.272 9.108 ;
  LAYER M3 ;
        RECT 2.304 6.6 2.336 9.108 ;
  LAYER M3 ;
        RECT 2.368 6.6 2.4 9.108 ;
  LAYER M3 ;
        RECT 2.432 6.6 2.464 9.108 ;
  LAYER M3 ;
        RECT 2.496 6.6 2.528 9.108 ;
  LAYER M3 ;
        RECT 2.56 6.6 2.592 9.108 ;
  LAYER M3 ;
        RECT 2.624 6.6 2.656 9.108 ;
  LAYER M3 ;
        RECT 2.688 6.6 2.72 9.108 ;
  LAYER M3 ;
        RECT 2.784 6.6 2.816 9.108 ;
  LAYER M1 ;
        RECT 0.399 6.636 0.401 9.072 ;
  LAYER M1 ;
        RECT 0.479 6.636 0.481 9.072 ;
  LAYER M1 ;
        RECT 0.559 6.636 0.561 9.072 ;
  LAYER M1 ;
        RECT 0.639 6.636 0.641 9.072 ;
  LAYER M1 ;
        RECT 0.719 6.636 0.721 9.072 ;
  LAYER M1 ;
        RECT 0.799 6.636 0.801 9.072 ;
  LAYER M1 ;
        RECT 0.879 6.636 0.881 9.072 ;
  LAYER M1 ;
        RECT 0.959 6.636 0.961 9.072 ;
  LAYER M1 ;
        RECT 1.039 6.636 1.041 9.072 ;
  LAYER M1 ;
        RECT 1.119 6.636 1.121 9.072 ;
  LAYER M1 ;
        RECT 1.199 6.636 1.201 9.072 ;
  LAYER M1 ;
        RECT 1.279 6.636 1.281 9.072 ;
  LAYER M1 ;
        RECT 1.359 6.636 1.361 9.072 ;
  LAYER M1 ;
        RECT 1.439 6.636 1.441 9.072 ;
  LAYER M1 ;
        RECT 1.519 6.636 1.521 9.072 ;
  LAYER M1 ;
        RECT 1.599 6.636 1.601 9.072 ;
  LAYER M1 ;
        RECT 1.679 6.636 1.681 9.072 ;
  LAYER M1 ;
        RECT 1.759 6.636 1.761 9.072 ;
  LAYER M1 ;
        RECT 1.839 6.636 1.841 9.072 ;
  LAYER M1 ;
        RECT 1.919 6.636 1.921 9.072 ;
  LAYER M1 ;
        RECT 1.999 6.636 2.001 9.072 ;
  LAYER M1 ;
        RECT 2.079 6.636 2.081 9.072 ;
  LAYER M1 ;
        RECT 2.159 6.636 2.161 9.072 ;
  LAYER M1 ;
        RECT 2.239 6.636 2.241 9.072 ;
  LAYER M1 ;
        RECT 2.319 6.636 2.321 9.072 ;
  LAYER M1 ;
        RECT 2.399 6.636 2.401 9.072 ;
  LAYER M1 ;
        RECT 2.479 6.636 2.481 9.072 ;
  LAYER M1 ;
        RECT 2.559 6.636 2.561 9.072 ;
  LAYER M1 ;
        RECT 2.639 6.636 2.641 9.072 ;
  LAYER M1 ;
        RECT 2.719 6.636 2.721 9.072 ;
  LAYER M2 ;
        RECT 0.4 6.635 2.8 6.637 ;
  LAYER M2 ;
        RECT 0.4 6.719 2.8 6.721 ;
  LAYER M2 ;
        RECT 0.4 6.803 2.8 6.805 ;
  LAYER M2 ;
        RECT 0.4 6.887 2.8 6.889 ;
  LAYER M2 ;
        RECT 0.4 6.971 2.8 6.973 ;
  LAYER M2 ;
        RECT 0.4 7.055 2.8 7.057 ;
  LAYER M2 ;
        RECT 0.4 7.139 2.8 7.141 ;
  LAYER M2 ;
        RECT 0.4 7.223 2.8 7.225 ;
  LAYER M2 ;
        RECT 0.4 7.307 2.8 7.309 ;
  LAYER M2 ;
        RECT 0.4 7.391 2.8 7.393 ;
  LAYER M2 ;
        RECT 0.4 7.475 2.8 7.477 ;
  LAYER M2 ;
        RECT 0.4 7.559 2.8 7.561 ;
  LAYER M2 ;
        RECT 0.4 7.6425 2.8 7.6445 ;
  LAYER M2 ;
        RECT 0.4 7.727 2.8 7.729 ;
  LAYER M2 ;
        RECT 0.4 7.811 2.8 7.813 ;
  LAYER M2 ;
        RECT 0.4 7.895 2.8 7.897 ;
  LAYER M2 ;
        RECT 0.4 7.979 2.8 7.981 ;
  LAYER M2 ;
        RECT 0.4 8.063 2.8 8.065 ;
  LAYER M2 ;
        RECT 0.4 8.147 2.8 8.149 ;
  LAYER M2 ;
        RECT 0.4 8.231 2.8 8.233 ;
  LAYER M2 ;
        RECT 0.4 8.315 2.8 8.317 ;
  LAYER M2 ;
        RECT 0.4 8.399 2.8 8.401 ;
  LAYER M2 ;
        RECT 0.4 8.483 2.8 8.485 ;
  LAYER M2 ;
        RECT 0.4 8.567 2.8 8.569 ;
  LAYER M2 ;
        RECT 0.4 8.651 2.8 8.653 ;
  LAYER M2 ;
        RECT 0.4 8.735 2.8 8.737 ;
  LAYER M2 ;
        RECT 0.4 8.819 2.8 8.821 ;
  LAYER M2 ;
        RECT 0.4 8.903 2.8 8.905 ;
  LAYER M2 ;
        RECT 0.4 8.987 2.8 8.989 ;
  LAYER M1 ;
        RECT 0.384 9.54 0.416 12.048 ;
  LAYER M1 ;
        RECT 0.448 9.54 0.48 12.048 ;
  LAYER M1 ;
        RECT 0.512 9.54 0.544 12.048 ;
  LAYER M1 ;
        RECT 0.576 9.54 0.608 12.048 ;
  LAYER M1 ;
        RECT 0.64 9.54 0.672 12.048 ;
  LAYER M1 ;
        RECT 0.704 9.54 0.736 12.048 ;
  LAYER M1 ;
        RECT 0.768 9.54 0.8 12.048 ;
  LAYER M1 ;
        RECT 0.832 9.54 0.864 12.048 ;
  LAYER M1 ;
        RECT 0.896 9.54 0.928 12.048 ;
  LAYER M1 ;
        RECT 0.96 9.54 0.992 12.048 ;
  LAYER M1 ;
        RECT 1.024 9.54 1.056 12.048 ;
  LAYER M1 ;
        RECT 1.088 9.54 1.12 12.048 ;
  LAYER M1 ;
        RECT 1.152 9.54 1.184 12.048 ;
  LAYER M1 ;
        RECT 1.216 9.54 1.248 12.048 ;
  LAYER M1 ;
        RECT 1.28 9.54 1.312 12.048 ;
  LAYER M1 ;
        RECT 1.344 9.54 1.376 12.048 ;
  LAYER M1 ;
        RECT 1.408 9.54 1.44 12.048 ;
  LAYER M1 ;
        RECT 1.472 9.54 1.504 12.048 ;
  LAYER M1 ;
        RECT 1.536 9.54 1.568 12.048 ;
  LAYER M1 ;
        RECT 1.6 9.54 1.632 12.048 ;
  LAYER M1 ;
        RECT 1.664 9.54 1.696 12.048 ;
  LAYER M1 ;
        RECT 1.728 9.54 1.76 12.048 ;
  LAYER M1 ;
        RECT 1.792 9.54 1.824 12.048 ;
  LAYER M1 ;
        RECT 1.856 9.54 1.888 12.048 ;
  LAYER M1 ;
        RECT 1.92 9.54 1.952 12.048 ;
  LAYER M1 ;
        RECT 1.984 9.54 2.016 12.048 ;
  LAYER M1 ;
        RECT 2.048 9.54 2.08 12.048 ;
  LAYER M1 ;
        RECT 2.112 9.54 2.144 12.048 ;
  LAYER M1 ;
        RECT 2.176 9.54 2.208 12.048 ;
  LAYER M1 ;
        RECT 2.24 9.54 2.272 12.048 ;
  LAYER M1 ;
        RECT 2.304 9.54 2.336 12.048 ;
  LAYER M1 ;
        RECT 2.368 9.54 2.4 12.048 ;
  LAYER M1 ;
        RECT 2.432 9.54 2.464 12.048 ;
  LAYER M1 ;
        RECT 2.496 9.54 2.528 12.048 ;
  LAYER M1 ;
        RECT 2.56 9.54 2.592 12.048 ;
  LAYER M1 ;
        RECT 2.624 9.54 2.656 12.048 ;
  LAYER M1 ;
        RECT 2.688 9.54 2.72 12.048 ;
  LAYER M2 ;
        RECT 0.364 9.624 2.836 9.656 ;
  LAYER M2 ;
        RECT 0.364 9.688 2.836 9.72 ;
  LAYER M2 ;
        RECT 0.364 9.752 2.836 9.784 ;
  LAYER M2 ;
        RECT 0.364 9.816 2.836 9.848 ;
  LAYER M2 ;
        RECT 0.364 9.88 2.836 9.912 ;
  LAYER M2 ;
        RECT 0.364 9.944 2.836 9.976 ;
  LAYER M2 ;
        RECT 0.364 10.008 2.836 10.04 ;
  LAYER M2 ;
        RECT 0.364 10.072 2.836 10.104 ;
  LAYER M2 ;
        RECT 0.364 10.136 2.836 10.168 ;
  LAYER M2 ;
        RECT 0.364 10.2 2.836 10.232 ;
  LAYER M2 ;
        RECT 0.364 10.264 2.836 10.296 ;
  LAYER M2 ;
        RECT 0.364 10.328 2.836 10.36 ;
  LAYER M2 ;
        RECT 0.364 10.392 2.836 10.424 ;
  LAYER M2 ;
        RECT 0.364 10.456 2.836 10.488 ;
  LAYER M2 ;
        RECT 0.364 10.52 2.836 10.552 ;
  LAYER M2 ;
        RECT 0.364 10.584 2.836 10.616 ;
  LAYER M2 ;
        RECT 0.364 10.648 2.836 10.68 ;
  LAYER M2 ;
        RECT 0.364 10.712 2.836 10.744 ;
  LAYER M2 ;
        RECT 0.364 10.776 2.836 10.808 ;
  LAYER M2 ;
        RECT 0.364 10.84 2.836 10.872 ;
  LAYER M2 ;
        RECT 0.364 10.904 2.836 10.936 ;
  LAYER M2 ;
        RECT 0.364 10.968 2.836 11 ;
  LAYER M2 ;
        RECT 0.364 11.032 2.836 11.064 ;
  LAYER M2 ;
        RECT 0.364 11.096 2.836 11.128 ;
  LAYER M2 ;
        RECT 0.364 11.16 2.836 11.192 ;
  LAYER M2 ;
        RECT 0.364 11.224 2.836 11.256 ;
  LAYER M2 ;
        RECT 0.364 11.288 2.836 11.32 ;
  LAYER M2 ;
        RECT 0.364 11.352 2.836 11.384 ;
  LAYER M2 ;
        RECT 0.364 11.416 2.836 11.448 ;
  LAYER M2 ;
        RECT 0.364 11.48 2.836 11.512 ;
  LAYER M2 ;
        RECT 0.364 11.544 2.836 11.576 ;
  LAYER M2 ;
        RECT 0.364 11.608 2.836 11.64 ;
  LAYER M2 ;
        RECT 0.364 11.672 2.836 11.704 ;
  LAYER M2 ;
        RECT 0.364 11.736 2.836 11.768 ;
  LAYER M2 ;
        RECT 0.364 11.8 2.836 11.832 ;
  LAYER M2 ;
        RECT 0.364 11.864 2.836 11.896 ;
  LAYER M3 ;
        RECT 0.384 9.54 0.416 12.048 ;
  LAYER M3 ;
        RECT 0.448 9.54 0.48 12.048 ;
  LAYER M3 ;
        RECT 0.512 9.54 0.544 12.048 ;
  LAYER M3 ;
        RECT 0.576 9.54 0.608 12.048 ;
  LAYER M3 ;
        RECT 0.64 9.54 0.672 12.048 ;
  LAYER M3 ;
        RECT 0.704 9.54 0.736 12.048 ;
  LAYER M3 ;
        RECT 0.768 9.54 0.8 12.048 ;
  LAYER M3 ;
        RECT 0.832 9.54 0.864 12.048 ;
  LAYER M3 ;
        RECT 0.896 9.54 0.928 12.048 ;
  LAYER M3 ;
        RECT 0.96 9.54 0.992 12.048 ;
  LAYER M3 ;
        RECT 1.024 9.54 1.056 12.048 ;
  LAYER M3 ;
        RECT 1.088 9.54 1.12 12.048 ;
  LAYER M3 ;
        RECT 1.152 9.54 1.184 12.048 ;
  LAYER M3 ;
        RECT 1.216 9.54 1.248 12.048 ;
  LAYER M3 ;
        RECT 1.28 9.54 1.312 12.048 ;
  LAYER M3 ;
        RECT 1.344 9.54 1.376 12.048 ;
  LAYER M3 ;
        RECT 1.408 9.54 1.44 12.048 ;
  LAYER M3 ;
        RECT 1.472 9.54 1.504 12.048 ;
  LAYER M3 ;
        RECT 1.536 9.54 1.568 12.048 ;
  LAYER M3 ;
        RECT 1.6 9.54 1.632 12.048 ;
  LAYER M3 ;
        RECT 1.664 9.54 1.696 12.048 ;
  LAYER M3 ;
        RECT 1.728 9.54 1.76 12.048 ;
  LAYER M3 ;
        RECT 1.792 9.54 1.824 12.048 ;
  LAYER M3 ;
        RECT 1.856 9.54 1.888 12.048 ;
  LAYER M3 ;
        RECT 1.92 9.54 1.952 12.048 ;
  LAYER M3 ;
        RECT 1.984 9.54 2.016 12.048 ;
  LAYER M3 ;
        RECT 2.048 9.54 2.08 12.048 ;
  LAYER M3 ;
        RECT 2.112 9.54 2.144 12.048 ;
  LAYER M3 ;
        RECT 2.176 9.54 2.208 12.048 ;
  LAYER M3 ;
        RECT 2.24 9.54 2.272 12.048 ;
  LAYER M3 ;
        RECT 2.304 9.54 2.336 12.048 ;
  LAYER M3 ;
        RECT 2.368 9.54 2.4 12.048 ;
  LAYER M3 ;
        RECT 2.432 9.54 2.464 12.048 ;
  LAYER M3 ;
        RECT 2.496 9.54 2.528 12.048 ;
  LAYER M3 ;
        RECT 2.56 9.54 2.592 12.048 ;
  LAYER M3 ;
        RECT 2.624 9.54 2.656 12.048 ;
  LAYER M3 ;
        RECT 2.688 9.54 2.72 12.048 ;
  LAYER M3 ;
        RECT 2.784 9.54 2.816 12.048 ;
  LAYER M1 ;
        RECT 0.399 9.576 0.401 12.012 ;
  LAYER M1 ;
        RECT 0.479 9.576 0.481 12.012 ;
  LAYER M1 ;
        RECT 0.559 9.576 0.561 12.012 ;
  LAYER M1 ;
        RECT 0.639 9.576 0.641 12.012 ;
  LAYER M1 ;
        RECT 0.719 9.576 0.721 12.012 ;
  LAYER M1 ;
        RECT 0.799 9.576 0.801 12.012 ;
  LAYER M1 ;
        RECT 0.879 9.576 0.881 12.012 ;
  LAYER M1 ;
        RECT 0.959 9.576 0.961 12.012 ;
  LAYER M1 ;
        RECT 1.039 9.576 1.041 12.012 ;
  LAYER M1 ;
        RECT 1.119 9.576 1.121 12.012 ;
  LAYER M1 ;
        RECT 1.199 9.576 1.201 12.012 ;
  LAYER M1 ;
        RECT 1.279 9.576 1.281 12.012 ;
  LAYER M1 ;
        RECT 1.359 9.576 1.361 12.012 ;
  LAYER M1 ;
        RECT 1.439 9.576 1.441 12.012 ;
  LAYER M1 ;
        RECT 1.519 9.576 1.521 12.012 ;
  LAYER M1 ;
        RECT 1.599 9.576 1.601 12.012 ;
  LAYER M1 ;
        RECT 1.679 9.576 1.681 12.012 ;
  LAYER M1 ;
        RECT 1.759 9.576 1.761 12.012 ;
  LAYER M1 ;
        RECT 1.839 9.576 1.841 12.012 ;
  LAYER M1 ;
        RECT 1.919 9.576 1.921 12.012 ;
  LAYER M1 ;
        RECT 1.999 9.576 2.001 12.012 ;
  LAYER M1 ;
        RECT 2.079 9.576 2.081 12.012 ;
  LAYER M1 ;
        RECT 2.159 9.576 2.161 12.012 ;
  LAYER M1 ;
        RECT 2.239 9.576 2.241 12.012 ;
  LAYER M1 ;
        RECT 2.319 9.576 2.321 12.012 ;
  LAYER M1 ;
        RECT 2.399 9.576 2.401 12.012 ;
  LAYER M1 ;
        RECT 2.479 9.576 2.481 12.012 ;
  LAYER M1 ;
        RECT 2.559 9.576 2.561 12.012 ;
  LAYER M1 ;
        RECT 2.639 9.576 2.641 12.012 ;
  LAYER M1 ;
        RECT 2.719 9.576 2.721 12.012 ;
  LAYER M2 ;
        RECT 0.4 9.575 2.8 9.577 ;
  LAYER M2 ;
        RECT 0.4 9.659 2.8 9.661 ;
  LAYER M2 ;
        RECT 0.4 9.743 2.8 9.745 ;
  LAYER M2 ;
        RECT 0.4 9.827 2.8 9.829 ;
  LAYER M2 ;
        RECT 0.4 9.911 2.8 9.913 ;
  LAYER M2 ;
        RECT 0.4 9.995 2.8 9.997 ;
  LAYER M2 ;
        RECT 0.4 10.079 2.8 10.081 ;
  LAYER M2 ;
        RECT 0.4 10.163 2.8 10.165 ;
  LAYER M2 ;
        RECT 0.4 10.247 2.8 10.249 ;
  LAYER M2 ;
        RECT 0.4 10.331 2.8 10.333 ;
  LAYER M2 ;
        RECT 0.4 10.415 2.8 10.417 ;
  LAYER M2 ;
        RECT 0.4 10.499 2.8 10.501 ;
  LAYER M2 ;
        RECT 0.4 10.5825 2.8 10.5845 ;
  LAYER M2 ;
        RECT 0.4 10.667 2.8 10.669 ;
  LAYER M2 ;
        RECT 0.4 10.751 2.8 10.753 ;
  LAYER M2 ;
        RECT 0.4 10.835 2.8 10.837 ;
  LAYER M2 ;
        RECT 0.4 10.919 2.8 10.921 ;
  LAYER M2 ;
        RECT 0.4 11.003 2.8 11.005 ;
  LAYER M2 ;
        RECT 0.4 11.087 2.8 11.089 ;
  LAYER M2 ;
        RECT 0.4 11.171 2.8 11.173 ;
  LAYER M2 ;
        RECT 0.4 11.255 2.8 11.257 ;
  LAYER M2 ;
        RECT 0.4 11.339 2.8 11.341 ;
  LAYER M2 ;
        RECT 0.4 11.423 2.8 11.425 ;
  LAYER M2 ;
        RECT 0.4 11.507 2.8 11.509 ;
  LAYER M2 ;
        RECT 0.4 11.591 2.8 11.593 ;
  LAYER M2 ;
        RECT 0.4 11.675 2.8 11.677 ;
  LAYER M2 ;
        RECT 0.4 11.759 2.8 11.761 ;
  LAYER M2 ;
        RECT 0.4 11.843 2.8 11.845 ;
  LAYER M2 ;
        RECT 0.4 11.927 2.8 11.929 ;
  LAYER M1 ;
        RECT 0.384 12.48 0.416 14.988 ;
  LAYER M1 ;
        RECT 0.448 12.48 0.48 14.988 ;
  LAYER M1 ;
        RECT 0.512 12.48 0.544 14.988 ;
  LAYER M1 ;
        RECT 0.576 12.48 0.608 14.988 ;
  LAYER M1 ;
        RECT 0.64 12.48 0.672 14.988 ;
  LAYER M1 ;
        RECT 0.704 12.48 0.736 14.988 ;
  LAYER M1 ;
        RECT 0.768 12.48 0.8 14.988 ;
  LAYER M1 ;
        RECT 0.832 12.48 0.864 14.988 ;
  LAYER M1 ;
        RECT 0.896 12.48 0.928 14.988 ;
  LAYER M1 ;
        RECT 0.96 12.48 0.992 14.988 ;
  LAYER M1 ;
        RECT 1.024 12.48 1.056 14.988 ;
  LAYER M1 ;
        RECT 1.088 12.48 1.12 14.988 ;
  LAYER M1 ;
        RECT 1.152 12.48 1.184 14.988 ;
  LAYER M1 ;
        RECT 1.216 12.48 1.248 14.988 ;
  LAYER M1 ;
        RECT 1.28 12.48 1.312 14.988 ;
  LAYER M1 ;
        RECT 1.344 12.48 1.376 14.988 ;
  LAYER M1 ;
        RECT 1.408 12.48 1.44 14.988 ;
  LAYER M1 ;
        RECT 1.472 12.48 1.504 14.988 ;
  LAYER M1 ;
        RECT 1.536 12.48 1.568 14.988 ;
  LAYER M1 ;
        RECT 1.6 12.48 1.632 14.988 ;
  LAYER M1 ;
        RECT 1.664 12.48 1.696 14.988 ;
  LAYER M1 ;
        RECT 1.728 12.48 1.76 14.988 ;
  LAYER M1 ;
        RECT 1.792 12.48 1.824 14.988 ;
  LAYER M1 ;
        RECT 1.856 12.48 1.888 14.988 ;
  LAYER M1 ;
        RECT 1.92 12.48 1.952 14.988 ;
  LAYER M1 ;
        RECT 1.984 12.48 2.016 14.988 ;
  LAYER M1 ;
        RECT 2.048 12.48 2.08 14.988 ;
  LAYER M1 ;
        RECT 2.112 12.48 2.144 14.988 ;
  LAYER M1 ;
        RECT 2.176 12.48 2.208 14.988 ;
  LAYER M1 ;
        RECT 2.24 12.48 2.272 14.988 ;
  LAYER M1 ;
        RECT 2.304 12.48 2.336 14.988 ;
  LAYER M1 ;
        RECT 2.368 12.48 2.4 14.988 ;
  LAYER M1 ;
        RECT 2.432 12.48 2.464 14.988 ;
  LAYER M1 ;
        RECT 2.496 12.48 2.528 14.988 ;
  LAYER M1 ;
        RECT 2.56 12.48 2.592 14.988 ;
  LAYER M1 ;
        RECT 2.624 12.48 2.656 14.988 ;
  LAYER M1 ;
        RECT 2.688 12.48 2.72 14.988 ;
  LAYER M2 ;
        RECT 0.364 12.564 2.836 12.596 ;
  LAYER M2 ;
        RECT 0.364 12.628 2.836 12.66 ;
  LAYER M2 ;
        RECT 0.364 12.692 2.836 12.724 ;
  LAYER M2 ;
        RECT 0.364 12.756 2.836 12.788 ;
  LAYER M2 ;
        RECT 0.364 12.82 2.836 12.852 ;
  LAYER M2 ;
        RECT 0.364 12.884 2.836 12.916 ;
  LAYER M2 ;
        RECT 0.364 12.948 2.836 12.98 ;
  LAYER M2 ;
        RECT 0.364 13.012 2.836 13.044 ;
  LAYER M2 ;
        RECT 0.364 13.076 2.836 13.108 ;
  LAYER M2 ;
        RECT 0.364 13.14 2.836 13.172 ;
  LAYER M2 ;
        RECT 0.364 13.204 2.836 13.236 ;
  LAYER M2 ;
        RECT 0.364 13.268 2.836 13.3 ;
  LAYER M2 ;
        RECT 0.364 13.332 2.836 13.364 ;
  LAYER M2 ;
        RECT 0.364 13.396 2.836 13.428 ;
  LAYER M2 ;
        RECT 0.364 13.46 2.836 13.492 ;
  LAYER M2 ;
        RECT 0.364 13.524 2.836 13.556 ;
  LAYER M2 ;
        RECT 0.364 13.588 2.836 13.62 ;
  LAYER M2 ;
        RECT 0.364 13.652 2.836 13.684 ;
  LAYER M2 ;
        RECT 0.364 13.716 2.836 13.748 ;
  LAYER M2 ;
        RECT 0.364 13.78 2.836 13.812 ;
  LAYER M2 ;
        RECT 0.364 13.844 2.836 13.876 ;
  LAYER M2 ;
        RECT 0.364 13.908 2.836 13.94 ;
  LAYER M2 ;
        RECT 0.364 13.972 2.836 14.004 ;
  LAYER M2 ;
        RECT 0.364 14.036 2.836 14.068 ;
  LAYER M2 ;
        RECT 0.364 14.1 2.836 14.132 ;
  LAYER M2 ;
        RECT 0.364 14.164 2.836 14.196 ;
  LAYER M2 ;
        RECT 0.364 14.228 2.836 14.26 ;
  LAYER M2 ;
        RECT 0.364 14.292 2.836 14.324 ;
  LAYER M2 ;
        RECT 0.364 14.356 2.836 14.388 ;
  LAYER M2 ;
        RECT 0.364 14.42 2.836 14.452 ;
  LAYER M2 ;
        RECT 0.364 14.484 2.836 14.516 ;
  LAYER M2 ;
        RECT 0.364 14.548 2.836 14.58 ;
  LAYER M2 ;
        RECT 0.364 14.612 2.836 14.644 ;
  LAYER M2 ;
        RECT 0.364 14.676 2.836 14.708 ;
  LAYER M2 ;
        RECT 0.364 14.74 2.836 14.772 ;
  LAYER M2 ;
        RECT 0.364 14.804 2.836 14.836 ;
  LAYER M3 ;
        RECT 0.384 12.48 0.416 14.988 ;
  LAYER M3 ;
        RECT 0.448 12.48 0.48 14.988 ;
  LAYER M3 ;
        RECT 0.512 12.48 0.544 14.988 ;
  LAYER M3 ;
        RECT 0.576 12.48 0.608 14.988 ;
  LAYER M3 ;
        RECT 0.64 12.48 0.672 14.988 ;
  LAYER M3 ;
        RECT 0.704 12.48 0.736 14.988 ;
  LAYER M3 ;
        RECT 0.768 12.48 0.8 14.988 ;
  LAYER M3 ;
        RECT 0.832 12.48 0.864 14.988 ;
  LAYER M3 ;
        RECT 0.896 12.48 0.928 14.988 ;
  LAYER M3 ;
        RECT 0.96 12.48 0.992 14.988 ;
  LAYER M3 ;
        RECT 1.024 12.48 1.056 14.988 ;
  LAYER M3 ;
        RECT 1.088 12.48 1.12 14.988 ;
  LAYER M3 ;
        RECT 1.152 12.48 1.184 14.988 ;
  LAYER M3 ;
        RECT 1.216 12.48 1.248 14.988 ;
  LAYER M3 ;
        RECT 1.28 12.48 1.312 14.988 ;
  LAYER M3 ;
        RECT 1.344 12.48 1.376 14.988 ;
  LAYER M3 ;
        RECT 1.408 12.48 1.44 14.988 ;
  LAYER M3 ;
        RECT 1.472 12.48 1.504 14.988 ;
  LAYER M3 ;
        RECT 1.536 12.48 1.568 14.988 ;
  LAYER M3 ;
        RECT 1.6 12.48 1.632 14.988 ;
  LAYER M3 ;
        RECT 1.664 12.48 1.696 14.988 ;
  LAYER M3 ;
        RECT 1.728 12.48 1.76 14.988 ;
  LAYER M3 ;
        RECT 1.792 12.48 1.824 14.988 ;
  LAYER M3 ;
        RECT 1.856 12.48 1.888 14.988 ;
  LAYER M3 ;
        RECT 1.92 12.48 1.952 14.988 ;
  LAYER M3 ;
        RECT 1.984 12.48 2.016 14.988 ;
  LAYER M3 ;
        RECT 2.048 12.48 2.08 14.988 ;
  LAYER M3 ;
        RECT 2.112 12.48 2.144 14.988 ;
  LAYER M3 ;
        RECT 2.176 12.48 2.208 14.988 ;
  LAYER M3 ;
        RECT 2.24 12.48 2.272 14.988 ;
  LAYER M3 ;
        RECT 2.304 12.48 2.336 14.988 ;
  LAYER M3 ;
        RECT 2.368 12.48 2.4 14.988 ;
  LAYER M3 ;
        RECT 2.432 12.48 2.464 14.988 ;
  LAYER M3 ;
        RECT 2.496 12.48 2.528 14.988 ;
  LAYER M3 ;
        RECT 2.56 12.48 2.592 14.988 ;
  LAYER M3 ;
        RECT 2.624 12.48 2.656 14.988 ;
  LAYER M3 ;
        RECT 2.688 12.48 2.72 14.988 ;
  LAYER M3 ;
        RECT 2.784 12.48 2.816 14.988 ;
  LAYER M1 ;
        RECT 0.399 12.516 0.401 14.952 ;
  LAYER M1 ;
        RECT 0.479 12.516 0.481 14.952 ;
  LAYER M1 ;
        RECT 0.559 12.516 0.561 14.952 ;
  LAYER M1 ;
        RECT 0.639 12.516 0.641 14.952 ;
  LAYER M1 ;
        RECT 0.719 12.516 0.721 14.952 ;
  LAYER M1 ;
        RECT 0.799 12.516 0.801 14.952 ;
  LAYER M1 ;
        RECT 0.879 12.516 0.881 14.952 ;
  LAYER M1 ;
        RECT 0.959 12.516 0.961 14.952 ;
  LAYER M1 ;
        RECT 1.039 12.516 1.041 14.952 ;
  LAYER M1 ;
        RECT 1.119 12.516 1.121 14.952 ;
  LAYER M1 ;
        RECT 1.199 12.516 1.201 14.952 ;
  LAYER M1 ;
        RECT 1.279 12.516 1.281 14.952 ;
  LAYER M1 ;
        RECT 1.359 12.516 1.361 14.952 ;
  LAYER M1 ;
        RECT 1.439 12.516 1.441 14.952 ;
  LAYER M1 ;
        RECT 1.519 12.516 1.521 14.952 ;
  LAYER M1 ;
        RECT 1.599 12.516 1.601 14.952 ;
  LAYER M1 ;
        RECT 1.679 12.516 1.681 14.952 ;
  LAYER M1 ;
        RECT 1.759 12.516 1.761 14.952 ;
  LAYER M1 ;
        RECT 1.839 12.516 1.841 14.952 ;
  LAYER M1 ;
        RECT 1.919 12.516 1.921 14.952 ;
  LAYER M1 ;
        RECT 1.999 12.516 2.001 14.952 ;
  LAYER M1 ;
        RECT 2.079 12.516 2.081 14.952 ;
  LAYER M1 ;
        RECT 2.159 12.516 2.161 14.952 ;
  LAYER M1 ;
        RECT 2.239 12.516 2.241 14.952 ;
  LAYER M1 ;
        RECT 2.319 12.516 2.321 14.952 ;
  LAYER M1 ;
        RECT 2.399 12.516 2.401 14.952 ;
  LAYER M1 ;
        RECT 2.479 12.516 2.481 14.952 ;
  LAYER M1 ;
        RECT 2.559 12.516 2.561 14.952 ;
  LAYER M1 ;
        RECT 2.639 12.516 2.641 14.952 ;
  LAYER M1 ;
        RECT 2.719 12.516 2.721 14.952 ;
  LAYER M2 ;
        RECT 0.4 12.515 2.8 12.517 ;
  LAYER M2 ;
        RECT 0.4 12.599 2.8 12.601 ;
  LAYER M2 ;
        RECT 0.4 12.683 2.8 12.685 ;
  LAYER M2 ;
        RECT 0.4 12.767 2.8 12.769 ;
  LAYER M2 ;
        RECT 0.4 12.851 2.8 12.853 ;
  LAYER M2 ;
        RECT 0.4 12.935 2.8 12.937 ;
  LAYER M2 ;
        RECT 0.4 13.019 2.8 13.021 ;
  LAYER M2 ;
        RECT 0.4 13.103 2.8 13.105 ;
  LAYER M2 ;
        RECT 0.4 13.187 2.8 13.189 ;
  LAYER M2 ;
        RECT 0.4 13.271 2.8 13.273 ;
  LAYER M2 ;
        RECT 0.4 13.355 2.8 13.357 ;
  LAYER M2 ;
        RECT 0.4 13.439 2.8 13.441 ;
  LAYER M2 ;
        RECT 0.4 13.5225 2.8 13.5245 ;
  LAYER M2 ;
        RECT 0.4 13.607 2.8 13.609 ;
  LAYER M2 ;
        RECT 0.4 13.691 2.8 13.693 ;
  LAYER M2 ;
        RECT 0.4 13.775 2.8 13.777 ;
  LAYER M2 ;
        RECT 0.4 13.859 2.8 13.861 ;
  LAYER M2 ;
        RECT 0.4 13.943 2.8 13.945 ;
  LAYER M2 ;
        RECT 0.4 14.027 2.8 14.029 ;
  LAYER M2 ;
        RECT 0.4 14.111 2.8 14.113 ;
  LAYER M2 ;
        RECT 0.4 14.195 2.8 14.197 ;
  LAYER M2 ;
        RECT 0.4 14.279 2.8 14.281 ;
  LAYER M2 ;
        RECT 0.4 14.363 2.8 14.365 ;
  LAYER M2 ;
        RECT 0.4 14.447 2.8 14.449 ;
  LAYER M2 ;
        RECT 0.4 14.531 2.8 14.533 ;
  LAYER M2 ;
        RECT 0.4 14.615 2.8 14.617 ;
  LAYER M2 ;
        RECT 0.4 14.699 2.8 14.701 ;
  LAYER M2 ;
        RECT 0.4 14.783 2.8 14.785 ;
  LAYER M2 ;
        RECT 0.4 14.867 2.8 14.869 ;
  LAYER M1 ;
        RECT 0.384 15.42 0.416 17.928 ;
  LAYER M1 ;
        RECT 0.448 15.42 0.48 17.928 ;
  LAYER M1 ;
        RECT 0.512 15.42 0.544 17.928 ;
  LAYER M1 ;
        RECT 0.576 15.42 0.608 17.928 ;
  LAYER M1 ;
        RECT 0.64 15.42 0.672 17.928 ;
  LAYER M1 ;
        RECT 0.704 15.42 0.736 17.928 ;
  LAYER M1 ;
        RECT 0.768 15.42 0.8 17.928 ;
  LAYER M1 ;
        RECT 0.832 15.42 0.864 17.928 ;
  LAYER M1 ;
        RECT 0.896 15.42 0.928 17.928 ;
  LAYER M1 ;
        RECT 0.96 15.42 0.992 17.928 ;
  LAYER M1 ;
        RECT 1.024 15.42 1.056 17.928 ;
  LAYER M1 ;
        RECT 1.088 15.42 1.12 17.928 ;
  LAYER M1 ;
        RECT 1.152 15.42 1.184 17.928 ;
  LAYER M1 ;
        RECT 1.216 15.42 1.248 17.928 ;
  LAYER M1 ;
        RECT 1.28 15.42 1.312 17.928 ;
  LAYER M1 ;
        RECT 1.344 15.42 1.376 17.928 ;
  LAYER M1 ;
        RECT 1.408 15.42 1.44 17.928 ;
  LAYER M1 ;
        RECT 1.472 15.42 1.504 17.928 ;
  LAYER M1 ;
        RECT 1.536 15.42 1.568 17.928 ;
  LAYER M1 ;
        RECT 1.6 15.42 1.632 17.928 ;
  LAYER M1 ;
        RECT 1.664 15.42 1.696 17.928 ;
  LAYER M1 ;
        RECT 1.728 15.42 1.76 17.928 ;
  LAYER M1 ;
        RECT 1.792 15.42 1.824 17.928 ;
  LAYER M1 ;
        RECT 1.856 15.42 1.888 17.928 ;
  LAYER M1 ;
        RECT 1.92 15.42 1.952 17.928 ;
  LAYER M1 ;
        RECT 1.984 15.42 2.016 17.928 ;
  LAYER M1 ;
        RECT 2.048 15.42 2.08 17.928 ;
  LAYER M1 ;
        RECT 2.112 15.42 2.144 17.928 ;
  LAYER M1 ;
        RECT 2.176 15.42 2.208 17.928 ;
  LAYER M1 ;
        RECT 2.24 15.42 2.272 17.928 ;
  LAYER M1 ;
        RECT 2.304 15.42 2.336 17.928 ;
  LAYER M1 ;
        RECT 2.368 15.42 2.4 17.928 ;
  LAYER M1 ;
        RECT 2.432 15.42 2.464 17.928 ;
  LAYER M1 ;
        RECT 2.496 15.42 2.528 17.928 ;
  LAYER M1 ;
        RECT 2.56 15.42 2.592 17.928 ;
  LAYER M1 ;
        RECT 2.624 15.42 2.656 17.928 ;
  LAYER M1 ;
        RECT 2.688 15.42 2.72 17.928 ;
  LAYER M2 ;
        RECT 0.364 15.504 2.836 15.536 ;
  LAYER M2 ;
        RECT 0.364 15.568 2.836 15.6 ;
  LAYER M2 ;
        RECT 0.364 15.632 2.836 15.664 ;
  LAYER M2 ;
        RECT 0.364 15.696 2.836 15.728 ;
  LAYER M2 ;
        RECT 0.364 15.76 2.836 15.792 ;
  LAYER M2 ;
        RECT 0.364 15.824 2.836 15.856 ;
  LAYER M2 ;
        RECT 0.364 15.888 2.836 15.92 ;
  LAYER M2 ;
        RECT 0.364 15.952 2.836 15.984 ;
  LAYER M2 ;
        RECT 0.364 16.016 2.836 16.048 ;
  LAYER M2 ;
        RECT 0.364 16.08 2.836 16.112 ;
  LAYER M2 ;
        RECT 0.364 16.144 2.836 16.176 ;
  LAYER M2 ;
        RECT 0.364 16.208 2.836 16.24 ;
  LAYER M2 ;
        RECT 0.364 16.272 2.836 16.304 ;
  LAYER M2 ;
        RECT 0.364 16.336 2.836 16.368 ;
  LAYER M2 ;
        RECT 0.364 16.4 2.836 16.432 ;
  LAYER M2 ;
        RECT 0.364 16.464 2.836 16.496 ;
  LAYER M2 ;
        RECT 0.364 16.528 2.836 16.56 ;
  LAYER M2 ;
        RECT 0.364 16.592 2.836 16.624 ;
  LAYER M2 ;
        RECT 0.364 16.656 2.836 16.688 ;
  LAYER M2 ;
        RECT 0.364 16.72 2.836 16.752 ;
  LAYER M2 ;
        RECT 0.364 16.784 2.836 16.816 ;
  LAYER M2 ;
        RECT 0.364 16.848 2.836 16.88 ;
  LAYER M2 ;
        RECT 0.364 16.912 2.836 16.944 ;
  LAYER M2 ;
        RECT 0.364 16.976 2.836 17.008 ;
  LAYER M2 ;
        RECT 0.364 17.04 2.836 17.072 ;
  LAYER M2 ;
        RECT 0.364 17.104 2.836 17.136 ;
  LAYER M2 ;
        RECT 0.364 17.168 2.836 17.2 ;
  LAYER M2 ;
        RECT 0.364 17.232 2.836 17.264 ;
  LAYER M2 ;
        RECT 0.364 17.296 2.836 17.328 ;
  LAYER M2 ;
        RECT 0.364 17.36 2.836 17.392 ;
  LAYER M2 ;
        RECT 0.364 17.424 2.836 17.456 ;
  LAYER M2 ;
        RECT 0.364 17.488 2.836 17.52 ;
  LAYER M2 ;
        RECT 0.364 17.552 2.836 17.584 ;
  LAYER M2 ;
        RECT 0.364 17.616 2.836 17.648 ;
  LAYER M2 ;
        RECT 0.364 17.68 2.836 17.712 ;
  LAYER M2 ;
        RECT 0.364 17.744 2.836 17.776 ;
  LAYER M3 ;
        RECT 0.384 15.42 0.416 17.928 ;
  LAYER M3 ;
        RECT 0.448 15.42 0.48 17.928 ;
  LAYER M3 ;
        RECT 0.512 15.42 0.544 17.928 ;
  LAYER M3 ;
        RECT 0.576 15.42 0.608 17.928 ;
  LAYER M3 ;
        RECT 0.64 15.42 0.672 17.928 ;
  LAYER M3 ;
        RECT 0.704 15.42 0.736 17.928 ;
  LAYER M3 ;
        RECT 0.768 15.42 0.8 17.928 ;
  LAYER M3 ;
        RECT 0.832 15.42 0.864 17.928 ;
  LAYER M3 ;
        RECT 0.896 15.42 0.928 17.928 ;
  LAYER M3 ;
        RECT 0.96 15.42 0.992 17.928 ;
  LAYER M3 ;
        RECT 1.024 15.42 1.056 17.928 ;
  LAYER M3 ;
        RECT 1.088 15.42 1.12 17.928 ;
  LAYER M3 ;
        RECT 1.152 15.42 1.184 17.928 ;
  LAYER M3 ;
        RECT 1.216 15.42 1.248 17.928 ;
  LAYER M3 ;
        RECT 1.28 15.42 1.312 17.928 ;
  LAYER M3 ;
        RECT 1.344 15.42 1.376 17.928 ;
  LAYER M3 ;
        RECT 1.408 15.42 1.44 17.928 ;
  LAYER M3 ;
        RECT 1.472 15.42 1.504 17.928 ;
  LAYER M3 ;
        RECT 1.536 15.42 1.568 17.928 ;
  LAYER M3 ;
        RECT 1.6 15.42 1.632 17.928 ;
  LAYER M3 ;
        RECT 1.664 15.42 1.696 17.928 ;
  LAYER M3 ;
        RECT 1.728 15.42 1.76 17.928 ;
  LAYER M3 ;
        RECT 1.792 15.42 1.824 17.928 ;
  LAYER M3 ;
        RECT 1.856 15.42 1.888 17.928 ;
  LAYER M3 ;
        RECT 1.92 15.42 1.952 17.928 ;
  LAYER M3 ;
        RECT 1.984 15.42 2.016 17.928 ;
  LAYER M3 ;
        RECT 2.048 15.42 2.08 17.928 ;
  LAYER M3 ;
        RECT 2.112 15.42 2.144 17.928 ;
  LAYER M3 ;
        RECT 2.176 15.42 2.208 17.928 ;
  LAYER M3 ;
        RECT 2.24 15.42 2.272 17.928 ;
  LAYER M3 ;
        RECT 2.304 15.42 2.336 17.928 ;
  LAYER M3 ;
        RECT 2.368 15.42 2.4 17.928 ;
  LAYER M3 ;
        RECT 2.432 15.42 2.464 17.928 ;
  LAYER M3 ;
        RECT 2.496 15.42 2.528 17.928 ;
  LAYER M3 ;
        RECT 2.56 15.42 2.592 17.928 ;
  LAYER M3 ;
        RECT 2.624 15.42 2.656 17.928 ;
  LAYER M3 ;
        RECT 2.688 15.42 2.72 17.928 ;
  LAYER M3 ;
        RECT 2.784 15.42 2.816 17.928 ;
  LAYER M1 ;
        RECT 0.399 15.456 0.401 17.892 ;
  LAYER M1 ;
        RECT 0.479 15.456 0.481 17.892 ;
  LAYER M1 ;
        RECT 0.559 15.456 0.561 17.892 ;
  LAYER M1 ;
        RECT 0.639 15.456 0.641 17.892 ;
  LAYER M1 ;
        RECT 0.719 15.456 0.721 17.892 ;
  LAYER M1 ;
        RECT 0.799 15.456 0.801 17.892 ;
  LAYER M1 ;
        RECT 0.879 15.456 0.881 17.892 ;
  LAYER M1 ;
        RECT 0.959 15.456 0.961 17.892 ;
  LAYER M1 ;
        RECT 1.039 15.456 1.041 17.892 ;
  LAYER M1 ;
        RECT 1.119 15.456 1.121 17.892 ;
  LAYER M1 ;
        RECT 1.199 15.456 1.201 17.892 ;
  LAYER M1 ;
        RECT 1.279 15.456 1.281 17.892 ;
  LAYER M1 ;
        RECT 1.359 15.456 1.361 17.892 ;
  LAYER M1 ;
        RECT 1.439 15.456 1.441 17.892 ;
  LAYER M1 ;
        RECT 1.519 15.456 1.521 17.892 ;
  LAYER M1 ;
        RECT 1.599 15.456 1.601 17.892 ;
  LAYER M1 ;
        RECT 1.679 15.456 1.681 17.892 ;
  LAYER M1 ;
        RECT 1.759 15.456 1.761 17.892 ;
  LAYER M1 ;
        RECT 1.839 15.456 1.841 17.892 ;
  LAYER M1 ;
        RECT 1.919 15.456 1.921 17.892 ;
  LAYER M1 ;
        RECT 1.999 15.456 2.001 17.892 ;
  LAYER M1 ;
        RECT 2.079 15.456 2.081 17.892 ;
  LAYER M1 ;
        RECT 2.159 15.456 2.161 17.892 ;
  LAYER M1 ;
        RECT 2.239 15.456 2.241 17.892 ;
  LAYER M1 ;
        RECT 2.319 15.456 2.321 17.892 ;
  LAYER M1 ;
        RECT 2.399 15.456 2.401 17.892 ;
  LAYER M1 ;
        RECT 2.479 15.456 2.481 17.892 ;
  LAYER M1 ;
        RECT 2.559 15.456 2.561 17.892 ;
  LAYER M1 ;
        RECT 2.639 15.456 2.641 17.892 ;
  LAYER M1 ;
        RECT 2.719 15.456 2.721 17.892 ;
  LAYER M2 ;
        RECT 0.4 15.455 2.8 15.457 ;
  LAYER M2 ;
        RECT 0.4 15.539 2.8 15.541 ;
  LAYER M2 ;
        RECT 0.4 15.623 2.8 15.625 ;
  LAYER M2 ;
        RECT 0.4 15.707 2.8 15.709 ;
  LAYER M2 ;
        RECT 0.4 15.791 2.8 15.793 ;
  LAYER M2 ;
        RECT 0.4 15.875 2.8 15.877 ;
  LAYER M2 ;
        RECT 0.4 15.959 2.8 15.961 ;
  LAYER M2 ;
        RECT 0.4 16.043 2.8 16.045 ;
  LAYER M2 ;
        RECT 0.4 16.127 2.8 16.129 ;
  LAYER M2 ;
        RECT 0.4 16.211 2.8 16.213 ;
  LAYER M2 ;
        RECT 0.4 16.295 2.8 16.297 ;
  LAYER M2 ;
        RECT 0.4 16.379 2.8 16.381 ;
  LAYER M2 ;
        RECT 0.4 16.4625 2.8 16.4645 ;
  LAYER M2 ;
        RECT 0.4 16.547 2.8 16.549 ;
  LAYER M2 ;
        RECT 0.4 16.631 2.8 16.633 ;
  LAYER M2 ;
        RECT 0.4 16.715 2.8 16.717 ;
  LAYER M2 ;
        RECT 0.4 16.799 2.8 16.801 ;
  LAYER M2 ;
        RECT 0.4 16.883 2.8 16.885 ;
  LAYER M2 ;
        RECT 0.4 16.967 2.8 16.969 ;
  LAYER M2 ;
        RECT 0.4 17.051 2.8 17.053 ;
  LAYER M2 ;
        RECT 0.4 17.135 2.8 17.137 ;
  LAYER M2 ;
        RECT 0.4 17.219 2.8 17.221 ;
  LAYER M2 ;
        RECT 0.4 17.303 2.8 17.305 ;
  LAYER M2 ;
        RECT 0.4 17.387 2.8 17.389 ;
  LAYER M2 ;
        RECT 0.4 17.471 2.8 17.473 ;
  LAYER M2 ;
        RECT 0.4 17.555 2.8 17.557 ;
  LAYER M2 ;
        RECT 0.4 17.639 2.8 17.641 ;
  LAYER M2 ;
        RECT 0.4 17.723 2.8 17.725 ;
  LAYER M2 ;
        RECT 0.4 17.807 2.8 17.809 ;
  LAYER M1 ;
        RECT 0.384 18.36 0.416 20.868 ;
  LAYER M1 ;
        RECT 0.448 18.36 0.48 20.868 ;
  LAYER M1 ;
        RECT 0.512 18.36 0.544 20.868 ;
  LAYER M1 ;
        RECT 0.576 18.36 0.608 20.868 ;
  LAYER M1 ;
        RECT 0.64 18.36 0.672 20.868 ;
  LAYER M1 ;
        RECT 0.704 18.36 0.736 20.868 ;
  LAYER M1 ;
        RECT 0.768 18.36 0.8 20.868 ;
  LAYER M1 ;
        RECT 0.832 18.36 0.864 20.868 ;
  LAYER M1 ;
        RECT 0.896 18.36 0.928 20.868 ;
  LAYER M1 ;
        RECT 0.96 18.36 0.992 20.868 ;
  LAYER M1 ;
        RECT 1.024 18.36 1.056 20.868 ;
  LAYER M1 ;
        RECT 1.088 18.36 1.12 20.868 ;
  LAYER M1 ;
        RECT 1.152 18.36 1.184 20.868 ;
  LAYER M1 ;
        RECT 1.216 18.36 1.248 20.868 ;
  LAYER M1 ;
        RECT 1.28 18.36 1.312 20.868 ;
  LAYER M1 ;
        RECT 1.344 18.36 1.376 20.868 ;
  LAYER M1 ;
        RECT 1.408 18.36 1.44 20.868 ;
  LAYER M1 ;
        RECT 1.472 18.36 1.504 20.868 ;
  LAYER M1 ;
        RECT 1.536 18.36 1.568 20.868 ;
  LAYER M1 ;
        RECT 1.6 18.36 1.632 20.868 ;
  LAYER M1 ;
        RECT 1.664 18.36 1.696 20.868 ;
  LAYER M1 ;
        RECT 1.728 18.36 1.76 20.868 ;
  LAYER M1 ;
        RECT 1.792 18.36 1.824 20.868 ;
  LAYER M1 ;
        RECT 1.856 18.36 1.888 20.868 ;
  LAYER M1 ;
        RECT 1.92 18.36 1.952 20.868 ;
  LAYER M1 ;
        RECT 1.984 18.36 2.016 20.868 ;
  LAYER M1 ;
        RECT 2.048 18.36 2.08 20.868 ;
  LAYER M1 ;
        RECT 2.112 18.36 2.144 20.868 ;
  LAYER M1 ;
        RECT 2.176 18.36 2.208 20.868 ;
  LAYER M1 ;
        RECT 2.24 18.36 2.272 20.868 ;
  LAYER M1 ;
        RECT 2.304 18.36 2.336 20.868 ;
  LAYER M1 ;
        RECT 2.368 18.36 2.4 20.868 ;
  LAYER M1 ;
        RECT 2.432 18.36 2.464 20.868 ;
  LAYER M1 ;
        RECT 2.496 18.36 2.528 20.868 ;
  LAYER M1 ;
        RECT 2.56 18.36 2.592 20.868 ;
  LAYER M1 ;
        RECT 2.624 18.36 2.656 20.868 ;
  LAYER M1 ;
        RECT 2.688 18.36 2.72 20.868 ;
  LAYER M2 ;
        RECT 0.364 18.444 2.836 18.476 ;
  LAYER M2 ;
        RECT 0.364 18.508 2.836 18.54 ;
  LAYER M2 ;
        RECT 0.364 18.572 2.836 18.604 ;
  LAYER M2 ;
        RECT 0.364 18.636 2.836 18.668 ;
  LAYER M2 ;
        RECT 0.364 18.7 2.836 18.732 ;
  LAYER M2 ;
        RECT 0.364 18.764 2.836 18.796 ;
  LAYER M2 ;
        RECT 0.364 18.828 2.836 18.86 ;
  LAYER M2 ;
        RECT 0.364 18.892 2.836 18.924 ;
  LAYER M2 ;
        RECT 0.364 18.956 2.836 18.988 ;
  LAYER M2 ;
        RECT 0.364 19.02 2.836 19.052 ;
  LAYER M2 ;
        RECT 0.364 19.084 2.836 19.116 ;
  LAYER M2 ;
        RECT 0.364 19.148 2.836 19.18 ;
  LAYER M2 ;
        RECT 0.364 19.212 2.836 19.244 ;
  LAYER M2 ;
        RECT 0.364 19.276 2.836 19.308 ;
  LAYER M2 ;
        RECT 0.364 19.34 2.836 19.372 ;
  LAYER M2 ;
        RECT 0.364 19.404 2.836 19.436 ;
  LAYER M2 ;
        RECT 0.364 19.468 2.836 19.5 ;
  LAYER M2 ;
        RECT 0.364 19.532 2.836 19.564 ;
  LAYER M2 ;
        RECT 0.364 19.596 2.836 19.628 ;
  LAYER M2 ;
        RECT 0.364 19.66 2.836 19.692 ;
  LAYER M2 ;
        RECT 0.364 19.724 2.836 19.756 ;
  LAYER M2 ;
        RECT 0.364 19.788 2.836 19.82 ;
  LAYER M2 ;
        RECT 0.364 19.852 2.836 19.884 ;
  LAYER M2 ;
        RECT 0.364 19.916 2.836 19.948 ;
  LAYER M2 ;
        RECT 0.364 19.98 2.836 20.012 ;
  LAYER M2 ;
        RECT 0.364 20.044 2.836 20.076 ;
  LAYER M2 ;
        RECT 0.364 20.108 2.836 20.14 ;
  LAYER M2 ;
        RECT 0.364 20.172 2.836 20.204 ;
  LAYER M2 ;
        RECT 0.364 20.236 2.836 20.268 ;
  LAYER M2 ;
        RECT 0.364 20.3 2.836 20.332 ;
  LAYER M2 ;
        RECT 0.364 20.364 2.836 20.396 ;
  LAYER M2 ;
        RECT 0.364 20.428 2.836 20.46 ;
  LAYER M2 ;
        RECT 0.364 20.492 2.836 20.524 ;
  LAYER M2 ;
        RECT 0.364 20.556 2.836 20.588 ;
  LAYER M2 ;
        RECT 0.364 20.62 2.836 20.652 ;
  LAYER M2 ;
        RECT 0.364 20.684 2.836 20.716 ;
  LAYER M3 ;
        RECT 0.384 18.36 0.416 20.868 ;
  LAYER M3 ;
        RECT 0.448 18.36 0.48 20.868 ;
  LAYER M3 ;
        RECT 0.512 18.36 0.544 20.868 ;
  LAYER M3 ;
        RECT 0.576 18.36 0.608 20.868 ;
  LAYER M3 ;
        RECT 0.64 18.36 0.672 20.868 ;
  LAYER M3 ;
        RECT 0.704 18.36 0.736 20.868 ;
  LAYER M3 ;
        RECT 0.768 18.36 0.8 20.868 ;
  LAYER M3 ;
        RECT 0.832 18.36 0.864 20.868 ;
  LAYER M3 ;
        RECT 0.896 18.36 0.928 20.868 ;
  LAYER M3 ;
        RECT 0.96 18.36 0.992 20.868 ;
  LAYER M3 ;
        RECT 1.024 18.36 1.056 20.868 ;
  LAYER M3 ;
        RECT 1.088 18.36 1.12 20.868 ;
  LAYER M3 ;
        RECT 1.152 18.36 1.184 20.868 ;
  LAYER M3 ;
        RECT 1.216 18.36 1.248 20.868 ;
  LAYER M3 ;
        RECT 1.28 18.36 1.312 20.868 ;
  LAYER M3 ;
        RECT 1.344 18.36 1.376 20.868 ;
  LAYER M3 ;
        RECT 1.408 18.36 1.44 20.868 ;
  LAYER M3 ;
        RECT 1.472 18.36 1.504 20.868 ;
  LAYER M3 ;
        RECT 1.536 18.36 1.568 20.868 ;
  LAYER M3 ;
        RECT 1.6 18.36 1.632 20.868 ;
  LAYER M3 ;
        RECT 1.664 18.36 1.696 20.868 ;
  LAYER M3 ;
        RECT 1.728 18.36 1.76 20.868 ;
  LAYER M3 ;
        RECT 1.792 18.36 1.824 20.868 ;
  LAYER M3 ;
        RECT 1.856 18.36 1.888 20.868 ;
  LAYER M3 ;
        RECT 1.92 18.36 1.952 20.868 ;
  LAYER M3 ;
        RECT 1.984 18.36 2.016 20.868 ;
  LAYER M3 ;
        RECT 2.048 18.36 2.08 20.868 ;
  LAYER M3 ;
        RECT 2.112 18.36 2.144 20.868 ;
  LAYER M3 ;
        RECT 2.176 18.36 2.208 20.868 ;
  LAYER M3 ;
        RECT 2.24 18.36 2.272 20.868 ;
  LAYER M3 ;
        RECT 2.304 18.36 2.336 20.868 ;
  LAYER M3 ;
        RECT 2.368 18.36 2.4 20.868 ;
  LAYER M3 ;
        RECT 2.432 18.36 2.464 20.868 ;
  LAYER M3 ;
        RECT 2.496 18.36 2.528 20.868 ;
  LAYER M3 ;
        RECT 2.56 18.36 2.592 20.868 ;
  LAYER M3 ;
        RECT 2.624 18.36 2.656 20.868 ;
  LAYER M3 ;
        RECT 2.688 18.36 2.72 20.868 ;
  LAYER M3 ;
        RECT 2.784 18.36 2.816 20.868 ;
  LAYER M1 ;
        RECT 0.399 18.396 0.401 20.832 ;
  LAYER M1 ;
        RECT 0.479 18.396 0.481 20.832 ;
  LAYER M1 ;
        RECT 0.559 18.396 0.561 20.832 ;
  LAYER M1 ;
        RECT 0.639 18.396 0.641 20.832 ;
  LAYER M1 ;
        RECT 0.719 18.396 0.721 20.832 ;
  LAYER M1 ;
        RECT 0.799 18.396 0.801 20.832 ;
  LAYER M1 ;
        RECT 0.879 18.396 0.881 20.832 ;
  LAYER M1 ;
        RECT 0.959 18.396 0.961 20.832 ;
  LAYER M1 ;
        RECT 1.039 18.396 1.041 20.832 ;
  LAYER M1 ;
        RECT 1.119 18.396 1.121 20.832 ;
  LAYER M1 ;
        RECT 1.199 18.396 1.201 20.832 ;
  LAYER M1 ;
        RECT 1.279 18.396 1.281 20.832 ;
  LAYER M1 ;
        RECT 1.359 18.396 1.361 20.832 ;
  LAYER M1 ;
        RECT 1.439 18.396 1.441 20.832 ;
  LAYER M1 ;
        RECT 1.519 18.396 1.521 20.832 ;
  LAYER M1 ;
        RECT 1.599 18.396 1.601 20.832 ;
  LAYER M1 ;
        RECT 1.679 18.396 1.681 20.832 ;
  LAYER M1 ;
        RECT 1.759 18.396 1.761 20.832 ;
  LAYER M1 ;
        RECT 1.839 18.396 1.841 20.832 ;
  LAYER M1 ;
        RECT 1.919 18.396 1.921 20.832 ;
  LAYER M1 ;
        RECT 1.999 18.396 2.001 20.832 ;
  LAYER M1 ;
        RECT 2.079 18.396 2.081 20.832 ;
  LAYER M1 ;
        RECT 2.159 18.396 2.161 20.832 ;
  LAYER M1 ;
        RECT 2.239 18.396 2.241 20.832 ;
  LAYER M1 ;
        RECT 2.319 18.396 2.321 20.832 ;
  LAYER M1 ;
        RECT 2.399 18.396 2.401 20.832 ;
  LAYER M1 ;
        RECT 2.479 18.396 2.481 20.832 ;
  LAYER M1 ;
        RECT 2.559 18.396 2.561 20.832 ;
  LAYER M1 ;
        RECT 2.639 18.396 2.641 20.832 ;
  LAYER M1 ;
        RECT 2.719 18.396 2.721 20.832 ;
  LAYER M2 ;
        RECT 0.4 18.395 2.8 18.397 ;
  LAYER M2 ;
        RECT 0.4 18.479 2.8 18.481 ;
  LAYER M2 ;
        RECT 0.4 18.563 2.8 18.565 ;
  LAYER M2 ;
        RECT 0.4 18.647 2.8 18.649 ;
  LAYER M2 ;
        RECT 0.4 18.731 2.8 18.733 ;
  LAYER M2 ;
        RECT 0.4 18.815 2.8 18.817 ;
  LAYER M2 ;
        RECT 0.4 18.899 2.8 18.901 ;
  LAYER M2 ;
        RECT 0.4 18.983 2.8 18.985 ;
  LAYER M2 ;
        RECT 0.4 19.067 2.8 19.069 ;
  LAYER M2 ;
        RECT 0.4 19.151 2.8 19.153 ;
  LAYER M2 ;
        RECT 0.4 19.235 2.8 19.237 ;
  LAYER M2 ;
        RECT 0.4 19.319 2.8 19.321 ;
  LAYER M2 ;
        RECT 0.4 19.4025 2.8 19.4045 ;
  LAYER M2 ;
        RECT 0.4 19.487 2.8 19.489 ;
  LAYER M2 ;
        RECT 0.4 19.571 2.8 19.573 ;
  LAYER M2 ;
        RECT 0.4 19.655 2.8 19.657 ;
  LAYER M2 ;
        RECT 0.4 19.739 2.8 19.741 ;
  LAYER M2 ;
        RECT 0.4 19.823 2.8 19.825 ;
  LAYER M2 ;
        RECT 0.4 19.907 2.8 19.909 ;
  LAYER M2 ;
        RECT 0.4 19.991 2.8 19.993 ;
  LAYER M2 ;
        RECT 0.4 20.075 2.8 20.077 ;
  LAYER M2 ;
        RECT 0.4 20.159 2.8 20.161 ;
  LAYER M2 ;
        RECT 0.4 20.243 2.8 20.245 ;
  LAYER M2 ;
        RECT 0.4 20.327 2.8 20.329 ;
  LAYER M2 ;
        RECT 0.4 20.411 2.8 20.413 ;
  LAYER M2 ;
        RECT 0.4 20.495 2.8 20.497 ;
  LAYER M2 ;
        RECT 0.4 20.579 2.8 20.581 ;
  LAYER M2 ;
        RECT 0.4 20.663 2.8 20.665 ;
  LAYER M2 ;
        RECT 0.4 20.747 2.8 20.749 ;
  LAYER M1 ;
        RECT 0.384 21.3 0.416 23.808 ;
  LAYER M1 ;
        RECT 0.448 21.3 0.48 23.808 ;
  LAYER M1 ;
        RECT 0.512 21.3 0.544 23.808 ;
  LAYER M1 ;
        RECT 0.576 21.3 0.608 23.808 ;
  LAYER M1 ;
        RECT 0.64 21.3 0.672 23.808 ;
  LAYER M1 ;
        RECT 0.704 21.3 0.736 23.808 ;
  LAYER M1 ;
        RECT 0.768 21.3 0.8 23.808 ;
  LAYER M1 ;
        RECT 0.832 21.3 0.864 23.808 ;
  LAYER M1 ;
        RECT 0.896 21.3 0.928 23.808 ;
  LAYER M1 ;
        RECT 0.96 21.3 0.992 23.808 ;
  LAYER M1 ;
        RECT 1.024 21.3 1.056 23.808 ;
  LAYER M1 ;
        RECT 1.088 21.3 1.12 23.808 ;
  LAYER M1 ;
        RECT 1.152 21.3 1.184 23.808 ;
  LAYER M1 ;
        RECT 1.216 21.3 1.248 23.808 ;
  LAYER M1 ;
        RECT 1.28 21.3 1.312 23.808 ;
  LAYER M1 ;
        RECT 1.344 21.3 1.376 23.808 ;
  LAYER M1 ;
        RECT 1.408 21.3 1.44 23.808 ;
  LAYER M1 ;
        RECT 1.472 21.3 1.504 23.808 ;
  LAYER M1 ;
        RECT 1.536 21.3 1.568 23.808 ;
  LAYER M1 ;
        RECT 1.6 21.3 1.632 23.808 ;
  LAYER M1 ;
        RECT 1.664 21.3 1.696 23.808 ;
  LAYER M1 ;
        RECT 1.728 21.3 1.76 23.808 ;
  LAYER M1 ;
        RECT 1.792 21.3 1.824 23.808 ;
  LAYER M1 ;
        RECT 1.856 21.3 1.888 23.808 ;
  LAYER M1 ;
        RECT 1.92 21.3 1.952 23.808 ;
  LAYER M1 ;
        RECT 1.984 21.3 2.016 23.808 ;
  LAYER M1 ;
        RECT 2.048 21.3 2.08 23.808 ;
  LAYER M1 ;
        RECT 2.112 21.3 2.144 23.808 ;
  LAYER M1 ;
        RECT 2.176 21.3 2.208 23.808 ;
  LAYER M1 ;
        RECT 2.24 21.3 2.272 23.808 ;
  LAYER M1 ;
        RECT 2.304 21.3 2.336 23.808 ;
  LAYER M1 ;
        RECT 2.368 21.3 2.4 23.808 ;
  LAYER M1 ;
        RECT 2.432 21.3 2.464 23.808 ;
  LAYER M1 ;
        RECT 2.496 21.3 2.528 23.808 ;
  LAYER M1 ;
        RECT 2.56 21.3 2.592 23.808 ;
  LAYER M1 ;
        RECT 2.624 21.3 2.656 23.808 ;
  LAYER M1 ;
        RECT 2.688 21.3 2.72 23.808 ;
  LAYER M2 ;
        RECT 0.364 21.384 2.836 21.416 ;
  LAYER M2 ;
        RECT 0.364 21.448 2.836 21.48 ;
  LAYER M2 ;
        RECT 0.364 21.512 2.836 21.544 ;
  LAYER M2 ;
        RECT 0.364 21.576 2.836 21.608 ;
  LAYER M2 ;
        RECT 0.364 21.64 2.836 21.672 ;
  LAYER M2 ;
        RECT 0.364 21.704 2.836 21.736 ;
  LAYER M2 ;
        RECT 0.364 21.768 2.836 21.8 ;
  LAYER M2 ;
        RECT 0.364 21.832 2.836 21.864 ;
  LAYER M2 ;
        RECT 0.364 21.896 2.836 21.928 ;
  LAYER M2 ;
        RECT 0.364 21.96 2.836 21.992 ;
  LAYER M2 ;
        RECT 0.364 22.024 2.836 22.056 ;
  LAYER M2 ;
        RECT 0.364 22.088 2.836 22.12 ;
  LAYER M2 ;
        RECT 0.364 22.152 2.836 22.184 ;
  LAYER M2 ;
        RECT 0.364 22.216 2.836 22.248 ;
  LAYER M2 ;
        RECT 0.364 22.28 2.836 22.312 ;
  LAYER M2 ;
        RECT 0.364 22.344 2.836 22.376 ;
  LAYER M2 ;
        RECT 0.364 22.408 2.836 22.44 ;
  LAYER M2 ;
        RECT 0.364 22.472 2.836 22.504 ;
  LAYER M2 ;
        RECT 0.364 22.536 2.836 22.568 ;
  LAYER M2 ;
        RECT 0.364 22.6 2.836 22.632 ;
  LAYER M2 ;
        RECT 0.364 22.664 2.836 22.696 ;
  LAYER M2 ;
        RECT 0.364 22.728 2.836 22.76 ;
  LAYER M2 ;
        RECT 0.364 22.792 2.836 22.824 ;
  LAYER M2 ;
        RECT 0.364 22.856 2.836 22.888 ;
  LAYER M2 ;
        RECT 0.364 22.92 2.836 22.952 ;
  LAYER M2 ;
        RECT 0.364 22.984 2.836 23.016 ;
  LAYER M2 ;
        RECT 0.364 23.048 2.836 23.08 ;
  LAYER M2 ;
        RECT 0.364 23.112 2.836 23.144 ;
  LAYER M2 ;
        RECT 0.364 23.176 2.836 23.208 ;
  LAYER M2 ;
        RECT 0.364 23.24 2.836 23.272 ;
  LAYER M2 ;
        RECT 0.364 23.304 2.836 23.336 ;
  LAYER M2 ;
        RECT 0.364 23.368 2.836 23.4 ;
  LAYER M2 ;
        RECT 0.364 23.432 2.836 23.464 ;
  LAYER M2 ;
        RECT 0.364 23.496 2.836 23.528 ;
  LAYER M2 ;
        RECT 0.364 23.56 2.836 23.592 ;
  LAYER M2 ;
        RECT 0.364 23.624 2.836 23.656 ;
  LAYER M3 ;
        RECT 0.384 21.3 0.416 23.808 ;
  LAYER M3 ;
        RECT 0.448 21.3 0.48 23.808 ;
  LAYER M3 ;
        RECT 0.512 21.3 0.544 23.808 ;
  LAYER M3 ;
        RECT 0.576 21.3 0.608 23.808 ;
  LAYER M3 ;
        RECT 0.64 21.3 0.672 23.808 ;
  LAYER M3 ;
        RECT 0.704 21.3 0.736 23.808 ;
  LAYER M3 ;
        RECT 0.768 21.3 0.8 23.808 ;
  LAYER M3 ;
        RECT 0.832 21.3 0.864 23.808 ;
  LAYER M3 ;
        RECT 0.896 21.3 0.928 23.808 ;
  LAYER M3 ;
        RECT 0.96 21.3 0.992 23.808 ;
  LAYER M3 ;
        RECT 1.024 21.3 1.056 23.808 ;
  LAYER M3 ;
        RECT 1.088 21.3 1.12 23.808 ;
  LAYER M3 ;
        RECT 1.152 21.3 1.184 23.808 ;
  LAYER M3 ;
        RECT 1.216 21.3 1.248 23.808 ;
  LAYER M3 ;
        RECT 1.28 21.3 1.312 23.808 ;
  LAYER M3 ;
        RECT 1.344 21.3 1.376 23.808 ;
  LAYER M3 ;
        RECT 1.408 21.3 1.44 23.808 ;
  LAYER M3 ;
        RECT 1.472 21.3 1.504 23.808 ;
  LAYER M3 ;
        RECT 1.536 21.3 1.568 23.808 ;
  LAYER M3 ;
        RECT 1.6 21.3 1.632 23.808 ;
  LAYER M3 ;
        RECT 1.664 21.3 1.696 23.808 ;
  LAYER M3 ;
        RECT 1.728 21.3 1.76 23.808 ;
  LAYER M3 ;
        RECT 1.792 21.3 1.824 23.808 ;
  LAYER M3 ;
        RECT 1.856 21.3 1.888 23.808 ;
  LAYER M3 ;
        RECT 1.92 21.3 1.952 23.808 ;
  LAYER M3 ;
        RECT 1.984 21.3 2.016 23.808 ;
  LAYER M3 ;
        RECT 2.048 21.3 2.08 23.808 ;
  LAYER M3 ;
        RECT 2.112 21.3 2.144 23.808 ;
  LAYER M3 ;
        RECT 2.176 21.3 2.208 23.808 ;
  LAYER M3 ;
        RECT 2.24 21.3 2.272 23.808 ;
  LAYER M3 ;
        RECT 2.304 21.3 2.336 23.808 ;
  LAYER M3 ;
        RECT 2.368 21.3 2.4 23.808 ;
  LAYER M3 ;
        RECT 2.432 21.3 2.464 23.808 ;
  LAYER M3 ;
        RECT 2.496 21.3 2.528 23.808 ;
  LAYER M3 ;
        RECT 2.56 21.3 2.592 23.808 ;
  LAYER M3 ;
        RECT 2.624 21.3 2.656 23.808 ;
  LAYER M3 ;
        RECT 2.688 21.3 2.72 23.808 ;
  LAYER M3 ;
        RECT 2.784 21.3 2.816 23.808 ;
  LAYER M1 ;
        RECT 0.399 21.336 0.401 23.772 ;
  LAYER M1 ;
        RECT 0.479 21.336 0.481 23.772 ;
  LAYER M1 ;
        RECT 0.559 21.336 0.561 23.772 ;
  LAYER M1 ;
        RECT 0.639 21.336 0.641 23.772 ;
  LAYER M1 ;
        RECT 0.719 21.336 0.721 23.772 ;
  LAYER M1 ;
        RECT 0.799 21.336 0.801 23.772 ;
  LAYER M1 ;
        RECT 0.879 21.336 0.881 23.772 ;
  LAYER M1 ;
        RECT 0.959 21.336 0.961 23.772 ;
  LAYER M1 ;
        RECT 1.039 21.336 1.041 23.772 ;
  LAYER M1 ;
        RECT 1.119 21.336 1.121 23.772 ;
  LAYER M1 ;
        RECT 1.199 21.336 1.201 23.772 ;
  LAYER M1 ;
        RECT 1.279 21.336 1.281 23.772 ;
  LAYER M1 ;
        RECT 1.359 21.336 1.361 23.772 ;
  LAYER M1 ;
        RECT 1.439 21.336 1.441 23.772 ;
  LAYER M1 ;
        RECT 1.519 21.336 1.521 23.772 ;
  LAYER M1 ;
        RECT 1.599 21.336 1.601 23.772 ;
  LAYER M1 ;
        RECT 1.679 21.336 1.681 23.772 ;
  LAYER M1 ;
        RECT 1.759 21.336 1.761 23.772 ;
  LAYER M1 ;
        RECT 1.839 21.336 1.841 23.772 ;
  LAYER M1 ;
        RECT 1.919 21.336 1.921 23.772 ;
  LAYER M1 ;
        RECT 1.999 21.336 2.001 23.772 ;
  LAYER M1 ;
        RECT 2.079 21.336 2.081 23.772 ;
  LAYER M1 ;
        RECT 2.159 21.336 2.161 23.772 ;
  LAYER M1 ;
        RECT 2.239 21.336 2.241 23.772 ;
  LAYER M1 ;
        RECT 2.319 21.336 2.321 23.772 ;
  LAYER M1 ;
        RECT 2.399 21.336 2.401 23.772 ;
  LAYER M1 ;
        RECT 2.479 21.336 2.481 23.772 ;
  LAYER M1 ;
        RECT 2.559 21.336 2.561 23.772 ;
  LAYER M1 ;
        RECT 2.639 21.336 2.641 23.772 ;
  LAYER M1 ;
        RECT 2.719 21.336 2.721 23.772 ;
  LAYER M2 ;
        RECT 0.4 21.335 2.8 21.337 ;
  LAYER M2 ;
        RECT 0.4 21.419 2.8 21.421 ;
  LAYER M2 ;
        RECT 0.4 21.503 2.8 21.505 ;
  LAYER M2 ;
        RECT 0.4 21.587 2.8 21.589 ;
  LAYER M2 ;
        RECT 0.4 21.671 2.8 21.673 ;
  LAYER M2 ;
        RECT 0.4 21.755 2.8 21.757 ;
  LAYER M2 ;
        RECT 0.4 21.839 2.8 21.841 ;
  LAYER M2 ;
        RECT 0.4 21.923 2.8 21.925 ;
  LAYER M2 ;
        RECT 0.4 22.007 2.8 22.009 ;
  LAYER M2 ;
        RECT 0.4 22.091 2.8 22.093 ;
  LAYER M2 ;
        RECT 0.4 22.175 2.8 22.177 ;
  LAYER M2 ;
        RECT 0.4 22.259 2.8 22.261 ;
  LAYER M2 ;
        RECT 0.4 22.3425 2.8 22.3445 ;
  LAYER M2 ;
        RECT 0.4 22.427 2.8 22.429 ;
  LAYER M2 ;
        RECT 0.4 22.511 2.8 22.513 ;
  LAYER M2 ;
        RECT 0.4 22.595 2.8 22.597 ;
  LAYER M2 ;
        RECT 0.4 22.679 2.8 22.681 ;
  LAYER M2 ;
        RECT 0.4 22.763 2.8 22.765 ;
  LAYER M2 ;
        RECT 0.4 22.847 2.8 22.849 ;
  LAYER M2 ;
        RECT 0.4 22.931 2.8 22.933 ;
  LAYER M2 ;
        RECT 0.4 23.015 2.8 23.017 ;
  LAYER M2 ;
        RECT 0.4 23.099 2.8 23.101 ;
  LAYER M2 ;
        RECT 0.4 23.183 2.8 23.185 ;
  LAYER M2 ;
        RECT 0.4 23.267 2.8 23.269 ;
  LAYER M2 ;
        RECT 0.4 23.351 2.8 23.353 ;
  LAYER M2 ;
        RECT 0.4 23.435 2.8 23.437 ;
  LAYER M2 ;
        RECT 0.4 23.519 2.8 23.521 ;
  LAYER M2 ;
        RECT 0.4 23.603 2.8 23.605 ;
  LAYER M2 ;
        RECT 0.4 23.687 2.8 23.689 ;
  LAYER M1 ;
        RECT 3.264 0.72 3.296 3.228 ;
  LAYER M1 ;
        RECT 3.328 0.72 3.36 3.228 ;
  LAYER M1 ;
        RECT 3.392 0.72 3.424 3.228 ;
  LAYER M1 ;
        RECT 3.456 0.72 3.488 3.228 ;
  LAYER M1 ;
        RECT 3.52 0.72 3.552 3.228 ;
  LAYER M1 ;
        RECT 3.584 0.72 3.616 3.228 ;
  LAYER M1 ;
        RECT 3.648 0.72 3.68 3.228 ;
  LAYER M1 ;
        RECT 3.712 0.72 3.744 3.228 ;
  LAYER M1 ;
        RECT 3.776 0.72 3.808 3.228 ;
  LAYER M1 ;
        RECT 3.84 0.72 3.872 3.228 ;
  LAYER M1 ;
        RECT 3.904 0.72 3.936 3.228 ;
  LAYER M1 ;
        RECT 3.968 0.72 4 3.228 ;
  LAYER M1 ;
        RECT 4.032 0.72 4.064 3.228 ;
  LAYER M1 ;
        RECT 4.096 0.72 4.128 3.228 ;
  LAYER M1 ;
        RECT 4.16 0.72 4.192 3.228 ;
  LAYER M1 ;
        RECT 4.224 0.72 4.256 3.228 ;
  LAYER M1 ;
        RECT 4.288 0.72 4.32 3.228 ;
  LAYER M1 ;
        RECT 4.352 0.72 4.384 3.228 ;
  LAYER M1 ;
        RECT 4.416 0.72 4.448 3.228 ;
  LAYER M1 ;
        RECT 4.48 0.72 4.512 3.228 ;
  LAYER M1 ;
        RECT 4.544 0.72 4.576 3.228 ;
  LAYER M1 ;
        RECT 4.608 0.72 4.64 3.228 ;
  LAYER M1 ;
        RECT 4.672 0.72 4.704 3.228 ;
  LAYER M1 ;
        RECT 4.736 0.72 4.768 3.228 ;
  LAYER M1 ;
        RECT 4.8 0.72 4.832 3.228 ;
  LAYER M1 ;
        RECT 4.864 0.72 4.896 3.228 ;
  LAYER M1 ;
        RECT 4.928 0.72 4.96 3.228 ;
  LAYER M1 ;
        RECT 4.992 0.72 5.024 3.228 ;
  LAYER M1 ;
        RECT 5.056 0.72 5.088 3.228 ;
  LAYER M1 ;
        RECT 5.12 0.72 5.152 3.228 ;
  LAYER M1 ;
        RECT 5.184 0.72 5.216 3.228 ;
  LAYER M1 ;
        RECT 5.248 0.72 5.28 3.228 ;
  LAYER M1 ;
        RECT 5.312 0.72 5.344 3.228 ;
  LAYER M1 ;
        RECT 5.376 0.72 5.408 3.228 ;
  LAYER M1 ;
        RECT 5.44 0.72 5.472 3.228 ;
  LAYER M1 ;
        RECT 5.504 0.72 5.536 3.228 ;
  LAYER M1 ;
        RECT 5.568 0.72 5.6 3.228 ;
  LAYER M2 ;
        RECT 3.244 0.804 5.716 0.836 ;
  LAYER M2 ;
        RECT 3.244 0.868 5.716 0.9 ;
  LAYER M2 ;
        RECT 3.244 0.932 5.716 0.964 ;
  LAYER M2 ;
        RECT 3.244 0.996 5.716 1.028 ;
  LAYER M2 ;
        RECT 3.244 1.06 5.716 1.092 ;
  LAYER M2 ;
        RECT 3.244 1.124 5.716 1.156 ;
  LAYER M2 ;
        RECT 3.244 1.188 5.716 1.22 ;
  LAYER M2 ;
        RECT 3.244 1.252 5.716 1.284 ;
  LAYER M2 ;
        RECT 3.244 1.316 5.716 1.348 ;
  LAYER M2 ;
        RECT 3.244 1.38 5.716 1.412 ;
  LAYER M2 ;
        RECT 3.244 1.444 5.716 1.476 ;
  LAYER M2 ;
        RECT 3.244 1.508 5.716 1.54 ;
  LAYER M2 ;
        RECT 3.244 1.572 5.716 1.604 ;
  LAYER M2 ;
        RECT 3.244 1.636 5.716 1.668 ;
  LAYER M2 ;
        RECT 3.244 1.7 5.716 1.732 ;
  LAYER M2 ;
        RECT 3.244 1.764 5.716 1.796 ;
  LAYER M2 ;
        RECT 3.244 1.828 5.716 1.86 ;
  LAYER M2 ;
        RECT 3.244 1.892 5.716 1.924 ;
  LAYER M2 ;
        RECT 3.244 1.956 5.716 1.988 ;
  LAYER M2 ;
        RECT 3.244 2.02 5.716 2.052 ;
  LAYER M2 ;
        RECT 3.244 2.084 5.716 2.116 ;
  LAYER M2 ;
        RECT 3.244 2.148 5.716 2.18 ;
  LAYER M2 ;
        RECT 3.244 2.212 5.716 2.244 ;
  LAYER M2 ;
        RECT 3.244 2.276 5.716 2.308 ;
  LAYER M2 ;
        RECT 3.244 2.34 5.716 2.372 ;
  LAYER M2 ;
        RECT 3.244 2.404 5.716 2.436 ;
  LAYER M2 ;
        RECT 3.244 2.468 5.716 2.5 ;
  LAYER M2 ;
        RECT 3.244 2.532 5.716 2.564 ;
  LAYER M2 ;
        RECT 3.244 2.596 5.716 2.628 ;
  LAYER M2 ;
        RECT 3.244 2.66 5.716 2.692 ;
  LAYER M2 ;
        RECT 3.244 2.724 5.716 2.756 ;
  LAYER M2 ;
        RECT 3.244 2.788 5.716 2.82 ;
  LAYER M2 ;
        RECT 3.244 2.852 5.716 2.884 ;
  LAYER M2 ;
        RECT 3.244 2.916 5.716 2.948 ;
  LAYER M2 ;
        RECT 3.244 2.98 5.716 3.012 ;
  LAYER M2 ;
        RECT 3.244 3.044 5.716 3.076 ;
  LAYER M3 ;
        RECT 3.264 0.72 3.296 3.228 ;
  LAYER M3 ;
        RECT 3.328 0.72 3.36 3.228 ;
  LAYER M3 ;
        RECT 3.392 0.72 3.424 3.228 ;
  LAYER M3 ;
        RECT 3.456 0.72 3.488 3.228 ;
  LAYER M3 ;
        RECT 3.52 0.72 3.552 3.228 ;
  LAYER M3 ;
        RECT 3.584 0.72 3.616 3.228 ;
  LAYER M3 ;
        RECT 3.648 0.72 3.68 3.228 ;
  LAYER M3 ;
        RECT 3.712 0.72 3.744 3.228 ;
  LAYER M3 ;
        RECT 3.776 0.72 3.808 3.228 ;
  LAYER M3 ;
        RECT 3.84 0.72 3.872 3.228 ;
  LAYER M3 ;
        RECT 3.904 0.72 3.936 3.228 ;
  LAYER M3 ;
        RECT 3.968 0.72 4 3.228 ;
  LAYER M3 ;
        RECT 4.032 0.72 4.064 3.228 ;
  LAYER M3 ;
        RECT 4.096 0.72 4.128 3.228 ;
  LAYER M3 ;
        RECT 4.16 0.72 4.192 3.228 ;
  LAYER M3 ;
        RECT 4.224 0.72 4.256 3.228 ;
  LAYER M3 ;
        RECT 4.288 0.72 4.32 3.228 ;
  LAYER M3 ;
        RECT 4.352 0.72 4.384 3.228 ;
  LAYER M3 ;
        RECT 4.416 0.72 4.448 3.228 ;
  LAYER M3 ;
        RECT 4.48 0.72 4.512 3.228 ;
  LAYER M3 ;
        RECT 4.544 0.72 4.576 3.228 ;
  LAYER M3 ;
        RECT 4.608 0.72 4.64 3.228 ;
  LAYER M3 ;
        RECT 4.672 0.72 4.704 3.228 ;
  LAYER M3 ;
        RECT 4.736 0.72 4.768 3.228 ;
  LAYER M3 ;
        RECT 4.8 0.72 4.832 3.228 ;
  LAYER M3 ;
        RECT 4.864 0.72 4.896 3.228 ;
  LAYER M3 ;
        RECT 4.928 0.72 4.96 3.228 ;
  LAYER M3 ;
        RECT 4.992 0.72 5.024 3.228 ;
  LAYER M3 ;
        RECT 5.056 0.72 5.088 3.228 ;
  LAYER M3 ;
        RECT 5.12 0.72 5.152 3.228 ;
  LAYER M3 ;
        RECT 5.184 0.72 5.216 3.228 ;
  LAYER M3 ;
        RECT 5.248 0.72 5.28 3.228 ;
  LAYER M3 ;
        RECT 5.312 0.72 5.344 3.228 ;
  LAYER M3 ;
        RECT 5.376 0.72 5.408 3.228 ;
  LAYER M3 ;
        RECT 5.44 0.72 5.472 3.228 ;
  LAYER M3 ;
        RECT 5.504 0.72 5.536 3.228 ;
  LAYER M3 ;
        RECT 5.568 0.72 5.6 3.228 ;
  LAYER M3 ;
        RECT 5.664 0.72 5.696 3.228 ;
  LAYER M1 ;
        RECT 3.279 0.756 3.281 3.192 ;
  LAYER M1 ;
        RECT 3.359 0.756 3.361 3.192 ;
  LAYER M1 ;
        RECT 3.439 0.756 3.441 3.192 ;
  LAYER M1 ;
        RECT 3.519 0.756 3.521 3.192 ;
  LAYER M1 ;
        RECT 3.599 0.756 3.601 3.192 ;
  LAYER M1 ;
        RECT 3.679 0.756 3.681 3.192 ;
  LAYER M1 ;
        RECT 3.759 0.756 3.761 3.192 ;
  LAYER M1 ;
        RECT 3.839 0.756 3.841 3.192 ;
  LAYER M1 ;
        RECT 3.919 0.756 3.921 3.192 ;
  LAYER M1 ;
        RECT 3.999 0.756 4.001 3.192 ;
  LAYER M1 ;
        RECT 4.079 0.756 4.081 3.192 ;
  LAYER M1 ;
        RECT 4.159 0.756 4.161 3.192 ;
  LAYER M1 ;
        RECT 4.239 0.756 4.241 3.192 ;
  LAYER M1 ;
        RECT 4.319 0.756 4.321 3.192 ;
  LAYER M1 ;
        RECT 4.399 0.756 4.401 3.192 ;
  LAYER M1 ;
        RECT 4.479 0.756 4.481 3.192 ;
  LAYER M1 ;
        RECT 4.559 0.756 4.561 3.192 ;
  LAYER M1 ;
        RECT 4.639 0.756 4.641 3.192 ;
  LAYER M1 ;
        RECT 4.719 0.756 4.721 3.192 ;
  LAYER M1 ;
        RECT 4.799 0.756 4.801 3.192 ;
  LAYER M1 ;
        RECT 4.879 0.756 4.881 3.192 ;
  LAYER M1 ;
        RECT 4.959 0.756 4.961 3.192 ;
  LAYER M1 ;
        RECT 5.039 0.756 5.041 3.192 ;
  LAYER M1 ;
        RECT 5.119 0.756 5.121 3.192 ;
  LAYER M1 ;
        RECT 5.199 0.756 5.201 3.192 ;
  LAYER M1 ;
        RECT 5.279 0.756 5.281 3.192 ;
  LAYER M1 ;
        RECT 5.359 0.756 5.361 3.192 ;
  LAYER M1 ;
        RECT 5.439 0.756 5.441 3.192 ;
  LAYER M1 ;
        RECT 5.519 0.756 5.521 3.192 ;
  LAYER M1 ;
        RECT 5.599 0.756 5.601 3.192 ;
  LAYER M2 ;
        RECT 3.28 0.755 5.68 0.757 ;
  LAYER M2 ;
        RECT 3.28 0.839 5.68 0.841 ;
  LAYER M2 ;
        RECT 3.28 0.923 5.68 0.925 ;
  LAYER M2 ;
        RECT 3.28 1.007 5.68 1.009 ;
  LAYER M2 ;
        RECT 3.28 1.091 5.68 1.093 ;
  LAYER M2 ;
        RECT 3.28 1.175 5.68 1.177 ;
  LAYER M2 ;
        RECT 3.28 1.259 5.68 1.261 ;
  LAYER M2 ;
        RECT 3.28 1.343 5.68 1.345 ;
  LAYER M2 ;
        RECT 3.28 1.427 5.68 1.429 ;
  LAYER M2 ;
        RECT 3.28 1.511 5.68 1.513 ;
  LAYER M2 ;
        RECT 3.28 1.595 5.68 1.597 ;
  LAYER M2 ;
        RECT 3.28 1.679 5.68 1.681 ;
  LAYER M2 ;
        RECT 3.28 1.7625 5.68 1.7645 ;
  LAYER M2 ;
        RECT 3.28 1.847 5.68 1.849 ;
  LAYER M2 ;
        RECT 3.28 1.931 5.68 1.933 ;
  LAYER M2 ;
        RECT 3.28 2.015 5.68 2.017 ;
  LAYER M2 ;
        RECT 3.28 2.099 5.68 2.101 ;
  LAYER M2 ;
        RECT 3.28 2.183 5.68 2.185 ;
  LAYER M2 ;
        RECT 3.28 2.267 5.68 2.269 ;
  LAYER M2 ;
        RECT 3.28 2.351 5.68 2.353 ;
  LAYER M2 ;
        RECT 3.28 2.435 5.68 2.437 ;
  LAYER M2 ;
        RECT 3.28 2.519 5.68 2.521 ;
  LAYER M2 ;
        RECT 3.28 2.603 5.68 2.605 ;
  LAYER M2 ;
        RECT 3.28 2.687 5.68 2.689 ;
  LAYER M2 ;
        RECT 3.28 2.771 5.68 2.773 ;
  LAYER M2 ;
        RECT 3.28 2.855 5.68 2.857 ;
  LAYER M2 ;
        RECT 3.28 2.939 5.68 2.941 ;
  LAYER M2 ;
        RECT 3.28 3.023 5.68 3.025 ;
  LAYER M2 ;
        RECT 3.28 3.107 5.68 3.109 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 6.168 ;
  LAYER M1 ;
        RECT 3.328 3.66 3.36 6.168 ;
  LAYER M1 ;
        RECT 3.392 3.66 3.424 6.168 ;
  LAYER M1 ;
        RECT 3.456 3.66 3.488 6.168 ;
  LAYER M1 ;
        RECT 3.52 3.66 3.552 6.168 ;
  LAYER M1 ;
        RECT 3.584 3.66 3.616 6.168 ;
  LAYER M1 ;
        RECT 3.648 3.66 3.68 6.168 ;
  LAYER M1 ;
        RECT 3.712 3.66 3.744 6.168 ;
  LAYER M1 ;
        RECT 3.776 3.66 3.808 6.168 ;
  LAYER M1 ;
        RECT 3.84 3.66 3.872 6.168 ;
  LAYER M1 ;
        RECT 3.904 3.66 3.936 6.168 ;
  LAYER M1 ;
        RECT 3.968 3.66 4 6.168 ;
  LAYER M1 ;
        RECT 4.032 3.66 4.064 6.168 ;
  LAYER M1 ;
        RECT 4.096 3.66 4.128 6.168 ;
  LAYER M1 ;
        RECT 4.16 3.66 4.192 6.168 ;
  LAYER M1 ;
        RECT 4.224 3.66 4.256 6.168 ;
  LAYER M1 ;
        RECT 4.288 3.66 4.32 6.168 ;
  LAYER M1 ;
        RECT 4.352 3.66 4.384 6.168 ;
  LAYER M1 ;
        RECT 4.416 3.66 4.448 6.168 ;
  LAYER M1 ;
        RECT 4.48 3.66 4.512 6.168 ;
  LAYER M1 ;
        RECT 4.544 3.66 4.576 6.168 ;
  LAYER M1 ;
        RECT 4.608 3.66 4.64 6.168 ;
  LAYER M1 ;
        RECT 4.672 3.66 4.704 6.168 ;
  LAYER M1 ;
        RECT 4.736 3.66 4.768 6.168 ;
  LAYER M1 ;
        RECT 4.8 3.66 4.832 6.168 ;
  LAYER M1 ;
        RECT 4.864 3.66 4.896 6.168 ;
  LAYER M1 ;
        RECT 4.928 3.66 4.96 6.168 ;
  LAYER M1 ;
        RECT 4.992 3.66 5.024 6.168 ;
  LAYER M1 ;
        RECT 5.056 3.66 5.088 6.168 ;
  LAYER M1 ;
        RECT 5.12 3.66 5.152 6.168 ;
  LAYER M1 ;
        RECT 5.184 3.66 5.216 6.168 ;
  LAYER M1 ;
        RECT 5.248 3.66 5.28 6.168 ;
  LAYER M1 ;
        RECT 5.312 3.66 5.344 6.168 ;
  LAYER M1 ;
        RECT 5.376 3.66 5.408 6.168 ;
  LAYER M1 ;
        RECT 5.44 3.66 5.472 6.168 ;
  LAYER M1 ;
        RECT 5.504 3.66 5.536 6.168 ;
  LAYER M1 ;
        RECT 5.568 3.66 5.6 6.168 ;
  LAYER M2 ;
        RECT 3.244 3.744 5.716 3.776 ;
  LAYER M2 ;
        RECT 3.244 3.808 5.716 3.84 ;
  LAYER M2 ;
        RECT 3.244 3.872 5.716 3.904 ;
  LAYER M2 ;
        RECT 3.244 3.936 5.716 3.968 ;
  LAYER M2 ;
        RECT 3.244 4 5.716 4.032 ;
  LAYER M2 ;
        RECT 3.244 4.064 5.716 4.096 ;
  LAYER M2 ;
        RECT 3.244 4.128 5.716 4.16 ;
  LAYER M2 ;
        RECT 3.244 4.192 5.716 4.224 ;
  LAYER M2 ;
        RECT 3.244 4.256 5.716 4.288 ;
  LAYER M2 ;
        RECT 3.244 4.32 5.716 4.352 ;
  LAYER M2 ;
        RECT 3.244 4.384 5.716 4.416 ;
  LAYER M2 ;
        RECT 3.244 4.448 5.716 4.48 ;
  LAYER M2 ;
        RECT 3.244 4.512 5.716 4.544 ;
  LAYER M2 ;
        RECT 3.244 4.576 5.716 4.608 ;
  LAYER M2 ;
        RECT 3.244 4.64 5.716 4.672 ;
  LAYER M2 ;
        RECT 3.244 4.704 5.716 4.736 ;
  LAYER M2 ;
        RECT 3.244 4.768 5.716 4.8 ;
  LAYER M2 ;
        RECT 3.244 4.832 5.716 4.864 ;
  LAYER M2 ;
        RECT 3.244 4.896 5.716 4.928 ;
  LAYER M2 ;
        RECT 3.244 4.96 5.716 4.992 ;
  LAYER M2 ;
        RECT 3.244 5.024 5.716 5.056 ;
  LAYER M2 ;
        RECT 3.244 5.088 5.716 5.12 ;
  LAYER M2 ;
        RECT 3.244 5.152 5.716 5.184 ;
  LAYER M2 ;
        RECT 3.244 5.216 5.716 5.248 ;
  LAYER M2 ;
        RECT 3.244 5.28 5.716 5.312 ;
  LAYER M2 ;
        RECT 3.244 5.344 5.716 5.376 ;
  LAYER M2 ;
        RECT 3.244 5.408 5.716 5.44 ;
  LAYER M2 ;
        RECT 3.244 5.472 5.716 5.504 ;
  LAYER M2 ;
        RECT 3.244 5.536 5.716 5.568 ;
  LAYER M2 ;
        RECT 3.244 5.6 5.716 5.632 ;
  LAYER M2 ;
        RECT 3.244 5.664 5.716 5.696 ;
  LAYER M2 ;
        RECT 3.244 5.728 5.716 5.76 ;
  LAYER M2 ;
        RECT 3.244 5.792 5.716 5.824 ;
  LAYER M2 ;
        RECT 3.244 5.856 5.716 5.888 ;
  LAYER M2 ;
        RECT 3.244 5.92 5.716 5.952 ;
  LAYER M2 ;
        RECT 3.244 5.984 5.716 6.016 ;
  LAYER M3 ;
        RECT 3.264 3.66 3.296 6.168 ;
  LAYER M3 ;
        RECT 3.328 3.66 3.36 6.168 ;
  LAYER M3 ;
        RECT 3.392 3.66 3.424 6.168 ;
  LAYER M3 ;
        RECT 3.456 3.66 3.488 6.168 ;
  LAYER M3 ;
        RECT 3.52 3.66 3.552 6.168 ;
  LAYER M3 ;
        RECT 3.584 3.66 3.616 6.168 ;
  LAYER M3 ;
        RECT 3.648 3.66 3.68 6.168 ;
  LAYER M3 ;
        RECT 3.712 3.66 3.744 6.168 ;
  LAYER M3 ;
        RECT 3.776 3.66 3.808 6.168 ;
  LAYER M3 ;
        RECT 3.84 3.66 3.872 6.168 ;
  LAYER M3 ;
        RECT 3.904 3.66 3.936 6.168 ;
  LAYER M3 ;
        RECT 3.968 3.66 4 6.168 ;
  LAYER M3 ;
        RECT 4.032 3.66 4.064 6.168 ;
  LAYER M3 ;
        RECT 4.096 3.66 4.128 6.168 ;
  LAYER M3 ;
        RECT 4.16 3.66 4.192 6.168 ;
  LAYER M3 ;
        RECT 4.224 3.66 4.256 6.168 ;
  LAYER M3 ;
        RECT 4.288 3.66 4.32 6.168 ;
  LAYER M3 ;
        RECT 4.352 3.66 4.384 6.168 ;
  LAYER M3 ;
        RECT 4.416 3.66 4.448 6.168 ;
  LAYER M3 ;
        RECT 4.48 3.66 4.512 6.168 ;
  LAYER M3 ;
        RECT 4.544 3.66 4.576 6.168 ;
  LAYER M3 ;
        RECT 4.608 3.66 4.64 6.168 ;
  LAYER M3 ;
        RECT 4.672 3.66 4.704 6.168 ;
  LAYER M3 ;
        RECT 4.736 3.66 4.768 6.168 ;
  LAYER M3 ;
        RECT 4.8 3.66 4.832 6.168 ;
  LAYER M3 ;
        RECT 4.864 3.66 4.896 6.168 ;
  LAYER M3 ;
        RECT 4.928 3.66 4.96 6.168 ;
  LAYER M3 ;
        RECT 4.992 3.66 5.024 6.168 ;
  LAYER M3 ;
        RECT 5.056 3.66 5.088 6.168 ;
  LAYER M3 ;
        RECT 5.12 3.66 5.152 6.168 ;
  LAYER M3 ;
        RECT 5.184 3.66 5.216 6.168 ;
  LAYER M3 ;
        RECT 5.248 3.66 5.28 6.168 ;
  LAYER M3 ;
        RECT 5.312 3.66 5.344 6.168 ;
  LAYER M3 ;
        RECT 5.376 3.66 5.408 6.168 ;
  LAYER M3 ;
        RECT 5.44 3.66 5.472 6.168 ;
  LAYER M3 ;
        RECT 5.504 3.66 5.536 6.168 ;
  LAYER M3 ;
        RECT 5.568 3.66 5.6 6.168 ;
  LAYER M3 ;
        RECT 5.664 3.66 5.696 6.168 ;
  LAYER M1 ;
        RECT 3.279 3.696 3.281 6.132 ;
  LAYER M1 ;
        RECT 3.359 3.696 3.361 6.132 ;
  LAYER M1 ;
        RECT 3.439 3.696 3.441 6.132 ;
  LAYER M1 ;
        RECT 3.519 3.696 3.521 6.132 ;
  LAYER M1 ;
        RECT 3.599 3.696 3.601 6.132 ;
  LAYER M1 ;
        RECT 3.679 3.696 3.681 6.132 ;
  LAYER M1 ;
        RECT 3.759 3.696 3.761 6.132 ;
  LAYER M1 ;
        RECT 3.839 3.696 3.841 6.132 ;
  LAYER M1 ;
        RECT 3.919 3.696 3.921 6.132 ;
  LAYER M1 ;
        RECT 3.999 3.696 4.001 6.132 ;
  LAYER M1 ;
        RECT 4.079 3.696 4.081 6.132 ;
  LAYER M1 ;
        RECT 4.159 3.696 4.161 6.132 ;
  LAYER M1 ;
        RECT 4.239 3.696 4.241 6.132 ;
  LAYER M1 ;
        RECT 4.319 3.696 4.321 6.132 ;
  LAYER M1 ;
        RECT 4.399 3.696 4.401 6.132 ;
  LAYER M1 ;
        RECT 4.479 3.696 4.481 6.132 ;
  LAYER M1 ;
        RECT 4.559 3.696 4.561 6.132 ;
  LAYER M1 ;
        RECT 4.639 3.696 4.641 6.132 ;
  LAYER M1 ;
        RECT 4.719 3.696 4.721 6.132 ;
  LAYER M1 ;
        RECT 4.799 3.696 4.801 6.132 ;
  LAYER M1 ;
        RECT 4.879 3.696 4.881 6.132 ;
  LAYER M1 ;
        RECT 4.959 3.696 4.961 6.132 ;
  LAYER M1 ;
        RECT 5.039 3.696 5.041 6.132 ;
  LAYER M1 ;
        RECT 5.119 3.696 5.121 6.132 ;
  LAYER M1 ;
        RECT 5.199 3.696 5.201 6.132 ;
  LAYER M1 ;
        RECT 5.279 3.696 5.281 6.132 ;
  LAYER M1 ;
        RECT 5.359 3.696 5.361 6.132 ;
  LAYER M1 ;
        RECT 5.439 3.696 5.441 6.132 ;
  LAYER M1 ;
        RECT 5.519 3.696 5.521 6.132 ;
  LAYER M1 ;
        RECT 5.599 3.696 5.601 6.132 ;
  LAYER M2 ;
        RECT 3.28 3.695 5.68 3.697 ;
  LAYER M2 ;
        RECT 3.28 3.779 5.68 3.781 ;
  LAYER M2 ;
        RECT 3.28 3.863 5.68 3.865 ;
  LAYER M2 ;
        RECT 3.28 3.947 5.68 3.949 ;
  LAYER M2 ;
        RECT 3.28 4.031 5.68 4.033 ;
  LAYER M2 ;
        RECT 3.28 4.115 5.68 4.117 ;
  LAYER M2 ;
        RECT 3.28 4.199 5.68 4.201 ;
  LAYER M2 ;
        RECT 3.28 4.283 5.68 4.285 ;
  LAYER M2 ;
        RECT 3.28 4.367 5.68 4.369 ;
  LAYER M2 ;
        RECT 3.28 4.451 5.68 4.453 ;
  LAYER M2 ;
        RECT 3.28 4.535 5.68 4.537 ;
  LAYER M2 ;
        RECT 3.28 4.619 5.68 4.621 ;
  LAYER M2 ;
        RECT 3.28 4.7025 5.68 4.7045 ;
  LAYER M2 ;
        RECT 3.28 4.787 5.68 4.789 ;
  LAYER M2 ;
        RECT 3.28 4.871 5.68 4.873 ;
  LAYER M2 ;
        RECT 3.28 4.955 5.68 4.957 ;
  LAYER M2 ;
        RECT 3.28 5.039 5.68 5.041 ;
  LAYER M2 ;
        RECT 3.28 5.123 5.68 5.125 ;
  LAYER M2 ;
        RECT 3.28 5.207 5.68 5.209 ;
  LAYER M2 ;
        RECT 3.28 5.291 5.68 5.293 ;
  LAYER M2 ;
        RECT 3.28 5.375 5.68 5.377 ;
  LAYER M2 ;
        RECT 3.28 5.459 5.68 5.461 ;
  LAYER M2 ;
        RECT 3.28 5.543 5.68 5.545 ;
  LAYER M2 ;
        RECT 3.28 5.627 5.68 5.629 ;
  LAYER M2 ;
        RECT 3.28 5.711 5.68 5.713 ;
  LAYER M2 ;
        RECT 3.28 5.795 5.68 5.797 ;
  LAYER M2 ;
        RECT 3.28 5.879 5.68 5.881 ;
  LAYER M2 ;
        RECT 3.28 5.963 5.68 5.965 ;
  LAYER M2 ;
        RECT 3.28 6.047 5.68 6.049 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 9.108 ;
  LAYER M1 ;
        RECT 3.328 6.6 3.36 9.108 ;
  LAYER M1 ;
        RECT 3.392 6.6 3.424 9.108 ;
  LAYER M1 ;
        RECT 3.456 6.6 3.488 9.108 ;
  LAYER M1 ;
        RECT 3.52 6.6 3.552 9.108 ;
  LAYER M1 ;
        RECT 3.584 6.6 3.616 9.108 ;
  LAYER M1 ;
        RECT 3.648 6.6 3.68 9.108 ;
  LAYER M1 ;
        RECT 3.712 6.6 3.744 9.108 ;
  LAYER M1 ;
        RECT 3.776 6.6 3.808 9.108 ;
  LAYER M1 ;
        RECT 3.84 6.6 3.872 9.108 ;
  LAYER M1 ;
        RECT 3.904 6.6 3.936 9.108 ;
  LAYER M1 ;
        RECT 3.968 6.6 4 9.108 ;
  LAYER M1 ;
        RECT 4.032 6.6 4.064 9.108 ;
  LAYER M1 ;
        RECT 4.096 6.6 4.128 9.108 ;
  LAYER M1 ;
        RECT 4.16 6.6 4.192 9.108 ;
  LAYER M1 ;
        RECT 4.224 6.6 4.256 9.108 ;
  LAYER M1 ;
        RECT 4.288 6.6 4.32 9.108 ;
  LAYER M1 ;
        RECT 4.352 6.6 4.384 9.108 ;
  LAYER M1 ;
        RECT 4.416 6.6 4.448 9.108 ;
  LAYER M1 ;
        RECT 4.48 6.6 4.512 9.108 ;
  LAYER M1 ;
        RECT 4.544 6.6 4.576 9.108 ;
  LAYER M1 ;
        RECT 4.608 6.6 4.64 9.108 ;
  LAYER M1 ;
        RECT 4.672 6.6 4.704 9.108 ;
  LAYER M1 ;
        RECT 4.736 6.6 4.768 9.108 ;
  LAYER M1 ;
        RECT 4.8 6.6 4.832 9.108 ;
  LAYER M1 ;
        RECT 4.864 6.6 4.896 9.108 ;
  LAYER M1 ;
        RECT 4.928 6.6 4.96 9.108 ;
  LAYER M1 ;
        RECT 4.992 6.6 5.024 9.108 ;
  LAYER M1 ;
        RECT 5.056 6.6 5.088 9.108 ;
  LAYER M1 ;
        RECT 5.12 6.6 5.152 9.108 ;
  LAYER M1 ;
        RECT 5.184 6.6 5.216 9.108 ;
  LAYER M1 ;
        RECT 5.248 6.6 5.28 9.108 ;
  LAYER M1 ;
        RECT 5.312 6.6 5.344 9.108 ;
  LAYER M1 ;
        RECT 5.376 6.6 5.408 9.108 ;
  LAYER M1 ;
        RECT 5.44 6.6 5.472 9.108 ;
  LAYER M1 ;
        RECT 5.504 6.6 5.536 9.108 ;
  LAYER M1 ;
        RECT 5.568 6.6 5.6 9.108 ;
  LAYER M2 ;
        RECT 3.244 6.684 5.716 6.716 ;
  LAYER M2 ;
        RECT 3.244 6.748 5.716 6.78 ;
  LAYER M2 ;
        RECT 3.244 6.812 5.716 6.844 ;
  LAYER M2 ;
        RECT 3.244 6.876 5.716 6.908 ;
  LAYER M2 ;
        RECT 3.244 6.94 5.716 6.972 ;
  LAYER M2 ;
        RECT 3.244 7.004 5.716 7.036 ;
  LAYER M2 ;
        RECT 3.244 7.068 5.716 7.1 ;
  LAYER M2 ;
        RECT 3.244 7.132 5.716 7.164 ;
  LAYER M2 ;
        RECT 3.244 7.196 5.716 7.228 ;
  LAYER M2 ;
        RECT 3.244 7.26 5.716 7.292 ;
  LAYER M2 ;
        RECT 3.244 7.324 5.716 7.356 ;
  LAYER M2 ;
        RECT 3.244 7.388 5.716 7.42 ;
  LAYER M2 ;
        RECT 3.244 7.452 5.716 7.484 ;
  LAYER M2 ;
        RECT 3.244 7.516 5.716 7.548 ;
  LAYER M2 ;
        RECT 3.244 7.58 5.716 7.612 ;
  LAYER M2 ;
        RECT 3.244 7.644 5.716 7.676 ;
  LAYER M2 ;
        RECT 3.244 7.708 5.716 7.74 ;
  LAYER M2 ;
        RECT 3.244 7.772 5.716 7.804 ;
  LAYER M2 ;
        RECT 3.244 7.836 5.716 7.868 ;
  LAYER M2 ;
        RECT 3.244 7.9 5.716 7.932 ;
  LAYER M2 ;
        RECT 3.244 7.964 5.716 7.996 ;
  LAYER M2 ;
        RECT 3.244 8.028 5.716 8.06 ;
  LAYER M2 ;
        RECT 3.244 8.092 5.716 8.124 ;
  LAYER M2 ;
        RECT 3.244 8.156 5.716 8.188 ;
  LAYER M2 ;
        RECT 3.244 8.22 5.716 8.252 ;
  LAYER M2 ;
        RECT 3.244 8.284 5.716 8.316 ;
  LAYER M2 ;
        RECT 3.244 8.348 5.716 8.38 ;
  LAYER M2 ;
        RECT 3.244 8.412 5.716 8.444 ;
  LAYER M2 ;
        RECT 3.244 8.476 5.716 8.508 ;
  LAYER M2 ;
        RECT 3.244 8.54 5.716 8.572 ;
  LAYER M2 ;
        RECT 3.244 8.604 5.716 8.636 ;
  LAYER M2 ;
        RECT 3.244 8.668 5.716 8.7 ;
  LAYER M2 ;
        RECT 3.244 8.732 5.716 8.764 ;
  LAYER M2 ;
        RECT 3.244 8.796 5.716 8.828 ;
  LAYER M2 ;
        RECT 3.244 8.86 5.716 8.892 ;
  LAYER M2 ;
        RECT 3.244 8.924 5.716 8.956 ;
  LAYER M3 ;
        RECT 3.264 6.6 3.296 9.108 ;
  LAYER M3 ;
        RECT 3.328 6.6 3.36 9.108 ;
  LAYER M3 ;
        RECT 3.392 6.6 3.424 9.108 ;
  LAYER M3 ;
        RECT 3.456 6.6 3.488 9.108 ;
  LAYER M3 ;
        RECT 3.52 6.6 3.552 9.108 ;
  LAYER M3 ;
        RECT 3.584 6.6 3.616 9.108 ;
  LAYER M3 ;
        RECT 3.648 6.6 3.68 9.108 ;
  LAYER M3 ;
        RECT 3.712 6.6 3.744 9.108 ;
  LAYER M3 ;
        RECT 3.776 6.6 3.808 9.108 ;
  LAYER M3 ;
        RECT 3.84 6.6 3.872 9.108 ;
  LAYER M3 ;
        RECT 3.904 6.6 3.936 9.108 ;
  LAYER M3 ;
        RECT 3.968 6.6 4 9.108 ;
  LAYER M3 ;
        RECT 4.032 6.6 4.064 9.108 ;
  LAYER M3 ;
        RECT 4.096 6.6 4.128 9.108 ;
  LAYER M3 ;
        RECT 4.16 6.6 4.192 9.108 ;
  LAYER M3 ;
        RECT 4.224 6.6 4.256 9.108 ;
  LAYER M3 ;
        RECT 4.288 6.6 4.32 9.108 ;
  LAYER M3 ;
        RECT 4.352 6.6 4.384 9.108 ;
  LAYER M3 ;
        RECT 4.416 6.6 4.448 9.108 ;
  LAYER M3 ;
        RECT 4.48 6.6 4.512 9.108 ;
  LAYER M3 ;
        RECT 4.544 6.6 4.576 9.108 ;
  LAYER M3 ;
        RECT 4.608 6.6 4.64 9.108 ;
  LAYER M3 ;
        RECT 4.672 6.6 4.704 9.108 ;
  LAYER M3 ;
        RECT 4.736 6.6 4.768 9.108 ;
  LAYER M3 ;
        RECT 4.8 6.6 4.832 9.108 ;
  LAYER M3 ;
        RECT 4.864 6.6 4.896 9.108 ;
  LAYER M3 ;
        RECT 4.928 6.6 4.96 9.108 ;
  LAYER M3 ;
        RECT 4.992 6.6 5.024 9.108 ;
  LAYER M3 ;
        RECT 5.056 6.6 5.088 9.108 ;
  LAYER M3 ;
        RECT 5.12 6.6 5.152 9.108 ;
  LAYER M3 ;
        RECT 5.184 6.6 5.216 9.108 ;
  LAYER M3 ;
        RECT 5.248 6.6 5.28 9.108 ;
  LAYER M3 ;
        RECT 5.312 6.6 5.344 9.108 ;
  LAYER M3 ;
        RECT 5.376 6.6 5.408 9.108 ;
  LAYER M3 ;
        RECT 5.44 6.6 5.472 9.108 ;
  LAYER M3 ;
        RECT 5.504 6.6 5.536 9.108 ;
  LAYER M3 ;
        RECT 5.568 6.6 5.6 9.108 ;
  LAYER M3 ;
        RECT 5.664 6.6 5.696 9.108 ;
  LAYER M1 ;
        RECT 3.279 6.636 3.281 9.072 ;
  LAYER M1 ;
        RECT 3.359 6.636 3.361 9.072 ;
  LAYER M1 ;
        RECT 3.439 6.636 3.441 9.072 ;
  LAYER M1 ;
        RECT 3.519 6.636 3.521 9.072 ;
  LAYER M1 ;
        RECT 3.599 6.636 3.601 9.072 ;
  LAYER M1 ;
        RECT 3.679 6.636 3.681 9.072 ;
  LAYER M1 ;
        RECT 3.759 6.636 3.761 9.072 ;
  LAYER M1 ;
        RECT 3.839 6.636 3.841 9.072 ;
  LAYER M1 ;
        RECT 3.919 6.636 3.921 9.072 ;
  LAYER M1 ;
        RECT 3.999 6.636 4.001 9.072 ;
  LAYER M1 ;
        RECT 4.079 6.636 4.081 9.072 ;
  LAYER M1 ;
        RECT 4.159 6.636 4.161 9.072 ;
  LAYER M1 ;
        RECT 4.239 6.636 4.241 9.072 ;
  LAYER M1 ;
        RECT 4.319 6.636 4.321 9.072 ;
  LAYER M1 ;
        RECT 4.399 6.636 4.401 9.072 ;
  LAYER M1 ;
        RECT 4.479 6.636 4.481 9.072 ;
  LAYER M1 ;
        RECT 4.559 6.636 4.561 9.072 ;
  LAYER M1 ;
        RECT 4.639 6.636 4.641 9.072 ;
  LAYER M1 ;
        RECT 4.719 6.636 4.721 9.072 ;
  LAYER M1 ;
        RECT 4.799 6.636 4.801 9.072 ;
  LAYER M1 ;
        RECT 4.879 6.636 4.881 9.072 ;
  LAYER M1 ;
        RECT 4.959 6.636 4.961 9.072 ;
  LAYER M1 ;
        RECT 5.039 6.636 5.041 9.072 ;
  LAYER M1 ;
        RECT 5.119 6.636 5.121 9.072 ;
  LAYER M1 ;
        RECT 5.199 6.636 5.201 9.072 ;
  LAYER M1 ;
        RECT 5.279 6.636 5.281 9.072 ;
  LAYER M1 ;
        RECT 5.359 6.636 5.361 9.072 ;
  LAYER M1 ;
        RECT 5.439 6.636 5.441 9.072 ;
  LAYER M1 ;
        RECT 5.519 6.636 5.521 9.072 ;
  LAYER M1 ;
        RECT 5.599 6.636 5.601 9.072 ;
  LAYER M2 ;
        RECT 3.28 6.635 5.68 6.637 ;
  LAYER M2 ;
        RECT 3.28 6.719 5.68 6.721 ;
  LAYER M2 ;
        RECT 3.28 6.803 5.68 6.805 ;
  LAYER M2 ;
        RECT 3.28 6.887 5.68 6.889 ;
  LAYER M2 ;
        RECT 3.28 6.971 5.68 6.973 ;
  LAYER M2 ;
        RECT 3.28 7.055 5.68 7.057 ;
  LAYER M2 ;
        RECT 3.28 7.139 5.68 7.141 ;
  LAYER M2 ;
        RECT 3.28 7.223 5.68 7.225 ;
  LAYER M2 ;
        RECT 3.28 7.307 5.68 7.309 ;
  LAYER M2 ;
        RECT 3.28 7.391 5.68 7.393 ;
  LAYER M2 ;
        RECT 3.28 7.475 5.68 7.477 ;
  LAYER M2 ;
        RECT 3.28 7.559 5.68 7.561 ;
  LAYER M2 ;
        RECT 3.28 7.6425 5.68 7.6445 ;
  LAYER M2 ;
        RECT 3.28 7.727 5.68 7.729 ;
  LAYER M2 ;
        RECT 3.28 7.811 5.68 7.813 ;
  LAYER M2 ;
        RECT 3.28 7.895 5.68 7.897 ;
  LAYER M2 ;
        RECT 3.28 7.979 5.68 7.981 ;
  LAYER M2 ;
        RECT 3.28 8.063 5.68 8.065 ;
  LAYER M2 ;
        RECT 3.28 8.147 5.68 8.149 ;
  LAYER M2 ;
        RECT 3.28 8.231 5.68 8.233 ;
  LAYER M2 ;
        RECT 3.28 8.315 5.68 8.317 ;
  LAYER M2 ;
        RECT 3.28 8.399 5.68 8.401 ;
  LAYER M2 ;
        RECT 3.28 8.483 5.68 8.485 ;
  LAYER M2 ;
        RECT 3.28 8.567 5.68 8.569 ;
  LAYER M2 ;
        RECT 3.28 8.651 5.68 8.653 ;
  LAYER M2 ;
        RECT 3.28 8.735 5.68 8.737 ;
  LAYER M2 ;
        RECT 3.28 8.819 5.68 8.821 ;
  LAYER M2 ;
        RECT 3.28 8.903 5.68 8.905 ;
  LAYER M2 ;
        RECT 3.28 8.987 5.68 8.989 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 12.048 ;
  LAYER M1 ;
        RECT 3.328 9.54 3.36 12.048 ;
  LAYER M1 ;
        RECT 3.392 9.54 3.424 12.048 ;
  LAYER M1 ;
        RECT 3.456 9.54 3.488 12.048 ;
  LAYER M1 ;
        RECT 3.52 9.54 3.552 12.048 ;
  LAYER M1 ;
        RECT 3.584 9.54 3.616 12.048 ;
  LAYER M1 ;
        RECT 3.648 9.54 3.68 12.048 ;
  LAYER M1 ;
        RECT 3.712 9.54 3.744 12.048 ;
  LAYER M1 ;
        RECT 3.776 9.54 3.808 12.048 ;
  LAYER M1 ;
        RECT 3.84 9.54 3.872 12.048 ;
  LAYER M1 ;
        RECT 3.904 9.54 3.936 12.048 ;
  LAYER M1 ;
        RECT 3.968 9.54 4 12.048 ;
  LAYER M1 ;
        RECT 4.032 9.54 4.064 12.048 ;
  LAYER M1 ;
        RECT 4.096 9.54 4.128 12.048 ;
  LAYER M1 ;
        RECT 4.16 9.54 4.192 12.048 ;
  LAYER M1 ;
        RECT 4.224 9.54 4.256 12.048 ;
  LAYER M1 ;
        RECT 4.288 9.54 4.32 12.048 ;
  LAYER M1 ;
        RECT 4.352 9.54 4.384 12.048 ;
  LAYER M1 ;
        RECT 4.416 9.54 4.448 12.048 ;
  LAYER M1 ;
        RECT 4.48 9.54 4.512 12.048 ;
  LAYER M1 ;
        RECT 4.544 9.54 4.576 12.048 ;
  LAYER M1 ;
        RECT 4.608 9.54 4.64 12.048 ;
  LAYER M1 ;
        RECT 4.672 9.54 4.704 12.048 ;
  LAYER M1 ;
        RECT 4.736 9.54 4.768 12.048 ;
  LAYER M1 ;
        RECT 4.8 9.54 4.832 12.048 ;
  LAYER M1 ;
        RECT 4.864 9.54 4.896 12.048 ;
  LAYER M1 ;
        RECT 4.928 9.54 4.96 12.048 ;
  LAYER M1 ;
        RECT 4.992 9.54 5.024 12.048 ;
  LAYER M1 ;
        RECT 5.056 9.54 5.088 12.048 ;
  LAYER M1 ;
        RECT 5.12 9.54 5.152 12.048 ;
  LAYER M1 ;
        RECT 5.184 9.54 5.216 12.048 ;
  LAYER M1 ;
        RECT 5.248 9.54 5.28 12.048 ;
  LAYER M1 ;
        RECT 5.312 9.54 5.344 12.048 ;
  LAYER M1 ;
        RECT 5.376 9.54 5.408 12.048 ;
  LAYER M1 ;
        RECT 5.44 9.54 5.472 12.048 ;
  LAYER M1 ;
        RECT 5.504 9.54 5.536 12.048 ;
  LAYER M1 ;
        RECT 5.568 9.54 5.6 12.048 ;
  LAYER M2 ;
        RECT 3.244 9.624 5.716 9.656 ;
  LAYER M2 ;
        RECT 3.244 9.688 5.716 9.72 ;
  LAYER M2 ;
        RECT 3.244 9.752 5.716 9.784 ;
  LAYER M2 ;
        RECT 3.244 9.816 5.716 9.848 ;
  LAYER M2 ;
        RECT 3.244 9.88 5.716 9.912 ;
  LAYER M2 ;
        RECT 3.244 9.944 5.716 9.976 ;
  LAYER M2 ;
        RECT 3.244 10.008 5.716 10.04 ;
  LAYER M2 ;
        RECT 3.244 10.072 5.716 10.104 ;
  LAYER M2 ;
        RECT 3.244 10.136 5.716 10.168 ;
  LAYER M2 ;
        RECT 3.244 10.2 5.716 10.232 ;
  LAYER M2 ;
        RECT 3.244 10.264 5.716 10.296 ;
  LAYER M2 ;
        RECT 3.244 10.328 5.716 10.36 ;
  LAYER M2 ;
        RECT 3.244 10.392 5.716 10.424 ;
  LAYER M2 ;
        RECT 3.244 10.456 5.716 10.488 ;
  LAYER M2 ;
        RECT 3.244 10.52 5.716 10.552 ;
  LAYER M2 ;
        RECT 3.244 10.584 5.716 10.616 ;
  LAYER M2 ;
        RECT 3.244 10.648 5.716 10.68 ;
  LAYER M2 ;
        RECT 3.244 10.712 5.716 10.744 ;
  LAYER M2 ;
        RECT 3.244 10.776 5.716 10.808 ;
  LAYER M2 ;
        RECT 3.244 10.84 5.716 10.872 ;
  LAYER M2 ;
        RECT 3.244 10.904 5.716 10.936 ;
  LAYER M2 ;
        RECT 3.244 10.968 5.716 11 ;
  LAYER M2 ;
        RECT 3.244 11.032 5.716 11.064 ;
  LAYER M2 ;
        RECT 3.244 11.096 5.716 11.128 ;
  LAYER M2 ;
        RECT 3.244 11.16 5.716 11.192 ;
  LAYER M2 ;
        RECT 3.244 11.224 5.716 11.256 ;
  LAYER M2 ;
        RECT 3.244 11.288 5.716 11.32 ;
  LAYER M2 ;
        RECT 3.244 11.352 5.716 11.384 ;
  LAYER M2 ;
        RECT 3.244 11.416 5.716 11.448 ;
  LAYER M2 ;
        RECT 3.244 11.48 5.716 11.512 ;
  LAYER M2 ;
        RECT 3.244 11.544 5.716 11.576 ;
  LAYER M2 ;
        RECT 3.244 11.608 5.716 11.64 ;
  LAYER M2 ;
        RECT 3.244 11.672 5.716 11.704 ;
  LAYER M2 ;
        RECT 3.244 11.736 5.716 11.768 ;
  LAYER M2 ;
        RECT 3.244 11.8 5.716 11.832 ;
  LAYER M2 ;
        RECT 3.244 11.864 5.716 11.896 ;
  LAYER M3 ;
        RECT 3.264 9.54 3.296 12.048 ;
  LAYER M3 ;
        RECT 3.328 9.54 3.36 12.048 ;
  LAYER M3 ;
        RECT 3.392 9.54 3.424 12.048 ;
  LAYER M3 ;
        RECT 3.456 9.54 3.488 12.048 ;
  LAYER M3 ;
        RECT 3.52 9.54 3.552 12.048 ;
  LAYER M3 ;
        RECT 3.584 9.54 3.616 12.048 ;
  LAYER M3 ;
        RECT 3.648 9.54 3.68 12.048 ;
  LAYER M3 ;
        RECT 3.712 9.54 3.744 12.048 ;
  LAYER M3 ;
        RECT 3.776 9.54 3.808 12.048 ;
  LAYER M3 ;
        RECT 3.84 9.54 3.872 12.048 ;
  LAYER M3 ;
        RECT 3.904 9.54 3.936 12.048 ;
  LAYER M3 ;
        RECT 3.968 9.54 4 12.048 ;
  LAYER M3 ;
        RECT 4.032 9.54 4.064 12.048 ;
  LAYER M3 ;
        RECT 4.096 9.54 4.128 12.048 ;
  LAYER M3 ;
        RECT 4.16 9.54 4.192 12.048 ;
  LAYER M3 ;
        RECT 4.224 9.54 4.256 12.048 ;
  LAYER M3 ;
        RECT 4.288 9.54 4.32 12.048 ;
  LAYER M3 ;
        RECT 4.352 9.54 4.384 12.048 ;
  LAYER M3 ;
        RECT 4.416 9.54 4.448 12.048 ;
  LAYER M3 ;
        RECT 4.48 9.54 4.512 12.048 ;
  LAYER M3 ;
        RECT 4.544 9.54 4.576 12.048 ;
  LAYER M3 ;
        RECT 4.608 9.54 4.64 12.048 ;
  LAYER M3 ;
        RECT 4.672 9.54 4.704 12.048 ;
  LAYER M3 ;
        RECT 4.736 9.54 4.768 12.048 ;
  LAYER M3 ;
        RECT 4.8 9.54 4.832 12.048 ;
  LAYER M3 ;
        RECT 4.864 9.54 4.896 12.048 ;
  LAYER M3 ;
        RECT 4.928 9.54 4.96 12.048 ;
  LAYER M3 ;
        RECT 4.992 9.54 5.024 12.048 ;
  LAYER M3 ;
        RECT 5.056 9.54 5.088 12.048 ;
  LAYER M3 ;
        RECT 5.12 9.54 5.152 12.048 ;
  LAYER M3 ;
        RECT 5.184 9.54 5.216 12.048 ;
  LAYER M3 ;
        RECT 5.248 9.54 5.28 12.048 ;
  LAYER M3 ;
        RECT 5.312 9.54 5.344 12.048 ;
  LAYER M3 ;
        RECT 5.376 9.54 5.408 12.048 ;
  LAYER M3 ;
        RECT 5.44 9.54 5.472 12.048 ;
  LAYER M3 ;
        RECT 5.504 9.54 5.536 12.048 ;
  LAYER M3 ;
        RECT 5.568 9.54 5.6 12.048 ;
  LAYER M3 ;
        RECT 5.664 9.54 5.696 12.048 ;
  LAYER M1 ;
        RECT 3.279 9.576 3.281 12.012 ;
  LAYER M1 ;
        RECT 3.359 9.576 3.361 12.012 ;
  LAYER M1 ;
        RECT 3.439 9.576 3.441 12.012 ;
  LAYER M1 ;
        RECT 3.519 9.576 3.521 12.012 ;
  LAYER M1 ;
        RECT 3.599 9.576 3.601 12.012 ;
  LAYER M1 ;
        RECT 3.679 9.576 3.681 12.012 ;
  LAYER M1 ;
        RECT 3.759 9.576 3.761 12.012 ;
  LAYER M1 ;
        RECT 3.839 9.576 3.841 12.012 ;
  LAYER M1 ;
        RECT 3.919 9.576 3.921 12.012 ;
  LAYER M1 ;
        RECT 3.999 9.576 4.001 12.012 ;
  LAYER M1 ;
        RECT 4.079 9.576 4.081 12.012 ;
  LAYER M1 ;
        RECT 4.159 9.576 4.161 12.012 ;
  LAYER M1 ;
        RECT 4.239 9.576 4.241 12.012 ;
  LAYER M1 ;
        RECT 4.319 9.576 4.321 12.012 ;
  LAYER M1 ;
        RECT 4.399 9.576 4.401 12.012 ;
  LAYER M1 ;
        RECT 4.479 9.576 4.481 12.012 ;
  LAYER M1 ;
        RECT 4.559 9.576 4.561 12.012 ;
  LAYER M1 ;
        RECT 4.639 9.576 4.641 12.012 ;
  LAYER M1 ;
        RECT 4.719 9.576 4.721 12.012 ;
  LAYER M1 ;
        RECT 4.799 9.576 4.801 12.012 ;
  LAYER M1 ;
        RECT 4.879 9.576 4.881 12.012 ;
  LAYER M1 ;
        RECT 4.959 9.576 4.961 12.012 ;
  LAYER M1 ;
        RECT 5.039 9.576 5.041 12.012 ;
  LAYER M1 ;
        RECT 5.119 9.576 5.121 12.012 ;
  LAYER M1 ;
        RECT 5.199 9.576 5.201 12.012 ;
  LAYER M1 ;
        RECT 5.279 9.576 5.281 12.012 ;
  LAYER M1 ;
        RECT 5.359 9.576 5.361 12.012 ;
  LAYER M1 ;
        RECT 5.439 9.576 5.441 12.012 ;
  LAYER M1 ;
        RECT 5.519 9.576 5.521 12.012 ;
  LAYER M1 ;
        RECT 5.599 9.576 5.601 12.012 ;
  LAYER M2 ;
        RECT 3.28 9.575 5.68 9.577 ;
  LAYER M2 ;
        RECT 3.28 9.659 5.68 9.661 ;
  LAYER M2 ;
        RECT 3.28 9.743 5.68 9.745 ;
  LAYER M2 ;
        RECT 3.28 9.827 5.68 9.829 ;
  LAYER M2 ;
        RECT 3.28 9.911 5.68 9.913 ;
  LAYER M2 ;
        RECT 3.28 9.995 5.68 9.997 ;
  LAYER M2 ;
        RECT 3.28 10.079 5.68 10.081 ;
  LAYER M2 ;
        RECT 3.28 10.163 5.68 10.165 ;
  LAYER M2 ;
        RECT 3.28 10.247 5.68 10.249 ;
  LAYER M2 ;
        RECT 3.28 10.331 5.68 10.333 ;
  LAYER M2 ;
        RECT 3.28 10.415 5.68 10.417 ;
  LAYER M2 ;
        RECT 3.28 10.499 5.68 10.501 ;
  LAYER M2 ;
        RECT 3.28 10.5825 5.68 10.5845 ;
  LAYER M2 ;
        RECT 3.28 10.667 5.68 10.669 ;
  LAYER M2 ;
        RECT 3.28 10.751 5.68 10.753 ;
  LAYER M2 ;
        RECT 3.28 10.835 5.68 10.837 ;
  LAYER M2 ;
        RECT 3.28 10.919 5.68 10.921 ;
  LAYER M2 ;
        RECT 3.28 11.003 5.68 11.005 ;
  LAYER M2 ;
        RECT 3.28 11.087 5.68 11.089 ;
  LAYER M2 ;
        RECT 3.28 11.171 5.68 11.173 ;
  LAYER M2 ;
        RECT 3.28 11.255 5.68 11.257 ;
  LAYER M2 ;
        RECT 3.28 11.339 5.68 11.341 ;
  LAYER M2 ;
        RECT 3.28 11.423 5.68 11.425 ;
  LAYER M2 ;
        RECT 3.28 11.507 5.68 11.509 ;
  LAYER M2 ;
        RECT 3.28 11.591 5.68 11.593 ;
  LAYER M2 ;
        RECT 3.28 11.675 5.68 11.677 ;
  LAYER M2 ;
        RECT 3.28 11.759 5.68 11.761 ;
  LAYER M2 ;
        RECT 3.28 11.843 5.68 11.845 ;
  LAYER M2 ;
        RECT 3.28 11.927 5.68 11.929 ;
  LAYER M1 ;
        RECT 3.264 12.48 3.296 14.988 ;
  LAYER M1 ;
        RECT 3.328 12.48 3.36 14.988 ;
  LAYER M1 ;
        RECT 3.392 12.48 3.424 14.988 ;
  LAYER M1 ;
        RECT 3.456 12.48 3.488 14.988 ;
  LAYER M1 ;
        RECT 3.52 12.48 3.552 14.988 ;
  LAYER M1 ;
        RECT 3.584 12.48 3.616 14.988 ;
  LAYER M1 ;
        RECT 3.648 12.48 3.68 14.988 ;
  LAYER M1 ;
        RECT 3.712 12.48 3.744 14.988 ;
  LAYER M1 ;
        RECT 3.776 12.48 3.808 14.988 ;
  LAYER M1 ;
        RECT 3.84 12.48 3.872 14.988 ;
  LAYER M1 ;
        RECT 3.904 12.48 3.936 14.988 ;
  LAYER M1 ;
        RECT 3.968 12.48 4 14.988 ;
  LAYER M1 ;
        RECT 4.032 12.48 4.064 14.988 ;
  LAYER M1 ;
        RECT 4.096 12.48 4.128 14.988 ;
  LAYER M1 ;
        RECT 4.16 12.48 4.192 14.988 ;
  LAYER M1 ;
        RECT 4.224 12.48 4.256 14.988 ;
  LAYER M1 ;
        RECT 4.288 12.48 4.32 14.988 ;
  LAYER M1 ;
        RECT 4.352 12.48 4.384 14.988 ;
  LAYER M1 ;
        RECT 4.416 12.48 4.448 14.988 ;
  LAYER M1 ;
        RECT 4.48 12.48 4.512 14.988 ;
  LAYER M1 ;
        RECT 4.544 12.48 4.576 14.988 ;
  LAYER M1 ;
        RECT 4.608 12.48 4.64 14.988 ;
  LAYER M1 ;
        RECT 4.672 12.48 4.704 14.988 ;
  LAYER M1 ;
        RECT 4.736 12.48 4.768 14.988 ;
  LAYER M1 ;
        RECT 4.8 12.48 4.832 14.988 ;
  LAYER M1 ;
        RECT 4.864 12.48 4.896 14.988 ;
  LAYER M1 ;
        RECT 4.928 12.48 4.96 14.988 ;
  LAYER M1 ;
        RECT 4.992 12.48 5.024 14.988 ;
  LAYER M1 ;
        RECT 5.056 12.48 5.088 14.988 ;
  LAYER M1 ;
        RECT 5.12 12.48 5.152 14.988 ;
  LAYER M1 ;
        RECT 5.184 12.48 5.216 14.988 ;
  LAYER M1 ;
        RECT 5.248 12.48 5.28 14.988 ;
  LAYER M1 ;
        RECT 5.312 12.48 5.344 14.988 ;
  LAYER M1 ;
        RECT 5.376 12.48 5.408 14.988 ;
  LAYER M1 ;
        RECT 5.44 12.48 5.472 14.988 ;
  LAYER M1 ;
        RECT 5.504 12.48 5.536 14.988 ;
  LAYER M1 ;
        RECT 5.568 12.48 5.6 14.988 ;
  LAYER M2 ;
        RECT 3.244 12.564 5.716 12.596 ;
  LAYER M2 ;
        RECT 3.244 12.628 5.716 12.66 ;
  LAYER M2 ;
        RECT 3.244 12.692 5.716 12.724 ;
  LAYER M2 ;
        RECT 3.244 12.756 5.716 12.788 ;
  LAYER M2 ;
        RECT 3.244 12.82 5.716 12.852 ;
  LAYER M2 ;
        RECT 3.244 12.884 5.716 12.916 ;
  LAYER M2 ;
        RECT 3.244 12.948 5.716 12.98 ;
  LAYER M2 ;
        RECT 3.244 13.012 5.716 13.044 ;
  LAYER M2 ;
        RECT 3.244 13.076 5.716 13.108 ;
  LAYER M2 ;
        RECT 3.244 13.14 5.716 13.172 ;
  LAYER M2 ;
        RECT 3.244 13.204 5.716 13.236 ;
  LAYER M2 ;
        RECT 3.244 13.268 5.716 13.3 ;
  LAYER M2 ;
        RECT 3.244 13.332 5.716 13.364 ;
  LAYER M2 ;
        RECT 3.244 13.396 5.716 13.428 ;
  LAYER M2 ;
        RECT 3.244 13.46 5.716 13.492 ;
  LAYER M2 ;
        RECT 3.244 13.524 5.716 13.556 ;
  LAYER M2 ;
        RECT 3.244 13.588 5.716 13.62 ;
  LAYER M2 ;
        RECT 3.244 13.652 5.716 13.684 ;
  LAYER M2 ;
        RECT 3.244 13.716 5.716 13.748 ;
  LAYER M2 ;
        RECT 3.244 13.78 5.716 13.812 ;
  LAYER M2 ;
        RECT 3.244 13.844 5.716 13.876 ;
  LAYER M2 ;
        RECT 3.244 13.908 5.716 13.94 ;
  LAYER M2 ;
        RECT 3.244 13.972 5.716 14.004 ;
  LAYER M2 ;
        RECT 3.244 14.036 5.716 14.068 ;
  LAYER M2 ;
        RECT 3.244 14.1 5.716 14.132 ;
  LAYER M2 ;
        RECT 3.244 14.164 5.716 14.196 ;
  LAYER M2 ;
        RECT 3.244 14.228 5.716 14.26 ;
  LAYER M2 ;
        RECT 3.244 14.292 5.716 14.324 ;
  LAYER M2 ;
        RECT 3.244 14.356 5.716 14.388 ;
  LAYER M2 ;
        RECT 3.244 14.42 5.716 14.452 ;
  LAYER M2 ;
        RECT 3.244 14.484 5.716 14.516 ;
  LAYER M2 ;
        RECT 3.244 14.548 5.716 14.58 ;
  LAYER M2 ;
        RECT 3.244 14.612 5.716 14.644 ;
  LAYER M2 ;
        RECT 3.244 14.676 5.716 14.708 ;
  LAYER M2 ;
        RECT 3.244 14.74 5.716 14.772 ;
  LAYER M2 ;
        RECT 3.244 14.804 5.716 14.836 ;
  LAYER M3 ;
        RECT 3.264 12.48 3.296 14.988 ;
  LAYER M3 ;
        RECT 3.328 12.48 3.36 14.988 ;
  LAYER M3 ;
        RECT 3.392 12.48 3.424 14.988 ;
  LAYER M3 ;
        RECT 3.456 12.48 3.488 14.988 ;
  LAYER M3 ;
        RECT 3.52 12.48 3.552 14.988 ;
  LAYER M3 ;
        RECT 3.584 12.48 3.616 14.988 ;
  LAYER M3 ;
        RECT 3.648 12.48 3.68 14.988 ;
  LAYER M3 ;
        RECT 3.712 12.48 3.744 14.988 ;
  LAYER M3 ;
        RECT 3.776 12.48 3.808 14.988 ;
  LAYER M3 ;
        RECT 3.84 12.48 3.872 14.988 ;
  LAYER M3 ;
        RECT 3.904 12.48 3.936 14.988 ;
  LAYER M3 ;
        RECT 3.968 12.48 4 14.988 ;
  LAYER M3 ;
        RECT 4.032 12.48 4.064 14.988 ;
  LAYER M3 ;
        RECT 4.096 12.48 4.128 14.988 ;
  LAYER M3 ;
        RECT 4.16 12.48 4.192 14.988 ;
  LAYER M3 ;
        RECT 4.224 12.48 4.256 14.988 ;
  LAYER M3 ;
        RECT 4.288 12.48 4.32 14.988 ;
  LAYER M3 ;
        RECT 4.352 12.48 4.384 14.988 ;
  LAYER M3 ;
        RECT 4.416 12.48 4.448 14.988 ;
  LAYER M3 ;
        RECT 4.48 12.48 4.512 14.988 ;
  LAYER M3 ;
        RECT 4.544 12.48 4.576 14.988 ;
  LAYER M3 ;
        RECT 4.608 12.48 4.64 14.988 ;
  LAYER M3 ;
        RECT 4.672 12.48 4.704 14.988 ;
  LAYER M3 ;
        RECT 4.736 12.48 4.768 14.988 ;
  LAYER M3 ;
        RECT 4.8 12.48 4.832 14.988 ;
  LAYER M3 ;
        RECT 4.864 12.48 4.896 14.988 ;
  LAYER M3 ;
        RECT 4.928 12.48 4.96 14.988 ;
  LAYER M3 ;
        RECT 4.992 12.48 5.024 14.988 ;
  LAYER M3 ;
        RECT 5.056 12.48 5.088 14.988 ;
  LAYER M3 ;
        RECT 5.12 12.48 5.152 14.988 ;
  LAYER M3 ;
        RECT 5.184 12.48 5.216 14.988 ;
  LAYER M3 ;
        RECT 5.248 12.48 5.28 14.988 ;
  LAYER M3 ;
        RECT 5.312 12.48 5.344 14.988 ;
  LAYER M3 ;
        RECT 5.376 12.48 5.408 14.988 ;
  LAYER M3 ;
        RECT 5.44 12.48 5.472 14.988 ;
  LAYER M3 ;
        RECT 5.504 12.48 5.536 14.988 ;
  LAYER M3 ;
        RECT 5.568 12.48 5.6 14.988 ;
  LAYER M3 ;
        RECT 5.664 12.48 5.696 14.988 ;
  LAYER M1 ;
        RECT 3.279 12.516 3.281 14.952 ;
  LAYER M1 ;
        RECT 3.359 12.516 3.361 14.952 ;
  LAYER M1 ;
        RECT 3.439 12.516 3.441 14.952 ;
  LAYER M1 ;
        RECT 3.519 12.516 3.521 14.952 ;
  LAYER M1 ;
        RECT 3.599 12.516 3.601 14.952 ;
  LAYER M1 ;
        RECT 3.679 12.516 3.681 14.952 ;
  LAYER M1 ;
        RECT 3.759 12.516 3.761 14.952 ;
  LAYER M1 ;
        RECT 3.839 12.516 3.841 14.952 ;
  LAYER M1 ;
        RECT 3.919 12.516 3.921 14.952 ;
  LAYER M1 ;
        RECT 3.999 12.516 4.001 14.952 ;
  LAYER M1 ;
        RECT 4.079 12.516 4.081 14.952 ;
  LAYER M1 ;
        RECT 4.159 12.516 4.161 14.952 ;
  LAYER M1 ;
        RECT 4.239 12.516 4.241 14.952 ;
  LAYER M1 ;
        RECT 4.319 12.516 4.321 14.952 ;
  LAYER M1 ;
        RECT 4.399 12.516 4.401 14.952 ;
  LAYER M1 ;
        RECT 4.479 12.516 4.481 14.952 ;
  LAYER M1 ;
        RECT 4.559 12.516 4.561 14.952 ;
  LAYER M1 ;
        RECT 4.639 12.516 4.641 14.952 ;
  LAYER M1 ;
        RECT 4.719 12.516 4.721 14.952 ;
  LAYER M1 ;
        RECT 4.799 12.516 4.801 14.952 ;
  LAYER M1 ;
        RECT 4.879 12.516 4.881 14.952 ;
  LAYER M1 ;
        RECT 4.959 12.516 4.961 14.952 ;
  LAYER M1 ;
        RECT 5.039 12.516 5.041 14.952 ;
  LAYER M1 ;
        RECT 5.119 12.516 5.121 14.952 ;
  LAYER M1 ;
        RECT 5.199 12.516 5.201 14.952 ;
  LAYER M1 ;
        RECT 5.279 12.516 5.281 14.952 ;
  LAYER M1 ;
        RECT 5.359 12.516 5.361 14.952 ;
  LAYER M1 ;
        RECT 5.439 12.516 5.441 14.952 ;
  LAYER M1 ;
        RECT 5.519 12.516 5.521 14.952 ;
  LAYER M1 ;
        RECT 5.599 12.516 5.601 14.952 ;
  LAYER M2 ;
        RECT 3.28 12.515 5.68 12.517 ;
  LAYER M2 ;
        RECT 3.28 12.599 5.68 12.601 ;
  LAYER M2 ;
        RECT 3.28 12.683 5.68 12.685 ;
  LAYER M2 ;
        RECT 3.28 12.767 5.68 12.769 ;
  LAYER M2 ;
        RECT 3.28 12.851 5.68 12.853 ;
  LAYER M2 ;
        RECT 3.28 12.935 5.68 12.937 ;
  LAYER M2 ;
        RECT 3.28 13.019 5.68 13.021 ;
  LAYER M2 ;
        RECT 3.28 13.103 5.68 13.105 ;
  LAYER M2 ;
        RECT 3.28 13.187 5.68 13.189 ;
  LAYER M2 ;
        RECT 3.28 13.271 5.68 13.273 ;
  LAYER M2 ;
        RECT 3.28 13.355 5.68 13.357 ;
  LAYER M2 ;
        RECT 3.28 13.439 5.68 13.441 ;
  LAYER M2 ;
        RECT 3.28 13.5225 5.68 13.5245 ;
  LAYER M2 ;
        RECT 3.28 13.607 5.68 13.609 ;
  LAYER M2 ;
        RECT 3.28 13.691 5.68 13.693 ;
  LAYER M2 ;
        RECT 3.28 13.775 5.68 13.777 ;
  LAYER M2 ;
        RECT 3.28 13.859 5.68 13.861 ;
  LAYER M2 ;
        RECT 3.28 13.943 5.68 13.945 ;
  LAYER M2 ;
        RECT 3.28 14.027 5.68 14.029 ;
  LAYER M2 ;
        RECT 3.28 14.111 5.68 14.113 ;
  LAYER M2 ;
        RECT 3.28 14.195 5.68 14.197 ;
  LAYER M2 ;
        RECT 3.28 14.279 5.68 14.281 ;
  LAYER M2 ;
        RECT 3.28 14.363 5.68 14.365 ;
  LAYER M2 ;
        RECT 3.28 14.447 5.68 14.449 ;
  LAYER M2 ;
        RECT 3.28 14.531 5.68 14.533 ;
  LAYER M2 ;
        RECT 3.28 14.615 5.68 14.617 ;
  LAYER M2 ;
        RECT 3.28 14.699 5.68 14.701 ;
  LAYER M2 ;
        RECT 3.28 14.783 5.68 14.785 ;
  LAYER M2 ;
        RECT 3.28 14.867 5.68 14.869 ;
  LAYER M1 ;
        RECT 3.264 15.42 3.296 17.928 ;
  LAYER M1 ;
        RECT 3.328 15.42 3.36 17.928 ;
  LAYER M1 ;
        RECT 3.392 15.42 3.424 17.928 ;
  LAYER M1 ;
        RECT 3.456 15.42 3.488 17.928 ;
  LAYER M1 ;
        RECT 3.52 15.42 3.552 17.928 ;
  LAYER M1 ;
        RECT 3.584 15.42 3.616 17.928 ;
  LAYER M1 ;
        RECT 3.648 15.42 3.68 17.928 ;
  LAYER M1 ;
        RECT 3.712 15.42 3.744 17.928 ;
  LAYER M1 ;
        RECT 3.776 15.42 3.808 17.928 ;
  LAYER M1 ;
        RECT 3.84 15.42 3.872 17.928 ;
  LAYER M1 ;
        RECT 3.904 15.42 3.936 17.928 ;
  LAYER M1 ;
        RECT 3.968 15.42 4 17.928 ;
  LAYER M1 ;
        RECT 4.032 15.42 4.064 17.928 ;
  LAYER M1 ;
        RECT 4.096 15.42 4.128 17.928 ;
  LAYER M1 ;
        RECT 4.16 15.42 4.192 17.928 ;
  LAYER M1 ;
        RECT 4.224 15.42 4.256 17.928 ;
  LAYER M1 ;
        RECT 4.288 15.42 4.32 17.928 ;
  LAYER M1 ;
        RECT 4.352 15.42 4.384 17.928 ;
  LAYER M1 ;
        RECT 4.416 15.42 4.448 17.928 ;
  LAYER M1 ;
        RECT 4.48 15.42 4.512 17.928 ;
  LAYER M1 ;
        RECT 4.544 15.42 4.576 17.928 ;
  LAYER M1 ;
        RECT 4.608 15.42 4.64 17.928 ;
  LAYER M1 ;
        RECT 4.672 15.42 4.704 17.928 ;
  LAYER M1 ;
        RECT 4.736 15.42 4.768 17.928 ;
  LAYER M1 ;
        RECT 4.8 15.42 4.832 17.928 ;
  LAYER M1 ;
        RECT 4.864 15.42 4.896 17.928 ;
  LAYER M1 ;
        RECT 4.928 15.42 4.96 17.928 ;
  LAYER M1 ;
        RECT 4.992 15.42 5.024 17.928 ;
  LAYER M1 ;
        RECT 5.056 15.42 5.088 17.928 ;
  LAYER M1 ;
        RECT 5.12 15.42 5.152 17.928 ;
  LAYER M1 ;
        RECT 5.184 15.42 5.216 17.928 ;
  LAYER M1 ;
        RECT 5.248 15.42 5.28 17.928 ;
  LAYER M1 ;
        RECT 5.312 15.42 5.344 17.928 ;
  LAYER M1 ;
        RECT 5.376 15.42 5.408 17.928 ;
  LAYER M1 ;
        RECT 5.44 15.42 5.472 17.928 ;
  LAYER M1 ;
        RECT 5.504 15.42 5.536 17.928 ;
  LAYER M1 ;
        RECT 5.568 15.42 5.6 17.928 ;
  LAYER M2 ;
        RECT 3.244 15.504 5.716 15.536 ;
  LAYER M2 ;
        RECT 3.244 15.568 5.716 15.6 ;
  LAYER M2 ;
        RECT 3.244 15.632 5.716 15.664 ;
  LAYER M2 ;
        RECT 3.244 15.696 5.716 15.728 ;
  LAYER M2 ;
        RECT 3.244 15.76 5.716 15.792 ;
  LAYER M2 ;
        RECT 3.244 15.824 5.716 15.856 ;
  LAYER M2 ;
        RECT 3.244 15.888 5.716 15.92 ;
  LAYER M2 ;
        RECT 3.244 15.952 5.716 15.984 ;
  LAYER M2 ;
        RECT 3.244 16.016 5.716 16.048 ;
  LAYER M2 ;
        RECT 3.244 16.08 5.716 16.112 ;
  LAYER M2 ;
        RECT 3.244 16.144 5.716 16.176 ;
  LAYER M2 ;
        RECT 3.244 16.208 5.716 16.24 ;
  LAYER M2 ;
        RECT 3.244 16.272 5.716 16.304 ;
  LAYER M2 ;
        RECT 3.244 16.336 5.716 16.368 ;
  LAYER M2 ;
        RECT 3.244 16.4 5.716 16.432 ;
  LAYER M2 ;
        RECT 3.244 16.464 5.716 16.496 ;
  LAYER M2 ;
        RECT 3.244 16.528 5.716 16.56 ;
  LAYER M2 ;
        RECT 3.244 16.592 5.716 16.624 ;
  LAYER M2 ;
        RECT 3.244 16.656 5.716 16.688 ;
  LAYER M2 ;
        RECT 3.244 16.72 5.716 16.752 ;
  LAYER M2 ;
        RECT 3.244 16.784 5.716 16.816 ;
  LAYER M2 ;
        RECT 3.244 16.848 5.716 16.88 ;
  LAYER M2 ;
        RECT 3.244 16.912 5.716 16.944 ;
  LAYER M2 ;
        RECT 3.244 16.976 5.716 17.008 ;
  LAYER M2 ;
        RECT 3.244 17.04 5.716 17.072 ;
  LAYER M2 ;
        RECT 3.244 17.104 5.716 17.136 ;
  LAYER M2 ;
        RECT 3.244 17.168 5.716 17.2 ;
  LAYER M2 ;
        RECT 3.244 17.232 5.716 17.264 ;
  LAYER M2 ;
        RECT 3.244 17.296 5.716 17.328 ;
  LAYER M2 ;
        RECT 3.244 17.36 5.716 17.392 ;
  LAYER M2 ;
        RECT 3.244 17.424 5.716 17.456 ;
  LAYER M2 ;
        RECT 3.244 17.488 5.716 17.52 ;
  LAYER M2 ;
        RECT 3.244 17.552 5.716 17.584 ;
  LAYER M2 ;
        RECT 3.244 17.616 5.716 17.648 ;
  LAYER M2 ;
        RECT 3.244 17.68 5.716 17.712 ;
  LAYER M2 ;
        RECT 3.244 17.744 5.716 17.776 ;
  LAYER M3 ;
        RECT 3.264 15.42 3.296 17.928 ;
  LAYER M3 ;
        RECT 3.328 15.42 3.36 17.928 ;
  LAYER M3 ;
        RECT 3.392 15.42 3.424 17.928 ;
  LAYER M3 ;
        RECT 3.456 15.42 3.488 17.928 ;
  LAYER M3 ;
        RECT 3.52 15.42 3.552 17.928 ;
  LAYER M3 ;
        RECT 3.584 15.42 3.616 17.928 ;
  LAYER M3 ;
        RECT 3.648 15.42 3.68 17.928 ;
  LAYER M3 ;
        RECT 3.712 15.42 3.744 17.928 ;
  LAYER M3 ;
        RECT 3.776 15.42 3.808 17.928 ;
  LAYER M3 ;
        RECT 3.84 15.42 3.872 17.928 ;
  LAYER M3 ;
        RECT 3.904 15.42 3.936 17.928 ;
  LAYER M3 ;
        RECT 3.968 15.42 4 17.928 ;
  LAYER M3 ;
        RECT 4.032 15.42 4.064 17.928 ;
  LAYER M3 ;
        RECT 4.096 15.42 4.128 17.928 ;
  LAYER M3 ;
        RECT 4.16 15.42 4.192 17.928 ;
  LAYER M3 ;
        RECT 4.224 15.42 4.256 17.928 ;
  LAYER M3 ;
        RECT 4.288 15.42 4.32 17.928 ;
  LAYER M3 ;
        RECT 4.352 15.42 4.384 17.928 ;
  LAYER M3 ;
        RECT 4.416 15.42 4.448 17.928 ;
  LAYER M3 ;
        RECT 4.48 15.42 4.512 17.928 ;
  LAYER M3 ;
        RECT 4.544 15.42 4.576 17.928 ;
  LAYER M3 ;
        RECT 4.608 15.42 4.64 17.928 ;
  LAYER M3 ;
        RECT 4.672 15.42 4.704 17.928 ;
  LAYER M3 ;
        RECT 4.736 15.42 4.768 17.928 ;
  LAYER M3 ;
        RECT 4.8 15.42 4.832 17.928 ;
  LAYER M3 ;
        RECT 4.864 15.42 4.896 17.928 ;
  LAYER M3 ;
        RECT 4.928 15.42 4.96 17.928 ;
  LAYER M3 ;
        RECT 4.992 15.42 5.024 17.928 ;
  LAYER M3 ;
        RECT 5.056 15.42 5.088 17.928 ;
  LAYER M3 ;
        RECT 5.12 15.42 5.152 17.928 ;
  LAYER M3 ;
        RECT 5.184 15.42 5.216 17.928 ;
  LAYER M3 ;
        RECT 5.248 15.42 5.28 17.928 ;
  LAYER M3 ;
        RECT 5.312 15.42 5.344 17.928 ;
  LAYER M3 ;
        RECT 5.376 15.42 5.408 17.928 ;
  LAYER M3 ;
        RECT 5.44 15.42 5.472 17.928 ;
  LAYER M3 ;
        RECT 5.504 15.42 5.536 17.928 ;
  LAYER M3 ;
        RECT 5.568 15.42 5.6 17.928 ;
  LAYER M3 ;
        RECT 5.664 15.42 5.696 17.928 ;
  LAYER M1 ;
        RECT 3.279 15.456 3.281 17.892 ;
  LAYER M1 ;
        RECT 3.359 15.456 3.361 17.892 ;
  LAYER M1 ;
        RECT 3.439 15.456 3.441 17.892 ;
  LAYER M1 ;
        RECT 3.519 15.456 3.521 17.892 ;
  LAYER M1 ;
        RECT 3.599 15.456 3.601 17.892 ;
  LAYER M1 ;
        RECT 3.679 15.456 3.681 17.892 ;
  LAYER M1 ;
        RECT 3.759 15.456 3.761 17.892 ;
  LAYER M1 ;
        RECT 3.839 15.456 3.841 17.892 ;
  LAYER M1 ;
        RECT 3.919 15.456 3.921 17.892 ;
  LAYER M1 ;
        RECT 3.999 15.456 4.001 17.892 ;
  LAYER M1 ;
        RECT 4.079 15.456 4.081 17.892 ;
  LAYER M1 ;
        RECT 4.159 15.456 4.161 17.892 ;
  LAYER M1 ;
        RECT 4.239 15.456 4.241 17.892 ;
  LAYER M1 ;
        RECT 4.319 15.456 4.321 17.892 ;
  LAYER M1 ;
        RECT 4.399 15.456 4.401 17.892 ;
  LAYER M1 ;
        RECT 4.479 15.456 4.481 17.892 ;
  LAYER M1 ;
        RECT 4.559 15.456 4.561 17.892 ;
  LAYER M1 ;
        RECT 4.639 15.456 4.641 17.892 ;
  LAYER M1 ;
        RECT 4.719 15.456 4.721 17.892 ;
  LAYER M1 ;
        RECT 4.799 15.456 4.801 17.892 ;
  LAYER M1 ;
        RECT 4.879 15.456 4.881 17.892 ;
  LAYER M1 ;
        RECT 4.959 15.456 4.961 17.892 ;
  LAYER M1 ;
        RECT 5.039 15.456 5.041 17.892 ;
  LAYER M1 ;
        RECT 5.119 15.456 5.121 17.892 ;
  LAYER M1 ;
        RECT 5.199 15.456 5.201 17.892 ;
  LAYER M1 ;
        RECT 5.279 15.456 5.281 17.892 ;
  LAYER M1 ;
        RECT 5.359 15.456 5.361 17.892 ;
  LAYER M1 ;
        RECT 5.439 15.456 5.441 17.892 ;
  LAYER M1 ;
        RECT 5.519 15.456 5.521 17.892 ;
  LAYER M1 ;
        RECT 5.599 15.456 5.601 17.892 ;
  LAYER M2 ;
        RECT 3.28 15.455 5.68 15.457 ;
  LAYER M2 ;
        RECT 3.28 15.539 5.68 15.541 ;
  LAYER M2 ;
        RECT 3.28 15.623 5.68 15.625 ;
  LAYER M2 ;
        RECT 3.28 15.707 5.68 15.709 ;
  LAYER M2 ;
        RECT 3.28 15.791 5.68 15.793 ;
  LAYER M2 ;
        RECT 3.28 15.875 5.68 15.877 ;
  LAYER M2 ;
        RECT 3.28 15.959 5.68 15.961 ;
  LAYER M2 ;
        RECT 3.28 16.043 5.68 16.045 ;
  LAYER M2 ;
        RECT 3.28 16.127 5.68 16.129 ;
  LAYER M2 ;
        RECT 3.28 16.211 5.68 16.213 ;
  LAYER M2 ;
        RECT 3.28 16.295 5.68 16.297 ;
  LAYER M2 ;
        RECT 3.28 16.379 5.68 16.381 ;
  LAYER M2 ;
        RECT 3.28 16.4625 5.68 16.4645 ;
  LAYER M2 ;
        RECT 3.28 16.547 5.68 16.549 ;
  LAYER M2 ;
        RECT 3.28 16.631 5.68 16.633 ;
  LAYER M2 ;
        RECT 3.28 16.715 5.68 16.717 ;
  LAYER M2 ;
        RECT 3.28 16.799 5.68 16.801 ;
  LAYER M2 ;
        RECT 3.28 16.883 5.68 16.885 ;
  LAYER M2 ;
        RECT 3.28 16.967 5.68 16.969 ;
  LAYER M2 ;
        RECT 3.28 17.051 5.68 17.053 ;
  LAYER M2 ;
        RECT 3.28 17.135 5.68 17.137 ;
  LAYER M2 ;
        RECT 3.28 17.219 5.68 17.221 ;
  LAYER M2 ;
        RECT 3.28 17.303 5.68 17.305 ;
  LAYER M2 ;
        RECT 3.28 17.387 5.68 17.389 ;
  LAYER M2 ;
        RECT 3.28 17.471 5.68 17.473 ;
  LAYER M2 ;
        RECT 3.28 17.555 5.68 17.557 ;
  LAYER M2 ;
        RECT 3.28 17.639 5.68 17.641 ;
  LAYER M2 ;
        RECT 3.28 17.723 5.68 17.725 ;
  LAYER M2 ;
        RECT 3.28 17.807 5.68 17.809 ;
  LAYER M1 ;
        RECT 3.264 18.36 3.296 20.868 ;
  LAYER M1 ;
        RECT 3.328 18.36 3.36 20.868 ;
  LAYER M1 ;
        RECT 3.392 18.36 3.424 20.868 ;
  LAYER M1 ;
        RECT 3.456 18.36 3.488 20.868 ;
  LAYER M1 ;
        RECT 3.52 18.36 3.552 20.868 ;
  LAYER M1 ;
        RECT 3.584 18.36 3.616 20.868 ;
  LAYER M1 ;
        RECT 3.648 18.36 3.68 20.868 ;
  LAYER M1 ;
        RECT 3.712 18.36 3.744 20.868 ;
  LAYER M1 ;
        RECT 3.776 18.36 3.808 20.868 ;
  LAYER M1 ;
        RECT 3.84 18.36 3.872 20.868 ;
  LAYER M1 ;
        RECT 3.904 18.36 3.936 20.868 ;
  LAYER M1 ;
        RECT 3.968 18.36 4 20.868 ;
  LAYER M1 ;
        RECT 4.032 18.36 4.064 20.868 ;
  LAYER M1 ;
        RECT 4.096 18.36 4.128 20.868 ;
  LAYER M1 ;
        RECT 4.16 18.36 4.192 20.868 ;
  LAYER M1 ;
        RECT 4.224 18.36 4.256 20.868 ;
  LAYER M1 ;
        RECT 4.288 18.36 4.32 20.868 ;
  LAYER M1 ;
        RECT 4.352 18.36 4.384 20.868 ;
  LAYER M1 ;
        RECT 4.416 18.36 4.448 20.868 ;
  LAYER M1 ;
        RECT 4.48 18.36 4.512 20.868 ;
  LAYER M1 ;
        RECT 4.544 18.36 4.576 20.868 ;
  LAYER M1 ;
        RECT 4.608 18.36 4.64 20.868 ;
  LAYER M1 ;
        RECT 4.672 18.36 4.704 20.868 ;
  LAYER M1 ;
        RECT 4.736 18.36 4.768 20.868 ;
  LAYER M1 ;
        RECT 4.8 18.36 4.832 20.868 ;
  LAYER M1 ;
        RECT 4.864 18.36 4.896 20.868 ;
  LAYER M1 ;
        RECT 4.928 18.36 4.96 20.868 ;
  LAYER M1 ;
        RECT 4.992 18.36 5.024 20.868 ;
  LAYER M1 ;
        RECT 5.056 18.36 5.088 20.868 ;
  LAYER M1 ;
        RECT 5.12 18.36 5.152 20.868 ;
  LAYER M1 ;
        RECT 5.184 18.36 5.216 20.868 ;
  LAYER M1 ;
        RECT 5.248 18.36 5.28 20.868 ;
  LAYER M1 ;
        RECT 5.312 18.36 5.344 20.868 ;
  LAYER M1 ;
        RECT 5.376 18.36 5.408 20.868 ;
  LAYER M1 ;
        RECT 5.44 18.36 5.472 20.868 ;
  LAYER M1 ;
        RECT 5.504 18.36 5.536 20.868 ;
  LAYER M1 ;
        RECT 5.568 18.36 5.6 20.868 ;
  LAYER M2 ;
        RECT 3.244 18.444 5.716 18.476 ;
  LAYER M2 ;
        RECT 3.244 18.508 5.716 18.54 ;
  LAYER M2 ;
        RECT 3.244 18.572 5.716 18.604 ;
  LAYER M2 ;
        RECT 3.244 18.636 5.716 18.668 ;
  LAYER M2 ;
        RECT 3.244 18.7 5.716 18.732 ;
  LAYER M2 ;
        RECT 3.244 18.764 5.716 18.796 ;
  LAYER M2 ;
        RECT 3.244 18.828 5.716 18.86 ;
  LAYER M2 ;
        RECT 3.244 18.892 5.716 18.924 ;
  LAYER M2 ;
        RECT 3.244 18.956 5.716 18.988 ;
  LAYER M2 ;
        RECT 3.244 19.02 5.716 19.052 ;
  LAYER M2 ;
        RECT 3.244 19.084 5.716 19.116 ;
  LAYER M2 ;
        RECT 3.244 19.148 5.716 19.18 ;
  LAYER M2 ;
        RECT 3.244 19.212 5.716 19.244 ;
  LAYER M2 ;
        RECT 3.244 19.276 5.716 19.308 ;
  LAYER M2 ;
        RECT 3.244 19.34 5.716 19.372 ;
  LAYER M2 ;
        RECT 3.244 19.404 5.716 19.436 ;
  LAYER M2 ;
        RECT 3.244 19.468 5.716 19.5 ;
  LAYER M2 ;
        RECT 3.244 19.532 5.716 19.564 ;
  LAYER M2 ;
        RECT 3.244 19.596 5.716 19.628 ;
  LAYER M2 ;
        RECT 3.244 19.66 5.716 19.692 ;
  LAYER M2 ;
        RECT 3.244 19.724 5.716 19.756 ;
  LAYER M2 ;
        RECT 3.244 19.788 5.716 19.82 ;
  LAYER M2 ;
        RECT 3.244 19.852 5.716 19.884 ;
  LAYER M2 ;
        RECT 3.244 19.916 5.716 19.948 ;
  LAYER M2 ;
        RECT 3.244 19.98 5.716 20.012 ;
  LAYER M2 ;
        RECT 3.244 20.044 5.716 20.076 ;
  LAYER M2 ;
        RECT 3.244 20.108 5.716 20.14 ;
  LAYER M2 ;
        RECT 3.244 20.172 5.716 20.204 ;
  LAYER M2 ;
        RECT 3.244 20.236 5.716 20.268 ;
  LAYER M2 ;
        RECT 3.244 20.3 5.716 20.332 ;
  LAYER M2 ;
        RECT 3.244 20.364 5.716 20.396 ;
  LAYER M2 ;
        RECT 3.244 20.428 5.716 20.46 ;
  LAYER M2 ;
        RECT 3.244 20.492 5.716 20.524 ;
  LAYER M2 ;
        RECT 3.244 20.556 5.716 20.588 ;
  LAYER M2 ;
        RECT 3.244 20.62 5.716 20.652 ;
  LAYER M2 ;
        RECT 3.244 20.684 5.716 20.716 ;
  LAYER M3 ;
        RECT 3.264 18.36 3.296 20.868 ;
  LAYER M3 ;
        RECT 3.328 18.36 3.36 20.868 ;
  LAYER M3 ;
        RECT 3.392 18.36 3.424 20.868 ;
  LAYER M3 ;
        RECT 3.456 18.36 3.488 20.868 ;
  LAYER M3 ;
        RECT 3.52 18.36 3.552 20.868 ;
  LAYER M3 ;
        RECT 3.584 18.36 3.616 20.868 ;
  LAYER M3 ;
        RECT 3.648 18.36 3.68 20.868 ;
  LAYER M3 ;
        RECT 3.712 18.36 3.744 20.868 ;
  LAYER M3 ;
        RECT 3.776 18.36 3.808 20.868 ;
  LAYER M3 ;
        RECT 3.84 18.36 3.872 20.868 ;
  LAYER M3 ;
        RECT 3.904 18.36 3.936 20.868 ;
  LAYER M3 ;
        RECT 3.968 18.36 4 20.868 ;
  LAYER M3 ;
        RECT 4.032 18.36 4.064 20.868 ;
  LAYER M3 ;
        RECT 4.096 18.36 4.128 20.868 ;
  LAYER M3 ;
        RECT 4.16 18.36 4.192 20.868 ;
  LAYER M3 ;
        RECT 4.224 18.36 4.256 20.868 ;
  LAYER M3 ;
        RECT 4.288 18.36 4.32 20.868 ;
  LAYER M3 ;
        RECT 4.352 18.36 4.384 20.868 ;
  LAYER M3 ;
        RECT 4.416 18.36 4.448 20.868 ;
  LAYER M3 ;
        RECT 4.48 18.36 4.512 20.868 ;
  LAYER M3 ;
        RECT 4.544 18.36 4.576 20.868 ;
  LAYER M3 ;
        RECT 4.608 18.36 4.64 20.868 ;
  LAYER M3 ;
        RECT 4.672 18.36 4.704 20.868 ;
  LAYER M3 ;
        RECT 4.736 18.36 4.768 20.868 ;
  LAYER M3 ;
        RECT 4.8 18.36 4.832 20.868 ;
  LAYER M3 ;
        RECT 4.864 18.36 4.896 20.868 ;
  LAYER M3 ;
        RECT 4.928 18.36 4.96 20.868 ;
  LAYER M3 ;
        RECT 4.992 18.36 5.024 20.868 ;
  LAYER M3 ;
        RECT 5.056 18.36 5.088 20.868 ;
  LAYER M3 ;
        RECT 5.12 18.36 5.152 20.868 ;
  LAYER M3 ;
        RECT 5.184 18.36 5.216 20.868 ;
  LAYER M3 ;
        RECT 5.248 18.36 5.28 20.868 ;
  LAYER M3 ;
        RECT 5.312 18.36 5.344 20.868 ;
  LAYER M3 ;
        RECT 5.376 18.36 5.408 20.868 ;
  LAYER M3 ;
        RECT 5.44 18.36 5.472 20.868 ;
  LAYER M3 ;
        RECT 5.504 18.36 5.536 20.868 ;
  LAYER M3 ;
        RECT 5.568 18.36 5.6 20.868 ;
  LAYER M3 ;
        RECT 5.664 18.36 5.696 20.868 ;
  LAYER M1 ;
        RECT 3.279 18.396 3.281 20.832 ;
  LAYER M1 ;
        RECT 3.359 18.396 3.361 20.832 ;
  LAYER M1 ;
        RECT 3.439 18.396 3.441 20.832 ;
  LAYER M1 ;
        RECT 3.519 18.396 3.521 20.832 ;
  LAYER M1 ;
        RECT 3.599 18.396 3.601 20.832 ;
  LAYER M1 ;
        RECT 3.679 18.396 3.681 20.832 ;
  LAYER M1 ;
        RECT 3.759 18.396 3.761 20.832 ;
  LAYER M1 ;
        RECT 3.839 18.396 3.841 20.832 ;
  LAYER M1 ;
        RECT 3.919 18.396 3.921 20.832 ;
  LAYER M1 ;
        RECT 3.999 18.396 4.001 20.832 ;
  LAYER M1 ;
        RECT 4.079 18.396 4.081 20.832 ;
  LAYER M1 ;
        RECT 4.159 18.396 4.161 20.832 ;
  LAYER M1 ;
        RECT 4.239 18.396 4.241 20.832 ;
  LAYER M1 ;
        RECT 4.319 18.396 4.321 20.832 ;
  LAYER M1 ;
        RECT 4.399 18.396 4.401 20.832 ;
  LAYER M1 ;
        RECT 4.479 18.396 4.481 20.832 ;
  LAYER M1 ;
        RECT 4.559 18.396 4.561 20.832 ;
  LAYER M1 ;
        RECT 4.639 18.396 4.641 20.832 ;
  LAYER M1 ;
        RECT 4.719 18.396 4.721 20.832 ;
  LAYER M1 ;
        RECT 4.799 18.396 4.801 20.832 ;
  LAYER M1 ;
        RECT 4.879 18.396 4.881 20.832 ;
  LAYER M1 ;
        RECT 4.959 18.396 4.961 20.832 ;
  LAYER M1 ;
        RECT 5.039 18.396 5.041 20.832 ;
  LAYER M1 ;
        RECT 5.119 18.396 5.121 20.832 ;
  LAYER M1 ;
        RECT 5.199 18.396 5.201 20.832 ;
  LAYER M1 ;
        RECT 5.279 18.396 5.281 20.832 ;
  LAYER M1 ;
        RECT 5.359 18.396 5.361 20.832 ;
  LAYER M1 ;
        RECT 5.439 18.396 5.441 20.832 ;
  LAYER M1 ;
        RECT 5.519 18.396 5.521 20.832 ;
  LAYER M1 ;
        RECT 5.599 18.396 5.601 20.832 ;
  LAYER M2 ;
        RECT 3.28 18.395 5.68 18.397 ;
  LAYER M2 ;
        RECT 3.28 18.479 5.68 18.481 ;
  LAYER M2 ;
        RECT 3.28 18.563 5.68 18.565 ;
  LAYER M2 ;
        RECT 3.28 18.647 5.68 18.649 ;
  LAYER M2 ;
        RECT 3.28 18.731 5.68 18.733 ;
  LAYER M2 ;
        RECT 3.28 18.815 5.68 18.817 ;
  LAYER M2 ;
        RECT 3.28 18.899 5.68 18.901 ;
  LAYER M2 ;
        RECT 3.28 18.983 5.68 18.985 ;
  LAYER M2 ;
        RECT 3.28 19.067 5.68 19.069 ;
  LAYER M2 ;
        RECT 3.28 19.151 5.68 19.153 ;
  LAYER M2 ;
        RECT 3.28 19.235 5.68 19.237 ;
  LAYER M2 ;
        RECT 3.28 19.319 5.68 19.321 ;
  LAYER M2 ;
        RECT 3.28 19.4025 5.68 19.4045 ;
  LAYER M2 ;
        RECT 3.28 19.487 5.68 19.489 ;
  LAYER M2 ;
        RECT 3.28 19.571 5.68 19.573 ;
  LAYER M2 ;
        RECT 3.28 19.655 5.68 19.657 ;
  LAYER M2 ;
        RECT 3.28 19.739 5.68 19.741 ;
  LAYER M2 ;
        RECT 3.28 19.823 5.68 19.825 ;
  LAYER M2 ;
        RECT 3.28 19.907 5.68 19.909 ;
  LAYER M2 ;
        RECT 3.28 19.991 5.68 19.993 ;
  LAYER M2 ;
        RECT 3.28 20.075 5.68 20.077 ;
  LAYER M2 ;
        RECT 3.28 20.159 5.68 20.161 ;
  LAYER M2 ;
        RECT 3.28 20.243 5.68 20.245 ;
  LAYER M2 ;
        RECT 3.28 20.327 5.68 20.329 ;
  LAYER M2 ;
        RECT 3.28 20.411 5.68 20.413 ;
  LAYER M2 ;
        RECT 3.28 20.495 5.68 20.497 ;
  LAYER M2 ;
        RECT 3.28 20.579 5.68 20.581 ;
  LAYER M2 ;
        RECT 3.28 20.663 5.68 20.665 ;
  LAYER M2 ;
        RECT 3.28 20.747 5.68 20.749 ;
  LAYER M1 ;
        RECT 3.264 21.3 3.296 23.808 ;
  LAYER M1 ;
        RECT 3.328 21.3 3.36 23.808 ;
  LAYER M1 ;
        RECT 3.392 21.3 3.424 23.808 ;
  LAYER M1 ;
        RECT 3.456 21.3 3.488 23.808 ;
  LAYER M1 ;
        RECT 3.52 21.3 3.552 23.808 ;
  LAYER M1 ;
        RECT 3.584 21.3 3.616 23.808 ;
  LAYER M1 ;
        RECT 3.648 21.3 3.68 23.808 ;
  LAYER M1 ;
        RECT 3.712 21.3 3.744 23.808 ;
  LAYER M1 ;
        RECT 3.776 21.3 3.808 23.808 ;
  LAYER M1 ;
        RECT 3.84 21.3 3.872 23.808 ;
  LAYER M1 ;
        RECT 3.904 21.3 3.936 23.808 ;
  LAYER M1 ;
        RECT 3.968 21.3 4 23.808 ;
  LAYER M1 ;
        RECT 4.032 21.3 4.064 23.808 ;
  LAYER M1 ;
        RECT 4.096 21.3 4.128 23.808 ;
  LAYER M1 ;
        RECT 4.16 21.3 4.192 23.808 ;
  LAYER M1 ;
        RECT 4.224 21.3 4.256 23.808 ;
  LAYER M1 ;
        RECT 4.288 21.3 4.32 23.808 ;
  LAYER M1 ;
        RECT 4.352 21.3 4.384 23.808 ;
  LAYER M1 ;
        RECT 4.416 21.3 4.448 23.808 ;
  LAYER M1 ;
        RECT 4.48 21.3 4.512 23.808 ;
  LAYER M1 ;
        RECT 4.544 21.3 4.576 23.808 ;
  LAYER M1 ;
        RECT 4.608 21.3 4.64 23.808 ;
  LAYER M1 ;
        RECT 4.672 21.3 4.704 23.808 ;
  LAYER M1 ;
        RECT 4.736 21.3 4.768 23.808 ;
  LAYER M1 ;
        RECT 4.8 21.3 4.832 23.808 ;
  LAYER M1 ;
        RECT 4.864 21.3 4.896 23.808 ;
  LAYER M1 ;
        RECT 4.928 21.3 4.96 23.808 ;
  LAYER M1 ;
        RECT 4.992 21.3 5.024 23.808 ;
  LAYER M1 ;
        RECT 5.056 21.3 5.088 23.808 ;
  LAYER M1 ;
        RECT 5.12 21.3 5.152 23.808 ;
  LAYER M1 ;
        RECT 5.184 21.3 5.216 23.808 ;
  LAYER M1 ;
        RECT 5.248 21.3 5.28 23.808 ;
  LAYER M1 ;
        RECT 5.312 21.3 5.344 23.808 ;
  LAYER M1 ;
        RECT 5.376 21.3 5.408 23.808 ;
  LAYER M1 ;
        RECT 5.44 21.3 5.472 23.808 ;
  LAYER M1 ;
        RECT 5.504 21.3 5.536 23.808 ;
  LAYER M1 ;
        RECT 5.568 21.3 5.6 23.808 ;
  LAYER M2 ;
        RECT 3.244 21.384 5.716 21.416 ;
  LAYER M2 ;
        RECT 3.244 21.448 5.716 21.48 ;
  LAYER M2 ;
        RECT 3.244 21.512 5.716 21.544 ;
  LAYER M2 ;
        RECT 3.244 21.576 5.716 21.608 ;
  LAYER M2 ;
        RECT 3.244 21.64 5.716 21.672 ;
  LAYER M2 ;
        RECT 3.244 21.704 5.716 21.736 ;
  LAYER M2 ;
        RECT 3.244 21.768 5.716 21.8 ;
  LAYER M2 ;
        RECT 3.244 21.832 5.716 21.864 ;
  LAYER M2 ;
        RECT 3.244 21.896 5.716 21.928 ;
  LAYER M2 ;
        RECT 3.244 21.96 5.716 21.992 ;
  LAYER M2 ;
        RECT 3.244 22.024 5.716 22.056 ;
  LAYER M2 ;
        RECT 3.244 22.088 5.716 22.12 ;
  LAYER M2 ;
        RECT 3.244 22.152 5.716 22.184 ;
  LAYER M2 ;
        RECT 3.244 22.216 5.716 22.248 ;
  LAYER M2 ;
        RECT 3.244 22.28 5.716 22.312 ;
  LAYER M2 ;
        RECT 3.244 22.344 5.716 22.376 ;
  LAYER M2 ;
        RECT 3.244 22.408 5.716 22.44 ;
  LAYER M2 ;
        RECT 3.244 22.472 5.716 22.504 ;
  LAYER M2 ;
        RECT 3.244 22.536 5.716 22.568 ;
  LAYER M2 ;
        RECT 3.244 22.6 5.716 22.632 ;
  LAYER M2 ;
        RECT 3.244 22.664 5.716 22.696 ;
  LAYER M2 ;
        RECT 3.244 22.728 5.716 22.76 ;
  LAYER M2 ;
        RECT 3.244 22.792 5.716 22.824 ;
  LAYER M2 ;
        RECT 3.244 22.856 5.716 22.888 ;
  LAYER M2 ;
        RECT 3.244 22.92 5.716 22.952 ;
  LAYER M2 ;
        RECT 3.244 22.984 5.716 23.016 ;
  LAYER M2 ;
        RECT 3.244 23.048 5.716 23.08 ;
  LAYER M2 ;
        RECT 3.244 23.112 5.716 23.144 ;
  LAYER M2 ;
        RECT 3.244 23.176 5.716 23.208 ;
  LAYER M2 ;
        RECT 3.244 23.24 5.716 23.272 ;
  LAYER M2 ;
        RECT 3.244 23.304 5.716 23.336 ;
  LAYER M2 ;
        RECT 3.244 23.368 5.716 23.4 ;
  LAYER M2 ;
        RECT 3.244 23.432 5.716 23.464 ;
  LAYER M2 ;
        RECT 3.244 23.496 5.716 23.528 ;
  LAYER M2 ;
        RECT 3.244 23.56 5.716 23.592 ;
  LAYER M2 ;
        RECT 3.244 23.624 5.716 23.656 ;
  LAYER M3 ;
        RECT 3.264 21.3 3.296 23.808 ;
  LAYER M3 ;
        RECT 3.328 21.3 3.36 23.808 ;
  LAYER M3 ;
        RECT 3.392 21.3 3.424 23.808 ;
  LAYER M3 ;
        RECT 3.456 21.3 3.488 23.808 ;
  LAYER M3 ;
        RECT 3.52 21.3 3.552 23.808 ;
  LAYER M3 ;
        RECT 3.584 21.3 3.616 23.808 ;
  LAYER M3 ;
        RECT 3.648 21.3 3.68 23.808 ;
  LAYER M3 ;
        RECT 3.712 21.3 3.744 23.808 ;
  LAYER M3 ;
        RECT 3.776 21.3 3.808 23.808 ;
  LAYER M3 ;
        RECT 3.84 21.3 3.872 23.808 ;
  LAYER M3 ;
        RECT 3.904 21.3 3.936 23.808 ;
  LAYER M3 ;
        RECT 3.968 21.3 4 23.808 ;
  LAYER M3 ;
        RECT 4.032 21.3 4.064 23.808 ;
  LAYER M3 ;
        RECT 4.096 21.3 4.128 23.808 ;
  LAYER M3 ;
        RECT 4.16 21.3 4.192 23.808 ;
  LAYER M3 ;
        RECT 4.224 21.3 4.256 23.808 ;
  LAYER M3 ;
        RECT 4.288 21.3 4.32 23.808 ;
  LAYER M3 ;
        RECT 4.352 21.3 4.384 23.808 ;
  LAYER M3 ;
        RECT 4.416 21.3 4.448 23.808 ;
  LAYER M3 ;
        RECT 4.48 21.3 4.512 23.808 ;
  LAYER M3 ;
        RECT 4.544 21.3 4.576 23.808 ;
  LAYER M3 ;
        RECT 4.608 21.3 4.64 23.808 ;
  LAYER M3 ;
        RECT 4.672 21.3 4.704 23.808 ;
  LAYER M3 ;
        RECT 4.736 21.3 4.768 23.808 ;
  LAYER M3 ;
        RECT 4.8 21.3 4.832 23.808 ;
  LAYER M3 ;
        RECT 4.864 21.3 4.896 23.808 ;
  LAYER M3 ;
        RECT 4.928 21.3 4.96 23.808 ;
  LAYER M3 ;
        RECT 4.992 21.3 5.024 23.808 ;
  LAYER M3 ;
        RECT 5.056 21.3 5.088 23.808 ;
  LAYER M3 ;
        RECT 5.12 21.3 5.152 23.808 ;
  LAYER M3 ;
        RECT 5.184 21.3 5.216 23.808 ;
  LAYER M3 ;
        RECT 5.248 21.3 5.28 23.808 ;
  LAYER M3 ;
        RECT 5.312 21.3 5.344 23.808 ;
  LAYER M3 ;
        RECT 5.376 21.3 5.408 23.808 ;
  LAYER M3 ;
        RECT 5.44 21.3 5.472 23.808 ;
  LAYER M3 ;
        RECT 5.504 21.3 5.536 23.808 ;
  LAYER M3 ;
        RECT 5.568 21.3 5.6 23.808 ;
  LAYER M3 ;
        RECT 5.664 21.3 5.696 23.808 ;
  LAYER M1 ;
        RECT 3.279 21.336 3.281 23.772 ;
  LAYER M1 ;
        RECT 3.359 21.336 3.361 23.772 ;
  LAYER M1 ;
        RECT 3.439 21.336 3.441 23.772 ;
  LAYER M1 ;
        RECT 3.519 21.336 3.521 23.772 ;
  LAYER M1 ;
        RECT 3.599 21.336 3.601 23.772 ;
  LAYER M1 ;
        RECT 3.679 21.336 3.681 23.772 ;
  LAYER M1 ;
        RECT 3.759 21.336 3.761 23.772 ;
  LAYER M1 ;
        RECT 3.839 21.336 3.841 23.772 ;
  LAYER M1 ;
        RECT 3.919 21.336 3.921 23.772 ;
  LAYER M1 ;
        RECT 3.999 21.336 4.001 23.772 ;
  LAYER M1 ;
        RECT 4.079 21.336 4.081 23.772 ;
  LAYER M1 ;
        RECT 4.159 21.336 4.161 23.772 ;
  LAYER M1 ;
        RECT 4.239 21.336 4.241 23.772 ;
  LAYER M1 ;
        RECT 4.319 21.336 4.321 23.772 ;
  LAYER M1 ;
        RECT 4.399 21.336 4.401 23.772 ;
  LAYER M1 ;
        RECT 4.479 21.336 4.481 23.772 ;
  LAYER M1 ;
        RECT 4.559 21.336 4.561 23.772 ;
  LAYER M1 ;
        RECT 4.639 21.336 4.641 23.772 ;
  LAYER M1 ;
        RECT 4.719 21.336 4.721 23.772 ;
  LAYER M1 ;
        RECT 4.799 21.336 4.801 23.772 ;
  LAYER M1 ;
        RECT 4.879 21.336 4.881 23.772 ;
  LAYER M1 ;
        RECT 4.959 21.336 4.961 23.772 ;
  LAYER M1 ;
        RECT 5.039 21.336 5.041 23.772 ;
  LAYER M1 ;
        RECT 5.119 21.336 5.121 23.772 ;
  LAYER M1 ;
        RECT 5.199 21.336 5.201 23.772 ;
  LAYER M1 ;
        RECT 5.279 21.336 5.281 23.772 ;
  LAYER M1 ;
        RECT 5.359 21.336 5.361 23.772 ;
  LAYER M1 ;
        RECT 5.439 21.336 5.441 23.772 ;
  LAYER M1 ;
        RECT 5.519 21.336 5.521 23.772 ;
  LAYER M1 ;
        RECT 5.599 21.336 5.601 23.772 ;
  LAYER M2 ;
        RECT 3.28 21.335 5.68 21.337 ;
  LAYER M2 ;
        RECT 3.28 21.419 5.68 21.421 ;
  LAYER M2 ;
        RECT 3.28 21.503 5.68 21.505 ;
  LAYER M2 ;
        RECT 3.28 21.587 5.68 21.589 ;
  LAYER M2 ;
        RECT 3.28 21.671 5.68 21.673 ;
  LAYER M2 ;
        RECT 3.28 21.755 5.68 21.757 ;
  LAYER M2 ;
        RECT 3.28 21.839 5.68 21.841 ;
  LAYER M2 ;
        RECT 3.28 21.923 5.68 21.925 ;
  LAYER M2 ;
        RECT 3.28 22.007 5.68 22.009 ;
  LAYER M2 ;
        RECT 3.28 22.091 5.68 22.093 ;
  LAYER M2 ;
        RECT 3.28 22.175 5.68 22.177 ;
  LAYER M2 ;
        RECT 3.28 22.259 5.68 22.261 ;
  LAYER M2 ;
        RECT 3.28 22.3425 5.68 22.3445 ;
  LAYER M2 ;
        RECT 3.28 22.427 5.68 22.429 ;
  LAYER M2 ;
        RECT 3.28 22.511 5.68 22.513 ;
  LAYER M2 ;
        RECT 3.28 22.595 5.68 22.597 ;
  LAYER M2 ;
        RECT 3.28 22.679 5.68 22.681 ;
  LAYER M2 ;
        RECT 3.28 22.763 5.68 22.765 ;
  LAYER M2 ;
        RECT 3.28 22.847 5.68 22.849 ;
  LAYER M2 ;
        RECT 3.28 22.931 5.68 22.933 ;
  LAYER M2 ;
        RECT 3.28 23.015 5.68 23.017 ;
  LAYER M2 ;
        RECT 3.28 23.099 5.68 23.101 ;
  LAYER M2 ;
        RECT 3.28 23.183 5.68 23.185 ;
  LAYER M2 ;
        RECT 3.28 23.267 5.68 23.269 ;
  LAYER M2 ;
        RECT 3.28 23.351 5.68 23.353 ;
  LAYER M2 ;
        RECT 3.28 23.435 5.68 23.437 ;
  LAYER M2 ;
        RECT 3.28 23.519 5.68 23.521 ;
  LAYER M2 ;
        RECT 3.28 23.603 5.68 23.605 ;
  LAYER M2 ;
        RECT 3.28 23.687 5.68 23.689 ;
  LAYER M1 ;
        RECT 6.144 0.72 6.176 3.228 ;
  LAYER M1 ;
        RECT 6.208 0.72 6.24 3.228 ;
  LAYER M1 ;
        RECT 6.272 0.72 6.304 3.228 ;
  LAYER M1 ;
        RECT 6.336 0.72 6.368 3.228 ;
  LAYER M1 ;
        RECT 6.4 0.72 6.432 3.228 ;
  LAYER M1 ;
        RECT 6.464 0.72 6.496 3.228 ;
  LAYER M1 ;
        RECT 6.528 0.72 6.56 3.228 ;
  LAYER M1 ;
        RECT 6.592 0.72 6.624 3.228 ;
  LAYER M1 ;
        RECT 6.656 0.72 6.688 3.228 ;
  LAYER M1 ;
        RECT 6.72 0.72 6.752 3.228 ;
  LAYER M1 ;
        RECT 6.784 0.72 6.816 3.228 ;
  LAYER M1 ;
        RECT 6.848 0.72 6.88 3.228 ;
  LAYER M1 ;
        RECT 6.912 0.72 6.944 3.228 ;
  LAYER M1 ;
        RECT 6.976 0.72 7.008 3.228 ;
  LAYER M1 ;
        RECT 7.04 0.72 7.072 3.228 ;
  LAYER M1 ;
        RECT 7.104 0.72 7.136 3.228 ;
  LAYER M1 ;
        RECT 7.168 0.72 7.2 3.228 ;
  LAYER M1 ;
        RECT 7.232 0.72 7.264 3.228 ;
  LAYER M1 ;
        RECT 7.296 0.72 7.328 3.228 ;
  LAYER M1 ;
        RECT 7.36 0.72 7.392 3.228 ;
  LAYER M1 ;
        RECT 7.424 0.72 7.456 3.228 ;
  LAYER M1 ;
        RECT 7.488 0.72 7.52 3.228 ;
  LAYER M1 ;
        RECT 7.552 0.72 7.584 3.228 ;
  LAYER M1 ;
        RECT 7.616 0.72 7.648 3.228 ;
  LAYER M1 ;
        RECT 7.68 0.72 7.712 3.228 ;
  LAYER M1 ;
        RECT 7.744 0.72 7.776 3.228 ;
  LAYER M1 ;
        RECT 7.808 0.72 7.84 3.228 ;
  LAYER M1 ;
        RECT 7.872 0.72 7.904 3.228 ;
  LAYER M1 ;
        RECT 7.936 0.72 7.968 3.228 ;
  LAYER M1 ;
        RECT 8 0.72 8.032 3.228 ;
  LAYER M1 ;
        RECT 8.064 0.72 8.096 3.228 ;
  LAYER M1 ;
        RECT 8.128 0.72 8.16 3.228 ;
  LAYER M1 ;
        RECT 8.192 0.72 8.224 3.228 ;
  LAYER M1 ;
        RECT 8.256 0.72 8.288 3.228 ;
  LAYER M1 ;
        RECT 8.32 0.72 8.352 3.228 ;
  LAYER M1 ;
        RECT 8.384 0.72 8.416 3.228 ;
  LAYER M1 ;
        RECT 8.448 0.72 8.48 3.228 ;
  LAYER M2 ;
        RECT 6.124 0.804 8.596 0.836 ;
  LAYER M2 ;
        RECT 6.124 0.868 8.596 0.9 ;
  LAYER M2 ;
        RECT 6.124 0.932 8.596 0.964 ;
  LAYER M2 ;
        RECT 6.124 0.996 8.596 1.028 ;
  LAYER M2 ;
        RECT 6.124 1.06 8.596 1.092 ;
  LAYER M2 ;
        RECT 6.124 1.124 8.596 1.156 ;
  LAYER M2 ;
        RECT 6.124 1.188 8.596 1.22 ;
  LAYER M2 ;
        RECT 6.124 1.252 8.596 1.284 ;
  LAYER M2 ;
        RECT 6.124 1.316 8.596 1.348 ;
  LAYER M2 ;
        RECT 6.124 1.38 8.596 1.412 ;
  LAYER M2 ;
        RECT 6.124 1.444 8.596 1.476 ;
  LAYER M2 ;
        RECT 6.124 1.508 8.596 1.54 ;
  LAYER M2 ;
        RECT 6.124 1.572 8.596 1.604 ;
  LAYER M2 ;
        RECT 6.124 1.636 8.596 1.668 ;
  LAYER M2 ;
        RECT 6.124 1.7 8.596 1.732 ;
  LAYER M2 ;
        RECT 6.124 1.764 8.596 1.796 ;
  LAYER M2 ;
        RECT 6.124 1.828 8.596 1.86 ;
  LAYER M2 ;
        RECT 6.124 1.892 8.596 1.924 ;
  LAYER M2 ;
        RECT 6.124 1.956 8.596 1.988 ;
  LAYER M2 ;
        RECT 6.124 2.02 8.596 2.052 ;
  LAYER M2 ;
        RECT 6.124 2.084 8.596 2.116 ;
  LAYER M2 ;
        RECT 6.124 2.148 8.596 2.18 ;
  LAYER M2 ;
        RECT 6.124 2.212 8.596 2.244 ;
  LAYER M2 ;
        RECT 6.124 2.276 8.596 2.308 ;
  LAYER M2 ;
        RECT 6.124 2.34 8.596 2.372 ;
  LAYER M2 ;
        RECT 6.124 2.404 8.596 2.436 ;
  LAYER M2 ;
        RECT 6.124 2.468 8.596 2.5 ;
  LAYER M2 ;
        RECT 6.124 2.532 8.596 2.564 ;
  LAYER M2 ;
        RECT 6.124 2.596 8.596 2.628 ;
  LAYER M2 ;
        RECT 6.124 2.66 8.596 2.692 ;
  LAYER M2 ;
        RECT 6.124 2.724 8.596 2.756 ;
  LAYER M2 ;
        RECT 6.124 2.788 8.596 2.82 ;
  LAYER M2 ;
        RECT 6.124 2.852 8.596 2.884 ;
  LAYER M2 ;
        RECT 6.124 2.916 8.596 2.948 ;
  LAYER M2 ;
        RECT 6.124 2.98 8.596 3.012 ;
  LAYER M2 ;
        RECT 6.124 3.044 8.596 3.076 ;
  LAYER M3 ;
        RECT 6.144 0.72 6.176 3.228 ;
  LAYER M3 ;
        RECT 6.208 0.72 6.24 3.228 ;
  LAYER M3 ;
        RECT 6.272 0.72 6.304 3.228 ;
  LAYER M3 ;
        RECT 6.336 0.72 6.368 3.228 ;
  LAYER M3 ;
        RECT 6.4 0.72 6.432 3.228 ;
  LAYER M3 ;
        RECT 6.464 0.72 6.496 3.228 ;
  LAYER M3 ;
        RECT 6.528 0.72 6.56 3.228 ;
  LAYER M3 ;
        RECT 6.592 0.72 6.624 3.228 ;
  LAYER M3 ;
        RECT 6.656 0.72 6.688 3.228 ;
  LAYER M3 ;
        RECT 6.72 0.72 6.752 3.228 ;
  LAYER M3 ;
        RECT 6.784 0.72 6.816 3.228 ;
  LAYER M3 ;
        RECT 6.848 0.72 6.88 3.228 ;
  LAYER M3 ;
        RECT 6.912 0.72 6.944 3.228 ;
  LAYER M3 ;
        RECT 6.976 0.72 7.008 3.228 ;
  LAYER M3 ;
        RECT 7.04 0.72 7.072 3.228 ;
  LAYER M3 ;
        RECT 7.104 0.72 7.136 3.228 ;
  LAYER M3 ;
        RECT 7.168 0.72 7.2 3.228 ;
  LAYER M3 ;
        RECT 7.232 0.72 7.264 3.228 ;
  LAYER M3 ;
        RECT 7.296 0.72 7.328 3.228 ;
  LAYER M3 ;
        RECT 7.36 0.72 7.392 3.228 ;
  LAYER M3 ;
        RECT 7.424 0.72 7.456 3.228 ;
  LAYER M3 ;
        RECT 7.488 0.72 7.52 3.228 ;
  LAYER M3 ;
        RECT 7.552 0.72 7.584 3.228 ;
  LAYER M3 ;
        RECT 7.616 0.72 7.648 3.228 ;
  LAYER M3 ;
        RECT 7.68 0.72 7.712 3.228 ;
  LAYER M3 ;
        RECT 7.744 0.72 7.776 3.228 ;
  LAYER M3 ;
        RECT 7.808 0.72 7.84 3.228 ;
  LAYER M3 ;
        RECT 7.872 0.72 7.904 3.228 ;
  LAYER M3 ;
        RECT 7.936 0.72 7.968 3.228 ;
  LAYER M3 ;
        RECT 8 0.72 8.032 3.228 ;
  LAYER M3 ;
        RECT 8.064 0.72 8.096 3.228 ;
  LAYER M3 ;
        RECT 8.128 0.72 8.16 3.228 ;
  LAYER M3 ;
        RECT 8.192 0.72 8.224 3.228 ;
  LAYER M3 ;
        RECT 8.256 0.72 8.288 3.228 ;
  LAYER M3 ;
        RECT 8.32 0.72 8.352 3.228 ;
  LAYER M3 ;
        RECT 8.384 0.72 8.416 3.228 ;
  LAYER M3 ;
        RECT 8.448 0.72 8.48 3.228 ;
  LAYER M3 ;
        RECT 8.544 0.72 8.576 3.228 ;
  LAYER M1 ;
        RECT 6.159 0.756 6.161 3.192 ;
  LAYER M1 ;
        RECT 6.239 0.756 6.241 3.192 ;
  LAYER M1 ;
        RECT 6.319 0.756 6.321 3.192 ;
  LAYER M1 ;
        RECT 6.399 0.756 6.401 3.192 ;
  LAYER M1 ;
        RECT 6.479 0.756 6.481 3.192 ;
  LAYER M1 ;
        RECT 6.559 0.756 6.561 3.192 ;
  LAYER M1 ;
        RECT 6.639 0.756 6.641 3.192 ;
  LAYER M1 ;
        RECT 6.719 0.756 6.721 3.192 ;
  LAYER M1 ;
        RECT 6.799 0.756 6.801 3.192 ;
  LAYER M1 ;
        RECT 6.879 0.756 6.881 3.192 ;
  LAYER M1 ;
        RECT 6.959 0.756 6.961 3.192 ;
  LAYER M1 ;
        RECT 7.039 0.756 7.041 3.192 ;
  LAYER M1 ;
        RECT 7.119 0.756 7.121 3.192 ;
  LAYER M1 ;
        RECT 7.199 0.756 7.201 3.192 ;
  LAYER M1 ;
        RECT 7.279 0.756 7.281 3.192 ;
  LAYER M1 ;
        RECT 7.359 0.756 7.361 3.192 ;
  LAYER M1 ;
        RECT 7.439 0.756 7.441 3.192 ;
  LAYER M1 ;
        RECT 7.519 0.756 7.521 3.192 ;
  LAYER M1 ;
        RECT 7.599 0.756 7.601 3.192 ;
  LAYER M1 ;
        RECT 7.679 0.756 7.681 3.192 ;
  LAYER M1 ;
        RECT 7.759 0.756 7.761 3.192 ;
  LAYER M1 ;
        RECT 7.839 0.756 7.841 3.192 ;
  LAYER M1 ;
        RECT 7.919 0.756 7.921 3.192 ;
  LAYER M1 ;
        RECT 7.999 0.756 8.001 3.192 ;
  LAYER M1 ;
        RECT 8.079 0.756 8.081 3.192 ;
  LAYER M1 ;
        RECT 8.159 0.756 8.161 3.192 ;
  LAYER M1 ;
        RECT 8.239 0.756 8.241 3.192 ;
  LAYER M1 ;
        RECT 8.319 0.756 8.321 3.192 ;
  LAYER M1 ;
        RECT 8.399 0.756 8.401 3.192 ;
  LAYER M1 ;
        RECT 8.479 0.756 8.481 3.192 ;
  LAYER M2 ;
        RECT 6.16 0.755 8.56 0.757 ;
  LAYER M2 ;
        RECT 6.16 0.839 8.56 0.841 ;
  LAYER M2 ;
        RECT 6.16 0.923 8.56 0.925 ;
  LAYER M2 ;
        RECT 6.16 1.007 8.56 1.009 ;
  LAYER M2 ;
        RECT 6.16 1.091 8.56 1.093 ;
  LAYER M2 ;
        RECT 6.16 1.175 8.56 1.177 ;
  LAYER M2 ;
        RECT 6.16 1.259 8.56 1.261 ;
  LAYER M2 ;
        RECT 6.16 1.343 8.56 1.345 ;
  LAYER M2 ;
        RECT 6.16 1.427 8.56 1.429 ;
  LAYER M2 ;
        RECT 6.16 1.511 8.56 1.513 ;
  LAYER M2 ;
        RECT 6.16 1.595 8.56 1.597 ;
  LAYER M2 ;
        RECT 6.16 1.679 8.56 1.681 ;
  LAYER M2 ;
        RECT 6.16 1.7625 8.56 1.7645 ;
  LAYER M2 ;
        RECT 6.16 1.847 8.56 1.849 ;
  LAYER M2 ;
        RECT 6.16 1.931 8.56 1.933 ;
  LAYER M2 ;
        RECT 6.16 2.015 8.56 2.017 ;
  LAYER M2 ;
        RECT 6.16 2.099 8.56 2.101 ;
  LAYER M2 ;
        RECT 6.16 2.183 8.56 2.185 ;
  LAYER M2 ;
        RECT 6.16 2.267 8.56 2.269 ;
  LAYER M2 ;
        RECT 6.16 2.351 8.56 2.353 ;
  LAYER M2 ;
        RECT 6.16 2.435 8.56 2.437 ;
  LAYER M2 ;
        RECT 6.16 2.519 8.56 2.521 ;
  LAYER M2 ;
        RECT 6.16 2.603 8.56 2.605 ;
  LAYER M2 ;
        RECT 6.16 2.687 8.56 2.689 ;
  LAYER M2 ;
        RECT 6.16 2.771 8.56 2.773 ;
  LAYER M2 ;
        RECT 6.16 2.855 8.56 2.857 ;
  LAYER M2 ;
        RECT 6.16 2.939 8.56 2.941 ;
  LAYER M2 ;
        RECT 6.16 3.023 8.56 3.025 ;
  LAYER M2 ;
        RECT 6.16 3.107 8.56 3.109 ;
  LAYER M1 ;
        RECT 6.144 3.66 6.176 6.168 ;
  LAYER M1 ;
        RECT 6.208 3.66 6.24 6.168 ;
  LAYER M1 ;
        RECT 6.272 3.66 6.304 6.168 ;
  LAYER M1 ;
        RECT 6.336 3.66 6.368 6.168 ;
  LAYER M1 ;
        RECT 6.4 3.66 6.432 6.168 ;
  LAYER M1 ;
        RECT 6.464 3.66 6.496 6.168 ;
  LAYER M1 ;
        RECT 6.528 3.66 6.56 6.168 ;
  LAYER M1 ;
        RECT 6.592 3.66 6.624 6.168 ;
  LAYER M1 ;
        RECT 6.656 3.66 6.688 6.168 ;
  LAYER M1 ;
        RECT 6.72 3.66 6.752 6.168 ;
  LAYER M1 ;
        RECT 6.784 3.66 6.816 6.168 ;
  LAYER M1 ;
        RECT 6.848 3.66 6.88 6.168 ;
  LAYER M1 ;
        RECT 6.912 3.66 6.944 6.168 ;
  LAYER M1 ;
        RECT 6.976 3.66 7.008 6.168 ;
  LAYER M1 ;
        RECT 7.04 3.66 7.072 6.168 ;
  LAYER M1 ;
        RECT 7.104 3.66 7.136 6.168 ;
  LAYER M1 ;
        RECT 7.168 3.66 7.2 6.168 ;
  LAYER M1 ;
        RECT 7.232 3.66 7.264 6.168 ;
  LAYER M1 ;
        RECT 7.296 3.66 7.328 6.168 ;
  LAYER M1 ;
        RECT 7.36 3.66 7.392 6.168 ;
  LAYER M1 ;
        RECT 7.424 3.66 7.456 6.168 ;
  LAYER M1 ;
        RECT 7.488 3.66 7.52 6.168 ;
  LAYER M1 ;
        RECT 7.552 3.66 7.584 6.168 ;
  LAYER M1 ;
        RECT 7.616 3.66 7.648 6.168 ;
  LAYER M1 ;
        RECT 7.68 3.66 7.712 6.168 ;
  LAYER M1 ;
        RECT 7.744 3.66 7.776 6.168 ;
  LAYER M1 ;
        RECT 7.808 3.66 7.84 6.168 ;
  LAYER M1 ;
        RECT 7.872 3.66 7.904 6.168 ;
  LAYER M1 ;
        RECT 7.936 3.66 7.968 6.168 ;
  LAYER M1 ;
        RECT 8 3.66 8.032 6.168 ;
  LAYER M1 ;
        RECT 8.064 3.66 8.096 6.168 ;
  LAYER M1 ;
        RECT 8.128 3.66 8.16 6.168 ;
  LAYER M1 ;
        RECT 8.192 3.66 8.224 6.168 ;
  LAYER M1 ;
        RECT 8.256 3.66 8.288 6.168 ;
  LAYER M1 ;
        RECT 8.32 3.66 8.352 6.168 ;
  LAYER M1 ;
        RECT 8.384 3.66 8.416 6.168 ;
  LAYER M1 ;
        RECT 8.448 3.66 8.48 6.168 ;
  LAYER M2 ;
        RECT 6.124 3.744 8.596 3.776 ;
  LAYER M2 ;
        RECT 6.124 3.808 8.596 3.84 ;
  LAYER M2 ;
        RECT 6.124 3.872 8.596 3.904 ;
  LAYER M2 ;
        RECT 6.124 3.936 8.596 3.968 ;
  LAYER M2 ;
        RECT 6.124 4 8.596 4.032 ;
  LAYER M2 ;
        RECT 6.124 4.064 8.596 4.096 ;
  LAYER M2 ;
        RECT 6.124 4.128 8.596 4.16 ;
  LAYER M2 ;
        RECT 6.124 4.192 8.596 4.224 ;
  LAYER M2 ;
        RECT 6.124 4.256 8.596 4.288 ;
  LAYER M2 ;
        RECT 6.124 4.32 8.596 4.352 ;
  LAYER M2 ;
        RECT 6.124 4.384 8.596 4.416 ;
  LAYER M2 ;
        RECT 6.124 4.448 8.596 4.48 ;
  LAYER M2 ;
        RECT 6.124 4.512 8.596 4.544 ;
  LAYER M2 ;
        RECT 6.124 4.576 8.596 4.608 ;
  LAYER M2 ;
        RECT 6.124 4.64 8.596 4.672 ;
  LAYER M2 ;
        RECT 6.124 4.704 8.596 4.736 ;
  LAYER M2 ;
        RECT 6.124 4.768 8.596 4.8 ;
  LAYER M2 ;
        RECT 6.124 4.832 8.596 4.864 ;
  LAYER M2 ;
        RECT 6.124 4.896 8.596 4.928 ;
  LAYER M2 ;
        RECT 6.124 4.96 8.596 4.992 ;
  LAYER M2 ;
        RECT 6.124 5.024 8.596 5.056 ;
  LAYER M2 ;
        RECT 6.124 5.088 8.596 5.12 ;
  LAYER M2 ;
        RECT 6.124 5.152 8.596 5.184 ;
  LAYER M2 ;
        RECT 6.124 5.216 8.596 5.248 ;
  LAYER M2 ;
        RECT 6.124 5.28 8.596 5.312 ;
  LAYER M2 ;
        RECT 6.124 5.344 8.596 5.376 ;
  LAYER M2 ;
        RECT 6.124 5.408 8.596 5.44 ;
  LAYER M2 ;
        RECT 6.124 5.472 8.596 5.504 ;
  LAYER M2 ;
        RECT 6.124 5.536 8.596 5.568 ;
  LAYER M2 ;
        RECT 6.124 5.6 8.596 5.632 ;
  LAYER M2 ;
        RECT 6.124 5.664 8.596 5.696 ;
  LAYER M2 ;
        RECT 6.124 5.728 8.596 5.76 ;
  LAYER M2 ;
        RECT 6.124 5.792 8.596 5.824 ;
  LAYER M2 ;
        RECT 6.124 5.856 8.596 5.888 ;
  LAYER M2 ;
        RECT 6.124 5.92 8.596 5.952 ;
  LAYER M2 ;
        RECT 6.124 5.984 8.596 6.016 ;
  LAYER M3 ;
        RECT 6.144 3.66 6.176 6.168 ;
  LAYER M3 ;
        RECT 6.208 3.66 6.24 6.168 ;
  LAYER M3 ;
        RECT 6.272 3.66 6.304 6.168 ;
  LAYER M3 ;
        RECT 6.336 3.66 6.368 6.168 ;
  LAYER M3 ;
        RECT 6.4 3.66 6.432 6.168 ;
  LAYER M3 ;
        RECT 6.464 3.66 6.496 6.168 ;
  LAYER M3 ;
        RECT 6.528 3.66 6.56 6.168 ;
  LAYER M3 ;
        RECT 6.592 3.66 6.624 6.168 ;
  LAYER M3 ;
        RECT 6.656 3.66 6.688 6.168 ;
  LAYER M3 ;
        RECT 6.72 3.66 6.752 6.168 ;
  LAYER M3 ;
        RECT 6.784 3.66 6.816 6.168 ;
  LAYER M3 ;
        RECT 6.848 3.66 6.88 6.168 ;
  LAYER M3 ;
        RECT 6.912 3.66 6.944 6.168 ;
  LAYER M3 ;
        RECT 6.976 3.66 7.008 6.168 ;
  LAYER M3 ;
        RECT 7.04 3.66 7.072 6.168 ;
  LAYER M3 ;
        RECT 7.104 3.66 7.136 6.168 ;
  LAYER M3 ;
        RECT 7.168 3.66 7.2 6.168 ;
  LAYER M3 ;
        RECT 7.232 3.66 7.264 6.168 ;
  LAYER M3 ;
        RECT 7.296 3.66 7.328 6.168 ;
  LAYER M3 ;
        RECT 7.36 3.66 7.392 6.168 ;
  LAYER M3 ;
        RECT 7.424 3.66 7.456 6.168 ;
  LAYER M3 ;
        RECT 7.488 3.66 7.52 6.168 ;
  LAYER M3 ;
        RECT 7.552 3.66 7.584 6.168 ;
  LAYER M3 ;
        RECT 7.616 3.66 7.648 6.168 ;
  LAYER M3 ;
        RECT 7.68 3.66 7.712 6.168 ;
  LAYER M3 ;
        RECT 7.744 3.66 7.776 6.168 ;
  LAYER M3 ;
        RECT 7.808 3.66 7.84 6.168 ;
  LAYER M3 ;
        RECT 7.872 3.66 7.904 6.168 ;
  LAYER M3 ;
        RECT 7.936 3.66 7.968 6.168 ;
  LAYER M3 ;
        RECT 8 3.66 8.032 6.168 ;
  LAYER M3 ;
        RECT 8.064 3.66 8.096 6.168 ;
  LAYER M3 ;
        RECT 8.128 3.66 8.16 6.168 ;
  LAYER M3 ;
        RECT 8.192 3.66 8.224 6.168 ;
  LAYER M3 ;
        RECT 8.256 3.66 8.288 6.168 ;
  LAYER M3 ;
        RECT 8.32 3.66 8.352 6.168 ;
  LAYER M3 ;
        RECT 8.384 3.66 8.416 6.168 ;
  LAYER M3 ;
        RECT 8.448 3.66 8.48 6.168 ;
  LAYER M3 ;
        RECT 8.544 3.66 8.576 6.168 ;
  LAYER M1 ;
        RECT 6.159 3.696 6.161 6.132 ;
  LAYER M1 ;
        RECT 6.239 3.696 6.241 6.132 ;
  LAYER M1 ;
        RECT 6.319 3.696 6.321 6.132 ;
  LAYER M1 ;
        RECT 6.399 3.696 6.401 6.132 ;
  LAYER M1 ;
        RECT 6.479 3.696 6.481 6.132 ;
  LAYER M1 ;
        RECT 6.559 3.696 6.561 6.132 ;
  LAYER M1 ;
        RECT 6.639 3.696 6.641 6.132 ;
  LAYER M1 ;
        RECT 6.719 3.696 6.721 6.132 ;
  LAYER M1 ;
        RECT 6.799 3.696 6.801 6.132 ;
  LAYER M1 ;
        RECT 6.879 3.696 6.881 6.132 ;
  LAYER M1 ;
        RECT 6.959 3.696 6.961 6.132 ;
  LAYER M1 ;
        RECT 7.039 3.696 7.041 6.132 ;
  LAYER M1 ;
        RECT 7.119 3.696 7.121 6.132 ;
  LAYER M1 ;
        RECT 7.199 3.696 7.201 6.132 ;
  LAYER M1 ;
        RECT 7.279 3.696 7.281 6.132 ;
  LAYER M1 ;
        RECT 7.359 3.696 7.361 6.132 ;
  LAYER M1 ;
        RECT 7.439 3.696 7.441 6.132 ;
  LAYER M1 ;
        RECT 7.519 3.696 7.521 6.132 ;
  LAYER M1 ;
        RECT 7.599 3.696 7.601 6.132 ;
  LAYER M1 ;
        RECT 7.679 3.696 7.681 6.132 ;
  LAYER M1 ;
        RECT 7.759 3.696 7.761 6.132 ;
  LAYER M1 ;
        RECT 7.839 3.696 7.841 6.132 ;
  LAYER M1 ;
        RECT 7.919 3.696 7.921 6.132 ;
  LAYER M1 ;
        RECT 7.999 3.696 8.001 6.132 ;
  LAYER M1 ;
        RECT 8.079 3.696 8.081 6.132 ;
  LAYER M1 ;
        RECT 8.159 3.696 8.161 6.132 ;
  LAYER M1 ;
        RECT 8.239 3.696 8.241 6.132 ;
  LAYER M1 ;
        RECT 8.319 3.696 8.321 6.132 ;
  LAYER M1 ;
        RECT 8.399 3.696 8.401 6.132 ;
  LAYER M1 ;
        RECT 8.479 3.696 8.481 6.132 ;
  LAYER M2 ;
        RECT 6.16 3.695 8.56 3.697 ;
  LAYER M2 ;
        RECT 6.16 3.779 8.56 3.781 ;
  LAYER M2 ;
        RECT 6.16 3.863 8.56 3.865 ;
  LAYER M2 ;
        RECT 6.16 3.947 8.56 3.949 ;
  LAYER M2 ;
        RECT 6.16 4.031 8.56 4.033 ;
  LAYER M2 ;
        RECT 6.16 4.115 8.56 4.117 ;
  LAYER M2 ;
        RECT 6.16 4.199 8.56 4.201 ;
  LAYER M2 ;
        RECT 6.16 4.283 8.56 4.285 ;
  LAYER M2 ;
        RECT 6.16 4.367 8.56 4.369 ;
  LAYER M2 ;
        RECT 6.16 4.451 8.56 4.453 ;
  LAYER M2 ;
        RECT 6.16 4.535 8.56 4.537 ;
  LAYER M2 ;
        RECT 6.16 4.619 8.56 4.621 ;
  LAYER M2 ;
        RECT 6.16 4.7025 8.56 4.7045 ;
  LAYER M2 ;
        RECT 6.16 4.787 8.56 4.789 ;
  LAYER M2 ;
        RECT 6.16 4.871 8.56 4.873 ;
  LAYER M2 ;
        RECT 6.16 4.955 8.56 4.957 ;
  LAYER M2 ;
        RECT 6.16 5.039 8.56 5.041 ;
  LAYER M2 ;
        RECT 6.16 5.123 8.56 5.125 ;
  LAYER M2 ;
        RECT 6.16 5.207 8.56 5.209 ;
  LAYER M2 ;
        RECT 6.16 5.291 8.56 5.293 ;
  LAYER M2 ;
        RECT 6.16 5.375 8.56 5.377 ;
  LAYER M2 ;
        RECT 6.16 5.459 8.56 5.461 ;
  LAYER M2 ;
        RECT 6.16 5.543 8.56 5.545 ;
  LAYER M2 ;
        RECT 6.16 5.627 8.56 5.629 ;
  LAYER M2 ;
        RECT 6.16 5.711 8.56 5.713 ;
  LAYER M2 ;
        RECT 6.16 5.795 8.56 5.797 ;
  LAYER M2 ;
        RECT 6.16 5.879 8.56 5.881 ;
  LAYER M2 ;
        RECT 6.16 5.963 8.56 5.965 ;
  LAYER M2 ;
        RECT 6.16 6.047 8.56 6.049 ;
  LAYER M1 ;
        RECT 6.144 6.6 6.176 9.108 ;
  LAYER M1 ;
        RECT 6.208 6.6 6.24 9.108 ;
  LAYER M1 ;
        RECT 6.272 6.6 6.304 9.108 ;
  LAYER M1 ;
        RECT 6.336 6.6 6.368 9.108 ;
  LAYER M1 ;
        RECT 6.4 6.6 6.432 9.108 ;
  LAYER M1 ;
        RECT 6.464 6.6 6.496 9.108 ;
  LAYER M1 ;
        RECT 6.528 6.6 6.56 9.108 ;
  LAYER M1 ;
        RECT 6.592 6.6 6.624 9.108 ;
  LAYER M1 ;
        RECT 6.656 6.6 6.688 9.108 ;
  LAYER M1 ;
        RECT 6.72 6.6 6.752 9.108 ;
  LAYER M1 ;
        RECT 6.784 6.6 6.816 9.108 ;
  LAYER M1 ;
        RECT 6.848 6.6 6.88 9.108 ;
  LAYER M1 ;
        RECT 6.912 6.6 6.944 9.108 ;
  LAYER M1 ;
        RECT 6.976 6.6 7.008 9.108 ;
  LAYER M1 ;
        RECT 7.04 6.6 7.072 9.108 ;
  LAYER M1 ;
        RECT 7.104 6.6 7.136 9.108 ;
  LAYER M1 ;
        RECT 7.168 6.6 7.2 9.108 ;
  LAYER M1 ;
        RECT 7.232 6.6 7.264 9.108 ;
  LAYER M1 ;
        RECT 7.296 6.6 7.328 9.108 ;
  LAYER M1 ;
        RECT 7.36 6.6 7.392 9.108 ;
  LAYER M1 ;
        RECT 7.424 6.6 7.456 9.108 ;
  LAYER M1 ;
        RECT 7.488 6.6 7.52 9.108 ;
  LAYER M1 ;
        RECT 7.552 6.6 7.584 9.108 ;
  LAYER M1 ;
        RECT 7.616 6.6 7.648 9.108 ;
  LAYER M1 ;
        RECT 7.68 6.6 7.712 9.108 ;
  LAYER M1 ;
        RECT 7.744 6.6 7.776 9.108 ;
  LAYER M1 ;
        RECT 7.808 6.6 7.84 9.108 ;
  LAYER M1 ;
        RECT 7.872 6.6 7.904 9.108 ;
  LAYER M1 ;
        RECT 7.936 6.6 7.968 9.108 ;
  LAYER M1 ;
        RECT 8 6.6 8.032 9.108 ;
  LAYER M1 ;
        RECT 8.064 6.6 8.096 9.108 ;
  LAYER M1 ;
        RECT 8.128 6.6 8.16 9.108 ;
  LAYER M1 ;
        RECT 8.192 6.6 8.224 9.108 ;
  LAYER M1 ;
        RECT 8.256 6.6 8.288 9.108 ;
  LAYER M1 ;
        RECT 8.32 6.6 8.352 9.108 ;
  LAYER M1 ;
        RECT 8.384 6.6 8.416 9.108 ;
  LAYER M1 ;
        RECT 8.448 6.6 8.48 9.108 ;
  LAYER M2 ;
        RECT 6.124 6.684 8.596 6.716 ;
  LAYER M2 ;
        RECT 6.124 6.748 8.596 6.78 ;
  LAYER M2 ;
        RECT 6.124 6.812 8.596 6.844 ;
  LAYER M2 ;
        RECT 6.124 6.876 8.596 6.908 ;
  LAYER M2 ;
        RECT 6.124 6.94 8.596 6.972 ;
  LAYER M2 ;
        RECT 6.124 7.004 8.596 7.036 ;
  LAYER M2 ;
        RECT 6.124 7.068 8.596 7.1 ;
  LAYER M2 ;
        RECT 6.124 7.132 8.596 7.164 ;
  LAYER M2 ;
        RECT 6.124 7.196 8.596 7.228 ;
  LAYER M2 ;
        RECT 6.124 7.26 8.596 7.292 ;
  LAYER M2 ;
        RECT 6.124 7.324 8.596 7.356 ;
  LAYER M2 ;
        RECT 6.124 7.388 8.596 7.42 ;
  LAYER M2 ;
        RECT 6.124 7.452 8.596 7.484 ;
  LAYER M2 ;
        RECT 6.124 7.516 8.596 7.548 ;
  LAYER M2 ;
        RECT 6.124 7.58 8.596 7.612 ;
  LAYER M2 ;
        RECT 6.124 7.644 8.596 7.676 ;
  LAYER M2 ;
        RECT 6.124 7.708 8.596 7.74 ;
  LAYER M2 ;
        RECT 6.124 7.772 8.596 7.804 ;
  LAYER M2 ;
        RECT 6.124 7.836 8.596 7.868 ;
  LAYER M2 ;
        RECT 6.124 7.9 8.596 7.932 ;
  LAYER M2 ;
        RECT 6.124 7.964 8.596 7.996 ;
  LAYER M2 ;
        RECT 6.124 8.028 8.596 8.06 ;
  LAYER M2 ;
        RECT 6.124 8.092 8.596 8.124 ;
  LAYER M2 ;
        RECT 6.124 8.156 8.596 8.188 ;
  LAYER M2 ;
        RECT 6.124 8.22 8.596 8.252 ;
  LAYER M2 ;
        RECT 6.124 8.284 8.596 8.316 ;
  LAYER M2 ;
        RECT 6.124 8.348 8.596 8.38 ;
  LAYER M2 ;
        RECT 6.124 8.412 8.596 8.444 ;
  LAYER M2 ;
        RECT 6.124 8.476 8.596 8.508 ;
  LAYER M2 ;
        RECT 6.124 8.54 8.596 8.572 ;
  LAYER M2 ;
        RECT 6.124 8.604 8.596 8.636 ;
  LAYER M2 ;
        RECT 6.124 8.668 8.596 8.7 ;
  LAYER M2 ;
        RECT 6.124 8.732 8.596 8.764 ;
  LAYER M2 ;
        RECT 6.124 8.796 8.596 8.828 ;
  LAYER M2 ;
        RECT 6.124 8.86 8.596 8.892 ;
  LAYER M2 ;
        RECT 6.124 8.924 8.596 8.956 ;
  LAYER M3 ;
        RECT 6.144 6.6 6.176 9.108 ;
  LAYER M3 ;
        RECT 6.208 6.6 6.24 9.108 ;
  LAYER M3 ;
        RECT 6.272 6.6 6.304 9.108 ;
  LAYER M3 ;
        RECT 6.336 6.6 6.368 9.108 ;
  LAYER M3 ;
        RECT 6.4 6.6 6.432 9.108 ;
  LAYER M3 ;
        RECT 6.464 6.6 6.496 9.108 ;
  LAYER M3 ;
        RECT 6.528 6.6 6.56 9.108 ;
  LAYER M3 ;
        RECT 6.592 6.6 6.624 9.108 ;
  LAYER M3 ;
        RECT 6.656 6.6 6.688 9.108 ;
  LAYER M3 ;
        RECT 6.72 6.6 6.752 9.108 ;
  LAYER M3 ;
        RECT 6.784 6.6 6.816 9.108 ;
  LAYER M3 ;
        RECT 6.848 6.6 6.88 9.108 ;
  LAYER M3 ;
        RECT 6.912 6.6 6.944 9.108 ;
  LAYER M3 ;
        RECT 6.976 6.6 7.008 9.108 ;
  LAYER M3 ;
        RECT 7.04 6.6 7.072 9.108 ;
  LAYER M3 ;
        RECT 7.104 6.6 7.136 9.108 ;
  LAYER M3 ;
        RECT 7.168 6.6 7.2 9.108 ;
  LAYER M3 ;
        RECT 7.232 6.6 7.264 9.108 ;
  LAYER M3 ;
        RECT 7.296 6.6 7.328 9.108 ;
  LAYER M3 ;
        RECT 7.36 6.6 7.392 9.108 ;
  LAYER M3 ;
        RECT 7.424 6.6 7.456 9.108 ;
  LAYER M3 ;
        RECT 7.488 6.6 7.52 9.108 ;
  LAYER M3 ;
        RECT 7.552 6.6 7.584 9.108 ;
  LAYER M3 ;
        RECT 7.616 6.6 7.648 9.108 ;
  LAYER M3 ;
        RECT 7.68 6.6 7.712 9.108 ;
  LAYER M3 ;
        RECT 7.744 6.6 7.776 9.108 ;
  LAYER M3 ;
        RECT 7.808 6.6 7.84 9.108 ;
  LAYER M3 ;
        RECT 7.872 6.6 7.904 9.108 ;
  LAYER M3 ;
        RECT 7.936 6.6 7.968 9.108 ;
  LAYER M3 ;
        RECT 8 6.6 8.032 9.108 ;
  LAYER M3 ;
        RECT 8.064 6.6 8.096 9.108 ;
  LAYER M3 ;
        RECT 8.128 6.6 8.16 9.108 ;
  LAYER M3 ;
        RECT 8.192 6.6 8.224 9.108 ;
  LAYER M3 ;
        RECT 8.256 6.6 8.288 9.108 ;
  LAYER M3 ;
        RECT 8.32 6.6 8.352 9.108 ;
  LAYER M3 ;
        RECT 8.384 6.6 8.416 9.108 ;
  LAYER M3 ;
        RECT 8.448 6.6 8.48 9.108 ;
  LAYER M3 ;
        RECT 8.544 6.6 8.576 9.108 ;
  LAYER M1 ;
        RECT 6.159 6.636 6.161 9.072 ;
  LAYER M1 ;
        RECT 6.239 6.636 6.241 9.072 ;
  LAYER M1 ;
        RECT 6.319 6.636 6.321 9.072 ;
  LAYER M1 ;
        RECT 6.399 6.636 6.401 9.072 ;
  LAYER M1 ;
        RECT 6.479 6.636 6.481 9.072 ;
  LAYER M1 ;
        RECT 6.559 6.636 6.561 9.072 ;
  LAYER M1 ;
        RECT 6.639 6.636 6.641 9.072 ;
  LAYER M1 ;
        RECT 6.719 6.636 6.721 9.072 ;
  LAYER M1 ;
        RECT 6.799 6.636 6.801 9.072 ;
  LAYER M1 ;
        RECT 6.879 6.636 6.881 9.072 ;
  LAYER M1 ;
        RECT 6.959 6.636 6.961 9.072 ;
  LAYER M1 ;
        RECT 7.039 6.636 7.041 9.072 ;
  LAYER M1 ;
        RECT 7.119 6.636 7.121 9.072 ;
  LAYER M1 ;
        RECT 7.199 6.636 7.201 9.072 ;
  LAYER M1 ;
        RECT 7.279 6.636 7.281 9.072 ;
  LAYER M1 ;
        RECT 7.359 6.636 7.361 9.072 ;
  LAYER M1 ;
        RECT 7.439 6.636 7.441 9.072 ;
  LAYER M1 ;
        RECT 7.519 6.636 7.521 9.072 ;
  LAYER M1 ;
        RECT 7.599 6.636 7.601 9.072 ;
  LAYER M1 ;
        RECT 7.679 6.636 7.681 9.072 ;
  LAYER M1 ;
        RECT 7.759 6.636 7.761 9.072 ;
  LAYER M1 ;
        RECT 7.839 6.636 7.841 9.072 ;
  LAYER M1 ;
        RECT 7.919 6.636 7.921 9.072 ;
  LAYER M1 ;
        RECT 7.999 6.636 8.001 9.072 ;
  LAYER M1 ;
        RECT 8.079 6.636 8.081 9.072 ;
  LAYER M1 ;
        RECT 8.159 6.636 8.161 9.072 ;
  LAYER M1 ;
        RECT 8.239 6.636 8.241 9.072 ;
  LAYER M1 ;
        RECT 8.319 6.636 8.321 9.072 ;
  LAYER M1 ;
        RECT 8.399 6.636 8.401 9.072 ;
  LAYER M1 ;
        RECT 8.479 6.636 8.481 9.072 ;
  LAYER M2 ;
        RECT 6.16 6.635 8.56 6.637 ;
  LAYER M2 ;
        RECT 6.16 6.719 8.56 6.721 ;
  LAYER M2 ;
        RECT 6.16 6.803 8.56 6.805 ;
  LAYER M2 ;
        RECT 6.16 6.887 8.56 6.889 ;
  LAYER M2 ;
        RECT 6.16 6.971 8.56 6.973 ;
  LAYER M2 ;
        RECT 6.16 7.055 8.56 7.057 ;
  LAYER M2 ;
        RECT 6.16 7.139 8.56 7.141 ;
  LAYER M2 ;
        RECT 6.16 7.223 8.56 7.225 ;
  LAYER M2 ;
        RECT 6.16 7.307 8.56 7.309 ;
  LAYER M2 ;
        RECT 6.16 7.391 8.56 7.393 ;
  LAYER M2 ;
        RECT 6.16 7.475 8.56 7.477 ;
  LAYER M2 ;
        RECT 6.16 7.559 8.56 7.561 ;
  LAYER M2 ;
        RECT 6.16 7.6425 8.56 7.6445 ;
  LAYER M2 ;
        RECT 6.16 7.727 8.56 7.729 ;
  LAYER M2 ;
        RECT 6.16 7.811 8.56 7.813 ;
  LAYER M2 ;
        RECT 6.16 7.895 8.56 7.897 ;
  LAYER M2 ;
        RECT 6.16 7.979 8.56 7.981 ;
  LAYER M2 ;
        RECT 6.16 8.063 8.56 8.065 ;
  LAYER M2 ;
        RECT 6.16 8.147 8.56 8.149 ;
  LAYER M2 ;
        RECT 6.16 8.231 8.56 8.233 ;
  LAYER M2 ;
        RECT 6.16 8.315 8.56 8.317 ;
  LAYER M2 ;
        RECT 6.16 8.399 8.56 8.401 ;
  LAYER M2 ;
        RECT 6.16 8.483 8.56 8.485 ;
  LAYER M2 ;
        RECT 6.16 8.567 8.56 8.569 ;
  LAYER M2 ;
        RECT 6.16 8.651 8.56 8.653 ;
  LAYER M2 ;
        RECT 6.16 8.735 8.56 8.737 ;
  LAYER M2 ;
        RECT 6.16 8.819 8.56 8.821 ;
  LAYER M2 ;
        RECT 6.16 8.903 8.56 8.905 ;
  LAYER M2 ;
        RECT 6.16 8.987 8.56 8.989 ;
  LAYER M1 ;
        RECT 6.144 9.54 6.176 12.048 ;
  LAYER M1 ;
        RECT 6.208 9.54 6.24 12.048 ;
  LAYER M1 ;
        RECT 6.272 9.54 6.304 12.048 ;
  LAYER M1 ;
        RECT 6.336 9.54 6.368 12.048 ;
  LAYER M1 ;
        RECT 6.4 9.54 6.432 12.048 ;
  LAYER M1 ;
        RECT 6.464 9.54 6.496 12.048 ;
  LAYER M1 ;
        RECT 6.528 9.54 6.56 12.048 ;
  LAYER M1 ;
        RECT 6.592 9.54 6.624 12.048 ;
  LAYER M1 ;
        RECT 6.656 9.54 6.688 12.048 ;
  LAYER M1 ;
        RECT 6.72 9.54 6.752 12.048 ;
  LAYER M1 ;
        RECT 6.784 9.54 6.816 12.048 ;
  LAYER M1 ;
        RECT 6.848 9.54 6.88 12.048 ;
  LAYER M1 ;
        RECT 6.912 9.54 6.944 12.048 ;
  LAYER M1 ;
        RECT 6.976 9.54 7.008 12.048 ;
  LAYER M1 ;
        RECT 7.04 9.54 7.072 12.048 ;
  LAYER M1 ;
        RECT 7.104 9.54 7.136 12.048 ;
  LAYER M1 ;
        RECT 7.168 9.54 7.2 12.048 ;
  LAYER M1 ;
        RECT 7.232 9.54 7.264 12.048 ;
  LAYER M1 ;
        RECT 7.296 9.54 7.328 12.048 ;
  LAYER M1 ;
        RECT 7.36 9.54 7.392 12.048 ;
  LAYER M1 ;
        RECT 7.424 9.54 7.456 12.048 ;
  LAYER M1 ;
        RECT 7.488 9.54 7.52 12.048 ;
  LAYER M1 ;
        RECT 7.552 9.54 7.584 12.048 ;
  LAYER M1 ;
        RECT 7.616 9.54 7.648 12.048 ;
  LAYER M1 ;
        RECT 7.68 9.54 7.712 12.048 ;
  LAYER M1 ;
        RECT 7.744 9.54 7.776 12.048 ;
  LAYER M1 ;
        RECT 7.808 9.54 7.84 12.048 ;
  LAYER M1 ;
        RECT 7.872 9.54 7.904 12.048 ;
  LAYER M1 ;
        RECT 7.936 9.54 7.968 12.048 ;
  LAYER M1 ;
        RECT 8 9.54 8.032 12.048 ;
  LAYER M1 ;
        RECT 8.064 9.54 8.096 12.048 ;
  LAYER M1 ;
        RECT 8.128 9.54 8.16 12.048 ;
  LAYER M1 ;
        RECT 8.192 9.54 8.224 12.048 ;
  LAYER M1 ;
        RECT 8.256 9.54 8.288 12.048 ;
  LAYER M1 ;
        RECT 8.32 9.54 8.352 12.048 ;
  LAYER M1 ;
        RECT 8.384 9.54 8.416 12.048 ;
  LAYER M1 ;
        RECT 8.448 9.54 8.48 12.048 ;
  LAYER M2 ;
        RECT 6.124 9.624 8.596 9.656 ;
  LAYER M2 ;
        RECT 6.124 9.688 8.596 9.72 ;
  LAYER M2 ;
        RECT 6.124 9.752 8.596 9.784 ;
  LAYER M2 ;
        RECT 6.124 9.816 8.596 9.848 ;
  LAYER M2 ;
        RECT 6.124 9.88 8.596 9.912 ;
  LAYER M2 ;
        RECT 6.124 9.944 8.596 9.976 ;
  LAYER M2 ;
        RECT 6.124 10.008 8.596 10.04 ;
  LAYER M2 ;
        RECT 6.124 10.072 8.596 10.104 ;
  LAYER M2 ;
        RECT 6.124 10.136 8.596 10.168 ;
  LAYER M2 ;
        RECT 6.124 10.2 8.596 10.232 ;
  LAYER M2 ;
        RECT 6.124 10.264 8.596 10.296 ;
  LAYER M2 ;
        RECT 6.124 10.328 8.596 10.36 ;
  LAYER M2 ;
        RECT 6.124 10.392 8.596 10.424 ;
  LAYER M2 ;
        RECT 6.124 10.456 8.596 10.488 ;
  LAYER M2 ;
        RECT 6.124 10.52 8.596 10.552 ;
  LAYER M2 ;
        RECT 6.124 10.584 8.596 10.616 ;
  LAYER M2 ;
        RECT 6.124 10.648 8.596 10.68 ;
  LAYER M2 ;
        RECT 6.124 10.712 8.596 10.744 ;
  LAYER M2 ;
        RECT 6.124 10.776 8.596 10.808 ;
  LAYER M2 ;
        RECT 6.124 10.84 8.596 10.872 ;
  LAYER M2 ;
        RECT 6.124 10.904 8.596 10.936 ;
  LAYER M2 ;
        RECT 6.124 10.968 8.596 11 ;
  LAYER M2 ;
        RECT 6.124 11.032 8.596 11.064 ;
  LAYER M2 ;
        RECT 6.124 11.096 8.596 11.128 ;
  LAYER M2 ;
        RECT 6.124 11.16 8.596 11.192 ;
  LAYER M2 ;
        RECT 6.124 11.224 8.596 11.256 ;
  LAYER M2 ;
        RECT 6.124 11.288 8.596 11.32 ;
  LAYER M2 ;
        RECT 6.124 11.352 8.596 11.384 ;
  LAYER M2 ;
        RECT 6.124 11.416 8.596 11.448 ;
  LAYER M2 ;
        RECT 6.124 11.48 8.596 11.512 ;
  LAYER M2 ;
        RECT 6.124 11.544 8.596 11.576 ;
  LAYER M2 ;
        RECT 6.124 11.608 8.596 11.64 ;
  LAYER M2 ;
        RECT 6.124 11.672 8.596 11.704 ;
  LAYER M2 ;
        RECT 6.124 11.736 8.596 11.768 ;
  LAYER M2 ;
        RECT 6.124 11.8 8.596 11.832 ;
  LAYER M2 ;
        RECT 6.124 11.864 8.596 11.896 ;
  LAYER M3 ;
        RECT 6.144 9.54 6.176 12.048 ;
  LAYER M3 ;
        RECT 6.208 9.54 6.24 12.048 ;
  LAYER M3 ;
        RECT 6.272 9.54 6.304 12.048 ;
  LAYER M3 ;
        RECT 6.336 9.54 6.368 12.048 ;
  LAYER M3 ;
        RECT 6.4 9.54 6.432 12.048 ;
  LAYER M3 ;
        RECT 6.464 9.54 6.496 12.048 ;
  LAYER M3 ;
        RECT 6.528 9.54 6.56 12.048 ;
  LAYER M3 ;
        RECT 6.592 9.54 6.624 12.048 ;
  LAYER M3 ;
        RECT 6.656 9.54 6.688 12.048 ;
  LAYER M3 ;
        RECT 6.72 9.54 6.752 12.048 ;
  LAYER M3 ;
        RECT 6.784 9.54 6.816 12.048 ;
  LAYER M3 ;
        RECT 6.848 9.54 6.88 12.048 ;
  LAYER M3 ;
        RECT 6.912 9.54 6.944 12.048 ;
  LAYER M3 ;
        RECT 6.976 9.54 7.008 12.048 ;
  LAYER M3 ;
        RECT 7.04 9.54 7.072 12.048 ;
  LAYER M3 ;
        RECT 7.104 9.54 7.136 12.048 ;
  LAYER M3 ;
        RECT 7.168 9.54 7.2 12.048 ;
  LAYER M3 ;
        RECT 7.232 9.54 7.264 12.048 ;
  LAYER M3 ;
        RECT 7.296 9.54 7.328 12.048 ;
  LAYER M3 ;
        RECT 7.36 9.54 7.392 12.048 ;
  LAYER M3 ;
        RECT 7.424 9.54 7.456 12.048 ;
  LAYER M3 ;
        RECT 7.488 9.54 7.52 12.048 ;
  LAYER M3 ;
        RECT 7.552 9.54 7.584 12.048 ;
  LAYER M3 ;
        RECT 7.616 9.54 7.648 12.048 ;
  LAYER M3 ;
        RECT 7.68 9.54 7.712 12.048 ;
  LAYER M3 ;
        RECT 7.744 9.54 7.776 12.048 ;
  LAYER M3 ;
        RECT 7.808 9.54 7.84 12.048 ;
  LAYER M3 ;
        RECT 7.872 9.54 7.904 12.048 ;
  LAYER M3 ;
        RECT 7.936 9.54 7.968 12.048 ;
  LAYER M3 ;
        RECT 8 9.54 8.032 12.048 ;
  LAYER M3 ;
        RECT 8.064 9.54 8.096 12.048 ;
  LAYER M3 ;
        RECT 8.128 9.54 8.16 12.048 ;
  LAYER M3 ;
        RECT 8.192 9.54 8.224 12.048 ;
  LAYER M3 ;
        RECT 8.256 9.54 8.288 12.048 ;
  LAYER M3 ;
        RECT 8.32 9.54 8.352 12.048 ;
  LAYER M3 ;
        RECT 8.384 9.54 8.416 12.048 ;
  LAYER M3 ;
        RECT 8.448 9.54 8.48 12.048 ;
  LAYER M3 ;
        RECT 8.544 9.54 8.576 12.048 ;
  LAYER M1 ;
        RECT 6.159 9.576 6.161 12.012 ;
  LAYER M1 ;
        RECT 6.239 9.576 6.241 12.012 ;
  LAYER M1 ;
        RECT 6.319 9.576 6.321 12.012 ;
  LAYER M1 ;
        RECT 6.399 9.576 6.401 12.012 ;
  LAYER M1 ;
        RECT 6.479 9.576 6.481 12.012 ;
  LAYER M1 ;
        RECT 6.559 9.576 6.561 12.012 ;
  LAYER M1 ;
        RECT 6.639 9.576 6.641 12.012 ;
  LAYER M1 ;
        RECT 6.719 9.576 6.721 12.012 ;
  LAYER M1 ;
        RECT 6.799 9.576 6.801 12.012 ;
  LAYER M1 ;
        RECT 6.879 9.576 6.881 12.012 ;
  LAYER M1 ;
        RECT 6.959 9.576 6.961 12.012 ;
  LAYER M1 ;
        RECT 7.039 9.576 7.041 12.012 ;
  LAYER M1 ;
        RECT 7.119 9.576 7.121 12.012 ;
  LAYER M1 ;
        RECT 7.199 9.576 7.201 12.012 ;
  LAYER M1 ;
        RECT 7.279 9.576 7.281 12.012 ;
  LAYER M1 ;
        RECT 7.359 9.576 7.361 12.012 ;
  LAYER M1 ;
        RECT 7.439 9.576 7.441 12.012 ;
  LAYER M1 ;
        RECT 7.519 9.576 7.521 12.012 ;
  LAYER M1 ;
        RECT 7.599 9.576 7.601 12.012 ;
  LAYER M1 ;
        RECT 7.679 9.576 7.681 12.012 ;
  LAYER M1 ;
        RECT 7.759 9.576 7.761 12.012 ;
  LAYER M1 ;
        RECT 7.839 9.576 7.841 12.012 ;
  LAYER M1 ;
        RECT 7.919 9.576 7.921 12.012 ;
  LAYER M1 ;
        RECT 7.999 9.576 8.001 12.012 ;
  LAYER M1 ;
        RECT 8.079 9.576 8.081 12.012 ;
  LAYER M1 ;
        RECT 8.159 9.576 8.161 12.012 ;
  LAYER M1 ;
        RECT 8.239 9.576 8.241 12.012 ;
  LAYER M1 ;
        RECT 8.319 9.576 8.321 12.012 ;
  LAYER M1 ;
        RECT 8.399 9.576 8.401 12.012 ;
  LAYER M1 ;
        RECT 8.479 9.576 8.481 12.012 ;
  LAYER M2 ;
        RECT 6.16 9.575 8.56 9.577 ;
  LAYER M2 ;
        RECT 6.16 9.659 8.56 9.661 ;
  LAYER M2 ;
        RECT 6.16 9.743 8.56 9.745 ;
  LAYER M2 ;
        RECT 6.16 9.827 8.56 9.829 ;
  LAYER M2 ;
        RECT 6.16 9.911 8.56 9.913 ;
  LAYER M2 ;
        RECT 6.16 9.995 8.56 9.997 ;
  LAYER M2 ;
        RECT 6.16 10.079 8.56 10.081 ;
  LAYER M2 ;
        RECT 6.16 10.163 8.56 10.165 ;
  LAYER M2 ;
        RECT 6.16 10.247 8.56 10.249 ;
  LAYER M2 ;
        RECT 6.16 10.331 8.56 10.333 ;
  LAYER M2 ;
        RECT 6.16 10.415 8.56 10.417 ;
  LAYER M2 ;
        RECT 6.16 10.499 8.56 10.501 ;
  LAYER M2 ;
        RECT 6.16 10.5825 8.56 10.5845 ;
  LAYER M2 ;
        RECT 6.16 10.667 8.56 10.669 ;
  LAYER M2 ;
        RECT 6.16 10.751 8.56 10.753 ;
  LAYER M2 ;
        RECT 6.16 10.835 8.56 10.837 ;
  LAYER M2 ;
        RECT 6.16 10.919 8.56 10.921 ;
  LAYER M2 ;
        RECT 6.16 11.003 8.56 11.005 ;
  LAYER M2 ;
        RECT 6.16 11.087 8.56 11.089 ;
  LAYER M2 ;
        RECT 6.16 11.171 8.56 11.173 ;
  LAYER M2 ;
        RECT 6.16 11.255 8.56 11.257 ;
  LAYER M2 ;
        RECT 6.16 11.339 8.56 11.341 ;
  LAYER M2 ;
        RECT 6.16 11.423 8.56 11.425 ;
  LAYER M2 ;
        RECT 6.16 11.507 8.56 11.509 ;
  LAYER M2 ;
        RECT 6.16 11.591 8.56 11.593 ;
  LAYER M2 ;
        RECT 6.16 11.675 8.56 11.677 ;
  LAYER M2 ;
        RECT 6.16 11.759 8.56 11.761 ;
  LAYER M2 ;
        RECT 6.16 11.843 8.56 11.845 ;
  LAYER M2 ;
        RECT 6.16 11.927 8.56 11.929 ;
  LAYER M1 ;
        RECT 6.144 12.48 6.176 14.988 ;
  LAYER M1 ;
        RECT 6.208 12.48 6.24 14.988 ;
  LAYER M1 ;
        RECT 6.272 12.48 6.304 14.988 ;
  LAYER M1 ;
        RECT 6.336 12.48 6.368 14.988 ;
  LAYER M1 ;
        RECT 6.4 12.48 6.432 14.988 ;
  LAYER M1 ;
        RECT 6.464 12.48 6.496 14.988 ;
  LAYER M1 ;
        RECT 6.528 12.48 6.56 14.988 ;
  LAYER M1 ;
        RECT 6.592 12.48 6.624 14.988 ;
  LAYER M1 ;
        RECT 6.656 12.48 6.688 14.988 ;
  LAYER M1 ;
        RECT 6.72 12.48 6.752 14.988 ;
  LAYER M1 ;
        RECT 6.784 12.48 6.816 14.988 ;
  LAYER M1 ;
        RECT 6.848 12.48 6.88 14.988 ;
  LAYER M1 ;
        RECT 6.912 12.48 6.944 14.988 ;
  LAYER M1 ;
        RECT 6.976 12.48 7.008 14.988 ;
  LAYER M1 ;
        RECT 7.04 12.48 7.072 14.988 ;
  LAYER M1 ;
        RECT 7.104 12.48 7.136 14.988 ;
  LAYER M1 ;
        RECT 7.168 12.48 7.2 14.988 ;
  LAYER M1 ;
        RECT 7.232 12.48 7.264 14.988 ;
  LAYER M1 ;
        RECT 7.296 12.48 7.328 14.988 ;
  LAYER M1 ;
        RECT 7.36 12.48 7.392 14.988 ;
  LAYER M1 ;
        RECT 7.424 12.48 7.456 14.988 ;
  LAYER M1 ;
        RECT 7.488 12.48 7.52 14.988 ;
  LAYER M1 ;
        RECT 7.552 12.48 7.584 14.988 ;
  LAYER M1 ;
        RECT 7.616 12.48 7.648 14.988 ;
  LAYER M1 ;
        RECT 7.68 12.48 7.712 14.988 ;
  LAYER M1 ;
        RECT 7.744 12.48 7.776 14.988 ;
  LAYER M1 ;
        RECT 7.808 12.48 7.84 14.988 ;
  LAYER M1 ;
        RECT 7.872 12.48 7.904 14.988 ;
  LAYER M1 ;
        RECT 7.936 12.48 7.968 14.988 ;
  LAYER M1 ;
        RECT 8 12.48 8.032 14.988 ;
  LAYER M1 ;
        RECT 8.064 12.48 8.096 14.988 ;
  LAYER M1 ;
        RECT 8.128 12.48 8.16 14.988 ;
  LAYER M1 ;
        RECT 8.192 12.48 8.224 14.988 ;
  LAYER M1 ;
        RECT 8.256 12.48 8.288 14.988 ;
  LAYER M1 ;
        RECT 8.32 12.48 8.352 14.988 ;
  LAYER M1 ;
        RECT 8.384 12.48 8.416 14.988 ;
  LAYER M1 ;
        RECT 8.448 12.48 8.48 14.988 ;
  LAYER M2 ;
        RECT 6.124 12.564 8.596 12.596 ;
  LAYER M2 ;
        RECT 6.124 12.628 8.596 12.66 ;
  LAYER M2 ;
        RECT 6.124 12.692 8.596 12.724 ;
  LAYER M2 ;
        RECT 6.124 12.756 8.596 12.788 ;
  LAYER M2 ;
        RECT 6.124 12.82 8.596 12.852 ;
  LAYER M2 ;
        RECT 6.124 12.884 8.596 12.916 ;
  LAYER M2 ;
        RECT 6.124 12.948 8.596 12.98 ;
  LAYER M2 ;
        RECT 6.124 13.012 8.596 13.044 ;
  LAYER M2 ;
        RECT 6.124 13.076 8.596 13.108 ;
  LAYER M2 ;
        RECT 6.124 13.14 8.596 13.172 ;
  LAYER M2 ;
        RECT 6.124 13.204 8.596 13.236 ;
  LAYER M2 ;
        RECT 6.124 13.268 8.596 13.3 ;
  LAYER M2 ;
        RECT 6.124 13.332 8.596 13.364 ;
  LAYER M2 ;
        RECT 6.124 13.396 8.596 13.428 ;
  LAYER M2 ;
        RECT 6.124 13.46 8.596 13.492 ;
  LAYER M2 ;
        RECT 6.124 13.524 8.596 13.556 ;
  LAYER M2 ;
        RECT 6.124 13.588 8.596 13.62 ;
  LAYER M2 ;
        RECT 6.124 13.652 8.596 13.684 ;
  LAYER M2 ;
        RECT 6.124 13.716 8.596 13.748 ;
  LAYER M2 ;
        RECT 6.124 13.78 8.596 13.812 ;
  LAYER M2 ;
        RECT 6.124 13.844 8.596 13.876 ;
  LAYER M2 ;
        RECT 6.124 13.908 8.596 13.94 ;
  LAYER M2 ;
        RECT 6.124 13.972 8.596 14.004 ;
  LAYER M2 ;
        RECT 6.124 14.036 8.596 14.068 ;
  LAYER M2 ;
        RECT 6.124 14.1 8.596 14.132 ;
  LAYER M2 ;
        RECT 6.124 14.164 8.596 14.196 ;
  LAYER M2 ;
        RECT 6.124 14.228 8.596 14.26 ;
  LAYER M2 ;
        RECT 6.124 14.292 8.596 14.324 ;
  LAYER M2 ;
        RECT 6.124 14.356 8.596 14.388 ;
  LAYER M2 ;
        RECT 6.124 14.42 8.596 14.452 ;
  LAYER M2 ;
        RECT 6.124 14.484 8.596 14.516 ;
  LAYER M2 ;
        RECT 6.124 14.548 8.596 14.58 ;
  LAYER M2 ;
        RECT 6.124 14.612 8.596 14.644 ;
  LAYER M2 ;
        RECT 6.124 14.676 8.596 14.708 ;
  LAYER M2 ;
        RECT 6.124 14.74 8.596 14.772 ;
  LAYER M2 ;
        RECT 6.124 14.804 8.596 14.836 ;
  LAYER M3 ;
        RECT 6.144 12.48 6.176 14.988 ;
  LAYER M3 ;
        RECT 6.208 12.48 6.24 14.988 ;
  LAYER M3 ;
        RECT 6.272 12.48 6.304 14.988 ;
  LAYER M3 ;
        RECT 6.336 12.48 6.368 14.988 ;
  LAYER M3 ;
        RECT 6.4 12.48 6.432 14.988 ;
  LAYER M3 ;
        RECT 6.464 12.48 6.496 14.988 ;
  LAYER M3 ;
        RECT 6.528 12.48 6.56 14.988 ;
  LAYER M3 ;
        RECT 6.592 12.48 6.624 14.988 ;
  LAYER M3 ;
        RECT 6.656 12.48 6.688 14.988 ;
  LAYER M3 ;
        RECT 6.72 12.48 6.752 14.988 ;
  LAYER M3 ;
        RECT 6.784 12.48 6.816 14.988 ;
  LAYER M3 ;
        RECT 6.848 12.48 6.88 14.988 ;
  LAYER M3 ;
        RECT 6.912 12.48 6.944 14.988 ;
  LAYER M3 ;
        RECT 6.976 12.48 7.008 14.988 ;
  LAYER M3 ;
        RECT 7.04 12.48 7.072 14.988 ;
  LAYER M3 ;
        RECT 7.104 12.48 7.136 14.988 ;
  LAYER M3 ;
        RECT 7.168 12.48 7.2 14.988 ;
  LAYER M3 ;
        RECT 7.232 12.48 7.264 14.988 ;
  LAYER M3 ;
        RECT 7.296 12.48 7.328 14.988 ;
  LAYER M3 ;
        RECT 7.36 12.48 7.392 14.988 ;
  LAYER M3 ;
        RECT 7.424 12.48 7.456 14.988 ;
  LAYER M3 ;
        RECT 7.488 12.48 7.52 14.988 ;
  LAYER M3 ;
        RECT 7.552 12.48 7.584 14.988 ;
  LAYER M3 ;
        RECT 7.616 12.48 7.648 14.988 ;
  LAYER M3 ;
        RECT 7.68 12.48 7.712 14.988 ;
  LAYER M3 ;
        RECT 7.744 12.48 7.776 14.988 ;
  LAYER M3 ;
        RECT 7.808 12.48 7.84 14.988 ;
  LAYER M3 ;
        RECT 7.872 12.48 7.904 14.988 ;
  LAYER M3 ;
        RECT 7.936 12.48 7.968 14.988 ;
  LAYER M3 ;
        RECT 8 12.48 8.032 14.988 ;
  LAYER M3 ;
        RECT 8.064 12.48 8.096 14.988 ;
  LAYER M3 ;
        RECT 8.128 12.48 8.16 14.988 ;
  LAYER M3 ;
        RECT 8.192 12.48 8.224 14.988 ;
  LAYER M3 ;
        RECT 8.256 12.48 8.288 14.988 ;
  LAYER M3 ;
        RECT 8.32 12.48 8.352 14.988 ;
  LAYER M3 ;
        RECT 8.384 12.48 8.416 14.988 ;
  LAYER M3 ;
        RECT 8.448 12.48 8.48 14.988 ;
  LAYER M3 ;
        RECT 8.544 12.48 8.576 14.988 ;
  LAYER M1 ;
        RECT 6.159 12.516 6.161 14.952 ;
  LAYER M1 ;
        RECT 6.239 12.516 6.241 14.952 ;
  LAYER M1 ;
        RECT 6.319 12.516 6.321 14.952 ;
  LAYER M1 ;
        RECT 6.399 12.516 6.401 14.952 ;
  LAYER M1 ;
        RECT 6.479 12.516 6.481 14.952 ;
  LAYER M1 ;
        RECT 6.559 12.516 6.561 14.952 ;
  LAYER M1 ;
        RECT 6.639 12.516 6.641 14.952 ;
  LAYER M1 ;
        RECT 6.719 12.516 6.721 14.952 ;
  LAYER M1 ;
        RECT 6.799 12.516 6.801 14.952 ;
  LAYER M1 ;
        RECT 6.879 12.516 6.881 14.952 ;
  LAYER M1 ;
        RECT 6.959 12.516 6.961 14.952 ;
  LAYER M1 ;
        RECT 7.039 12.516 7.041 14.952 ;
  LAYER M1 ;
        RECT 7.119 12.516 7.121 14.952 ;
  LAYER M1 ;
        RECT 7.199 12.516 7.201 14.952 ;
  LAYER M1 ;
        RECT 7.279 12.516 7.281 14.952 ;
  LAYER M1 ;
        RECT 7.359 12.516 7.361 14.952 ;
  LAYER M1 ;
        RECT 7.439 12.516 7.441 14.952 ;
  LAYER M1 ;
        RECT 7.519 12.516 7.521 14.952 ;
  LAYER M1 ;
        RECT 7.599 12.516 7.601 14.952 ;
  LAYER M1 ;
        RECT 7.679 12.516 7.681 14.952 ;
  LAYER M1 ;
        RECT 7.759 12.516 7.761 14.952 ;
  LAYER M1 ;
        RECT 7.839 12.516 7.841 14.952 ;
  LAYER M1 ;
        RECT 7.919 12.516 7.921 14.952 ;
  LAYER M1 ;
        RECT 7.999 12.516 8.001 14.952 ;
  LAYER M1 ;
        RECT 8.079 12.516 8.081 14.952 ;
  LAYER M1 ;
        RECT 8.159 12.516 8.161 14.952 ;
  LAYER M1 ;
        RECT 8.239 12.516 8.241 14.952 ;
  LAYER M1 ;
        RECT 8.319 12.516 8.321 14.952 ;
  LAYER M1 ;
        RECT 8.399 12.516 8.401 14.952 ;
  LAYER M1 ;
        RECT 8.479 12.516 8.481 14.952 ;
  LAYER M2 ;
        RECT 6.16 12.515 8.56 12.517 ;
  LAYER M2 ;
        RECT 6.16 12.599 8.56 12.601 ;
  LAYER M2 ;
        RECT 6.16 12.683 8.56 12.685 ;
  LAYER M2 ;
        RECT 6.16 12.767 8.56 12.769 ;
  LAYER M2 ;
        RECT 6.16 12.851 8.56 12.853 ;
  LAYER M2 ;
        RECT 6.16 12.935 8.56 12.937 ;
  LAYER M2 ;
        RECT 6.16 13.019 8.56 13.021 ;
  LAYER M2 ;
        RECT 6.16 13.103 8.56 13.105 ;
  LAYER M2 ;
        RECT 6.16 13.187 8.56 13.189 ;
  LAYER M2 ;
        RECT 6.16 13.271 8.56 13.273 ;
  LAYER M2 ;
        RECT 6.16 13.355 8.56 13.357 ;
  LAYER M2 ;
        RECT 6.16 13.439 8.56 13.441 ;
  LAYER M2 ;
        RECT 6.16 13.5225 8.56 13.5245 ;
  LAYER M2 ;
        RECT 6.16 13.607 8.56 13.609 ;
  LAYER M2 ;
        RECT 6.16 13.691 8.56 13.693 ;
  LAYER M2 ;
        RECT 6.16 13.775 8.56 13.777 ;
  LAYER M2 ;
        RECT 6.16 13.859 8.56 13.861 ;
  LAYER M2 ;
        RECT 6.16 13.943 8.56 13.945 ;
  LAYER M2 ;
        RECT 6.16 14.027 8.56 14.029 ;
  LAYER M2 ;
        RECT 6.16 14.111 8.56 14.113 ;
  LAYER M2 ;
        RECT 6.16 14.195 8.56 14.197 ;
  LAYER M2 ;
        RECT 6.16 14.279 8.56 14.281 ;
  LAYER M2 ;
        RECT 6.16 14.363 8.56 14.365 ;
  LAYER M2 ;
        RECT 6.16 14.447 8.56 14.449 ;
  LAYER M2 ;
        RECT 6.16 14.531 8.56 14.533 ;
  LAYER M2 ;
        RECT 6.16 14.615 8.56 14.617 ;
  LAYER M2 ;
        RECT 6.16 14.699 8.56 14.701 ;
  LAYER M2 ;
        RECT 6.16 14.783 8.56 14.785 ;
  LAYER M2 ;
        RECT 6.16 14.867 8.56 14.869 ;
  LAYER M1 ;
        RECT 6.144 15.42 6.176 17.928 ;
  LAYER M1 ;
        RECT 6.208 15.42 6.24 17.928 ;
  LAYER M1 ;
        RECT 6.272 15.42 6.304 17.928 ;
  LAYER M1 ;
        RECT 6.336 15.42 6.368 17.928 ;
  LAYER M1 ;
        RECT 6.4 15.42 6.432 17.928 ;
  LAYER M1 ;
        RECT 6.464 15.42 6.496 17.928 ;
  LAYER M1 ;
        RECT 6.528 15.42 6.56 17.928 ;
  LAYER M1 ;
        RECT 6.592 15.42 6.624 17.928 ;
  LAYER M1 ;
        RECT 6.656 15.42 6.688 17.928 ;
  LAYER M1 ;
        RECT 6.72 15.42 6.752 17.928 ;
  LAYER M1 ;
        RECT 6.784 15.42 6.816 17.928 ;
  LAYER M1 ;
        RECT 6.848 15.42 6.88 17.928 ;
  LAYER M1 ;
        RECT 6.912 15.42 6.944 17.928 ;
  LAYER M1 ;
        RECT 6.976 15.42 7.008 17.928 ;
  LAYER M1 ;
        RECT 7.04 15.42 7.072 17.928 ;
  LAYER M1 ;
        RECT 7.104 15.42 7.136 17.928 ;
  LAYER M1 ;
        RECT 7.168 15.42 7.2 17.928 ;
  LAYER M1 ;
        RECT 7.232 15.42 7.264 17.928 ;
  LAYER M1 ;
        RECT 7.296 15.42 7.328 17.928 ;
  LAYER M1 ;
        RECT 7.36 15.42 7.392 17.928 ;
  LAYER M1 ;
        RECT 7.424 15.42 7.456 17.928 ;
  LAYER M1 ;
        RECT 7.488 15.42 7.52 17.928 ;
  LAYER M1 ;
        RECT 7.552 15.42 7.584 17.928 ;
  LAYER M1 ;
        RECT 7.616 15.42 7.648 17.928 ;
  LAYER M1 ;
        RECT 7.68 15.42 7.712 17.928 ;
  LAYER M1 ;
        RECT 7.744 15.42 7.776 17.928 ;
  LAYER M1 ;
        RECT 7.808 15.42 7.84 17.928 ;
  LAYER M1 ;
        RECT 7.872 15.42 7.904 17.928 ;
  LAYER M1 ;
        RECT 7.936 15.42 7.968 17.928 ;
  LAYER M1 ;
        RECT 8 15.42 8.032 17.928 ;
  LAYER M1 ;
        RECT 8.064 15.42 8.096 17.928 ;
  LAYER M1 ;
        RECT 8.128 15.42 8.16 17.928 ;
  LAYER M1 ;
        RECT 8.192 15.42 8.224 17.928 ;
  LAYER M1 ;
        RECT 8.256 15.42 8.288 17.928 ;
  LAYER M1 ;
        RECT 8.32 15.42 8.352 17.928 ;
  LAYER M1 ;
        RECT 8.384 15.42 8.416 17.928 ;
  LAYER M1 ;
        RECT 8.448 15.42 8.48 17.928 ;
  LAYER M2 ;
        RECT 6.124 15.504 8.596 15.536 ;
  LAYER M2 ;
        RECT 6.124 15.568 8.596 15.6 ;
  LAYER M2 ;
        RECT 6.124 15.632 8.596 15.664 ;
  LAYER M2 ;
        RECT 6.124 15.696 8.596 15.728 ;
  LAYER M2 ;
        RECT 6.124 15.76 8.596 15.792 ;
  LAYER M2 ;
        RECT 6.124 15.824 8.596 15.856 ;
  LAYER M2 ;
        RECT 6.124 15.888 8.596 15.92 ;
  LAYER M2 ;
        RECT 6.124 15.952 8.596 15.984 ;
  LAYER M2 ;
        RECT 6.124 16.016 8.596 16.048 ;
  LAYER M2 ;
        RECT 6.124 16.08 8.596 16.112 ;
  LAYER M2 ;
        RECT 6.124 16.144 8.596 16.176 ;
  LAYER M2 ;
        RECT 6.124 16.208 8.596 16.24 ;
  LAYER M2 ;
        RECT 6.124 16.272 8.596 16.304 ;
  LAYER M2 ;
        RECT 6.124 16.336 8.596 16.368 ;
  LAYER M2 ;
        RECT 6.124 16.4 8.596 16.432 ;
  LAYER M2 ;
        RECT 6.124 16.464 8.596 16.496 ;
  LAYER M2 ;
        RECT 6.124 16.528 8.596 16.56 ;
  LAYER M2 ;
        RECT 6.124 16.592 8.596 16.624 ;
  LAYER M2 ;
        RECT 6.124 16.656 8.596 16.688 ;
  LAYER M2 ;
        RECT 6.124 16.72 8.596 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.784 8.596 16.816 ;
  LAYER M2 ;
        RECT 6.124 16.848 8.596 16.88 ;
  LAYER M2 ;
        RECT 6.124 16.912 8.596 16.944 ;
  LAYER M2 ;
        RECT 6.124 16.976 8.596 17.008 ;
  LAYER M2 ;
        RECT 6.124 17.04 8.596 17.072 ;
  LAYER M2 ;
        RECT 6.124 17.104 8.596 17.136 ;
  LAYER M2 ;
        RECT 6.124 17.168 8.596 17.2 ;
  LAYER M2 ;
        RECT 6.124 17.232 8.596 17.264 ;
  LAYER M2 ;
        RECT 6.124 17.296 8.596 17.328 ;
  LAYER M2 ;
        RECT 6.124 17.36 8.596 17.392 ;
  LAYER M2 ;
        RECT 6.124 17.424 8.596 17.456 ;
  LAYER M2 ;
        RECT 6.124 17.488 8.596 17.52 ;
  LAYER M2 ;
        RECT 6.124 17.552 8.596 17.584 ;
  LAYER M2 ;
        RECT 6.124 17.616 8.596 17.648 ;
  LAYER M2 ;
        RECT 6.124 17.68 8.596 17.712 ;
  LAYER M2 ;
        RECT 6.124 17.744 8.596 17.776 ;
  LAYER M3 ;
        RECT 6.144 15.42 6.176 17.928 ;
  LAYER M3 ;
        RECT 6.208 15.42 6.24 17.928 ;
  LAYER M3 ;
        RECT 6.272 15.42 6.304 17.928 ;
  LAYER M3 ;
        RECT 6.336 15.42 6.368 17.928 ;
  LAYER M3 ;
        RECT 6.4 15.42 6.432 17.928 ;
  LAYER M3 ;
        RECT 6.464 15.42 6.496 17.928 ;
  LAYER M3 ;
        RECT 6.528 15.42 6.56 17.928 ;
  LAYER M3 ;
        RECT 6.592 15.42 6.624 17.928 ;
  LAYER M3 ;
        RECT 6.656 15.42 6.688 17.928 ;
  LAYER M3 ;
        RECT 6.72 15.42 6.752 17.928 ;
  LAYER M3 ;
        RECT 6.784 15.42 6.816 17.928 ;
  LAYER M3 ;
        RECT 6.848 15.42 6.88 17.928 ;
  LAYER M3 ;
        RECT 6.912 15.42 6.944 17.928 ;
  LAYER M3 ;
        RECT 6.976 15.42 7.008 17.928 ;
  LAYER M3 ;
        RECT 7.04 15.42 7.072 17.928 ;
  LAYER M3 ;
        RECT 7.104 15.42 7.136 17.928 ;
  LAYER M3 ;
        RECT 7.168 15.42 7.2 17.928 ;
  LAYER M3 ;
        RECT 7.232 15.42 7.264 17.928 ;
  LAYER M3 ;
        RECT 7.296 15.42 7.328 17.928 ;
  LAYER M3 ;
        RECT 7.36 15.42 7.392 17.928 ;
  LAYER M3 ;
        RECT 7.424 15.42 7.456 17.928 ;
  LAYER M3 ;
        RECT 7.488 15.42 7.52 17.928 ;
  LAYER M3 ;
        RECT 7.552 15.42 7.584 17.928 ;
  LAYER M3 ;
        RECT 7.616 15.42 7.648 17.928 ;
  LAYER M3 ;
        RECT 7.68 15.42 7.712 17.928 ;
  LAYER M3 ;
        RECT 7.744 15.42 7.776 17.928 ;
  LAYER M3 ;
        RECT 7.808 15.42 7.84 17.928 ;
  LAYER M3 ;
        RECT 7.872 15.42 7.904 17.928 ;
  LAYER M3 ;
        RECT 7.936 15.42 7.968 17.928 ;
  LAYER M3 ;
        RECT 8 15.42 8.032 17.928 ;
  LAYER M3 ;
        RECT 8.064 15.42 8.096 17.928 ;
  LAYER M3 ;
        RECT 8.128 15.42 8.16 17.928 ;
  LAYER M3 ;
        RECT 8.192 15.42 8.224 17.928 ;
  LAYER M3 ;
        RECT 8.256 15.42 8.288 17.928 ;
  LAYER M3 ;
        RECT 8.32 15.42 8.352 17.928 ;
  LAYER M3 ;
        RECT 8.384 15.42 8.416 17.928 ;
  LAYER M3 ;
        RECT 8.448 15.42 8.48 17.928 ;
  LAYER M3 ;
        RECT 8.544 15.42 8.576 17.928 ;
  LAYER M1 ;
        RECT 6.159 15.456 6.161 17.892 ;
  LAYER M1 ;
        RECT 6.239 15.456 6.241 17.892 ;
  LAYER M1 ;
        RECT 6.319 15.456 6.321 17.892 ;
  LAYER M1 ;
        RECT 6.399 15.456 6.401 17.892 ;
  LAYER M1 ;
        RECT 6.479 15.456 6.481 17.892 ;
  LAYER M1 ;
        RECT 6.559 15.456 6.561 17.892 ;
  LAYER M1 ;
        RECT 6.639 15.456 6.641 17.892 ;
  LAYER M1 ;
        RECT 6.719 15.456 6.721 17.892 ;
  LAYER M1 ;
        RECT 6.799 15.456 6.801 17.892 ;
  LAYER M1 ;
        RECT 6.879 15.456 6.881 17.892 ;
  LAYER M1 ;
        RECT 6.959 15.456 6.961 17.892 ;
  LAYER M1 ;
        RECT 7.039 15.456 7.041 17.892 ;
  LAYER M1 ;
        RECT 7.119 15.456 7.121 17.892 ;
  LAYER M1 ;
        RECT 7.199 15.456 7.201 17.892 ;
  LAYER M1 ;
        RECT 7.279 15.456 7.281 17.892 ;
  LAYER M1 ;
        RECT 7.359 15.456 7.361 17.892 ;
  LAYER M1 ;
        RECT 7.439 15.456 7.441 17.892 ;
  LAYER M1 ;
        RECT 7.519 15.456 7.521 17.892 ;
  LAYER M1 ;
        RECT 7.599 15.456 7.601 17.892 ;
  LAYER M1 ;
        RECT 7.679 15.456 7.681 17.892 ;
  LAYER M1 ;
        RECT 7.759 15.456 7.761 17.892 ;
  LAYER M1 ;
        RECT 7.839 15.456 7.841 17.892 ;
  LAYER M1 ;
        RECT 7.919 15.456 7.921 17.892 ;
  LAYER M1 ;
        RECT 7.999 15.456 8.001 17.892 ;
  LAYER M1 ;
        RECT 8.079 15.456 8.081 17.892 ;
  LAYER M1 ;
        RECT 8.159 15.456 8.161 17.892 ;
  LAYER M1 ;
        RECT 8.239 15.456 8.241 17.892 ;
  LAYER M1 ;
        RECT 8.319 15.456 8.321 17.892 ;
  LAYER M1 ;
        RECT 8.399 15.456 8.401 17.892 ;
  LAYER M1 ;
        RECT 8.479 15.456 8.481 17.892 ;
  LAYER M2 ;
        RECT 6.16 15.455 8.56 15.457 ;
  LAYER M2 ;
        RECT 6.16 15.539 8.56 15.541 ;
  LAYER M2 ;
        RECT 6.16 15.623 8.56 15.625 ;
  LAYER M2 ;
        RECT 6.16 15.707 8.56 15.709 ;
  LAYER M2 ;
        RECT 6.16 15.791 8.56 15.793 ;
  LAYER M2 ;
        RECT 6.16 15.875 8.56 15.877 ;
  LAYER M2 ;
        RECT 6.16 15.959 8.56 15.961 ;
  LAYER M2 ;
        RECT 6.16 16.043 8.56 16.045 ;
  LAYER M2 ;
        RECT 6.16 16.127 8.56 16.129 ;
  LAYER M2 ;
        RECT 6.16 16.211 8.56 16.213 ;
  LAYER M2 ;
        RECT 6.16 16.295 8.56 16.297 ;
  LAYER M2 ;
        RECT 6.16 16.379 8.56 16.381 ;
  LAYER M2 ;
        RECT 6.16 16.4625 8.56 16.4645 ;
  LAYER M2 ;
        RECT 6.16 16.547 8.56 16.549 ;
  LAYER M2 ;
        RECT 6.16 16.631 8.56 16.633 ;
  LAYER M2 ;
        RECT 6.16 16.715 8.56 16.717 ;
  LAYER M2 ;
        RECT 6.16 16.799 8.56 16.801 ;
  LAYER M2 ;
        RECT 6.16 16.883 8.56 16.885 ;
  LAYER M2 ;
        RECT 6.16 16.967 8.56 16.969 ;
  LAYER M2 ;
        RECT 6.16 17.051 8.56 17.053 ;
  LAYER M2 ;
        RECT 6.16 17.135 8.56 17.137 ;
  LAYER M2 ;
        RECT 6.16 17.219 8.56 17.221 ;
  LAYER M2 ;
        RECT 6.16 17.303 8.56 17.305 ;
  LAYER M2 ;
        RECT 6.16 17.387 8.56 17.389 ;
  LAYER M2 ;
        RECT 6.16 17.471 8.56 17.473 ;
  LAYER M2 ;
        RECT 6.16 17.555 8.56 17.557 ;
  LAYER M2 ;
        RECT 6.16 17.639 8.56 17.641 ;
  LAYER M2 ;
        RECT 6.16 17.723 8.56 17.725 ;
  LAYER M2 ;
        RECT 6.16 17.807 8.56 17.809 ;
  LAYER M1 ;
        RECT 6.144 18.36 6.176 20.868 ;
  LAYER M1 ;
        RECT 6.208 18.36 6.24 20.868 ;
  LAYER M1 ;
        RECT 6.272 18.36 6.304 20.868 ;
  LAYER M1 ;
        RECT 6.336 18.36 6.368 20.868 ;
  LAYER M1 ;
        RECT 6.4 18.36 6.432 20.868 ;
  LAYER M1 ;
        RECT 6.464 18.36 6.496 20.868 ;
  LAYER M1 ;
        RECT 6.528 18.36 6.56 20.868 ;
  LAYER M1 ;
        RECT 6.592 18.36 6.624 20.868 ;
  LAYER M1 ;
        RECT 6.656 18.36 6.688 20.868 ;
  LAYER M1 ;
        RECT 6.72 18.36 6.752 20.868 ;
  LAYER M1 ;
        RECT 6.784 18.36 6.816 20.868 ;
  LAYER M1 ;
        RECT 6.848 18.36 6.88 20.868 ;
  LAYER M1 ;
        RECT 6.912 18.36 6.944 20.868 ;
  LAYER M1 ;
        RECT 6.976 18.36 7.008 20.868 ;
  LAYER M1 ;
        RECT 7.04 18.36 7.072 20.868 ;
  LAYER M1 ;
        RECT 7.104 18.36 7.136 20.868 ;
  LAYER M1 ;
        RECT 7.168 18.36 7.2 20.868 ;
  LAYER M1 ;
        RECT 7.232 18.36 7.264 20.868 ;
  LAYER M1 ;
        RECT 7.296 18.36 7.328 20.868 ;
  LAYER M1 ;
        RECT 7.36 18.36 7.392 20.868 ;
  LAYER M1 ;
        RECT 7.424 18.36 7.456 20.868 ;
  LAYER M1 ;
        RECT 7.488 18.36 7.52 20.868 ;
  LAYER M1 ;
        RECT 7.552 18.36 7.584 20.868 ;
  LAYER M1 ;
        RECT 7.616 18.36 7.648 20.868 ;
  LAYER M1 ;
        RECT 7.68 18.36 7.712 20.868 ;
  LAYER M1 ;
        RECT 7.744 18.36 7.776 20.868 ;
  LAYER M1 ;
        RECT 7.808 18.36 7.84 20.868 ;
  LAYER M1 ;
        RECT 7.872 18.36 7.904 20.868 ;
  LAYER M1 ;
        RECT 7.936 18.36 7.968 20.868 ;
  LAYER M1 ;
        RECT 8 18.36 8.032 20.868 ;
  LAYER M1 ;
        RECT 8.064 18.36 8.096 20.868 ;
  LAYER M1 ;
        RECT 8.128 18.36 8.16 20.868 ;
  LAYER M1 ;
        RECT 8.192 18.36 8.224 20.868 ;
  LAYER M1 ;
        RECT 8.256 18.36 8.288 20.868 ;
  LAYER M1 ;
        RECT 8.32 18.36 8.352 20.868 ;
  LAYER M1 ;
        RECT 8.384 18.36 8.416 20.868 ;
  LAYER M1 ;
        RECT 8.448 18.36 8.48 20.868 ;
  LAYER M2 ;
        RECT 6.124 18.444 8.596 18.476 ;
  LAYER M2 ;
        RECT 6.124 18.508 8.596 18.54 ;
  LAYER M2 ;
        RECT 6.124 18.572 8.596 18.604 ;
  LAYER M2 ;
        RECT 6.124 18.636 8.596 18.668 ;
  LAYER M2 ;
        RECT 6.124 18.7 8.596 18.732 ;
  LAYER M2 ;
        RECT 6.124 18.764 8.596 18.796 ;
  LAYER M2 ;
        RECT 6.124 18.828 8.596 18.86 ;
  LAYER M2 ;
        RECT 6.124 18.892 8.596 18.924 ;
  LAYER M2 ;
        RECT 6.124 18.956 8.596 18.988 ;
  LAYER M2 ;
        RECT 6.124 19.02 8.596 19.052 ;
  LAYER M2 ;
        RECT 6.124 19.084 8.596 19.116 ;
  LAYER M2 ;
        RECT 6.124 19.148 8.596 19.18 ;
  LAYER M2 ;
        RECT 6.124 19.212 8.596 19.244 ;
  LAYER M2 ;
        RECT 6.124 19.276 8.596 19.308 ;
  LAYER M2 ;
        RECT 6.124 19.34 8.596 19.372 ;
  LAYER M2 ;
        RECT 6.124 19.404 8.596 19.436 ;
  LAYER M2 ;
        RECT 6.124 19.468 8.596 19.5 ;
  LAYER M2 ;
        RECT 6.124 19.532 8.596 19.564 ;
  LAYER M2 ;
        RECT 6.124 19.596 8.596 19.628 ;
  LAYER M2 ;
        RECT 6.124 19.66 8.596 19.692 ;
  LAYER M2 ;
        RECT 6.124 19.724 8.596 19.756 ;
  LAYER M2 ;
        RECT 6.124 19.788 8.596 19.82 ;
  LAYER M2 ;
        RECT 6.124 19.852 8.596 19.884 ;
  LAYER M2 ;
        RECT 6.124 19.916 8.596 19.948 ;
  LAYER M2 ;
        RECT 6.124 19.98 8.596 20.012 ;
  LAYER M2 ;
        RECT 6.124 20.044 8.596 20.076 ;
  LAYER M2 ;
        RECT 6.124 20.108 8.596 20.14 ;
  LAYER M2 ;
        RECT 6.124 20.172 8.596 20.204 ;
  LAYER M2 ;
        RECT 6.124 20.236 8.596 20.268 ;
  LAYER M2 ;
        RECT 6.124 20.3 8.596 20.332 ;
  LAYER M2 ;
        RECT 6.124 20.364 8.596 20.396 ;
  LAYER M2 ;
        RECT 6.124 20.428 8.596 20.46 ;
  LAYER M2 ;
        RECT 6.124 20.492 8.596 20.524 ;
  LAYER M2 ;
        RECT 6.124 20.556 8.596 20.588 ;
  LAYER M2 ;
        RECT 6.124 20.62 8.596 20.652 ;
  LAYER M2 ;
        RECT 6.124 20.684 8.596 20.716 ;
  LAYER M3 ;
        RECT 6.144 18.36 6.176 20.868 ;
  LAYER M3 ;
        RECT 6.208 18.36 6.24 20.868 ;
  LAYER M3 ;
        RECT 6.272 18.36 6.304 20.868 ;
  LAYER M3 ;
        RECT 6.336 18.36 6.368 20.868 ;
  LAYER M3 ;
        RECT 6.4 18.36 6.432 20.868 ;
  LAYER M3 ;
        RECT 6.464 18.36 6.496 20.868 ;
  LAYER M3 ;
        RECT 6.528 18.36 6.56 20.868 ;
  LAYER M3 ;
        RECT 6.592 18.36 6.624 20.868 ;
  LAYER M3 ;
        RECT 6.656 18.36 6.688 20.868 ;
  LAYER M3 ;
        RECT 6.72 18.36 6.752 20.868 ;
  LAYER M3 ;
        RECT 6.784 18.36 6.816 20.868 ;
  LAYER M3 ;
        RECT 6.848 18.36 6.88 20.868 ;
  LAYER M3 ;
        RECT 6.912 18.36 6.944 20.868 ;
  LAYER M3 ;
        RECT 6.976 18.36 7.008 20.868 ;
  LAYER M3 ;
        RECT 7.04 18.36 7.072 20.868 ;
  LAYER M3 ;
        RECT 7.104 18.36 7.136 20.868 ;
  LAYER M3 ;
        RECT 7.168 18.36 7.2 20.868 ;
  LAYER M3 ;
        RECT 7.232 18.36 7.264 20.868 ;
  LAYER M3 ;
        RECT 7.296 18.36 7.328 20.868 ;
  LAYER M3 ;
        RECT 7.36 18.36 7.392 20.868 ;
  LAYER M3 ;
        RECT 7.424 18.36 7.456 20.868 ;
  LAYER M3 ;
        RECT 7.488 18.36 7.52 20.868 ;
  LAYER M3 ;
        RECT 7.552 18.36 7.584 20.868 ;
  LAYER M3 ;
        RECT 7.616 18.36 7.648 20.868 ;
  LAYER M3 ;
        RECT 7.68 18.36 7.712 20.868 ;
  LAYER M3 ;
        RECT 7.744 18.36 7.776 20.868 ;
  LAYER M3 ;
        RECT 7.808 18.36 7.84 20.868 ;
  LAYER M3 ;
        RECT 7.872 18.36 7.904 20.868 ;
  LAYER M3 ;
        RECT 7.936 18.36 7.968 20.868 ;
  LAYER M3 ;
        RECT 8 18.36 8.032 20.868 ;
  LAYER M3 ;
        RECT 8.064 18.36 8.096 20.868 ;
  LAYER M3 ;
        RECT 8.128 18.36 8.16 20.868 ;
  LAYER M3 ;
        RECT 8.192 18.36 8.224 20.868 ;
  LAYER M3 ;
        RECT 8.256 18.36 8.288 20.868 ;
  LAYER M3 ;
        RECT 8.32 18.36 8.352 20.868 ;
  LAYER M3 ;
        RECT 8.384 18.36 8.416 20.868 ;
  LAYER M3 ;
        RECT 8.448 18.36 8.48 20.868 ;
  LAYER M3 ;
        RECT 8.544 18.36 8.576 20.868 ;
  LAYER M1 ;
        RECT 6.159 18.396 6.161 20.832 ;
  LAYER M1 ;
        RECT 6.239 18.396 6.241 20.832 ;
  LAYER M1 ;
        RECT 6.319 18.396 6.321 20.832 ;
  LAYER M1 ;
        RECT 6.399 18.396 6.401 20.832 ;
  LAYER M1 ;
        RECT 6.479 18.396 6.481 20.832 ;
  LAYER M1 ;
        RECT 6.559 18.396 6.561 20.832 ;
  LAYER M1 ;
        RECT 6.639 18.396 6.641 20.832 ;
  LAYER M1 ;
        RECT 6.719 18.396 6.721 20.832 ;
  LAYER M1 ;
        RECT 6.799 18.396 6.801 20.832 ;
  LAYER M1 ;
        RECT 6.879 18.396 6.881 20.832 ;
  LAYER M1 ;
        RECT 6.959 18.396 6.961 20.832 ;
  LAYER M1 ;
        RECT 7.039 18.396 7.041 20.832 ;
  LAYER M1 ;
        RECT 7.119 18.396 7.121 20.832 ;
  LAYER M1 ;
        RECT 7.199 18.396 7.201 20.832 ;
  LAYER M1 ;
        RECT 7.279 18.396 7.281 20.832 ;
  LAYER M1 ;
        RECT 7.359 18.396 7.361 20.832 ;
  LAYER M1 ;
        RECT 7.439 18.396 7.441 20.832 ;
  LAYER M1 ;
        RECT 7.519 18.396 7.521 20.832 ;
  LAYER M1 ;
        RECT 7.599 18.396 7.601 20.832 ;
  LAYER M1 ;
        RECT 7.679 18.396 7.681 20.832 ;
  LAYER M1 ;
        RECT 7.759 18.396 7.761 20.832 ;
  LAYER M1 ;
        RECT 7.839 18.396 7.841 20.832 ;
  LAYER M1 ;
        RECT 7.919 18.396 7.921 20.832 ;
  LAYER M1 ;
        RECT 7.999 18.396 8.001 20.832 ;
  LAYER M1 ;
        RECT 8.079 18.396 8.081 20.832 ;
  LAYER M1 ;
        RECT 8.159 18.396 8.161 20.832 ;
  LAYER M1 ;
        RECT 8.239 18.396 8.241 20.832 ;
  LAYER M1 ;
        RECT 8.319 18.396 8.321 20.832 ;
  LAYER M1 ;
        RECT 8.399 18.396 8.401 20.832 ;
  LAYER M1 ;
        RECT 8.479 18.396 8.481 20.832 ;
  LAYER M2 ;
        RECT 6.16 18.395 8.56 18.397 ;
  LAYER M2 ;
        RECT 6.16 18.479 8.56 18.481 ;
  LAYER M2 ;
        RECT 6.16 18.563 8.56 18.565 ;
  LAYER M2 ;
        RECT 6.16 18.647 8.56 18.649 ;
  LAYER M2 ;
        RECT 6.16 18.731 8.56 18.733 ;
  LAYER M2 ;
        RECT 6.16 18.815 8.56 18.817 ;
  LAYER M2 ;
        RECT 6.16 18.899 8.56 18.901 ;
  LAYER M2 ;
        RECT 6.16 18.983 8.56 18.985 ;
  LAYER M2 ;
        RECT 6.16 19.067 8.56 19.069 ;
  LAYER M2 ;
        RECT 6.16 19.151 8.56 19.153 ;
  LAYER M2 ;
        RECT 6.16 19.235 8.56 19.237 ;
  LAYER M2 ;
        RECT 6.16 19.319 8.56 19.321 ;
  LAYER M2 ;
        RECT 6.16 19.4025 8.56 19.4045 ;
  LAYER M2 ;
        RECT 6.16 19.487 8.56 19.489 ;
  LAYER M2 ;
        RECT 6.16 19.571 8.56 19.573 ;
  LAYER M2 ;
        RECT 6.16 19.655 8.56 19.657 ;
  LAYER M2 ;
        RECT 6.16 19.739 8.56 19.741 ;
  LAYER M2 ;
        RECT 6.16 19.823 8.56 19.825 ;
  LAYER M2 ;
        RECT 6.16 19.907 8.56 19.909 ;
  LAYER M2 ;
        RECT 6.16 19.991 8.56 19.993 ;
  LAYER M2 ;
        RECT 6.16 20.075 8.56 20.077 ;
  LAYER M2 ;
        RECT 6.16 20.159 8.56 20.161 ;
  LAYER M2 ;
        RECT 6.16 20.243 8.56 20.245 ;
  LAYER M2 ;
        RECT 6.16 20.327 8.56 20.329 ;
  LAYER M2 ;
        RECT 6.16 20.411 8.56 20.413 ;
  LAYER M2 ;
        RECT 6.16 20.495 8.56 20.497 ;
  LAYER M2 ;
        RECT 6.16 20.579 8.56 20.581 ;
  LAYER M2 ;
        RECT 6.16 20.663 8.56 20.665 ;
  LAYER M2 ;
        RECT 6.16 20.747 8.56 20.749 ;
  LAYER M1 ;
        RECT 6.144 21.3 6.176 23.808 ;
  LAYER M1 ;
        RECT 6.208 21.3 6.24 23.808 ;
  LAYER M1 ;
        RECT 6.272 21.3 6.304 23.808 ;
  LAYER M1 ;
        RECT 6.336 21.3 6.368 23.808 ;
  LAYER M1 ;
        RECT 6.4 21.3 6.432 23.808 ;
  LAYER M1 ;
        RECT 6.464 21.3 6.496 23.808 ;
  LAYER M1 ;
        RECT 6.528 21.3 6.56 23.808 ;
  LAYER M1 ;
        RECT 6.592 21.3 6.624 23.808 ;
  LAYER M1 ;
        RECT 6.656 21.3 6.688 23.808 ;
  LAYER M1 ;
        RECT 6.72 21.3 6.752 23.808 ;
  LAYER M1 ;
        RECT 6.784 21.3 6.816 23.808 ;
  LAYER M1 ;
        RECT 6.848 21.3 6.88 23.808 ;
  LAYER M1 ;
        RECT 6.912 21.3 6.944 23.808 ;
  LAYER M1 ;
        RECT 6.976 21.3 7.008 23.808 ;
  LAYER M1 ;
        RECT 7.04 21.3 7.072 23.808 ;
  LAYER M1 ;
        RECT 7.104 21.3 7.136 23.808 ;
  LAYER M1 ;
        RECT 7.168 21.3 7.2 23.808 ;
  LAYER M1 ;
        RECT 7.232 21.3 7.264 23.808 ;
  LAYER M1 ;
        RECT 7.296 21.3 7.328 23.808 ;
  LAYER M1 ;
        RECT 7.36 21.3 7.392 23.808 ;
  LAYER M1 ;
        RECT 7.424 21.3 7.456 23.808 ;
  LAYER M1 ;
        RECT 7.488 21.3 7.52 23.808 ;
  LAYER M1 ;
        RECT 7.552 21.3 7.584 23.808 ;
  LAYER M1 ;
        RECT 7.616 21.3 7.648 23.808 ;
  LAYER M1 ;
        RECT 7.68 21.3 7.712 23.808 ;
  LAYER M1 ;
        RECT 7.744 21.3 7.776 23.808 ;
  LAYER M1 ;
        RECT 7.808 21.3 7.84 23.808 ;
  LAYER M1 ;
        RECT 7.872 21.3 7.904 23.808 ;
  LAYER M1 ;
        RECT 7.936 21.3 7.968 23.808 ;
  LAYER M1 ;
        RECT 8 21.3 8.032 23.808 ;
  LAYER M1 ;
        RECT 8.064 21.3 8.096 23.808 ;
  LAYER M1 ;
        RECT 8.128 21.3 8.16 23.808 ;
  LAYER M1 ;
        RECT 8.192 21.3 8.224 23.808 ;
  LAYER M1 ;
        RECT 8.256 21.3 8.288 23.808 ;
  LAYER M1 ;
        RECT 8.32 21.3 8.352 23.808 ;
  LAYER M1 ;
        RECT 8.384 21.3 8.416 23.808 ;
  LAYER M1 ;
        RECT 8.448 21.3 8.48 23.808 ;
  LAYER M2 ;
        RECT 6.124 21.384 8.596 21.416 ;
  LAYER M2 ;
        RECT 6.124 21.448 8.596 21.48 ;
  LAYER M2 ;
        RECT 6.124 21.512 8.596 21.544 ;
  LAYER M2 ;
        RECT 6.124 21.576 8.596 21.608 ;
  LAYER M2 ;
        RECT 6.124 21.64 8.596 21.672 ;
  LAYER M2 ;
        RECT 6.124 21.704 8.596 21.736 ;
  LAYER M2 ;
        RECT 6.124 21.768 8.596 21.8 ;
  LAYER M2 ;
        RECT 6.124 21.832 8.596 21.864 ;
  LAYER M2 ;
        RECT 6.124 21.896 8.596 21.928 ;
  LAYER M2 ;
        RECT 6.124 21.96 8.596 21.992 ;
  LAYER M2 ;
        RECT 6.124 22.024 8.596 22.056 ;
  LAYER M2 ;
        RECT 6.124 22.088 8.596 22.12 ;
  LAYER M2 ;
        RECT 6.124 22.152 8.596 22.184 ;
  LAYER M2 ;
        RECT 6.124 22.216 8.596 22.248 ;
  LAYER M2 ;
        RECT 6.124 22.28 8.596 22.312 ;
  LAYER M2 ;
        RECT 6.124 22.344 8.596 22.376 ;
  LAYER M2 ;
        RECT 6.124 22.408 8.596 22.44 ;
  LAYER M2 ;
        RECT 6.124 22.472 8.596 22.504 ;
  LAYER M2 ;
        RECT 6.124 22.536 8.596 22.568 ;
  LAYER M2 ;
        RECT 6.124 22.6 8.596 22.632 ;
  LAYER M2 ;
        RECT 6.124 22.664 8.596 22.696 ;
  LAYER M2 ;
        RECT 6.124 22.728 8.596 22.76 ;
  LAYER M2 ;
        RECT 6.124 22.792 8.596 22.824 ;
  LAYER M2 ;
        RECT 6.124 22.856 8.596 22.888 ;
  LAYER M2 ;
        RECT 6.124 22.92 8.596 22.952 ;
  LAYER M2 ;
        RECT 6.124 22.984 8.596 23.016 ;
  LAYER M2 ;
        RECT 6.124 23.048 8.596 23.08 ;
  LAYER M2 ;
        RECT 6.124 23.112 8.596 23.144 ;
  LAYER M2 ;
        RECT 6.124 23.176 8.596 23.208 ;
  LAYER M2 ;
        RECT 6.124 23.24 8.596 23.272 ;
  LAYER M2 ;
        RECT 6.124 23.304 8.596 23.336 ;
  LAYER M2 ;
        RECT 6.124 23.368 8.596 23.4 ;
  LAYER M2 ;
        RECT 6.124 23.432 8.596 23.464 ;
  LAYER M2 ;
        RECT 6.124 23.496 8.596 23.528 ;
  LAYER M2 ;
        RECT 6.124 23.56 8.596 23.592 ;
  LAYER M2 ;
        RECT 6.124 23.624 8.596 23.656 ;
  LAYER M3 ;
        RECT 6.144 21.3 6.176 23.808 ;
  LAYER M3 ;
        RECT 6.208 21.3 6.24 23.808 ;
  LAYER M3 ;
        RECT 6.272 21.3 6.304 23.808 ;
  LAYER M3 ;
        RECT 6.336 21.3 6.368 23.808 ;
  LAYER M3 ;
        RECT 6.4 21.3 6.432 23.808 ;
  LAYER M3 ;
        RECT 6.464 21.3 6.496 23.808 ;
  LAYER M3 ;
        RECT 6.528 21.3 6.56 23.808 ;
  LAYER M3 ;
        RECT 6.592 21.3 6.624 23.808 ;
  LAYER M3 ;
        RECT 6.656 21.3 6.688 23.808 ;
  LAYER M3 ;
        RECT 6.72 21.3 6.752 23.808 ;
  LAYER M3 ;
        RECT 6.784 21.3 6.816 23.808 ;
  LAYER M3 ;
        RECT 6.848 21.3 6.88 23.808 ;
  LAYER M3 ;
        RECT 6.912 21.3 6.944 23.808 ;
  LAYER M3 ;
        RECT 6.976 21.3 7.008 23.808 ;
  LAYER M3 ;
        RECT 7.04 21.3 7.072 23.808 ;
  LAYER M3 ;
        RECT 7.104 21.3 7.136 23.808 ;
  LAYER M3 ;
        RECT 7.168 21.3 7.2 23.808 ;
  LAYER M3 ;
        RECT 7.232 21.3 7.264 23.808 ;
  LAYER M3 ;
        RECT 7.296 21.3 7.328 23.808 ;
  LAYER M3 ;
        RECT 7.36 21.3 7.392 23.808 ;
  LAYER M3 ;
        RECT 7.424 21.3 7.456 23.808 ;
  LAYER M3 ;
        RECT 7.488 21.3 7.52 23.808 ;
  LAYER M3 ;
        RECT 7.552 21.3 7.584 23.808 ;
  LAYER M3 ;
        RECT 7.616 21.3 7.648 23.808 ;
  LAYER M3 ;
        RECT 7.68 21.3 7.712 23.808 ;
  LAYER M3 ;
        RECT 7.744 21.3 7.776 23.808 ;
  LAYER M3 ;
        RECT 7.808 21.3 7.84 23.808 ;
  LAYER M3 ;
        RECT 7.872 21.3 7.904 23.808 ;
  LAYER M3 ;
        RECT 7.936 21.3 7.968 23.808 ;
  LAYER M3 ;
        RECT 8 21.3 8.032 23.808 ;
  LAYER M3 ;
        RECT 8.064 21.3 8.096 23.808 ;
  LAYER M3 ;
        RECT 8.128 21.3 8.16 23.808 ;
  LAYER M3 ;
        RECT 8.192 21.3 8.224 23.808 ;
  LAYER M3 ;
        RECT 8.256 21.3 8.288 23.808 ;
  LAYER M3 ;
        RECT 8.32 21.3 8.352 23.808 ;
  LAYER M3 ;
        RECT 8.384 21.3 8.416 23.808 ;
  LAYER M3 ;
        RECT 8.448 21.3 8.48 23.808 ;
  LAYER M3 ;
        RECT 8.544 21.3 8.576 23.808 ;
  LAYER M1 ;
        RECT 6.159 21.336 6.161 23.772 ;
  LAYER M1 ;
        RECT 6.239 21.336 6.241 23.772 ;
  LAYER M1 ;
        RECT 6.319 21.336 6.321 23.772 ;
  LAYER M1 ;
        RECT 6.399 21.336 6.401 23.772 ;
  LAYER M1 ;
        RECT 6.479 21.336 6.481 23.772 ;
  LAYER M1 ;
        RECT 6.559 21.336 6.561 23.772 ;
  LAYER M1 ;
        RECT 6.639 21.336 6.641 23.772 ;
  LAYER M1 ;
        RECT 6.719 21.336 6.721 23.772 ;
  LAYER M1 ;
        RECT 6.799 21.336 6.801 23.772 ;
  LAYER M1 ;
        RECT 6.879 21.336 6.881 23.772 ;
  LAYER M1 ;
        RECT 6.959 21.336 6.961 23.772 ;
  LAYER M1 ;
        RECT 7.039 21.336 7.041 23.772 ;
  LAYER M1 ;
        RECT 7.119 21.336 7.121 23.772 ;
  LAYER M1 ;
        RECT 7.199 21.336 7.201 23.772 ;
  LAYER M1 ;
        RECT 7.279 21.336 7.281 23.772 ;
  LAYER M1 ;
        RECT 7.359 21.336 7.361 23.772 ;
  LAYER M1 ;
        RECT 7.439 21.336 7.441 23.772 ;
  LAYER M1 ;
        RECT 7.519 21.336 7.521 23.772 ;
  LAYER M1 ;
        RECT 7.599 21.336 7.601 23.772 ;
  LAYER M1 ;
        RECT 7.679 21.336 7.681 23.772 ;
  LAYER M1 ;
        RECT 7.759 21.336 7.761 23.772 ;
  LAYER M1 ;
        RECT 7.839 21.336 7.841 23.772 ;
  LAYER M1 ;
        RECT 7.919 21.336 7.921 23.772 ;
  LAYER M1 ;
        RECT 7.999 21.336 8.001 23.772 ;
  LAYER M1 ;
        RECT 8.079 21.336 8.081 23.772 ;
  LAYER M1 ;
        RECT 8.159 21.336 8.161 23.772 ;
  LAYER M1 ;
        RECT 8.239 21.336 8.241 23.772 ;
  LAYER M1 ;
        RECT 8.319 21.336 8.321 23.772 ;
  LAYER M1 ;
        RECT 8.399 21.336 8.401 23.772 ;
  LAYER M1 ;
        RECT 8.479 21.336 8.481 23.772 ;
  LAYER M2 ;
        RECT 6.16 21.335 8.56 21.337 ;
  LAYER M2 ;
        RECT 6.16 21.419 8.56 21.421 ;
  LAYER M2 ;
        RECT 6.16 21.503 8.56 21.505 ;
  LAYER M2 ;
        RECT 6.16 21.587 8.56 21.589 ;
  LAYER M2 ;
        RECT 6.16 21.671 8.56 21.673 ;
  LAYER M2 ;
        RECT 6.16 21.755 8.56 21.757 ;
  LAYER M2 ;
        RECT 6.16 21.839 8.56 21.841 ;
  LAYER M2 ;
        RECT 6.16 21.923 8.56 21.925 ;
  LAYER M2 ;
        RECT 6.16 22.007 8.56 22.009 ;
  LAYER M2 ;
        RECT 6.16 22.091 8.56 22.093 ;
  LAYER M2 ;
        RECT 6.16 22.175 8.56 22.177 ;
  LAYER M2 ;
        RECT 6.16 22.259 8.56 22.261 ;
  LAYER M2 ;
        RECT 6.16 22.3425 8.56 22.3445 ;
  LAYER M2 ;
        RECT 6.16 22.427 8.56 22.429 ;
  LAYER M2 ;
        RECT 6.16 22.511 8.56 22.513 ;
  LAYER M2 ;
        RECT 6.16 22.595 8.56 22.597 ;
  LAYER M2 ;
        RECT 6.16 22.679 8.56 22.681 ;
  LAYER M2 ;
        RECT 6.16 22.763 8.56 22.765 ;
  LAYER M2 ;
        RECT 6.16 22.847 8.56 22.849 ;
  LAYER M2 ;
        RECT 6.16 22.931 8.56 22.933 ;
  LAYER M2 ;
        RECT 6.16 23.015 8.56 23.017 ;
  LAYER M2 ;
        RECT 6.16 23.099 8.56 23.101 ;
  LAYER M2 ;
        RECT 6.16 23.183 8.56 23.185 ;
  LAYER M2 ;
        RECT 6.16 23.267 8.56 23.269 ;
  LAYER M2 ;
        RECT 6.16 23.351 8.56 23.353 ;
  LAYER M2 ;
        RECT 6.16 23.435 8.56 23.437 ;
  LAYER M2 ;
        RECT 6.16 23.519 8.56 23.521 ;
  LAYER M2 ;
        RECT 6.16 23.603 8.56 23.605 ;
  LAYER M2 ;
        RECT 6.16 23.687 8.56 23.689 ;
  END 
END Cap_60fF
