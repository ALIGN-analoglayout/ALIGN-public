MACRO cap_test
  ORIGIN 0 0 ;
  FOREIGN cap_test 0 0 ;
  SIZE 2.3680 BY 2.4360 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 2.3400 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 2.3360 2.3400 2.3680 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.0480 0.0480 0.0800 2.3880 ;
    LAYER M3 ;
      RECT 0.0480 0.0480 0.0800 2.3880 ;
    LAYER V1 ;
      RECT 0.0480 2.3360 0.0800 2.3680 ;
    LAYER V1 ;
      RECT 0.0480 2.3360 0.0800 2.3680 ;
    LAYER M1 ;
      RECT 0.1120 0.0480 0.1440 2.3880 ;
    LAYER M3 ;
      RECT 0.1120 0.0480 0.1440 2.3880 ;
    LAYER V1 ;
      RECT 0.1120 0.0680 0.1440 0.1000 ;
    LAYER V1 ;
      RECT 0.1120 0.0680 0.1440 0.1000 ;
    LAYER M1 ;
      RECT 0.1760 0.0480 0.2080 2.3880 ;
    LAYER M3 ;
      RECT 0.1760 0.0480 0.2080 2.3880 ;
    LAYER V1 ;
      RECT 0.1760 2.3360 0.2080 2.3680 ;
    LAYER V1 ;
      RECT 0.1760 2.3360 0.2080 2.3680 ;
    LAYER M1 ;
      RECT 0.2400 0.0480 0.2720 2.3880 ;
    LAYER M3 ;
      RECT 0.2400 0.0480 0.2720 2.3880 ;
    LAYER V1 ;
      RECT 0.2400 0.0680 0.2720 0.1000 ;
    LAYER V1 ;
      RECT 0.2400 0.0680 0.2720 0.1000 ;
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 2.3880 ;
    LAYER M3 ;
      RECT 0.3040 0.0480 0.3360 2.3880 ;
    LAYER V1 ;
      RECT 0.3040 2.3360 0.3360 2.3680 ;
    LAYER V1 ;
      RECT 0.3040 2.3360 0.3360 2.3680 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 2.3880 ;
    LAYER M3 ;
      RECT 0.3680 0.0480 0.4000 2.3880 ;
    LAYER V1 ;
      RECT 0.3680 0.0680 0.4000 0.1000 ;
    LAYER V1 ;
      RECT 0.3680 0.0680 0.4000 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 2.3880 ;
    LAYER M3 ;
      RECT 0.4320 0.0480 0.4640 2.3880 ;
    LAYER V1 ;
      RECT 0.4320 2.3360 0.4640 2.3680 ;
    LAYER V1 ;
      RECT 0.4320 2.3360 0.4640 2.3680 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 2.3880 ;
    LAYER M3 ;
      RECT 0.4960 0.0480 0.5280 2.3880 ;
    LAYER V1 ;
      RECT 0.4960 0.0680 0.5280 0.1000 ;
    LAYER V1 ;
      RECT 0.4960 0.0680 0.5280 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 2.3880 ;
    LAYER M3 ;
      RECT 0.5600 0.0480 0.5920 2.3880 ;
    LAYER V1 ;
      RECT 0.5600 2.3360 0.5920 2.3680 ;
    LAYER V1 ;
      RECT 0.5600 2.3360 0.5920 2.3680 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 2.3880 ;
    LAYER M3 ;
      RECT 0.6240 0.0480 0.6560 2.3880 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER M1 ;
      RECT 0.6880 0.0480 0.7200 2.3880 ;
    LAYER M3 ;
      RECT 0.6880 0.0480 0.7200 2.3880 ;
    LAYER V1 ;
      RECT 0.6880 2.3360 0.7200 2.3680 ;
    LAYER V1 ;
      RECT 0.6880 2.3360 0.7200 2.3680 ;
    LAYER M1 ;
      RECT 0.7520 0.0480 0.7840 2.3880 ;
    LAYER M3 ;
      RECT 0.7520 0.0480 0.7840 2.3880 ;
    LAYER V1 ;
      RECT 0.7520 0.0680 0.7840 0.1000 ;
    LAYER V1 ;
      RECT 0.7520 0.0680 0.7840 0.1000 ;
    LAYER M1 ;
      RECT 0.8160 0.0480 0.8480 2.3880 ;
    LAYER M3 ;
      RECT 0.8160 0.0480 0.8480 2.3880 ;
    LAYER V1 ;
      RECT 0.8160 2.3360 0.8480 2.3680 ;
    LAYER V1 ;
      RECT 0.8160 2.3360 0.8480 2.3680 ;
    LAYER M1 ;
      RECT 0.8800 0.0480 0.9120 2.3880 ;
    LAYER M3 ;
      RECT 0.8800 0.0480 0.9120 2.3880 ;
    LAYER V1 ;
      RECT 0.8800 0.0680 0.9120 0.1000 ;
    LAYER V1 ;
      RECT 0.8800 0.0680 0.9120 0.1000 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 2.3880 ;
    LAYER M3 ;
      RECT 0.9440 0.0480 0.9760 2.3880 ;
    LAYER V1 ;
      RECT 0.9440 2.3360 0.9760 2.3680 ;
    LAYER V1 ;
      RECT 0.9440 2.3360 0.9760 2.3680 ;
    LAYER M1 ;
      RECT 1.0080 0.0480 1.0400 2.3880 ;
    LAYER M3 ;
      RECT 1.0080 0.0480 1.0400 2.3880 ;
    LAYER V1 ;
      RECT 1.0080 0.0680 1.0400 0.1000 ;
    LAYER V1 ;
      RECT 1.0080 0.0680 1.0400 0.1000 ;
    LAYER M1 ;
      RECT 1.0720 0.0480 1.1040 2.3880 ;
    LAYER M3 ;
      RECT 1.0720 0.0480 1.1040 2.3880 ;
    LAYER V1 ;
      RECT 1.0720 2.3360 1.1040 2.3680 ;
    LAYER V1 ;
      RECT 1.0720 2.3360 1.1040 2.3680 ;
    LAYER M1 ;
      RECT 1.1360 0.0480 1.1680 2.3880 ;
    LAYER M3 ;
      RECT 1.1360 0.0480 1.1680 2.3880 ;
    LAYER V1 ;
      RECT 1.1360 0.0680 1.1680 0.1000 ;
    LAYER V1 ;
      RECT 1.1360 0.0680 1.1680 0.1000 ;
    LAYER M1 ;
      RECT 1.2000 0.0480 1.2320 2.3880 ;
    LAYER M3 ;
      RECT 1.2000 0.0480 1.2320 2.3880 ;
    LAYER V1 ;
      RECT 1.2000 2.3360 1.2320 2.3680 ;
    LAYER V1 ;
      RECT 1.2000 2.3360 1.2320 2.3680 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 2.3880 ;
    LAYER M3 ;
      RECT 1.2640 0.0480 1.2960 2.3880 ;
    LAYER V1 ;
      RECT 1.2640 0.0680 1.2960 0.1000 ;
    LAYER V1 ;
      RECT 1.2640 0.0680 1.2960 0.1000 ;
    LAYER M1 ;
      RECT 1.3280 0.0480 1.3600 2.3880 ;
    LAYER M3 ;
      RECT 1.3280 0.0480 1.3600 2.3880 ;
    LAYER V1 ;
      RECT 1.3280 2.3360 1.3600 2.3680 ;
    LAYER V1 ;
      RECT 1.3280 2.3360 1.3600 2.3680 ;
    LAYER M1 ;
      RECT 1.3920 0.0480 1.4240 2.3880 ;
    LAYER M3 ;
      RECT 1.3920 0.0480 1.4240 2.3880 ;
    LAYER V1 ;
      RECT 1.3920 0.0680 1.4240 0.1000 ;
    LAYER V1 ;
      RECT 1.3920 0.0680 1.4240 0.1000 ;
    LAYER M1 ;
      RECT 1.4560 0.0480 1.4880 2.3880 ;
    LAYER M3 ;
      RECT 1.4560 0.0480 1.4880 2.3880 ;
    LAYER V1 ;
      RECT 1.4560 2.3360 1.4880 2.3680 ;
    LAYER V1 ;
      RECT 1.4560 2.3360 1.4880 2.3680 ;
    LAYER M1 ;
      RECT 1.5200 0.0480 1.5520 2.3880 ;
    LAYER M3 ;
      RECT 1.5200 0.0480 1.5520 2.3880 ;
    LAYER V1 ;
      RECT 1.5200 0.0680 1.5520 0.1000 ;
    LAYER V1 ;
      RECT 1.5200 0.0680 1.5520 0.1000 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 2.3880 ;
    LAYER M3 ;
      RECT 1.5840 0.0480 1.6160 2.3880 ;
    LAYER V1 ;
      RECT 1.5840 2.3360 1.6160 2.3680 ;
    LAYER V1 ;
      RECT 1.5840 2.3360 1.6160 2.3680 ;
    LAYER M1 ;
      RECT 1.6480 0.0480 1.6800 2.3880 ;
    LAYER M3 ;
      RECT 1.6480 0.0480 1.6800 2.3880 ;
    LAYER V1 ;
      RECT 1.6480 0.0680 1.6800 0.1000 ;
    LAYER V1 ;
      RECT 1.6480 0.0680 1.6800 0.1000 ;
    LAYER M1 ;
      RECT 1.7120 0.0480 1.7440 2.3880 ;
    LAYER M3 ;
      RECT 1.7120 0.0480 1.7440 2.3880 ;
    LAYER V1 ;
      RECT 1.7120 2.3360 1.7440 2.3680 ;
    LAYER V1 ;
      RECT 1.7120 2.3360 1.7440 2.3680 ;
    LAYER M1 ;
      RECT 1.7760 0.0480 1.8080 2.3880 ;
    LAYER M3 ;
      RECT 1.7760 0.0480 1.8080 2.3880 ;
    LAYER V1 ;
      RECT 1.7760 0.0680 1.8080 0.1000 ;
    LAYER V1 ;
      RECT 1.7760 0.0680 1.8080 0.1000 ;
    LAYER M1 ;
      RECT 1.8400 0.0480 1.8720 2.3880 ;
    LAYER M3 ;
      RECT 1.8400 0.0480 1.8720 2.3880 ;
    LAYER V1 ;
      RECT 1.8400 2.3360 1.8720 2.3680 ;
    LAYER V1 ;
      RECT 1.8400 2.3360 1.8720 2.3680 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 2.3880 ;
    LAYER M3 ;
      RECT 1.9040 0.0480 1.9360 2.3880 ;
    LAYER V1 ;
      RECT 1.9040 0.0680 1.9360 0.1000 ;
    LAYER V1 ;
      RECT 1.9040 0.0680 1.9360 0.1000 ;
    LAYER M1 ;
      RECT 1.9680 0.0480 2.0000 2.3880 ;
    LAYER M3 ;
      RECT 1.9680 0.0480 2.0000 2.3880 ;
    LAYER V1 ;
      RECT 1.9680 2.3360 2.0000 2.3680 ;
    LAYER V1 ;
      RECT 1.9680 2.3360 2.0000 2.3680 ;
    LAYER M1 ;
      RECT 2.0320 0.0480 2.0640 2.3880 ;
    LAYER M3 ;
      RECT 2.0320 0.0480 2.0640 2.3880 ;
    LAYER V1 ;
      RECT 2.0320 0.0680 2.0640 0.1000 ;
    LAYER V1 ;
      RECT 2.0320 0.0680 2.0640 0.1000 ;
    LAYER M1 ;
      RECT 2.0960 0.0480 2.1280 2.3880 ;
    LAYER M3 ;
      RECT 2.0960 0.0480 2.1280 2.3880 ;
    LAYER V1 ;
      RECT 2.0960 2.3360 2.1280 2.3680 ;
    LAYER V1 ;
      RECT 2.0960 2.3360 2.1280 2.3680 ;
    LAYER M1 ;
      RECT 2.1600 0.0480 2.1920 2.3880 ;
    LAYER M3 ;
      RECT 2.1600 0.0480 2.1920 2.3880 ;
    LAYER V1 ;
      RECT 2.1600 0.0680 2.1920 0.1000 ;
    LAYER V1 ;
      RECT 2.1600 0.0680 2.1920 0.1000 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 2.3880 ;
    LAYER M3 ;
      RECT 2.2240 0.0480 2.2560 2.3880 ;
    LAYER V1 ;
      RECT 2.2240 2.3360 2.2560 2.3680 ;
    LAYER V1 ;
      RECT 2.2240 2.3360 2.2560 2.3680 ;
    LAYER M1 ;
      RECT 2.2880 0.0480 2.3200 2.3880 ;
    LAYER M3 ;
      RECT 2.2880 0.0480 2.3200 2.3880 ;
    LAYER V1 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER V1 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER V1 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER V2 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER V1 ;
      RECT 0.0480 0.1320 0.0800 0.1640 ;
    LAYER V2 ;
      RECT 0.0480 0.1320 0.0800 0.1640 ;
    LAYER M2 ;
      RECT 0.0280 0.1320 2.3400 0.1640 ;
    LAYER V1 ;
      RECT 2.2880 0.1960 2.3200 0.2280 ;
    LAYER V2 ;
      RECT 2.2880 0.1960 2.3200 0.2280 ;
    LAYER M2 ;
      RECT 0.0280 0.1960 2.3400 0.2280 ;
    LAYER V1 ;
      RECT 0.0480 0.2600 0.0800 0.2920 ;
    LAYER V2 ;
      RECT 0.0480 0.2600 0.0800 0.2920 ;
    LAYER M2 ;
      RECT 0.0280 0.2600 2.3400 0.2920 ;
    LAYER V1 ;
      RECT 2.2880 0.3240 2.3200 0.3560 ;
    LAYER V2 ;
      RECT 2.2880 0.3240 2.3200 0.3560 ;
    LAYER M2 ;
      RECT 0.0280 0.3240 2.3400 0.3560 ;
    LAYER V1 ;
      RECT 0.0480 0.3880 0.0800 0.4200 ;
    LAYER V2 ;
      RECT 0.0480 0.3880 0.0800 0.4200 ;
    LAYER M2 ;
      RECT 0.0280 0.3880 2.3400 0.4200 ;
    LAYER V1 ;
      RECT 2.2880 0.4520 2.3200 0.4840 ;
    LAYER V2 ;
      RECT 2.2880 0.4520 2.3200 0.4840 ;
    LAYER M2 ;
      RECT 0.0280 0.4520 2.3400 0.4840 ;
    LAYER V1 ;
      RECT 0.0480 0.5160 0.0800 0.5480 ;
    LAYER V2 ;
      RECT 0.0480 0.5160 0.0800 0.5480 ;
    LAYER M2 ;
      RECT 0.0280 0.5160 2.3400 0.5480 ;
    LAYER V1 ;
      RECT 2.2880 0.5800 2.3200 0.6120 ;
    LAYER V2 ;
      RECT 2.2880 0.5800 2.3200 0.6120 ;
    LAYER M2 ;
      RECT 0.0280 0.5800 2.3400 0.6120 ;
    LAYER V1 ;
      RECT 0.0480 0.6440 0.0800 0.6760 ;
    LAYER V2 ;
      RECT 0.0480 0.6440 0.0800 0.6760 ;
    LAYER M2 ;
      RECT 0.0280 0.6440 2.3400 0.6760 ;
    LAYER V1 ;
      RECT 2.2880 0.7080 2.3200 0.7400 ;
    LAYER V2 ;
      RECT 2.2880 0.7080 2.3200 0.7400 ;
    LAYER M2 ;
      RECT 0.0280 0.7080 2.3400 0.7400 ;
    LAYER V1 ;
      RECT 0.0480 0.7720 0.0800 0.8040 ;
    LAYER V2 ;
      RECT 0.0480 0.7720 0.0800 0.8040 ;
    LAYER M2 ;
      RECT 0.0280 0.7720 2.3400 0.8040 ;
    LAYER V1 ;
      RECT 2.2880 0.8360 2.3200 0.8680 ;
    LAYER V2 ;
      RECT 2.2880 0.8360 2.3200 0.8680 ;
    LAYER M2 ;
      RECT 0.0280 0.8360 2.3400 0.8680 ;
    LAYER V1 ;
      RECT 0.0480 0.9000 0.0800 0.9320 ;
    LAYER V2 ;
      RECT 0.0480 0.9000 0.0800 0.9320 ;
    LAYER M2 ;
      RECT 0.0280 0.9000 2.3400 0.9320 ;
    LAYER V1 ;
      RECT 2.2880 0.9640 2.3200 0.9960 ;
    LAYER V2 ;
      RECT 2.2880 0.9640 2.3200 0.9960 ;
    LAYER M2 ;
      RECT 0.0280 0.9640 2.3400 0.9960 ;
    LAYER V1 ;
      RECT 0.0480 1.0280 0.0800 1.0600 ;
    LAYER V2 ;
      RECT 0.0480 1.0280 0.0800 1.0600 ;
    LAYER M2 ;
      RECT 0.0280 1.0280 2.3400 1.0600 ;
    LAYER V1 ;
      RECT 2.2880 1.0920 2.3200 1.1240 ;
    LAYER V2 ;
      RECT 2.2880 1.0920 2.3200 1.1240 ;
    LAYER M2 ;
      RECT 0.0280 1.0920 2.3400 1.1240 ;
    LAYER V1 ;
      RECT 0.0480 1.1560 0.0800 1.1880 ;
    LAYER V2 ;
      RECT 0.0480 1.1560 0.0800 1.1880 ;
    LAYER M2 ;
      RECT 0.0280 1.1560 2.3400 1.1880 ;
    LAYER V1 ;
      RECT 2.2880 1.2200 2.3200 1.2520 ;
    LAYER V2 ;
      RECT 2.2880 1.2200 2.3200 1.2520 ;
    LAYER M2 ;
      RECT 0.0280 1.2200 2.3400 1.2520 ;
    LAYER V1 ;
      RECT 0.0480 1.2840 0.0800 1.3160 ;
    LAYER V2 ;
      RECT 0.0480 1.2840 0.0800 1.3160 ;
    LAYER M2 ;
      RECT 0.0280 1.2840 2.3400 1.3160 ;
    LAYER V1 ;
      RECT 2.2880 1.3480 2.3200 1.3800 ;
    LAYER V2 ;
      RECT 2.2880 1.3480 2.3200 1.3800 ;
    LAYER M2 ;
      RECT 0.0280 1.3480 2.3400 1.3800 ;
    LAYER V1 ;
      RECT 0.0480 1.4120 0.0800 1.4440 ;
    LAYER V2 ;
      RECT 0.0480 1.4120 0.0800 1.4440 ;
    LAYER M2 ;
      RECT 0.0280 1.4120 2.3400 1.4440 ;
    LAYER V1 ;
      RECT 2.2880 1.4760 2.3200 1.5080 ;
    LAYER V2 ;
      RECT 2.2880 1.4760 2.3200 1.5080 ;
    LAYER M2 ;
      RECT 0.0280 1.4760 2.3400 1.5080 ;
    LAYER V1 ;
      RECT 0.0480 1.5400 0.0800 1.5720 ;
    LAYER V2 ;
      RECT 0.0480 1.5400 0.0800 1.5720 ;
    LAYER M2 ;
      RECT 0.0280 1.5400 2.3400 1.5720 ;
    LAYER V1 ;
      RECT 2.2880 1.6040 2.3200 1.6360 ;
    LAYER V2 ;
      RECT 2.2880 1.6040 2.3200 1.6360 ;
    LAYER M2 ;
      RECT 0.0280 1.6040 2.3400 1.6360 ;
    LAYER V1 ;
      RECT 0.0480 1.6680 0.0800 1.7000 ;
    LAYER V2 ;
      RECT 0.0480 1.6680 0.0800 1.7000 ;
    LAYER M2 ;
      RECT 0.0280 1.6680 2.3400 1.7000 ;
    LAYER V1 ;
      RECT 2.2880 1.7320 2.3200 1.7640 ;
    LAYER V2 ;
      RECT 2.2880 1.7320 2.3200 1.7640 ;
    LAYER M2 ;
      RECT 0.0280 1.7320 2.3400 1.7640 ;
    LAYER V1 ;
      RECT 0.0480 1.7960 0.0800 1.8280 ;
    LAYER V2 ;
      RECT 0.0480 1.7960 0.0800 1.8280 ;
    LAYER M2 ;
      RECT 0.0280 1.7960 2.3400 1.8280 ;
    LAYER V1 ;
      RECT 2.2880 1.8600 2.3200 1.8920 ;
    LAYER V2 ;
      RECT 2.2880 1.8600 2.3200 1.8920 ;
    LAYER M2 ;
      RECT 0.0280 1.8600 2.3400 1.8920 ;
    LAYER V1 ;
      RECT 0.0480 1.9240 0.0800 1.9560 ;
    LAYER V2 ;
      RECT 0.0480 1.9240 0.0800 1.9560 ;
    LAYER M2 ;
      RECT 0.0280 1.9240 2.3400 1.9560 ;
    LAYER V1 ;
      RECT 2.2880 1.9880 2.3200 2.0200 ;
    LAYER V2 ;
      RECT 2.2880 1.9880 2.3200 2.0200 ;
    LAYER M2 ;
      RECT 0.0280 1.9880 2.3400 2.0200 ;
    LAYER V1 ;
      RECT 0.0480 2.0520 0.0800 2.0840 ;
    LAYER V2 ;
      RECT 0.0480 2.0520 0.0800 2.0840 ;
    LAYER M2 ;
      RECT 0.0280 2.0520 2.3400 2.0840 ;
    LAYER V1 ;
      RECT 2.2880 2.1160 2.3200 2.1480 ;
    LAYER V2 ;
      RECT 2.2880 2.1160 2.3200 2.1480 ;
    LAYER M2 ;
      RECT 0.0280 2.1160 2.3400 2.1480 ;
    LAYER V1 ;
      RECT 0.0480 2.1800 0.0800 2.2120 ;
    LAYER V2 ;
      RECT 0.0480 2.1800 0.0800 2.2120 ;
    LAYER M2 ;
      RECT 0.0280 2.1800 2.3400 2.2120 ;
    LAYER V1 ;
      RECT 2.2880 2.2440 2.3200 2.2760 ;
    LAYER V2 ;
      RECT 2.2880 2.2440 2.3200 2.2760 ;
    LAYER M2 ;
      RECT 0.0280 2.2440 2.3400 2.2760 ;
    LAYER boundary ;
      RECT 0.0000 0.0000 2.3680 2.4360 ;
  END
END cap_test
