MACRO switched_capacitor_filter
  ORIGIN 0 0 ;
  FOREIGN switched_capacitor_filter 0 0 ;
  SIZE 46.08 BY 37.8 ;
  PIN id
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.184 -0.016 23.216 0.016 ;
      LAYER M3 ;
        RECT 23.18 0.3 23.22 0.708 ;
      LAYER M3 ;
        RECT 22.86 0.3 22.9 0.708 ;
      LAYER M3 ;
        RECT 23.18 0.399 23.22 0.609 ;
      LAYER M4 ;
        RECT 23.2 0.484 23.68 0.524 ;
      LAYER M3 ;
        RECT 23.66 0 23.7 0.504 ;
      LAYER M2 ;
        RECT 23.2 -0.016 23.68 0.016 ;
    END
  END id
  PIN voutn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.264 37.784 15.296 37.816 ;
      LAYER M2 ;
        RECT 22.124 4.436 23.956 4.468 ;
      LAYER M2 ;
        RECT 21.964 3.008 24.596 3.04 ;
      LAYER M2 ;
        RECT 22.46 4.436 22.66 4.468 ;
      LAYER M3 ;
        RECT 22.54 3.192 22.58 4.452 ;
      LAYER M4 ;
        RECT 22.49 3.172 22.63 3.212 ;
      LAYER M5 ;
        RECT 22.528 3.024 22.592 3.192 ;
      LAYER M4 ;
        RECT 22.49 3.004 22.63 3.044 ;
      LAYER M3 ;
        RECT 22.54 2.919 22.58 3.129 ;
      LAYER M2 ;
        RECT 22.46 3.008 22.66 3.04 ;
      LAYER M2 ;
        RECT 7.244 0.824 7.476 0.856 ;
      LAYER M1 ;
        RECT 11.744 1.308 11.776 1.38 ;
      LAYER M2 ;
        RECT 11.724 1.328 11.796 1.36 ;
      LAYER M1 ;
        RECT 3.104 1.308 3.136 1.38 ;
      LAYER M2 ;
        RECT 3.084 1.328 3.156 1.36 ;
      LAYER M2 ;
        RECT 3.12 1.328 11.76 1.36 ;
      LAYER M2 ;
        RECT 7.18 0.824 7.38 0.856 ;
      LAYER M3 ;
        RECT 7.26 0.84 7.3 1.344 ;
      LAYER M2 ;
        RECT 7.18 1.328 7.38 1.36 ;
      LAYER M1 ;
        RECT 21.504 37.344 21.536 37.416 ;
      LAYER M2 ;
        RECT 21.484 37.364 21.556 37.396 ;
      LAYER M1 ;
        RECT 24.384 37.344 24.416 37.416 ;
      LAYER M2 ;
        RECT 24.364 37.364 24.436 37.396 ;
      LAYER M2 ;
        RECT 21.52 37.364 24.4 37.396 ;
      LAYER M2 ;
        RECT 21.04 3.008 22 3.04 ;
      LAYER M3 ;
        RECT 21.02 2.919 21.06 3.129 ;
      LAYER M4 ;
        RECT 20.88 3.004 21.04 3.044 ;
      LAYER M5 ;
        RECT 20.848 3.024 20.912 3.36 ;
      LAYER M4 ;
        RECT 12.816 3.34 20.88 3.38 ;
      LAYER M5 ;
        RECT 12.784 1.596 12.848 3.36 ;
      LAYER M4 ;
        RECT 12.24 1.576 12.816 1.616 ;
      LAYER M3 ;
        RECT 12.22 1.344 12.26 1.596 ;
      LAYER M2 ;
        RECT 11.76 1.328 12.24 1.36 ;
      LAYER M2 ;
        RECT 23.66 4.436 23.86 4.468 ;
      LAYER M3 ;
        RECT 23.74 4.452 23.78 4.956 ;
      LAYER M4 ;
        RECT 23.76 4.936 25.632 4.976 ;
      LAYER M5 ;
        RECT 25.6 4.956 25.664 37.38 ;
      LAYER M4 ;
        RECT 25.2 37.36 25.632 37.4 ;
      LAYER M3 ;
        RECT 25.18 37.275 25.22 37.485 ;
      LAYER M2 ;
        RECT 24.72 37.364 25.2 37.396 ;
      LAYER M3 ;
        RECT 24.7 37.275 24.74 37.485 ;
      LAYER M4 ;
        RECT 24.4 37.36 24.72 37.4 ;
      LAYER M3 ;
        RECT 24.38 37.275 24.42 37.485 ;
      LAYER M2 ;
        RECT 24.3 37.364 24.5 37.396 ;
      LAYER M2 ;
        RECT 19.6 37.364 21.52 37.396 ;
      LAYER M3 ;
        RECT 19.58 37.275 19.62 37.485 ;
      LAYER M4 ;
        RECT 19.296 37.36 19.6 37.4 ;
      LAYER M5 ;
        RECT 19.264 35.28 19.328 37.38 ;
      LAYER M6 ;
        RECT 15.84 35.248 19.296 35.312 ;
      LAYER M5 ;
        RECT 15.808 35.28 15.872 37.548 ;
      LAYER M4 ;
        RECT 15.77 37.528 15.91 37.568 ;
      LAYER M3 ;
        RECT 15.82 37.443 15.86 37.653 ;
      LAYER M2 ;
        RECT 15.6 37.532 15.84 37.564 ;
      LAYER M3 ;
        RECT 15.58 37.548 15.62 37.8 ;
      LAYER M4 ;
        RECT 15.28 37.78 15.6 37.82 ;
      LAYER M3 ;
        RECT 15.26 37.695 15.3 37.905 ;
      LAYER M2 ;
        RECT 15.18 37.784 15.38 37.816 ;
    END
  END voutn
  PIN voutp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 30.704 37.784 30.736 37.816 ;
      LAYER M2 ;
        RECT 22.764 4.268 23.316 4.3 ;
      LAYER M2 ;
        RECT 21.324 3.176 23.956 3.208 ;
      LAYER M2 ;
        RECT 23.18 4.268 23.38 4.3 ;
      LAYER M3 ;
        RECT 23.26 4.032 23.3 4.284 ;
      LAYER M4 ;
        RECT 23.21 4.012 23.35 4.052 ;
      LAYER M5 ;
        RECT 23.248 3.696 23.312 4.032 ;
      LAYER M4 ;
        RECT 23.21 3.676 23.35 3.716 ;
      LAYER M3 ;
        RECT 23.26 3.192 23.3 3.696 ;
      LAYER M2 ;
        RECT 23.18 3.176 23.38 3.208 ;
      LAYER M2 ;
        RECT 38.604 0.824 38.836 0.856 ;
      LAYER M1 ;
        RECT 34.304 1.308 34.336 1.38 ;
      LAYER M2 ;
        RECT 34.284 1.328 34.356 1.36 ;
      LAYER M1 ;
        RECT 42.944 1.308 42.976 1.38 ;
      LAYER M2 ;
        RECT 42.924 1.328 42.996 1.36 ;
      LAYER M2 ;
        RECT 34.32 1.328 42.96 1.36 ;
      LAYER M2 ;
        RECT 38.7 0.824 38.9 0.856 ;
      LAYER M3 ;
        RECT 38.78 0.84 38.82 1.344 ;
      LAYER M2 ;
        RECT 38.7 1.328 38.9 1.36 ;
      LAYER M1 ;
        RECT 18.624 37.512 18.656 37.584 ;
      LAYER M2 ;
        RECT 18.604 37.532 18.676 37.564 ;
      LAYER M1 ;
        RECT 27.264 37.512 27.296 37.584 ;
      LAYER M2 ;
        RECT 27.244 37.532 27.316 37.564 ;
      LAYER M2 ;
        RECT 18.64 37.532 27.28 37.564 ;
      LAYER M2 ;
        RECT 23.92 3.176 25.36 3.208 ;
      LAYER M3 ;
        RECT 25.34 3.087 25.38 3.297 ;
      LAYER M4 ;
        RECT 25.354 3.172 25.494 3.212 ;
      LAYER M5 ;
        RECT 25.456 3.192 25.52 3.36 ;
      LAYER M4 ;
        RECT 25.488 3.34 33.552 3.38 ;
      LAYER M5 ;
        RECT 33.52 1.596 33.584 3.36 ;
      LAYER M4 ;
        RECT 33.552 1.576 34.32 1.616 ;
      LAYER M3 ;
        RECT 34.3 1.344 34.34 1.596 ;
      LAYER M2 ;
        RECT 34.22 1.328 34.42 1.36 ;
      LAYER M4 ;
        RECT 25.85 3.34 25.99 3.38 ;
      LAYER M3 ;
        RECT 25.9 3.36 25.94 5.628 ;
      LAYER M4 ;
        RECT 25.85 5.608 25.99 5.648 ;
      LAYER M5 ;
        RECT 25.888 5.628 25.952 37.548 ;
      LAYER M4 ;
        RECT 25.85 37.528 25.99 37.568 ;
      LAYER M3 ;
        RECT 25.9 37.443 25.94 37.653 ;
      LAYER M2 ;
        RECT 25.82 37.532 26.02 37.564 ;
      LAYER M2 ;
        RECT 27.28 37.532 30.4 37.564 ;
      LAYER M3 ;
        RECT 30.38 37.548 30.42 37.8 ;
      LAYER M4 ;
        RECT 30.4 37.78 30.72 37.82 ;
      LAYER M3 ;
        RECT 30.7 37.695 30.74 37.905 ;
      LAYER M2 ;
        RECT 30.62 37.784 30.82 37.816 ;
    END
  END voutp
  PIN vss
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 22.784 -0.016 22.816 0.016 ;
      LAYER M3 ;
        RECT 23.26 0.216 23.3 0.624 ;
      LAYER M3 ;
        RECT 22.94 0.216 22.98 0.624 ;
      LAYER M1 ;
        RECT 21.664 19.2 21.696 19.272 ;
      LAYER M2 ;
        RECT 21.644 19.22 21.716 19.252 ;
      LAYER M1 ;
        RECT 24.544 19.2 24.576 19.272 ;
      LAYER M2 ;
        RECT 24.524 19.22 24.596 19.252 ;
      LAYER M2 ;
        RECT 21.68 19.22 24.56 19.252 ;
      LAYER M1 ;
        RECT 18.784 19.032 18.816 19.104 ;
      LAYER M2 ;
        RECT 18.764 19.052 18.836 19.084 ;
      LAYER M1 ;
        RECT 27.424 19.032 27.456 19.104 ;
      LAYER M2 ;
        RECT 27.404 19.052 27.476 19.084 ;
      LAYER M2 ;
        RECT 18.8 19.052 27.44 19.084 ;
      LAYER M3 ;
        RECT 22.94 0 22.98 0.252 ;
      LAYER M2 ;
        RECT 22.72 -0.016 22.96 0.016 ;
      LAYER M3 ;
        RECT 22.7 0 22.74 0.252 ;
      LAYER M4 ;
        RECT 22.56 0.232 22.72 0.272 ;
      LAYER M3 ;
        RECT 22.54 0 22.58 0.252 ;
      LAYER M2 ;
        RECT 22.56 -0.016 22.8 0.016 ;
      LAYER M3 ;
        RECT 23.26 0.588 23.3 1.344 ;
      LAYER M2 ;
        RECT 23.28 1.328 23.76 1.36 ;
      LAYER M3 ;
        RECT 23.74 1.344 23.78 1.596 ;
      LAYER M4 ;
        RECT 23.76 1.576 25.776 1.616 ;
      LAYER M5 ;
        RECT 25.744 1.596 25.808 19.236 ;
      LAYER M4 ;
        RECT 24.48 19.216 25.776 19.256 ;
      LAYER M3 ;
        RECT 24.46 19.131 24.5 19.341 ;
      LAYER M2 ;
        RECT 24.38 19.22 24.58 19.252 ;
      LAYER M5 ;
        RECT 25.744 19.018 25.808 19.118 ;
      LAYER M4 ;
        RECT 25.776 19.048 25.92 19.088 ;
      LAYER M3 ;
        RECT 25.9 18.963 25.94 19.173 ;
      LAYER M2 ;
        RECT 25.82 19.052 26.02 19.084 ;
    END
  END vss
  PIN vinn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.024 -0.016 15.056 0.016 ;
      LAYER M3 ;
        RECT 15.02 17.688 15.06 18.012 ;
      LAYER M3 ;
        RECT 15.26 17.688 15.3 18.012 ;
      LAYER M1 ;
        RECT 27.424 18.444 27.456 18.516 ;
      LAYER M2 ;
        RECT 27.404 18.464 27.476 18.496 ;
      LAYER M1 ;
        RECT 18.784 18.444 18.816 18.516 ;
      LAYER M2 ;
        RECT 18.764 18.464 18.836 18.496 ;
      LAYER M2 ;
        RECT 18.8 18.464 27.44 18.496 ;
      LAYER M3 ;
        RECT 15.26 17.976 15.3 18.48 ;
      LAYER M4 ;
        RECT 15.28 18.46 15.92 18.5 ;
      LAYER M3 ;
        RECT 15.9 18.375 15.94 18.585 ;
      LAYER M2 ;
        RECT 15.92 18.464 18.8 18.496 ;
      LAYER M3 ;
        RECT 15.02 16.968 15.06 17.724 ;
      LAYER M4 ;
        RECT 14.4 16.948 15.04 16.988 ;
      LAYER M5 ;
        RECT 14.368 0.756 14.432 16.968 ;
      LAYER M4 ;
        RECT 14.4 0.736 14.56 0.776 ;
      LAYER M3 ;
        RECT 14.54 0.504 14.58 0.756 ;
      LAYER M2 ;
        RECT 14.56 0.488 14.8 0.52 ;
      LAYER M3 ;
        RECT 14.78 0 14.82 0.504 ;
      LAYER M2 ;
        RECT 14.8 -0.016 15.04 0.016 ;
    END
  END vinn
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.344 -0.016 15.376 0.016 ;
      LAYER M3 ;
        RECT 4.94 0.636 4.98 0.96 ;
      LAYER M3 ;
        RECT 5.18 0.636 5.22 0.96 ;
      LAYER M2 ;
        RECT 5.724 0.74 5.956 0.772 ;
      LAYER M2 ;
        RECT 7.724 0.74 7.956 0.772 ;
      LAYER M3 ;
        RECT 5.18 0.504 5.22 0.756 ;
      LAYER M4 ;
        RECT 5.2 0.484 5.52 0.524 ;
      LAYER M3 ;
        RECT 5.5 0.504 5.54 0.756 ;
      LAYER M2 ;
        RECT 5.52 0.74 5.76 0.772 ;
      LAYER M2 ;
        RECT 5.92 0.74 7.84 0.772 ;
      LAYER M3 ;
        RECT 41.1 0.636 41.14 0.96 ;
      LAYER M3 ;
        RECT 40.86 0.636 40.9 0.96 ;
      LAYER M2 ;
        RECT 40.124 0.74 40.356 0.772 ;
      LAYER M2 ;
        RECT 38.124 0.74 38.356 0.772 ;
      LAYER M3 ;
        RECT 40.86 0.504 40.9 0.756 ;
      LAYER M4 ;
        RECT 40.56 0.484 40.88 0.524 ;
      LAYER M3 ;
        RECT 40.54 0.504 40.58 0.756 ;
      LAYER M2 ;
        RECT 40.32 0.74 40.56 0.772 ;
      LAYER M2 ;
        RECT 38.24 0.74 40.16 0.772 ;
      LAYER M2 ;
        RECT 15.36 -0.016 15.6 0.016 ;
      LAYER M3 ;
        RECT 15.58 0 15.62 1.008 ;
      LAYER M4 ;
        RECT 14.256 0.988 15.6 1.028 ;
      LAYER M5 ;
        RECT 14.224 1.008 14.288 5.208 ;
      LAYER M4 ;
        RECT 14.256 5.188 17.568 5.228 ;
      LAYER M5 ;
        RECT 17.536 5.208 17.6 6.72 ;
      LAYER M4 ;
        RECT 17.568 6.7 38.16 6.74 ;
      LAYER M5 ;
        RECT 38.128 0.756 38.192 6.72 ;
      LAYER M4 ;
        RECT 38.09 0.736 38.23 0.776 ;
      LAYER M3 ;
        RECT 38.14 0.651 38.18 0.861 ;
      LAYER M2 ;
        RECT 38.06 0.74 38.26 0.772 ;
    END
  END agnd
  PIN vinp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.024 -0.016 31.056 0.016 ;
      LAYER M3 ;
        RECT 31.02 17.688 31.06 18.012 ;
      LAYER M3 ;
        RECT 30.78 17.688 30.82 18.012 ;
      LAYER M1 ;
        RECT 24.544 18.276 24.576 18.348 ;
      LAYER M2 ;
        RECT 24.524 18.296 24.596 18.328 ;
      LAYER M1 ;
        RECT 21.664 18.276 21.696 18.348 ;
      LAYER M2 ;
        RECT 21.644 18.296 21.716 18.328 ;
      LAYER M2 ;
        RECT 21.68 18.296 24.56 18.328 ;
      LAYER M3 ;
        RECT 30.78 17.976 30.82 18.48 ;
      LAYER M2 ;
        RECT 27.68 18.464 30.8 18.496 ;
      LAYER M3 ;
        RECT 27.66 18.375 27.7 18.585 ;
      LAYER M4 ;
        RECT 24.624 18.46 27.68 18.5 ;
      LAYER M5 ;
        RECT 24.592 18.312 24.656 18.48 ;
      LAYER M4 ;
        RECT 24.48 18.292 24.624 18.332 ;
      LAYER M3 ;
        RECT 24.46 18.207 24.5 18.417 ;
      LAYER M2 ;
        RECT 24.38 18.296 24.58 18.328 ;
      LAYER M3 ;
        RECT 31.02 16.968 31.06 17.724 ;
      LAYER M4 ;
        RECT 31.04 16.948 31.2 16.988 ;
      LAYER M3 ;
        RECT 31.18 16.863 31.22 17.073 ;
      LAYER M2 ;
        RECT 31.2 16.952 31.68 16.984 ;
      LAYER M3 ;
        RECT 31.66 16.863 31.7 17.073 ;
      LAYER M4 ;
        RECT 31.68 16.948 32.112 16.988 ;
      LAYER M5 ;
        RECT 32.08 0.756 32.144 16.968 ;
      LAYER M4 ;
        RECT 31.68 0.736 32.112 0.776 ;
      LAYER M3 ;
        RECT 31.66 0.504 31.7 0.756 ;
      LAYER M2 ;
        RECT 31.2 0.488 31.68 0.52 ;
      LAYER M3 ;
        RECT 31.18 0.252 31.22 0.504 ;
      LAYER M4 ;
        RECT 31.04 0.232 31.2 0.272 ;
      LAYER M3 ;
        RECT 31.02 0.147 31.06 0.357 ;
      LAYER M2 ;
        RECT 30.8 0.236 31.04 0.268 ;
      LAYER M3 ;
        RECT 30.78 0 30.82 0.252 ;
      LAYER M2 ;
        RECT 30.8 -0.016 31.04 0.016 ;
    END
  END vinp
  OBS 
  LAYER M2 ;
        RECT 21.404 3.26 24.676 3.292 ;
  LAYER M3 ;
        RECT 23.02 0.468 23.06 0.876 ;
  LAYER M3 ;
        RECT 22.7 0.468 22.74 0.876 ;
  LAYER M3 ;
        RECT 23.02 5.004 23.06 5.412 ;
  LAYER M3 ;
        RECT 22.7 5.004 22.74 5.412 ;
  LAYER M2 ;
        RECT 22.044 4.184 24.036 4.216 ;
  LAYER M3 ;
        RECT 23.26 4.752 23.3 5.16 ;
  LAYER M3 ;
        RECT 22.94 4.752 22.98 5.16 ;
  LAYER M3 ;
        RECT 23.1 1.56 23.14 2.472 ;
  LAYER M2 ;
        RECT 39.644 0.824 39.876 0.856 ;
  LAYER M1 ;
        RECT 34.144 16.848 34.176 16.92 ;
  LAYER M2 ;
        RECT 34.124 16.868 34.196 16.9 ;
  LAYER M1 ;
        RECT 42.784 16.848 42.816 16.92 ;
  LAYER M2 ;
        RECT 42.764 16.868 42.836 16.9 ;
  LAYER M2 ;
        RECT 34.16 16.868 42.8 16.9 ;
  LAYER M2 ;
        RECT 39.44 0.824 39.68 0.856 ;
  LAYER M3 ;
        RECT 39.42 0.84 39.46 1.848 ;
  LAYER M4 ;
        RECT 39.12 1.828 39.44 1.868 ;
  LAYER M5 ;
        RECT 39.088 1.848 39.152 16.632 ;
  LAYER M4 ;
        RECT 39.05 16.612 39.19 16.652 ;
  LAYER M3 ;
        RECT 39.1 16.632 39.14 16.884 ;
  LAYER M2 ;
        RECT 39.02 16.868 39.22 16.9 ;
  LAYER M1 ;
        RECT 27.264 5.844 27.296 5.916 ;
  LAYER M2 ;
        RECT 27.244 5.864 27.316 5.896 ;
  LAYER M1 ;
        RECT 18.624 5.844 18.656 5.916 ;
  LAYER M2 ;
        RECT 18.604 5.864 18.676 5.896 ;
  LAYER M2 ;
        RECT 18.64 5.864 27.28 5.896 ;
  LAYER M3 ;
        RECT 23.1 1.428 23.14 1.68 ;
  LAYER M2 ;
        RECT 23.12 1.412 39.44 1.444 ;
  LAYER M3 ;
        RECT 39.42 1.323 39.46 1.533 ;
  LAYER M3 ;
        RECT 23.1 2.352 23.14 4.62 ;
  LAYER M2 ;
        RECT 23.12 4.604 23.36 4.636 ;
  LAYER M3 ;
        RECT 23.34 4.62 23.38 5.88 ;
  LAYER M2 ;
        RECT 23.26 5.864 23.46 5.896 ;
  LAYER M3 ;
        RECT 23.18 1.476 23.22 2.388 ;
  LAYER M2 ;
        RECT 6.204 0.824 6.436 0.856 ;
  LAYER M1 ;
        RECT 11.904 16.848 11.936 16.92 ;
  LAYER M2 ;
        RECT 11.884 16.868 11.956 16.9 ;
  LAYER M1 ;
        RECT 3.264 16.848 3.296 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.868 3.316 16.9 ;
  LAYER M2 ;
        RECT 3.28 16.868 11.92 16.9 ;
  LAYER M2 ;
        RECT 6.4 0.824 6.64 0.856 ;
  LAYER M3 ;
        RECT 6.62 0.84 6.66 1.848 ;
  LAYER M4 ;
        RECT 6.64 1.828 6.96 1.868 ;
  LAYER M5 ;
        RECT 6.928 1.848 6.992 16.632 ;
  LAYER M4 ;
        RECT 6.89 16.612 7.03 16.652 ;
  LAYER M3 ;
        RECT 6.94 16.632 6.98 16.884 ;
  LAYER M2 ;
        RECT 6.86 16.868 7.06 16.9 ;
  LAYER M1 ;
        RECT 24.384 6.012 24.416 6.084 ;
  LAYER M2 ;
        RECT 24.364 6.032 24.436 6.064 ;
  LAYER M1 ;
        RECT 21.504 6.012 21.536 6.084 ;
  LAYER M2 ;
        RECT 21.484 6.032 21.556 6.064 ;
  LAYER M2 ;
        RECT 21.52 6.032 24.4 6.064 ;
  LAYER M3 ;
        RECT 23.18 2.352 23.22 2.604 ;
  LAYER M4 ;
        RECT 22.464 2.584 23.2 2.624 ;
  LAYER M5 ;
        RECT 22.432 2.604 22.496 5.04 ;
  LAYER M4 ;
        RECT 7.056 5.02 22.464 5.06 ;
  LAYER M5 ;
        RECT 7.024 4.99 7.088 5.09 ;
  LAYER M5 ;
        RECT 7.024 1.848 7.088 5.04 ;
  LAYER M5 ;
        RECT 6.928 1.878 7.088 1.882 ;
  LAYER M4 ;
        RECT 21.45 5.02 21.59 5.06 ;
  LAYER M3 ;
        RECT 21.5 5.04 21.54 6.048 ;
  LAYER M2 ;
        RECT 21.42 6.032 21.62 6.064 ;
  LAYER M3 ;
        RECT 15.18 17.52 15.22 17.844 ;
  LAYER M3 ;
        RECT 15.42 17.52 15.46 17.844 ;
  LAYER M2 ;
        RECT 6.284 0.656 6.516 0.688 ;
  LAYER M2 ;
        RECT 7.164 0.656 7.396 0.688 ;
  LAYER M3 ;
        RECT 15.18 10.5 15.22 17.556 ;
  LAYER M2 ;
        RECT 8.96 10.484 15.2 10.516 ;
  LAYER M3 ;
        RECT 8.94 8.484 8.98 10.5 ;
  LAYER M4 ;
        RECT 7.392 8.464 8.96 8.504 ;
  LAYER M5 ;
        RECT 7.36 0.672 7.424 8.484 ;
  LAYER M4 ;
        RECT 6.96 0.652 7.392 0.692 ;
  LAYER M3 ;
        RECT 6.94 0.567 6.98 0.777 ;
  LAYER M2 ;
        RECT 6.96 0.656 7.2 0.688 ;
  LAYER M2 ;
        RECT 6.48 0.656 6.96 0.688 ;
  LAYER M3 ;
        RECT 30.86 17.52 30.9 17.844 ;
  LAYER M3 ;
        RECT 30.62 17.52 30.66 17.844 ;
  LAYER M2 ;
        RECT 39.564 0.656 39.796 0.688 ;
  LAYER M2 ;
        RECT 38.684 0.656 38.916 0.688 ;
  LAYER M3 ;
        RECT 30.86 10.5 30.9 17.556 ;
  LAYER M2 ;
        RECT 30.88 10.484 37.12 10.516 ;
  LAYER M3 ;
        RECT 37.1 8.484 37.14 10.5 ;
  LAYER M4 ;
        RECT 37.12 8.464 38.688 8.504 ;
  LAYER M5 ;
        RECT 38.656 0.672 38.72 8.484 ;
  LAYER M4 ;
        RECT 38.688 0.652 39.12 0.692 ;
  LAYER M3 ;
        RECT 39.1 0.567 39.14 0.777 ;
  LAYER M2 ;
        RECT 38.88 0.656 39.12 0.688 ;
  LAYER M2 ;
        RECT 39.12 0.656 39.6 0.688 ;
  LAYER M3 ;
        RECT 15.18 14.847 15.22 15.057 ;
  LAYER M4 ;
        RECT 15.2 14.932 15.52 14.972 ;
  LAYER M3 ;
        RECT 15.5 14.847 15.54 15.057 ;
  LAYER M2 ;
        RECT 15.52 14.936 30.88 14.968 ;
  LAYER M3 ;
        RECT 30.86 14.847 30.9 15.057 ;
  LAYER M3 ;
        RECT 5.1 0.468 5.14 0.792 ;
  LAYER M3 ;
        RECT 5.34 0.468 5.38 0.792 ;
  LAYER M2 ;
        RECT 5.804 0.572 6.036 0.604 ;
  LAYER M2 ;
        RECT 7.644 0.572 7.876 0.604 ;
  LAYER M3 ;
        RECT 5.34 0.336 5.38 0.588 ;
  LAYER M2 ;
        RECT 5.36 0.32 5.84 0.352 ;
  LAYER M3 ;
        RECT 5.82 0.336 5.86 0.588 ;
  LAYER M2 ;
        RECT 5.74 0.572 5.94 0.604 ;
  LAYER M2 ;
        RECT 6 0.572 7.68 0.604 ;
  LAYER M3 ;
        RECT 40.94 0.468 40.98 0.792 ;
  LAYER M3 ;
        RECT 40.7 0.468 40.74 0.792 ;
  LAYER M2 ;
        RECT 40.044 0.572 40.276 0.604 ;
  LAYER M2 ;
        RECT 38.204 0.572 38.436 0.604 ;
  LAYER M3 ;
        RECT 40.7 0.336 40.74 0.588 ;
  LAYER M2 ;
        RECT 40.24 0.32 40.72 0.352 ;
  LAYER M3 ;
        RECT 40.22 0.336 40.26 0.588 ;
  LAYER M2 ;
        RECT 40.14 0.572 40.34 0.604 ;
  LAYER M2 ;
        RECT 38.4 0.572 40.08 0.604 ;
  LAYER M2 ;
        RECT 7.84 0.572 20.32 0.604 ;
  LAYER M3 ;
        RECT 20.3 0.483 20.34 0.693 ;
  LAYER M4 ;
        RECT 20.32 0.568 38.24 0.608 ;
  LAYER M3 ;
        RECT 38.22 0.483 38.26 0.693 ;
  LAYER M2 ;
        RECT 38.14 0.572 38.34 0.604 ;
  LAYER M3 ;
        RECT 23.18 4.836 23.22 5.244 ;
  LAYER M3 ;
        RECT 22.86 4.836 22.9 5.244 ;
  LAYER M2 ;
        RECT 22.604 4.352 23.476 4.384 ;
  LAYER M3 ;
        RECT 22.86 4.368 22.9 4.872 ;
  LAYER M2 ;
        RECT 22.78 4.352 22.98 4.384 ;
  LAYER M3 ;
        RECT 23.1 4.92 23.14 5.328 ;
  LAYER M3 ;
        RECT 22.78 4.92 22.82 5.328 ;
  LAYER M2 ;
        RECT 21.964 4.52 24.116 4.552 ;
  LAYER M3 ;
        RECT 22.78 4.536 22.82 5.04 ;
  LAYER M2 ;
        RECT 22.7 4.52 22.9 4.552 ;
  LAYER M3 ;
        RECT 22.94 1.728 22.98 2.64 ;
  LAYER M2 ;
        RECT 21.484 3.092 24.116 3.124 ;
  LAYER M3 ;
        RECT 22.94 2.604 22.98 3.108 ;
  LAYER M2 ;
        RECT 22.86 3.092 23.06 3.124 ;
  LAYER M3 ;
        RECT 22.86 1.812 22.9 2.724 ;
  LAYER M3 ;
        RECT 23.1 0.384 23.14 0.792 ;
  LAYER M3 ;
        RECT 22.78 0.384 22.82 0.792 ;
  LAYER M3 ;
        RECT 22.86 0.924 22.9 1.932 ;
  LAYER M2 ;
        RECT 22.88 0.908 23.12 0.94 ;
  LAYER M3 ;
        RECT 23.1 0.672 23.14 0.924 ;
  LAYER M3 ;
        RECT 23.02 1.644 23.06 2.556 ;
  LAYER M2 ;
        RECT 22.124 2.924 24.756 2.956 ;
  LAYER M3 ;
        RECT 23.02 2.436 23.06 2.94 ;
  LAYER M2 ;
        RECT 22.94 2.924 23.14 2.956 ;
  LAYER M1 ;
        RECT 23.344 4.752 23.376 5.412 ;
  LAYER M1 ;
        RECT 23.424 4.752 23.456 5.412 ;
  LAYER M1 ;
        RECT 23.264 4.752 23.296 5.412 ;
  LAYER M1 ;
        RECT 22.704 4.752 22.736 5.412 ;
  LAYER M1 ;
        RECT 22.784 4.752 22.816 5.412 ;
  LAYER M1 ;
        RECT 22.624 4.752 22.656 5.412 ;
  LAYER M2 ;
        RECT 22.764 4.772 23.476 4.804 ;
  LAYER M2 ;
        RECT 22.764 5.108 23.476 5.14 ;
  LAYER M2 ;
        RECT 22.844 4.856 23.316 4.888 ;
  LAYER M2 ;
        RECT 22.844 5.192 23.316 5.224 ;
  LAYER M2 ;
        RECT 22.604 4.94 23.156 4.972 ;
  LAYER M2 ;
        RECT 22.604 5.276 23.156 5.308 ;
  LAYER M2 ;
        RECT 22.684 5.024 23.396 5.056 ;
  LAYER M2 ;
        RECT 22.684 5.36 23.396 5.392 ;
  LAYER M1 ;
        RECT 21.424 2.064 21.456 2.724 ;
  LAYER M1 ;
        RECT 21.424 1.224 21.456 1.884 ;
  LAYER M1 ;
        RECT 21.344 2.064 21.376 2.724 ;
  LAYER M1 ;
        RECT 21.344 1.224 21.376 1.884 ;
  LAYER M1 ;
        RECT 21.504 2.064 21.536 2.724 ;
  LAYER M1 ;
        RECT 21.504 1.224 21.536 1.884 ;
  LAYER M1 ;
        RECT 22.064 2.064 22.096 2.724 ;
  LAYER M1 ;
        RECT 22.064 1.224 22.096 1.884 ;
  LAYER M1 ;
        RECT 21.984 2.064 22.016 2.724 ;
  LAYER M1 ;
        RECT 21.984 1.224 22.016 1.884 ;
  LAYER M1 ;
        RECT 22.144 2.064 22.176 2.724 ;
  LAYER M1 ;
        RECT 22.144 1.224 22.176 1.884 ;
  LAYER M1 ;
        RECT 22.704 2.064 22.736 2.724 ;
  LAYER M1 ;
        RECT 22.704 1.224 22.736 1.884 ;
  LAYER M1 ;
        RECT 22.624 2.064 22.656 2.724 ;
  LAYER M1 ;
        RECT 22.624 1.224 22.656 1.884 ;
  LAYER M1 ;
        RECT 22.784 2.064 22.816 2.724 ;
  LAYER M1 ;
        RECT 22.784 1.224 22.816 1.884 ;
  LAYER M1 ;
        RECT 23.344 2.064 23.376 2.724 ;
  LAYER M1 ;
        RECT 23.344 1.224 23.376 1.884 ;
  LAYER M1 ;
        RECT 23.264 2.064 23.296 2.724 ;
  LAYER M1 ;
        RECT 23.264 1.224 23.296 1.884 ;
  LAYER M1 ;
        RECT 23.424 2.064 23.456 2.724 ;
  LAYER M1 ;
        RECT 23.424 1.224 23.456 1.884 ;
  LAYER M1 ;
        RECT 23.984 2.064 24.016 2.724 ;
  LAYER M1 ;
        RECT 23.984 1.224 24.016 1.884 ;
  LAYER M1 ;
        RECT 23.904 2.064 23.936 2.724 ;
  LAYER M1 ;
        RECT 23.904 1.224 23.936 1.884 ;
  LAYER M1 ;
        RECT 24.064 2.064 24.096 2.724 ;
  LAYER M1 ;
        RECT 24.064 1.224 24.096 1.884 ;
  LAYER M1 ;
        RECT 24.624 2.064 24.656 2.724 ;
  LAYER M1 ;
        RECT 24.624 1.224 24.656 1.884 ;
  LAYER M1 ;
        RECT 24.544 2.064 24.576 2.724 ;
  LAYER M1 ;
        RECT 24.544 1.224 24.576 1.884 ;
  LAYER M1 ;
        RECT 24.704 2.064 24.736 2.724 ;
  LAYER M1 ;
        RECT 24.704 1.224 24.736 1.884 ;
  LAYER M2 ;
        RECT 21.324 2.672 24.596 2.704 ;
  LAYER M2 ;
        RECT 21.484 2.588 24.116 2.62 ;
  LAYER M2 ;
        RECT 22.124 2.504 24.756 2.536 ;
  LAYER M2 ;
        RECT 21.404 2.42 24.036 2.452 ;
  LAYER M2 ;
        RECT 22.044 2.336 24.676 2.368 ;
  LAYER M2 ;
        RECT 21.324 1.832 24.596 1.864 ;
  LAYER M2 ;
        RECT 22.124 1.748 24.756 1.78 ;
  LAYER M2 ;
        RECT 21.484 1.664 24.116 1.696 ;
  LAYER M2 ;
        RECT 22.044 1.58 24.676 1.612 ;
  LAYER M2 ;
        RECT 21.404 1.496 24.036 1.528 ;
  LAYER M1 ;
        RECT 25.264 0.216 25.296 0.876 ;
  LAYER M1 ;
        RECT 25.344 0.216 25.376 0.876 ;
  LAYER M1 ;
        RECT 25.184 0.216 25.216 0.876 ;
  LAYER M1 ;
        RECT 24.624 0.216 24.656 0.876 ;
  LAYER M1 ;
        RECT 24.704 0.216 24.736 0.876 ;
  LAYER M1 ;
        RECT 24.544 0.216 24.576 0.876 ;
  LAYER M1 ;
        RECT 23.984 0.216 24.016 0.876 ;
  LAYER M1 ;
        RECT 24.064 0.216 24.096 0.876 ;
  LAYER M1 ;
        RECT 23.904 0.216 23.936 0.876 ;
  LAYER M1 ;
        RECT 23.344 0.216 23.376 0.876 ;
  LAYER M1 ;
        RECT 23.424 0.216 23.456 0.876 ;
  LAYER M1 ;
        RECT 23.264 0.216 23.296 0.876 ;
  LAYER M1 ;
        RECT 22.704 0.216 22.736 0.876 ;
  LAYER M1 ;
        RECT 22.784 0.216 22.816 0.876 ;
  LAYER M1 ;
        RECT 22.624 0.216 22.656 0.876 ;
  LAYER M1 ;
        RECT 22.064 0.216 22.096 0.876 ;
  LAYER M1 ;
        RECT 22.144 0.216 22.176 0.876 ;
  LAYER M1 ;
        RECT 21.984 0.216 22.016 0.876 ;
  LAYER M1 ;
        RECT 21.424 0.216 21.456 0.876 ;
  LAYER M1 ;
        RECT 21.504 0.216 21.536 0.876 ;
  LAYER M1 ;
        RECT 21.344 0.216 21.376 0.876 ;
  LAYER M1 ;
        RECT 20.784 0.216 20.816 0.876 ;
  LAYER M1 ;
        RECT 20.864 0.216 20.896 0.876 ;
  LAYER M1 ;
        RECT 20.704 0.216 20.736 0.876 ;
  LAYER M2 ;
        RECT 20.844 0.236 25.396 0.268 ;
  LAYER M2 ;
        RECT 20.844 0.572 25.396 0.604 ;
  LAYER M2 ;
        RECT 22.604 0.32 23.396 0.352 ;
  LAYER M2 ;
        RECT 22.604 0.656 23.396 0.688 ;
  LAYER M2 ;
        RECT 20.684 0.404 25.236 0.436 ;
  LAYER M2 ;
        RECT 20.684 0.74 25.236 0.772 ;
  LAYER M2 ;
        RECT 20.764 0.488 25.316 0.52 ;
  LAYER M2 ;
        RECT 20.764 0.824 25.316 0.856 ;
  LAYER M1 ;
        RECT 22.064 3.912 22.096 4.572 ;
  LAYER M1 ;
        RECT 21.984 3.912 22.016 4.572 ;
  LAYER M1 ;
        RECT 22.144 3.912 22.176 4.572 ;
  LAYER M1 ;
        RECT 22.704 3.912 22.736 4.572 ;
  LAYER M1 ;
        RECT 22.624 3.912 22.656 4.572 ;
  LAYER M1 ;
        RECT 22.784 3.912 22.816 4.572 ;
  LAYER M1 ;
        RECT 23.344 3.912 23.376 4.572 ;
  LAYER M1 ;
        RECT 23.424 3.912 23.456 4.572 ;
  LAYER M1 ;
        RECT 23.264 3.912 23.296 4.572 ;
  LAYER M1 ;
        RECT 23.984 3.912 24.016 4.572 ;
  LAYER M1 ;
        RECT 24.064 3.912 24.096 4.572 ;
  LAYER M1 ;
        RECT 23.904 3.912 23.936 4.572 ;
  LAYER M1 ;
        RECT 24.624 2.904 24.656 3.564 ;
  LAYER M1 ;
        RECT 24.704 2.904 24.736 3.564 ;
  LAYER M1 ;
        RECT 24.544 2.904 24.576 3.564 ;
  LAYER M1 ;
        RECT 23.984 2.904 24.016 3.564 ;
  LAYER M1 ;
        RECT 24.064 2.904 24.096 3.564 ;
  LAYER M1 ;
        RECT 23.904 2.904 23.936 3.564 ;
  LAYER M1 ;
        RECT 23.344 2.904 23.376 3.564 ;
  LAYER M1 ;
        RECT 23.424 2.904 23.456 3.564 ;
  LAYER M1 ;
        RECT 23.264 2.904 23.296 3.564 ;
  LAYER M1 ;
        RECT 22.704 2.904 22.736 3.564 ;
  LAYER M1 ;
        RECT 22.784 2.904 22.816 3.564 ;
  LAYER M1 ;
        RECT 22.624 2.904 22.656 3.564 ;
  LAYER M1 ;
        RECT 22.064 2.904 22.096 3.564 ;
  LAYER M1 ;
        RECT 22.144 2.904 22.176 3.564 ;
  LAYER M1 ;
        RECT 21.984 2.904 22.016 3.564 ;
  LAYER M1 ;
        RECT 21.424 2.904 21.456 3.564 ;
  LAYER M1 ;
        RECT 21.504 2.904 21.536 3.564 ;
  LAYER M1 ;
        RECT 21.344 2.904 21.376 3.564 ;
  LAYER M1 ;
        RECT 6.224 29.7 6.256 29.772 ;
  LAYER M2 ;
        RECT 6.204 29.72 6.276 29.752 ;
  LAYER M1 ;
        RECT 9.104 29.7 9.136 29.772 ;
  LAYER M2 ;
        RECT 9.084 29.72 9.156 29.752 ;
  LAYER M2 ;
        RECT 6.24 29.72 9.12 29.752 ;
  LAYER M2 ;
        RECT 5.884 0.908 6.596 0.94 ;
  LAYER M1 ;
        RECT 9.024 16.68 9.056 16.752 ;
  LAYER M2 ;
        RECT 9.004 16.7 9.076 16.732 ;
  LAYER M1 ;
        RECT 6.144 16.68 6.176 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.7 6.196 16.732 ;
  LAYER M2 ;
        RECT 6.16 16.7 9.04 16.732 ;
  LAYER M2 ;
        RECT 8.3 29.72 8.5 29.752 ;
  LAYER M3 ;
        RECT 8.38 29.484 8.42 29.736 ;
  LAYER M4 ;
        RECT 8.33 29.464 8.47 29.504 ;
  LAYER M5 ;
        RECT 8.368 16.968 8.432 29.484 ;
  LAYER M4 ;
        RECT 8.33 16.948 8.47 16.988 ;
  LAYER M3 ;
        RECT 8.38 16.716 8.42 16.968 ;
  LAYER M2 ;
        RECT 8.3 16.7 8.5 16.732 ;
  LAYER M2 ;
        RECT 6.14 16.7 6.34 16.732 ;
  LAYER M3 ;
        RECT 6.22 1.596 6.26 16.716 ;
  LAYER M4 ;
        RECT 6.17 1.576 6.31 1.616 ;
  LAYER M5 ;
        RECT 6.208 1.428 6.272 1.596 ;
  LAYER M4 ;
        RECT 6.17 1.408 6.31 1.448 ;
  LAYER M3 ;
        RECT 6.22 0.924 6.26 1.428 ;
  LAYER M2 ;
        RECT 6.14 0.908 6.34 0.94 ;
  LAYER M1 ;
        RECT 6.064 17.436 6.096 17.508 ;
  LAYER M2 ;
        RECT 6.044 17.456 6.116 17.488 ;
  LAYER M1 ;
        RECT 8.944 17.436 8.976 17.508 ;
  LAYER M2 ;
        RECT 8.924 17.456 8.996 17.488 ;
  LAYER M2 ;
        RECT 6.08 17.456 8.96 17.488 ;
  LAYER M3 ;
        RECT 5.02 0.552 5.06 0.876 ;
  LAYER M3 ;
        RECT 5.26 0.552 5.3 0.876 ;
  LAYER M3 ;
        RECT 15.1 17.604 15.14 17.928 ;
  LAYER M3 ;
        RECT 15.34 17.604 15.38 17.928 ;
  LAYER M2 ;
        RECT 8.96 17.456 14.96 17.488 ;
  LAYER M3 ;
        RECT 14.94 17.367 14.98 17.577 ;
  LAYER M4 ;
        RECT 14.96 17.452 15.12 17.492 ;
  LAYER M3 ;
        RECT 15.1 17.472 15.14 17.724 ;
  LAYER M2 ;
        RECT 5.98 17.456 6.18 17.488 ;
  LAYER M3 ;
        RECT 6.06 0.84 6.1 17.472 ;
  LAYER M4 ;
        RECT 5.28 0.82 6.08 0.86 ;
  LAYER M3 ;
        RECT 5.26 0.735 5.3 0.945 ;
  LAYER M2 ;
        RECT 7.084 0.908 7.796 0.94 ;
  LAYER M1 ;
        RECT 8.864 1.476 8.896 1.548 ;
  LAYER M2 ;
        RECT 8.844 1.496 8.916 1.528 ;
  LAYER M1 ;
        RECT 5.984 1.476 6.016 1.548 ;
  LAYER M2 ;
        RECT 5.964 1.496 6.036 1.528 ;
  LAYER M2 ;
        RECT 6 1.496 8.88 1.528 ;
  LAYER M2 ;
        RECT 7.42 0.908 7.62 0.94 ;
  LAYER M3 ;
        RECT 7.5 0.924 7.54 1.428 ;
  LAYER M4 ;
        RECT 7.52 1.408 7.68 1.448 ;
  LAYER M5 ;
        RECT 7.648 1.42 7.712 1.52 ;
  LAYER M4 ;
        RECT 7.61 1.492 7.75 1.532 ;
  LAYER M3 ;
        RECT 7.66 1.407 7.7 1.617 ;
  LAYER M2 ;
        RECT 7.58 1.496 7.78 1.528 ;
  LAYER M1 ;
        RECT 8.784 20.88 8.816 20.952 ;
  LAYER M2 ;
        RECT 8.764 20.9 8.836 20.932 ;
  LAYER M2 ;
        RECT 6.08 20.9 8.8 20.932 ;
  LAYER M1 ;
        RECT 6.064 20.88 6.096 20.952 ;
  LAYER M2 ;
        RECT 6.044 20.9 6.116 20.932 ;
  LAYER M1 ;
        RECT 8.784 23.82 8.816 23.892 ;
  LAYER M2 ;
        RECT 8.764 23.84 8.836 23.872 ;
  LAYER M2 ;
        RECT 6.08 23.84 8.8 23.872 ;
  LAYER M1 ;
        RECT 6.064 23.82 6.096 23.892 ;
  LAYER M2 ;
        RECT 6.044 23.84 6.116 23.872 ;
  LAYER M1 ;
        RECT 5.904 20.88 5.936 20.952 ;
  LAYER M2 ;
        RECT 5.884 20.9 5.956 20.932 ;
  LAYER M1 ;
        RECT 5.904 20.748 5.936 20.916 ;
  LAYER M1 ;
        RECT 5.904 20.712 5.936 20.784 ;
  LAYER M2 ;
        RECT 5.884 20.732 5.956 20.764 ;
  LAYER M2 ;
        RECT 5.92 20.732 6.08 20.764 ;
  LAYER M1 ;
        RECT 6.064 20.712 6.096 20.784 ;
  LAYER M2 ;
        RECT 6.044 20.732 6.116 20.764 ;
  LAYER M1 ;
        RECT 5.904 23.82 5.936 23.892 ;
  LAYER M2 ;
        RECT 5.884 23.84 5.956 23.872 ;
  LAYER M1 ;
        RECT 5.904 23.688 5.936 23.856 ;
  LAYER M1 ;
        RECT 5.904 23.652 5.936 23.724 ;
  LAYER M2 ;
        RECT 5.884 23.672 5.956 23.704 ;
  LAYER M2 ;
        RECT 5.92 23.672 6.08 23.704 ;
  LAYER M1 ;
        RECT 6.064 23.652 6.096 23.724 ;
  LAYER M2 ;
        RECT 6.044 23.672 6.116 23.704 ;
  LAYER M1 ;
        RECT 6.064 17.436 6.096 17.508 ;
  LAYER M2 ;
        RECT 6.044 17.456 6.116 17.488 ;
  LAYER M1 ;
        RECT 6.064 17.472 6.096 17.64 ;
  LAYER M1 ;
        RECT 6.064 17.64 6.096 23.856 ;
  LAYER M1 ;
        RECT 11.664 23.82 11.696 23.892 ;
  LAYER M2 ;
        RECT 11.644 23.84 11.716 23.872 ;
  LAYER M2 ;
        RECT 8.96 23.84 11.68 23.872 ;
  LAYER M1 ;
        RECT 8.944 23.82 8.976 23.892 ;
  LAYER M2 ;
        RECT 8.924 23.84 8.996 23.872 ;
  LAYER M1 ;
        RECT 11.664 20.88 11.696 20.952 ;
  LAYER M2 ;
        RECT 11.644 20.9 11.716 20.932 ;
  LAYER M2 ;
        RECT 8.96 20.9 11.68 20.932 ;
  LAYER M1 ;
        RECT 8.944 20.88 8.976 20.952 ;
  LAYER M2 ;
        RECT 8.924 20.9 8.996 20.932 ;
  LAYER M1 ;
        RECT 8.944 17.436 8.976 17.508 ;
  LAYER M2 ;
        RECT 8.924 17.456 8.996 17.488 ;
  LAYER M1 ;
        RECT 8.944 17.472 8.976 17.64 ;
  LAYER M1 ;
        RECT 8.944 17.64 8.976 23.856 ;
  LAYER M2 ;
        RECT 6.08 17.456 8.96 17.488 ;
  LAYER M1 ;
        RECT 3.024 17.94 3.056 18.012 ;
  LAYER M2 ;
        RECT 3.004 17.96 3.076 17.992 ;
  LAYER M1 ;
        RECT 3.024 17.808 3.056 17.976 ;
  LAYER M1 ;
        RECT 3.024 17.772 3.056 17.844 ;
  LAYER M2 ;
        RECT 3.004 17.792 3.076 17.824 ;
  LAYER M2 ;
        RECT 3.04 17.792 3.2 17.824 ;
  LAYER M1 ;
        RECT 3.184 17.772 3.216 17.844 ;
  LAYER M2 ;
        RECT 3.164 17.792 3.236 17.824 ;
  LAYER M1 ;
        RECT 3.024 20.88 3.056 20.952 ;
  LAYER M2 ;
        RECT 3.004 20.9 3.076 20.932 ;
  LAYER M1 ;
        RECT 3.024 20.748 3.056 20.916 ;
  LAYER M1 ;
        RECT 3.024 20.712 3.056 20.784 ;
  LAYER M2 ;
        RECT 3.004 20.732 3.076 20.764 ;
  LAYER M2 ;
        RECT 3.04 20.732 3.2 20.764 ;
  LAYER M1 ;
        RECT 3.184 20.712 3.216 20.784 ;
  LAYER M2 ;
        RECT 3.164 20.732 3.236 20.764 ;
  LAYER M1 ;
        RECT 3.024 23.82 3.056 23.892 ;
  LAYER M2 ;
        RECT 3.004 23.84 3.076 23.872 ;
  LAYER M1 ;
        RECT 3.024 23.688 3.056 23.856 ;
  LAYER M1 ;
        RECT 3.024 23.652 3.056 23.724 ;
  LAYER M2 ;
        RECT 3.004 23.672 3.076 23.704 ;
  LAYER M2 ;
        RECT 3.04 23.672 3.2 23.704 ;
  LAYER M1 ;
        RECT 3.184 23.652 3.216 23.724 ;
  LAYER M2 ;
        RECT 3.164 23.672 3.236 23.704 ;
  LAYER M1 ;
        RECT 3.024 26.76 3.056 26.832 ;
  LAYER M2 ;
        RECT 3.004 26.78 3.076 26.812 ;
  LAYER M1 ;
        RECT 3.024 26.628 3.056 26.796 ;
  LAYER M1 ;
        RECT 3.024 26.592 3.056 26.664 ;
  LAYER M2 ;
        RECT 3.004 26.612 3.076 26.644 ;
  LAYER M2 ;
        RECT 3.04 26.612 3.2 26.644 ;
  LAYER M1 ;
        RECT 3.184 26.592 3.216 26.664 ;
  LAYER M2 ;
        RECT 3.164 26.612 3.236 26.644 ;
  LAYER M1 ;
        RECT 5.904 17.94 5.936 18.012 ;
  LAYER M2 ;
        RECT 5.884 17.96 5.956 17.992 ;
  LAYER M2 ;
        RECT 3.2 17.96 5.92 17.992 ;
  LAYER M1 ;
        RECT 3.184 17.94 3.216 18.012 ;
  LAYER M2 ;
        RECT 3.164 17.96 3.236 17.992 ;
  LAYER M1 ;
        RECT 5.904 26.76 5.936 26.832 ;
  LAYER M2 ;
        RECT 5.884 26.78 5.956 26.812 ;
  LAYER M2 ;
        RECT 3.2 26.78 5.92 26.812 ;
  LAYER M1 ;
        RECT 3.184 26.76 3.216 26.832 ;
  LAYER M2 ;
        RECT 3.164 26.78 3.236 26.812 ;
  LAYER M1 ;
        RECT 3.184 17.268 3.216 17.34 ;
  LAYER M2 ;
        RECT 3.164 17.288 3.236 17.32 ;
  LAYER M1 ;
        RECT 3.184 17.304 3.216 17.64 ;
  LAYER M1 ;
        RECT 3.184 17.64 3.216 26.796 ;
  LAYER M1 ;
        RECT 11.664 17.94 11.696 18.012 ;
  LAYER M2 ;
        RECT 11.644 17.96 11.716 17.992 ;
  LAYER M1 ;
        RECT 11.664 17.808 11.696 17.976 ;
  LAYER M1 ;
        RECT 11.664 17.772 11.696 17.844 ;
  LAYER M2 ;
        RECT 11.644 17.792 11.716 17.824 ;
  LAYER M2 ;
        RECT 11.68 17.792 11.84 17.824 ;
  LAYER M1 ;
        RECT 11.824 17.772 11.856 17.844 ;
  LAYER M2 ;
        RECT 11.804 17.792 11.876 17.824 ;
  LAYER M1 ;
        RECT 11.664 26.76 11.696 26.832 ;
  LAYER M2 ;
        RECT 11.644 26.78 11.716 26.812 ;
  LAYER M1 ;
        RECT 11.664 26.628 11.696 26.796 ;
  LAYER M1 ;
        RECT 11.664 26.592 11.696 26.664 ;
  LAYER M2 ;
        RECT 11.644 26.612 11.716 26.644 ;
  LAYER M2 ;
        RECT 11.68 26.612 11.84 26.644 ;
  LAYER M1 ;
        RECT 11.824 26.592 11.856 26.664 ;
  LAYER M2 ;
        RECT 11.804 26.612 11.876 26.644 ;
  LAYER M1 ;
        RECT 14.544 17.94 14.576 18.012 ;
  LAYER M2 ;
        RECT 14.524 17.96 14.596 17.992 ;
  LAYER M2 ;
        RECT 11.84 17.96 14.56 17.992 ;
  LAYER M1 ;
        RECT 11.824 17.94 11.856 18.012 ;
  LAYER M2 ;
        RECT 11.804 17.96 11.876 17.992 ;
  LAYER M1 ;
        RECT 14.544 20.88 14.576 20.952 ;
  LAYER M2 ;
        RECT 14.524 20.9 14.596 20.932 ;
  LAYER M2 ;
        RECT 11.84 20.9 14.56 20.932 ;
  LAYER M1 ;
        RECT 11.824 20.88 11.856 20.952 ;
  LAYER M2 ;
        RECT 11.804 20.9 11.876 20.932 ;
  LAYER M1 ;
        RECT 14.544 23.82 14.576 23.892 ;
  LAYER M2 ;
        RECT 14.524 23.84 14.596 23.872 ;
  LAYER M2 ;
        RECT 11.84 23.84 14.56 23.872 ;
  LAYER M1 ;
        RECT 11.824 23.82 11.856 23.892 ;
  LAYER M2 ;
        RECT 11.804 23.84 11.876 23.872 ;
  LAYER M1 ;
        RECT 14.544 26.76 14.576 26.832 ;
  LAYER M2 ;
        RECT 14.524 26.78 14.596 26.812 ;
  LAYER M2 ;
        RECT 11.84 26.78 14.56 26.812 ;
  LAYER M1 ;
        RECT 11.824 26.76 11.856 26.832 ;
  LAYER M2 ;
        RECT 11.804 26.78 11.876 26.812 ;
  LAYER M1 ;
        RECT 11.824 17.268 11.856 17.34 ;
  LAYER M2 ;
        RECT 11.804 17.288 11.876 17.32 ;
  LAYER M1 ;
        RECT 11.824 17.304 11.856 17.64 ;
  LAYER M1 ;
        RECT 11.824 17.64 11.856 26.796 ;
  LAYER M2 ;
        RECT 3.2 17.288 11.84 17.32 ;
  LAYER M1 ;
        RECT 8.784 26.76 8.816 26.832 ;
  LAYER M2 ;
        RECT 8.764 26.78 8.836 26.812 ;
  LAYER M2 ;
        RECT 5.92 26.78 8.8 26.812 ;
  LAYER M1 ;
        RECT 5.904 26.76 5.936 26.832 ;
  LAYER M2 ;
        RECT 5.884 26.78 5.956 26.812 ;
  LAYER M1 ;
        RECT 8.784 17.94 8.816 18.012 ;
  LAYER M2 ;
        RECT 8.764 17.96 8.836 17.992 ;
  LAYER M2 ;
        RECT 8.8 17.96 11.68 17.992 ;
  LAYER M1 ;
        RECT 11.664 17.94 11.696 18.012 ;
  LAYER M2 ;
        RECT 11.644 17.96 11.716 17.992 ;
  LAYER M1 ;
        RECT 6.384 23.316 6.416 23.388 ;
  LAYER M2 ;
        RECT 6.364 23.336 6.436 23.368 ;
  LAYER M2 ;
        RECT 6.24 23.336 6.4 23.368 ;
  LAYER M1 ;
        RECT 6.224 23.316 6.256 23.388 ;
  LAYER M2 ;
        RECT 6.204 23.336 6.276 23.368 ;
  LAYER M1 ;
        RECT 6.384 26.256 6.416 26.328 ;
  LAYER M2 ;
        RECT 6.364 26.276 6.436 26.308 ;
  LAYER M2 ;
        RECT 6.24 26.276 6.4 26.308 ;
  LAYER M1 ;
        RECT 6.224 26.256 6.256 26.328 ;
  LAYER M2 ;
        RECT 6.204 26.276 6.276 26.308 ;
  LAYER M1 ;
        RECT 3.504 23.316 3.536 23.388 ;
  LAYER M2 ;
        RECT 3.484 23.336 3.556 23.368 ;
  LAYER M1 ;
        RECT 3.504 23.352 3.536 23.52 ;
  LAYER M1 ;
        RECT 3.504 23.484 3.536 23.556 ;
  LAYER M2 ;
        RECT 3.484 23.504 3.556 23.536 ;
  LAYER M2 ;
        RECT 3.52 23.504 6.24 23.536 ;
  LAYER M1 ;
        RECT 6.224 23.484 6.256 23.556 ;
  LAYER M2 ;
        RECT 6.204 23.504 6.276 23.536 ;
  LAYER M1 ;
        RECT 3.504 26.256 3.536 26.328 ;
  LAYER M2 ;
        RECT 3.484 26.276 3.556 26.308 ;
  LAYER M1 ;
        RECT 3.504 26.292 3.536 26.46 ;
  LAYER M1 ;
        RECT 3.504 26.424 3.536 26.496 ;
  LAYER M2 ;
        RECT 3.484 26.444 3.556 26.476 ;
  LAYER M2 ;
        RECT 3.52 26.444 6.24 26.476 ;
  LAYER M1 ;
        RECT 6.224 26.424 6.256 26.496 ;
  LAYER M2 ;
        RECT 6.204 26.444 6.276 26.476 ;
  LAYER M1 ;
        RECT 6.224 29.7 6.256 29.772 ;
  LAYER M2 ;
        RECT 6.204 29.72 6.276 29.752 ;
  LAYER M1 ;
        RECT 6.224 29.568 6.256 29.736 ;
  LAYER M1 ;
        RECT 6.224 23.352 6.256 29.568 ;
  LAYER M1 ;
        RECT 9.264 26.256 9.296 26.328 ;
  LAYER M2 ;
        RECT 9.244 26.276 9.316 26.308 ;
  LAYER M2 ;
        RECT 9.12 26.276 9.28 26.308 ;
  LAYER M1 ;
        RECT 9.104 26.256 9.136 26.328 ;
  LAYER M2 ;
        RECT 9.084 26.276 9.156 26.308 ;
  LAYER M1 ;
        RECT 9.264 23.316 9.296 23.388 ;
  LAYER M2 ;
        RECT 9.244 23.336 9.316 23.368 ;
  LAYER M2 ;
        RECT 9.12 23.336 9.28 23.368 ;
  LAYER M1 ;
        RECT 9.104 23.316 9.136 23.388 ;
  LAYER M2 ;
        RECT 9.084 23.336 9.156 23.368 ;
  LAYER M1 ;
        RECT 9.104 29.7 9.136 29.772 ;
  LAYER M2 ;
        RECT 9.084 29.72 9.156 29.752 ;
  LAYER M1 ;
        RECT 9.104 29.568 9.136 29.736 ;
  LAYER M1 ;
        RECT 9.104 23.352 9.136 29.568 ;
  LAYER M2 ;
        RECT 6.24 29.72 9.12 29.752 ;
  LAYER M1 ;
        RECT 0.624 20.376 0.656 20.448 ;
  LAYER M2 ;
        RECT 0.604 20.396 0.676 20.428 ;
  LAYER M2 ;
        RECT 0.32 20.396 0.64 20.428 ;
  LAYER M1 ;
        RECT 0.304 20.376 0.336 20.448 ;
  LAYER M2 ;
        RECT 0.284 20.396 0.356 20.428 ;
  LAYER M1 ;
        RECT 0.624 23.316 0.656 23.388 ;
  LAYER M2 ;
        RECT 0.604 23.336 0.676 23.368 ;
  LAYER M2 ;
        RECT 0.32 23.336 0.64 23.368 ;
  LAYER M1 ;
        RECT 0.304 23.316 0.336 23.388 ;
  LAYER M2 ;
        RECT 0.284 23.336 0.356 23.368 ;
  LAYER M1 ;
        RECT 0.624 26.256 0.656 26.328 ;
  LAYER M2 ;
        RECT 0.604 26.276 0.676 26.308 ;
  LAYER M2 ;
        RECT 0.32 26.276 0.64 26.308 ;
  LAYER M1 ;
        RECT 0.304 26.256 0.336 26.328 ;
  LAYER M2 ;
        RECT 0.284 26.276 0.356 26.308 ;
  LAYER M1 ;
        RECT 0.624 29.196 0.656 29.268 ;
  LAYER M2 ;
        RECT 0.604 29.216 0.676 29.248 ;
  LAYER M2 ;
        RECT 0.32 29.216 0.64 29.248 ;
  LAYER M1 ;
        RECT 0.304 29.196 0.336 29.268 ;
  LAYER M2 ;
        RECT 0.284 29.216 0.356 29.248 ;
  LAYER M1 ;
        RECT 0.304 29.868 0.336 29.94 ;
  LAYER M2 ;
        RECT 0.284 29.888 0.356 29.92 ;
  LAYER M1 ;
        RECT 0.304 29.568 0.336 29.904 ;
  LAYER M1 ;
        RECT 0.304 20.412 0.336 29.568 ;
  LAYER M1 ;
        RECT 12.144 20.376 12.176 20.448 ;
  LAYER M2 ;
        RECT 12.124 20.396 12.196 20.428 ;
  LAYER M1 ;
        RECT 12.144 20.412 12.176 20.58 ;
  LAYER M1 ;
        RECT 12.144 20.544 12.176 20.616 ;
  LAYER M2 ;
        RECT 12.124 20.564 12.196 20.596 ;
  LAYER M2 ;
        RECT 12.16 20.564 14.72 20.596 ;
  LAYER M1 ;
        RECT 14.704 20.544 14.736 20.616 ;
  LAYER M2 ;
        RECT 14.684 20.564 14.756 20.596 ;
  LAYER M1 ;
        RECT 12.144 23.316 12.176 23.388 ;
  LAYER M2 ;
        RECT 12.124 23.336 12.196 23.368 ;
  LAYER M1 ;
        RECT 12.144 23.352 12.176 23.52 ;
  LAYER M1 ;
        RECT 12.144 23.484 12.176 23.556 ;
  LAYER M2 ;
        RECT 12.124 23.504 12.196 23.536 ;
  LAYER M2 ;
        RECT 12.16 23.504 14.72 23.536 ;
  LAYER M1 ;
        RECT 14.704 23.484 14.736 23.556 ;
  LAYER M2 ;
        RECT 14.684 23.504 14.756 23.536 ;
  LAYER M1 ;
        RECT 12.144 26.256 12.176 26.328 ;
  LAYER M2 ;
        RECT 12.124 26.276 12.196 26.308 ;
  LAYER M1 ;
        RECT 12.144 26.292 12.176 26.46 ;
  LAYER M1 ;
        RECT 12.144 26.424 12.176 26.496 ;
  LAYER M2 ;
        RECT 12.124 26.444 12.196 26.476 ;
  LAYER M2 ;
        RECT 12.16 26.444 14.72 26.476 ;
  LAYER M1 ;
        RECT 14.704 26.424 14.736 26.496 ;
  LAYER M2 ;
        RECT 14.684 26.444 14.756 26.476 ;
  LAYER M1 ;
        RECT 12.144 29.196 12.176 29.268 ;
  LAYER M2 ;
        RECT 12.124 29.216 12.196 29.248 ;
  LAYER M1 ;
        RECT 12.144 29.232 12.176 29.4 ;
  LAYER M1 ;
        RECT 12.144 29.364 12.176 29.436 ;
  LAYER M2 ;
        RECT 12.124 29.384 12.196 29.416 ;
  LAYER M2 ;
        RECT 12.16 29.384 14.72 29.416 ;
  LAYER M1 ;
        RECT 14.704 29.364 14.736 29.436 ;
  LAYER M2 ;
        RECT 14.684 29.384 14.756 29.416 ;
  LAYER M1 ;
        RECT 14.704 29.868 14.736 29.94 ;
  LAYER M2 ;
        RECT 14.684 29.888 14.756 29.92 ;
  LAYER M1 ;
        RECT 14.704 29.568 14.736 29.904 ;
  LAYER M1 ;
        RECT 14.704 20.58 14.736 29.568 ;
  LAYER M2 ;
        RECT 0.32 29.888 14.72 29.92 ;
  LAYER M1 ;
        RECT 3.504 20.376 3.536 20.448 ;
  LAYER M2 ;
        RECT 3.484 20.396 3.556 20.428 ;
  LAYER M2 ;
        RECT 0.64 20.396 3.52 20.428 ;
  LAYER M1 ;
        RECT 0.624 20.376 0.656 20.448 ;
  LAYER M2 ;
        RECT 0.604 20.396 0.676 20.428 ;
  LAYER M1 ;
        RECT 3.504 29.196 3.536 29.268 ;
  LAYER M2 ;
        RECT 3.484 29.216 3.556 29.248 ;
  LAYER M2 ;
        RECT 0.64 29.216 3.52 29.248 ;
  LAYER M1 ;
        RECT 0.624 29.196 0.656 29.268 ;
  LAYER M2 ;
        RECT 0.604 29.216 0.676 29.248 ;
  LAYER M1 ;
        RECT 6.384 29.196 6.416 29.268 ;
  LAYER M2 ;
        RECT 6.364 29.216 6.436 29.248 ;
  LAYER M2 ;
        RECT 3.52 29.216 6.4 29.248 ;
  LAYER M1 ;
        RECT 3.504 29.196 3.536 29.268 ;
  LAYER M2 ;
        RECT 3.484 29.216 3.556 29.248 ;
  LAYER M1 ;
        RECT 9.264 29.196 9.296 29.268 ;
  LAYER M2 ;
        RECT 9.244 29.216 9.316 29.248 ;
  LAYER M2 ;
        RECT 6.4 29.216 9.28 29.248 ;
  LAYER M1 ;
        RECT 6.384 29.196 6.416 29.268 ;
  LAYER M2 ;
        RECT 6.364 29.216 6.436 29.248 ;
  LAYER M1 ;
        RECT 9.264 20.376 9.296 20.448 ;
  LAYER M2 ;
        RECT 9.244 20.396 9.316 20.428 ;
  LAYER M2 ;
        RECT 9.28 20.396 12.16 20.428 ;
  LAYER M1 ;
        RECT 12.144 20.376 12.176 20.448 ;
  LAYER M2 ;
        RECT 12.124 20.396 12.196 20.428 ;
  LAYER M1 ;
        RECT 6.384 20.376 6.416 20.448 ;
  LAYER M2 ;
        RECT 6.364 20.396 6.436 20.428 ;
  LAYER M2 ;
        RECT 6.4 20.396 9.28 20.428 ;
  LAYER M1 ;
        RECT 9.264 20.376 9.296 20.448 ;
  LAYER M2 ;
        RECT 9.244 20.396 9.316 20.428 ;
  LAYER M1 ;
        RECT 0.64 17.976 3.04 20.412 ;
  LAYER M2 ;
        RECT 0.64 17.976 3.04 20.412 ;
  LAYER M3 ;
        RECT 0.64 17.976 3.04 20.412 ;
  LAYER M1 ;
        RECT 0.64 20.916 3.04 23.352 ;
  LAYER M2 ;
        RECT 0.64 20.916 3.04 23.352 ;
  LAYER M3 ;
        RECT 0.64 20.916 3.04 23.352 ;
  LAYER M1 ;
        RECT 0.64 23.856 3.04 26.292 ;
  LAYER M2 ;
        RECT 0.64 23.856 3.04 26.292 ;
  LAYER M3 ;
        RECT 0.64 23.856 3.04 26.292 ;
  LAYER M1 ;
        RECT 0.64 26.796 3.04 29.232 ;
  LAYER M2 ;
        RECT 0.64 26.796 3.04 29.232 ;
  LAYER M3 ;
        RECT 0.64 26.796 3.04 29.232 ;
  LAYER M1 ;
        RECT 3.52 17.976 5.92 20.412 ;
  LAYER M2 ;
        RECT 3.52 17.976 5.92 20.412 ;
  LAYER M3 ;
        RECT 3.52 17.976 5.92 20.412 ;
  LAYER M1 ;
        RECT 3.52 20.916 5.92 23.352 ;
  LAYER M2 ;
        RECT 3.52 20.916 5.92 23.352 ;
  LAYER M3 ;
        RECT 3.52 20.916 5.92 23.352 ;
  LAYER M1 ;
        RECT 3.52 23.856 5.92 26.292 ;
  LAYER M2 ;
        RECT 3.52 23.856 5.92 26.292 ;
  LAYER M3 ;
        RECT 3.52 23.856 5.92 26.292 ;
  LAYER M1 ;
        RECT 3.52 26.796 5.92 29.232 ;
  LAYER M2 ;
        RECT 3.52 26.796 5.92 29.232 ;
  LAYER M3 ;
        RECT 3.52 26.796 5.92 29.232 ;
  LAYER M1 ;
        RECT 6.4 17.976 8.8 20.412 ;
  LAYER M2 ;
        RECT 6.4 17.976 8.8 20.412 ;
  LAYER M3 ;
        RECT 6.4 17.976 8.8 20.412 ;
  LAYER M1 ;
        RECT 6.4 20.916 8.8 23.352 ;
  LAYER M2 ;
        RECT 6.4 20.916 8.8 23.352 ;
  LAYER M3 ;
        RECT 6.4 20.916 8.8 23.352 ;
  LAYER M1 ;
        RECT 6.4 23.856 8.8 26.292 ;
  LAYER M2 ;
        RECT 6.4 23.856 8.8 26.292 ;
  LAYER M3 ;
        RECT 6.4 23.856 8.8 26.292 ;
  LAYER M1 ;
        RECT 6.4 26.796 8.8 29.232 ;
  LAYER M2 ;
        RECT 6.4 26.796 8.8 29.232 ;
  LAYER M3 ;
        RECT 6.4 26.796 8.8 29.232 ;
  LAYER M1 ;
        RECT 9.28 17.976 11.68 20.412 ;
  LAYER M2 ;
        RECT 9.28 17.976 11.68 20.412 ;
  LAYER M3 ;
        RECT 9.28 17.976 11.68 20.412 ;
  LAYER M1 ;
        RECT 9.28 20.916 11.68 23.352 ;
  LAYER M2 ;
        RECT 9.28 20.916 11.68 23.352 ;
  LAYER M3 ;
        RECT 9.28 20.916 11.68 23.352 ;
  LAYER M1 ;
        RECT 9.28 23.856 11.68 26.292 ;
  LAYER M2 ;
        RECT 9.28 23.856 11.68 26.292 ;
  LAYER M3 ;
        RECT 9.28 23.856 11.68 26.292 ;
  LAYER M1 ;
        RECT 9.28 26.796 11.68 29.232 ;
  LAYER M2 ;
        RECT 9.28 26.796 11.68 29.232 ;
  LAYER M3 ;
        RECT 9.28 26.796 11.68 29.232 ;
  LAYER M1 ;
        RECT 12.16 17.976 14.56 20.412 ;
  LAYER M2 ;
        RECT 12.16 17.976 14.56 20.412 ;
  LAYER M3 ;
        RECT 12.16 17.976 14.56 20.412 ;
  LAYER M1 ;
        RECT 12.16 20.916 14.56 23.352 ;
  LAYER M2 ;
        RECT 12.16 20.916 14.56 23.352 ;
  LAYER M3 ;
        RECT 12.16 20.916 14.56 23.352 ;
  LAYER M1 ;
        RECT 12.16 23.856 14.56 26.292 ;
  LAYER M2 ;
        RECT 12.16 23.856 14.56 26.292 ;
  LAYER M3 ;
        RECT 12.16 23.856 14.56 26.292 ;
  LAYER M1 ;
        RECT 12.16 26.796 14.56 29.232 ;
  LAYER M2 ;
        RECT 12.16 26.796 14.56 29.232 ;
  LAYER M3 ;
        RECT 12.16 26.796 14.56 29.232 ;
  LAYER M1 ;
        RECT 5.104 0.3 5.136 0.96 ;
  LAYER M1 ;
        RECT 5.024 0.3 5.056 0.96 ;
  LAYER M1 ;
        RECT 5.184 0.3 5.216 0.96 ;
  LAYER M2 ;
        RECT 4.924 0.908 5.236 0.94 ;
  LAYER M2 ;
        RECT 4.924 0.656 5.236 0.688 ;
  LAYER M2 ;
        RECT 5.004 0.824 5.316 0.856 ;
  LAYER M2 ;
        RECT 5.004 0.572 5.316 0.604 ;
  LAYER M2 ;
        RECT 5.004 0.74 5.396 0.772 ;
  LAYER M2 ;
        RECT 5.004 0.488 5.396 0.52 ;
  LAYER M1 ;
        RECT 15.184 17.352 15.216 18.012 ;
  LAYER M1 ;
        RECT 15.104 17.352 15.136 18.012 ;
  LAYER M1 ;
        RECT 15.264 17.352 15.296 18.012 ;
  LAYER M2 ;
        RECT 15.004 17.96 15.316 17.992 ;
  LAYER M2 ;
        RECT 15.004 17.708 15.316 17.74 ;
  LAYER M2 ;
        RECT 15.084 17.876 15.396 17.908 ;
  LAYER M2 ;
        RECT 15.084 17.624 15.396 17.656 ;
  LAYER M2 ;
        RECT 15.084 17.792 15.476 17.824 ;
  LAYER M2 ;
        RECT 15.084 17.54 15.476 17.572 ;
  LAYER M1 ;
        RECT 6.464 0.3 6.496 0.96 ;
  LAYER M1 ;
        RECT 6.544 0.3 6.576 0.96 ;
  LAYER M1 ;
        RECT 6.384 0.3 6.416 0.96 ;
  LAYER M1 ;
        RECT 5.824 0.3 5.856 0.96 ;
  LAYER M1 ;
        RECT 5.904 0.3 5.936 0.96 ;
  LAYER M1 ;
        RECT 5.744 0.3 5.776 0.96 ;
  LAYER M1 ;
        RECT 7.184 0.3 7.216 0.96 ;
  LAYER M1 ;
        RECT 7.104 0.3 7.136 0.96 ;
  LAYER M1 ;
        RECT 7.264 0.3 7.296 0.96 ;
  LAYER M1 ;
        RECT 7.824 0.3 7.856 0.96 ;
  LAYER M1 ;
        RECT 7.744 0.3 7.776 0.96 ;
  LAYER M1 ;
        RECT 7.904 0.3 7.936 0.96 ;
  LAYER M1 ;
        RECT 6.304 10.296 6.336 10.368 ;
  LAYER M2 ;
        RECT 6.284 10.316 6.356 10.348 ;
  LAYER M2 ;
        RECT 6.32 10.316 9.04 10.348 ;
  LAYER M1 ;
        RECT 9.024 10.296 9.056 10.368 ;
  LAYER M2 ;
        RECT 9.004 10.316 9.076 10.348 ;
  LAYER M1 ;
        RECT 9.184 7.356 9.216 7.428 ;
  LAYER M2 ;
        RECT 9.164 7.376 9.236 7.408 ;
  LAYER M1 ;
        RECT 9.184 7.392 9.216 7.56 ;
  LAYER M1 ;
        RECT 9.184 7.524 9.216 7.596 ;
  LAYER M2 ;
        RECT 9.164 7.544 9.236 7.576 ;
  LAYER M2 ;
        RECT 9.04 7.544 9.2 7.576 ;
  LAYER M1 ;
        RECT 9.024 7.524 9.056 7.596 ;
  LAYER M2 ;
        RECT 9.004 7.544 9.076 7.576 ;
  LAYER M1 ;
        RECT 9.024 16.68 9.056 16.752 ;
  LAYER M2 ;
        RECT 9.004 16.7 9.076 16.732 ;
  LAYER M1 ;
        RECT 9.024 16.548 9.056 16.716 ;
  LAYER M1 ;
        RECT 9.024 7.56 9.056 16.548 ;
  LAYER M1 ;
        RECT 3.424 13.236 3.456 13.308 ;
  LAYER M2 ;
        RECT 3.404 13.256 3.476 13.288 ;
  LAYER M2 ;
        RECT 3.44 13.256 6.16 13.288 ;
  LAYER M1 ;
        RECT 6.144 13.236 6.176 13.308 ;
  LAYER M2 ;
        RECT 6.124 13.256 6.196 13.288 ;
  LAYER M1 ;
        RECT 6.144 16.68 6.176 16.752 ;
  LAYER M2 ;
        RECT 6.124 16.7 6.196 16.732 ;
  LAYER M1 ;
        RECT 6.144 16.548 6.176 16.716 ;
  LAYER M1 ;
        RECT 6.144 13.272 6.176 16.548 ;
  LAYER M2 ;
        RECT 6.16 16.7 9.04 16.732 ;
  LAYER M1 ;
        RECT 9.184 10.296 9.216 10.368 ;
  LAYER M2 ;
        RECT 9.164 10.316 9.236 10.348 ;
  LAYER M2 ;
        RECT 9.2 10.316 11.92 10.348 ;
  LAYER M1 ;
        RECT 11.904 10.296 11.936 10.368 ;
  LAYER M2 ;
        RECT 11.884 10.316 11.956 10.348 ;
  LAYER M1 ;
        RECT 9.184 13.236 9.216 13.308 ;
  LAYER M2 ;
        RECT 9.164 13.256 9.236 13.288 ;
  LAYER M2 ;
        RECT 9.2 13.256 11.92 13.288 ;
  LAYER M1 ;
        RECT 11.904 13.236 11.936 13.308 ;
  LAYER M2 ;
        RECT 11.884 13.256 11.956 13.288 ;
  LAYER M1 ;
        RECT 11.904 16.848 11.936 16.92 ;
  LAYER M2 ;
        RECT 11.884 16.868 11.956 16.9 ;
  LAYER M1 ;
        RECT 11.904 16.548 11.936 16.884 ;
  LAYER M1 ;
        RECT 11.904 10.332 11.936 16.548 ;
  LAYER M1 ;
        RECT 3.424 10.296 3.456 10.368 ;
  LAYER M2 ;
        RECT 3.404 10.316 3.476 10.348 ;
  LAYER M1 ;
        RECT 3.424 10.332 3.456 10.5 ;
  LAYER M1 ;
        RECT 3.424 10.464 3.456 10.536 ;
  LAYER M2 ;
        RECT 3.404 10.484 3.476 10.516 ;
  LAYER M2 ;
        RECT 3.28 10.484 3.44 10.516 ;
  LAYER M1 ;
        RECT 3.264 10.464 3.296 10.536 ;
  LAYER M2 ;
        RECT 3.244 10.484 3.316 10.516 ;
  LAYER M1 ;
        RECT 3.424 7.356 3.456 7.428 ;
  LAYER M2 ;
        RECT 3.404 7.376 3.476 7.408 ;
  LAYER M1 ;
        RECT 3.424 7.392 3.456 7.56 ;
  LAYER M1 ;
        RECT 3.424 7.524 3.456 7.596 ;
  LAYER M2 ;
        RECT 3.404 7.544 3.476 7.576 ;
  LAYER M2 ;
        RECT 3.28 7.544 3.44 7.576 ;
  LAYER M1 ;
        RECT 3.264 7.524 3.296 7.596 ;
  LAYER M2 ;
        RECT 3.244 7.544 3.316 7.576 ;
  LAYER M1 ;
        RECT 3.264 16.848 3.296 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.868 3.316 16.9 ;
  LAYER M1 ;
        RECT 3.264 16.548 3.296 16.884 ;
  LAYER M1 ;
        RECT 3.264 7.56 3.296 16.548 ;
  LAYER M2 ;
        RECT 3.28 16.868 11.92 16.9 ;
  LAYER M1 ;
        RECT 6.304 13.236 6.336 13.308 ;
  LAYER M2 ;
        RECT 6.284 13.256 6.356 13.288 ;
  LAYER M2 ;
        RECT 6.32 13.256 9.2 13.288 ;
  LAYER M1 ;
        RECT 9.184 13.236 9.216 13.308 ;
  LAYER M2 ;
        RECT 9.164 13.256 9.236 13.288 ;
  LAYER M1 ;
        RECT 6.304 7.356 6.336 7.428 ;
  LAYER M2 ;
        RECT 6.284 7.376 6.356 7.408 ;
  LAYER M2 ;
        RECT 3.44 7.376 6.32 7.408 ;
  LAYER M1 ;
        RECT 3.424 7.356 3.456 7.428 ;
  LAYER M2 ;
        RECT 3.404 7.376 3.476 7.408 ;
  LAYER M1 ;
        RECT 12.064 16.176 12.096 16.248 ;
  LAYER M2 ;
        RECT 12.044 16.196 12.116 16.228 ;
  LAYER M2 ;
        RECT 12.08 16.196 14.8 16.228 ;
  LAYER M1 ;
        RECT 14.784 16.176 14.816 16.248 ;
  LAYER M2 ;
        RECT 14.764 16.196 14.836 16.228 ;
  LAYER M1 ;
        RECT 12.064 13.236 12.096 13.308 ;
  LAYER M2 ;
        RECT 12.044 13.256 12.116 13.288 ;
  LAYER M2 ;
        RECT 12.08 13.256 14.8 13.288 ;
  LAYER M1 ;
        RECT 14.784 13.236 14.816 13.308 ;
  LAYER M2 ;
        RECT 14.764 13.256 14.836 13.288 ;
  LAYER M1 ;
        RECT 12.064 10.296 12.096 10.368 ;
  LAYER M2 ;
        RECT 12.044 10.316 12.116 10.348 ;
  LAYER M2 ;
        RECT 12.08 10.316 14.8 10.348 ;
  LAYER M1 ;
        RECT 14.784 10.296 14.816 10.368 ;
  LAYER M2 ;
        RECT 14.764 10.316 14.836 10.348 ;
  LAYER M1 ;
        RECT 12.064 7.356 12.096 7.428 ;
  LAYER M2 ;
        RECT 12.044 7.376 12.116 7.408 ;
  LAYER M2 ;
        RECT 12.08 7.376 14.8 7.408 ;
  LAYER M1 ;
        RECT 14.784 7.356 14.816 7.428 ;
  LAYER M2 ;
        RECT 14.764 7.376 14.836 7.408 ;
  LAYER M1 ;
        RECT 12.064 4.416 12.096 4.488 ;
  LAYER M2 ;
        RECT 12.044 4.436 12.116 4.468 ;
  LAYER M2 ;
        RECT 12.08 4.436 14.8 4.468 ;
  LAYER M1 ;
        RECT 14.784 4.416 14.816 4.488 ;
  LAYER M2 ;
        RECT 14.764 4.436 14.836 4.468 ;
  LAYER M1 ;
        RECT 14.784 17.016 14.816 17.088 ;
  LAYER M2 ;
        RECT 14.764 17.036 14.836 17.068 ;
  LAYER M1 ;
        RECT 14.784 16.548 14.816 17.052 ;
  LAYER M1 ;
        RECT 14.784 4.452 14.816 16.548 ;
  LAYER M1 ;
        RECT 0.544 16.176 0.576 16.248 ;
  LAYER M2 ;
        RECT 0.524 16.196 0.596 16.228 ;
  LAYER M1 ;
        RECT 0.544 16.212 0.576 16.38 ;
  LAYER M1 ;
        RECT 0.544 16.344 0.576 16.416 ;
  LAYER M2 ;
        RECT 0.524 16.364 0.596 16.396 ;
  LAYER M2 ;
        RECT 0.4 16.364 0.56 16.396 ;
  LAYER M1 ;
        RECT 0.384 16.344 0.416 16.416 ;
  LAYER M2 ;
        RECT 0.364 16.364 0.436 16.396 ;
  LAYER M1 ;
        RECT 0.544 13.236 0.576 13.308 ;
  LAYER M2 ;
        RECT 0.524 13.256 0.596 13.288 ;
  LAYER M1 ;
        RECT 0.544 13.272 0.576 13.44 ;
  LAYER M1 ;
        RECT 0.544 13.404 0.576 13.476 ;
  LAYER M2 ;
        RECT 0.524 13.424 0.596 13.456 ;
  LAYER M2 ;
        RECT 0.4 13.424 0.56 13.456 ;
  LAYER M1 ;
        RECT 0.384 13.404 0.416 13.476 ;
  LAYER M2 ;
        RECT 0.364 13.424 0.436 13.456 ;
  LAYER M1 ;
        RECT 0.544 10.296 0.576 10.368 ;
  LAYER M2 ;
        RECT 0.524 10.316 0.596 10.348 ;
  LAYER M1 ;
        RECT 0.544 10.332 0.576 10.5 ;
  LAYER M1 ;
        RECT 0.544 10.464 0.576 10.536 ;
  LAYER M2 ;
        RECT 0.524 10.484 0.596 10.516 ;
  LAYER M2 ;
        RECT 0.4 10.484 0.56 10.516 ;
  LAYER M1 ;
        RECT 0.384 10.464 0.416 10.536 ;
  LAYER M2 ;
        RECT 0.364 10.484 0.436 10.516 ;
  LAYER M1 ;
        RECT 0.544 7.356 0.576 7.428 ;
  LAYER M2 ;
        RECT 0.524 7.376 0.596 7.408 ;
  LAYER M1 ;
        RECT 0.544 7.392 0.576 7.56 ;
  LAYER M1 ;
        RECT 0.544 7.524 0.576 7.596 ;
  LAYER M2 ;
        RECT 0.524 7.544 0.596 7.576 ;
  LAYER M2 ;
        RECT 0.4 7.544 0.56 7.576 ;
  LAYER M1 ;
        RECT 0.384 7.524 0.416 7.596 ;
  LAYER M2 ;
        RECT 0.364 7.544 0.436 7.576 ;
  LAYER M1 ;
        RECT 0.544 4.416 0.576 4.488 ;
  LAYER M2 ;
        RECT 0.524 4.436 0.596 4.468 ;
  LAYER M1 ;
        RECT 0.544 4.452 0.576 4.62 ;
  LAYER M1 ;
        RECT 0.544 4.584 0.576 4.656 ;
  LAYER M2 ;
        RECT 0.524 4.604 0.596 4.636 ;
  LAYER M2 ;
        RECT 0.4 4.604 0.56 4.636 ;
  LAYER M1 ;
        RECT 0.384 4.584 0.416 4.656 ;
  LAYER M2 ;
        RECT 0.364 4.604 0.436 4.636 ;
  LAYER M1 ;
        RECT 0.384 17.016 0.416 17.088 ;
  LAYER M2 ;
        RECT 0.364 17.036 0.436 17.068 ;
  LAYER M1 ;
        RECT 0.384 16.548 0.416 17.052 ;
  LAYER M1 ;
        RECT 0.384 4.62 0.416 16.548 ;
  LAYER M2 ;
        RECT 0.4 17.036 14.8 17.068 ;
  LAYER M1 ;
        RECT 9.184 16.176 9.216 16.248 ;
  LAYER M2 ;
        RECT 9.164 16.196 9.236 16.228 ;
  LAYER M2 ;
        RECT 9.2 16.196 12.08 16.228 ;
  LAYER M1 ;
        RECT 12.064 16.176 12.096 16.248 ;
  LAYER M2 ;
        RECT 12.044 16.196 12.116 16.228 ;
  LAYER M1 ;
        RECT 9.184 4.416 9.216 4.488 ;
  LAYER M2 ;
        RECT 9.164 4.436 9.236 4.468 ;
  LAYER M2 ;
        RECT 9.2 4.436 12.08 4.468 ;
  LAYER M1 ;
        RECT 12.064 4.416 12.096 4.488 ;
  LAYER M2 ;
        RECT 12.044 4.436 12.116 4.468 ;
  LAYER M1 ;
        RECT 6.304 4.416 6.336 4.488 ;
  LAYER M2 ;
        RECT 6.284 4.436 6.356 4.468 ;
  LAYER M2 ;
        RECT 6.32 4.436 9.2 4.468 ;
  LAYER M1 ;
        RECT 9.184 4.416 9.216 4.488 ;
  LAYER M2 ;
        RECT 9.164 4.436 9.236 4.468 ;
  LAYER M1 ;
        RECT 3.424 4.416 3.456 4.488 ;
  LAYER M2 ;
        RECT 3.404 4.436 3.476 4.468 ;
  LAYER M2 ;
        RECT 3.44 4.436 6.32 4.468 ;
  LAYER M1 ;
        RECT 6.304 4.416 6.336 4.488 ;
  LAYER M2 ;
        RECT 6.284 4.436 6.356 4.468 ;
  LAYER M1 ;
        RECT 3.424 16.176 3.456 16.248 ;
  LAYER M2 ;
        RECT 3.404 16.196 3.476 16.228 ;
  LAYER M2 ;
        RECT 0.56 16.196 3.44 16.228 ;
  LAYER M1 ;
        RECT 0.544 16.176 0.576 16.248 ;
  LAYER M2 ;
        RECT 0.524 16.196 0.596 16.228 ;
  LAYER M1 ;
        RECT 6.304 16.176 6.336 16.248 ;
  LAYER M2 ;
        RECT 6.284 16.196 6.356 16.228 ;
  LAYER M2 ;
        RECT 3.44 16.196 6.32 16.228 ;
  LAYER M1 ;
        RECT 3.424 16.176 3.456 16.248 ;
  LAYER M2 ;
        RECT 3.404 16.196 3.476 16.228 ;
  LAYER M1 ;
        RECT 8.704 7.86 8.736 7.932 ;
  LAYER M2 ;
        RECT 8.684 7.88 8.756 7.912 ;
  LAYER M2 ;
        RECT 8.72 7.88 8.88 7.912 ;
  LAYER M1 ;
        RECT 8.864 7.86 8.896 7.932 ;
  LAYER M2 ;
        RECT 8.844 7.88 8.916 7.912 ;
  LAYER M1 ;
        RECT 11.584 4.92 11.616 4.992 ;
  LAYER M2 ;
        RECT 11.564 4.94 11.636 4.972 ;
  LAYER M1 ;
        RECT 11.584 4.788 11.616 4.956 ;
  LAYER M1 ;
        RECT 11.584 4.752 11.616 4.824 ;
  LAYER M2 ;
        RECT 11.564 4.772 11.636 4.804 ;
  LAYER M2 ;
        RECT 8.88 4.772 11.6 4.804 ;
  LAYER M1 ;
        RECT 8.864 4.752 8.896 4.824 ;
  LAYER M2 ;
        RECT 8.844 4.772 8.916 4.804 ;
  LAYER M1 ;
        RECT 8.864 1.476 8.896 1.548 ;
  LAYER M2 ;
        RECT 8.844 1.496 8.916 1.528 ;
  LAYER M1 ;
        RECT 8.864 1.512 8.896 1.68 ;
  LAYER M1 ;
        RECT 8.864 1.68 8.896 7.896 ;
  LAYER M1 ;
        RECT 5.824 10.8 5.856 10.872 ;
  LAYER M2 ;
        RECT 5.804 10.82 5.876 10.852 ;
  LAYER M2 ;
        RECT 5.84 10.82 6 10.852 ;
  LAYER M1 ;
        RECT 5.984 10.8 6.016 10.872 ;
  LAYER M2 ;
        RECT 5.964 10.82 6.036 10.852 ;
  LAYER M1 ;
        RECT 5.984 1.476 6.016 1.548 ;
  LAYER M2 ;
        RECT 5.964 1.496 6.036 1.528 ;
  LAYER M1 ;
        RECT 5.984 1.512 6.016 1.68 ;
  LAYER M1 ;
        RECT 5.984 1.68 6.016 10.836 ;
  LAYER M2 ;
        RECT 6 1.496 8.88 1.528 ;
  LAYER M1 ;
        RECT 11.584 7.86 11.616 7.932 ;
  LAYER M2 ;
        RECT 11.564 7.88 11.636 7.912 ;
  LAYER M2 ;
        RECT 11.6 7.88 11.76 7.912 ;
  LAYER M1 ;
        RECT 11.744 7.86 11.776 7.932 ;
  LAYER M2 ;
        RECT 11.724 7.88 11.796 7.912 ;
  LAYER M1 ;
        RECT 11.584 10.8 11.616 10.872 ;
  LAYER M2 ;
        RECT 11.564 10.82 11.636 10.852 ;
  LAYER M2 ;
        RECT 11.6 10.82 11.76 10.852 ;
  LAYER M1 ;
        RECT 11.744 10.8 11.776 10.872 ;
  LAYER M2 ;
        RECT 11.724 10.82 11.796 10.852 ;
  LAYER M1 ;
        RECT 11.744 1.308 11.776 1.38 ;
  LAYER M2 ;
        RECT 11.724 1.328 11.796 1.36 ;
  LAYER M1 ;
        RECT 11.744 1.344 11.776 1.68 ;
  LAYER M1 ;
        RECT 11.744 1.68 11.776 10.836 ;
  LAYER M1 ;
        RECT 5.824 7.86 5.856 7.932 ;
  LAYER M2 ;
        RECT 5.804 7.88 5.876 7.912 ;
  LAYER M1 ;
        RECT 5.824 7.728 5.856 7.896 ;
  LAYER M1 ;
        RECT 5.824 7.692 5.856 7.764 ;
  LAYER M2 ;
        RECT 5.804 7.712 5.876 7.744 ;
  LAYER M2 ;
        RECT 3.12 7.712 5.84 7.744 ;
  LAYER M1 ;
        RECT 3.104 7.692 3.136 7.764 ;
  LAYER M2 ;
        RECT 3.084 7.712 3.156 7.744 ;
  LAYER M1 ;
        RECT 5.824 4.92 5.856 4.992 ;
  LAYER M2 ;
        RECT 5.804 4.94 5.876 4.972 ;
  LAYER M1 ;
        RECT 5.824 4.788 5.856 4.956 ;
  LAYER M1 ;
        RECT 5.824 4.752 5.856 4.824 ;
  LAYER M2 ;
        RECT 5.804 4.772 5.876 4.804 ;
  LAYER M2 ;
        RECT 3.12 4.772 5.84 4.804 ;
  LAYER M1 ;
        RECT 3.104 4.752 3.136 4.824 ;
  LAYER M2 ;
        RECT 3.084 4.772 3.156 4.804 ;
  LAYER M1 ;
        RECT 3.104 1.308 3.136 1.38 ;
  LAYER M2 ;
        RECT 3.084 1.328 3.156 1.36 ;
  LAYER M1 ;
        RECT 3.104 1.344 3.136 1.68 ;
  LAYER M1 ;
        RECT 3.104 1.68 3.136 7.728 ;
  LAYER M2 ;
        RECT 3.12 1.328 11.76 1.36 ;
  LAYER M1 ;
        RECT 8.704 10.8 8.736 10.872 ;
  LAYER M2 ;
        RECT 8.684 10.82 8.756 10.852 ;
  LAYER M2 ;
        RECT 8.72 10.82 11.6 10.852 ;
  LAYER M1 ;
        RECT 11.584 10.8 11.616 10.872 ;
  LAYER M2 ;
        RECT 11.564 10.82 11.636 10.852 ;
  LAYER M1 ;
        RECT 8.704 4.92 8.736 4.992 ;
  LAYER M2 ;
        RECT 8.684 4.94 8.756 4.972 ;
  LAYER M2 ;
        RECT 5.84 4.94 8.72 4.972 ;
  LAYER M1 ;
        RECT 5.824 4.92 5.856 4.992 ;
  LAYER M2 ;
        RECT 5.804 4.94 5.876 4.972 ;
  LAYER M1 ;
        RECT 14.464 13.74 14.496 13.812 ;
  LAYER M2 ;
        RECT 14.444 13.76 14.516 13.792 ;
  LAYER M2 ;
        RECT 14.48 13.76 14.64 13.792 ;
  LAYER M1 ;
        RECT 14.624 13.74 14.656 13.812 ;
  LAYER M2 ;
        RECT 14.604 13.76 14.676 13.792 ;
  LAYER M1 ;
        RECT 14.464 10.8 14.496 10.872 ;
  LAYER M2 ;
        RECT 14.444 10.82 14.516 10.852 ;
  LAYER M2 ;
        RECT 14.48 10.82 14.64 10.852 ;
  LAYER M1 ;
        RECT 14.624 10.8 14.656 10.872 ;
  LAYER M2 ;
        RECT 14.604 10.82 14.676 10.852 ;
  LAYER M1 ;
        RECT 14.464 7.86 14.496 7.932 ;
  LAYER M2 ;
        RECT 14.444 7.88 14.516 7.912 ;
  LAYER M2 ;
        RECT 14.48 7.88 14.64 7.912 ;
  LAYER M1 ;
        RECT 14.624 7.86 14.656 7.932 ;
  LAYER M2 ;
        RECT 14.604 7.88 14.676 7.912 ;
  LAYER M1 ;
        RECT 14.464 4.92 14.496 4.992 ;
  LAYER M2 ;
        RECT 14.444 4.94 14.516 4.972 ;
  LAYER M2 ;
        RECT 14.48 4.94 14.64 4.972 ;
  LAYER M1 ;
        RECT 14.624 4.92 14.656 4.992 ;
  LAYER M2 ;
        RECT 14.604 4.94 14.676 4.972 ;
  LAYER M1 ;
        RECT 14.464 1.98 14.496 2.052 ;
  LAYER M2 ;
        RECT 14.444 2 14.516 2.032 ;
  LAYER M2 ;
        RECT 14.48 2 14.64 2.032 ;
  LAYER M1 ;
        RECT 14.624 1.98 14.656 2.052 ;
  LAYER M2 ;
        RECT 14.604 2 14.676 2.032 ;
  LAYER M1 ;
        RECT 14.624 1.14 14.656 1.212 ;
  LAYER M2 ;
        RECT 14.604 1.16 14.676 1.192 ;
  LAYER M1 ;
        RECT 14.624 1.176 14.656 1.68 ;
  LAYER M1 ;
        RECT 14.624 1.68 14.656 13.776 ;
  LAYER M1 ;
        RECT 2.944 13.74 2.976 13.812 ;
  LAYER M2 ;
        RECT 2.924 13.76 2.996 13.792 ;
  LAYER M1 ;
        RECT 2.944 13.608 2.976 13.776 ;
  LAYER M1 ;
        RECT 2.944 13.572 2.976 13.644 ;
  LAYER M2 ;
        RECT 2.924 13.592 2.996 13.624 ;
  LAYER M2 ;
        RECT 0.24 13.592 2.96 13.624 ;
  LAYER M1 ;
        RECT 0.224 13.572 0.256 13.644 ;
  LAYER M2 ;
        RECT 0.204 13.592 0.276 13.624 ;
  LAYER M1 ;
        RECT 2.944 10.8 2.976 10.872 ;
  LAYER M2 ;
        RECT 2.924 10.82 2.996 10.852 ;
  LAYER M1 ;
        RECT 2.944 10.668 2.976 10.836 ;
  LAYER M1 ;
        RECT 2.944 10.632 2.976 10.704 ;
  LAYER M2 ;
        RECT 2.924 10.652 2.996 10.684 ;
  LAYER M2 ;
        RECT 0.24 10.652 2.96 10.684 ;
  LAYER M1 ;
        RECT 0.224 10.632 0.256 10.704 ;
  LAYER M2 ;
        RECT 0.204 10.652 0.276 10.684 ;
  LAYER M1 ;
        RECT 2.944 7.86 2.976 7.932 ;
  LAYER M2 ;
        RECT 2.924 7.88 2.996 7.912 ;
  LAYER M1 ;
        RECT 2.944 7.728 2.976 7.896 ;
  LAYER M1 ;
        RECT 2.944 7.692 2.976 7.764 ;
  LAYER M2 ;
        RECT 2.924 7.712 2.996 7.744 ;
  LAYER M2 ;
        RECT 0.24 7.712 2.96 7.744 ;
  LAYER M1 ;
        RECT 0.224 7.692 0.256 7.764 ;
  LAYER M2 ;
        RECT 0.204 7.712 0.276 7.744 ;
  LAYER M1 ;
        RECT 2.944 4.92 2.976 4.992 ;
  LAYER M2 ;
        RECT 2.924 4.94 2.996 4.972 ;
  LAYER M1 ;
        RECT 2.944 4.788 2.976 4.956 ;
  LAYER M1 ;
        RECT 2.944 4.752 2.976 4.824 ;
  LAYER M2 ;
        RECT 2.924 4.772 2.996 4.804 ;
  LAYER M2 ;
        RECT 0.24 4.772 2.96 4.804 ;
  LAYER M1 ;
        RECT 0.224 4.752 0.256 4.824 ;
  LAYER M2 ;
        RECT 0.204 4.772 0.276 4.804 ;
  LAYER M1 ;
        RECT 2.944 1.98 2.976 2.052 ;
  LAYER M2 ;
        RECT 2.924 2 2.996 2.032 ;
  LAYER M1 ;
        RECT 2.944 1.848 2.976 2.016 ;
  LAYER M1 ;
        RECT 2.944 1.812 2.976 1.884 ;
  LAYER M2 ;
        RECT 2.924 1.832 2.996 1.864 ;
  LAYER M2 ;
        RECT 0.24 1.832 2.96 1.864 ;
  LAYER M1 ;
        RECT 0.224 1.812 0.256 1.884 ;
  LAYER M2 ;
        RECT 0.204 1.832 0.276 1.864 ;
  LAYER M1 ;
        RECT 0.224 1.14 0.256 1.212 ;
  LAYER M2 ;
        RECT 0.204 1.16 0.276 1.192 ;
  LAYER M1 ;
        RECT 0.224 1.176 0.256 1.68 ;
  LAYER M1 ;
        RECT 0.224 1.68 0.256 13.608 ;
  LAYER M2 ;
        RECT 0.24 1.16 14.64 1.192 ;
  LAYER M1 ;
        RECT 11.584 13.74 11.616 13.812 ;
  LAYER M2 ;
        RECT 11.564 13.76 11.636 13.792 ;
  LAYER M2 ;
        RECT 11.6 13.76 14.48 13.792 ;
  LAYER M1 ;
        RECT 14.464 13.74 14.496 13.812 ;
  LAYER M2 ;
        RECT 14.444 13.76 14.516 13.792 ;
  LAYER M1 ;
        RECT 11.584 1.98 11.616 2.052 ;
  LAYER M2 ;
        RECT 11.564 2 11.636 2.032 ;
  LAYER M2 ;
        RECT 11.6 2 14.48 2.032 ;
  LAYER M1 ;
        RECT 14.464 1.98 14.496 2.052 ;
  LAYER M2 ;
        RECT 14.444 2 14.516 2.032 ;
  LAYER M1 ;
        RECT 8.704 1.98 8.736 2.052 ;
  LAYER M2 ;
        RECT 8.684 2 8.756 2.032 ;
  LAYER M2 ;
        RECT 8.72 2 11.6 2.032 ;
  LAYER M1 ;
        RECT 11.584 1.98 11.616 2.052 ;
  LAYER M2 ;
        RECT 11.564 2 11.636 2.032 ;
  LAYER M1 ;
        RECT 5.824 1.98 5.856 2.052 ;
  LAYER M2 ;
        RECT 5.804 2 5.876 2.032 ;
  LAYER M2 ;
        RECT 5.84 2 8.72 2.032 ;
  LAYER M1 ;
        RECT 8.704 1.98 8.736 2.052 ;
  LAYER M2 ;
        RECT 8.684 2 8.756 2.032 ;
  LAYER M1 ;
        RECT 5.824 13.74 5.856 13.812 ;
  LAYER M2 ;
        RECT 5.804 13.76 5.876 13.792 ;
  LAYER M2 ;
        RECT 2.96 13.76 5.84 13.792 ;
  LAYER M1 ;
        RECT 2.944 13.74 2.976 13.812 ;
  LAYER M2 ;
        RECT 2.924 13.76 2.996 13.792 ;
  LAYER M1 ;
        RECT 8.704 13.74 8.736 13.812 ;
  LAYER M2 ;
        RECT 8.684 13.76 8.756 13.792 ;
  LAYER M2 ;
        RECT 5.84 13.76 8.72 13.792 ;
  LAYER M1 ;
        RECT 5.824 13.74 5.856 13.812 ;
  LAYER M2 ;
        RECT 5.804 13.76 5.876 13.792 ;
  LAYER M1 ;
        RECT 12.08 13.776 14.48 16.212 ;
  LAYER M2 ;
        RECT 12.08 13.776 14.48 16.212 ;
  LAYER M3 ;
        RECT 12.08 13.776 14.48 16.212 ;
  LAYER M1 ;
        RECT 12.08 10.836 14.48 13.272 ;
  LAYER M2 ;
        RECT 12.08 10.836 14.48 13.272 ;
  LAYER M3 ;
        RECT 12.08 10.836 14.48 13.272 ;
  LAYER M1 ;
        RECT 12.08 7.896 14.48 10.332 ;
  LAYER M2 ;
        RECT 12.08 7.896 14.48 10.332 ;
  LAYER M3 ;
        RECT 12.08 7.896 14.48 10.332 ;
  LAYER M1 ;
        RECT 12.08 4.956 14.48 7.392 ;
  LAYER M2 ;
        RECT 12.08 4.956 14.48 7.392 ;
  LAYER M3 ;
        RECT 12.08 4.956 14.48 7.392 ;
  LAYER M1 ;
        RECT 12.08 2.016 14.48 4.452 ;
  LAYER M2 ;
        RECT 12.08 2.016 14.48 4.452 ;
  LAYER M3 ;
        RECT 12.08 2.016 14.48 4.452 ;
  LAYER M1 ;
        RECT 9.2 13.776 11.6 16.212 ;
  LAYER M2 ;
        RECT 9.2 13.776 11.6 16.212 ;
  LAYER M3 ;
        RECT 9.2 13.776 11.6 16.212 ;
  LAYER M1 ;
        RECT 9.2 10.836 11.6 13.272 ;
  LAYER M2 ;
        RECT 9.2 10.836 11.6 13.272 ;
  LAYER M3 ;
        RECT 9.2 10.836 11.6 13.272 ;
  LAYER M1 ;
        RECT 9.2 7.896 11.6 10.332 ;
  LAYER M2 ;
        RECT 9.2 7.896 11.6 10.332 ;
  LAYER M3 ;
        RECT 9.2 7.896 11.6 10.332 ;
  LAYER M1 ;
        RECT 9.2 4.956 11.6 7.392 ;
  LAYER M2 ;
        RECT 9.2 4.956 11.6 7.392 ;
  LAYER M3 ;
        RECT 9.2 4.956 11.6 7.392 ;
  LAYER M1 ;
        RECT 9.2 2.016 11.6 4.452 ;
  LAYER M2 ;
        RECT 9.2 2.016 11.6 4.452 ;
  LAYER M3 ;
        RECT 9.2 2.016 11.6 4.452 ;
  LAYER M1 ;
        RECT 6.32 13.776 8.72 16.212 ;
  LAYER M2 ;
        RECT 6.32 13.776 8.72 16.212 ;
  LAYER M3 ;
        RECT 6.32 13.776 8.72 16.212 ;
  LAYER M1 ;
        RECT 6.32 10.836 8.72 13.272 ;
  LAYER M2 ;
        RECT 6.32 10.836 8.72 13.272 ;
  LAYER M3 ;
        RECT 6.32 10.836 8.72 13.272 ;
  LAYER M1 ;
        RECT 6.32 7.896 8.72 10.332 ;
  LAYER M2 ;
        RECT 6.32 7.896 8.72 10.332 ;
  LAYER M3 ;
        RECT 6.32 7.896 8.72 10.332 ;
  LAYER M1 ;
        RECT 6.32 4.956 8.72 7.392 ;
  LAYER M2 ;
        RECT 6.32 4.956 8.72 7.392 ;
  LAYER M3 ;
        RECT 6.32 4.956 8.72 7.392 ;
  LAYER M1 ;
        RECT 6.32 2.016 8.72 4.452 ;
  LAYER M2 ;
        RECT 6.32 2.016 8.72 4.452 ;
  LAYER M3 ;
        RECT 6.32 2.016 8.72 4.452 ;
  LAYER M1 ;
        RECT 3.44 13.776 5.84 16.212 ;
  LAYER M2 ;
        RECT 3.44 13.776 5.84 16.212 ;
  LAYER M3 ;
        RECT 3.44 13.776 5.84 16.212 ;
  LAYER M1 ;
        RECT 3.44 10.836 5.84 13.272 ;
  LAYER M2 ;
        RECT 3.44 10.836 5.84 13.272 ;
  LAYER M3 ;
        RECT 3.44 10.836 5.84 13.272 ;
  LAYER M1 ;
        RECT 3.44 7.896 5.84 10.332 ;
  LAYER M2 ;
        RECT 3.44 7.896 5.84 10.332 ;
  LAYER M3 ;
        RECT 3.44 7.896 5.84 10.332 ;
  LAYER M1 ;
        RECT 3.44 4.956 5.84 7.392 ;
  LAYER M2 ;
        RECT 3.44 4.956 5.84 7.392 ;
  LAYER M3 ;
        RECT 3.44 4.956 5.84 7.392 ;
  LAYER M1 ;
        RECT 3.44 2.016 5.84 4.452 ;
  LAYER M2 ;
        RECT 3.44 2.016 5.84 4.452 ;
  LAYER M3 ;
        RECT 3.44 2.016 5.84 4.452 ;
  LAYER M1 ;
        RECT 0.56 13.776 2.96 16.212 ;
  LAYER M2 ;
        RECT 0.56 13.776 2.96 16.212 ;
  LAYER M3 ;
        RECT 0.56 13.776 2.96 16.212 ;
  LAYER M1 ;
        RECT 0.56 10.836 2.96 13.272 ;
  LAYER M2 ;
        RECT 0.56 10.836 2.96 13.272 ;
  LAYER M3 ;
        RECT 0.56 10.836 2.96 13.272 ;
  LAYER M1 ;
        RECT 0.56 7.896 2.96 10.332 ;
  LAYER M2 ;
        RECT 0.56 7.896 2.96 10.332 ;
  LAYER M3 ;
        RECT 0.56 7.896 2.96 10.332 ;
  LAYER M1 ;
        RECT 0.56 4.956 2.96 7.392 ;
  LAYER M2 ;
        RECT 0.56 4.956 2.96 7.392 ;
  LAYER M3 ;
        RECT 0.56 4.956 2.96 7.392 ;
  LAYER M1 ;
        RECT 0.56 2.016 2.96 4.452 ;
  LAYER M2 ;
        RECT 0.56 2.016 2.96 4.452 ;
  LAYER M3 ;
        RECT 0.56 2.016 2.96 4.452 ;
  LAYER M1 ;
        RECT 39.824 29.7 39.856 29.772 ;
  LAYER M2 ;
        RECT 39.804 29.72 39.876 29.752 ;
  LAYER M1 ;
        RECT 36.944 29.7 36.976 29.772 ;
  LAYER M2 ;
        RECT 36.924 29.72 36.996 29.752 ;
  LAYER M2 ;
        RECT 36.96 29.72 39.84 29.752 ;
  LAYER M2 ;
        RECT 39.484 0.908 40.196 0.94 ;
  LAYER M1 ;
        RECT 37.024 16.68 37.056 16.752 ;
  LAYER M2 ;
        RECT 37.004 16.7 37.076 16.732 ;
  LAYER M1 ;
        RECT 39.904 16.68 39.936 16.752 ;
  LAYER M2 ;
        RECT 39.884 16.7 39.956 16.732 ;
  LAYER M2 ;
        RECT 37.04 16.7 39.92 16.732 ;
  LAYER M2 ;
        RECT 37.58 29.72 37.78 29.752 ;
  LAYER M3 ;
        RECT 37.66 29.484 37.7 29.736 ;
  LAYER M4 ;
        RECT 37.61 29.464 37.75 29.504 ;
  LAYER M5 ;
        RECT 37.648 16.968 37.712 29.484 ;
  LAYER M4 ;
        RECT 37.61 16.948 37.75 16.988 ;
  LAYER M3 ;
        RECT 37.66 16.716 37.7 16.968 ;
  LAYER M2 ;
        RECT 37.58 16.7 37.78 16.732 ;
  LAYER M2 ;
        RECT 39.74 16.7 39.94 16.732 ;
  LAYER M3 ;
        RECT 39.82 1.596 39.86 16.716 ;
  LAYER M4 ;
        RECT 39.77 1.576 39.91 1.616 ;
  LAYER M5 ;
        RECT 39.808 1.428 39.872 1.596 ;
  LAYER M4 ;
        RECT 39.77 1.408 39.91 1.448 ;
  LAYER M3 ;
        RECT 39.82 0.924 39.86 1.428 ;
  LAYER M2 ;
        RECT 39.74 0.908 39.94 0.94 ;
  LAYER M1 ;
        RECT 39.984 17.436 40.016 17.508 ;
  LAYER M2 ;
        RECT 39.964 17.456 40.036 17.488 ;
  LAYER M1 ;
        RECT 37.104 17.436 37.136 17.508 ;
  LAYER M2 ;
        RECT 37.084 17.456 37.156 17.488 ;
  LAYER M2 ;
        RECT 37.12 17.456 40 17.488 ;
  LAYER M3 ;
        RECT 41.02 0.552 41.06 0.876 ;
  LAYER M3 ;
        RECT 40.78 0.552 40.82 0.876 ;
  LAYER M3 ;
        RECT 30.94 17.604 30.98 17.928 ;
  LAYER M3 ;
        RECT 30.7 17.604 30.74 17.928 ;
  LAYER M2 ;
        RECT 31.12 17.456 37.12 17.488 ;
  LAYER M3 ;
        RECT 31.1 17.367 31.14 17.577 ;
  LAYER M4 ;
        RECT 30.96 17.452 31.12 17.492 ;
  LAYER M3 ;
        RECT 30.94 17.472 30.98 17.724 ;
  LAYER M2 ;
        RECT 39.9 17.456 40.1 17.488 ;
  LAYER M3 ;
        RECT 39.98 0.84 40.02 17.472 ;
  LAYER M4 ;
        RECT 40 0.82 40.8 0.86 ;
  LAYER M3 ;
        RECT 40.78 0.735 40.82 0.945 ;
  LAYER M2 ;
        RECT 38.284 0.908 38.996 0.94 ;
  LAYER M1 ;
        RECT 37.184 1.476 37.216 1.548 ;
  LAYER M2 ;
        RECT 37.164 1.496 37.236 1.528 ;
  LAYER M1 ;
        RECT 40.064 1.476 40.096 1.548 ;
  LAYER M2 ;
        RECT 40.044 1.496 40.116 1.528 ;
  LAYER M2 ;
        RECT 37.2 1.496 40.08 1.528 ;
  LAYER M2 ;
        RECT 38.46 0.908 38.66 0.94 ;
  LAYER M3 ;
        RECT 38.54 0.924 38.58 1.428 ;
  LAYER M4 ;
        RECT 38.4 1.408 38.56 1.448 ;
  LAYER M5 ;
        RECT 38.368 1.42 38.432 1.52 ;
  LAYER M4 ;
        RECT 38.33 1.492 38.47 1.532 ;
  LAYER M3 ;
        RECT 38.38 1.407 38.42 1.617 ;
  LAYER M2 ;
        RECT 38.3 1.496 38.5 1.528 ;
  LAYER M1 ;
        RECT 37.264 20.88 37.296 20.952 ;
  LAYER M2 ;
        RECT 37.244 20.9 37.316 20.932 ;
  LAYER M2 ;
        RECT 37.28 20.9 40 20.932 ;
  LAYER M1 ;
        RECT 39.984 20.88 40.016 20.952 ;
  LAYER M2 ;
        RECT 39.964 20.9 40.036 20.932 ;
  LAYER M1 ;
        RECT 37.264 23.82 37.296 23.892 ;
  LAYER M2 ;
        RECT 37.244 23.84 37.316 23.872 ;
  LAYER M2 ;
        RECT 37.28 23.84 40 23.872 ;
  LAYER M1 ;
        RECT 39.984 23.82 40.016 23.892 ;
  LAYER M2 ;
        RECT 39.964 23.84 40.036 23.872 ;
  LAYER M1 ;
        RECT 40.144 20.88 40.176 20.952 ;
  LAYER M2 ;
        RECT 40.124 20.9 40.196 20.932 ;
  LAYER M1 ;
        RECT 40.144 20.748 40.176 20.916 ;
  LAYER M1 ;
        RECT 40.144 20.712 40.176 20.784 ;
  LAYER M2 ;
        RECT 40.124 20.732 40.196 20.764 ;
  LAYER M2 ;
        RECT 40 20.732 40.16 20.764 ;
  LAYER M1 ;
        RECT 39.984 20.712 40.016 20.784 ;
  LAYER M2 ;
        RECT 39.964 20.732 40.036 20.764 ;
  LAYER M1 ;
        RECT 40.144 23.82 40.176 23.892 ;
  LAYER M2 ;
        RECT 40.124 23.84 40.196 23.872 ;
  LAYER M1 ;
        RECT 40.144 23.688 40.176 23.856 ;
  LAYER M1 ;
        RECT 40.144 23.652 40.176 23.724 ;
  LAYER M2 ;
        RECT 40.124 23.672 40.196 23.704 ;
  LAYER M2 ;
        RECT 40 23.672 40.16 23.704 ;
  LAYER M1 ;
        RECT 39.984 23.652 40.016 23.724 ;
  LAYER M2 ;
        RECT 39.964 23.672 40.036 23.704 ;
  LAYER M1 ;
        RECT 39.984 17.436 40.016 17.508 ;
  LAYER M2 ;
        RECT 39.964 17.456 40.036 17.488 ;
  LAYER M1 ;
        RECT 39.984 17.472 40.016 17.64 ;
  LAYER M1 ;
        RECT 39.984 17.64 40.016 23.856 ;
  LAYER M1 ;
        RECT 34.384 23.82 34.416 23.892 ;
  LAYER M2 ;
        RECT 34.364 23.84 34.436 23.872 ;
  LAYER M2 ;
        RECT 34.4 23.84 37.12 23.872 ;
  LAYER M1 ;
        RECT 37.104 23.82 37.136 23.892 ;
  LAYER M2 ;
        RECT 37.084 23.84 37.156 23.872 ;
  LAYER M1 ;
        RECT 34.384 20.88 34.416 20.952 ;
  LAYER M2 ;
        RECT 34.364 20.9 34.436 20.932 ;
  LAYER M2 ;
        RECT 34.4 20.9 37.12 20.932 ;
  LAYER M1 ;
        RECT 37.104 20.88 37.136 20.952 ;
  LAYER M2 ;
        RECT 37.084 20.9 37.156 20.932 ;
  LAYER M1 ;
        RECT 37.104 17.436 37.136 17.508 ;
  LAYER M2 ;
        RECT 37.084 17.456 37.156 17.488 ;
  LAYER M1 ;
        RECT 37.104 17.472 37.136 17.64 ;
  LAYER M1 ;
        RECT 37.104 17.64 37.136 23.856 ;
  LAYER M2 ;
        RECT 37.12 17.456 40 17.488 ;
  LAYER M1 ;
        RECT 43.024 17.94 43.056 18.012 ;
  LAYER M2 ;
        RECT 43.004 17.96 43.076 17.992 ;
  LAYER M1 ;
        RECT 43.024 17.808 43.056 17.976 ;
  LAYER M1 ;
        RECT 43.024 17.772 43.056 17.844 ;
  LAYER M2 ;
        RECT 43.004 17.792 43.076 17.824 ;
  LAYER M2 ;
        RECT 42.88 17.792 43.04 17.824 ;
  LAYER M1 ;
        RECT 42.864 17.772 42.896 17.844 ;
  LAYER M2 ;
        RECT 42.844 17.792 42.916 17.824 ;
  LAYER M1 ;
        RECT 43.024 20.88 43.056 20.952 ;
  LAYER M2 ;
        RECT 43.004 20.9 43.076 20.932 ;
  LAYER M1 ;
        RECT 43.024 20.748 43.056 20.916 ;
  LAYER M1 ;
        RECT 43.024 20.712 43.056 20.784 ;
  LAYER M2 ;
        RECT 43.004 20.732 43.076 20.764 ;
  LAYER M2 ;
        RECT 42.88 20.732 43.04 20.764 ;
  LAYER M1 ;
        RECT 42.864 20.712 42.896 20.784 ;
  LAYER M2 ;
        RECT 42.844 20.732 42.916 20.764 ;
  LAYER M1 ;
        RECT 43.024 23.82 43.056 23.892 ;
  LAYER M2 ;
        RECT 43.004 23.84 43.076 23.872 ;
  LAYER M1 ;
        RECT 43.024 23.688 43.056 23.856 ;
  LAYER M1 ;
        RECT 43.024 23.652 43.056 23.724 ;
  LAYER M2 ;
        RECT 43.004 23.672 43.076 23.704 ;
  LAYER M2 ;
        RECT 42.88 23.672 43.04 23.704 ;
  LAYER M1 ;
        RECT 42.864 23.652 42.896 23.724 ;
  LAYER M2 ;
        RECT 42.844 23.672 42.916 23.704 ;
  LAYER M1 ;
        RECT 43.024 26.76 43.056 26.832 ;
  LAYER M2 ;
        RECT 43.004 26.78 43.076 26.812 ;
  LAYER M1 ;
        RECT 43.024 26.628 43.056 26.796 ;
  LAYER M1 ;
        RECT 43.024 26.592 43.056 26.664 ;
  LAYER M2 ;
        RECT 43.004 26.612 43.076 26.644 ;
  LAYER M2 ;
        RECT 42.88 26.612 43.04 26.644 ;
  LAYER M1 ;
        RECT 42.864 26.592 42.896 26.664 ;
  LAYER M2 ;
        RECT 42.844 26.612 42.916 26.644 ;
  LAYER M1 ;
        RECT 40.144 17.94 40.176 18.012 ;
  LAYER M2 ;
        RECT 40.124 17.96 40.196 17.992 ;
  LAYER M2 ;
        RECT 40.16 17.96 42.88 17.992 ;
  LAYER M1 ;
        RECT 42.864 17.94 42.896 18.012 ;
  LAYER M2 ;
        RECT 42.844 17.96 42.916 17.992 ;
  LAYER M1 ;
        RECT 40.144 26.76 40.176 26.832 ;
  LAYER M2 ;
        RECT 40.124 26.78 40.196 26.812 ;
  LAYER M2 ;
        RECT 40.16 26.78 42.88 26.812 ;
  LAYER M1 ;
        RECT 42.864 26.76 42.896 26.832 ;
  LAYER M2 ;
        RECT 42.844 26.78 42.916 26.812 ;
  LAYER M1 ;
        RECT 42.864 17.268 42.896 17.34 ;
  LAYER M2 ;
        RECT 42.844 17.288 42.916 17.32 ;
  LAYER M1 ;
        RECT 42.864 17.304 42.896 17.64 ;
  LAYER M1 ;
        RECT 42.864 17.64 42.896 26.796 ;
  LAYER M1 ;
        RECT 34.384 17.94 34.416 18.012 ;
  LAYER M2 ;
        RECT 34.364 17.96 34.436 17.992 ;
  LAYER M1 ;
        RECT 34.384 17.808 34.416 17.976 ;
  LAYER M1 ;
        RECT 34.384 17.772 34.416 17.844 ;
  LAYER M2 ;
        RECT 34.364 17.792 34.436 17.824 ;
  LAYER M2 ;
        RECT 34.24 17.792 34.4 17.824 ;
  LAYER M1 ;
        RECT 34.224 17.772 34.256 17.844 ;
  LAYER M2 ;
        RECT 34.204 17.792 34.276 17.824 ;
  LAYER M1 ;
        RECT 34.384 26.76 34.416 26.832 ;
  LAYER M2 ;
        RECT 34.364 26.78 34.436 26.812 ;
  LAYER M1 ;
        RECT 34.384 26.628 34.416 26.796 ;
  LAYER M1 ;
        RECT 34.384 26.592 34.416 26.664 ;
  LAYER M2 ;
        RECT 34.364 26.612 34.436 26.644 ;
  LAYER M2 ;
        RECT 34.24 26.612 34.4 26.644 ;
  LAYER M1 ;
        RECT 34.224 26.592 34.256 26.664 ;
  LAYER M2 ;
        RECT 34.204 26.612 34.276 26.644 ;
  LAYER M1 ;
        RECT 31.504 17.94 31.536 18.012 ;
  LAYER M2 ;
        RECT 31.484 17.96 31.556 17.992 ;
  LAYER M2 ;
        RECT 31.52 17.96 34.24 17.992 ;
  LAYER M1 ;
        RECT 34.224 17.94 34.256 18.012 ;
  LAYER M2 ;
        RECT 34.204 17.96 34.276 17.992 ;
  LAYER M1 ;
        RECT 31.504 20.88 31.536 20.952 ;
  LAYER M2 ;
        RECT 31.484 20.9 31.556 20.932 ;
  LAYER M2 ;
        RECT 31.52 20.9 34.24 20.932 ;
  LAYER M1 ;
        RECT 34.224 20.88 34.256 20.952 ;
  LAYER M2 ;
        RECT 34.204 20.9 34.276 20.932 ;
  LAYER M1 ;
        RECT 31.504 23.82 31.536 23.892 ;
  LAYER M2 ;
        RECT 31.484 23.84 31.556 23.872 ;
  LAYER M2 ;
        RECT 31.52 23.84 34.24 23.872 ;
  LAYER M1 ;
        RECT 34.224 23.82 34.256 23.892 ;
  LAYER M2 ;
        RECT 34.204 23.84 34.276 23.872 ;
  LAYER M1 ;
        RECT 31.504 26.76 31.536 26.832 ;
  LAYER M2 ;
        RECT 31.484 26.78 31.556 26.812 ;
  LAYER M2 ;
        RECT 31.52 26.78 34.24 26.812 ;
  LAYER M1 ;
        RECT 34.224 26.76 34.256 26.832 ;
  LAYER M2 ;
        RECT 34.204 26.78 34.276 26.812 ;
  LAYER M1 ;
        RECT 34.224 17.268 34.256 17.34 ;
  LAYER M2 ;
        RECT 34.204 17.288 34.276 17.32 ;
  LAYER M1 ;
        RECT 34.224 17.304 34.256 17.64 ;
  LAYER M1 ;
        RECT 34.224 17.64 34.256 26.796 ;
  LAYER M2 ;
        RECT 34.24 17.288 42.88 17.32 ;
  LAYER M1 ;
        RECT 37.264 26.76 37.296 26.832 ;
  LAYER M2 ;
        RECT 37.244 26.78 37.316 26.812 ;
  LAYER M2 ;
        RECT 37.28 26.78 40.16 26.812 ;
  LAYER M1 ;
        RECT 40.144 26.76 40.176 26.832 ;
  LAYER M2 ;
        RECT 40.124 26.78 40.196 26.812 ;
  LAYER M1 ;
        RECT 37.264 17.94 37.296 18.012 ;
  LAYER M2 ;
        RECT 37.244 17.96 37.316 17.992 ;
  LAYER M2 ;
        RECT 34.4 17.96 37.28 17.992 ;
  LAYER M1 ;
        RECT 34.384 17.94 34.416 18.012 ;
  LAYER M2 ;
        RECT 34.364 17.96 34.436 17.992 ;
  LAYER M1 ;
        RECT 39.664 23.316 39.696 23.388 ;
  LAYER M2 ;
        RECT 39.644 23.336 39.716 23.368 ;
  LAYER M2 ;
        RECT 39.68 23.336 39.84 23.368 ;
  LAYER M1 ;
        RECT 39.824 23.316 39.856 23.388 ;
  LAYER M2 ;
        RECT 39.804 23.336 39.876 23.368 ;
  LAYER M1 ;
        RECT 39.664 26.256 39.696 26.328 ;
  LAYER M2 ;
        RECT 39.644 26.276 39.716 26.308 ;
  LAYER M2 ;
        RECT 39.68 26.276 39.84 26.308 ;
  LAYER M1 ;
        RECT 39.824 26.256 39.856 26.328 ;
  LAYER M2 ;
        RECT 39.804 26.276 39.876 26.308 ;
  LAYER M1 ;
        RECT 42.544 23.316 42.576 23.388 ;
  LAYER M2 ;
        RECT 42.524 23.336 42.596 23.368 ;
  LAYER M1 ;
        RECT 42.544 23.352 42.576 23.52 ;
  LAYER M1 ;
        RECT 42.544 23.484 42.576 23.556 ;
  LAYER M2 ;
        RECT 42.524 23.504 42.596 23.536 ;
  LAYER M2 ;
        RECT 39.84 23.504 42.56 23.536 ;
  LAYER M1 ;
        RECT 39.824 23.484 39.856 23.556 ;
  LAYER M2 ;
        RECT 39.804 23.504 39.876 23.536 ;
  LAYER M1 ;
        RECT 42.544 26.256 42.576 26.328 ;
  LAYER M2 ;
        RECT 42.524 26.276 42.596 26.308 ;
  LAYER M1 ;
        RECT 42.544 26.292 42.576 26.46 ;
  LAYER M1 ;
        RECT 42.544 26.424 42.576 26.496 ;
  LAYER M2 ;
        RECT 42.524 26.444 42.596 26.476 ;
  LAYER M2 ;
        RECT 39.84 26.444 42.56 26.476 ;
  LAYER M1 ;
        RECT 39.824 26.424 39.856 26.496 ;
  LAYER M2 ;
        RECT 39.804 26.444 39.876 26.476 ;
  LAYER M1 ;
        RECT 39.824 29.7 39.856 29.772 ;
  LAYER M2 ;
        RECT 39.804 29.72 39.876 29.752 ;
  LAYER M1 ;
        RECT 39.824 29.568 39.856 29.736 ;
  LAYER M1 ;
        RECT 39.824 23.352 39.856 29.568 ;
  LAYER M1 ;
        RECT 36.784 26.256 36.816 26.328 ;
  LAYER M2 ;
        RECT 36.764 26.276 36.836 26.308 ;
  LAYER M2 ;
        RECT 36.8 26.276 36.96 26.308 ;
  LAYER M1 ;
        RECT 36.944 26.256 36.976 26.328 ;
  LAYER M2 ;
        RECT 36.924 26.276 36.996 26.308 ;
  LAYER M1 ;
        RECT 36.784 23.316 36.816 23.388 ;
  LAYER M2 ;
        RECT 36.764 23.336 36.836 23.368 ;
  LAYER M2 ;
        RECT 36.8 23.336 36.96 23.368 ;
  LAYER M1 ;
        RECT 36.944 23.316 36.976 23.388 ;
  LAYER M2 ;
        RECT 36.924 23.336 36.996 23.368 ;
  LAYER M1 ;
        RECT 36.944 29.7 36.976 29.772 ;
  LAYER M2 ;
        RECT 36.924 29.72 36.996 29.752 ;
  LAYER M1 ;
        RECT 36.944 29.568 36.976 29.736 ;
  LAYER M1 ;
        RECT 36.944 23.352 36.976 29.568 ;
  LAYER M2 ;
        RECT 36.96 29.72 39.84 29.752 ;
  LAYER M1 ;
        RECT 45.424 20.376 45.456 20.448 ;
  LAYER M2 ;
        RECT 45.404 20.396 45.476 20.428 ;
  LAYER M2 ;
        RECT 45.44 20.396 45.76 20.428 ;
  LAYER M1 ;
        RECT 45.744 20.376 45.776 20.448 ;
  LAYER M2 ;
        RECT 45.724 20.396 45.796 20.428 ;
  LAYER M1 ;
        RECT 45.424 23.316 45.456 23.388 ;
  LAYER M2 ;
        RECT 45.404 23.336 45.476 23.368 ;
  LAYER M2 ;
        RECT 45.44 23.336 45.76 23.368 ;
  LAYER M1 ;
        RECT 45.744 23.316 45.776 23.388 ;
  LAYER M2 ;
        RECT 45.724 23.336 45.796 23.368 ;
  LAYER M1 ;
        RECT 45.424 26.256 45.456 26.328 ;
  LAYER M2 ;
        RECT 45.404 26.276 45.476 26.308 ;
  LAYER M2 ;
        RECT 45.44 26.276 45.76 26.308 ;
  LAYER M1 ;
        RECT 45.744 26.256 45.776 26.328 ;
  LAYER M2 ;
        RECT 45.724 26.276 45.796 26.308 ;
  LAYER M1 ;
        RECT 45.424 29.196 45.456 29.268 ;
  LAYER M2 ;
        RECT 45.404 29.216 45.476 29.248 ;
  LAYER M2 ;
        RECT 45.44 29.216 45.76 29.248 ;
  LAYER M1 ;
        RECT 45.744 29.196 45.776 29.268 ;
  LAYER M2 ;
        RECT 45.724 29.216 45.796 29.248 ;
  LAYER M1 ;
        RECT 45.744 29.868 45.776 29.94 ;
  LAYER M2 ;
        RECT 45.724 29.888 45.796 29.92 ;
  LAYER M1 ;
        RECT 45.744 29.568 45.776 29.904 ;
  LAYER M1 ;
        RECT 45.744 20.412 45.776 29.568 ;
  LAYER M1 ;
        RECT 33.904 20.376 33.936 20.448 ;
  LAYER M2 ;
        RECT 33.884 20.396 33.956 20.428 ;
  LAYER M1 ;
        RECT 33.904 20.412 33.936 20.58 ;
  LAYER M1 ;
        RECT 33.904 20.544 33.936 20.616 ;
  LAYER M2 ;
        RECT 33.884 20.564 33.956 20.596 ;
  LAYER M2 ;
        RECT 31.36 20.564 33.92 20.596 ;
  LAYER M1 ;
        RECT 31.344 20.544 31.376 20.616 ;
  LAYER M2 ;
        RECT 31.324 20.564 31.396 20.596 ;
  LAYER M1 ;
        RECT 33.904 23.316 33.936 23.388 ;
  LAYER M2 ;
        RECT 33.884 23.336 33.956 23.368 ;
  LAYER M1 ;
        RECT 33.904 23.352 33.936 23.52 ;
  LAYER M1 ;
        RECT 33.904 23.484 33.936 23.556 ;
  LAYER M2 ;
        RECT 33.884 23.504 33.956 23.536 ;
  LAYER M2 ;
        RECT 31.36 23.504 33.92 23.536 ;
  LAYER M1 ;
        RECT 31.344 23.484 31.376 23.556 ;
  LAYER M2 ;
        RECT 31.324 23.504 31.396 23.536 ;
  LAYER M1 ;
        RECT 33.904 26.256 33.936 26.328 ;
  LAYER M2 ;
        RECT 33.884 26.276 33.956 26.308 ;
  LAYER M1 ;
        RECT 33.904 26.292 33.936 26.46 ;
  LAYER M1 ;
        RECT 33.904 26.424 33.936 26.496 ;
  LAYER M2 ;
        RECT 33.884 26.444 33.956 26.476 ;
  LAYER M2 ;
        RECT 31.36 26.444 33.92 26.476 ;
  LAYER M1 ;
        RECT 31.344 26.424 31.376 26.496 ;
  LAYER M2 ;
        RECT 31.324 26.444 31.396 26.476 ;
  LAYER M1 ;
        RECT 33.904 29.196 33.936 29.268 ;
  LAYER M2 ;
        RECT 33.884 29.216 33.956 29.248 ;
  LAYER M1 ;
        RECT 33.904 29.232 33.936 29.4 ;
  LAYER M1 ;
        RECT 33.904 29.364 33.936 29.436 ;
  LAYER M2 ;
        RECT 33.884 29.384 33.956 29.416 ;
  LAYER M2 ;
        RECT 31.36 29.384 33.92 29.416 ;
  LAYER M1 ;
        RECT 31.344 29.364 31.376 29.436 ;
  LAYER M2 ;
        RECT 31.324 29.384 31.396 29.416 ;
  LAYER M1 ;
        RECT 31.344 29.868 31.376 29.94 ;
  LAYER M2 ;
        RECT 31.324 29.888 31.396 29.92 ;
  LAYER M1 ;
        RECT 31.344 29.568 31.376 29.904 ;
  LAYER M1 ;
        RECT 31.344 20.58 31.376 29.568 ;
  LAYER M2 ;
        RECT 31.36 29.888 45.76 29.92 ;
  LAYER M1 ;
        RECT 42.544 20.376 42.576 20.448 ;
  LAYER M2 ;
        RECT 42.524 20.396 42.596 20.428 ;
  LAYER M2 ;
        RECT 42.56 20.396 45.44 20.428 ;
  LAYER M1 ;
        RECT 45.424 20.376 45.456 20.448 ;
  LAYER M2 ;
        RECT 45.404 20.396 45.476 20.428 ;
  LAYER M1 ;
        RECT 42.544 29.196 42.576 29.268 ;
  LAYER M2 ;
        RECT 42.524 29.216 42.596 29.248 ;
  LAYER M2 ;
        RECT 42.56 29.216 45.44 29.248 ;
  LAYER M1 ;
        RECT 45.424 29.196 45.456 29.268 ;
  LAYER M2 ;
        RECT 45.404 29.216 45.476 29.248 ;
  LAYER M1 ;
        RECT 39.664 29.196 39.696 29.268 ;
  LAYER M2 ;
        RECT 39.644 29.216 39.716 29.248 ;
  LAYER M2 ;
        RECT 39.68 29.216 42.56 29.248 ;
  LAYER M1 ;
        RECT 42.544 29.196 42.576 29.268 ;
  LAYER M2 ;
        RECT 42.524 29.216 42.596 29.248 ;
  LAYER M1 ;
        RECT 36.784 29.196 36.816 29.268 ;
  LAYER M2 ;
        RECT 36.764 29.216 36.836 29.248 ;
  LAYER M2 ;
        RECT 36.8 29.216 39.68 29.248 ;
  LAYER M1 ;
        RECT 39.664 29.196 39.696 29.268 ;
  LAYER M2 ;
        RECT 39.644 29.216 39.716 29.248 ;
  LAYER M1 ;
        RECT 36.784 20.376 36.816 20.448 ;
  LAYER M2 ;
        RECT 36.764 20.396 36.836 20.428 ;
  LAYER M2 ;
        RECT 33.92 20.396 36.8 20.428 ;
  LAYER M1 ;
        RECT 33.904 20.376 33.936 20.448 ;
  LAYER M2 ;
        RECT 33.884 20.396 33.956 20.428 ;
  LAYER M1 ;
        RECT 39.664 20.376 39.696 20.448 ;
  LAYER M2 ;
        RECT 39.644 20.396 39.716 20.428 ;
  LAYER M2 ;
        RECT 36.8 20.396 39.68 20.428 ;
  LAYER M1 ;
        RECT 36.784 20.376 36.816 20.448 ;
  LAYER M2 ;
        RECT 36.764 20.396 36.836 20.428 ;
  LAYER M1 ;
        RECT 43.04 17.976 45.44 20.412 ;
  LAYER M2 ;
        RECT 43.04 17.976 45.44 20.412 ;
  LAYER M3 ;
        RECT 43.04 17.976 45.44 20.412 ;
  LAYER M1 ;
        RECT 43.04 20.916 45.44 23.352 ;
  LAYER M2 ;
        RECT 43.04 20.916 45.44 23.352 ;
  LAYER M3 ;
        RECT 43.04 20.916 45.44 23.352 ;
  LAYER M1 ;
        RECT 43.04 23.856 45.44 26.292 ;
  LAYER M2 ;
        RECT 43.04 23.856 45.44 26.292 ;
  LAYER M3 ;
        RECT 43.04 23.856 45.44 26.292 ;
  LAYER M1 ;
        RECT 43.04 26.796 45.44 29.232 ;
  LAYER M2 ;
        RECT 43.04 26.796 45.44 29.232 ;
  LAYER M3 ;
        RECT 43.04 26.796 45.44 29.232 ;
  LAYER M1 ;
        RECT 40.16 17.976 42.56 20.412 ;
  LAYER M2 ;
        RECT 40.16 17.976 42.56 20.412 ;
  LAYER M3 ;
        RECT 40.16 17.976 42.56 20.412 ;
  LAYER M1 ;
        RECT 40.16 20.916 42.56 23.352 ;
  LAYER M2 ;
        RECT 40.16 20.916 42.56 23.352 ;
  LAYER M3 ;
        RECT 40.16 20.916 42.56 23.352 ;
  LAYER M1 ;
        RECT 40.16 23.856 42.56 26.292 ;
  LAYER M2 ;
        RECT 40.16 23.856 42.56 26.292 ;
  LAYER M3 ;
        RECT 40.16 23.856 42.56 26.292 ;
  LAYER M1 ;
        RECT 40.16 26.796 42.56 29.232 ;
  LAYER M2 ;
        RECT 40.16 26.796 42.56 29.232 ;
  LAYER M3 ;
        RECT 40.16 26.796 42.56 29.232 ;
  LAYER M1 ;
        RECT 37.28 17.976 39.68 20.412 ;
  LAYER M2 ;
        RECT 37.28 17.976 39.68 20.412 ;
  LAYER M3 ;
        RECT 37.28 17.976 39.68 20.412 ;
  LAYER M1 ;
        RECT 37.28 20.916 39.68 23.352 ;
  LAYER M2 ;
        RECT 37.28 20.916 39.68 23.352 ;
  LAYER M3 ;
        RECT 37.28 20.916 39.68 23.352 ;
  LAYER M1 ;
        RECT 37.28 23.856 39.68 26.292 ;
  LAYER M2 ;
        RECT 37.28 23.856 39.68 26.292 ;
  LAYER M3 ;
        RECT 37.28 23.856 39.68 26.292 ;
  LAYER M1 ;
        RECT 37.28 26.796 39.68 29.232 ;
  LAYER M2 ;
        RECT 37.28 26.796 39.68 29.232 ;
  LAYER M3 ;
        RECT 37.28 26.796 39.68 29.232 ;
  LAYER M1 ;
        RECT 34.4 17.976 36.8 20.412 ;
  LAYER M2 ;
        RECT 34.4 17.976 36.8 20.412 ;
  LAYER M3 ;
        RECT 34.4 17.976 36.8 20.412 ;
  LAYER M1 ;
        RECT 34.4 20.916 36.8 23.352 ;
  LAYER M2 ;
        RECT 34.4 20.916 36.8 23.352 ;
  LAYER M3 ;
        RECT 34.4 20.916 36.8 23.352 ;
  LAYER M1 ;
        RECT 34.4 23.856 36.8 26.292 ;
  LAYER M2 ;
        RECT 34.4 23.856 36.8 26.292 ;
  LAYER M3 ;
        RECT 34.4 23.856 36.8 26.292 ;
  LAYER M1 ;
        RECT 34.4 26.796 36.8 29.232 ;
  LAYER M2 ;
        RECT 34.4 26.796 36.8 29.232 ;
  LAYER M3 ;
        RECT 34.4 26.796 36.8 29.232 ;
  LAYER M1 ;
        RECT 31.52 17.976 33.92 20.412 ;
  LAYER M2 ;
        RECT 31.52 17.976 33.92 20.412 ;
  LAYER M3 ;
        RECT 31.52 17.976 33.92 20.412 ;
  LAYER M1 ;
        RECT 31.52 20.916 33.92 23.352 ;
  LAYER M2 ;
        RECT 31.52 20.916 33.92 23.352 ;
  LAYER M3 ;
        RECT 31.52 20.916 33.92 23.352 ;
  LAYER M1 ;
        RECT 31.52 23.856 33.92 26.292 ;
  LAYER M2 ;
        RECT 31.52 23.856 33.92 26.292 ;
  LAYER M3 ;
        RECT 31.52 23.856 33.92 26.292 ;
  LAYER M1 ;
        RECT 31.52 26.796 33.92 29.232 ;
  LAYER M2 ;
        RECT 31.52 26.796 33.92 29.232 ;
  LAYER M3 ;
        RECT 31.52 26.796 33.92 29.232 ;
  LAYER M1 ;
        RECT 40.944 0.3 40.976 0.96 ;
  LAYER M1 ;
        RECT 41.024 0.3 41.056 0.96 ;
  LAYER M1 ;
        RECT 40.864 0.3 40.896 0.96 ;
  LAYER M2 ;
        RECT 40.844 0.908 41.156 0.94 ;
  LAYER M2 ;
        RECT 40.844 0.656 41.156 0.688 ;
  LAYER M2 ;
        RECT 40.764 0.824 41.076 0.856 ;
  LAYER M2 ;
        RECT 40.764 0.572 41.076 0.604 ;
  LAYER M2 ;
        RECT 40.684 0.74 41.076 0.772 ;
  LAYER M2 ;
        RECT 40.684 0.488 41.076 0.52 ;
  LAYER M1 ;
        RECT 30.864 17.352 30.896 18.012 ;
  LAYER M1 ;
        RECT 30.944 17.352 30.976 18.012 ;
  LAYER M1 ;
        RECT 30.784 17.352 30.816 18.012 ;
  LAYER M2 ;
        RECT 30.764 17.96 31.076 17.992 ;
  LAYER M2 ;
        RECT 30.764 17.708 31.076 17.74 ;
  LAYER M2 ;
        RECT 30.684 17.876 30.996 17.908 ;
  LAYER M2 ;
        RECT 30.684 17.624 30.996 17.656 ;
  LAYER M2 ;
        RECT 30.604 17.792 30.996 17.824 ;
  LAYER M2 ;
        RECT 30.604 17.54 30.996 17.572 ;
  LAYER M1 ;
        RECT 39.584 0.3 39.616 0.96 ;
  LAYER M1 ;
        RECT 39.504 0.3 39.536 0.96 ;
  LAYER M1 ;
        RECT 39.664 0.3 39.696 0.96 ;
  LAYER M1 ;
        RECT 40.224 0.3 40.256 0.96 ;
  LAYER M1 ;
        RECT 40.144 0.3 40.176 0.96 ;
  LAYER M1 ;
        RECT 40.304 0.3 40.336 0.96 ;
  LAYER M1 ;
        RECT 38.864 0.3 38.896 0.96 ;
  LAYER M1 ;
        RECT 38.944 0.3 38.976 0.96 ;
  LAYER M1 ;
        RECT 38.784 0.3 38.816 0.96 ;
  LAYER M1 ;
        RECT 38.224 0.3 38.256 0.96 ;
  LAYER M1 ;
        RECT 38.304 0.3 38.336 0.96 ;
  LAYER M1 ;
        RECT 38.144 0.3 38.176 0.96 ;
  LAYER M1 ;
        RECT 39.744 10.296 39.776 10.368 ;
  LAYER M2 ;
        RECT 39.724 10.316 39.796 10.348 ;
  LAYER M2 ;
        RECT 37.04 10.316 39.76 10.348 ;
  LAYER M1 ;
        RECT 37.024 10.296 37.056 10.368 ;
  LAYER M2 ;
        RECT 37.004 10.316 37.076 10.348 ;
  LAYER M1 ;
        RECT 36.864 7.356 36.896 7.428 ;
  LAYER M2 ;
        RECT 36.844 7.376 36.916 7.408 ;
  LAYER M1 ;
        RECT 36.864 7.392 36.896 7.56 ;
  LAYER M1 ;
        RECT 36.864 7.524 36.896 7.596 ;
  LAYER M2 ;
        RECT 36.844 7.544 36.916 7.576 ;
  LAYER M2 ;
        RECT 36.88 7.544 37.04 7.576 ;
  LAYER M1 ;
        RECT 37.024 7.524 37.056 7.596 ;
  LAYER M2 ;
        RECT 37.004 7.544 37.076 7.576 ;
  LAYER M1 ;
        RECT 37.024 16.68 37.056 16.752 ;
  LAYER M2 ;
        RECT 37.004 16.7 37.076 16.732 ;
  LAYER M1 ;
        RECT 37.024 16.548 37.056 16.716 ;
  LAYER M1 ;
        RECT 37.024 7.56 37.056 16.548 ;
  LAYER M1 ;
        RECT 42.624 13.236 42.656 13.308 ;
  LAYER M2 ;
        RECT 42.604 13.256 42.676 13.288 ;
  LAYER M2 ;
        RECT 39.92 13.256 42.64 13.288 ;
  LAYER M1 ;
        RECT 39.904 13.236 39.936 13.308 ;
  LAYER M2 ;
        RECT 39.884 13.256 39.956 13.288 ;
  LAYER M1 ;
        RECT 39.904 16.68 39.936 16.752 ;
  LAYER M2 ;
        RECT 39.884 16.7 39.956 16.732 ;
  LAYER M1 ;
        RECT 39.904 16.548 39.936 16.716 ;
  LAYER M1 ;
        RECT 39.904 13.272 39.936 16.548 ;
  LAYER M2 ;
        RECT 37.04 16.7 39.92 16.732 ;
  LAYER M1 ;
        RECT 36.864 10.296 36.896 10.368 ;
  LAYER M2 ;
        RECT 36.844 10.316 36.916 10.348 ;
  LAYER M2 ;
        RECT 34.16 10.316 36.88 10.348 ;
  LAYER M1 ;
        RECT 34.144 10.296 34.176 10.368 ;
  LAYER M2 ;
        RECT 34.124 10.316 34.196 10.348 ;
  LAYER M1 ;
        RECT 36.864 13.236 36.896 13.308 ;
  LAYER M2 ;
        RECT 36.844 13.256 36.916 13.288 ;
  LAYER M2 ;
        RECT 34.16 13.256 36.88 13.288 ;
  LAYER M1 ;
        RECT 34.144 13.236 34.176 13.308 ;
  LAYER M2 ;
        RECT 34.124 13.256 34.196 13.288 ;
  LAYER M1 ;
        RECT 34.144 16.848 34.176 16.92 ;
  LAYER M2 ;
        RECT 34.124 16.868 34.196 16.9 ;
  LAYER M1 ;
        RECT 34.144 16.548 34.176 16.884 ;
  LAYER M1 ;
        RECT 34.144 10.332 34.176 16.548 ;
  LAYER M1 ;
        RECT 42.624 10.296 42.656 10.368 ;
  LAYER M2 ;
        RECT 42.604 10.316 42.676 10.348 ;
  LAYER M1 ;
        RECT 42.624 10.332 42.656 10.5 ;
  LAYER M1 ;
        RECT 42.624 10.464 42.656 10.536 ;
  LAYER M2 ;
        RECT 42.604 10.484 42.676 10.516 ;
  LAYER M2 ;
        RECT 42.64 10.484 42.8 10.516 ;
  LAYER M1 ;
        RECT 42.784 10.464 42.816 10.536 ;
  LAYER M2 ;
        RECT 42.764 10.484 42.836 10.516 ;
  LAYER M1 ;
        RECT 42.624 7.356 42.656 7.428 ;
  LAYER M2 ;
        RECT 42.604 7.376 42.676 7.408 ;
  LAYER M1 ;
        RECT 42.624 7.392 42.656 7.56 ;
  LAYER M1 ;
        RECT 42.624 7.524 42.656 7.596 ;
  LAYER M2 ;
        RECT 42.604 7.544 42.676 7.576 ;
  LAYER M2 ;
        RECT 42.64 7.544 42.8 7.576 ;
  LAYER M1 ;
        RECT 42.784 7.524 42.816 7.596 ;
  LAYER M2 ;
        RECT 42.764 7.544 42.836 7.576 ;
  LAYER M1 ;
        RECT 42.784 16.848 42.816 16.92 ;
  LAYER M2 ;
        RECT 42.764 16.868 42.836 16.9 ;
  LAYER M1 ;
        RECT 42.784 16.548 42.816 16.884 ;
  LAYER M1 ;
        RECT 42.784 7.56 42.816 16.548 ;
  LAYER M2 ;
        RECT 34.16 16.868 42.8 16.9 ;
  LAYER M1 ;
        RECT 39.744 13.236 39.776 13.308 ;
  LAYER M2 ;
        RECT 39.724 13.256 39.796 13.288 ;
  LAYER M2 ;
        RECT 36.88 13.256 39.76 13.288 ;
  LAYER M1 ;
        RECT 36.864 13.236 36.896 13.308 ;
  LAYER M2 ;
        RECT 36.844 13.256 36.916 13.288 ;
  LAYER M1 ;
        RECT 39.744 7.356 39.776 7.428 ;
  LAYER M2 ;
        RECT 39.724 7.376 39.796 7.408 ;
  LAYER M2 ;
        RECT 39.76 7.376 42.64 7.408 ;
  LAYER M1 ;
        RECT 42.624 7.356 42.656 7.428 ;
  LAYER M2 ;
        RECT 42.604 7.376 42.676 7.408 ;
  LAYER M1 ;
        RECT 33.984 16.176 34.016 16.248 ;
  LAYER M2 ;
        RECT 33.964 16.196 34.036 16.228 ;
  LAYER M2 ;
        RECT 31.28 16.196 34 16.228 ;
  LAYER M1 ;
        RECT 31.264 16.176 31.296 16.248 ;
  LAYER M2 ;
        RECT 31.244 16.196 31.316 16.228 ;
  LAYER M1 ;
        RECT 33.984 13.236 34.016 13.308 ;
  LAYER M2 ;
        RECT 33.964 13.256 34.036 13.288 ;
  LAYER M2 ;
        RECT 31.28 13.256 34 13.288 ;
  LAYER M1 ;
        RECT 31.264 13.236 31.296 13.308 ;
  LAYER M2 ;
        RECT 31.244 13.256 31.316 13.288 ;
  LAYER M1 ;
        RECT 33.984 10.296 34.016 10.368 ;
  LAYER M2 ;
        RECT 33.964 10.316 34.036 10.348 ;
  LAYER M2 ;
        RECT 31.28 10.316 34 10.348 ;
  LAYER M1 ;
        RECT 31.264 10.296 31.296 10.368 ;
  LAYER M2 ;
        RECT 31.244 10.316 31.316 10.348 ;
  LAYER M1 ;
        RECT 33.984 7.356 34.016 7.428 ;
  LAYER M2 ;
        RECT 33.964 7.376 34.036 7.408 ;
  LAYER M2 ;
        RECT 31.28 7.376 34 7.408 ;
  LAYER M1 ;
        RECT 31.264 7.356 31.296 7.428 ;
  LAYER M2 ;
        RECT 31.244 7.376 31.316 7.408 ;
  LAYER M1 ;
        RECT 33.984 4.416 34.016 4.488 ;
  LAYER M2 ;
        RECT 33.964 4.436 34.036 4.468 ;
  LAYER M2 ;
        RECT 31.28 4.436 34 4.468 ;
  LAYER M1 ;
        RECT 31.264 4.416 31.296 4.488 ;
  LAYER M2 ;
        RECT 31.244 4.436 31.316 4.468 ;
  LAYER M1 ;
        RECT 31.264 17.016 31.296 17.088 ;
  LAYER M2 ;
        RECT 31.244 17.036 31.316 17.068 ;
  LAYER M1 ;
        RECT 31.264 16.548 31.296 17.052 ;
  LAYER M1 ;
        RECT 31.264 4.452 31.296 16.548 ;
  LAYER M1 ;
        RECT 45.504 16.176 45.536 16.248 ;
  LAYER M2 ;
        RECT 45.484 16.196 45.556 16.228 ;
  LAYER M1 ;
        RECT 45.504 16.212 45.536 16.38 ;
  LAYER M1 ;
        RECT 45.504 16.344 45.536 16.416 ;
  LAYER M2 ;
        RECT 45.484 16.364 45.556 16.396 ;
  LAYER M2 ;
        RECT 45.52 16.364 45.68 16.396 ;
  LAYER M1 ;
        RECT 45.664 16.344 45.696 16.416 ;
  LAYER M2 ;
        RECT 45.644 16.364 45.716 16.396 ;
  LAYER M1 ;
        RECT 45.504 13.236 45.536 13.308 ;
  LAYER M2 ;
        RECT 45.484 13.256 45.556 13.288 ;
  LAYER M1 ;
        RECT 45.504 13.272 45.536 13.44 ;
  LAYER M1 ;
        RECT 45.504 13.404 45.536 13.476 ;
  LAYER M2 ;
        RECT 45.484 13.424 45.556 13.456 ;
  LAYER M2 ;
        RECT 45.52 13.424 45.68 13.456 ;
  LAYER M1 ;
        RECT 45.664 13.404 45.696 13.476 ;
  LAYER M2 ;
        RECT 45.644 13.424 45.716 13.456 ;
  LAYER M1 ;
        RECT 45.504 10.296 45.536 10.368 ;
  LAYER M2 ;
        RECT 45.484 10.316 45.556 10.348 ;
  LAYER M1 ;
        RECT 45.504 10.332 45.536 10.5 ;
  LAYER M1 ;
        RECT 45.504 10.464 45.536 10.536 ;
  LAYER M2 ;
        RECT 45.484 10.484 45.556 10.516 ;
  LAYER M2 ;
        RECT 45.52 10.484 45.68 10.516 ;
  LAYER M1 ;
        RECT 45.664 10.464 45.696 10.536 ;
  LAYER M2 ;
        RECT 45.644 10.484 45.716 10.516 ;
  LAYER M1 ;
        RECT 45.504 7.356 45.536 7.428 ;
  LAYER M2 ;
        RECT 45.484 7.376 45.556 7.408 ;
  LAYER M1 ;
        RECT 45.504 7.392 45.536 7.56 ;
  LAYER M1 ;
        RECT 45.504 7.524 45.536 7.596 ;
  LAYER M2 ;
        RECT 45.484 7.544 45.556 7.576 ;
  LAYER M2 ;
        RECT 45.52 7.544 45.68 7.576 ;
  LAYER M1 ;
        RECT 45.664 7.524 45.696 7.596 ;
  LAYER M2 ;
        RECT 45.644 7.544 45.716 7.576 ;
  LAYER M1 ;
        RECT 45.504 4.416 45.536 4.488 ;
  LAYER M2 ;
        RECT 45.484 4.436 45.556 4.468 ;
  LAYER M1 ;
        RECT 45.504 4.452 45.536 4.62 ;
  LAYER M1 ;
        RECT 45.504 4.584 45.536 4.656 ;
  LAYER M2 ;
        RECT 45.484 4.604 45.556 4.636 ;
  LAYER M2 ;
        RECT 45.52 4.604 45.68 4.636 ;
  LAYER M1 ;
        RECT 45.664 4.584 45.696 4.656 ;
  LAYER M2 ;
        RECT 45.644 4.604 45.716 4.636 ;
  LAYER M1 ;
        RECT 45.664 17.016 45.696 17.088 ;
  LAYER M2 ;
        RECT 45.644 17.036 45.716 17.068 ;
  LAYER M1 ;
        RECT 45.664 16.548 45.696 17.052 ;
  LAYER M1 ;
        RECT 45.664 4.62 45.696 16.548 ;
  LAYER M2 ;
        RECT 31.28 17.036 45.68 17.068 ;
  LAYER M1 ;
        RECT 36.864 16.176 36.896 16.248 ;
  LAYER M2 ;
        RECT 36.844 16.196 36.916 16.228 ;
  LAYER M2 ;
        RECT 34 16.196 36.88 16.228 ;
  LAYER M1 ;
        RECT 33.984 16.176 34.016 16.248 ;
  LAYER M2 ;
        RECT 33.964 16.196 34.036 16.228 ;
  LAYER M1 ;
        RECT 36.864 4.416 36.896 4.488 ;
  LAYER M2 ;
        RECT 36.844 4.436 36.916 4.468 ;
  LAYER M2 ;
        RECT 34 4.436 36.88 4.468 ;
  LAYER M1 ;
        RECT 33.984 4.416 34.016 4.488 ;
  LAYER M2 ;
        RECT 33.964 4.436 34.036 4.468 ;
  LAYER M1 ;
        RECT 39.744 4.416 39.776 4.488 ;
  LAYER M2 ;
        RECT 39.724 4.436 39.796 4.468 ;
  LAYER M2 ;
        RECT 36.88 4.436 39.76 4.468 ;
  LAYER M1 ;
        RECT 36.864 4.416 36.896 4.488 ;
  LAYER M2 ;
        RECT 36.844 4.436 36.916 4.468 ;
  LAYER M1 ;
        RECT 42.624 4.416 42.656 4.488 ;
  LAYER M2 ;
        RECT 42.604 4.436 42.676 4.468 ;
  LAYER M2 ;
        RECT 39.76 4.436 42.64 4.468 ;
  LAYER M1 ;
        RECT 39.744 4.416 39.776 4.488 ;
  LAYER M2 ;
        RECT 39.724 4.436 39.796 4.468 ;
  LAYER M1 ;
        RECT 42.624 16.176 42.656 16.248 ;
  LAYER M2 ;
        RECT 42.604 16.196 42.676 16.228 ;
  LAYER M2 ;
        RECT 42.64 16.196 45.52 16.228 ;
  LAYER M1 ;
        RECT 45.504 16.176 45.536 16.248 ;
  LAYER M2 ;
        RECT 45.484 16.196 45.556 16.228 ;
  LAYER M1 ;
        RECT 39.744 16.176 39.776 16.248 ;
  LAYER M2 ;
        RECT 39.724 16.196 39.796 16.228 ;
  LAYER M2 ;
        RECT 39.76 16.196 42.64 16.228 ;
  LAYER M1 ;
        RECT 42.624 16.176 42.656 16.248 ;
  LAYER M2 ;
        RECT 42.604 16.196 42.676 16.228 ;
  LAYER M1 ;
        RECT 37.344 7.86 37.376 7.932 ;
  LAYER M2 ;
        RECT 37.324 7.88 37.396 7.912 ;
  LAYER M2 ;
        RECT 37.2 7.88 37.36 7.912 ;
  LAYER M1 ;
        RECT 37.184 7.86 37.216 7.932 ;
  LAYER M2 ;
        RECT 37.164 7.88 37.236 7.912 ;
  LAYER M1 ;
        RECT 34.464 4.92 34.496 4.992 ;
  LAYER M2 ;
        RECT 34.444 4.94 34.516 4.972 ;
  LAYER M1 ;
        RECT 34.464 4.788 34.496 4.956 ;
  LAYER M1 ;
        RECT 34.464 4.752 34.496 4.824 ;
  LAYER M2 ;
        RECT 34.444 4.772 34.516 4.804 ;
  LAYER M2 ;
        RECT 34.48 4.772 37.2 4.804 ;
  LAYER M1 ;
        RECT 37.184 4.752 37.216 4.824 ;
  LAYER M2 ;
        RECT 37.164 4.772 37.236 4.804 ;
  LAYER M1 ;
        RECT 37.184 1.476 37.216 1.548 ;
  LAYER M2 ;
        RECT 37.164 1.496 37.236 1.528 ;
  LAYER M1 ;
        RECT 37.184 1.512 37.216 1.68 ;
  LAYER M1 ;
        RECT 37.184 1.68 37.216 7.896 ;
  LAYER M1 ;
        RECT 40.224 10.8 40.256 10.872 ;
  LAYER M2 ;
        RECT 40.204 10.82 40.276 10.852 ;
  LAYER M2 ;
        RECT 40.08 10.82 40.24 10.852 ;
  LAYER M1 ;
        RECT 40.064 10.8 40.096 10.872 ;
  LAYER M2 ;
        RECT 40.044 10.82 40.116 10.852 ;
  LAYER M1 ;
        RECT 40.064 1.476 40.096 1.548 ;
  LAYER M2 ;
        RECT 40.044 1.496 40.116 1.528 ;
  LAYER M1 ;
        RECT 40.064 1.512 40.096 1.68 ;
  LAYER M1 ;
        RECT 40.064 1.68 40.096 10.836 ;
  LAYER M2 ;
        RECT 37.2 1.496 40.08 1.528 ;
  LAYER M1 ;
        RECT 34.464 7.86 34.496 7.932 ;
  LAYER M2 ;
        RECT 34.444 7.88 34.516 7.912 ;
  LAYER M2 ;
        RECT 34.32 7.88 34.48 7.912 ;
  LAYER M1 ;
        RECT 34.304 7.86 34.336 7.932 ;
  LAYER M2 ;
        RECT 34.284 7.88 34.356 7.912 ;
  LAYER M1 ;
        RECT 34.464 10.8 34.496 10.872 ;
  LAYER M2 ;
        RECT 34.444 10.82 34.516 10.852 ;
  LAYER M2 ;
        RECT 34.32 10.82 34.48 10.852 ;
  LAYER M1 ;
        RECT 34.304 10.8 34.336 10.872 ;
  LAYER M2 ;
        RECT 34.284 10.82 34.356 10.852 ;
  LAYER M1 ;
        RECT 34.304 1.308 34.336 1.38 ;
  LAYER M2 ;
        RECT 34.284 1.328 34.356 1.36 ;
  LAYER M1 ;
        RECT 34.304 1.344 34.336 1.68 ;
  LAYER M1 ;
        RECT 34.304 1.68 34.336 10.836 ;
  LAYER M1 ;
        RECT 40.224 7.86 40.256 7.932 ;
  LAYER M2 ;
        RECT 40.204 7.88 40.276 7.912 ;
  LAYER M1 ;
        RECT 40.224 7.728 40.256 7.896 ;
  LAYER M1 ;
        RECT 40.224 7.692 40.256 7.764 ;
  LAYER M2 ;
        RECT 40.204 7.712 40.276 7.744 ;
  LAYER M2 ;
        RECT 40.24 7.712 42.96 7.744 ;
  LAYER M1 ;
        RECT 42.944 7.692 42.976 7.764 ;
  LAYER M2 ;
        RECT 42.924 7.712 42.996 7.744 ;
  LAYER M1 ;
        RECT 40.224 4.92 40.256 4.992 ;
  LAYER M2 ;
        RECT 40.204 4.94 40.276 4.972 ;
  LAYER M1 ;
        RECT 40.224 4.788 40.256 4.956 ;
  LAYER M1 ;
        RECT 40.224 4.752 40.256 4.824 ;
  LAYER M2 ;
        RECT 40.204 4.772 40.276 4.804 ;
  LAYER M2 ;
        RECT 40.24 4.772 42.96 4.804 ;
  LAYER M1 ;
        RECT 42.944 4.752 42.976 4.824 ;
  LAYER M2 ;
        RECT 42.924 4.772 42.996 4.804 ;
  LAYER M1 ;
        RECT 42.944 1.308 42.976 1.38 ;
  LAYER M2 ;
        RECT 42.924 1.328 42.996 1.36 ;
  LAYER M1 ;
        RECT 42.944 1.344 42.976 1.68 ;
  LAYER M1 ;
        RECT 42.944 1.68 42.976 7.728 ;
  LAYER M2 ;
        RECT 34.32 1.328 42.96 1.36 ;
  LAYER M1 ;
        RECT 37.344 10.8 37.376 10.872 ;
  LAYER M2 ;
        RECT 37.324 10.82 37.396 10.852 ;
  LAYER M2 ;
        RECT 34.48 10.82 37.36 10.852 ;
  LAYER M1 ;
        RECT 34.464 10.8 34.496 10.872 ;
  LAYER M2 ;
        RECT 34.444 10.82 34.516 10.852 ;
  LAYER M1 ;
        RECT 37.344 4.92 37.376 4.992 ;
  LAYER M2 ;
        RECT 37.324 4.94 37.396 4.972 ;
  LAYER M2 ;
        RECT 37.36 4.94 40.24 4.972 ;
  LAYER M1 ;
        RECT 40.224 4.92 40.256 4.992 ;
  LAYER M2 ;
        RECT 40.204 4.94 40.276 4.972 ;
  LAYER M1 ;
        RECT 31.584 13.74 31.616 13.812 ;
  LAYER M2 ;
        RECT 31.564 13.76 31.636 13.792 ;
  LAYER M2 ;
        RECT 31.44 13.76 31.6 13.792 ;
  LAYER M1 ;
        RECT 31.424 13.74 31.456 13.812 ;
  LAYER M2 ;
        RECT 31.404 13.76 31.476 13.792 ;
  LAYER M1 ;
        RECT 31.584 10.8 31.616 10.872 ;
  LAYER M2 ;
        RECT 31.564 10.82 31.636 10.852 ;
  LAYER M2 ;
        RECT 31.44 10.82 31.6 10.852 ;
  LAYER M1 ;
        RECT 31.424 10.8 31.456 10.872 ;
  LAYER M2 ;
        RECT 31.404 10.82 31.476 10.852 ;
  LAYER M1 ;
        RECT 31.584 7.86 31.616 7.932 ;
  LAYER M2 ;
        RECT 31.564 7.88 31.636 7.912 ;
  LAYER M2 ;
        RECT 31.44 7.88 31.6 7.912 ;
  LAYER M1 ;
        RECT 31.424 7.86 31.456 7.932 ;
  LAYER M2 ;
        RECT 31.404 7.88 31.476 7.912 ;
  LAYER M1 ;
        RECT 31.584 4.92 31.616 4.992 ;
  LAYER M2 ;
        RECT 31.564 4.94 31.636 4.972 ;
  LAYER M2 ;
        RECT 31.44 4.94 31.6 4.972 ;
  LAYER M1 ;
        RECT 31.424 4.92 31.456 4.992 ;
  LAYER M2 ;
        RECT 31.404 4.94 31.476 4.972 ;
  LAYER M1 ;
        RECT 31.584 1.98 31.616 2.052 ;
  LAYER M2 ;
        RECT 31.564 2 31.636 2.032 ;
  LAYER M2 ;
        RECT 31.44 2 31.6 2.032 ;
  LAYER M1 ;
        RECT 31.424 1.98 31.456 2.052 ;
  LAYER M2 ;
        RECT 31.404 2 31.476 2.032 ;
  LAYER M1 ;
        RECT 31.424 1.14 31.456 1.212 ;
  LAYER M2 ;
        RECT 31.404 1.16 31.476 1.192 ;
  LAYER M1 ;
        RECT 31.424 1.176 31.456 1.68 ;
  LAYER M1 ;
        RECT 31.424 1.68 31.456 13.776 ;
  LAYER M1 ;
        RECT 43.104 13.74 43.136 13.812 ;
  LAYER M2 ;
        RECT 43.084 13.76 43.156 13.792 ;
  LAYER M1 ;
        RECT 43.104 13.608 43.136 13.776 ;
  LAYER M1 ;
        RECT 43.104 13.572 43.136 13.644 ;
  LAYER M2 ;
        RECT 43.084 13.592 43.156 13.624 ;
  LAYER M2 ;
        RECT 43.12 13.592 45.84 13.624 ;
  LAYER M1 ;
        RECT 45.824 13.572 45.856 13.644 ;
  LAYER M2 ;
        RECT 45.804 13.592 45.876 13.624 ;
  LAYER M1 ;
        RECT 43.104 10.8 43.136 10.872 ;
  LAYER M2 ;
        RECT 43.084 10.82 43.156 10.852 ;
  LAYER M1 ;
        RECT 43.104 10.668 43.136 10.836 ;
  LAYER M1 ;
        RECT 43.104 10.632 43.136 10.704 ;
  LAYER M2 ;
        RECT 43.084 10.652 43.156 10.684 ;
  LAYER M2 ;
        RECT 43.12 10.652 45.84 10.684 ;
  LAYER M1 ;
        RECT 45.824 10.632 45.856 10.704 ;
  LAYER M2 ;
        RECT 45.804 10.652 45.876 10.684 ;
  LAYER M1 ;
        RECT 43.104 7.86 43.136 7.932 ;
  LAYER M2 ;
        RECT 43.084 7.88 43.156 7.912 ;
  LAYER M1 ;
        RECT 43.104 7.728 43.136 7.896 ;
  LAYER M1 ;
        RECT 43.104 7.692 43.136 7.764 ;
  LAYER M2 ;
        RECT 43.084 7.712 43.156 7.744 ;
  LAYER M2 ;
        RECT 43.12 7.712 45.84 7.744 ;
  LAYER M1 ;
        RECT 45.824 7.692 45.856 7.764 ;
  LAYER M2 ;
        RECT 45.804 7.712 45.876 7.744 ;
  LAYER M1 ;
        RECT 43.104 4.92 43.136 4.992 ;
  LAYER M2 ;
        RECT 43.084 4.94 43.156 4.972 ;
  LAYER M1 ;
        RECT 43.104 4.788 43.136 4.956 ;
  LAYER M1 ;
        RECT 43.104 4.752 43.136 4.824 ;
  LAYER M2 ;
        RECT 43.084 4.772 43.156 4.804 ;
  LAYER M2 ;
        RECT 43.12 4.772 45.84 4.804 ;
  LAYER M1 ;
        RECT 45.824 4.752 45.856 4.824 ;
  LAYER M2 ;
        RECT 45.804 4.772 45.876 4.804 ;
  LAYER M1 ;
        RECT 43.104 1.98 43.136 2.052 ;
  LAYER M2 ;
        RECT 43.084 2 43.156 2.032 ;
  LAYER M1 ;
        RECT 43.104 1.848 43.136 2.016 ;
  LAYER M1 ;
        RECT 43.104 1.812 43.136 1.884 ;
  LAYER M2 ;
        RECT 43.084 1.832 43.156 1.864 ;
  LAYER M2 ;
        RECT 43.12 1.832 45.84 1.864 ;
  LAYER M1 ;
        RECT 45.824 1.812 45.856 1.884 ;
  LAYER M2 ;
        RECT 45.804 1.832 45.876 1.864 ;
  LAYER M1 ;
        RECT 45.824 1.14 45.856 1.212 ;
  LAYER M2 ;
        RECT 45.804 1.16 45.876 1.192 ;
  LAYER M1 ;
        RECT 45.824 1.176 45.856 1.68 ;
  LAYER M1 ;
        RECT 45.824 1.68 45.856 13.608 ;
  LAYER M2 ;
        RECT 31.44 1.16 45.84 1.192 ;
  LAYER M1 ;
        RECT 34.464 13.74 34.496 13.812 ;
  LAYER M2 ;
        RECT 34.444 13.76 34.516 13.792 ;
  LAYER M2 ;
        RECT 31.6 13.76 34.48 13.792 ;
  LAYER M1 ;
        RECT 31.584 13.74 31.616 13.812 ;
  LAYER M2 ;
        RECT 31.564 13.76 31.636 13.792 ;
  LAYER M1 ;
        RECT 34.464 1.98 34.496 2.052 ;
  LAYER M2 ;
        RECT 34.444 2 34.516 2.032 ;
  LAYER M2 ;
        RECT 31.6 2 34.48 2.032 ;
  LAYER M1 ;
        RECT 31.584 1.98 31.616 2.052 ;
  LAYER M2 ;
        RECT 31.564 2 31.636 2.032 ;
  LAYER M1 ;
        RECT 37.344 1.98 37.376 2.052 ;
  LAYER M2 ;
        RECT 37.324 2 37.396 2.032 ;
  LAYER M2 ;
        RECT 34.48 2 37.36 2.032 ;
  LAYER M1 ;
        RECT 34.464 1.98 34.496 2.052 ;
  LAYER M2 ;
        RECT 34.444 2 34.516 2.032 ;
  LAYER M1 ;
        RECT 40.224 1.98 40.256 2.052 ;
  LAYER M2 ;
        RECT 40.204 2 40.276 2.032 ;
  LAYER M2 ;
        RECT 37.36 2 40.24 2.032 ;
  LAYER M1 ;
        RECT 37.344 1.98 37.376 2.052 ;
  LAYER M2 ;
        RECT 37.324 2 37.396 2.032 ;
  LAYER M1 ;
        RECT 40.224 13.74 40.256 13.812 ;
  LAYER M2 ;
        RECT 40.204 13.76 40.276 13.792 ;
  LAYER M2 ;
        RECT 40.24 13.76 43.12 13.792 ;
  LAYER M1 ;
        RECT 43.104 13.74 43.136 13.812 ;
  LAYER M2 ;
        RECT 43.084 13.76 43.156 13.792 ;
  LAYER M1 ;
        RECT 37.344 13.74 37.376 13.812 ;
  LAYER M2 ;
        RECT 37.324 13.76 37.396 13.792 ;
  LAYER M2 ;
        RECT 37.36 13.76 40.24 13.792 ;
  LAYER M1 ;
        RECT 40.224 13.74 40.256 13.812 ;
  LAYER M2 ;
        RECT 40.204 13.76 40.276 13.792 ;
  LAYER M1 ;
        RECT 31.6 13.776 34 16.212 ;
  LAYER M2 ;
        RECT 31.6 13.776 34 16.212 ;
  LAYER M3 ;
        RECT 31.6 13.776 34 16.212 ;
  LAYER M1 ;
        RECT 31.6 10.836 34 13.272 ;
  LAYER M2 ;
        RECT 31.6 10.836 34 13.272 ;
  LAYER M3 ;
        RECT 31.6 10.836 34 13.272 ;
  LAYER M1 ;
        RECT 31.6 7.896 34 10.332 ;
  LAYER M2 ;
        RECT 31.6 7.896 34 10.332 ;
  LAYER M3 ;
        RECT 31.6 7.896 34 10.332 ;
  LAYER M1 ;
        RECT 31.6 4.956 34 7.392 ;
  LAYER M2 ;
        RECT 31.6 4.956 34 7.392 ;
  LAYER M3 ;
        RECT 31.6 4.956 34 7.392 ;
  LAYER M1 ;
        RECT 31.6 2.016 34 4.452 ;
  LAYER M2 ;
        RECT 31.6 2.016 34 4.452 ;
  LAYER M3 ;
        RECT 31.6 2.016 34 4.452 ;
  LAYER M1 ;
        RECT 34.48 13.776 36.88 16.212 ;
  LAYER M2 ;
        RECT 34.48 13.776 36.88 16.212 ;
  LAYER M3 ;
        RECT 34.48 13.776 36.88 16.212 ;
  LAYER M1 ;
        RECT 34.48 10.836 36.88 13.272 ;
  LAYER M2 ;
        RECT 34.48 10.836 36.88 13.272 ;
  LAYER M3 ;
        RECT 34.48 10.836 36.88 13.272 ;
  LAYER M1 ;
        RECT 34.48 7.896 36.88 10.332 ;
  LAYER M2 ;
        RECT 34.48 7.896 36.88 10.332 ;
  LAYER M3 ;
        RECT 34.48 7.896 36.88 10.332 ;
  LAYER M1 ;
        RECT 34.48 4.956 36.88 7.392 ;
  LAYER M2 ;
        RECT 34.48 4.956 36.88 7.392 ;
  LAYER M3 ;
        RECT 34.48 4.956 36.88 7.392 ;
  LAYER M1 ;
        RECT 34.48 2.016 36.88 4.452 ;
  LAYER M2 ;
        RECT 34.48 2.016 36.88 4.452 ;
  LAYER M3 ;
        RECT 34.48 2.016 36.88 4.452 ;
  LAYER M1 ;
        RECT 37.36 13.776 39.76 16.212 ;
  LAYER M2 ;
        RECT 37.36 13.776 39.76 16.212 ;
  LAYER M3 ;
        RECT 37.36 13.776 39.76 16.212 ;
  LAYER M1 ;
        RECT 37.36 10.836 39.76 13.272 ;
  LAYER M2 ;
        RECT 37.36 10.836 39.76 13.272 ;
  LAYER M3 ;
        RECT 37.36 10.836 39.76 13.272 ;
  LAYER M1 ;
        RECT 37.36 7.896 39.76 10.332 ;
  LAYER M2 ;
        RECT 37.36 7.896 39.76 10.332 ;
  LAYER M3 ;
        RECT 37.36 7.896 39.76 10.332 ;
  LAYER M1 ;
        RECT 37.36 4.956 39.76 7.392 ;
  LAYER M2 ;
        RECT 37.36 4.956 39.76 7.392 ;
  LAYER M3 ;
        RECT 37.36 4.956 39.76 7.392 ;
  LAYER M1 ;
        RECT 37.36 2.016 39.76 4.452 ;
  LAYER M2 ;
        RECT 37.36 2.016 39.76 4.452 ;
  LAYER M3 ;
        RECT 37.36 2.016 39.76 4.452 ;
  LAYER M1 ;
        RECT 40.24 13.776 42.64 16.212 ;
  LAYER M2 ;
        RECT 40.24 13.776 42.64 16.212 ;
  LAYER M3 ;
        RECT 40.24 13.776 42.64 16.212 ;
  LAYER M1 ;
        RECT 40.24 10.836 42.64 13.272 ;
  LAYER M2 ;
        RECT 40.24 10.836 42.64 13.272 ;
  LAYER M3 ;
        RECT 40.24 10.836 42.64 13.272 ;
  LAYER M1 ;
        RECT 40.24 7.896 42.64 10.332 ;
  LAYER M2 ;
        RECT 40.24 7.896 42.64 10.332 ;
  LAYER M3 ;
        RECT 40.24 7.896 42.64 10.332 ;
  LAYER M1 ;
        RECT 40.24 4.956 42.64 7.392 ;
  LAYER M2 ;
        RECT 40.24 4.956 42.64 7.392 ;
  LAYER M3 ;
        RECT 40.24 4.956 42.64 7.392 ;
  LAYER M1 ;
        RECT 40.24 2.016 42.64 4.452 ;
  LAYER M2 ;
        RECT 40.24 2.016 42.64 4.452 ;
  LAYER M3 ;
        RECT 40.24 2.016 42.64 4.452 ;
  LAYER M1 ;
        RECT 43.12 13.776 45.52 16.212 ;
  LAYER M2 ;
        RECT 43.12 13.776 45.52 16.212 ;
  LAYER M3 ;
        RECT 43.12 13.776 45.52 16.212 ;
  LAYER M1 ;
        RECT 43.12 10.836 45.52 13.272 ;
  LAYER M2 ;
        RECT 43.12 10.836 45.52 13.272 ;
  LAYER M3 ;
        RECT 43.12 10.836 45.52 13.272 ;
  LAYER M1 ;
        RECT 43.12 7.896 45.52 10.332 ;
  LAYER M2 ;
        RECT 43.12 7.896 45.52 10.332 ;
  LAYER M3 ;
        RECT 43.12 7.896 45.52 10.332 ;
  LAYER M1 ;
        RECT 43.12 4.956 45.52 7.392 ;
  LAYER M2 ;
        RECT 43.12 4.956 45.52 7.392 ;
  LAYER M3 ;
        RECT 43.12 4.956 45.52 7.392 ;
  LAYER M1 ;
        RECT 43.12 2.016 45.52 4.452 ;
  LAYER M2 ;
        RECT 43.12 2.016 45.52 4.452 ;
  LAYER M3 ;
        RECT 43.12 2.016 45.52 4.452 ;
  LAYER M1 ;
        RECT 21.824 11.892 21.856 11.964 ;
  LAYER M2 ;
        RECT 21.804 11.912 21.876 11.944 ;
  LAYER M2 ;
        RECT 21.84 11.912 24.56 11.944 ;
  LAYER M1 ;
        RECT 24.544 11.892 24.576 11.964 ;
  LAYER M2 ;
        RECT 24.524 11.912 24.596 11.944 ;
  LAYER M1 ;
        RECT 24.704 14.832 24.736 14.904 ;
  LAYER M2 ;
        RECT 24.684 14.852 24.756 14.884 ;
  LAYER M1 ;
        RECT 24.704 14.868 24.736 15.036 ;
  LAYER M1 ;
        RECT 24.704 15 24.736 15.072 ;
  LAYER M2 ;
        RECT 24.684 15.02 24.756 15.052 ;
  LAYER M2 ;
        RECT 24.56 15.02 24.72 15.052 ;
  LAYER M1 ;
        RECT 24.544 15 24.576 15.072 ;
  LAYER M2 ;
        RECT 24.524 15.02 24.596 15.052 ;
  LAYER M1 ;
        RECT 24.544 18.276 24.576 18.348 ;
  LAYER M2 ;
        RECT 24.524 18.296 24.596 18.328 ;
  LAYER M1 ;
        RECT 24.544 18.144 24.576 18.312 ;
  LAYER M1 ;
        RECT 24.544 11.928 24.576 18.144 ;
  LAYER M1 ;
        RECT 18.944 11.892 18.976 11.964 ;
  LAYER M2 ;
        RECT 18.924 11.912 18.996 11.944 ;
  LAYER M2 ;
        RECT 18.96 11.912 21.68 11.944 ;
  LAYER M1 ;
        RECT 21.664 11.892 21.696 11.964 ;
  LAYER M2 ;
        RECT 21.644 11.912 21.716 11.944 ;
  LAYER M1 ;
        RECT 21.664 18.276 21.696 18.348 ;
  LAYER M2 ;
        RECT 21.644 18.296 21.716 18.328 ;
  LAYER M1 ;
        RECT 21.664 18.144 21.696 18.312 ;
  LAYER M1 ;
        RECT 21.664 11.928 21.696 18.144 ;
  LAYER M2 ;
        RECT 21.68 18.296 24.56 18.328 ;
  LAYER M1 ;
        RECT 24.704 11.892 24.736 11.964 ;
  LAYER M2 ;
        RECT 24.684 11.912 24.756 11.944 ;
  LAYER M2 ;
        RECT 24.72 11.912 27.44 11.944 ;
  LAYER M1 ;
        RECT 27.424 11.892 27.456 11.964 ;
  LAYER M2 ;
        RECT 27.404 11.912 27.476 11.944 ;
  LAYER M1 ;
        RECT 27.424 18.444 27.456 18.516 ;
  LAYER M2 ;
        RECT 27.404 18.464 27.476 18.496 ;
  LAYER M1 ;
        RECT 27.424 18.144 27.456 18.48 ;
  LAYER M1 ;
        RECT 27.424 11.928 27.456 18.144 ;
  LAYER M1 ;
        RECT 18.944 14.832 18.976 14.904 ;
  LAYER M2 ;
        RECT 18.924 14.852 18.996 14.884 ;
  LAYER M1 ;
        RECT 18.944 14.868 18.976 15.036 ;
  LAYER M1 ;
        RECT 18.944 15 18.976 15.072 ;
  LAYER M2 ;
        RECT 18.924 15.02 18.996 15.052 ;
  LAYER M2 ;
        RECT 18.8 15.02 18.96 15.052 ;
  LAYER M1 ;
        RECT 18.784 15 18.816 15.072 ;
  LAYER M2 ;
        RECT 18.764 15.02 18.836 15.052 ;
  LAYER M1 ;
        RECT 18.784 18.444 18.816 18.516 ;
  LAYER M2 ;
        RECT 18.764 18.464 18.836 18.496 ;
  LAYER M1 ;
        RECT 18.784 18.144 18.816 18.48 ;
  LAYER M1 ;
        RECT 18.784 15.036 18.816 18.144 ;
  LAYER M2 ;
        RECT 18.8 18.464 27.44 18.496 ;
  LAYER M1 ;
        RECT 21.824 14.832 21.856 14.904 ;
  LAYER M2 ;
        RECT 21.804 14.852 21.876 14.884 ;
  LAYER M2 ;
        RECT 18.96 14.852 21.84 14.884 ;
  LAYER M1 ;
        RECT 18.944 14.832 18.976 14.904 ;
  LAYER M2 ;
        RECT 18.924 14.852 18.996 14.884 ;
  LAYER M1 ;
        RECT 27.584 17.772 27.616 17.844 ;
  LAYER M2 ;
        RECT 27.564 17.792 27.636 17.824 ;
  LAYER M2 ;
        RECT 27.6 17.792 30.32 17.824 ;
  LAYER M1 ;
        RECT 30.304 17.772 30.336 17.844 ;
  LAYER M2 ;
        RECT 30.284 17.792 30.356 17.824 ;
  LAYER M1 ;
        RECT 27.584 14.832 27.616 14.904 ;
  LAYER M2 ;
        RECT 27.564 14.852 27.636 14.884 ;
  LAYER M2 ;
        RECT 27.6 14.852 30.32 14.884 ;
  LAYER M1 ;
        RECT 30.304 14.832 30.336 14.904 ;
  LAYER M2 ;
        RECT 30.284 14.852 30.356 14.884 ;
  LAYER M1 ;
        RECT 27.584 11.892 27.616 11.964 ;
  LAYER M2 ;
        RECT 27.564 11.912 27.636 11.944 ;
  LAYER M2 ;
        RECT 27.6 11.912 30.32 11.944 ;
  LAYER M1 ;
        RECT 30.304 11.892 30.336 11.964 ;
  LAYER M2 ;
        RECT 30.284 11.912 30.356 11.944 ;
  LAYER M1 ;
        RECT 27.584 8.952 27.616 9.024 ;
  LAYER M2 ;
        RECT 27.564 8.972 27.636 9.004 ;
  LAYER M2 ;
        RECT 27.6 8.972 30.32 9.004 ;
  LAYER M1 ;
        RECT 30.304 8.952 30.336 9.024 ;
  LAYER M2 ;
        RECT 30.284 8.972 30.356 9.004 ;
  LAYER M1 ;
        RECT 30.304 18.612 30.336 18.684 ;
  LAYER M2 ;
        RECT 30.284 18.632 30.356 18.664 ;
  LAYER M1 ;
        RECT 30.304 18.144 30.336 18.648 ;
  LAYER M1 ;
        RECT 30.304 8.988 30.336 18.144 ;
  LAYER M1 ;
        RECT 16.064 17.772 16.096 17.844 ;
  LAYER M2 ;
        RECT 16.044 17.792 16.116 17.824 ;
  LAYER M1 ;
        RECT 16.064 17.808 16.096 17.976 ;
  LAYER M1 ;
        RECT 16.064 17.94 16.096 18.012 ;
  LAYER M2 ;
        RECT 16.044 17.96 16.116 17.992 ;
  LAYER M2 ;
        RECT 15.92 17.96 16.08 17.992 ;
  LAYER M1 ;
        RECT 15.904 17.94 15.936 18.012 ;
  LAYER M2 ;
        RECT 15.884 17.96 15.956 17.992 ;
  LAYER M1 ;
        RECT 16.064 14.832 16.096 14.904 ;
  LAYER M2 ;
        RECT 16.044 14.852 16.116 14.884 ;
  LAYER M1 ;
        RECT 16.064 14.868 16.096 15.036 ;
  LAYER M1 ;
        RECT 16.064 15 16.096 15.072 ;
  LAYER M2 ;
        RECT 16.044 15.02 16.116 15.052 ;
  LAYER M2 ;
        RECT 15.92 15.02 16.08 15.052 ;
  LAYER M1 ;
        RECT 15.904 15 15.936 15.072 ;
  LAYER M2 ;
        RECT 15.884 15.02 15.956 15.052 ;
  LAYER M1 ;
        RECT 16.064 11.892 16.096 11.964 ;
  LAYER M2 ;
        RECT 16.044 11.912 16.116 11.944 ;
  LAYER M1 ;
        RECT 16.064 11.928 16.096 12.096 ;
  LAYER M1 ;
        RECT 16.064 12.06 16.096 12.132 ;
  LAYER M2 ;
        RECT 16.044 12.08 16.116 12.112 ;
  LAYER M2 ;
        RECT 15.92 12.08 16.08 12.112 ;
  LAYER M1 ;
        RECT 15.904 12.06 15.936 12.132 ;
  LAYER M2 ;
        RECT 15.884 12.08 15.956 12.112 ;
  LAYER M1 ;
        RECT 16.064 8.952 16.096 9.024 ;
  LAYER M2 ;
        RECT 16.044 8.972 16.116 9.004 ;
  LAYER M1 ;
        RECT 16.064 8.988 16.096 9.156 ;
  LAYER M1 ;
        RECT 16.064 9.12 16.096 9.192 ;
  LAYER M2 ;
        RECT 16.044 9.14 16.116 9.172 ;
  LAYER M2 ;
        RECT 15.92 9.14 16.08 9.172 ;
  LAYER M1 ;
        RECT 15.904 9.12 15.936 9.192 ;
  LAYER M2 ;
        RECT 15.884 9.14 15.956 9.172 ;
  LAYER M1 ;
        RECT 15.904 18.612 15.936 18.684 ;
  LAYER M2 ;
        RECT 15.884 18.632 15.956 18.664 ;
  LAYER M1 ;
        RECT 15.904 18.144 15.936 18.648 ;
  LAYER M1 ;
        RECT 15.904 9.156 15.936 18.144 ;
  LAYER M2 ;
        RECT 15.92 18.632 30.32 18.664 ;
  LAYER M1 ;
        RECT 24.704 17.772 24.736 17.844 ;
  LAYER M2 ;
        RECT 24.684 17.792 24.756 17.824 ;
  LAYER M2 ;
        RECT 24.72 17.792 27.6 17.824 ;
  LAYER M1 ;
        RECT 27.584 17.772 27.616 17.844 ;
  LAYER M2 ;
        RECT 27.564 17.792 27.636 17.824 ;
  LAYER M1 ;
        RECT 24.704 8.952 24.736 9.024 ;
  LAYER M2 ;
        RECT 24.684 8.972 24.756 9.004 ;
  LAYER M2 ;
        RECT 24.72 8.972 27.6 9.004 ;
  LAYER M1 ;
        RECT 27.584 8.952 27.616 9.024 ;
  LAYER M2 ;
        RECT 27.564 8.972 27.636 9.004 ;
  LAYER M1 ;
        RECT 21.824 8.952 21.856 9.024 ;
  LAYER M2 ;
        RECT 21.804 8.972 21.876 9.004 ;
  LAYER M2 ;
        RECT 21.84 8.972 24.72 9.004 ;
  LAYER M1 ;
        RECT 24.704 8.952 24.736 9.024 ;
  LAYER M2 ;
        RECT 24.684 8.972 24.756 9.004 ;
  LAYER M1 ;
        RECT 18.944 8.952 18.976 9.024 ;
  LAYER M2 ;
        RECT 18.924 8.972 18.996 9.004 ;
  LAYER M2 ;
        RECT 18.96 8.972 21.84 9.004 ;
  LAYER M1 ;
        RECT 21.824 8.952 21.856 9.024 ;
  LAYER M2 ;
        RECT 21.804 8.972 21.876 9.004 ;
  LAYER M1 ;
        RECT 18.944 17.772 18.976 17.844 ;
  LAYER M2 ;
        RECT 18.924 17.792 18.996 17.824 ;
  LAYER M2 ;
        RECT 16.08 17.792 18.96 17.824 ;
  LAYER M1 ;
        RECT 16.064 17.772 16.096 17.844 ;
  LAYER M2 ;
        RECT 16.044 17.792 16.116 17.824 ;
  LAYER M1 ;
        RECT 21.824 17.772 21.856 17.844 ;
  LAYER M2 ;
        RECT 21.804 17.792 21.876 17.824 ;
  LAYER M2 ;
        RECT 18.96 17.792 21.84 17.824 ;
  LAYER M1 ;
        RECT 18.944 17.772 18.976 17.844 ;
  LAYER M2 ;
        RECT 18.924 17.792 18.996 17.824 ;
  LAYER M1 ;
        RECT 24.224 9.456 24.256 9.528 ;
  LAYER M2 ;
        RECT 24.204 9.476 24.276 9.508 ;
  LAYER M2 ;
        RECT 24.24 9.476 24.4 9.508 ;
  LAYER M1 ;
        RECT 24.384 9.456 24.416 9.528 ;
  LAYER M2 ;
        RECT 24.364 9.476 24.436 9.508 ;
  LAYER M1 ;
        RECT 27.104 12.396 27.136 12.468 ;
  LAYER M2 ;
        RECT 27.084 12.416 27.156 12.448 ;
  LAYER M1 ;
        RECT 27.104 12.264 27.136 12.432 ;
  LAYER M1 ;
        RECT 27.104 12.228 27.136 12.3 ;
  LAYER M2 ;
        RECT 27.084 12.248 27.156 12.28 ;
  LAYER M2 ;
        RECT 24.4 12.248 27.12 12.28 ;
  LAYER M1 ;
        RECT 24.384 12.228 24.416 12.3 ;
  LAYER M2 ;
        RECT 24.364 12.248 24.436 12.28 ;
  LAYER M1 ;
        RECT 24.384 6.012 24.416 6.084 ;
  LAYER M2 ;
        RECT 24.364 6.032 24.436 6.064 ;
  LAYER M1 ;
        RECT 24.384 6.048 24.416 6.216 ;
  LAYER M1 ;
        RECT 24.384 6.216 24.416 12.264 ;
  LAYER M1 ;
        RECT 21.344 9.456 21.376 9.528 ;
  LAYER M2 ;
        RECT 21.324 9.476 21.396 9.508 ;
  LAYER M2 ;
        RECT 21.36 9.476 21.52 9.508 ;
  LAYER M1 ;
        RECT 21.504 9.456 21.536 9.528 ;
  LAYER M2 ;
        RECT 21.484 9.476 21.556 9.508 ;
  LAYER M1 ;
        RECT 21.504 6.012 21.536 6.084 ;
  LAYER M2 ;
        RECT 21.484 6.032 21.556 6.064 ;
  LAYER M1 ;
        RECT 21.504 6.048 21.536 6.216 ;
  LAYER M1 ;
        RECT 21.504 6.216 21.536 9.492 ;
  LAYER M2 ;
        RECT 21.52 6.032 24.4 6.064 ;
  LAYER M1 ;
        RECT 27.104 9.456 27.136 9.528 ;
  LAYER M2 ;
        RECT 27.084 9.476 27.156 9.508 ;
  LAYER M2 ;
        RECT 27.12 9.476 27.28 9.508 ;
  LAYER M1 ;
        RECT 27.264 9.456 27.296 9.528 ;
  LAYER M2 ;
        RECT 27.244 9.476 27.316 9.508 ;
  LAYER M1 ;
        RECT 27.264 5.844 27.296 5.916 ;
  LAYER M2 ;
        RECT 27.244 5.864 27.316 5.896 ;
  LAYER M1 ;
        RECT 27.264 5.88 27.296 6.216 ;
  LAYER M1 ;
        RECT 27.264 6.216 27.296 9.492 ;
  LAYER M1 ;
        RECT 21.344 12.396 21.376 12.468 ;
  LAYER M2 ;
        RECT 21.324 12.416 21.396 12.448 ;
  LAYER M1 ;
        RECT 21.344 12.264 21.376 12.432 ;
  LAYER M1 ;
        RECT 21.344 12.228 21.376 12.3 ;
  LAYER M2 ;
        RECT 21.324 12.248 21.396 12.28 ;
  LAYER M2 ;
        RECT 18.64 12.248 21.36 12.28 ;
  LAYER M1 ;
        RECT 18.624 12.228 18.656 12.3 ;
  LAYER M2 ;
        RECT 18.604 12.248 18.676 12.28 ;
  LAYER M1 ;
        RECT 18.624 5.844 18.656 5.916 ;
  LAYER M2 ;
        RECT 18.604 5.864 18.676 5.896 ;
  LAYER M1 ;
        RECT 18.624 5.88 18.656 6.216 ;
  LAYER M1 ;
        RECT 18.624 6.216 18.656 12.264 ;
  LAYER M2 ;
        RECT 18.64 5.864 27.28 5.896 ;
  LAYER M1 ;
        RECT 24.224 12.396 24.256 12.468 ;
  LAYER M2 ;
        RECT 24.204 12.416 24.276 12.448 ;
  LAYER M2 ;
        RECT 21.36 12.416 24.24 12.448 ;
  LAYER M1 ;
        RECT 21.344 12.396 21.376 12.468 ;
  LAYER M2 ;
        RECT 21.324 12.416 21.396 12.448 ;
  LAYER M1 ;
        RECT 29.984 15.336 30.016 15.408 ;
  LAYER M2 ;
        RECT 29.964 15.356 30.036 15.388 ;
  LAYER M2 ;
        RECT 30 15.356 30.16 15.388 ;
  LAYER M1 ;
        RECT 30.144 15.336 30.176 15.408 ;
  LAYER M2 ;
        RECT 30.124 15.356 30.196 15.388 ;
  LAYER M1 ;
        RECT 29.984 12.396 30.016 12.468 ;
  LAYER M2 ;
        RECT 29.964 12.416 30.036 12.448 ;
  LAYER M2 ;
        RECT 30 12.416 30.16 12.448 ;
  LAYER M1 ;
        RECT 30.144 12.396 30.176 12.468 ;
  LAYER M2 ;
        RECT 30.124 12.416 30.196 12.448 ;
  LAYER M1 ;
        RECT 29.984 9.456 30.016 9.528 ;
  LAYER M2 ;
        RECT 29.964 9.476 30.036 9.508 ;
  LAYER M2 ;
        RECT 30 9.476 30.16 9.508 ;
  LAYER M1 ;
        RECT 30.144 9.456 30.176 9.528 ;
  LAYER M2 ;
        RECT 30.124 9.476 30.196 9.508 ;
  LAYER M1 ;
        RECT 29.984 6.516 30.016 6.588 ;
  LAYER M2 ;
        RECT 29.964 6.536 30.036 6.568 ;
  LAYER M2 ;
        RECT 30 6.536 30.16 6.568 ;
  LAYER M1 ;
        RECT 30.144 6.516 30.176 6.588 ;
  LAYER M2 ;
        RECT 30.124 6.536 30.196 6.568 ;
  LAYER M1 ;
        RECT 30.144 5.676 30.176 5.748 ;
  LAYER M2 ;
        RECT 30.124 5.696 30.196 5.728 ;
  LAYER M1 ;
        RECT 30.144 5.712 30.176 6.216 ;
  LAYER M1 ;
        RECT 30.144 6.216 30.176 15.372 ;
  LAYER M1 ;
        RECT 18.464 15.336 18.496 15.408 ;
  LAYER M2 ;
        RECT 18.444 15.356 18.516 15.388 ;
  LAYER M1 ;
        RECT 18.464 15.204 18.496 15.372 ;
  LAYER M1 ;
        RECT 18.464 15.168 18.496 15.24 ;
  LAYER M2 ;
        RECT 18.444 15.188 18.516 15.22 ;
  LAYER M2 ;
        RECT 15.76 15.188 18.48 15.22 ;
  LAYER M1 ;
        RECT 15.744 15.168 15.776 15.24 ;
  LAYER M2 ;
        RECT 15.724 15.188 15.796 15.22 ;
  LAYER M1 ;
        RECT 18.464 12.396 18.496 12.468 ;
  LAYER M2 ;
        RECT 18.444 12.416 18.516 12.448 ;
  LAYER M1 ;
        RECT 18.464 12.264 18.496 12.432 ;
  LAYER M1 ;
        RECT 18.464 12.228 18.496 12.3 ;
  LAYER M2 ;
        RECT 18.444 12.248 18.516 12.28 ;
  LAYER M2 ;
        RECT 15.76 12.248 18.48 12.28 ;
  LAYER M1 ;
        RECT 15.744 12.228 15.776 12.3 ;
  LAYER M2 ;
        RECT 15.724 12.248 15.796 12.28 ;
  LAYER M1 ;
        RECT 18.464 9.456 18.496 9.528 ;
  LAYER M2 ;
        RECT 18.444 9.476 18.516 9.508 ;
  LAYER M1 ;
        RECT 18.464 9.324 18.496 9.492 ;
  LAYER M1 ;
        RECT 18.464 9.288 18.496 9.36 ;
  LAYER M2 ;
        RECT 18.444 9.308 18.516 9.34 ;
  LAYER M2 ;
        RECT 15.76 9.308 18.48 9.34 ;
  LAYER M1 ;
        RECT 15.744 9.288 15.776 9.36 ;
  LAYER M2 ;
        RECT 15.724 9.308 15.796 9.34 ;
  LAYER M1 ;
        RECT 18.464 6.516 18.496 6.588 ;
  LAYER M2 ;
        RECT 18.444 6.536 18.516 6.568 ;
  LAYER M1 ;
        RECT 18.464 6.384 18.496 6.552 ;
  LAYER M1 ;
        RECT 18.464 6.348 18.496 6.42 ;
  LAYER M2 ;
        RECT 18.444 6.368 18.516 6.4 ;
  LAYER M2 ;
        RECT 15.76 6.368 18.48 6.4 ;
  LAYER M1 ;
        RECT 15.744 6.348 15.776 6.42 ;
  LAYER M2 ;
        RECT 15.724 6.368 15.796 6.4 ;
  LAYER M1 ;
        RECT 15.744 5.676 15.776 5.748 ;
  LAYER M2 ;
        RECT 15.724 5.696 15.796 5.728 ;
  LAYER M1 ;
        RECT 15.744 5.712 15.776 6.216 ;
  LAYER M1 ;
        RECT 15.744 6.216 15.776 15.204 ;
  LAYER M2 ;
        RECT 15.76 5.696 30.16 5.728 ;
  LAYER M1 ;
        RECT 27.104 15.336 27.136 15.408 ;
  LAYER M2 ;
        RECT 27.084 15.356 27.156 15.388 ;
  LAYER M2 ;
        RECT 27.12 15.356 30 15.388 ;
  LAYER M1 ;
        RECT 29.984 15.336 30.016 15.408 ;
  LAYER M2 ;
        RECT 29.964 15.356 30.036 15.388 ;
  LAYER M1 ;
        RECT 27.104 6.516 27.136 6.588 ;
  LAYER M2 ;
        RECT 27.084 6.536 27.156 6.568 ;
  LAYER M2 ;
        RECT 27.12 6.536 30 6.568 ;
  LAYER M1 ;
        RECT 29.984 6.516 30.016 6.588 ;
  LAYER M2 ;
        RECT 29.964 6.536 30.036 6.568 ;
  LAYER M1 ;
        RECT 24.224 6.516 24.256 6.588 ;
  LAYER M2 ;
        RECT 24.204 6.536 24.276 6.568 ;
  LAYER M2 ;
        RECT 24.24 6.536 27.12 6.568 ;
  LAYER M1 ;
        RECT 27.104 6.516 27.136 6.588 ;
  LAYER M2 ;
        RECT 27.084 6.536 27.156 6.568 ;
  LAYER M1 ;
        RECT 21.344 6.516 21.376 6.588 ;
  LAYER M2 ;
        RECT 21.324 6.536 21.396 6.568 ;
  LAYER M2 ;
        RECT 21.36 6.536 24.24 6.568 ;
  LAYER M1 ;
        RECT 24.224 6.516 24.256 6.588 ;
  LAYER M2 ;
        RECT 24.204 6.536 24.276 6.568 ;
  LAYER M1 ;
        RECT 21.344 15.336 21.376 15.408 ;
  LAYER M2 ;
        RECT 21.324 15.356 21.396 15.388 ;
  LAYER M2 ;
        RECT 18.48 15.356 21.36 15.388 ;
  LAYER M1 ;
        RECT 18.464 15.336 18.496 15.408 ;
  LAYER M2 ;
        RECT 18.444 15.356 18.516 15.388 ;
  LAYER M1 ;
        RECT 24.224 15.336 24.256 15.408 ;
  LAYER M2 ;
        RECT 24.204 15.356 24.276 15.388 ;
  LAYER M2 ;
        RECT 21.36 15.356 24.24 15.388 ;
  LAYER M1 ;
        RECT 21.344 15.336 21.376 15.408 ;
  LAYER M2 ;
        RECT 21.324 15.356 21.396 15.388 ;
  LAYER M1 ;
        RECT 27.6 15.372 30 17.808 ;
  LAYER M2 ;
        RECT 27.6 15.372 30 17.808 ;
  LAYER M3 ;
        RECT 27.6 15.372 30 17.808 ;
  LAYER M1 ;
        RECT 27.6 12.432 30 14.868 ;
  LAYER M2 ;
        RECT 27.6 12.432 30 14.868 ;
  LAYER M3 ;
        RECT 27.6 12.432 30 14.868 ;
  LAYER M1 ;
        RECT 27.6 9.492 30 11.928 ;
  LAYER M2 ;
        RECT 27.6 9.492 30 11.928 ;
  LAYER M3 ;
        RECT 27.6 9.492 30 11.928 ;
  LAYER M1 ;
        RECT 27.6 6.552 30 8.988 ;
  LAYER M2 ;
        RECT 27.6 6.552 30 8.988 ;
  LAYER M3 ;
        RECT 27.6 6.552 30 8.988 ;
  LAYER M1 ;
        RECT 24.72 15.372 27.12 17.808 ;
  LAYER M2 ;
        RECT 24.72 15.372 27.12 17.808 ;
  LAYER M3 ;
        RECT 24.72 15.372 27.12 17.808 ;
  LAYER M1 ;
        RECT 24.72 12.432 27.12 14.868 ;
  LAYER M2 ;
        RECT 24.72 12.432 27.12 14.868 ;
  LAYER M3 ;
        RECT 24.72 12.432 27.12 14.868 ;
  LAYER M1 ;
        RECT 24.72 9.492 27.12 11.928 ;
  LAYER M2 ;
        RECT 24.72 9.492 27.12 11.928 ;
  LAYER M3 ;
        RECT 24.72 9.492 27.12 11.928 ;
  LAYER M1 ;
        RECT 24.72 6.552 27.12 8.988 ;
  LAYER M2 ;
        RECT 24.72 6.552 27.12 8.988 ;
  LAYER M3 ;
        RECT 24.72 6.552 27.12 8.988 ;
  LAYER M1 ;
        RECT 21.84 15.372 24.24 17.808 ;
  LAYER M2 ;
        RECT 21.84 15.372 24.24 17.808 ;
  LAYER M3 ;
        RECT 21.84 15.372 24.24 17.808 ;
  LAYER M1 ;
        RECT 21.84 12.432 24.24 14.868 ;
  LAYER M2 ;
        RECT 21.84 12.432 24.24 14.868 ;
  LAYER M3 ;
        RECT 21.84 12.432 24.24 14.868 ;
  LAYER M1 ;
        RECT 21.84 9.492 24.24 11.928 ;
  LAYER M2 ;
        RECT 21.84 9.492 24.24 11.928 ;
  LAYER M3 ;
        RECT 21.84 9.492 24.24 11.928 ;
  LAYER M1 ;
        RECT 21.84 6.552 24.24 8.988 ;
  LAYER M2 ;
        RECT 21.84 6.552 24.24 8.988 ;
  LAYER M3 ;
        RECT 21.84 6.552 24.24 8.988 ;
  LAYER M1 ;
        RECT 18.96 15.372 21.36 17.808 ;
  LAYER M2 ;
        RECT 18.96 15.372 21.36 17.808 ;
  LAYER M3 ;
        RECT 18.96 15.372 21.36 17.808 ;
  LAYER M1 ;
        RECT 18.96 12.432 21.36 14.868 ;
  LAYER M2 ;
        RECT 18.96 12.432 21.36 14.868 ;
  LAYER M3 ;
        RECT 18.96 12.432 21.36 14.868 ;
  LAYER M1 ;
        RECT 18.96 9.492 21.36 11.928 ;
  LAYER M2 ;
        RECT 18.96 9.492 21.36 11.928 ;
  LAYER M3 ;
        RECT 18.96 9.492 21.36 11.928 ;
  LAYER M1 ;
        RECT 18.96 6.552 21.36 8.988 ;
  LAYER M2 ;
        RECT 18.96 6.552 21.36 8.988 ;
  LAYER M3 ;
        RECT 18.96 6.552 21.36 8.988 ;
  LAYER M1 ;
        RECT 16.08 15.372 18.48 17.808 ;
  LAYER M2 ;
        RECT 16.08 15.372 18.48 17.808 ;
  LAYER M3 ;
        RECT 16.08 15.372 18.48 17.808 ;
  LAYER M1 ;
        RECT 16.08 12.432 18.48 14.868 ;
  LAYER M2 ;
        RECT 16.08 12.432 18.48 14.868 ;
  LAYER M3 ;
        RECT 16.08 12.432 18.48 14.868 ;
  LAYER M1 ;
        RECT 16.08 9.492 18.48 11.928 ;
  LAYER M2 ;
        RECT 16.08 9.492 18.48 11.928 ;
  LAYER M3 ;
        RECT 16.08 9.492 18.48 11.928 ;
  LAYER M1 ;
        RECT 16.08 6.552 18.48 8.988 ;
  LAYER M2 ;
        RECT 16.08 6.552 18.48 8.988 ;
  LAYER M3 ;
        RECT 16.08 6.552 18.48 8.988 ;
  LAYER M1 ;
        RECT 24.224 30.96 24.256 31.032 ;
  LAYER M2 ;
        RECT 24.204 30.98 24.276 31.012 ;
  LAYER M2 ;
        RECT 21.52 30.98 24.24 31.012 ;
  LAYER M1 ;
        RECT 21.504 30.96 21.536 31.032 ;
  LAYER M2 ;
        RECT 21.484 30.98 21.556 31.012 ;
  LAYER M1 ;
        RECT 24.224 28.02 24.256 28.092 ;
  LAYER M2 ;
        RECT 24.204 28.04 24.276 28.072 ;
  LAYER M2 ;
        RECT 21.52 28.04 24.24 28.072 ;
  LAYER M1 ;
        RECT 21.504 28.02 21.536 28.092 ;
  LAYER M2 ;
        RECT 21.484 28.04 21.556 28.072 ;
  LAYER M1 ;
        RECT 21.344 30.96 21.376 31.032 ;
  LAYER M2 ;
        RECT 21.324 30.98 21.396 31.012 ;
  LAYER M1 ;
        RECT 21.344 30.996 21.376 31.164 ;
  LAYER M1 ;
        RECT 21.344 31.128 21.376 31.2 ;
  LAYER M2 ;
        RECT 21.324 31.148 21.396 31.18 ;
  LAYER M2 ;
        RECT 21.36 31.148 21.52 31.18 ;
  LAYER M1 ;
        RECT 21.504 31.128 21.536 31.2 ;
  LAYER M2 ;
        RECT 21.484 31.148 21.556 31.18 ;
  LAYER M1 ;
        RECT 21.344 28.02 21.376 28.092 ;
  LAYER M2 ;
        RECT 21.324 28.04 21.396 28.072 ;
  LAYER M1 ;
        RECT 21.344 28.056 21.376 28.224 ;
  LAYER M1 ;
        RECT 21.344 28.188 21.376 28.26 ;
  LAYER M2 ;
        RECT 21.324 28.208 21.396 28.24 ;
  LAYER M2 ;
        RECT 21.36 28.208 21.52 28.24 ;
  LAYER M1 ;
        RECT 21.504 28.188 21.536 28.26 ;
  LAYER M2 ;
        RECT 21.484 28.208 21.556 28.24 ;
  LAYER M1 ;
        RECT 21.504 37.344 21.536 37.416 ;
  LAYER M2 ;
        RECT 21.484 37.364 21.556 37.396 ;
  LAYER M1 ;
        RECT 21.504 37.212 21.536 37.38 ;
  LAYER M1 ;
        RECT 21.504 28.056 21.536 37.212 ;
  LAYER M1 ;
        RECT 27.104 28.02 27.136 28.092 ;
  LAYER M2 ;
        RECT 27.084 28.04 27.156 28.072 ;
  LAYER M2 ;
        RECT 24.4 28.04 27.12 28.072 ;
  LAYER M1 ;
        RECT 24.384 28.02 24.416 28.092 ;
  LAYER M2 ;
        RECT 24.364 28.04 24.436 28.072 ;
  LAYER M1 ;
        RECT 27.104 30.96 27.136 31.032 ;
  LAYER M2 ;
        RECT 27.084 30.98 27.156 31.012 ;
  LAYER M2 ;
        RECT 24.4 30.98 27.12 31.012 ;
  LAYER M1 ;
        RECT 24.384 30.96 24.416 31.032 ;
  LAYER M2 ;
        RECT 24.364 30.98 24.436 31.012 ;
  LAYER M1 ;
        RECT 24.384 37.344 24.416 37.416 ;
  LAYER M2 ;
        RECT 24.364 37.364 24.436 37.396 ;
  LAYER M1 ;
        RECT 24.384 37.212 24.416 37.38 ;
  LAYER M1 ;
        RECT 24.384 28.056 24.416 37.212 ;
  LAYER M2 ;
        RECT 21.52 37.364 24.4 37.396 ;
  LAYER M1 ;
        RECT 21.344 25.08 21.376 25.152 ;
  LAYER M2 ;
        RECT 21.324 25.1 21.396 25.132 ;
  LAYER M2 ;
        RECT 18.64 25.1 21.36 25.132 ;
  LAYER M1 ;
        RECT 18.624 25.08 18.656 25.152 ;
  LAYER M2 ;
        RECT 18.604 25.1 18.676 25.132 ;
  LAYER M1 ;
        RECT 21.344 33.9 21.376 33.972 ;
  LAYER M2 ;
        RECT 21.324 33.92 21.396 33.952 ;
  LAYER M2 ;
        RECT 18.64 33.92 21.36 33.952 ;
  LAYER M1 ;
        RECT 18.624 33.9 18.656 33.972 ;
  LAYER M2 ;
        RECT 18.604 33.92 18.676 33.952 ;
  LAYER M1 ;
        RECT 18.624 37.512 18.656 37.584 ;
  LAYER M2 ;
        RECT 18.604 37.532 18.676 37.564 ;
  LAYER M1 ;
        RECT 18.624 37.212 18.656 37.548 ;
  LAYER M1 ;
        RECT 18.624 25.116 18.656 37.212 ;
  LAYER M1 ;
        RECT 27.104 33.9 27.136 33.972 ;
  LAYER M2 ;
        RECT 27.084 33.92 27.156 33.952 ;
  LAYER M1 ;
        RECT 27.104 33.936 27.136 34.104 ;
  LAYER M1 ;
        RECT 27.104 34.068 27.136 34.14 ;
  LAYER M2 ;
        RECT 27.084 34.088 27.156 34.12 ;
  LAYER M2 ;
        RECT 27.12 34.088 27.28 34.12 ;
  LAYER M1 ;
        RECT 27.264 34.068 27.296 34.14 ;
  LAYER M2 ;
        RECT 27.244 34.088 27.316 34.12 ;
  LAYER M1 ;
        RECT 27.104 25.08 27.136 25.152 ;
  LAYER M2 ;
        RECT 27.084 25.1 27.156 25.132 ;
  LAYER M1 ;
        RECT 27.104 25.116 27.136 25.284 ;
  LAYER M1 ;
        RECT 27.104 25.248 27.136 25.32 ;
  LAYER M2 ;
        RECT 27.084 25.268 27.156 25.3 ;
  LAYER M2 ;
        RECT 27.12 25.268 27.28 25.3 ;
  LAYER M1 ;
        RECT 27.264 25.248 27.296 25.32 ;
  LAYER M2 ;
        RECT 27.244 25.268 27.316 25.3 ;
  LAYER M1 ;
        RECT 27.264 37.512 27.296 37.584 ;
  LAYER M2 ;
        RECT 27.244 37.532 27.316 37.564 ;
  LAYER M1 ;
        RECT 27.264 37.212 27.296 37.548 ;
  LAYER M1 ;
        RECT 27.264 25.284 27.296 37.212 ;
  LAYER M2 ;
        RECT 18.64 37.532 27.28 37.564 ;
  LAYER M1 ;
        RECT 24.224 33.9 24.256 33.972 ;
  LAYER M2 ;
        RECT 24.204 33.92 24.276 33.952 ;
  LAYER M2 ;
        RECT 24.24 33.92 27.12 33.952 ;
  LAYER M1 ;
        RECT 27.104 33.9 27.136 33.972 ;
  LAYER M2 ;
        RECT 27.084 33.92 27.156 33.952 ;
  LAYER M1 ;
        RECT 24.224 25.08 24.256 25.152 ;
  LAYER M2 ;
        RECT 24.204 25.1 24.276 25.132 ;
  LAYER M2 ;
        RECT 21.36 25.1 24.24 25.132 ;
  LAYER M1 ;
        RECT 21.344 25.08 21.376 25.152 ;
  LAYER M2 ;
        RECT 21.324 25.1 21.396 25.132 ;
  LAYER M1 ;
        RECT 18.464 36.84 18.496 36.912 ;
  LAYER M2 ;
        RECT 18.444 36.86 18.516 36.892 ;
  LAYER M2 ;
        RECT 15.76 36.86 18.48 36.892 ;
  LAYER M1 ;
        RECT 15.744 36.84 15.776 36.912 ;
  LAYER M2 ;
        RECT 15.724 36.86 15.796 36.892 ;
  LAYER M1 ;
        RECT 18.464 33.9 18.496 33.972 ;
  LAYER M2 ;
        RECT 18.444 33.92 18.516 33.952 ;
  LAYER M2 ;
        RECT 15.76 33.92 18.48 33.952 ;
  LAYER M1 ;
        RECT 15.744 33.9 15.776 33.972 ;
  LAYER M2 ;
        RECT 15.724 33.92 15.796 33.952 ;
  LAYER M1 ;
        RECT 18.464 30.96 18.496 31.032 ;
  LAYER M2 ;
        RECT 18.444 30.98 18.516 31.012 ;
  LAYER M2 ;
        RECT 15.76 30.98 18.48 31.012 ;
  LAYER M1 ;
        RECT 15.744 30.96 15.776 31.032 ;
  LAYER M2 ;
        RECT 15.724 30.98 15.796 31.012 ;
  LAYER M1 ;
        RECT 18.464 28.02 18.496 28.092 ;
  LAYER M2 ;
        RECT 18.444 28.04 18.516 28.072 ;
  LAYER M2 ;
        RECT 15.76 28.04 18.48 28.072 ;
  LAYER M1 ;
        RECT 15.744 28.02 15.776 28.092 ;
  LAYER M2 ;
        RECT 15.724 28.04 15.796 28.072 ;
  LAYER M1 ;
        RECT 18.464 25.08 18.496 25.152 ;
  LAYER M2 ;
        RECT 18.444 25.1 18.516 25.132 ;
  LAYER M2 ;
        RECT 15.76 25.1 18.48 25.132 ;
  LAYER M1 ;
        RECT 15.744 25.08 15.776 25.152 ;
  LAYER M2 ;
        RECT 15.724 25.1 15.796 25.132 ;
  LAYER M1 ;
        RECT 18.464 22.14 18.496 22.212 ;
  LAYER M2 ;
        RECT 18.444 22.16 18.516 22.192 ;
  LAYER M2 ;
        RECT 15.76 22.16 18.48 22.192 ;
  LAYER M1 ;
        RECT 15.744 22.14 15.776 22.212 ;
  LAYER M2 ;
        RECT 15.724 22.16 15.796 22.192 ;
  LAYER M1 ;
        RECT 15.744 37.68 15.776 37.752 ;
  LAYER M2 ;
        RECT 15.724 37.7 15.796 37.732 ;
  LAYER M1 ;
        RECT 15.744 37.212 15.776 37.716 ;
  LAYER M1 ;
        RECT 15.744 22.176 15.776 37.212 ;
  LAYER M1 ;
        RECT 29.984 36.84 30.016 36.912 ;
  LAYER M2 ;
        RECT 29.964 36.86 30.036 36.892 ;
  LAYER M1 ;
        RECT 29.984 36.876 30.016 37.044 ;
  LAYER M1 ;
        RECT 29.984 37.008 30.016 37.08 ;
  LAYER M2 ;
        RECT 29.964 37.028 30.036 37.06 ;
  LAYER M2 ;
        RECT 30 37.028 30.16 37.06 ;
  LAYER M1 ;
        RECT 30.144 37.008 30.176 37.08 ;
  LAYER M2 ;
        RECT 30.124 37.028 30.196 37.06 ;
  LAYER M1 ;
        RECT 29.984 33.9 30.016 33.972 ;
  LAYER M2 ;
        RECT 29.964 33.92 30.036 33.952 ;
  LAYER M1 ;
        RECT 29.984 33.936 30.016 34.104 ;
  LAYER M1 ;
        RECT 29.984 34.068 30.016 34.14 ;
  LAYER M2 ;
        RECT 29.964 34.088 30.036 34.12 ;
  LAYER M2 ;
        RECT 30 34.088 30.16 34.12 ;
  LAYER M1 ;
        RECT 30.144 34.068 30.176 34.14 ;
  LAYER M2 ;
        RECT 30.124 34.088 30.196 34.12 ;
  LAYER M1 ;
        RECT 29.984 30.96 30.016 31.032 ;
  LAYER M2 ;
        RECT 29.964 30.98 30.036 31.012 ;
  LAYER M1 ;
        RECT 29.984 30.996 30.016 31.164 ;
  LAYER M1 ;
        RECT 29.984 31.128 30.016 31.2 ;
  LAYER M2 ;
        RECT 29.964 31.148 30.036 31.18 ;
  LAYER M2 ;
        RECT 30 31.148 30.16 31.18 ;
  LAYER M1 ;
        RECT 30.144 31.128 30.176 31.2 ;
  LAYER M2 ;
        RECT 30.124 31.148 30.196 31.18 ;
  LAYER M1 ;
        RECT 29.984 28.02 30.016 28.092 ;
  LAYER M2 ;
        RECT 29.964 28.04 30.036 28.072 ;
  LAYER M1 ;
        RECT 29.984 28.056 30.016 28.224 ;
  LAYER M1 ;
        RECT 29.984 28.188 30.016 28.26 ;
  LAYER M2 ;
        RECT 29.964 28.208 30.036 28.24 ;
  LAYER M2 ;
        RECT 30 28.208 30.16 28.24 ;
  LAYER M1 ;
        RECT 30.144 28.188 30.176 28.26 ;
  LAYER M2 ;
        RECT 30.124 28.208 30.196 28.24 ;
  LAYER M1 ;
        RECT 29.984 25.08 30.016 25.152 ;
  LAYER M2 ;
        RECT 29.964 25.1 30.036 25.132 ;
  LAYER M1 ;
        RECT 29.984 25.116 30.016 25.284 ;
  LAYER M1 ;
        RECT 29.984 25.248 30.016 25.32 ;
  LAYER M2 ;
        RECT 29.964 25.268 30.036 25.3 ;
  LAYER M2 ;
        RECT 30 25.268 30.16 25.3 ;
  LAYER M1 ;
        RECT 30.144 25.248 30.176 25.32 ;
  LAYER M2 ;
        RECT 30.124 25.268 30.196 25.3 ;
  LAYER M1 ;
        RECT 29.984 22.14 30.016 22.212 ;
  LAYER M2 ;
        RECT 29.964 22.16 30.036 22.192 ;
  LAYER M1 ;
        RECT 29.984 22.176 30.016 22.344 ;
  LAYER M1 ;
        RECT 29.984 22.308 30.016 22.38 ;
  LAYER M2 ;
        RECT 29.964 22.328 30.036 22.36 ;
  LAYER M2 ;
        RECT 30 22.328 30.16 22.36 ;
  LAYER M1 ;
        RECT 30.144 22.308 30.176 22.38 ;
  LAYER M2 ;
        RECT 30.124 22.328 30.196 22.36 ;
  LAYER M1 ;
        RECT 30.144 37.68 30.176 37.752 ;
  LAYER M2 ;
        RECT 30.124 37.7 30.196 37.732 ;
  LAYER M1 ;
        RECT 30.144 37.212 30.176 37.716 ;
  LAYER M1 ;
        RECT 30.144 22.344 30.176 37.212 ;
  LAYER M2 ;
        RECT 15.76 37.7 30.16 37.732 ;
  LAYER M1 ;
        RECT 21.344 36.84 21.376 36.912 ;
  LAYER M2 ;
        RECT 21.324 36.86 21.396 36.892 ;
  LAYER M2 ;
        RECT 18.48 36.86 21.36 36.892 ;
  LAYER M1 ;
        RECT 18.464 36.84 18.496 36.912 ;
  LAYER M2 ;
        RECT 18.444 36.86 18.516 36.892 ;
  LAYER M1 ;
        RECT 21.344 22.14 21.376 22.212 ;
  LAYER M2 ;
        RECT 21.324 22.16 21.396 22.192 ;
  LAYER M2 ;
        RECT 18.48 22.16 21.36 22.192 ;
  LAYER M1 ;
        RECT 18.464 22.14 18.496 22.212 ;
  LAYER M2 ;
        RECT 18.444 22.16 18.516 22.192 ;
  LAYER M1 ;
        RECT 24.224 22.14 24.256 22.212 ;
  LAYER M2 ;
        RECT 24.204 22.16 24.276 22.192 ;
  LAYER M2 ;
        RECT 21.36 22.16 24.24 22.192 ;
  LAYER M1 ;
        RECT 21.344 22.14 21.376 22.212 ;
  LAYER M2 ;
        RECT 21.324 22.16 21.396 22.192 ;
  LAYER M1 ;
        RECT 27.104 22.14 27.136 22.212 ;
  LAYER M2 ;
        RECT 27.084 22.16 27.156 22.192 ;
  LAYER M2 ;
        RECT 24.24 22.16 27.12 22.192 ;
  LAYER M1 ;
        RECT 24.224 22.14 24.256 22.212 ;
  LAYER M2 ;
        RECT 24.204 22.16 24.276 22.192 ;
  LAYER M1 ;
        RECT 27.104 36.84 27.136 36.912 ;
  LAYER M2 ;
        RECT 27.084 36.86 27.156 36.892 ;
  LAYER M2 ;
        RECT 27.12 36.86 30 36.892 ;
  LAYER M1 ;
        RECT 29.984 36.84 30.016 36.912 ;
  LAYER M2 ;
        RECT 29.964 36.86 30.036 36.892 ;
  LAYER M1 ;
        RECT 24.224 36.84 24.256 36.912 ;
  LAYER M2 ;
        RECT 24.204 36.86 24.276 36.892 ;
  LAYER M2 ;
        RECT 24.24 36.86 27.12 36.892 ;
  LAYER M1 ;
        RECT 27.104 36.84 27.136 36.912 ;
  LAYER M2 ;
        RECT 27.084 36.86 27.156 36.892 ;
  LAYER M1 ;
        RECT 21.824 28.524 21.856 28.596 ;
  LAYER M2 ;
        RECT 21.804 28.544 21.876 28.576 ;
  LAYER M2 ;
        RECT 21.68 28.544 21.84 28.576 ;
  LAYER M1 ;
        RECT 21.664 28.524 21.696 28.596 ;
  LAYER M2 ;
        RECT 21.644 28.544 21.716 28.576 ;
  LAYER M1 ;
        RECT 21.824 25.584 21.856 25.656 ;
  LAYER M2 ;
        RECT 21.804 25.604 21.876 25.636 ;
  LAYER M2 ;
        RECT 21.68 25.604 21.84 25.636 ;
  LAYER M1 ;
        RECT 21.664 25.584 21.696 25.656 ;
  LAYER M2 ;
        RECT 21.644 25.604 21.716 25.636 ;
  LAYER M1 ;
        RECT 18.944 28.524 18.976 28.596 ;
  LAYER M2 ;
        RECT 18.924 28.544 18.996 28.576 ;
  LAYER M1 ;
        RECT 18.944 28.392 18.976 28.56 ;
  LAYER M1 ;
        RECT 18.944 28.356 18.976 28.428 ;
  LAYER M2 ;
        RECT 18.924 28.376 18.996 28.408 ;
  LAYER M2 ;
        RECT 18.96 28.376 21.68 28.408 ;
  LAYER M1 ;
        RECT 21.664 28.356 21.696 28.428 ;
  LAYER M2 ;
        RECT 21.644 28.376 21.716 28.408 ;
  LAYER M1 ;
        RECT 18.944 25.584 18.976 25.656 ;
  LAYER M2 ;
        RECT 18.924 25.604 18.996 25.636 ;
  LAYER M1 ;
        RECT 18.944 25.452 18.976 25.62 ;
  LAYER M1 ;
        RECT 18.944 25.416 18.976 25.488 ;
  LAYER M2 ;
        RECT 18.924 25.436 18.996 25.468 ;
  LAYER M2 ;
        RECT 18.96 25.436 21.68 25.468 ;
  LAYER M1 ;
        RECT 21.664 25.416 21.696 25.488 ;
  LAYER M2 ;
        RECT 21.644 25.436 21.716 25.468 ;
  LAYER M1 ;
        RECT 21.664 19.2 21.696 19.272 ;
  LAYER M2 ;
        RECT 21.644 19.22 21.716 19.252 ;
  LAYER M1 ;
        RECT 21.664 19.236 21.696 19.404 ;
  LAYER M1 ;
        RECT 21.664 19.404 21.696 28.56 ;
  LAYER M1 ;
        RECT 24.704 25.584 24.736 25.656 ;
  LAYER M2 ;
        RECT 24.684 25.604 24.756 25.636 ;
  LAYER M2 ;
        RECT 24.56 25.604 24.72 25.636 ;
  LAYER M1 ;
        RECT 24.544 25.584 24.576 25.656 ;
  LAYER M2 ;
        RECT 24.524 25.604 24.596 25.636 ;
  LAYER M1 ;
        RECT 24.704 28.524 24.736 28.596 ;
  LAYER M2 ;
        RECT 24.684 28.544 24.756 28.576 ;
  LAYER M2 ;
        RECT 24.56 28.544 24.72 28.576 ;
  LAYER M1 ;
        RECT 24.544 28.524 24.576 28.596 ;
  LAYER M2 ;
        RECT 24.524 28.544 24.596 28.576 ;
  LAYER M1 ;
        RECT 24.544 19.2 24.576 19.272 ;
  LAYER M2 ;
        RECT 24.524 19.22 24.596 19.252 ;
  LAYER M1 ;
        RECT 24.544 19.236 24.576 19.404 ;
  LAYER M1 ;
        RECT 24.544 19.404 24.576 28.56 ;
  LAYER M2 ;
        RECT 21.68 19.22 24.56 19.252 ;
  LAYER M1 ;
        RECT 18.944 22.644 18.976 22.716 ;
  LAYER M2 ;
        RECT 18.924 22.664 18.996 22.696 ;
  LAYER M2 ;
        RECT 18.8 22.664 18.96 22.696 ;
  LAYER M1 ;
        RECT 18.784 22.644 18.816 22.716 ;
  LAYER M2 ;
        RECT 18.764 22.664 18.836 22.696 ;
  LAYER M1 ;
        RECT 18.944 31.464 18.976 31.536 ;
  LAYER M2 ;
        RECT 18.924 31.484 18.996 31.516 ;
  LAYER M2 ;
        RECT 18.8 31.484 18.96 31.516 ;
  LAYER M1 ;
        RECT 18.784 31.464 18.816 31.536 ;
  LAYER M2 ;
        RECT 18.764 31.484 18.836 31.516 ;
  LAYER M1 ;
        RECT 18.784 19.032 18.816 19.104 ;
  LAYER M2 ;
        RECT 18.764 19.052 18.836 19.084 ;
  LAYER M1 ;
        RECT 18.784 19.068 18.816 19.404 ;
  LAYER M1 ;
        RECT 18.784 19.404 18.816 31.5 ;
  LAYER M1 ;
        RECT 24.704 31.464 24.736 31.536 ;
  LAYER M2 ;
        RECT 24.684 31.484 24.756 31.516 ;
  LAYER M1 ;
        RECT 24.704 31.332 24.736 31.5 ;
  LAYER M1 ;
        RECT 24.704 31.296 24.736 31.368 ;
  LAYER M2 ;
        RECT 24.684 31.316 24.756 31.348 ;
  LAYER M2 ;
        RECT 24.72 31.316 27.44 31.348 ;
  LAYER M1 ;
        RECT 27.424 31.296 27.456 31.368 ;
  LAYER M2 ;
        RECT 27.404 31.316 27.476 31.348 ;
  LAYER M1 ;
        RECT 24.704 22.644 24.736 22.716 ;
  LAYER M2 ;
        RECT 24.684 22.664 24.756 22.696 ;
  LAYER M1 ;
        RECT 24.704 22.512 24.736 22.68 ;
  LAYER M1 ;
        RECT 24.704 22.476 24.736 22.548 ;
  LAYER M2 ;
        RECT 24.684 22.496 24.756 22.528 ;
  LAYER M2 ;
        RECT 24.72 22.496 27.44 22.528 ;
  LAYER M1 ;
        RECT 27.424 22.476 27.456 22.548 ;
  LAYER M2 ;
        RECT 27.404 22.496 27.476 22.528 ;
  LAYER M1 ;
        RECT 27.424 19.032 27.456 19.104 ;
  LAYER M2 ;
        RECT 27.404 19.052 27.476 19.084 ;
  LAYER M1 ;
        RECT 27.424 19.068 27.456 19.404 ;
  LAYER M1 ;
        RECT 27.424 19.404 27.456 31.332 ;
  LAYER M2 ;
        RECT 18.8 19.052 27.44 19.084 ;
  LAYER M1 ;
        RECT 21.824 31.464 21.856 31.536 ;
  LAYER M2 ;
        RECT 21.804 31.484 21.876 31.516 ;
  LAYER M2 ;
        RECT 21.84 31.484 24.72 31.516 ;
  LAYER M1 ;
        RECT 24.704 31.464 24.736 31.536 ;
  LAYER M2 ;
        RECT 24.684 31.484 24.756 31.516 ;
  LAYER M1 ;
        RECT 21.824 22.644 21.856 22.716 ;
  LAYER M2 ;
        RECT 21.804 22.664 21.876 22.696 ;
  LAYER M2 ;
        RECT 18.96 22.664 21.84 22.696 ;
  LAYER M1 ;
        RECT 18.944 22.644 18.976 22.716 ;
  LAYER M2 ;
        RECT 18.924 22.664 18.996 22.696 ;
  LAYER M1 ;
        RECT 16.064 34.404 16.096 34.476 ;
  LAYER M2 ;
        RECT 16.044 34.424 16.116 34.456 ;
  LAYER M2 ;
        RECT 15.92 34.424 16.08 34.456 ;
  LAYER M1 ;
        RECT 15.904 34.404 15.936 34.476 ;
  LAYER M2 ;
        RECT 15.884 34.424 15.956 34.456 ;
  LAYER M1 ;
        RECT 16.064 31.464 16.096 31.536 ;
  LAYER M2 ;
        RECT 16.044 31.484 16.116 31.516 ;
  LAYER M2 ;
        RECT 15.92 31.484 16.08 31.516 ;
  LAYER M1 ;
        RECT 15.904 31.464 15.936 31.536 ;
  LAYER M2 ;
        RECT 15.884 31.484 15.956 31.516 ;
  LAYER M1 ;
        RECT 16.064 28.524 16.096 28.596 ;
  LAYER M2 ;
        RECT 16.044 28.544 16.116 28.576 ;
  LAYER M2 ;
        RECT 15.92 28.544 16.08 28.576 ;
  LAYER M1 ;
        RECT 15.904 28.524 15.936 28.596 ;
  LAYER M2 ;
        RECT 15.884 28.544 15.956 28.576 ;
  LAYER M1 ;
        RECT 16.064 25.584 16.096 25.656 ;
  LAYER M2 ;
        RECT 16.044 25.604 16.116 25.636 ;
  LAYER M2 ;
        RECT 15.92 25.604 16.08 25.636 ;
  LAYER M1 ;
        RECT 15.904 25.584 15.936 25.656 ;
  LAYER M2 ;
        RECT 15.884 25.604 15.956 25.636 ;
  LAYER M1 ;
        RECT 16.064 22.644 16.096 22.716 ;
  LAYER M2 ;
        RECT 16.044 22.664 16.116 22.696 ;
  LAYER M2 ;
        RECT 15.92 22.664 16.08 22.696 ;
  LAYER M1 ;
        RECT 15.904 22.644 15.936 22.716 ;
  LAYER M2 ;
        RECT 15.884 22.664 15.956 22.696 ;
  LAYER M1 ;
        RECT 16.064 19.704 16.096 19.776 ;
  LAYER M2 ;
        RECT 16.044 19.724 16.116 19.756 ;
  LAYER M2 ;
        RECT 15.92 19.724 16.08 19.756 ;
  LAYER M1 ;
        RECT 15.904 19.704 15.936 19.776 ;
  LAYER M2 ;
        RECT 15.884 19.724 15.956 19.756 ;
  LAYER M1 ;
        RECT 15.904 18.864 15.936 18.936 ;
  LAYER M2 ;
        RECT 15.884 18.884 15.956 18.916 ;
  LAYER M1 ;
        RECT 15.904 18.9 15.936 19.404 ;
  LAYER M1 ;
        RECT 15.904 19.404 15.936 34.44 ;
  LAYER M1 ;
        RECT 27.584 34.404 27.616 34.476 ;
  LAYER M2 ;
        RECT 27.564 34.424 27.636 34.456 ;
  LAYER M1 ;
        RECT 27.584 34.272 27.616 34.44 ;
  LAYER M1 ;
        RECT 27.584 34.236 27.616 34.308 ;
  LAYER M2 ;
        RECT 27.564 34.256 27.636 34.288 ;
  LAYER M2 ;
        RECT 27.6 34.256 30.32 34.288 ;
  LAYER M1 ;
        RECT 30.304 34.236 30.336 34.308 ;
  LAYER M2 ;
        RECT 30.284 34.256 30.356 34.288 ;
  LAYER M1 ;
        RECT 27.584 31.464 27.616 31.536 ;
  LAYER M2 ;
        RECT 27.564 31.484 27.636 31.516 ;
  LAYER M1 ;
        RECT 27.584 31.332 27.616 31.5 ;
  LAYER M1 ;
        RECT 27.584 31.296 27.616 31.368 ;
  LAYER M2 ;
        RECT 27.564 31.316 27.636 31.348 ;
  LAYER M2 ;
        RECT 27.6 31.316 30.32 31.348 ;
  LAYER M1 ;
        RECT 30.304 31.296 30.336 31.368 ;
  LAYER M2 ;
        RECT 30.284 31.316 30.356 31.348 ;
  LAYER M1 ;
        RECT 27.584 28.524 27.616 28.596 ;
  LAYER M2 ;
        RECT 27.564 28.544 27.636 28.576 ;
  LAYER M1 ;
        RECT 27.584 28.392 27.616 28.56 ;
  LAYER M1 ;
        RECT 27.584 28.356 27.616 28.428 ;
  LAYER M2 ;
        RECT 27.564 28.376 27.636 28.408 ;
  LAYER M2 ;
        RECT 27.6 28.376 30.32 28.408 ;
  LAYER M1 ;
        RECT 30.304 28.356 30.336 28.428 ;
  LAYER M2 ;
        RECT 30.284 28.376 30.356 28.408 ;
  LAYER M1 ;
        RECT 27.584 25.584 27.616 25.656 ;
  LAYER M2 ;
        RECT 27.564 25.604 27.636 25.636 ;
  LAYER M1 ;
        RECT 27.584 25.452 27.616 25.62 ;
  LAYER M1 ;
        RECT 27.584 25.416 27.616 25.488 ;
  LAYER M2 ;
        RECT 27.564 25.436 27.636 25.468 ;
  LAYER M2 ;
        RECT 27.6 25.436 30.32 25.468 ;
  LAYER M1 ;
        RECT 30.304 25.416 30.336 25.488 ;
  LAYER M2 ;
        RECT 30.284 25.436 30.356 25.468 ;
  LAYER M1 ;
        RECT 27.584 22.644 27.616 22.716 ;
  LAYER M2 ;
        RECT 27.564 22.664 27.636 22.696 ;
  LAYER M1 ;
        RECT 27.584 22.512 27.616 22.68 ;
  LAYER M1 ;
        RECT 27.584 22.476 27.616 22.548 ;
  LAYER M2 ;
        RECT 27.564 22.496 27.636 22.528 ;
  LAYER M2 ;
        RECT 27.6 22.496 30.32 22.528 ;
  LAYER M1 ;
        RECT 30.304 22.476 30.336 22.548 ;
  LAYER M2 ;
        RECT 30.284 22.496 30.356 22.528 ;
  LAYER M1 ;
        RECT 27.584 19.704 27.616 19.776 ;
  LAYER M2 ;
        RECT 27.564 19.724 27.636 19.756 ;
  LAYER M1 ;
        RECT 27.584 19.572 27.616 19.74 ;
  LAYER M1 ;
        RECT 27.584 19.536 27.616 19.608 ;
  LAYER M2 ;
        RECT 27.564 19.556 27.636 19.588 ;
  LAYER M2 ;
        RECT 27.6 19.556 30.32 19.588 ;
  LAYER M1 ;
        RECT 30.304 19.536 30.336 19.608 ;
  LAYER M2 ;
        RECT 30.284 19.556 30.356 19.588 ;
  LAYER M1 ;
        RECT 30.304 18.864 30.336 18.936 ;
  LAYER M2 ;
        RECT 30.284 18.884 30.356 18.916 ;
  LAYER M1 ;
        RECT 30.304 18.9 30.336 19.404 ;
  LAYER M1 ;
        RECT 30.304 19.404 30.336 34.272 ;
  LAYER M2 ;
        RECT 15.92 18.884 30.32 18.916 ;
  LAYER M1 ;
        RECT 18.944 34.404 18.976 34.476 ;
  LAYER M2 ;
        RECT 18.924 34.424 18.996 34.456 ;
  LAYER M2 ;
        RECT 16.08 34.424 18.96 34.456 ;
  LAYER M1 ;
        RECT 16.064 34.404 16.096 34.476 ;
  LAYER M2 ;
        RECT 16.044 34.424 16.116 34.456 ;
  LAYER M1 ;
        RECT 18.944 19.704 18.976 19.776 ;
  LAYER M2 ;
        RECT 18.924 19.724 18.996 19.756 ;
  LAYER M2 ;
        RECT 16.08 19.724 18.96 19.756 ;
  LAYER M1 ;
        RECT 16.064 19.704 16.096 19.776 ;
  LAYER M2 ;
        RECT 16.044 19.724 16.116 19.756 ;
  LAYER M1 ;
        RECT 21.824 19.704 21.856 19.776 ;
  LAYER M2 ;
        RECT 21.804 19.724 21.876 19.756 ;
  LAYER M2 ;
        RECT 18.96 19.724 21.84 19.756 ;
  LAYER M1 ;
        RECT 18.944 19.704 18.976 19.776 ;
  LAYER M2 ;
        RECT 18.924 19.724 18.996 19.756 ;
  LAYER M1 ;
        RECT 24.704 19.704 24.736 19.776 ;
  LAYER M2 ;
        RECT 24.684 19.724 24.756 19.756 ;
  LAYER M2 ;
        RECT 21.84 19.724 24.72 19.756 ;
  LAYER M1 ;
        RECT 21.824 19.704 21.856 19.776 ;
  LAYER M2 ;
        RECT 21.804 19.724 21.876 19.756 ;
  LAYER M1 ;
        RECT 24.704 34.404 24.736 34.476 ;
  LAYER M2 ;
        RECT 24.684 34.424 24.756 34.456 ;
  LAYER M2 ;
        RECT 24.72 34.424 27.6 34.456 ;
  LAYER M1 ;
        RECT 27.584 34.404 27.616 34.476 ;
  LAYER M2 ;
        RECT 27.564 34.424 27.636 34.456 ;
  LAYER M1 ;
        RECT 21.824 34.404 21.856 34.476 ;
  LAYER M2 ;
        RECT 21.804 34.424 21.876 34.456 ;
  LAYER M2 ;
        RECT 21.84 34.424 24.72 34.456 ;
  LAYER M1 ;
        RECT 24.704 34.404 24.736 34.476 ;
  LAYER M2 ;
        RECT 24.684 34.424 24.756 34.456 ;
  LAYER M1 ;
        RECT 16.08 34.44 18.48 36.876 ;
  LAYER M2 ;
        RECT 16.08 34.44 18.48 36.876 ;
  LAYER M3 ;
        RECT 16.08 34.44 18.48 36.876 ;
  LAYER M1 ;
        RECT 16.08 31.5 18.48 33.936 ;
  LAYER M2 ;
        RECT 16.08 31.5 18.48 33.936 ;
  LAYER M3 ;
        RECT 16.08 31.5 18.48 33.936 ;
  LAYER M1 ;
        RECT 16.08 28.56 18.48 30.996 ;
  LAYER M2 ;
        RECT 16.08 28.56 18.48 30.996 ;
  LAYER M3 ;
        RECT 16.08 28.56 18.48 30.996 ;
  LAYER M1 ;
        RECT 16.08 25.62 18.48 28.056 ;
  LAYER M2 ;
        RECT 16.08 25.62 18.48 28.056 ;
  LAYER M3 ;
        RECT 16.08 25.62 18.48 28.056 ;
  LAYER M1 ;
        RECT 16.08 22.68 18.48 25.116 ;
  LAYER M2 ;
        RECT 16.08 22.68 18.48 25.116 ;
  LAYER M3 ;
        RECT 16.08 22.68 18.48 25.116 ;
  LAYER M1 ;
        RECT 16.08 19.74 18.48 22.176 ;
  LAYER M2 ;
        RECT 16.08 19.74 18.48 22.176 ;
  LAYER M3 ;
        RECT 16.08 19.74 18.48 22.176 ;
  LAYER M1 ;
        RECT 18.96 34.44 21.36 36.876 ;
  LAYER M2 ;
        RECT 18.96 34.44 21.36 36.876 ;
  LAYER M3 ;
        RECT 18.96 34.44 21.36 36.876 ;
  LAYER M1 ;
        RECT 18.96 31.5 21.36 33.936 ;
  LAYER M2 ;
        RECT 18.96 31.5 21.36 33.936 ;
  LAYER M3 ;
        RECT 18.96 31.5 21.36 33.936 ;
  LAYER M1 ;
        RECT 18.96 28.56 21.36 30.996 ;
  LAYER M2 ;
        RECT 18.96 28.56 21.36 30.996 ;
  LAYER M3 ;
        RECT 18.96 28.56 21.36 30.996 ;
  LAYER M1 ;
        RECT 18.96 25.62 21.36 28.056 ;
  LAYER M2 ;
        RECT 18.96 25.62 21.36 28.056 ;
  LAYER M3 ;
        RECT 18.96 25.62 21.36 28.056 ;
  LAYER M1 ;
        RECT 18.96 22.68 21.36 25.116 ;
  LAYER M2 ;
        RECT 18.96 22.68 21.36 25.116 ;
  LAYER M3 ;
        RECT 18.96 22.68 21.36 25.116 ;
  LAYER M1 ;
        RECT 18.96 19.74 21.36 22.176 ;
  LAYER M2 ;
        RECT 18.96 19.74 21.36 22.176 ;
  LAYER M3 ;
        RECT 18.96 19.74 21.36 22.176 ;
  LAYER M1 ;
        RECT 21.84 34.44 24.24 36.876 ;
  LAYER M2 ;
        RECT 21.84 34.44 24.24 36.876 ;
  LAYER M3 ;
        RECT 21.84 34.44 24.24 36.876 ;
  LAYER M1 ;
        RECT 21.84 31.5 24.24 33.936 ;
  LAYER M2 ;
        RECT 21.84 31.5 24.24 33.936 ;
  LAYER M3 ;
        RECT 21.84 31.5 24.24 33.936 ;
  LAYER M1 ;
        RECT 21.84 28.56 24.24 30.996 ;
  LAYER M2 ;
        RECT 21.84 28.56 24.24 30.996 ;
  LAYER M3 ;
        RECT 21.84 28.56 24.24 30.996 ;
  LAYER M1 ;
        RECT 21.84 25.62 24.24 28.056 ;
  LAYER M2 ;
        RECT 21.84 25.62 24.24 28.056 ;
  LAYER M3 ;
        RECT 21.84 25.62 24.24 28.056 ;
  LAYER M1 ;
        RECT 21.84 22.68 24.24 25.116 ;
  LAYER M2 ;
        RECT 21.84 22.68 24.24 25.116 ;
  LAYER M3 ;
        RECT 21.84 22.68 24.24 25.116 ;
  LAYER M1 ;
        RECT 21.84 19.74 24.24 22.176 ;
  LAYER M2 ;
        RECT 21.84 19.74 24.24 22.176 ;
  LAYER M3 ;
        RECT 21.84 19.74 24.24 22.176 ;
  LAYER M1 ;
        RECT 24.72 34.44 27.12 36.876 ;
  LAYER M2 ;
        RECT 24.72 34.44 27.12 36.876 ;
  LAYER M3 ;
        RECT 24.72 34.44 27.12 36.876 ;
  LAYER M1 ;
        RECT 24.72 31.5 27.12 33.936 ;
  LAYER M2 ;
        RECT 24.72 31.5 27.12 33.936 ;
  LAYER M3 ;
        RECT 24.72 31.5 27.12 33.936 ;
  LAYER M1 ;
        RECT 24.72 28.56 27.12 30.996 ;
  LAYER M2 ;
        RECT 24.72 28.56 27.12 30.996 ;
  LAYER M3 ;
        RECT 24.72 28.56 27.12 30.996 ;
  LAYER M1 ;
        RECT 24.72 25.62 27.12 28.056 ;
  LAYER M2 ;
        RECT 24.72 25.62 27.12 28.056 ;
  LAYER M3 ;
        RECT 24.72 25.62 27.12 28.056 ;
  LAYER M1 ;
        RECT 24.72 22.68 27.12 25.116 ;
  LAYER M2 ;
        RECT 24.72 22.68 27.12 25.116 ;
  LAYER M3 ;
        RECT 24.72 22.68 27.12 25.116 ;
  LAYER M1 ;
        RECT 24.72 19.74 27.12 22.176 ;
  LAYER M2 ;
        RECT 24.72 19.74 27.12 22.176 ;
  LAYER M3 ;
        RECT 24.72 19.74 27.12 22.176 ;
  LAYER M1 ;
        RECT 27.6 34.44 30 36.876 ;
  LAYER M2 ;
        RECT 27.6 34.44 30 36.876 ;
  LAYER M3 ;
        RECT 27.6 34.44 30 36.876 ;
  LAYER M1 ;
        RECT 27.6 31.5 30 33.936 ;
  LAYER M2 ;
        RECT 27.6 31.5 30 33.936 ;
  LAYER M3 ;
        RECT 27.6 31.5 30 33.936 ;
  LAYER M1 ;
        RECT 27.6 28.56 30 30.996 ;
  LAYER M2 ;
        RECT 27.6 28.56 30 30.996 ;
  LAYER M3 ;
        RECT 27.6 28.56 30 30.996 ;
  LAYER M1 ;
        RECT 27.6 25.62 30 28.056 ;
  LAYER M2 ;
        RECT 27.6 25.62 30 28.056 ;
  LAYER M3 ;
        RECT 27.6 25.62 30 28.056 ;
  LAYER M1 ;
        RECT 27.6 22.68 30 25.116 ;
  LAYER M2 ;
        RECT 27.6 22.68 30 25.116 ;
  LAYER M3 ;
        RECT 27.6 22.68 30 25.116 ;
  LAYER M1 ;
        RECT 27.6 19.74 30 22.176 ;
  LAYER M2 ;
        RECT 27.6 19.74 30 22.176 ;
  LAYER M3 ;
        RECT 27.6 19.74 30 22.176 ;
  END 
END switched_capacitor_filter
