.subckt BUFFER_VREFP_FINAL2 gnd ibias sw<2> sw<1> sw<0> vdd vref vrefp
xm58 vrefp net459 net0129 vdd pfet_lvt w=w0 l=l0
xm43 net0125 net431 vrefp vdd pfet_lvt w=w1 l=l0
xm15 vfb net450 net0115 vdd pfet_lvt w=w2 l=l0
xm28 vrefp net459 net0127 vdd pfet_lvt w=w3 l=l0
xm27 net431 net431 vfb vdd pfet_lvt w=w4 l=l0
xm29 net459 net431 vrefp vdd pfet_lvt w=w5 l=l0
xm106 vdd net431 vdd vdd pfet_lvt w=w6 l=l1
xm32 net0132 net431 vrefp vdd pfet_lvt w=w5 l=l0
xm33 vrefp net459 net0113 vdd pfet_lvt w=w7 l=l0
xm34 vrefp net459 net0135 vdd pfet_lvt w=w8 l=l0
xm35 net0134 net431 vrefp vdd pfet_lvt w=w9 l=l0
xm62 swn2 swp2 gnd gnd nfet w=w10 l=l2
xm59 swp2 sw<2> gnd gnd nfet w=w10 l=l2
xm57 net0125 ibias net468 gnd nfet w=w11 l=l0
xm55 net468 swn2 gnd gnd nfet w=w12 l=l2
xm54 swn1 swp1 gnd gnd nfet w=w10 l=l2
xm51 swp1 sw<1> gnd gnd nfet w=w10 l=l2
xm50 swn0 swp0 gnd gnd nfet w=w10 l=l2
xm48 swp0 sw<0> gnd gnd nfet w=w10 l=l2
xm20 net469 swn1 gnd gnd nfet w=w13 l=l2
xm19 net470 swn0 gnd gnd nfet w=w13 l=l2
xm18 net463 vdd gnd gnd nfet w=w14 l=l2
xm17 net427 vdd gnd gnd nfet w=w15 l=l2
xm16 net462 vdd gnd gnd nfet w=w15 l=l2
xm9 net466 vdd gnd gnd nfet w=w15 l=l2
xm7 net467 vdd gnd gnd nfet w=w15 l=l2
xm2 net465 vdd gnd gnd nfet w=w15 l=l2
xm0 net464 vdd gnd gnd nfet w=w16 l=l2
xm6 net450 net412 net462 gnd nfet w=w17 l=l2
xm1 net412 net412 net467 gnd nfet w=w17 l=l2
xm3 net418 ibias net466 gnd nfet w=w18 l=l0
xm4 ibias ibias net464 gnd nfet w=w19 l=l0
xm5 net411 ibias net465 gnd nfet w=w19 l=l0
xm8 net423 vfb net418 gnd nfet w=w20 l=l0
xm10 net412 vfb net418 gnd nfet w=w20 l=l0
xm11 net417 vref net418 gnd nfet w=w20 l=l0
xm12 net450 vref net418 gnd nfet w=w20 l=l0
xm21 net431 ibias net427 net427 nfet w=w19 l=l0
xm30 net459 ibias net463 gnd nfet w=w21 l=l0
xm31 net0132 ibias net470 gnd nfet w=w21 l=l0
xm36 net0134 ibias net469 gnd nfet w=w22 l=l0
xm61 swn2 swp2 vdd vdd pfet w=w23 l=l2
xm60 swp2 sw<2> vdd vdd pfet w=w23 l=l2
xm53 swn1 swp1 vdd vdd pfet w=w23 l=l2
xm52 swp1 sw<1> vdd vdd pfet w=w23 l=l2
xm49 swn0 swp0 vdd vdd pfet w=w23 l=l2
xm47 swp0 sw<0> vdd vdd pfet w=w23 l=l2
xm46 net0135 swp1 vdd vdd pfet w=w24 l=l2
xm45 net0113 swp0 vdd vdd pfet w=w25 l=l2
xm44 net0127 gnd vdd vdd pfet w=w25 l=l2
xm56 net0129 swp2 vdd vdd pfet w=w26 l=l2
xm42 net0115 gnd vdd vdd pfet w=w27 l=l2
xm41 net0124 gnd vdd vdd pfet w=w27 l=l2
xm40 net0119 gnd vdd vdd pfet w=w27 l=l2
xm39 net0114 gnd vdd vdd pfet w=w27 l=l2
xm38 net0128 gnd vdd vdd pfet w=w27 l=l2
xm37 net0121 gnd vdd vdd pfet w=w13 l=l2
xm13 net450 net411 net0137 vdd pfet w=w28 l=l0
xm14 net412 net411 net0122 vdd pfet w=w28 l=l0
xm22 net411 net411 net0121 vdd pfet w=w17 l=l0
xm23 net423 net423 net0114 vdd pfet w=w29 l=l0
xm24 net0137 net423 net0124 vdd pfet w=w11 l=l0
xm25 net417 net417 net0119 vdd pfet w=w29 l=l0
xm26 net0122 net417 net0128 vdd pfet w=w11 l=l0
.ends BUFFER_VREFP_FINAL2

