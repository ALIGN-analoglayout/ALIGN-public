VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

VIA M4_M3_0
  VIARULE M4_M3 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M3 VIA3 M4 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 1 ;
END M4_M3_0

VIA M4_M3_1
  VIARULE M4_M3 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M3 VIA3 M4 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 20 ;
END M4_M3_1

VIA M3_M2_2
  VIARULE M3_M2 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M2 VIA2 M3 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 1 ;
END M3_M2_2

VIA M3_M2_3
  VIARULE M3_M2 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M2 VIA2 M3 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 20 ;
END M3_M2_3

VIA M2_M1_4
  VIARULE M2_M1 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M1 VIA1 M2 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 1 ;
END M2_M1_4

VIA M2_M1_5
  VIARULE M2_M1 ;
  CUTSIZE 0.1 0.1 ;
  LAYERS M1 VIA1 M2 ;
  CUTSPACING 0.1 0.1 ;
  ENCLOSURE 0.04 0.04 0.04 0.04 ;
  ROWCOL 1 20 ;
END M2_M1_5

MACRO SW_NMOS_wr2u_lr60n_nr16
  ORIGIN 0 0 ;
  FOREIGN SW_NMOS_wr2u_lr60n_nr16 0 0 ;
  SIZE 10 BY 7.54 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2.435 2.24 7.565 4.41 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8.02 2.695 8.2 4.78 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.65 5.24 7.35 6.54 ;
    END
  END D
  PIN DNWP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.76 1.03 8.97 6.29 ;
    END
  END DNWP
  OBS
    LAYER M1 ;
      RECT 1 1 8.61 6.51 ;
    LAYER M2 ;
      RECT 1.785 1.53 8.2 5.04 ;
    LAYER M3 ;
      RECT 1.785 2.5 7.93 5.04 ;
  END
END SW_NMOS_wr2u_lr60n_nr16

END LIBRARY
