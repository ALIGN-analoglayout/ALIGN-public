
.subckt dummy_hier_CK<10> CK<11> VALIDC CK<10> CKSBTB DVSS DVDD CK<9>
XI213 DVSS DVDD CK<11> CK<10> VALIDC CKSBTB DFFRB_B_V6_HVT
XI214 DVSS DVDD CK<10> VALIDC CKSBTB CK<9> DFFRB_B_V6_HVT
.ends dummy_hier_CK<10>

.subckt dummy_hier_TGC<8> TGC<8> SWC<8> CKSBT DVSS DVDD CK<8>
XI101 DVSS DVDD SWC<8> TGC<8> CKSBT NR2D1LVT
XI156 DVSS DVDD TGC<8> CKSBT CK<8> NR2D1LVT
.ends dummy_hier_TGC<8>

.subckt dummy_hier_TGC<10> SWC<10> CKSBT DVSS DVDD TGC<10> CK<10>
XI105 DVSS DVDD SWC<10> TGC<10> CKSBT NR2D1LVT
XI171 DVSS DVDD TGC<10> CKSBT CK<10> NR2D1LVT
.ends dummy_hier_TGC<10>

.subckt dummy_hier_TGC<11> CK<11> TGC<11> CKSBT DVSS DVDD SWC<11>
XI175 DVSS DVDD CK<11> TGC<11> CKSBT NR2D1LVT
XI107 DVSS DVDD TGC<11> CKSBT SWC<11> NR2D1LVT
.ends dummy_hier_TGC<11>

.subckt dummy_hier_TGC<9> TGC<9> CKSBT DVSS DVDD CK<9> SWC<9>
XI159 DVSS DVDD CK<9> TGC<9> CKSBT NR2D1LVT
XI39 DVSS DVDD TGC<9> CKSBT SWC<9> NR2D1LVT
.ends dummy_hier_TGC<9>

.subckt Sanitized_Coarse_SAR_Logic CPY OUTNC DVSS DVDD CK<8> DB<8> D<8> CK<11> OUTPC D<11> DB<11> CK<10> D<10> DB<10> CK<9> DB<9> D<9> DFB<7> DF<7> DF<8> DFB<8> DFB<9> DF<9> DF<10> DFB<10> TGC<11> TGCB<11> SWC<11> SWCB<11> SWC<10> SWCB<10> TGC<10> TGCB<10> TGC<9> TGCB<9> SWC<9> SWCB<9> SWC<8> SWCB<8> TGC<8> TGCB<8> DFB<11> DF<11> CKSBT VALIDC ST_FINE CKSBTB
XI228 CPY OUTNC DVSS DVDD net057 net018 DFF_HVT_Coarse
XI227 CK<8> OUTNC DVSS DVDD DB<8> D<8> DFF_HVT_Coarse
XI229 CK<11> OUTPC DVSS DVDD D<11> DB<11> DFF_HVT_Coarse
XI230 CK<10> OUTPC DVSS DVDD D<10> DB<10> DFF_HVT_Coarse
XI231 CK<9> OUTNC DVSS DVDD DB<9> D<9> DFF_HVT_Coarse
XI18 net018 DFB<7> DVDD DVSS INVD1LVT
XI17 net057 DF<7> DVDD DVSS INVD1LVT
XI16 DB<8> DF<8> DVDD DVSS INVD1LVT
XI15 D<8> DFB<8> DVDD DVSS INVD1LVT
XI14 D<9> DFB<9> DVDD DVSS INVD1LVT
XI13 DB<9> DF<9> DVDD DVSS INVD1LVT
XI12 DB<10> DF<10> DVDD DVSS INVD1LVT
XI11 D<10> DFB<10> DVDD DVSS INVD1LVT
XI173 TGC<11> TGCB<11> DVDD DVSS INVD1LVT
XI31 SWC<11> SWCB<11> DVDD DVSS INVD1LVT
XI104 SWC<10> SWCB<10> DVDD DVSS INVD1LVT
XI170 TGC<10> TGCB<10> DVDD DVSS INVD1LVT
XI158 TGC<9> TGCB<9> DVDD DVSS INVD1LVT
XI102 SWC<9> SWCB<9> DVDD DVSS INVD1LVT
XI100 SWC<8> SWCB<8> DVDD DVSS INVD1LVT
XI155 TGC<8> TGCB<8> DVDD DVSS INVD1LVT
XI9 D<11> DFB<11> DVDD DVSS INVD1LVT
XI10 DB<11> DF<11> DVDD DVSS INVD1LVT
XI8 net054 DVDD DVSS TIEHLVT
XI53 VALIDC net133 DVDD DVSS ST_FINE CKSBTB DFFRB_B_V6_HVT
XI54 VALIDC CPY DVDD DVSS net133 CKSBTB DFFRB_B_V6_HVT
XI212 VALIDC net054 DVDD DVSS CK<11> CKSBTB DFFRB_B_V6_HVT
XI215 VALIDC CK<9> DVDD DVSS CK<8> CKSBTB DFFRB_B_V6_HVT
XI216 VALIDC CK<8> DVDD DVSS CPY CKSBTB DFFRB_B_V6_HVT
XI213_XI214 VALIDC CK<10> CKSBTB DVSS DVDD CK<9> CK<11> dummy_hier_CK<10>
XI101_XI156 SWC<8> CKSBT DVSS DVDD CK<8> TGC<8> dummy_hier_TGC<8>
XI105_XI171 CKSBT DVSS DVDD TGC<10> CK<10> SWC<10> dummy_hier_TGC<10>
XI175_XI107 TGC<11> CKSBT DVSS DVDD SWC<11> CK<11> dummy_hier_TGC<11>
XI159_XI39 CKSBT DVSS DVDD CK<9> SWC<9> TGC<9> dummy_hier_TGC<9>
.ends Sanitized_Coarse_SAR_Logic

.subckt DP_NMOS_n12_X1_Y1 B DA GA S DB GB
xM0 DA GA S B Switch_NMOS_n12_X1_Y1
xM1 DB GB S B Switch_NMOS_n12_X1_Y1
.ends DP_NMOS_n12_X1_Y1

.subckt Switch_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_NMOS_n12_X1_Y1

.subckt DP_PMOS_n12_X1_Y1 B DA GA S DB GB
xM0 DA GA S B Switch_PMOS_n12_X1_Y1
xM1 DB GB S B Switch_PMOS_n12_X1_Y1
.ends DP_PMOS_n12_X1_Y1

.subckt Switch_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_PMOS_n12_X1_Y1

.subckt DFF_HVT_Coarse CK D DGND DVDD Q QN
xMM2 QN CK NET4 DGND Switch_NMOS_n12_X1_Y1
xMM7 Q QN DGND DGND Switch_NMOS_n12_X1_Y1
xMM4 NET2 N1 NET3 DGND Switch_NMOS_n12_X1_Y1
xMM3 NET4 NET2 DGND DGND Switch_NMOS_n12_X1_Y1
xMM12 Q QN DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM11 QN NET2 DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM15 N1 CK NET1 DVDD Switch_PMOS_n12_X1_Y1
xMM13_MM14 N1 D DGND NET3 CK DGND DP_NMOS_n12_X1_Y1
xMM8_MM9 NET1 D DVDD NET2 CK DVDD DP_PMOS_n12_X1_Y1
.ends DFF_HVT_Coarse

.subckt DP_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends DP_NMOS_n12_X1_Y1

.subckt DP_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends DP_PMOS_n12_X1_Y1

.subckt INVD1LVT I ZN VDD VSS
xMMU1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD1LVT

.subckt TIEHLVT Z VDD VSS
xMM_u2 net7 net7 VSS VSS DCL_NMOS_n12_X1_Y1
xMM_u1 Z net7 VDD VDD Switch_PMOS_n12_X1_Y1
.ends TIEHLVT

.subckt DCL_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends DCL_NMOS_n12_X1_Y1

.subckt NR2D1LVT A1 A2 ZN VDD VSS
xMMI1_M_u3 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u4 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI1_M_u1 net13 A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMI1_M_u2 ZN A1 net13 VDD Switch_PMOS_n12_X1_Y1
.ends NR2D1LVT

.subckt DFFRB_B_V6_HVT CK D DVDD DVSS Q RST
xMM8 NET1 D DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM10 NET2 CK net58 DVDD Switch_PMOS_n12_X1_Y1
xMM19 net58 RSTB DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM15 net06 RST DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM9 M1 CK NET1 DVDD Switch_PMOS_n12_X1_Y1
xMM14 Q net06 DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM12 net06 NET2 DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM0 RSTB RST DVDD DVDD Switch_PMOS_n12_X1_Y1
xMM16 NET3 CK DVSS DVSS Switch_NMOS_n12_X1_Y1
xMM13 NET4 NET2 DVSS DVSS Switch_NMOS_n12_X1_Y1
xMM7 Q net06 DVSS DVSS Switch_NMOS_n12_X1_Y1
xMM6 net06 CK NET4 DVSS Switch_NMOS_n12_X1_Y1
xMM17 M1 D DVSS DVSS Switch_NMOS_n12_X1_Y1
xMM5 NET2 RSTB DVSS DVSS Switch_NMOS_n12_X1_Y1
xMM4 NET2 M1 NET3 DVSS Switch_NMOS_n12_X1_Y1
xMM18 RSTB RST DVSS DVSS Switch_NMOS_n12_X1_Y1
.ends DFFRB_B_V6_HVT
