MACRO cap_12f
  ORIGIN 0 0 ;
  FOREIGN cap_12f 0 0 ;
  SIZE 2.4960 BY 2.6040 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 0.0680 2.4680 0.1000 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0280 2.5040 2.4680 2.5360 ;
    END
  END MINUS
  OBS
    LAYER M1 ;
      RECT 0.0480 0.0480 0.0800 2.5560 ;
    LAYER M3 ;
      RECT 0.0480 0.0480 0.0800 2.5560 ;
    LAYER V1 ;
      RECT 0.0480 2.5040 0.0800 2.5360 ;
    LAYER V1 ;
      RECT 0.0480 2.5040 0.0800 2.5360 ;
    LAYER M1 ;
      RECT 0.1120 0.0480 0.1440 2.5560 ;
    LAYER M3 ;
      RECT 0.1120 0.0480 0.1440 2.5560 ;
    LAYER V1 ;
      RECT 0.1120 0.0680 0.1440 0.1000 ;
    LAYER V1 ;
      RECT 0.1120 0.0680 0.1440 0.1000 ;
    LAYER M1 ;
      RECT 0.1760 0.0480 0.2080 2.5560 ;
    LAYER M3 ;
      RECT 0.1760 0.0480 0.2080 2.5560 ;
    LAYER V1 ;
      RECT 0.1760 2.5040 0.2080 2.5360 ;
    LAYER V1 ;
      RECT 0.1760 2.5040 0.2080 2.5360 ;
    LAYER M1 ;
      RECT 0.2400 0.0480 0.2720 2.5560 ;
    LAYER M3 ;
      RECT 0.2400 0.0480 0.2720 2.5560 ;
    LAYER V1 ;
      RECT 0.2400 0.0680 0.2720 0.1000 ;
    LAYER V1 ;
      RECT 0.2400 0.0680 0.2720 0.1000 ;
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 2.5560 ;
    LAYER M3 ;
      RECT 0.3040 0.0480 0.3360 2.5560 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER V1 ;
      RECT 0.3040 2.5040 0.3360 2.5360 ;
    LAYER M1 ;
      RECT 0.3680 0.0480 0.4000 2.5560 ;
    LAYER M3 ;
      RECT 0.3680 0.0480 0.4000 2.5560 ;
    LAYER V1 ;
      RECT 0.3680 0.0680 0.4000 0.1000 ;
    LAYER V1 ;
      RECT 0.3680 0.0680 0.4000 0.1000 ;
    LAYER M1 ;
      RECT 0.4320 0.0480 0.4640 2.5560 ;
    LAYER M3 ;
      RECT 0.4320 0.0480 0.4640 2.5560 ;
    LAYER V1 ;
      RECT 0.4320 2.5040 0.4640 2.5360 ;
    LAYER V1 ;
      RECT 0.4320 2.5040 0.4640 2.5360 ;
    LAYER M1 ;
      RECT 0.4960 0.0480 0.5280 2.5560 ;
    LAYER M3 ;
      RECT 0.4960 0.0480 0.5280 2.5560 ;
    LAYER V1 ;
      RECT 0.4960 0.0680 0.5280 0.1000 ;
    LAYER V1 ;
      RECT 0.4960 0.0680 0.5280 0.1000 ;
    LAYER M1 ;
      RECT 0.5600 0.0480 0.5920 2.5560 ;
    LAYER M3 ;
      RECT 0.5600 0.0480 0.5920 2.5560 ;
    LAYER V1 ;
      RECT 0.5600 2.5040 0.5920 2.5360 ;
    LAYER V1 ;
      RECT 0.5600 2.5040 0.5920 2.5360 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 2.5560 ;
    LAYER M3 ;
      RECT 0.6240 0.0480 0.6560 2.5560 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER M1 ;
      RECT 0.6880 0.0480 0.7200 2.5560 ;
    LAYER M3 ;
      RECT 0.6880 0.0480 0.7200 2.5560 ;
    LAYER V1 ;
      RECT 0.6880 2.5040 0.7200 2.5360 ;
    LAYER V1 ;
      RECT 0.6880 2.5040 0.7200 2.5360 ;
    LAYER M1 ;
      RECT 0.7520 0.0480 0.7840 2.5560 ;
    LAYER M3 ;
      RECT 0.7520 0.0480 0.7840 2.5560 ;
    LAYER V1 ;
      RECT 0.7520 0.0680 0.7840 0.1000 ;
    LAYER V1 ;
      RECT 0.7520 0.0680 0.7840 0.1000 ;
    LAYER M1 ;
      RECT 0.8160 0.0480 0.8480 2.5560 ;
    LAYER M3 ;
      RECT 0.8160 0.0480 0.8480 2.5560 ;
    LAYER V1 ;
      RECT 0.8160 2.5040 0.8480 2.5360 ;
    LAYER V1 ;
      RECT 0.8160 2.5040 0.8480 2.5360 ;
    LAYER M1 ;
      RECT 0.8800 0.0480 0.9120 2.5560 ;
    LAYER M3 ;
      RECT 0.8800 0.0480 0.9120 2.5560 ;
    LAYER V1 ;
      RECT 0.8800 0.0680 0.9120 0.1000 ;
    LAYER V1 ;
      RECT 0.8800 0.0680 0.9120 0.1000 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 2.5560 ;
    LAYER M3 ;
      RECT 0.9440 0.0480 0.9760 2.5560 ;
    LAYER V1 ;
      RECT 0.9440 2.5040 0.9760 2.5360 ;
    LAYER V1 ;
      RECT 0.9440 2.5040 0.9760 2.5360 ;
    LAYER M1 ;
      RECT 1.0080 0.0480 1.0400 2.5560 ;
    LAYER M3 ;
      RECT 1.0080 0.0480 1.0400 2.5560 ;
    LAYER V1 ;
      RECT 1.0080 0.0680 1.0400 0.1000 ;
    LAYER V1 ;
      RECT 1.0080 0.0680 1.0400 0.1000 ;
    LAYER M1 ;
      RECT 1.0720 0.0480 1.1040 2.5560 ;
    LAYER M3 ;
      RECT 1.0720 0.0480 1.1040 2.5560 ;
    LAYER V1 ;
      RECT 1.0720 2.5040 1.1040 2.5360 ;
    LAYER V1 ;
      RECT 1.0720 2.5040 1.1040 2.5360 ;
    LAYER M1 ;
      RECT 1.1360 0.0480 1.1680 2.5560 ;
    LAYER M3 ;
      RECT 1.1360 0.0480 1.1680 2.5560 ;
    LAYER V1 ;
      RECT 1.1360 0.0680 1.1680 0.1000 ;
    LAYER V1 ;
      RECT 1.1360 0.0680 1.1680 0.1000 ;
    LAYER M1 ;
      RECT 1.2000 0.0480 1.2320 2.5560 ;
    LAYER M3 ;
      RECT 1.2000 0.0480 1.2320 2.5560 ;
    LAYER V1 ;
      RECT 1.2000 2.5040 1.2320 2.5360 ;
    LAYER V1 ;
      RECT 1.2000 2.5040 1.2320 2.5360 ;
    LAYER M1 ;
      RECT 1.2640 0.0480 1.2960 2.5560 ;
    LAYER M3 ;
      RECT 1.2640 0.0480 1.2960 2.5560 ;
    LAYER V1 ;
      RECT 1.2640 0.0680 1.2960 0.1000 ;
    LAYER V1 ;
      RECT 1.2640 0.0680 1.2960 0.1000 ;
    LAYER M1 ;
      RECT 1.3280 0.0480 1.3600 2.5560 ;
    LAYER M3 ;
      RECT 1.3280 0.0480 1.3600 2.5560 ;
    LAYER V1 ;
      RECT 1.3280 2.5040 1.3600 2.5360 ;
    LAYER V1 ;
      RECT 1.3280 2.5040 1.3600 2.5360 ;
    LAYER M1 ;
      RECT 1.3920 0.0480 1.4240 2.5560 ;
    LAYER M3 ;
      RECT 1.3920 0.0480 1.4240 2.5560 ;
    LAYER V1 ;
      RECT 1.3920 0.0680 1.4240 0.1000 ;
    LAYER V1 ;
      RECT 1.3920 0.0680 1.4240 0.1000 ;
    LAYER M1 ;
      RECT 1.4560 0.0480 1.4880 2.5560 ;
    LAYER M3 ;
      RECT 1.4560 0.0480 1.4880 2.5560 ;
    LAYER V1 ;
      RECT 1.4560 2.5040 1.4880 2.5360 ;
    LAYER V1 ;
      RECT 1.4560 2.5040 1.4880 2.5360 ;
    LAYER M1 ;
      RECT 1.5200 0.0480 1.5520 2.5560 ;
    LAYER M3 ;
      RECT 1.5200 0.0480 1.5520 2.5560 ;
    LAYER V1 ;
      RECT 1.5200 0.0680 1.5520 0.1000 ;
    LAYER V1 ;
      RECT 1.5200 0.0680 1.5520 0.1000 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 2.5560 ;
    LAYER M3 ;
      RECT 1.5840 0.0480 1.6160 2.5560 ;
    LAYER V1 ;
      RECT 1.5840 2.5040 1.6160 2.5360 ;
    LAYER V1 ;
      RECT 1.5840 2.5040 1.6160 2.5360 ;
    LAYER M1 ;
      RECT 1.6480 0.0480 1.6800 2.5560 ;
    LAYER M3 ;
      RECT 1.6480 0.0480 1.6800 2.5560 ;
    LAYER V1 ;
      RECT 1.6480 0.0680 1.6800 0.1000 ;
    LAYER V1 ;
      RECT 1.6480 0.0680 1.6800 0.1000 ;
    LAYER M1 ;
      RECT 1.7120 0.0480 1.7440 2.5560 ;
    LAYER M3 ;
      RECT 1.7120 0.0480 1.7440 2.5560 ;
    LAYER V1 ;
      RECT 1.7120 2.5040 1.7440 2.5360 ;
    LAYER V1 ;
      RECT 1.7120 2.5040 1.7440 2.5360 ;
    LAYER M1 ;
      RECT 1.7760 0.0480 1.8080 2.5560 ;
    LAYER M3 ;
      RECT 1.7760 0.0480 1.8080 2.5560 ;
    LAYER V1 ;
      RECT 1.7760 0.0680 1.8080 0.1000 ;
    LAYER V1 ;
      RECT 1.7760 0.0680 1.8080 0.1000 ;
    LAYER M1 ;
      RECT 1.8400 0.0480 1.8720 2.5560 ;
    LAYER M3 ;
      RECT 1.8400 0.0480 1.8720 2.5560 ;
    LAYER V1 ;
      RECT 1.8400 2.5040 1.8720 2.5360 ;
    LAYER V1 ;
      RECT 1.8400 2.5040 1.8720 2.5360 ;
    LAYER M1 ;
      RECT 1.9040 0.0480 1.9360 2.5560 ;
    LAYER M3 ;
      RECT 1.9040 0.0480 1.9360 2.5560 ;
    LAYER V1 ;
      RECT 1.9040 0.0680 1.9360 0.1000 ;
    LAYER V1 ;
      RECT 1.9040 0.0680 1.9360 0.1000 ;
    LAYER M1 ;
      RECT 1.9680 0.0480 2.0000 2.5560 ;
    LAYER M3 ;
      RECT 1.9680 0.0480 2.0000 2.5560 ;
    LAYER V1 ;
      RECT 1.9680 2.5040 2.0000 2.5360 ;
    LAYER V1 ;
      RECT 1.9680 2.5040 2.0000 2.5360 ;
    LAYER M1 ;
      RECT 2.0320 0.0480 2.0640 2.5560 ;
    LAYER M3 ;
      RECT 2.0320 0.0480 2.0640 2.5560 ;
    LAYER V1 ;
      RECT 2.0320 0.0680 2.0640 0.1000 ;
    LAYER V1 ;
      RECT 2.0320 0.0680 2.0640 0.1000 ;
    LAYER M1 ;
      RECT 2.0960 0.0480 2.1280 2.5560 ;
    LAYER M3 ;
      RECT 2.0960 0.0480 2.1280 2.5560 ;
    LAYER V1 ;
      RECT 2.0960 2.5040 2.1280 2.5360 ;
    LAYER V1 ;
      RECT 2.0960 2.5040 2.1280 2.5360 ;
    LAYER M1 ;
      RECT 2.1600 0.0480 2.1920 2.5560 ;
    LAYER M3 ;
      RECT 2.1600 0.0480 2.1920 2.5560 ;
    LAYER V1 ;
      RECT 2.1600 0.0680 2.1920 0.1000 ;
    LAYER V1 ;
      RECT 2.1600 0.0680 2.1920 0.1000 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 2.5560 ;
    LAYER M3 ;
      RECT 2.2240 0.0480 2.2560 2.5560 ;
    LAYER V1 ;
      RECT 2.2240 2.5040 2.2560 2.5360 ;
    LAYER V1 ;
      RECT 2.2240 2.5040 2.2560 2.5360 ;
    LAYER M1 ;
      RECT 2.2880 0.0480 2.3200 2.5560 ;
    LAYER M3 ;
      RECT 2.2880 0.0480 2.3200 2.5560 ;
    LAYER V1 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER V1 ;
      RECT 2.2880 0.0680 2.3200 0.1000 ;
    LAYER M1 ;
      RECT 2.3520 0.0480 2.3840 2.5560 ;
    LAYER M3 ;
      RECT 2.3520 0.0480 2.3840 2.5560 ;
    LAYER V1 ;
      RECT 2.3520 2.5040 2.3840 2.5360 ;
    LAYER V1 ;
      RECT 2.3520 2.5040 2.3840 2.5360 ;
    LAYER M1 ;
      RECT 2.4160 0.0480 2.4480 2.5560 ;
    LAYER M3 ;
      RECT 2.4160 0.0480 2.4480 2.5560 ;
    LAYER V1 ;
      RECT 2.4160 0.0680 2.4480 0.1000 ;
    LAYER V1 ;
      RECT 2.4160 0.0680 2.4480 0.1000 ;
    LAYER V1 ;
      RECT 2.4160 0.0680 2.4480 0.1000 ;
    LAYER V2 ;
      RECT 2.4160 0.0680 2.4480 0.1000 ;
    LAYER V1 ;
      RECT 0.0480 0.1320 0.0800 0.1640 ;
    LAYER V2 ;
      RECT 0.0480 0.1320 0.0800 0.1640 ;
    LAYER M2 ;
      RECT 0.0280 0.1320 2.4680 0.1640 ;
    LAYER V1 ;
      RECT 2.4160 0.1960 2.4480 0.2280 ;
    LAYER V2 ;
      RECT 2.4160 0.1960 2.4480 0.2280 ;
    LAYER M2 ;
      RECT 0.0280 0.1960 2.4680 0.2280 ;
    LAYER V1 ;
      RECT 0.0480 0.2600 0.0800 0.2920 ;
    LAYER V2 ;
      RECT 0.0480 0.2600 0.0800 0.2920 ;
    LAYER M2 ;
      RECT 0.0280 0.2600 2.4680 0.2920 ;
    LAYER V1 ;
      RECT 2.4160 0.3240 2.4480 0.3560 ;
    LAYER V2 ;
      RECT 2.4160 0.3240 2.4480 0.3560 ;
    LAYER M2 ;
      RECT 0.0280 0.3240 2.4680 0.3560 ;
    LAYER V1 ;
      RECT 0.0480 0.3880 0.0800 0.4200 ;
    LAYER V2 ;
      RECT 0.0480 0.3880 0.0800 0.4200 ;
    LAYER M2 ;
      RECT 0.0280 0.3880 2.4680 0.4200 ;
    LAYER V1 ;
      RECT 2.4160 0.4520 2.4480 0.4840 ;
    LAYER V2 ;
      RECT 2.4160 0.4520 2.4480 0.4840 ;
    LAYER M2 ;
      RECT 0.0280 0.4520 2.4680 0.4840 ;
    LAYER V1 ;
      RECT 0.0480 0.5160 0.0800 0.5480 ;
    LAYER V2 ;
      RECT 0.0480 0.5160 0.0800 0.5480 ;
    LAYER M2 ;
      RECT 0.0280 0.5160 2.4680 0.5480 ;
    LAYER V1 ;
      RECT 2.4160 0.5800 2.4480 0.6120 ;
    LAYER V2 ;
      RECT 2.4160 0.5800 2.4480 0.6120 ;
    LAYER M2 ;
      RECT 0.0280 0.5800 2.4680 0.6120 ;
    LAYER V1 ;
      RECT 0.0480 0.6440 0.0800 0.6760 ;
    LAYER V2 ;
      RECT 0.0480 0.6440 0.0800 0.6760 ;
    LAYER M2 ;
      RECT 0.0280 0.6440 2.4680 0.6760 ;
    LAYER V1 ;
      RECT 2.4160 0.7080 2.4480 0.7400 ;
    LAYER V2 ;
      RECT 2.4160 0.7080 2.4480 0.7400 ;
    LAYER M2 ;
      RECT 0.0280 0.7080 2.4680 0.7400 ;
    LAYER V1 ;
      RECT 0.0480 0.7720 0.0800 0.8040 ;
    LAYER V2 ;
      RECT 0.0480 0.7720 0.0800 0.8040 ;
    LAYER M2 ;
      RECT 0.0280 0.7720 2.4680 0.8040 ;
    LAYER V1 ;
      RECT 2.4160 0.8360 2.4480 0.8680 ;
    LAYER V2 ;
      RECT 2.4160 0.8360 2.4480 0.8680 ;
    LAYER M2 ;
      RECT 0.0280 0.8360 2.4680 0.8680 ;
    LAYER V1 ;
      RECT 0.0480 0.9000 0.0800 0.9320 ;
    LAYER V2 ;
      RECT 0.0480 0.9000 0.0800 0.9320 ;
    LAYER M2 ;
      RECT 0.0280 0.9000 2.4680 0.9320 ;
    LAYER V1 ;
      RECT 2.4160 0.9640 2.4480 0.9960 ;
    LAYER V2 ;
      RECT 2.4160 0.9640 2.4480 0.9960 ;
    LAYER M2 ;
      RECT 0.0280 0.9640 2.4680 0.9960 ;
    LAYER V1 ;
      RECT 0.0480 1.0280 0.0800 1.0600 ;
    LAYER V2 ;
      RECT 0.0480 1.0280 0.0800 1.0600 ;
    LAYER M2 ;
      RECT 0.0280 1.0280 2.4680 1.0600 ;
    LAYER V1 ;
      RECT 2.4160 1.0920 2.4480 1.1240 ;
    LAYER V2 ;
      RECT 2.4160 1.0920 2.4480 1.1240 ;
    LAYER M2 ;
      RECT 0.0280 1.0920 2.4680 1.1240 ;
    LAYER V1 ;
      RECT 0.0480 1.1560 0.0800 1.1880 ;
    LAYER V2 ;
      RECT 0.0480 1.1560 0.0800 1.1880 ;
    LAYER M2 ;
      RECT 0.0280 1.1560 2.4680 1.1880 ;
    LAYER V1 ;
      RECT 2.4160 1.2200 2.4480 1.2520 ;
    LAYER V2 ;
      RECT 2.4160 1.2200 2.4480 1.2520 ;
    LAYER M2 ;
      RECT 0.0280 1.2200 2.4680 1.2520 ;
    LAYER V1 ;
      RECT 0.0480 1.2840 0.0800 1.3160 ;
    LAYER V2 ;
      RECT 0.0480 1.2840 0.0800 1.3160 ;
    LAYER M2 ;
      RECT 0.0280 1.2840 2.4680 1.3160 ;
    LAYER V1 ;
      RECT 2.4160 1.3480 2.4480 1.3800 ;
    LAYER V2 ;
      RECT 2.4160 1.3480 2.4480 1.3800 ;
    LAYER M2 ;
      RECT 0.0280 1.3480 2.4680 1.3800 ;
    LAYER V1 ;
      RECT 0.0480 1.4120 0.0800 1.4440 ;
    LAYER V2 ;
      RECT 0.0480 1.4120 0.0800 1.4440 ;
    LAYER M2 ;
      RECT 0.0280 1.4120 2.4680 1.4440 ;
    LAYER V1 ;
      RECT 2.4160 1.4760 2.4480 1.5080 ;
    LAYER V2 ;
      RECT 2.4160 1.4760 2.4480 1.5080 ;
    LAYER M2 ;
      RECT 0.0280 1.4760 2.4680 1.5080 ;
    LAYER V1 ;
      RECT 0.0480 1.5400 0.0800 1.5720 ;
    LAYER V2 ;
      RECT 0.0480 1.5400 0.0800 1.5720 ;
    LAYER M2 ;
      RECT 0.0280 1.5400 2.4680 1.5720 ;
    LAYER V1 ;
      RECT 2.4160 1.6040 2.4480 1.6360 ;
    LAYER V2 ;
      RECT 2.4160 1.6040 2.4480 1.6360 ;
    LAYER M2 ;
      RECT 0.0280 1.6040 2.4680 1.6360 ;
    LAYER V1 ;
      RECT 0.0480 1.6680 0.0800 1.7000 ;
    LAYER V2 ;
      RECT 0.0480 1.6680 0.0800 1.7000 ;
    LAYER M2 ;
      RECT 0.0280 1.6680 2.4680 1.7000 ;
    LAYER V1 ;
      RECT 2.4160 1.7320 2.4480 1.7640 ;
    LAYER V2 ;
      RECT 2.4160 1.7320 2.4480 1.7640 ;
    LAYER M2 ;
      RECT 0.0280 1.7320 2.4680 1.7640 ;
    LAYER V1 ;
      RECT 0.0480 1.7960 0.0800 1.8280 ;
    LAYER V2 ;
      RECT 0.0480 1.7960 0.0800 1.8280 ;
    LAYER M2 ;
      RECT 0.0280 1.7960 2.4680 1.8280 ;
    LAYER V1 ;
      RECT 2.4160 1.8600 2.4480 1.8920 ;
    LAYER V2 ;
      RECT 2.4160 1.8600 2.4480 1.8920 ;
    LAYER M2 ;
      RECT 0.0280 1.8600 2.4680 1.8920 ;
    LAYER V1 ;
      RECT 0.0480 1.9240 0.0800 1.9560 ;
    LAYER V2 ;
      RECT 0.0480 1.9240 0.0800 1.9560 ;
    LAYER M2 ;
      RECT 0.0280 1.9240 2.4680 1.9560 ;
    LAYER V1 ;
      RECT 2.4160 1.9880 2.4480 2.0200 ;
    LAYER V2 ;
      RECT 2.4160 1.9880 2.4480 2.0200 ;
    LAYER M2 ;
      RECT 0.0280 1.9880 2.4680 2.0200 ;
    LAYER V1 ;
      RECT 0.0480 2.0520 0.0800 2.0840 ;
    LAYER V2 ;
      RECT 0.0480 2.0520 0.0800 2.0840 ;
    LAYER M2 ;
      RECT 0.0280 2.0520 2.4680 2.0840 ;
    LAYER V1 ;
      RECT 2.4160 2.1160 2.4480 2.1480 ;
    LAYER V2 ;
      RECT 2.4160 2.1160 2.4480 2.1480 ;
    LAYER M2 ;
      RECT 0.0280 2.1160 2.4680 2.1480 ;
    LAYER V1 ;
      RECT 0.0480 2.1800 0.0800 2.2120 ;
    LAYER V2 ;
      RECT 0.0480 2.1800 0.0800 2.2120 ;
    LAYER M2 ;
      RECT 0.0280 2.1800 2.4680 2.2120 ;
    LAYER V1 ;
      RECT 2.4160 2.2440 2.4480 2.2760 ;
    LAYER V2 ;
      RECT 2.4160 2.2440 2.4480 2.2760 ;
    LAYER M2 ;
      RECT 0.0280 2.2440 2.4680 2.2760 ;
    LAYER V1 ;
      RECT 0.0480 2.3080 0.0800 2.3400 ;
    LAYER V2 ;
      RECT 0.0480 2.3080 0.0800 2.3400 ;
    LAYER M2 ;
      RECT 0.0280 2.3080 2.4680 2.3400 ;
    LAYER V1 ;
      RECT 2.4160 2.3720 2.4480 2.4040 ;
    LAYER V2 ;
      RECT 2.4160 2.3720 2.4480 2.4040 ;
    LAYER M2 ;
      RECT 0.0280 2.3720 2.4680 2.4040 ;
    LAYER boundary ;
      RECT 0.0000 0.0000 2.4960 2.6040 ;
  END
END cap_12f
MACRO CMC_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2780 1.5560 0.3100 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3620 1.7160 0.3940 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4460 2.2760 0.4780 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V1 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V1 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V1 ;
      RECT 0.3040 0.4460 0.3360 0.4780 ;
    LAYER V1 ;
      RECT 2.2240 0.4460 2.2560 0.4780 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END CMC_NMOS_n12_X2_Y1
MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2780 1.5560 0.3100 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3620 1.7160 0.3940 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4460 2.2760 0.4780 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V1 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V1 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V1 ;
      RECT 0.3040 0.4460 0.3360 0.4780 ;
    LAYER V1 ;
      RECT 2.2240 0.4460 2.2560 0.4780 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END CMC_PMOS_n12_X2_Y1
MACRO CMC_PMOS_S_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 2.2760 0.3940 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 2.2240 0.3620 2.2560 0.3940 ;
    LAYER V1 ;
      RECT 0.9440 0.3620 0.9760 0.3940 ;
    LAYER V1 ;
      RECT 1.5840 0.3620 1.6160 0.3940 ;
  END
END CMC_PMOS_S_n12_X2_Y1
MACRO CMFB_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMFB_NMOS_n12_X2_Y1 0 0 ;
  SIZE 3.8400 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 3.4760 0.1420 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.5640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.2780 3.6360 0.3100 ;
    END
  END DB
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 3.5560 0.3940 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 2.8640 0.0900 2.8960 0.7500 ;
    LAYER M1 ;
      RECT 3.5040 0.0900 3.5360 0.7500 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 2.7840 0.0900 2.8160 0.7500 ;
    LAYER V0 ;
      RECT 2.7840 0.2780 2.8160 0.3100 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER M1 ;
      RECT 3.4240 0.0900 3.4560 0.7500 ;
    LAYER V0 ;
      RECT 3.4240 0.2780 3.4560 0.3100 ;
    LAYER V0 ;
      RECT 3.4240 0.4040 3.4560 0.4360 ;
    LAYER V0 ;
      RECT 3.4240 0.5300 3.4560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 2.9440 0.0900 2.9760 0.7500 ;
    LAYER V0 ;
      RECT 2.9440 0.2780 2.9760 0.3100 ;
    LAYER V0 ;
      RECT 2.9440 0.4040 2.9760 0.4360 ;
    LAYER V0 ;
      RECT 2.9440 0.5300 2.9760 0.5620 ;
    LAYER M1 ;
      RECT 3.5840 0.0900 3.6160 0.7500 ;
    LAYER V0 ;
      RECT 3.5840 0.2780 3.6160 0.3100 ;
    LAYER V0 ;
      RECT 3.5840 0.4040 3.6160 0.4360 ;
    LAYER V0 ;
      RECT 3.5840 0.5300 3.6160 0.5620 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 2.7840 0.1100 2.8160 0.1420 ;
    LAYER V1 ;
      RECT 3.4240 0.1100 3.4560 0.1420 ;
    LAYER V1 ;
      RECT 1.6640 0.1940 1.6960 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 1.5840 0.1940 1.6160 0.2260 ;
    LAYER V1 ;
      RECT 2.2240 0.1940 2.2560 0.2260 ;
    LAYER V1 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 2.9440 0.2780 2.9760 0.3100 ;
    LAYER V1 ;
      RECT 3.5840 0.2780 3.6160 0.3100 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 0.9440 0.3620 0.9760 0.3940 ;
    LAYER V1 ;
      RECT 2.8640 0.3620 2.8960 0.3940 ;
    LAYER V1 ;
      RECT 3.5040 0.3620 3.5360 0.3940 ;
  END
END CMFB_NMOS_n12_X2_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3040 0.1940 0.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.9440 0.1940 0.9760 0.2260 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DP_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 2.2760 0.3940 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4460 1.6360 0.4780 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 2.2240 0.3620 2.2560 0.3940 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END DP_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2780 0.9960 0.3100 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
    LAYER V1 ;
      RECT 0.3040 0.2780 0.3360 0.3100 ;
    LAYER V1 ;
      RECT 0.9440 0.2780 0.9760 0.3100 ;
  END
END Switch_NMOS_n12_X2_Y1
MACRO Switch_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2780 0.9960 0.3100 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
    LAYER V1 ;
      RECT 0.3040 0.2780 0.3360 0.3100 ;
    LAYER V1 ;
      RECT 0.9440 0.2780 0.9760 0.3100 ;
  END
END Switch_PMOS_n12_X2_Y1
MACRO CMC_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2780 1.5560 0.3100 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3620 1.7160 0.3940 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4460 2.2760 0.4780 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V1 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V1 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V1 ;
      RECT 0.3040 0.4460 0.3360 0.4780 ;
    LAYER V1 ;
      RECT 2.2240 0.4460 2.2560 0.4780 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END CMC_NMOS_n12_X2_Y1
MACRO CMC_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2780 1.5560 0.3100 ;
    END
  END SB
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3620 1.7160 0.3940 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4460 2.2760 0.4780 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V1 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V1 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V1 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V1 ;
      RECT 0.3040 0.4460 0.3360 0.4780 ;
    LAYER V1 ;
      RECT 2.2240 0.4460 2.2560 0.4780 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END CMC_PMOS_n12_X2_Y1
MACRO CMC_PMOS_S_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_S_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 2.2760 0.3940 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 2.2240 0.3620 2.2560 0.3940 ;
    LAYER V1 ;
      RECT 0.9440 0.3620 0.9760 0.3940 ;
    LAYER V1 ;
      RECT 1.5840 0.3620 1.6160 0.3940 ;
  END
END CMC_PMOS_S_n12_X2_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3040 0.1940 0.3360 0.2260 ;
    LAYER V1 ;
      RECT 0.9440 0.1940 0.9760 0.2260 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DP_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 2.1960 0.1420 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 2.3560 0.2260 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2780 1.7160 0.3100 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3620 2.2760 0.3940 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4460 1.6360 0.4780 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 2.2240 0.0900 2.2560 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 1.5840 0.0900 1.6160 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 2.1440 0.0900 2.1760 0.7500 ;
    LAYER V0 ;
      RECT 2.1440 0.2780 2.1760 0.3100 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 1.5040 0.0900 1.5360 0.7500 ;
    LAYER V0 ;
      RECT 1.5040 0.2780 1.5360 0.3100 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 2.3040 0.0900 2.3360 0.7500 ;
    LAYER V0 ;
      RECT 2.3040 0.2780 2.3360 0.3100 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER M1 ;
      RECT 1.6640 0.0900 1.6960 0.7500 ;
    LAYER V0 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 2.1440 0.1100 2.1760 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 1.5040 0.1100 1.5360 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 2.3040 0.1940 2.3360 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V1 ;
      RECT 1.6640 0.2780 1.6960 0.3100 ;
    LAYER V1 ;
      RECT 0.3040 0.3620 0.3360 0.3940 ;
    LAYER V1 ;
      RECT 2.2240 0.3620 2.2560 0.3940 ;
    LAYER V1 ;
      RECT 0.9440 0.4460 0.9760 0.4780 ;
    LAYER V1 ;
      RECT 1.5840 0.4460 1.6160 0.4780 ;
  END
END DP_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2780 0.9960 0.3100 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
    LAYER V1 ;
      RECT 0.3040 0.2780 0.3360 0.3100 ;
    LAYER V1 ;
      RECT 0.9440 0.2780 0.9760 0.3100 ;
  END
END Switch_NMOS_n12_X2_Y1
MACRO Switch_PMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 0.9240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.1100 0.9160 0.1420 ;
    END
  END S
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2780 0.9960 0.3100 ;
    END
  END G
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1940 1.0760 0.2260 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0900 0.3360 0.7500 ;
    LAYER M1 ;
      RECT 0.9440 0.0900 0.9760 0.7500 ;
    LAYER M1 ;
      RECT 0.2240 0.0900 0.2560 0.7500 ;
    LAYER V0 ;
      RECT 0.2240 0.2780 0.2560 0.3100 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER M1 ;
      RECT 0.8640 0.0900 0.8960 0.7500 ;
    LAYER V0 ;
      RECT 0.8640 0.2780 0.8960 0.3100 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER M1 ;
      RECT 0.3840 0.0900 0.4160 0.7500 ;
    LAYER V0 ;
      RECT 0.3840 0.2780 0.4160 0.3100 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER M1 ;
      RECT 1.0240 0.0900 1.0560 0.7500 ;
    LAYER V0 ;
      RECT 1.0240 0.2780 1.0560 0.3100 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V1 ;
      RECT 0.2240 0.1100 0.2560 0.1420 ;
    LAYER V1 ;
      RECT 0.8640 0.1100 0.8960 0.1420 ;
    LAYER V1 ;
      RECT 0.3840 0.1940 0.4160 0.2260 ;
    LAYER V1 ;
      RECT 1.0240 0.1940 1.0560 0.2260 ;
    LAYER V1 ;
      RECT 0.3040 0.2780 0.3360 0.3100 ;
    LAYER V1 ;
      RECT 0.9440 0.2780 0.9760 0.3100 ;
  END
END Switch_PMOS_n12_X2_Y1
