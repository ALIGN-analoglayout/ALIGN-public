.subckt cap_pair vip vin vop von vss vdd
c0 vip vop 30e-15
c1 vin von 60e-15
.ends cap_pair
