MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 10.24 BY 26.208 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.68 25.752 3.712 25.824 ;
      LAYER M2 ;
        RECT 3.66 25.772 3.732 25.804 ;
      LAYER M1 ;
        RECT 6.976 25.752 7.008 25.824 ;
      LAYER M2 ;
        RECT 6.956 25.772 7.028 25.804 ;
      LAYER M2 ;
        RECT 3.696 25.772 6.992 25.804 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
      LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
      LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
      LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
      LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.84 25.92 3.872 25.992 ;
      LAYER M2 ;
        RECT 3.82 25.94 3.892 25.972 ;
      LAYER M1 ;
        RECT 7.136 25.92 7.168 25.992 ;
      LAYER M2 ;
        RECT 7.116 25.94 7.188 25.972 ;
      LAYER M2 ;
        RECT 3.856 25.94 7.152 25.972 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
      LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
      LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
      LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
      LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M2 ;
        RECT 3.376 13.424 6.448 13.456 ;
  LAYER M1 ;
        RECT 3.36 13.404 3.392 13.476 ;
  LAYER M2 ;
        RECT 3.34 13.424 3.412 13.456 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M2 ;
        RECT 3.376 7.208 6.448 7.24 ;
  LAYER M1 ;
        RECT 3.36 7.188 3.392 7.26 ;
  LAYER M2 ;
        RECT 3.34 7.208 3.412 7.24 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M2 ;
        RECT 3.376 16.532 6.448 16.564 ;
  LAYER M1 ;
        RECT 3.36 16.512 3.392 16.584 ;
  LAYER M2 ;
        RECT 3.34 16.532 3.412 16.564 ;
  LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
  LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
  LAYER M1 ;
        RECT 3.36 0.42 3.392 0.672 ;
  LAYER M1 ;
        RECT 3.36 0.672 3.392 16.548 ;
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M1 ;
        RECT 6.432 13.272 6.464 13.44 ;
  LAYER M1 ;
        RECT 6.432 13.236 6.464 13.308 ;
  LAYER M2 ;
        RECT 6.412 13.256 6.484 13.288 ;
  LAYER M2 ;
        RECT 6.448 13.256 6.672 13.288 ;
  LAYER M1 ;
        RECT 6.656 13.236 6.688 13.308 ;
  LAYER M2 ;
        RECT 6.636 13.256 6.708 13.288 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M1 ;
        RECT 6.432 7.056 6.464 7.224 ;
  LAYER M1 ;
        RECT 6.432 7.02 6.464 7.092 ;
  LAYER M2 ;
        RECT 6.412 7.04 6.484 7.072 ;
  LAYER M2 ;
        RECT 6.448 7.04 6.672 7.072 ;
  LAYER M1 ;
        RECT 6.656 7.02 6.688 7.092 ;
  LAYER M2 ;
        RECT 6.636 7.04 6.708 7.072 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M1 ;
        RECT 6.432 16.38 6.464 16.548 ;
  LAYER M1 ;
        RECT 6.432 16.344 6.464 16.416 ;
  LAYER M2 ;
        RECT 6.412 16.364 6.484 16.396 ;
  LAYER M2 ;
        RECT 6.448 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 16.416 ;
  LAYER M2 ;
        RECT 6.636 16.364 6.708 16.396 ;
  LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
  LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
  LAYER M1 ;
        RECT 6.656 0.42 6.688 0.672 ;
  LAYER M1 ;
        RECT 6.656 0.672 6.688 16.38 ;
  LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M2 ;
        RECT 3.536 10.316 6.448 10.348 ;
  LAYER M1 ;
        RECT 3.52 10.296 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.5 10.316 3.572 10.348 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M2 ;
        RECT 3.536 4.1 6.448 4.132 ;
  LAYER M1 ;
        RECT 3.52 4.08 3.552 4.152 ;
  LAYER M2 ;
        RECT 3.5 4.1 3.572 4.132 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M2 ;
        RECT 3.536 19.64 6.448 19.672 ;
  LAYER M1 ;
        RECT 3.52 19.62 3.552 19.692 ;
  LAYER M2 ;
        RECT 3.5 19.64 3.572 19.672 ;
  LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
  LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
  LAYER M1 ;
        RECT 3.52 0.252 3.552 0.672 ;
  LAYER M1 ;
        RECT 3.52 0.672 3.552 19.656 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M1 ;
        RECT 6.432 10.164 6.464 10.332 ;
  LAYER M1 ;
        RECT 6.432 10.128 6.464 10.2 ;
  LAYER M2 ;
        RECT 6.412 10.148 6.484 10.18 ;
  LAYER M2 ;
        RECT 6.448 10.148 6.832 10.18 ;
  LAYER M1 ;
        RECT 6.816 10.128 6.848 10.2 ;
  LAYER M2 ;
        RECT 6.796 10.148 6.868 10.18 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M1 ;
        RECT 6.432 3.948 6.464 4.116 ;
  LAYER M1 ;
        RECT 6.432 3.912 6.464 3.984 ;
  LAYER M2 ;
        RECT 6.412 3.932 6.484 3.964 ;
  LAYER M2 ;
        RECT 6.448 3.932 6.832 3.964 ;
  LAYER M1 ;
        RECT 6.816 3.912 6.848 3.984 ;
  LAYER M2 ;
        RECT 6.796 3.932 6.868 3.964 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M1 ;
        RECT 6.432 19.488 6.464 19.656 ;
  LAYER M1 ;
        RECT 6.432 19.452 6.464 19.524 ;
  LAYER M2 ;
        RECT 6.412 19.472 6.484 19.504 ;
  LAYER M2 ;
        RECT 6.448 19.472 6.832 19.504 ;
  LAYER M1 ;
        RECT 6.816 19.452 6.848 19.524 ;
  LAYER M2 ;
        RECT 6.796 19.472 6.868 19.504 ;
  LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
  LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
  LAYER M1 ;
        RECT 6.816 0.252 6.848 0.672 ;
  LAYER M1 ;
        RECT 6.816 0.672 6.848 19.488 ;
  LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 3.152 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 3.136 4.08 3.168 4.152 ;
  LAYER M2 ;
        RECT 3.116 4.1 3.188 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 3.152 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 3.136 7.188 3.168 7.26 ;
  LAYER M2 ;
        RECT 3.116 7.208 3.188 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 3.152 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 3.136 10.296 3.168 10.368 ;
  LAYER M2 ;
        RECT 3.116 10.316 3.188 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 3.152 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 3.136 13.404 3.168 13.476 ;
  LAYER M2 ;
        RECT 3.116 13.424 3.188 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 3.152 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 3.136 16.512 3.168 16.584 ;
  LAYER M2 ;
        RECT 3.116 16.532 3.188 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 3.152 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 3.136 19.62 3.168 19.692 ;
  LAYER M2 ;
        RECT 3.116 19.64 3.188 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 3.152 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 22.8 ;
  LAYER M2 ;
        RECT 3.116 22.748 3.188 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 3.152 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 22.764 ;
  LAYER M1 ;
        RECT 9.728 0.972 9.76 1.044 ;
  LAYER M2 ;
        RECT 9.708 0.992 9.78 1.024 ;
  LAYER M1 ;
        RECT 9.728 0.84 9.76 1.008 ;
  LAYER M1 ;
        RECT 9.728 0.804 9.76 0.876 ;
  LAYER M2 ;
        RECT 9.708 0.824 9.78 0.856 ;
  LAYER M2 ;
        RECT 9.744 0.824 9.968 0.856 ;
  LAYER M1 ;
        RECT 9.952 0.804 9.984 0.876 ;
  LAYER M2 ;
        RECT 9.932 0.824 10.004 0.856 ;
  LAYER M1 ;
        RECT 9.728 4.08 9.76 4.152 ;
  LAYER M2 ;
        RECT 9.708 4.1 9.78 4.132 ;
  LAYER M1 ;
        RECT 9.728 3.948 9.76 4.116 ;
  LAYER M1 ;
        RECT 9.728 3.912 9.76 3.984 ;
  LAYER M2 ;
        RECT 9.708 3.932 9.78 3.964 ;
  LAYER M2 ;
        RECT 9.744 3.932 9.968 3.964 ;
  LAYER M1 ;
        RECT 9.952 3.912 9.984 3.984 ;
  LAYER M2 ;
        RECT 9.932 3.932 10.004 3.964 ;
  LAYER M1 ;
        RECT 9.728 7.188 9.76 7.26 ;
  LAYER M2 ;
        RECT 9.708 7.208 9.78 7.24 ;
  LAYER M1 ;
        RECT 9.728 7.056 9.76 7.224 ;
  LAYER M1 ;
        RECT 9.728 7.02 9.76 7.092 ;
  LAYER M2 ;
        RECT 9.708 7.04 9.78 7.072 ;
  LAYER M2 ;
        RECT 9.744 7.04 9.968 7.072 ;
  LAYER M1 ;
        RECT 9.952 7.02 9.984 7.092 ;
  LAYER M2 ;
        RECT 9.932 7.04 10.004 7.072 ;
  LAYER M1 ;
        RECT 9.728 10.296 9.76 10.368 ;
  LAYER M2 ;
        RECT 9.708 10.316 9.78 10.348 ;
  LAYER M1 ;
        RECT 9.728 10.164 9.76 10.332 ;
  LAYER M1 ;
        RECT 9.728 10.128 9.76 10.2 ;
  LAYER M2 ;
        RECT 9.708 10.148 9.78 10.18 ;
  LAYER M2 ;
        RECT 9.744 10.148 9.968 10.18 ;
  LAYER M1 ;
        RECT 9.952 10.128 9.984 10.2 ;
  LAYER M2 ;
        RECT 9.932 10.148 10.004 10.18 ;
  LAYER M1 ;
        RECT 9.728 13.404 9.76 13.476 ;
  LAYER M2 ;
        RECT 9.708 13.424 9.78 13.456 ;
  LAYER M1 ;
        RECT 9.728 13.272 9.76 13.44 ;
  LAYER M1 ;
        RECT 9.728 13.236 9.76 13.308 ;
  LAYER M2 ;
        RECT 9.708 13.256 9.78 13.288 ;
  LAYER M2 ;
        RECT 9.744 13.256 9.968 13.288 ;
  LAYER M1 ;
        RECT 9.952 13.236 9.984 13.308 ;
  LAYER M2 ;
        RECT 9.932 13.256 10.004 13.288 ;
  LAYER M1 ;
        RECT 9.728 16.512 9.76 16.584 ;
  LAYER M2 ;
        RECT 9.708 16.532 9.78 16.564 ;
  LAYER M1 ;
        RECT 9.728 16.38 9.76 16.548 ;
  LAYER M1 ;
        RECT 9.728 16.344 9.76 16.416 ;
  LAYER M2 ;
        RECT 9.708 16.364 9.78 16.396 ;
  LAYER M2 ;
        RECT 9.744 16.364 9.968 16.396 ;
  LAYER M1 ;
        RECT 9.952 16.344 9.984 16.416 ;
  LAYER M2 ;
        RECT 9.932 16.364 10.004 16.396 ;
  LAYER M1 ;
        RECT 9.728 19.62 9.76 19.692 ;
  LAYER M2 ;
        RECT 9.708 19.64 9.78 19.672 ;
  LAYER M1 ;
        RECT 9.728 19.488 9.76 19.656 ;
  LAYER M1 ;
        RECT 9.728 19.452 9.76 19.524 ;
  LAYER M2 ;
        RECT 9.708 19.472 9.78 19.504 ;
  LAYER M2 ;
        RECT 9.744 19.472 9.968 19.504 ;
  LAYER M1 ;
        RECT 9.952 19.452 9.984 19.524 ;
  LAYER M2 ;
        RECT 9.932 19.472 10.004 19.504 ;
  LAYER M1 ;
        RECT 9.728 22.728 9.76 22.8 ;
  LAYER M2 ;
        RECT 9.708 22.748 9.78 22.78 ;
  LAYER M1 ;
        RECT 9.728 22.596 9.76 22.764 ;
  LAYER M1 ;
        RECT 9.728 22.56 9.76 22.632 ;
  LAYER M2 ;
        RECT 9.708 22.58 9.78 22.612 ;
  LAYER M2 ;
        RECT 9.744 22.58 9.968 22.612 ;
  LAYER M1 ;
        RECT 9.952 22.56 9.984 22.632 ;
  LAYER M2 ;
        RECT 9.932 22.58 10.004 22.612 ;
  LAYER M1 ;
        RECT 9.952 0.048 9.984 0.12 ;
  LAYER M2 ;
        RECT 9.932 0.068 10.004 0.1 ;
  LAYER M1 ;
        RECT 9.952 0.084 9.984 0.672 ;
  LAYER M1 ;
        RECT 9.952 0.672 9.984 22.596 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.968 0.1 ;
  LAYER M1 ;
        RECT 6.432 0.972 6.464 1.044 ;
  LAYER M2 ;
        RECT 6.412 0.992 6.484 1.024 ;
  LAYER M2 ;
        RECT 3.152 0.992 6.448 1.024 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M1 ;
        RECT 6.432 22.728 6.464 22.8 ;
  LAYER M2 ;
        RECT 6.412 22.748 6.484 22.78 ;
  LAYER M2 ;
        RECT 3.152 22.748 6.448 22.78 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 22.8 ;
  LAYER M2 ;
        RECT 3.116 22.748 3.188 22.78 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M2 ;
        RECT 3.696 15.86 4.08 15.892 ;
  LAYER M1 ;
        RECT 3.68 15.84 3.712 15.912 ;
  LAYER M2 ;
        RECT 3.66 15.86 3.732 15.892 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M2 ;
        RECT 3.696 9.644 4.08 9.676 ;
  LAYER M1 ;
        RECT 3.68 9.624 3.712 9.696 ;
  LAYER M2 ;
        RECT 3.66 9.644 3.732 9.676 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M2 ;
        RECT 3.696 18.968 4.08 19 ;
  LAYER M1 ;
        RECT 3.68 18.948 3.712 19.02 ;
  LAYER M2 ;
        RECT 3.66 18.968 3.732 19 ;
  LAYER M1 ;
        RECT 3.68 25.752 3.712 25.824 ;
  LAYER M2 ;
        RECT 3.66 25.772 3.732 25.804 ;
  LAYER M1 ;
        RECT 3.68 25.536 3.712 25.788 ;
  LAYER M1 ;
        RECT 3.68 9.66 3.712 25.536 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M1 ;
        RECT 4.064 15.876 4.096 16.044 ;
  LAYER M1 ;
        RECT 4.064 16.008 4.096 16.08 ;
  LAYER M2 ;
        RECT 4.044 16.028 4.116 16.06 ;
  LAYER M2 ;
        RECT 4.08 16.028 6.992 16.06 ;
  LAYER M1 ;
        RECT 6.976 16.008 7.008 16.08 ;
  LAYER M2 ;
        RECT 6.956 16.028 7.028 16.06 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M1 ;
        RECT 4.064 9.66 4.096 9.828 ;
  LAYER M1 ;
        RECT 4.064 9.792 4.096 9.864 ;
  LAYER M2 ;
        RECT 4.044 9.812 4.116 9.844 ;
  LAYER M2 ;
        RECT 4.08 9.812 6.992 9.844 ;
  LAYER M1 ;
        RECT 6.976 9.792 7.008 9.864 ;
  LAYER M2 ;
        RECT 6.956 9.812 7.028 9.844 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M1 ;
        RECT 4.064 18.984 4.096 19.152 ;
  LAYER M1 ;
        RECT 4.064 19.116 4.096 19.188 ;
  LAYER M2 ;
        RECT 4.044 19.136 4.116 19.168 ;
  LAYER M2 ;
        RECT 4.08 19.136 6.992 19.168 ;
  LAYER M1 ;
        RECT 6.976 19.116 7.008 19.188 ;
  LAYER M2 ;
        RECT 6.956 19.136 7.028 19.168 ;
  LAYER M1 ;
        RECT 6.976 25.752 7.008 25.824 ;
  LAYER M2 ;
        RECT 6.956 25.772 7.028 25.804 ;
  LAYER M1 ;
        RECT 6.976 25.536 7.008 25.788 ;
  LAYER M1 ;
        RECT 6.976 9.828 7.008 25.536 ;
  LAYER M2 ;
        RECT 3.696 25.772 6.992 25.804 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M2 ;
        RECT 3.856 12.752 4.08 12.784 ;
  LAYER M1 ;
        RECT 3.84 12.732 3.872 12.804 ;
  LAYER M2 ;
        RECT 3.82 12.752 3.892 12.784 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M2 ;
        RECT 3.856 6.536 4.08 6.568 ;
  LAYER M1 ;
        RECT 3.84 6.516 3.872 6.588 ;
  LAYER M2 ;
        RECT 3.82 6.536 3.892 6.568 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M2 ;
        RECT 3.856 22.076 4.08 22.108 ;
  LAYER M1 ;
        RECT 3.84 22.056 3.872 22.128 ;
  LAYER M2 ;
        RECT 3.82 22.076 3.892 22.108 ;
  LAYER M1 ;
        RECT 3.84 25.92 3.872 25.992 ;
  LAYER M2 ;
        RECT 3.82 25.94 3.892 25.972 ;
  LAYER M1 ;
        RECT 3.84 25.536 3.872 25.956 ;
  LAYER M1 ;
        RECT 3.84 6.552 3.872 25.536 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M1 ;
        RECT 4.064 12.768 4.096 12.936 ;
  LAYER M1 ;
        RECT 4.064 12.9 4.096 12.972 ;
  LAYER M2 ;
        RECT 4.044 12.92 4.116 12.952 ;
  LAYER M2 ;
        RECT 4.08 12.92 7.152 12.952 ;
  LAYER M1 ;
        RECT 7.136 12.9 7.168 12.972 ;
  LAYER M2 ;
        RECT 7.116 12.92 7.188 12.952 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M1 ;
        RECT 4.064 6.552 4.096 6.72 ;
  LAYER M1 ;
        RECT 4.064 6.684 4.096 6.756 ;
  LAYER M2 ;
        RECT 4.044 6.704 4.116 6.736 ;
  LAYER M2 ;
        RECT 4.08 6.704 7.152 6.736 ;
  LAYER M1 ;
        RECT 7.136 6.684 7.168 6.756 ;
  LAYER M2 ;
        RECT 7.116 6.704 7.188 6.736 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M1 ;
        RECT 4.064 22.092 4.096 22.26 ;
  LAYER M1 ;
        RECT 4.064 22.224 4.096 22.296 ;
  LAYER M2 ;
        RECT 4.044 22.244 4.116 22.276 ;
  LAYER M2 ;
        RECT 4.08 22.244 7.152 22.276 ;
  LAYER M1 ;
        RECT 7.136 22.224 7.168 22.296 ;
  LAYER M2 ;
        RECT 7.116 22.244 7.188 22.276 ;
  LAYER M1 ;
        RECT 7.136 25.92 7.168 25.992 ;
  LAYER M2 ;
        RECT 7.116 25.94 7.188 25.972 ;
  LAYER M1 ;
        RECT 7.136 25.536 7.168 25.956 ;
  LAYER M1 ;
        RECT 7.136 6.72 7.168 25.536 ;
  LAYER M2 ;
        RECT 3.856 25.94 7.152 25.972 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.784 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.768 6.516 0.8 6.588 ;
  LAYER M2 ;
        RECT 0.748 6.536 0.82 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.784 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.768 9.624 0.8 9.696 ;
  LAYER M2 ;
        RECT 0.748 9.644 0.82 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.784 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.768 12.732 0.8 12.804 ;
  LAYER M2 ;
        RECT 0.748 12.752 0.82 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.784 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.768 15.84 0.8 15.912 ;
  LAYER M2 ;
        RECT 0.748 15.86 0.82 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.784 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.768 18.948 0.8 19.02 ;
  LAYER M2 ;
        RECT 0.748 18.968 0.82 19 ;
  LAYER M2 ;
        RECT 0.24 18.968 0.784 19 ;
  LAYER M1 ;
        RECT 0.224 18.948 0.256 19.02 ;
  LAYER M2 ;
        RECT 0.204 18.968 0.276 19 ;
  LAYER M1 ;
        RECT 0.768 22.056 0.8 22.128 ;
  LAYER M2 ;
        RECT 0.748 22.076 0.82 22.108 ;
  LAYER M2 ;
        RECT 0.24 22.076 0.784 22.108 ;
  LAYER M1 ;
        RECT 0.224 22.056 0.256 22.128 ;
  LAYER M2 ;
        RECT 0.204 22.076 0.276 22.108 ;
  LAYER M1 ;
        RECT 0.768 25.164 0.8 25.236 ;
  LAYER M2 ;
        RECT 0.748 25.184 0.82 25.216 ;
  LAYER M2 ;
        RECT 0.24 25.184 0.784 25.216 ;
  LAYER M1 ;
        RECT 0.224 25.164 0.256 25.236 ;
  LAYER M2 ;
        RECT 0.204 25.184 0.276 25.216 ;
  LAYER M1 ;
        RECT 0.224 26.088 0.256 26.16 ;
  LAYER M2 ;
        RECT 0.204 26.108 0.276 26.14 ;
  LAYER M1 ;
        RECT 0.224 25.536 0.256 26.124 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 25.536 ;
  LAYER M1 ;
        RECT 7.36 3.408 7.392 3.48 ;
  LAYER M2 ;
        RECT 7.34 3.428 7.412 3.46 ;
  LAYER M1 ;
        RECT 7.376 3.428 10.128 3.46 ;
  LAYER M1 ;
        RECT 10.112 3.408 10.144 3.48 ;
  LAYER M2 ;
        RECT 10.092 3.428 10.164 3.46 ;
  LAYER M2 ;
        RECT 10.128 3.428 10.192 3.46 ;
  LAYER M1 ;
        RECT 10.176 3.408 10.208 3.48 ;
  LAYER M2 ;
        RECT 10.156 3.428 10.228 3.46 ;
  LAYER M1 ;
        RECT 7.36 6.516 7.392 6.588 ;
  LAYER M2 ;
        RECT 7.34 6.536 7.412 6.568 ;
  LAYER M1 ;
        RECT 7.376 6.536 10.128 6.568 ;
  LAYER M1 ;
        RECT 10.112 6.516 10.144 6.588 ;
  LAYER M2 ;
        RECT 10.092 6.536 10.164 6.568 ;
  LAYER M2 ;
        RECT 10.128 6.536 10.192 6.568 ;
  LAYER M1 ;
        RECT 10.176 6.516 10.208 6.588 ;
  LAYER M2 ;
        RECT 10.156 6.536 10.228 6.568 ;
  LAYER M1 ;
        RECT 7.36 9.624 7.392 9.696 ;
  LAYER M2 ;
        RECT 7.34 9.644 7.412 9.676 ;
  LAYER M1 ;
        RECT 7.376 9.644 10.128 9.676 ;
  LAYER M1 ;
        RECT 10.112 9.624 10.144 9.696 ;
  LAYER M2 ;
        RECT 10.092 9.644 10.164 9.676 ;
  LAYER M2 ;
        RECT 10.128 9.644 10.192 9.676 ;
  LAYER M1 ;
        RECT 10.176 9.624 10.208 9.696 ;
  LAYER M2 ;
        RECT 10.156 9.644 10.228 9.676 ;
  LAYER M1 ;
        RECT 7.36 12.732 7.392 12.804 ;
  LAYER M2 ;
        RECT 7.34 12.752 7.412 12.784 ;
  LAYER M1 ;
        RECT 7.376 12.752 10.128 12.784 ;
  LAYER M1 ;
        RECT 10.112 12.732 10.144 12.804 ;
  LAYER M2 ;
        RECT 10.092 12.752 10.164 12.784 ;
  LAYER M2 ;
        RECT 10.128 12.752 10.192 12.784 ;
  LAYER M1 ;
        RECT 10.176 12.732 10.208 12.804 ;
  LAYER M2 ;
        RECT 10.156 12.752 10.228 12.784 ;
  LAYER M1 ;
        RECT 7.36 15.84 7.392 15.912 ;
  LAYER M2 ;
        RECT 7.34 15.86 7.412 15.892 ;
  LAYER M1 ;
        RECT 7.376 15.86 10.128 15.892 ;
  LAYER M1 ;
        RECT 10.112 15.84 10.144 15.912 ;
  LAYER M2 ;
        RECT 10.092 15.86 10.164 15.892 ;
  LAYER M2 ;
        RECT 10.128 15.86 10.192 15.892 ;
  LAYER M1 ;
        RECT 10.176 15.84 10.208 15.912 ;
  LAYER M2 ;
        RECT 10.156 15.86 10.228 15.892 ;
  LAYER M1 ;
        RECT 7.36 18.948 7.392 19.02 ;
  LAYER M2 ;
        RECT 7.34 18.968 7.412 19 ;
  LAYER M1 ;
        RECT 7.376 18.968 10.128 19 ;
  LAYER M1 ;
        RECT 10.112 18.948 10.144 19.02 ;
  LAYER M2 ;
        RECT 10.092 18.968 10.164 19 ;
  LAYER M2 ;
        RECT 10.128 18.968 10.192 19 ;
  LAYER M1 ;
        RECT 10.176 18.948 10.208 19.02 ;
  LAYER M2 ;
        RECT 10.156 18.968 10.228 19 ;
  LAYER M1 ;
        RECT 7.36 22.056 7.392 22.128 ;
  LAYER M2 ;
        RECT 7.34 22.076 7.412 22.108 ;
  LAYER M1 ;
        RECT 7.376 22.076 10.128 22.108 ;
  LAYER M1 ;
        RECT 10.112 22.056 10.144 22.128 ;
  LAYER M2 ;
        RECT 10.092 22.076 10.164 22.108 ;
  LAYER M2 ;
        RECT 10.128 22.076 10.192 22.108 ;
  LAYER M1 ;
        RECT 10.176 22.056 10.208 22.128 ;
  LAYER M2 ;
        RECT 10.156 22.076 10.228 22.108 ;
  LAYER M1 ;
        RECT 7.36 25.164 7.392 25.236 ;
  LAYER M2 ;
        RECT 7.34 25.184 7.412 25.216 ;
  LAYER M1 ;
        RECT 7.376 25.184 10.128 25.216 ;
  LAYER M1 ;
        RECT 10.112 25.164 10.144 25.236 ;
  LAYER M2 ;
        RECT 10.092 25.184 10.164 25.216 ;
  LAYER M2 ;
        RECT 10.128 25.184 10.192 25.216 ;
  LAYER M1 ;
        RECT 10.176 25.164 10.208 25.236 ;
  LAYER M2 ;
        RECT 10.156 25.184 10.228 25.216 ;
  LAYER M1 ;
        RECT 10.176 26.088 10.208 26.16 ;
  LAYER M2 ;
        RECT 10.156 26.108 10.228 26.14 ;
  LAYER M1 ;
        RECT 10.176 25.536 10.208 26.124 ;
  LAYER M1 ;
        RECT 10.176 3.612 10.208 25.536 ;
  LAYER M2 ;
        RECT 0.24 26.108 10.192 26.14 ;
  LAYER M1 ;
        RECT 4.064 3.408 4.096 3.48 ;
  LAYER M2 ;
        RECT 4.044 3.428 4.116 3.46 ;
  LAYER M2 ;
        RECT 0.784 3.428 4.08 3.46 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M1 ;
        RECT 4.064 25.164 4.096 25.236 ;
  LAYER M2 ;
        RECT 4.044 25.184 4.116 25.216 ;
  LAYER M2 ;
        RECT 0.784 25.184 4.08 25.216 ;
  LAYER M1 ;
        RECT 0.768 25.164 0.8 25.236 ;
  LAYER M2 ;
        RECT 0.748 25.184 0.82 25.216 ;
  LAYER M1 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M3 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M2 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M1 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M3 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M2 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M1 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M3 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M2 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M1 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M3 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M2 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M1 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M3 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M2 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M1 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M3 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M2 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M1 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M3 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M2 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M1 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M3 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M2 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M1 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M3 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M2 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M1 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M3 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M2 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M1 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M3 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M2 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M1 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M3 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M2 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M1 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M3 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M2 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M1 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M3 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M2 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M1 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M3 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M2 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M1 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M3 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M2 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M1 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M3 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M2 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M1 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M3 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M2 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M1 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M3 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M2 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M1 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M3 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M2 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M1 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M3 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M2 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M1 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M3 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M2 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M1 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M3 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M2 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M1 ;
        RECT 7.312 22.68 9.808 25.284 ;
  LAYER M3 ;
        RECT 7.312 22.68 9.808 25.284 ;
  LAYER M2 ;
        RECT 7.312 22.68 9.808 25.284 ;
  END 
END Cap_30fF_Cap_30fF
