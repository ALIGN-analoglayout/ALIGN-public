MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 15.36 BY 21.924 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
      LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
      LAYER M1 ;
        RECT 12.384 21.468 12.416 21.54 ;
      LAYER M2 ;
        RECT 12.364 21.488 12.436 21.52 ;
      LAYER M2 ;
        RECT 2.8 21.488 12.4 21.52 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
      LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
      LAYER M1 ;
        RECT 9.024 0.384 9.056 0.456 ;
      LAYER M2 ;
        RECT 9.004 0.404 9.076 0.436 ;
      LAYER M2 ;
        RECT 5.84 0.404 9.04 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.144 21.636 6.176 21.708 ;
      LAYER M2 ;
        RECT 6.124 21.656 6.196 21.688 ;
      LAYER M1 ;
        RECT 9.344 21.636 9.376 21.708 ;
      LAYER M2 ;
        RECT 9.324 21.656 9.396 21.688 ;
      LAYER M2 ;
        RECT 6.16 21.656 9.36 21.688 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.624 0.216 2.656 0.288 ;
      LAYER M2 ;
        RECT 2.604 0.236 2.676 0.268 ;
      LAYER M1 ;
        RECT 12.224 0.216 12.256 0.288 ;
      LAYER M2 ;
        RECT 12.204 0.236 12.276 0.268 ;
      LAYER M2 ;
        RECT 2.64 0.236 12.24 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.464 6.768 6.496 6.84 ;
  LAYER M2 ;
        RECT 6.444 6.788 6.516 6.82 ;
  LAYER M2 ;
        RECT 5.84 6.788 6.48 6.82 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 6.84 ;
  LAYER M2 ;
        RECT 5.804 6.788 5.876 6.82 ;
  LAYER M1 ;
        RECT 6.464 12.648 6.496 12.72 ;
  LAYER M2 ;
        RECT 6.444 12.668 6.516 12.7 ;
  LAYER M2 ;
        RECT 5.84 12.668 6.48 12.7 ;
  LAYER M1 ;
        RECT 5.824 12.648 5.856 12.72 ;
  LAYER M2 ;
        RECT 5.804 12.668 5.876 12.7 ;
  LAYER M1 ;
        RECT 3.264 9.708 3.296 9.78 ;
  LAYER M2 ;
        RECT 3.244 9.728 3.316 9.76 ;
  LAYER M1 ;
        RECT 3.264 9.576 3.296 9.744 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 9.612 ;
  LAYER M2 ;
        RECT 3.244 9.56 3.316 9.592 ;
  LAYER M2 ;
        RECT 3.28 9.56 5.84 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 3.264 6.768 3.296 6.84 ;
  LAYER M2 ;
        RECT 3.244 6.788 3.316 6.82 ;
  LAYER M1 ;
        RECT 3.264 6.636 3.296 6.804 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 6.672 ;
  LAYER M2 ;
        RECT 3.244 6.62 3.316 6.652 ;
  LAYER M2 ;
        RECT 3.28 6.62 5.84 6.652 ;
  LAYER M1 ;
        RECT 5.824 6.6 5.856 6.672 ;
  LAYER M2 ;
        RECT 5.804 6.62 5.876 6.652 ;
  LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
  LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 0.588 ;
  LAYER M1 ;
        RECT 5.824 0.588 5.856 12.684 ;
  LAYER M1 ;
        RECT 9.664 9.708 9.696 9.78 ;
  LAYER M2 ;
        RECT 9.644 9.728 9.716 9.76 ;
  LAYER M2 ;
        RECT 9.04 9.728 9.68 9.76 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 9.78 ;
  LAYER M2 ;
        RECT 9.004 9.728 9.076 9.76 ;
  LAYER M1 ;
        RECT 9.664 12.648 9.696 12.72 ;
  LAYER M2 ;
        RECT 9.644 12.668 9.716 12.7 ;
  LAYER M2 ;
        RECT 9.04 12.668 9.68 12.7 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 12.72 ;
  LAYER M2 ;
        RECT 9.004 12.668 9.076 12.7 ;
  LAYER M1 ;
        RECT 9.024 0.384 9.056 0.456 ;
  LAYER M2 ;
        RECT 9.004 0.404 9.076 0.436 ;
  LAYER M1 ;
        RECT 9.024 0.42 9.056 0.588 ;
  LAYER M1 ;
        RECT 9.024 0.588 9.056 12.684 ;
  LAYER M2 ;
        RECT 5.84 0.404 9.04 0.436 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 12.72 ;
  LAYER M2 ;
        RECT 3.244 12.668 3.316 12.7 ;
  LAYER M2 ;
        RECT 2.64 12.668 3.28 12.7 ;
  LAYER M1 ;
        RECT 2.624 12.648 2.656 12.72 ;
  LAYER M2 ;
        RECT 2.604 12.668 2.676 12.7 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M2 ;
        RECT 2.64 15.608 3.28 15.64 ;
  LAYER M1 ;
        RECT 2.624 15.588 2.656 15.66 ;
  LAYER M2 ;
        RECT 2.604 15.608 2.676 15.64 ;
  LAYER M1 ;
        RECT 2.624 0.216 2.656 0.288 ;
  LAYER M2 ;
        RECT 2.604 0.236 2.676 0.268 ;
  LAYER M1 ;
        RECT 2.624 0.252 2.656 0.588 ;
  LAYER M1 ;
        RECT 2.624 0.588 2.656 15.624 ;
  LAYER M1 ;
        RECT 9.664 6.768 9.696 6.84 ;
  LAYER M2 ;
        RECT 9.644 6.788 9.716 6.82 ;
  LAYER M1 ;
        RECT 9.664 6.636 9.696 6.804 ;
  LAYER M1 ;
        RECT 9.664 6.6 9.696 6.672 ;
  LAYER M2 ;
        RECT 9.644 6.62 9.716 6.652 ;
  LAYER M2 ;
        RECT 9.68 6.62 12.24 6.652 ;
  LAYER M1 ;
        RECT 12.224 6.6 12.256 6.672 ;
  LAYER M2 ;
        RECT 12.204 6.62 12.276 6.652 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 3.9 ;
  LAYER M2 ;
        RECT 9.644 3.848 9.716 3.88 ;
  LAYER M1 ;
        RECT 9.664 3.696 9.696 3.864 ;
  LAYER M1 ;
        RECT 9.664 3.66 9.696 3.732 ;
  LAYER M2 ;
        RECT 9.644 3.68 9.716 3.712 ;
  LAYER M2 ;
        RECT 9.68 3.68 12.24 3.712 ;
  LAYER M1 ;
        RECT 12.224 3.66 12.256 3.732 ;
  LAYER M2 ;
        RECT 12.204 3.68 12.276 3.712 ;
  LAYER M1 ;
        RECT 12.224 0.216 12.256 0.288 ;
  LAYER M2 ;
        RECT 12.204 0.236 12.276 0.268 ;
  LAYER M1 ;
        RECT 12.224 0.252 12.256 0.588 ;
  LAYER M1 ;
        RECT 12.224 0.588 12.256 6.636 ;
  LAYER M2 ;
        RECT 2.64 0.236 12.24 0.268 ;
  LAYER M1 ;
        RECT 6.464 15.588 6.496 15.66 ;
  LAYER M2 ;
        RECT 6.444 15.608 6.516 15.64 ;
  LAYER M2 ;
        RECT 3.28 15.608 6.48 15.64 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M1 ;
        RECT 6.464 3.828 6.496 3.9 ;
  LAYER M2 ;
        RECT 6.444 3.848 6.516 3.88 ;
  LAYER M2 ;
        RECT 6.48 3.848 9.68 3.88 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 3.9 ;
  LAYER M2 ;
        RECT 9.644 3.848 9.716 3.88 ;
  LAYER M1 ;
        RECT 3.264 0.888 3.296 0.96 ;
  LAYER M2 ;
        RECT 3.244 0.908 3.316 0.94 ;
  LAYER M1 ;
        RECT 3.264 0.756 3.296 0.924 ;
  LAYER M1 ;
        RECT 3.264 0.72 3.296 0.792 ;
  LAYER M2 ;
        RECT 3.244 0.74 3.316 0.772 ;
  LAYER M2 ;
        RECT 3.28 0.74 6 0.772 ;
  LAYER M1 ;
        RECT 5.984 0.72 6.016 0.792 ;
  LAYER M2 ;
        RECT 5.964 0.74 6.036 0.772 ;
  LAYER M1 ;
        RECT 3.264 3.828 3.296 3.9 ;
  LAYER M2 ;
        RECT 3.244 3.848 3.316 3.88 ;
  LAYER M1 ;
        RECT 3.264 3.696 3.296 3.864 ;
  LAYER M1 ;
        RECT 3.264 3.66 3.296 3.732 ;
  LAYER M2 ;
        RECT 3.244 3.68 3.316 3.712 ;
  LAYER M2 ;
        RECT 3.28 3.68 6 3.712 ;
  LAYER M1 ;
        RECT 5.984 3.66 6.016 3.732 ;
  LAYER M2 ;
        RECT 5.964 3.68 6.036 3.712 ;
  LAYER M1 ;
        RECT 3.264 18.528 3.296 18.6 ;
  LAYER M2 ;
        RECT 3.244 18.548 3.316 18.58 ;
  LAYER M1 ;
        RECT 3.264 18.396 3.296 18.564 ;
  LAYER M1 ;
        RECT 3.264 18.36 3.296 18.432 ;
  LAYER M2 ;
        RECT 3.244 18.38 3.316 18.412 ;
  LAYER M2 ;
        RECT 3.28 18.38 6 18.412 ;
  LAYER M1 ;
        RECT 5.984 18.36 6.016 18.432 ;
  LAYER M2 ;
        RECT 5.964 18.38 6.036 18.412 ;
  LAYER M1 ;
        RECT 6.464 0.888 6.496 0.96 ;
  LAYER M2 ;
        RECT 6.444 0.908 6.516 0.94 ;
  LAYER M2 ;
        RECT 6 0.908 6.48 0.94 ;
  LAYER M1 ;
        RECT 5.984 0.888 6.016 0.96 ;
  LAYER M2 ;
        RECT 5.964 0.908 6.036 0.94 ;
  LAYER M1 ;
        RECT 6.464 9.708 6.496 9.78 ;
  LAYER M2 ;
        RECT 6.444 9.728 6.516 9.76 ;
  LAYER M2 ;
        RECT 6 9.728 6.48 9.76 ;
  LAYER M1 ;
        RECT 5.984 9.708 6.016 9.78 ;
  LAYER M2 ;
        RECT 5.964 9.728 6.036 9.76 ;
  LAYER M1 ;
        RECT 6.464 18.528 6.496 18.6 ;
  LAYER M2 ;
        RECT 6.444 18.548 6.516 18.58 ;
  LAYER M2 ;
        RECT 6 18.548 6.48 18.58 ;
  LAYER M1 ;
        RECT 5.984 18.528 6.016 18.6 ;
  LAYER M2 ;
        RECT 5.964 18.548 6.036 18.58 ;
  LAYER M1 ;
        RECT 5.984 0.048 6.016 0.12 ;
  LAYER M2 ;
        RECT 5.964 0.068 6.036 0.1 ;
  LAYER M1 ;
        RECT 5.984 0.084 6.016 0.588 ;
  LAYER M1 ;
        RECT 5.984 0.588 6.016 18.564 ;
  LAYER M1 ;
        RECT 9.664 0.888 9.696 0.96 ;
  LAYER M2 ;
        RECT 9.644 0.908 9.716 0.94 ;
  LAYER M2 ;
        RECT 9.2 0.908 9.68 0.94 ;
  LAYER M1 ;
        RECT 9.184 0.888 9.216 0.96 ;
  LAYER M2 ;
        RECT 9.164 0.908 9.236 0.94 ;
  LAYER M1 ;
        RECT 9.664 15.588 9.696 15.66 ;
  LAYER M2 ;
        RECT 9.644 15.608 9.716 15.64 ;
  LAYER M2 ;
        RECT 9.2 15.608 9.68 15.64 ;
  LAYER M1 ;
        RECT 9.184 15.588 9.216 15.66 ;
  LAYER M2 ;
        RECT 9.164 15.608 9.236 15.64 ;
  LAYER M1 ;
        RECT 9.664 18.528 9.696 18.6 ;
  LAYER M2 ;
        RECT 9.644 18.548 9.716 18.58 ;
  LAYER M2 ;
        RECT 9.2 18.548 9.68 18.58 ;
  LAYER M1 ;
        RECT 9.184 18.528 9.216 18.6 ;
  LAYER M2 ;
        RECT 9.164 18.548 9.236 18.58 ;
  LAYER M1 ;
        RECT 9.184 0.048 9.216 0.12 ;
  LAYER M2 ;
        RECT 9.164 0.068 9.236 0.1 ;
  LAYER M1 ;
        RECT 9.184 0.084 9.216 0.588 ;
  LAYER M1 ;
        RECT 9.184 0.588 9.216 18.564 ;
  LAYER M2 ;
        RECT 6 0.068 9.2 0.1 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M2 ;
        RECT 0.08 18.548 3.28 18.58 ;
  LAYER M1 ;
        RECT 3.264 18.528 3.296 18.6 ;
  LAYER M2 ;
        RECT 3.244 18.548 3.316 18.58 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.624 0.096 18.564 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.684 0.096 15.624 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.744 0.096 12.684 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.804 0.096 9.744 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.864 0.096 6.804 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.924 0.096 3.864 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 12.864 18.528 12.896 18.6 ;
  LAYER M2 ;
        RECT 12.844 18.548 12.916 18.58 ;
  LAYER M2 ;
        RECT 9.68 18.548 12.88 18.58 ;
  LAYER M1 ;
        RECT 9.664 18.528 9.696 18.6 ;
  LAYER M2 ;
        RECT 9.644 18.548 9.716 18.58 ;
  LAYER M1 ;
        RECT 12.864 15.588 12.896 15.66 ;
  LAYER M2 ;
        RECT 12.844 15.608 12.916 15.64 ;
  LAYER M2 ;
        RECT 9.68 15.608 12.88 15.64 ;
  LAYER M1 ;
        RECT 9.664 15.588 9.696 15.66 ;
  LAYER M2 ;
        RECT 9.644 15.608 9.716 15.64 ;
  LAYER M1 ;
        RECT 12.864 12.648 12.896 12.72 ;
  LAYER M2 ;
        RECT 12.844 12.668 12.916 12.7 ;
  LAYER M1 ;
        RECT 12.864 12.684 12.896 15.624 ;
  LAYER M1 ;
        RECT 12.864 15.588 12.896 15.66 ;
  LAYER M2 ;
        RECT 12.844 15.608 12.916 15.64 ;
  LAYER M1 ;
        RECT 12.864 9.708 12.896 9.78 ;
  LAYER M2 ;
        RECT 12.844 9.728 12.916 9.76 ;
  LAYER M1 ;
        RECT 12.864 9.744 12.896 12.684 ;
  LAYER M1 ;
        RECT 12.864 12.648 12.896 12.72 ;
  LAYER M2 ;
        RECT 12.844 12.668 12.916 12.7 ;
  LAYER M1 ;
        RECT 12.864 6.768 12.896 6.84 ;
  LAYER M2 ;
        RECT 12.844 6.788 12.916 6.82 ;
  LAYER M1 ;
        RECT 12.864 6.804 12.896 9.744 ;
  LAYER M1 ;
        RECT 12.864 9.708 12.896 9.78 ;
  LAYER M2 ;
        RECT 12.844 9.728 12.916 9.76 ;
  LAYER M1 ;
        RECT 12.864 3.828 12.896 3.9 ;
  LAYER M2 ;
        RECT 12.844 3.848 12.916 3.88 ;
  LAYER M1 ;
        RECT 12.864 3.864 12.896 6.804 ;
  LAYER M1 ;
        RECT 12.864 6.768 12.896 6.84 ;
  LAYER M2 ;
        RECT 12.844 6.788 12.916 6.82 ;
  LAYER M1 ;
        RECT 12.864 0.888 12.896 0.96 ;
  LAYER M2 ;
        RECT 12.844 0.908 12.916 0.94 ;
  LAYER M1 ;
        RECT 12.864 0.924 12.896 3.864 ;
  LAYER M1 ;
        RECT 12.864 3.828 12.896 3.9 ;
  LAYER M2 ;
        RECT 12.844 3.848 12.916 3.88 ;
  LAYER M1 ;
        RECT 5.664 12.144 5.696 12.216 ;
  LAYER M2 ;
        RECT 5.644 12.164 5.716 12.196 ;
  LAYER M2 ;
        RECT 2.8 12.164 5.68 12.196 ;
  LAYER M1 ;
        RECT 2.784 12.144 2.816 12.216 ;
  LAYER M2 ;
        RECT 2.764 12.164 2.836 12.196 ;
  LAYER M1 ;
        RECT 5.664 9.204 5.696 9.276 ;
  LAYER M2 ;
        RECT 5.644 9.224 5.716 9.256 ;
  LAYER M2 ;
        RECT 2.8 9.224 5.68 9.256 ;
  LAYER M1 ;
        RECT 2.784 9.204 2.816 9.276 ;
  LAYER M2 ;
        RECT 2.764 9.224 2.836 9.256 ;
  LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
  LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
  LAYER M1 ;
        RECT 2.784 21.336 2.816 21.504 ;
  LAYER M1 ;
        RECT 2.784 9.24 2.816 21.336 ;
  LAYER M1 ;
        RECT 12.064 12.144 12.096 12.216 ;
  LAYER M2 ;
        RECT 12.044 12.164 12.116 12.196 ;
  LAYER M1 ;
        RECT 12.064 12.18 12.096 12.348 ;
  LAYER M1 ;
        RECT 12.064 12.312 12.096 12.384 ;
  LAYER M2 ;
        RECT 12.044 12.332 12.116 12.364 ;
  LAYER M2 ;
        RECT 12.08 12.332 12.4 12.364 ;
  LAYER M1 ;
        RECT 12.384 12.312 12.416 12.384 ;
  LAYER M2 ;
        RECT 12.364 12.332 12.436 12.364 ;
  LAYER M1 ;
        RECT 12.064 15.084 12.096 15.156 ;
  LAYER M2 ;
        RECT 12.044 15.104 12.116 15.136 ;
  LAYER M1 ;
        RECT 12.064 15.12 12.096 15.288 ;
  LAYER M1 ;
        RECT 12.064 15.252 12.096 15.324 ;
  LAYER M2 ;
        RECT 12.044 15.272 12.116 15.304 ;
  LAYER M2 ;
        RECT 12.08 15.272 12.4 15.304 ;
  LAYER M1 ;
        RECT 12.384 15.252 12.416 15.324 ;
  LAYER M2 ;
        RECT 12.364 15.272 12.436 15.304 ;
  LAYER M1 ;
        RECT 12.384 21.468 12.416 21.54 ;
  LAYER M2 ;
        RECT 12.364 21.488 12.436 21.52 ;
  LAYER M1 ;
        RECT 12.384 21.336 12.416 21.504 ;
  LAYER M1 ;
        RECT 12.384 12.348 12.416 21.336 ;
  LAYER M2 ;
        RECT 2.8 21.488 12.4 21.52 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M2 ;
        RECT 5.68 9.224 8.88 9.256 ;
  LAYER M1 ;
        RECT 5.664 9.204 5.696 9.276 ;
  LAYER M2 ;
        RECT 5.644 9.224 5.716 9.256 ;
  LAYER M1 ;
        RECT 8.864 15.084 8.896 15.156 ;
  LAYER M2 ;
        RECT 8.844 15.104 8.916 15.136 ;
  LAYER M2 ;
        RECT 8.88 15.104 12.08 15.136 ;
  LAYER M1 ;
        RECT 12.064 15.084 12.096 15.156 ;
  LAYER M2 ;
        RECT 12.044 15.104 12.116 15.136 ;
  LAYER M1 ;
        RECT 5.664 15.084 5.696 15.156 ;
  LAYER M2 ;
        RECT 5.644 15.104 5.716 15.136 ;
  LAYER M1 ;
        RECT 5.664 15.12 5.696 15.288 ;
  LAYER M1 ;
        RECT 5.664 15.252 5.696 15.324 ;
  LAYER M2 ;
        RECT 5.644 15.272 5.716 15.304 ;
  LAYER M2 ;
        RECT 5.68 15.272 6.16 15.304 ;
  LAYER M1 ;
        RECT 6.144 15.252 6.176 15.324 ;
  LAYER M2 ;
        RECT 6.124 15.272 6.196 15.304 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M2 ;
        RECT 6.16 6.284 8.88 6.316 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M1 ;
        RECT 8.864 18.024 8.896 18.096 ;
  LAYER M2 ;
        RECT 8.844 18.044 8.916 18.076 ;
  LAYER M2 ;
        RECT 6.16 18.044 8.88 18.076 ;
  LAYER M1 ;
        RECT 6.144 18.024 6.176 18.096 ;
  LAYER M2 ;
        RECT 6.124 18.044 6.196 18.076 ;
  LAYER M1 ;
        RECT 5.664 18.024 5.696 18.096 ;
  LAYER M2 ;
        RECT 5.644 18.044 5.716 18.076 ;
  LAYER M1 ;
        RECT 5.664 18.06 5.696 18.228 ;
  LAYER M1 ;
        RECT 5.664 18.192 5.696 18.264 ;
  LAYER M2 ;
        RECT 5.644 18.212 5.716 18.244 ;
  LAYER M2 ;
        RECT 5.68 18.212 6.16 18.244 ;
  LAYER M1 ;
        RECT 6.144 18.192 6.176 18.264 ;
  LAYER M2 ;
        RECT 6.124 18.212 6.196 18.244 ;
  LAYER M1 ;
        RECT 6.144 21.636 6.176 21.708 ;
  LAYER M2 ;
        RECT 6.124 21.656 6.196 21.688 ;
  LAYER M1 ;
        RECT 6.144 21.336 6.176 21.672 ;
  LAYER M1 ;
        RECT 6.144 6.3 6.176 21.336 ;
  LAYER M1 ;
        RECT 12.064 9.204 12.096 9.276 ;
  LAYER M2 ;
        RECT 12.044 9.224 12.116 9.256 ;
  LAYER M2 ;
        RECT 9.36 9.224 12.08 9.256 ;
  LAYER M1 ;
        RECT 9.344 9.204 9.376 9.276 ;
  LAYER M2 ;
        RECT 9.324 9.224 9.396 9.256 ;
  LAYER M1 ;
        RECT 12.064 6.264 12.096 6.336 ;
  LAYER M2 ;
        RECT 12.044 6.284 12.116 6.316 ;
  LAYER M2 ;
        RECT 9.36 6.284 12.08 6.316 ;
  LAYER M1 ;
        RECT 9.344 6.264 9.376 6.336 ;
  LAYER M2 ;
        RECT 9.324 6.284 9.396 6.316 ;
  LAYER M1 ;
        RECT 9.344 21.636 9.376 21.708 ;
  LAYER M2 ;
        RECT 9.324 21.656 9.396 21.688 ;
  LAYER M1 ;
        RECT 9.344 21.336 9.376 21.672 ;
  LAYER M1 ;
        RECT 9.344 6.3 9.376 21.336 ;
  LAYER M2 ;
        RECT 6.16 21.656 9.36 21.688 ;
  LAYER M1 ;
        RECT 5.664 3.324 5.696 3.396 ;
  LAYER M2 ;
        RECT 5.644 3.344 5.716 3.376 ;
  LAYER M1 ;
        RECT 5.664 3.36 5.696 3.528 ;
  LAYER M1 ;
        RECT 5.664 3.492 5.696 3.564 ;
  LAYER M2 ;
        RECT 5.644 3.512 5.716 3.544 ;
  LAYER M2 ;
        RECT 5.68 3.512 6.32 3.544 ;
  LAYER M1 ;
        RECT 6.304 3.492 6.336 3.564 ;
  LAYER M2 ;
        RECT 6.284 3.512 6.356 3.544 ;
  LAYER M1 ;
        RECT 5.664 6.264 5.696 6.336 ;
  LAYER M2 ;
        RECT 5.644 6.284 5.716 6.316 ;
  LAYER M1 ;
        RECT 5.664 6.3 5.696 6.468 ;
  LAYER M1 ;
        RECT 5.664 6.432 5.696 6.504 ;
  LAYER M2 ;
        RECT 5.644 6.452 5.716 6.484 ;
  LAYER M2 ;
        RECT 5.68 6.452 6.32 6.484 ;
  LAYER M1 ;
        RECT 6.304 6.432 6.336 6.504 ;
  LAYER M2 ;
        RECT 6.284 6.452 6.356 6.484 ;
  LAYER M1 ;
        RECT 5.664 20.964 5.696 21.036 ;
  LAYER M2 ;
        RECT 5.644 20.984 5.716 21.016 ;
  LAYER M1 ;
        RECT 5.664 21 5.696 21.168 ;
  LAYER M1 ;
        RECT 5.664 21.132 5.696 21.204 ;
  LAYER M2 ;
        RECT 5.644 21.152 5.716 21.184 ;
  LAYER M2 ;
        RECT 5.68 21.152 6.32 21.184 ;
  LAYER M1 ;
        RECT 6.304 21.132 6.336 21.204 ;
  LAYER M2 ;
        RECT 6.284 21.152 6.356 21.184 ;
  LAYER M1 ;
        RECT 8.864 3.324 8.896 3.396 ;
  LAYER M2 ;
        RECT 8.844 3.344 8.916 3.376 ;
  LAYER M2 ;
        RECT 6.32 3.344 8.88 3.376 ;
  LAYER M1 ;
        RECT 6.304 3.324 6.336 3.396 ;
  LAYER M2 ;
        RECT 6.284 3.344 6.356 3.376 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M2 ;
        RECT 6.32 12.164 8.88 12.196 ;
  LAYER M1 ;
        RECT 6.304 12.144 6.336 12.216 ;
  LAYER M2 ;
        RECT 6.284 12.164 6.356 12.196 ;
  LAYER M1 ;
        RECT 8.864 20.964 8.896 21.036 ;
  LAYER M2 ;
        RECT 8.844 20.984 8.916 21.016 ;
  LAYER M2 ;
        RECT 6.32 20.984 8.88 21.016 ;
  LAYER M1 ;
        RECT 6.304 20.964 6.336 21.036 ;
  LAYER M2 ;
        RECT 6.284 20.984 6.356 21.016 ;
  LAYER M1 ;
        RECT 6.304 21.804 6.336 21.876 ;
  LAYER M2 ;
        RECT 6.284 21.824 6.356 21.856 ;
  LAYER M1 ;
        RECT 6.304 21.336 6.336 21.84 ;
  LAYER M1 ;
        RECT 6.304 3.36 6.336 21.336 ;
  LAYER M1 ;
        RECT 12.064 3.324 12.096 3.396 ;
  LAYER M2 ;
        RECT 12.044 3.344 12.116 3.376 ;
  LAYER M2 ;
        RECT 9.52 3.344 12.08 3.376 ;
  LAYER M1 ;
        RECT 9.504 3.324 9.536 3.396 ;
  LAYER M2 ;
        RECT 9.484 3.344 9.556 3.376 ;
  LAYER M1 ;
        RECT 12.064 18.024 12.096 18.096 ;
  LAYER M2 ;
        RECT 12.044 18.044 12.116 18.076 ;
  LAYER M2 ;
        RECT 9.52 18.044 12.08 18.076 ;
  LAYER M1 ;
        RECT 9.504 18.024 9.536 18.096 ;
  LAYER M2 ;
        RECT 9.484 18.044 9.556 18.076 ;
  LAYER M1 ;
        RECT 12.064 20.964 12.096 21.036 ;
  LAYER M2 ;
        RECT 12.044 20.984 12.116 21.016 ;
  LAYER M2 ;
        RECT 9.52 20.984 12.08 21.016 ;
  LAYER M1 ;
        RECT 9.504 20.964 9.536 21.036 ;
  LAYER M2 ;
        RECT 9.484 20.984 9.556 21.016 ;
  LAYER M1 ;
        RECT 9.504 21.804 9.536 21.876 ;
  LAYER M2 ;
        RECT 9.484 21.824 9.556 21.856 ;
  LAYER M1 ;
        RECT 9.504 21.336 9.536 21.84 ;
  LAYER M1 ;
        RECT 9.504 3.36 9.536 21.336 ;
  LAYER M2 ;
        RECT 6.32 21.824 9.52 21.856 ;
  LAYER M1 ;
        RECT 2.464 20.964 2.496 21.036 ;
  LAYER M2 ;
        RECT 2.444 20.984 2.516 21.016 ;
  LAYER M2 ;
        RECT 2.48 20.984 5.68 21.016 ;
  LAYER M1 ;
        RECT 5.664 20.964 5.696 21.036 ;
  LAYER M2 ;
        RECT 5.644 20.984 5.716 21.016 ;
  LAYER M1 ;
        RECT 2.464 18.024 2.496 18.096 ;
  LAYER M2 ;
        RECT 2.444 18.044 2.516 18.076 ;
  LAYER M1 ;
        RECT 2.464 18.06 2.496 21 ;
  LAYER M1 ;
        RECT 2.464 20.964 2.496 21.036 ;
  LAYER M2 ;
        RECT 2.444 20.984 2.516 21.016 ;
  LAYER M1 ;
        RECT 2.464 15.084 2.496 15.156 ;
  LAYER M2 ;
        RECT 2.444 15.104 2.516 15.136 ;
  LAYER M1 ;
        RECT 2.464 15.12 2.496 18.06 ;
  LAYER M1 ;
        RECT 2.464 18.024 2.496 18.096 ;
  LAYER M2 ;
        RECT 2.444 18.044 2.516 18.076 ;
  LAYER M1 ;
        RECT 2.464 12.144 2.496 12.216 ;
  LAYER M2 ;
        RECT 2.444 12.164 2.516 12.196 ;
  LAYER M1 ;
        RECT 2.464 12.18 2.496 15.12 ;
  LAYER M1 ;
        RECT 2.464 15.084 2.496 15.156 ;
  LAYER M2 ;
        RECT 2.444 15.104 2.516 15.136 ;
  LAYER M1 ;
        RECT 2.464 9.204 2.496 9.276 ;
  LAYER M2 ;
        RECT 2.444 9.224 2.516 9.256 ;
  LAYER M1 ;
        RECT 2.464 9.24 2.496 12.18 ;
  LAYER M1 ;
        RECT 2.464 12.144 2.496 12.216 ;
  LAYER M2 ;
        RECT 2.444 12.164 2.516 12.196 ;
  LAYER M1 ;
        RECT 2.464 6.264 2.496 6.336 ;
  LAYER M2 ;
        RECT 2.444 6.284 2.516 6.316 ;
  LAYER M1 ;
        RECT 2.464 6.3 2.496 9.24 ;
  LAYER M1 ;
        RECT 2.464 9.204 2.496 9.276 ;
  LAYER M2 ;
        RECT 2.444 9.224 2.516 9.256 ;
  LAYER M1 ;
        RECT 2.464 3.324 2.496 3.396 ;
  LAYER M2 ;
        RECT 2.444 3.344 2.516 3.376 ;
  LAYER M1 ;
        RECT 2.464 3.36 2.496 6.3 ;
  LAYER M1 ;
        RECT 2.464 6.264 2.496 6.336 ;
  LAYER M2 ;
        RECT 2.444 6.284 2.516 6.316 ;
  LAYER M1 ;
        RECT 15.264 20.964 15.296 21.036 ;
  LAYER M2 ;
        RECT 15.244 20.984 15.316 21.016 ;
  LAYER M2 ;
        RECT 12.08 20.984 15.28 21.016 ;
  LAYER M1 ;
        RECT 12.064 20.964 12.096 21.036 ;
  LAYER M2 ;
        RECT 12.044 20.984 12.116 21.016 ;
  LAYER M1 ;
        RECT 15.264 18.024 15.296 18.096 ;
  LAYER M2 ;
        RECT 15.244 18.044 15.316 18.076 ;
  LAYER M2 ;
        RECT 12.08 18.044 15.28 18.076 ;
  LAYER M1 ;
        RECT 12.064 18.024 12.096 18.096 ;
  LAYER M2 ;
        RECT 12.044 18.044 12.116 18.076 ;
  LAYER M1 ;
        RECT 15.264 15.084 15.296 15.156 ;
  LAYER M2 ;
        RECT 15.244 15.104 15.316 15.136 ;
  LAYER M1 ;
        RECT 15.264 15.12 15.296 18.06 ;
  LAYER M1 ;
        RECT 15.264 18.024 15.296 18.096 ;
  LAYER M2 ;
        RECT 15.244 18.044 15.316 18.076 ;
  LAYER M1 ;
        RECT 15.264 12.144 15.296 12.216 ;
  LAYER M2 ;
        RECT 15.244 12.164 15.316 12.196 ;
  LAYER M1 ;
        RECT 15.264 12.18 15.296 15.12 ;
  LAYER M1 ;
        RECT 15.264 15.084 15.296 15.156 ;
  LAYER M2 ;
        RECT 15.244 15.104 15.316 15.136 ;
  LAYER M1 ;
        RECT 15.264 9.204 15.296 9.276 ;
  LAYER M2 ;
        RECT 15.244 9.224 15.316 9.256 ;
  LAYER M1 ;
        RECT 15.264 9.24 15.296 12.18 ;
  LAYER M1 ;
        RECT 15.264 12.144 15.296 12.216 ;
  LAYER M2 ;
        RECT 15.244 12.164 15.316 12.196 ;
  LAYER M1 ;
        RECT 15.264 6.264 15.296 6.336 ;
  LAYER M2 ;
        RECT 15.244 6.284 15.316 6.316 ;
  LAYER M1 ;
        RECT 15.264 6.3 15.296 9.24 ;
  LAYER M1 ;
        RECT 15.264 9.204 15.296 9.276 ;
  LAYER M2 ;
        RECT 15.244 9.224 15.316 9.256 ;
  LAYER M1 ;
        RECT 15.264 3.324 15.296 3.396 ;
  LAYER M2 ;
        RECT 15.244 3.344 15.316 3.376 ;
  LAYER M1 ;
        RECT 15.264 3.36 15.296 6.3 ;
  LAYER M1 ;
        RECT 15.264 6.264 15.296 6.336 ;
  LAYER M2 ;
        RECT 15.244 6.284 15.316 6.316 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 3.396 ;
  LAYER M1 ;
        RECT 0.128 0.888 0.16 3.396 ;
  LAYER M1 ;
        RECT 0.192 0.888 0.224 3.396 ;
  LAYER M1 ;
        RECT 0.256 0.888 0.288 3.396 ;
  LAYER M1 ;
        RECT 0.32 0.888 0.352 3.396 ;
  LAYER M1 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M1 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M1 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M1 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M1 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M1 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M1 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M1 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M1 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M1 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M1 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M1 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M1 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M1 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M1 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M1 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M1 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M1 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M1 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M1 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M1 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M1 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M1 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M1 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M1 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M1 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M1 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M1 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M1 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M1 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M1 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M2 ;
        RECT 0.044 0.972 2.516 1.004 ;
  LAYER M2 ;
        RECT 0.044 1.036 2.516 1.068 ;
  LAYER M2 ;
        RECT 0.044 1.1 2.516 1.132 ;
  LAYER M2 ;
        RECT 0.044 1.164 2.516 1.196 ;
  LAYER M2 ;
        RECT 0.044 1.228 2.516 1.26 ;
  LAYER M2 ;
        RECT 0.044 1.292 2.516 1.324 ;
  LAYER M2 ;
        RECT 0.044 1.356 2.516 1.388 ;
  LAYER M2 ;
        RECT 0.044 1.42 2.516 1.452 ;
  LAYER M2 ;
        RECT 0.044 1.484 2.516 1.516 ;
  LAYER M2 ;
        RECT 0.044 1.548 2.516 1.58 ;
  LAYER M2 ;
        RECT 0.044 1.612 2.516 1.644 ;
  LAYER M2 ;
        RECT 0.044 1.676 2.516 1.708 ;
  LAYER M2 ;
        RECT 0.044 1.74 2.516 1.772 ;
  LAYER M2 ;
        RECT 0.044 1.804 2.516 1.836 ;
  LAYER M2 ;
        RECT 0.044 1.868 2.516 1.9 ;
  LAYER M2 ;
        RECT 0.044 1.932 2.516 1.964 ;
  LAYER M2 ;
        RECT 0.044 1.996 2.516 2.028 ;
  LAYER M2 ;
        RECT 0.044 2.06 2.516 2.092 ;
  LAYER M2 ;
        RECT 0.044 2.124 2.516 2.156 ;
  LAYER M2 ;
        RECT 0.044 2.188 2.516 2.22 ;
  LAYER M2 ;
        RECT 0.044 2.252 2.516 2.284 ;
  LAYER M2 ;
        RECT 0.044 2.316 2.516 2.348 ;
  LAYER M2 ;
        RECT 0.044 2.38 2.516 2.412 ;
  LAYER M2 ;
        RECT 0.044 2.444 2.516 2.476 ;
  LAYER M2 ;
        RECT 0.044 2.508 2.516 2.54 ;
  LAYER M2 ;
        RECT 0.044 2.572 2.516 2.604 ;
  LAYER M2 ;
        RECT 0.044 2.636 2.516 2.668 ;
  LAYER M2 ;
        RECT 0.044 2.7 2.516 2.732 ;
  LAYER M2 ;
        RECT 0.044 2.764 2.516 2.796 ;
  LAYER M2 ;
        RECT 0.044 2.828 2.516 2.86 ;
  LAYER M2 ;
        RECT 0.044 2.892 2.516 2.924 ;
  LAYER M2 ;
        RECT 0.044 2.956 2.516 2.988 ;
  LAYER M2 ;
        RECT 0.044 3.02 2.516 3.052 ;
  LAYER M2 ;
        RECT 0.044 3.084 2.516 3.116 ;
  LAYER M2 ;
        RECT 0.044 3.148 2.516 3.18 ;
  LAYER M2 ;
        RECT 0.044 3.212 2.516 3.244 ;
  LAYER M3 ;
        RECT 0.064 0.888 0.096 3.396 ;
  LAYER M3 ;
        RECT 0.128 0.888 0.16 3.396 ;
  LAYER M3 ;
        RECT 0.192 0.888 0.224 3.396 ;
  LAYER M3 ;
        RECT 0.256 0.888 0.288 3.396 ;
  LAYER M3 ;
        RECT 0.32 0.888 0.352 3.396 ;
  LAYER M3 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M3 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M3 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M3 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M3 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M3 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M3 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M3 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M3 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M3 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M3 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M3 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M3 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M3 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M3 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M3 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M3 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M3 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M3 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M3 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M3 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M3 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M3 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M3 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M3 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M3 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M3 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M3 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M3 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M3 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M3 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M3 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M3 ;
        RECT 2.464 0.888 2.496 3.396 ;
  LAYER M1 ;
        RECT 0.079 0.924 0.081 3.36 ;
  LAYER M1 ;
        RECT 0.159 0.924 0.161 3.36 ;
  LAYER M1 ;
        RECT 0.239 0.924 0.241 3.36 ;
  LAYER M1 ;
        RECT 0.319 0.924 0.321 3.36 ;
  LAYER M1 ;
        RECT 0.399 0.924 0.401 3.36 ;
  LAYER M1 ;
        RECT 0.479 0.924 0.481 3.36 ;
  LAYER M1 ;
        RECT 0.559 0.924 0.561 3.36 ;
  LAYER M1 ;
        RECT 0.639 0.924 0.641 3.36 ;
  LAYER M1 ;
        RECT 0.719 0.924 0.721 3.36 ;
  LAYER M1 ;
        RECT 0.799 0.924 0.801 3.36 ;
  LAYER M1 ;
        RECT 0.879 0.924 0.881 3.36 ;
  LAYER M1 ;
        RECT 0.959 0.924 0.961 3.36 ;
  LAYER M1 ;
        RECT 1.039 0.924 1.041 3.36 ;
  LAYER M1 ;
        RECT 1.119 0.924 1.121 3.36 ;
  LAYER M1 ;
        RECT 1.199 0.924 1.201 3.36 ;
  LAYER M1 ;
        RECT 1.279 0.924 1.281 3.36 ;
  LAYER M1 ;
        RECT 1.359 0.924 1.361 3.36 ;
  LAYER M1 ;
        RECT 1.439 0.924 1.441 3.36 ;
  LAYER M1 ;
        RECT 1.519 0.924 1.521 3.36 ;
  LAYER M1 ;
        RECT 1.599 0.924 1.601 3.36 ;
  LAYER M1 ;
        RECT 1.679 0.924 1.681 3.36 ;
  LAYER M1 ;
        RECT 1.759 0.924 1.761 3.36 ;
  LAYER M1 ;
        RECT 1.839 0.924 1.841 3.36 ;
  LAYER M1 ;
        RECT 1.919 0.924 1.921 3.36 ;
  LAYER M1 ;
        RECT 1.999 0.924 2.001 3.36 ;
  LAYER M1 ;
        RECT 2.079 0.924 2.081 3.36 ;
  LAYER M1 ;
        RECT 2.159 0.924 2.161 3.36 ;
  LAYER M1 ;
        RECT 2.239 0.924 2.241 3.36 ;
  LAYER M1 ;
        RECT 2.319 0.924 2.321 3.36 ;
  LAYER M1 ;
        RECT 2.399 0.924 2.401 3.36 ;
  LAYER M2 ;
        RECT 0.08 0.923 2.48 0.925 ;
  LAYER M2 ;
        RECT 0.08 1.007 2.48 1.009 ;
  LAYER M2 ;
        RECT 0.08 1.091 2.48 1.093 ;
  LAYER M2 ;
        RECT 0.08 1.175 2.48 1.177 ;
  LAYER M2 ;
        RECT 0.08 1.259 2.48 1.261 ;
  LAYER M2 ;
        RECT 0.08 1.343 2.48 1.345 ;
  LAYER M2 ;
        RECT 0.08 1.427 2.48 1.429 ;
  LAYER M2 ;
        RECT 0.08 1.511 2.48 1.513 ;
  LAYER M2 ;
        RECT 0.08 1.595 2.48 1.597 ;
  LAYER M2 ;
        RECT 0.08 1.679 2.48 1.681 ;
  LAYER M2 ;
        RECT 0.08 1.763 2.48 1.765 ;
  LAYER M2 ;
        RECT 0.08 1.847 2.48 1.849 ;
  LAYER M2 ;
        RECT 0.08 1.9305 2.48 1.9325 ;
  LAYER M2 ;
        RECT 0.08 2.015 2.48 2.017 ;
  LAYER M2 ;
        RECT 0.08 2.099 2.48 2.101 ;
  LAYER M2 ;
        RECT 0.08 2.183 2.48 2.185 ;
  LAYER M2 ;
        RECT 0.08 2.267 2.48 2.269 ;
  LAYER M2 ;
        RECT 0.08 2.351 2.48 2.353 ;
  LAYER M2 ;
        RECT 0.08 2.435 2.48 2.437 ;
  LAYER M2 ;
        RECT 0.08 2.519 2.48 2.521 ;
  LAYER M2 ;
        RECT 0.08 2.603 2.48 2.605 ;
  LAYER M2 ;
        RECT 0.08 2.687 2.48 2.689 ;
  LAYER M2 ;
        RECT 0.08 2.771 2.48 2.773 ;
  LAYER M2 ;
        RECT 0.08 2.855 2.48 2.857 ;
  LAYER M2 ;
        RECT 0.08 2.939 2.48 2.941 ;
  LAYER M2 ;
        RECT 0.08 3.023 2.48 3.025 ;
  LAYER M2 ;
        RECT 0.08 3.107 2.48 3.109 ;
  LAYER M2 ;
        RECT 0.08 3.191 2.48 3.193 ;
  LAYER M2 ;
        RECT 0.08 3.275 2.48 3.277 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 6.336 ;
  LAYER M1 ;
        RECT 0.128 3.828 0.16 6.336 ;
  LAYER M1 ;
        RECT 0.192 3.828 0.224 6.336 ;
  LAYER M1 ;
        RECT 0.256 3.828 0.288 6.336 ;
  LAYER M1 ;
        RECT 0.32 3.828 0.352 6.336 ;
  LAYER M1 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M1 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M1 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M1 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M1 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M1 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M1 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M1 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M1 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M1 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M1 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M1 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M1 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M1 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M1 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M1 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M1 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M1 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M1 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M1 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M1 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M1 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M1 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M1 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M1 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M1 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M1 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M1 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M1 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M1 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M1 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M1 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M2 ;
        RECT 0.044 3.912 2.516 3.944 ;
  LAYER M2 ;
        RECT 0.044 3.976 2.516 4.008 ;
  LAYER M2 ;
        RECT 0.044 4.04 2.516 4.072 ;
  LAYER M2 ;
        RECT 0.044 4.104 2.516 4.136 ;
  LAYER M2 ;
        RECT 0.044 4.168 2.516 4.2 ;
  LAYER M2 ;
        RECT 0.044 4.232 2.516 4.264 ;
  LAYER M2 ;
        RECT 0.044 4.296 2.516 4.328 ;
  LAYER M2 ;
        RECT 0.044 4.36 2.516 4.392 ;
  LAYER M2 ;
        RECT 0.044 4.424 2.516 4.456 ;
  LAYER M2 ;
        RECT 0.044 4.488 2.516 4.52 ;
  LAYER M2 ;
        RECT 0.044 4.552 2.516 4.584 ;
  LAYER M2 ;
        RECT 0.044 4.616 2.516 4.648 ;
  LAYER M2 ;
        RECT 0.044 4.68 2.516 4.712 ;
  LAYER M2 ;
        RECT 0.044 4.744 2.516 4.776 ;
  LAYER M2 ;
        RECT 0.044 4.808 2.516 4.84 ;
  LAYER M2 ;
        RECT 0.044 4.872 2.516 4.904 ;
  LAYER M2 ;
        RECT 0.044 4.936 2.516 4.968 ;
  LAYER M2 ;
        RECT 0.044 5 2.516 5.032 ;
  LAYER M2 ;
        RECT 0.044 5.064 2.516 5.096 ;
  LAYER M2 ;
        RECT 0.044 5.128 2.516 5.16 ;
  LAYER M2 ;
        RECT 0.044 5.192 2.516 5.224 ;
  LAYER M2 ;
        RECT 0.044 5.256 2.516 5.288 ;
  LAYER M2 ;
        RECT 0.044 5.32 2.516 5.352 ;
  LAYER M2 ;
        RECT 0.044 5.384 2.516 5.416 ;
  LAYER M2 ;
        RECT 0.044 5.448 2.516 5.48 ;
  LAYER M2 ;
        RECT 0.044 5.512 2.516 5.544 ;
  LAYER M2 ;
        RECT 0.044 5.576 2.516 5.608 ;
  LAYER M2 ;
        RECT 0.044 5.64 2.516 5.672 ;
  LAYER M2 ;
        RECT 0.044 5.704 2.516 5.736 ;
  LAYER M2 ;
        RECT 0.044 5.768 2.516 5.8 ;
  LAYER M2 ;
        RECT 0.044 5.832 2.516 5.864 ;
  LAYER M2 ;
        RECT 0.044 5.896 2.516 5.928 ;
  LAYER M2 ;
        RECT 0.044 5.96 2.516 5.992 ;
  LAYER M2 ;
        RECT 0.044 6.024 2.516 6.056 ;
  LAYER M2 ;
        RECT 0.044 6.088 2.516 6.12 ;
  LAYER M2 ;
        RECT 0.044 6.152 2.516 6.184 ;
  LAYER M3 ;
        RECT 0.064 3.828 0.096 6.336 ;
  LAYER M3 ;
        RECT 0.128 3.828 0.16 6.336 ;
  LAYER M3 ;
        RECT 0.192 3.828 0.224 6.336 ;
  LAYER M3 ;
        RECT 0.256 3.828 0.288 6.336 ;
  LAYER M3 ;
        RECT 0.32 3.828 0.352 6.336 ;
  LAYER M3 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M3 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M3 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M3 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M3 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M3 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M3 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M3 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M3 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M3 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M3 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M3 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M3 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M3 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M3 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M3 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M3 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M3 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M3 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M3 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M3 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M3 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M3 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M3 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M3 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M3 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M3 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M3 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M3 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M3 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M3 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M3 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M3 ;
        RECT 2.464 3.828 2.496 6.336 ;
  LAYER M1 ;
        RECT 0.079 3.864 0.081 6.3 ;
  LAYER M1 ;
        RECT 0.159 3.864 0.161 6.3 ;
  LAYER M1 ;
        RECT 0.239 3.864 0.241 6.3 ;
  LAYER M1 ;
        RECT 0.319 3.864 0.321 6.3 ;
  LAYER M1 ;
        RECT 0.399 3.864 0.401 6.3 ;
  LAYER M1 ;
        RECT 0.479 3.864 0.481 6.3 ;
  LAYER M1 ;
        RECT 0.559 3.864 0.561 6.3 ;
  LAYER M1 ;
        RECT 0.639 3.864 0.641 6.3 ;
  LAYER M1 ;
        RECT 0.719 3.864 0.721 6.3 ;
  LAYER M1 ;
        RECT 0.799 3.864 0.801 6.3 ;
  LAYER M1 ;
        RECT 0.879 3.864 0.881 6.3 ;
  LAYER M1 ;
        RECT 0.959 3.864 0.961 6.3 ;
  LAYER M1 ;
        RECT 1.039 3.864 1.041 6.3 ;
  LAYER M1 ;
        RECT 1.119 3.864 1.121 6.3 ;
  LAYER M1 ;
        RECT 1.199 3.864 1.201 6.3 ;
  LAYER M1 ;
        RECT 1.279 3.864 1.281 6.3 ;
  LAYER M1 ;
        RECT 1.359 3.864 1.361 6.3 ;
  LAYER M1 ;
        RECT 1.439 3.864 1.441 6.3 ;
  LAYER M1 ;
        RECT 1.519 3.864 1.521 6.3 ;
  LAYER M1 ;
        RECT 1.599 3.864 1.601 6.3 ;
  LAYER M1 ;
        RECT 1.679 3.864 1.681 6.3 ;
  LAYER M1 ;
        RECT 1.759 3.864 1.761 6.3 ;
  LAYER M1 ;
        RECT 1.839 3.864 1.841 6.3 ;
  LAYER M1 ;
        RECT 1.919 3.864 1.921 6.3 ;
  LAYER M1 ;
        RECT 1.999 3.864 2.001 6.3 ;
  LAYER M1 ;
        RECT 2.079 3.864 2.081 6.3 ;
  LAYER M1 ;
        RECT 2.159 3.864 2.161 6.3 ;
  LAYER M1 ;
        RECT 2.239 3.864 2.241 6.3 ;
  LAYER M1 ;
        RECT 2.319 3.864 2.321 6.3 ;
  LAYER M1 ;
        RECT 2.399 3.864 2.401 6.3 ;
  LAYER M2 ;
        RECT 0.08 3.863 2.48 3.865 ;
  LAYER M2 ;
        RECT 0.08 3.947 2.48 3.949 ;
  LAYER M2 ;
        RECT 0.08 4.031 2.48 4.033 ;
  LAYER M2 ;
        RECT 0.08 4.115 2.48 4.117 ;
  LAYER M2 ;
        RECT 0.08 4.199 2.48 4.201 ;
  LAYER M2 ;
        RECT 0.08 4.283 2.48 4.285 ;
  LAYER M2 ;
        RECT 0.08 4.367 2.48 4.369 ;
  LAYER M2 ;
        RECT 0.08 4.451 2.48 4.453 ;
  LAYER M2 ;
        RECT 0.08 4.535 2.48 4.537 ;
  LAYER M2 ;
        RECT 0.08 4.619 2.48 4.621 ;
  LAYER M2 ;
        RECT 0.08 4.703 2.48 4.705 ;
  LAYER M2 ;
        RECT 0.08 4.787 2.48 4.789 ;
  LAYER M2 ;
        RECT 0.08 4.8705 2.48 4.8725 ;
  LAYER M2 ;
        RECT 0.08 4.955 2.48 4.957 ;
  LAYER M2 ;
        RECT 0.08 5.039 2.48 5.041 ;
  LAYER M2 ;
        RECT 0.08 5.123 2.48 5.125 ;
  LAYER M2 ;
        RECT 0.08 5.207 2.48 5.209 ;
  LAYER M2 ;
        RECT 0.08 5.291 2.48 5.293 ;
  LAYER M2 ;
        RECT 0.08 5.375 2.48 5.377 ;
  LAYER M2 ;
        RECT 0.08 5.459 2.48 5.461 ;
  LAYER M2 ;
        RECT 0.08 5.543 2.48 5.545 ;
  LAYER M2 ;
        RECT 0.08 5.627 2.48 5.629 ;
  LAYER M2 ;
        RECT 0.08 5.711 2.48 5.713 ;
  LAYER M2 ;
        RECT 0.08 5.795 2.48 5.797 ;
  LAYER M2 ;
        RECT 0.08 5.879 2.48 5.881 ;
  LAYER M2 ;
        RECT 0.08 5.963 2.48 5.965 ;
  LAYER M2 ;
        RECT 0.08 6.047 2.48 6.049 ;
  LAYER M2 ;
        RECT 0.08 6.131 2.48 6.133 ;
  LAYER M2 ;
        RECT 0.08 6.215 2.48 6.217 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 9.276 ;
  LAYER M1 ;
        RECT 0.128 6.768 0.16 9.276 ;
  LAYER M1 ;
        RECT 0.192 6.768 0.224 9.276 ;
  LAYER M1 ;
        RECT 0.256 6.768 0.288 9.276 ;
  LAYER M1 ;
        RECT 0.32 6.768 0.352 9.276 ;
  LAYER M1 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M1 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M1 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M1 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M1 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M1 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M1 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M1 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M1 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M1 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M1 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M1 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M1 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M1 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M1 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M1 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M1 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M1 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M1 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M1 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M1 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M1 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M1 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M1 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M1 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M1 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M1 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M1 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M1 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M1 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M1 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M1 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M2 ;
        RECT 0.044 6.852 2.516 6.884 ;
  LAYER M2 ;
        RECT 0.044 6.916 2.516 6.948 ;
  LAYER M2 ;
        RECT 0.044 6.98 2.516 7.012 ;
  LAYER M2 ;
        RECT 0.044 7.044 2.516 7.076 ;
  LAYER M2 ;
        RECT 0.044 7.108 2.516 7.14 ;
  LAYER M2 ;
        RECT 0.044 7.172 2.516 7.204 ;
  LAYER M2 ;
        RECT 0.044 7.236 2.516 7.268 ;
  LAYER M2 ;
        RECT 0.044 7.3 2.516 7.332 ;
  LAYER M2 ;
        RECT 0.044 7.364 2.516 7.396 ;
  LAYER M2 ;
        RECT 0.044 7.428 2.516 7.46 ;
  LAYER M2 ;
        RECT 0.044 7.492 2.516 7.524 ;
  LAYER M2 ;
        RECT 0.044 7.556 2.516 7.588 ;
  LAYER M2 ;
        RECT 0.044 7.62 2.516 7.652 ;
  LAYER M2 ;
        RECT 0.044 7.684 2.516 7.716 ;
  LAYER M2 ;
        RECT 0.044 7.748 2.516 7.78 ;
  LAYER M2 ;
        RECT 0.044 7.812 2.516 7.844 ;
  LAYER M2 ;
        RECT 0.044 7.876 2.516 7.908 ;
  LAYER M2 ;
        RECT 0.044 7.94 2.516 7.972 ;
  LAYER M2 ;
        RECT 0.044 8.004 2.516 8.036 ;
  LAYER M2 ;
        RECT 0.044 8.068 2.516 8.1 ;
  LAYER M2 ;
        RECT 0.044 8.132 2.516 8.164 ;
  LAYER M2 ;
        RECT 0.044 8.196 2.516 8.228 ;
  LAYER M2 ;
        RECT 0.044 8.26 2.516 8.292 ;
  LAYER M2 ;
        RECT 0.044 8.324 2.516 8.356 ;
  LAYER M2 ;
        RECT 0.044 8.388 2.516 8.42 ;
  LAYER M2 ;
        RECT 0.044 8.452 2.516 8.484 ;
  LAYER M2 ;
        RECT 0.044 8.516 2.516 8.548 ;
  LAYER M2 ;
        RECT 0.044 8.58 2.516 8.612 ;
  LAYER M2 ;
        RECT 0.044 8.644 2.516 8.676 ;
  LAYER M2 ;
        RECT 0.044 8.708 2.516 8.74 ;
  LAYER M2 ;
        RECT 0.044 8.772 2.516 8.804 ;
  LAYER M2 ;
        RECT 0.044 8.836 2.516 8.868 ;
  LAYER M2 ;
        RECT 0.044 8.9 2.516 8.932 ;
  LAYER M2 ;
        RECT 0.044 8.964 2.516 8.996 ;
  LAYER M2 ;
        RECT 0.044 9.028 2.516 9.06 ;
  LAYER M2 ;
        RECT 0.044 9.092 2.516 9.124 ;
  LAYER M3 ;
        RECT 0.064 6.768 0.096 9.276 ;
  LAYER M3 ;
        RECT 0.128 6.768 0.16 9.276 ;
  LAYER M3 ;
        RECT 0.192 6.768 0.224 9.276 ;
  LAYER M3 ;
        RECT 0.256 6.768 0.288 9.276 ;
  LAYER M3 ;
        RECT 0.32 6.768 0.352 9.276 ;
  LAYER M3 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M3 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M3 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M3 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M3 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M3 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M3 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M3 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M3 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M3 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M3 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M3 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M3 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M3 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M3 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M3 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M3 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M3 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M3 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M3 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M3 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M3 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M3 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M3 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M3 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M3 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M3 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M3 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M3 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M3 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M3 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M3 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M3 ;
        RECT 2.464 6.768 2.496 9.276 ;
  LAYER M1 ;
        RECT 0.079 6.804 0.081 9.24 ;
  LAYER M1 ;
        RECT 0.159 6.804 0.161 9.24 ;
  LAYER M1 ;
        RECT 0.239 6.804 0.241 9.24 ;
  LAYER M1 ;
        RECT 0.319 6.804 0.321 9.24 ;
  LAYER M1 ;
        RECT 0.399 6.804 0.401 9.24 ;
  LAYER M1 ;
        RECT 0.479 6.804 0.481 9.24 ;
  LAYER M1 ;
        RECT 0.559 6.804 0.561 9.24 ;
  LAYER M1 ;
        RECT 0.639 6.804 0.641 9.24 ;
  LAYER M1 ;
        RECT 0.719 6.804 0.721 9.24 ;
  LAYER M1 ;
        RECT 0.799 6.804 0.801 9.24 ;
  LAYER M1 ;
        RECT 0.879 6.804 0.881 9.24 ;
  LAYER M1 ;
        RECT 0.959 6.804 0.961 9.24 ;
  LAYER M1 ;
        RECT 1.039 6.804 1.041 9.24 ;
  LAYER M1 ;
        RECT 1.119 6.804 1.121 9.24 ;
  LAYER M1 ;
        RECT 1.199 6.804 1.201 9.24 ;
  LAYER M1 ;
        RECT 1.279 6.804 1.281 9.24 ;
  LAYER M1 ;
        RECT 1.359 6.804 1.361 9.24 ;
  LAYER M1 ;
        RECT 1.439 6.804 1.441 9.24 ;
  LAYER M1 ;
        RECT 1.519 6.804 1.521 9.24 ;
  LAYER M1 ;
        RECT 1.599 6.804 1.601 9.24 ;
  LAYER M1 ;
        RECT 1.679 6.804 1.681 9.24 ;
  LAYER M1 ;
        RECT 1.759 6.804 1.761 9.24 ;
  LAYER M1 ;
        RECT 1.839 6.804 1.841 9.24 ;
  LAYER M1 ;
        RECT 1.919 6.804 1.921 9.24 ;
  LAYER M1 ;
        RECT 1.999 6.804 2.001 9.24 ;
  LAYER M1 ;
        RECT 2.079 6.804 2.081 9.24 ;
  LAYER M1 ;
        RECT 2.159 6.804 2.161 9.24 ;
  LAYER M1 ;
        RECT 2.239 6.804 2.241 9.24 ;
  LAYER M1 ;
        RECT 2.319 6.804 2.321 9.24 ;
  LAYER M1 ;
        RECT 2.399 6.804 2.401 9.24 ;
  LAYER M2 ;
        RECT 0.08 6.803 2.48 6.805 ;
  LAYER M2 ;
        RECT 0.08 6.887 2.48 6.889 ;
  LAYER M2 ;
        RECT 0.08 6.971 2.48 6.973 ;
  LAYER M2 ;
        RECT 0.08 7.055 2.48 7.057 ;
  LAYER M2 ;
        RECT 0.08 7.139 2.48 7.141 ;
  LAYER M2 ;
        RECT 0.08 7.223 2.48 7.225 ;
  LAYER M2 ;
        RECT 0.08 7.307 2.48 7.309 ;
  LAYER M2 ;
        RECT 0.08 7.391 2.48 7.393 ;
  LAYER M2 ;
        RECT 0.08 7.475 2.48 7.477 ;
  LAYER M2 ;
        RECT 0.08 7.559 2.48 7.561 ;
  LAYER M2 ;
        RECT 0.08 7.643 2.48 7.645 ;
  LAYER M2 ;
        RECT 0.08 7.727 2.48 7.729 ;
  LAYER M2 ;
        RECT 0.08 7.8105 2.48 7.8125 ;
  LAYER M2 ;
        RECT 0.08 7.895 2.48 7.897 ;
  LAYER M2 ;
        RECT 0.08 7.979 2.48 7.981 ;
  LAYER M2 ;
        RECT 0.08 8.063 2.48 8.065 ;
  LAYER M2 ;
        RECT 0.08 8.147 2.48 8.149 ;
  LAYER M2 ;
        RECT 0.08 8.231 2.48 8.233 ;
  LAYER M2 ;
        RECT 0.08 8.315 2.48 8.317 ;
  LAYER M2 ;
        RECT 0.08 8.399 2.48 8.401 ;
  LAYER M2 ;
        RECT 0.08 8.483 2.48 8.485 ;
  LAYER M2 ;
        RECT 0.08 8.567 2.48 8.569 ;
  LAYER M2 ;
        RECT 0.08 8.651 2.48 8.653 ;
  LAYER M2 ;
        RECT 0.08 8.735 2.48 8.737 ;
  LAYER M2 ;
        RECT 0.08 8.819 2.48 8.821 ;
  LAYER M2 ;
        RECT 0.08 8.903 2.48 8.905 ;
  LAYER M2 ;
        RECT 0.08 8.987 2.48 8.989 ;
  LAYER M2 ;
        RECT 0.08 9.071 2.48 9.073 ;
  LAYER M2 ;
        RECT 0.08 9.155 2.48 9.157 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 12.216 ;
  LAYER M1 ;
        RECT 0.128 9.708 0.16 12.216 ;
  LAYER M1 ;
        RECT 0.192 9.708 0.224 12.216 ;
  LAYER M1 ;
        RECT 0.256 9.708 0.288 12.216 ;
  LAYER M1 ;
        RECT 0.32 9.708 0.352 12.216 ;
  LAYER M1 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M1 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M1 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M1 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M1 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M1 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M1 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M1 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M1 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M1 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M1 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M1 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M1 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M1 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M1 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M1 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M1 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M1 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M1 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M1 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M1 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M1 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M1 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M1 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M1 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M1 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M1 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M1 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M1 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M1 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M1 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M1 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M2 ;
        RECT 0.044 9.792 2.516 9.824 ;
  LAYER M2 ;
        RECT 0.044 9.856 2.516 9.888 ;
  LAYER M2 ;
        RECT 0.044 9.92 2.516 9.952 ;
  LAYER M2 ;
        RECT 0.044 9.984 2.516 10.016 ;
  LAYER M2 ;
        RECT 0.044 10.048 2.516 10.08 ;
  LAYER M2 ;
        RECT 0.044 10.112 2.516 10.144 ;
  LAYER M2 ;
        RECT 0.044 10.176 2.516 10.208 ;
  LAYER M2 ;
        RECT 0.044 10.24 2.516 10.272 ;
  LAYER M2 ;
        RECT 0.044 10.304 2.516 10.336 ;
  LAYER M2 ;
        RECT 0.044 10.368 2.516 10.4 ;
  LAYER M2 ;
        RECT 0.044 10.432 2.516 10.464 ;
  LAYER M2 ;
        RECT 0.044 10.496 2.516 10.528 ;
  LAYER M2 ;
        RECT 0.044 10.56 2.516 10.592 ;
  LAYER M2 ;
        RECT 0.044 10.624 2.516 10.656 ;
  LAYER M2 ;
        RECT 0.044 10.688 2.516 10.72 ;
  LAYER M2 ;
        RECT 0.044 10.752 2.516 10.784 ;
  LAYER M2 ;
        RECT 0.044 10.816 2.516 10.848 ;
  LAYER M2 ;
        RECT 0.044 10.88 2.516 10.912 ;
  LAYER M2 ;
        RECT 0.044 10.944 2.516 10.976 ;
  LAYER M2 ;
        RECT 0.044 11.008 2.516 11.04 ;
  LAYER M2 ;
        RECT 0.044 11.072 2.516 11.104 ;
  LAYER M2 ;
        RECT 0.044 11.136 2.516 11.168 ;
  LAYER M2 ;
        RECT 0.044 11.2 2.516 11.232 ;
  LAYER M2 ;
        RECT 0.044 11.264 2.516 11.296 ;
  LAYER M2 ;
        RECT 0.044 11.328 2.516 11.36 ;
  LAYER M2 ;
        RECT 0.044 11.392 2.516 11.424 ;
  LAYER M2 ;
        RECT 0.044 11.456 2.516 11.488 ;
  LAYER M2 ;
        RECT 0.044 11.52 2.516 11.552 ;
  LAYER M2 ;
        RECT 0.044 11.584 2.516 11.616 ;
  LAYER M2 ;
        RECT 0.044 11.648 2.516 11.68 ;
  LAYER M2 ;
        RECT 0.044 11.712 2.516 11.744 ;
  LAYER M2 ;
        RECT 0.044 11.776 2.516 11.808 ;
  LAYER M2 ;
        RECT 0.044 11.84 2.516 11.872 ;
  LAYER M2 ;
        RECT 0.044 11.904 2.516 11.936 ;
  LAYER M2 ;
        RECT 0.044 11.968 2.516 12 ;
  LAYER M2 ;
        RECT 0.044 12.032 2.516 12.064 ;
  LAYER M3 ;
        RECT 0.064 9.708 0.096 12.216 ;
  LAYER M3 ;
        RECT 0.128 9.708 0.16 12.216 ;
  LAYER M3 ;
        RECT 0.192 9.708 0.224 12.216 ;
  LAYER M3 ;
        RECT 0.256 9.708 0.288 12.216 ;
  LAYER M3 ;
        RECT 0.32 9.708 0.352 12.216 ;
  LAYER M3 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M3 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M3 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M3 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M3 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M3 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M3 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M3 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M3 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M3 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M3 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M3 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M3 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M3 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M3 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M3 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M3 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M3 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M3 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M3 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M3 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M3 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M3 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M3 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M3 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M3 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M3 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M3 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M3 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M3 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M3 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M3 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M3 ;
        RECT 2.464 9.708 2.496 12.216 ;
  LAYER M1 ;
        RECT 0.079 9.744 0.081 12.18 ;
  LAYER M1 ;
        RECT 0.159 9.744 0.161 12.18 ;
  LAYER M1 ;
        RECT 0.239 9.744 0.241 12.18 ;
  LAYER M1 ;
        RECT 0.319 9.744 0.321 12.18 ;
  LAYER M1 ;
        RECT 0.399 9.744 0.401 12.18 ;
  LAYER M1 ;
        RECT 0.479 9.744 0.481 12.18 ;
  LAYER M1 ;
        RECT 0.559 9.744 0.561 12.18 ;
  LAYER M1 ;
        RECT 0.639 9.744 0.641 12.18 ;
  LAYER M1 ;
        RECT 0.719 9.744 0.721 12.18 ;
  LAYER M1 ;
        RECT 0.799 9.744 0.801 12.18 ;
  LAYER M1 ;
        RECT 0.879 9.744 0.881 12.18 ;
  LAYER M1 ;
        RECT 0.959 9.744 0.961 12.18 ;
  LAYER M1 ;
        RECT 1.039 9.744 1.041 12.18 ;
  LAYER M1 ;
        RECT 1.119 9.744 1.121 12.18 ;
  LAYER M1 ;
        RECT 1.199 9.744 1.201 12.18 ;
  LAYER M1 ;
        RECT 1.279 9.744 1.281 12.18 ;
  LAYER M1 ;
        RECT 1.359 9.744 1.361 12.18 ;
  LAYER M1 ;
        RECT 1.439 9.744 1.441 12.18 ;
  LAYER M1 ;
        RECT 1.519 9.744 1.521 12.18 ;
  LAYER M1 ;
        RECT 1.599 9.744 1.601 12.18 ;
  LAYER M1 ;
        RECT 1.679 9.744 1.681 12.18 ;
  LAYER M1 ;
        RECT 1.759 9.744 1.761 12.18 ;
  LAYER M1 ;
        RECT 1.839 9.744 1.841 12.18 ;
  LAYER M1 ;
        RECT 1.919 9.744 1.921 12.18 ;
  LAYER M1 ;
        RECT 1.999 9.744 2.001 12.18 ;
  LAYER M1 ;
        RECT 2.079 9.744 2.081 12.18 ;
  LAYER M1 ;
        RECT 2.159 9.744 2.161 12.18 ;
  LAYER M1 ;
        RECT 2.239 9.744 2.241 12.18 ;
  LAYER M1 ;
        RECT 2.319 9.744 2.321 12.18 ;
  LAYER M1 ;
        RECT 2.399 9.744 2.401 12.18 ;
  LAYER M2 ;
        RECT 0.08 9.743 2.48 9.745 ;
  LAYER M2 ;
        RECT 0.08 9.827 2.48 9.829 ;
  LAYER M2 ;
        RECT 0.08 9.911 2.48 9.913 ;
  LAYER M2 ;
        RECT 0.08 9.995 2.48 9.997 ;
  LAYER M2 ;
        RECT 0.08 10.079 2.48 10.081 ;
  LAYER M2 ;
        RECT 0.08 10.163 2.48 10.165 ;
  LAYER M2 ;
        RECT 0.08 10.247 2.48 10.249 ;
  LAYER M2 ;
        RECT 0.08 10.331 2.48 10.333 ;
  LAYER M2 ;
        RECT 0.08 10.415 2.48 10.417 ;
  LAYER M2 ;
        RECT 0.08 10.499 2.48 10.501 ;
  LAYER M2 ;
        RECT 0.08 10.583 2.48 10.585 ;
  LAYER M2 ;
        RECT 0.08 10.667 2.48 10.669 ;
  LAYER M2 ;
        RECT 0.08 10.7505 2.48 10.7525 ;
  LAYER M2 ;
        RECT 0.08 10.835 2.48 10.837 ;
  LAYER M2 ;
        RECT 0.08 10.919 2.48 10.921 ;
  LAYER M2 ;
        RECT 0.08 11.003 2.48 11.005 ;
  LAYER M2 ;
        RECT 0.08 11.087 2.48 11.089 ;
  LAYER M2 ;
        RECT 0.08 11.171 2.48 11.173 ;
  LAYER M2 ;
        RECT 0.08 11.255 2.48 11.257 ;
  LAYER M2 ;
        RECT 0.08 11.339 2.48 11.341 ;
  LAYER M2 ;
        RECT 0.08 11.423 2.48 11.425 ;
  LAYER M2 ;
        RECT 0.08 11.507 2.48 11.509 ;
  LAYER M2 ;
        RECT 0.08 11.591 2.48 11.593 ;
  LAYER M2 ;
        RECT 0.08 11.675 2.48 11.677 ;
  LAYER M2 ;
        RECT 0.08 11.759 2.48 11.761 ;
  LAYER M2 ;
        RECT 0.08 11.843 2.48 11.845 ;
  LAYER M2 ;
        RECT 0.08 11.927 2.48 11.929 ;
  LAYER M2 ;
        RECT 0.08 12.011 2.48 12.013 ;
  LAYER M2 ;
        RECT 0.08 12.095 2.48 12.097 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 15.156 ;
  LAYER M1 ;
        RECT 0.128 12.648 0.16 15.156 ;
  LAYER M1 ;
        RECT 0.192 12.648 0.224 15.156 ;
  LAYER M1 ;
        RECT 0.256 12.648 0.288 15.156 ;
  LAYER M1 ;
        RECT 0.32 12.648 0.352 15.156 ;
  LAYER M1 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M1 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M1 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M1 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M1 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M1 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M1 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M1 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M1 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M1 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M1 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M1 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M1 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M1 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M1 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M1 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M1 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M1 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M1 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M1 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M1 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M1 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M1 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M1 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M1 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M1 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M1 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M1 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M1 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M1 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M1 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M1 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M2 ;
        RECT 0.044 12.732 2.516 12.764 ;
  LAYER M2 ;
        RECT 0.044 12.796 2.516 12.828 ;
  LAYER M2 ;
        RECT 0.044 12.86 2.516 12.892 ;
  LAYER M2 ;
        RECT 0.044 12.924 2.516 12.956 ;
  LAYER M2 ;
        RECT 0.044 12.988 2.516 13.02 ;
  LAYER M2 ;
        RECT 0.044 13.052 2.516 13.084 ;
  LAYER M2 ;
        RECT 0.044 13.116 2.516 13.148 ;
  LAYER M2 ;
        RECT 0.044 13.18 2.516 13.212 ;
  LAYER M2 ;
        RECT 0.044 13.244 2.516 13.276 ;
  LAYER M2 ;
        RECT 0.044 13.308 2.516 13.34 ;
  LAYER M2 ;
        RECT 0.044 13.372 2.516 13.404 ;
  LAYER M2 ;
        RECT 0.044 13.436 2.516 13.468 ;
  LAYER M2 ;
        RECT 0.044 13.5 2.516 13.532 ;
  LAYER M2 ;
        RECT 0.044 13.564 2.516 13.596 ;
  LAYER M2 ;
        RECT 0.044 13.628 2.516 13.66 ;
  LAYER M2 ;
        RECT 0.044 13.692 2.516 13.724 ;
  LAYER M2 ;
        RECT 0.044 13.756 2.516 13.788 ;
  LAYER M2 ;
        RECT 0.044 13.82 2.516 13.852 ;
  LAYER M2 ;
        RECT 0.044 13.884 2.516 13.916 ;
  LAYER M2 ;
        RECT 0.044 13.948 2.516 13.98 ;
  LAYER M2 ;
        RECT 0.044 14.012 2.516 14.044 ;
  LAYER M2 ;
        RECT 0.044 14.076 2.516 14.108 ;
  LAYER M2 ;
        RECT 0.044 14.14 2.516 14.172 ;
  LAYER M2 ;
        RECT 0.044 14.204 2.516 14.236 ;
  LAYER M2 ;
        RECT 0.044 14.268 2.516 14.3 ;
  LAYER M2 ;
        RECT 0.044 14.332 2.516 14.364 ;
  LAYER M2 ;
        RECT 0.044 14.396 2.516 14.428 ;
  LAYER M2 ;
        RECT 0.044 14.46 2.516 14.492 ;
  LAYER M2 ;
        RECT 0.044 14.524 2.516 14.556 ;
  LAYER M2 ;
        RECT 0.044 14.588 2.516 14.62 ;
  LAYER M2 ;
        RECT 0.044 14.652 2.516 14.684 ;
  LAYER M2 ;
        RECT 0.044 14.716 2.516 14.748 ;
  LAYER M2 ;
        RECT 0.044 14.78 2.516 14.812 ;
  LAYER M2 ;
        RECT 0.044 14.844 2.516 14.876 ;
  LAYER M2 ;
        RECT 0.044 14.908 2.516 14.94 ;
  LAYER M2 ;
        RECT 0.044 14.972 2.516 15.004 ;
  LAYER M3 ;
        RECT 0.064 12.648 0.096 15.156 ;
  LAYER M3 ;
        RECT 0.128 12.648 0.16 15.156 ;
  LAYER M3 ;
        RECT 0.192 12.648 0.224 15.156 ;
  LAYER M3 ;
        RECT 0.256 12.648 0.288 15.156 ;
  LAYER M3 ;
        RECT 0.32 12.648 0.352 15.156 ;
  LAYER M3 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M3 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M3 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M3 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M3 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M3 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M3 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M3 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M3 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M3 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M3 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M3 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M3 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M3 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M3 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M3 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M3 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M3 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M3 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M3 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M3 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M3 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M3 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M3 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M3 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M3 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M3 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M3 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M3 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M3 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M3 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M3 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M3 ;
        RECT 2.464 12.648 2.496 15.156 ;
  LAYER M1 ;
        RECT 0.079 12.684 0.081 15.12 ;
  LAYER M1 ;
        RECT 0.159 12.684 0.161 15.12 ;
  LAYER M1 ;
        RECT 0.239 12.684 0.241 15.12 ;
  LAYER M1 ;
        RECT 0.319 12.684 0.321 15.12 ;
  LAYER M1 ;
        RECT 0.399 12.684 0.401 15.12 ;
  LAYER M1 ;
        RECT 0.479 12.684 0.481 15.12 ;
  LAYER M1 ;
        RECT 0.559 12.684 0.561 15.12 ;
  LAYER M1 ;
        RECT 0.639 12.684 0.641 15.12 ;
  LAYER M1 ;
        RECT 0.719 12.684 0.721 15.12 ;
  LAYER M1 ;
        RECT 0.799 12.684 0.801 15.12 ;
  LAYER M1 ;
        RECT 0.879 12.684 0.881 15.12 ;
  LAYER M1 ;
        RECT 0.959 12.684 0.961 15.12 ;
  LAYER M1 ;
        RECT 1.039 12.684 1.041 15.12 ;
  LAYER M1 ;
        RECT 1.119 12.684 1.121 15.12 ;
  LAYER M1 ;
        RECT 1.199 12.684 1.201 15.12 ;
  LAYER M1 ;
        RECT 1.279 12.684 1.281 15.12 ;
  LAYER M1 ;
        RECT 1.359 12.684 1.361 15.12 ;
  LAYER M1 ;
        RECT 1.439 12.684 1.441 15.12 ;
  LAYER M1 ;
        RECT 1.519 12.684 1.521 15.12 ;
  LAYER M1 ;
        RECT 1.599 12.684 1.601 15.12 ;
  LAYER M1 ;
        RECT 1.679 12.684 1.681 15.12 ;
  LAYER M1 ;
        RECT 1.759 12.684 1.761 15.12 ;
  LAYER M1 ;
        RECT 1.839 12.684 1.841 15.12 ;
  LAYER M1 ;
        RECT 1.919 12.684 1.921 15.12 ;
  LAYER M1 ;
        RECT 1.999 12.684 2.001 15.12 ;
  LAYER M1 ;
        RECT 2.079 12.684 2.081 15.12 ;
  LAYER M1 ;
        RECT 2.159 12.684 2.161 15.12 ;
  LAYER M1 ;
        RECT 2.239 12.684 2.241 15.12 ;
  LAYER M1 ;
        RECT 2.319 12.684 2.321 15.12 ;
  LAYER M1 ;
        RECT 2.399 12.684 2.401 15.12 ;
  LAYER M2 ;
        RECT 0.08 12.683 2.48 12.685 ;
  LAYER M2 ;
        RECT 0.08 12.767 2.48 12.769 ;
  LAYER M2 ;
        RECT 0.08 12.851 2.48 12.853 ;
  LAYER M2 ;
        RECT 0.08 12.935 2.48 12.937 ;
  LAYER M2 ;
        RECT 0.08 13.019 2.48 13.021 ;
  LAYER M2 ;
        RECT 0.08 13.103 2.48 13.105 ;
  LAYER M2 ;
        RECT 0.08 13.187 2.48 13.189 ;
  LAYER M2 ;
        RECT 0.08 13.271 2.48 13.273 ;
  LAYER M2 ;
        RECT 0.08 13.355 2.48 13.357 ;
  LAYER M2 ;
        RECT 0.08 13.439 2.48 13.441 ;
  LAYER M2 ;
        RECT 0.08 13.523 2.48 13.525 ;
  LAYER M2 ;
        RECT 0.08 13.607 2.48 13.609 ;
  LAYER M2 ;
        RECT 0.08 13.6905 2.48 13.6925 ;
  LAYER M2 ;
        RECT 0.08 13.775 2.48 13.777 ;
  LAYER M2 ;
        RECT 0.08 13.859 2.48 13.861 ;
  LAYER M2 ;
        RECT 0.08 13.943 2.48 13.945 ;
  LAYER M2 ;
        RECT 0.08 14.027 2.48 14.029 ;
  LAYER M2 ;
        RECT 0.08 14.111 2.48 14.113 ;
  LAYER M2 ;
        RECT 0.08 14.195 2.48 14.197 ;
  LAYER M2 ;
        RECT 0.08 14.279 2.48 14.281 ;
  LAYER M2 ;
        RECT 0.08 14.363 2.48 14.365 ;
  LAYER M2 ;
        RECT 0.08 14.447 2.48 14.449 ;
  LAYER M2 ;
        RECT 0.08 14.531 2.48 14.533 ;
  LAYER M2 ;
        RECT 0.08 14.615 2.48 14.617 ;
  LAYER M2 ;
        RECT 0.08 14.699 2.48 14.701 ;
  LAYER M2 ;
        RECT 0.08 14.783 2.48 14.785 ;
  LAYER M2 ;
        RECT 0.08 14.867 2.48 14.869 ;
  LAYER M2 ;
        RECT 0.08 14.951 2.48 14.953 ;
  LAYER M2 ;
        RECT 0.08 15.035 2.48 15.037 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 18.096 ;
  LAYER M1 ;
        RECT 0.128 15.588 0.16 18.096 ;
  LAYER M1 ;
        RECT 0.192 15.588 0.224 18.096 ;
  LAYER M1 ;
        RECT 0.256 15.588 0.288 18.096 ;
  LAYER M1 ;
        RECT 0.32 15.588 0.352 18.096 ;
  LAYER M1 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M1 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M1 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M1 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M1 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M1 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M1 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M1 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M1 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M1 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M1 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M1 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M1 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M1 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M1 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M1 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M1 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M1 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M1 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M1 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M1 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M1 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M1 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M1 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M1 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M1 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M1 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M1 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M1 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M1 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M1 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M1 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M2 ;
        RECT 0.044 15.672 2.516 15.704 ;
  LAYER M2 ;
        RECT 0.044 15.736 2.516 15.768 ;
  LAYER M2 ;
        RECT 0.044 15.8 2.516 15.832 ;
  LAYER M2 ;
        RECT 0.044 15.864 2.516 15.896 ;
  LAYER M2 ;
        RECT 0.044 15.928 2.516 15.96 ;
  LAYER M2 ;
        RECT 0.044 15.992 2.516 16.024 ;
  LAYER M2 ;
        RECT 0.044 16.056 2.516 16.088 ;
  LAYER M2 ;
        RECT 0.044 16.12 2.516 16.152 ;
  LAYER M2 ;
        RECT 0.044 16.184 2.516 16.216 ;
  LAYER M2 ;
        RECT 0.044 16.248 2.516 16.28 ;
  LAYER M2 ;
        RECT 0.044 16.312 2.516 16.344 ;
  LAYER M2 ;
        RECT 0.044 16.376 2.516 16.408 ;
  LAYER M2 ;
        RECT 0.044 16.44 2.516 16.472 ;
  LAYER M2 ;
        RECT 0.044 16.504 2.516 16.536 ;
  LAYER M2 ;
        RECT 0.044 16.568 2.516 16.6 ;
  LAYER M2 ;
        RECT 0.044 16.632 2.516 16.664 ;
  LAYER M2 ;
        RECT 0.044 16.696 2.516 16.728 ;
  LAYER M2 ;
        RECT 0.044 16.76 2.516 16.792 ;
  LAYER M2 ;
        RECT 0.044 16.824 2.516 16.856 ;
  LAYER M2 ;
        RECT 0.044 16.888 2.516 16.92 ;
  LAYER M2 ;
        RECT 0.044 16.952 2.516 16.984 ;
  LAYER M2 ;
        RECT 0.044 17.016 2.516 17.048 ;
  LAYER M2 ;
        RECT 0.044 17.08 2.516 17.112 ;
  LAYER M2 ;
        RECT 0.044 17.144 2.516 17.176 ;
  LAYER M2 ;
        RECT 0.044 17.208 2.516 17.24 ;
  LAYER M2 ;
        RECT 0.044 17.272 2.516 17.304 ;
  LAYER M2 ;
        RECT 0.044 17.336 2.516 17.368 ;
  LAYER M2 ;
        RECT 0.044 17.4 2.516 17.432 ;
  LAYER M2 ;
        RECT 0.044 17.464 2.516 17.496 ;
  LAYER M2 ;
        RECT 0.044 17.528 2.516 17.56 ;
  LAYER M2 ;
        RECT 0.044 17.592 2.516 17.624 ;
  LAYER M2 ;
        RECT 0.044 17.656 2.516 17.688 ;
  LAYER M2 ;
        RECT 0.044 17.72 2.516 17.752 ;
  LAYER M2 ;
        RECT 0.044 17.784 2.516 17.816 ;
  LAYER M2 ;
        RECT 0.044 17.848 2.516 17.88 ;
  LAYER M2 ;
        RECT 0.044 17.912 2.516 17.944 ;
  LAYER M3 ;
        RECT 0.064 15.588 0.096 18.096 ;
  LAYER M3 ;
        RECT 0.128 15.588 0.16 18.096 ;
  LAYER M3 ;
        RECT 0.192 15.588 0.224 18.096 ;
  LAYER M3 ;
        RECT 0.256 15.588 0.288 18.096 ;
  LAYER M3 ;
        RECT 0.32 15.588 0.352 18.096 ;
  LAYER M3 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M3 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M3 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M3 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M3 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M3 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M3 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M3 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M3 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M3 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M3 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M3 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M3 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M3 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M3 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M3 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M3 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M3 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M3 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M3 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M3 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M3 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M3 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M3 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M3 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M3 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M3 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M3 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M3 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M3 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M3 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M3 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M3 ;
        RECT 2.464 15.588 2.496 18.096 ;
  LAYER M1 ;
        RECT 0.079 15.624 0.081 18.06 ;
  LAYER M1 ;
        RECT 0.159 15.624 0.161 18.06 ;
  LAYER M1 ;
        RECT 0.239 15.624 0.241 18.06 ;
  LAYER M1 ;
        RECT 0.319 15.624 0.321 18.06 ;
  LAYER M1 ;
        RECT 0.399 15.624 0.401 18.06 ;
  LAYER M1 ;
        RECT 0.479 15.624 0.481 18.06 ;
  LAYER M1 ;
        RECT 0.559 15.624 0.561 18.06 ;
  LAYER M1 ;
        RECT 0.639 15.624 0.641 18.06 ;
  LAYER M1 ;
        RECT 0.719 15.624 0.721 18.06 ;
  LAYER M1 ;
        RECT 0.799 15.624 0.801 18.06 ;
  LAYER M1 ;
        RECT 0.879 15.624 0.881 18.06 ;
  LAYER M1 ;
        RECT 0.959 15.624 0.961 18.06 ;
  LAYER M1 ;
        RECT 1.039 15.624 1.041 18.06 ;
  LAYER M1 ;
        RECT 1.119 15.624 1.121 18.06 ;
  LAYER M1 ;
        RECT 1.199 15.624 1.201 18.06 ;
  LAYER M1 ;
        RECT 1.279 15.624 1.281 18.06 ;
  LAYER M1 ;
        RECT 1.359 15.624 1.361 18.06 ;
  LAYER M1 ;
        RECT 1.439 15.624 1.441 18.06 ;
  LAYER M1 ;
        RECT 1.519 15.624 1.521 18.06 ;
  LAYER M1 ;
        RECT 1.599 15.624 1.601 18.06 ;
  LAYER M1 ;
        RECT 1.679 15.624 1.681 18.06 ;
  LAYER M1 ;
        RECT 1.759 15.624 1.761 18.06 ;
  LAYER M1 ;
        RECT 1.839 15.624 1.841 18.06 ;
  LAYER M1 ;
        RECT 1.919 15.624 1.921 18.06 ;
  LAYER M1 ;
        RECT 1.999 15.624 2.001 18.06 ;
  LAYER M1 ;
        RECT 2.079 15.624 2.081 18.06 ;
  LAYER M1 ;
        RECT 2.159 15.624 2.161 18.06 ;
  LAYER M1 ;
        RECT 2.239 15.624 2.241 18.06 ;
  LAYER M1 ;
        RECT 2.319 15.624 2.321 18.06 ;
  LAYER M1 ;
        RECT 2.399 15.624 2.401 18.06 ;
  LAYER M2 ;
        RECT 0.08 15.623 2.48 15.625 ;
  LAYER M2 ;
        RECT 0.08 15.707 2.48 15.709 ;
  LAYER M2 ;
        RECT 0.08 15.791 2.48 15.793 ;
  LAYER M2 ;
        RECT 0.08 15.875 2.48 15.877 ;
  LAYER M2 ;
        RECT 0.08 15.959 2.48 15.961 ;
  LAYER M2 ;
        RECT 0.08 16.043 2.48 16.045 ;
  LAYER M2 ;
        RECT 0.08 16.127 2.48 16.129 ;
  LAYER M2 ;
        RECT 0.08 16.211 2.48 16.213 ;
  LAYER M2 ;
        RECT 0.08 16.295 2.48 16.297 ;
  LAYER M2 ;
        RECT 0.08 16.379 2.48 16.381 ;
  LAYER M2 ;
        RECT 0.08 16.463 2.48 16.465 ;
  LAYER M2 ;
        RECT 0.08 16.547 2.48 16.549 ;
  LAYER M2 ;
        RECT 0.08 16.6305 2.48 16.6325 ;
  LAYER M2 ;
        RECT 0.08 16.715 2.48 16.717 ;
  LAYER M2 ;
        RECT 0.08 16.799 2.48 16.801 ;
  LAYER M2 ;
        RECT 0.08 16.883 2.48 16.885 ;
  LAYER M2 ;
        RECT 0.08 16.967 2.48 16.969 ;
  LAYER M2 ;
        RECT 0.08 17.051 2.48 17.053 ;
  LAYER M2 ;
        RECT 0.08 17.135 2.48 17.137 ;
  LAYER M2 ;
        RECT 0.08 17.219 2.48 17.221 ;
  LAYER M2 ;
        RECT 0.08 17.303 2.48 17.305 ;
  LAYER M2 ;
        RECT 0.08 17.387 2.48 17.389 ;
  LAYER M2 ;
        RECT 0.08 17.471 2.48 17.473 ;
  LAYER M2 ;
        RECT 0.08 17.555 2.48 17.557 ;
  LAYER M2 ;
        RECT 0.08 17.639 2.48 17.641 ;
  LAYER M2 ;
        RECT 0.08 17.723 2.48 17.725 ;
  LAYER M2 ;
        RECT 0.08 17.807 2.48 17.809 ;
  LAYER M2 ;
        RECT 0.08 17.891 2.48 17.893 ;
  LAYER M2 ;
        RECT 0.08 17.975 2.48 17.977 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 21.036 ;
  LAYER M1 ;
        RECT 0.128 18.528 0.16 21.036 ;
  LAYER M1 ;
        RECT 0.192 18.528 0.224 21.036 ;
  LAYER M1 ;
        RECT 0.256 18.528 0.288 21.036 ;
  LAYER M1 ;
        RECT 0.32 18.528 0.352 21.036 ;
  LAYER M1 ;
        RECT 0.384 18.528 0.416 21.036 ;
  LAYER M1 ;
        RECT 0.448 18.528 0.48 21.036 ;
  LAYER M1 ;
        RECT 0.512 18.528 0.544 21.036 ;
  LAYER M1 ;
        RECT 0.576 18.528 0.608 21.036 ;
  LAYER M1 ;
        RECT 0.64 18.528 0.672 21.036 ;
  LAYER M1 ;
        RECT 0.704 18.528 0.736 21.036 ;
  LAYER M1 ;
        RECT 0.768 18.528 0.8 21.036 ;
  LAYER M1 ;
        RECT 0.832 18.528 0.864 21.036 ;
  LAYER M1 ;
        RECT 0.896 18.528 0.928 21.036 ;
  LAYER M1 ;
        RECT 0.96 18.528 0.992 21.036 ;
  LAYER M1 ;
        RECT 1.024 18.528 1.056 21.036 ;
  LAYER M1 ;
        RECT 1.088 18.528 1.12 21.036 ;
  LAYER M1 ;
        RECT 1.152 18.528 1.184 21.036 ;
  LAYER M1 ;
        RECT 1.216 18.528 1.248 21.036 ;
  LAYER M1 ;
        RECT 1.28 18.528 1.312 21.036 ;
  LAYER M1 ;
        RECT 1.344 18.528 1.376 21.036 ;
  LAYER M1 ;
        RECT 1.408 18.528 1.44 21.036 ;
  LAYER M1 ;
        RECT 1.472 18.528 1.504 21.036 ;
  LAYER M1 ;
        RECT 1.536 18.528 1.568 21.036 ;
  LAYER M1 ;
        RECT 1.6 18.528 1.632 21.036 ;
  LAYER M1 ;
        RECT 1.664 18.528 1.696 21.036 ;
  LAYER M1 ;
        RECT 1.728 18.528 1.76 21.036 ;
  LAYER M1 ;
        RECT 1.792 18.528 1.824 21.036 ;
  LAYER M1 ;
        RECT 1.856 18.528 1.888 21.036 ;
  LAYER M1 ;
        RECT 1.92 18.528 1.952 21.036 ;
  LAYER M1 ;
        RECT 1.984 18.528 2.016 21.036 ;
  LAYER M1 ;
        RECT 2.048 18.528 2.08 21.036 ;
  LAYER M1 ;
        RECT 2.112 18.528 2.144 21.036 ;
  LAYER M1 ;
        RECT 2.176 18.528 2.208 21.036 ;
  LAYER M1 ;
        RECT 2.24 18.528 2.272 21.036 ;
  LAYER M1 ;
        RECT 2.304 18.528 2.336 21.036 ;
  LAYER M1 ;
        RECT 2.368 18.528 2.4 21.036 ;
  LAYER M2 ;
        RECT 0.044 18.612 2.516 18.644 ;
  LAYER M2 ;
        RECT 0.044 18.676 2.516 18.708 ;
  LAYER M2 ;
        RECT 0.044 18.74 2.516 18.772 ;
  LAYER M2 ;
        RECT 0.044 18.804 2.516 18.836 ;
  LAYER M2 ;
        RECT 0.044 18.868 2.516 18.9 ;
  LAYER M2 ;
        RECT 0.044 18.932 2.516 18.964 ;
  LAYER M2 ;
        RECT 0.044 18.996 2.516 19.028 ;
  LAYER M2 ;
        RECT 0.044 19.06 2.516 19.092 ;
  LAYER M2 ;
        RECT 0.044 19.124 2.516 19.156 ;
  LAYER M2 ;
        RECT 0.044 19.188 2.516 19.22 ;
  LAYER M2 ;
        RECT 0.044 19.252 2.516 19.284 ;
  LAYER M2 ;
        RECT 0.044 19.316 2.516 19.348 ;
  LAYER M2 ;
        RECT 0.044 19.38 2.516 19.412 ;
  LAYER M2 ;
        RECT 0.044 19.444 2.516 19.476 ;
  LAYER M2 ;
        RECT 0.044 19.508 2.516 19.54 ;
  LAYER M2 ;
        RECT 0.044 19.572 2.516 19.604 ;
  LAYER M2 ;
        RECT 0.044 19.636 2.516 19.668 ;
  LAYER M2 ;
        RECT 0.044 19.7 2.516 19.732 ;
  LAYER M2 ;
        RECT 0.044 19.764 2.516 19.796 ;
  LAYER M2 ;
        RECT 0.044 19.828 2.516 19.86 ;
  LAYER M2 ;
        RECT 0.044 19.892 2.516 19.924 ;
  LAYER M2 ;
        RECT 0.044 19.956 2.516 19.988 ;
  LAYER M2 ;
        RECT 0.044 20.02 2.516 20.052 ;
  LAYER M2 ;
        RECT 0.044 20.084 2.516 20.116 ;
  LAYER M2 ;
        RECT 0.044 20.148 2.516 20.18 ;
  LAYER M2 ;
        RECT 0.044 20.212 2.516 20.244 ;
  LAYER M2 ;
        RECT 0.044 20.276 2.516 20.308 ;
  LAYER M2 ;
        RECT 0.044 20.34 2.516 20.372 ;
  LAYER M2 ;
        RECT 0.044 20.404 2.516 20.436 ;
  LAYER M2 ;
        RECT 0.044 20.468 2.516 20.5 ;
  LAYER M2 ;
        RECT 0.044 20.532 2.516 20.564 ;
  LAYER M2 ;
        RECT 0.044 20.596 2.516 20.628 ;
  LAYER M2 ;
        RECT 0.044 20.66 2.516 20.692 ;
  LAYER M2 ;
        RECT 0.044 20.724 2.516 20.756 ;
  LAYER M2 ;
        RECT 0.044 20.788 2.516 20.82 ;
  LAYER M2 ;
        RECT 0.044 20.852 2.516 20.884 ;
  LAYER M3 ;
        RECT 0.064 18.528 0.096 21.036 ;
  LAYER M3 ;
        RECT 0.128 18.528 0.16 21.036 ;
  LAYER M3 ;
        RECT 0.192 18.528 0.224 21.036 ;
  LAYER M3 ;
        RECT 0.256 18.528 0.288 21.036 ;
  LAYER M3 ;
        RECT 0.32 18.528 0.352 21.036 ;
  LAYER M3 ;
        RECT 0.384 18.528 0.416 21.036 ;
  LAYER M3 ;
        RECT 0.448 18.528 0.48 21.036 ;
  LAYER M3 ;
        RECT 0.512 18.528 0.544 21.036 ;
  LAYER M3 ;
        RECT 0.576 18.528 0.608 21.036 ;
  LAYER M3 ;
        RECT 0.64 18.528 0.672 21.036 ;
  LAYER M3 ;
        RECT 0.704 18.528 0.736 21.036 ;
  LAYER M3 ;
        RECT 0.768 18.528 0.8 21.036 ;
  LAYER M3 ;
        RECT 0.832 18.528 0.864 21.036 ;
  LAYER M3 ;
        RECT 0.896 18.528 0.928 21.036 ;
  LAYER M3 ;
        RECT 0.96 18.528 0.992 21.036 ;
  LAYER M3 ;
        RECT 1.024 18.528 1.056 21.036 ;
  LAYER M3 ;
        RECT 1.088 18.528 1.12 21.036 ;
  LAYER M3 ;
        RECT 1.152 18.528 1.184 21.036 ;
  LAYER M3 ;
        RECT 1.216 18.528 1.248 21.036 ;
  LAYER M3 ;
        RECT 1.28 18.528 1.312 21.036 ;
  LAYER M3 ;
        RECT 1.344 18.528 1.376 21.036 ;
  LAYER M3 ;
        RECT 1.408 18.528 1.44 21.036 ;
  LAYER M3 ;
        RECT 1.472 18.528 1.504 21.036 ;
  LAYER M3 ;
        RECT 1.536 18.528 1.568 21.036 ;
  LAYER M3 ;
        RECT 1.6 18.528 1.632 21.036 ;
  LAYER M3 ;
        RECT 1.664 18.528 1.696 21.036 ;
  LAYER M3 ;
        RECT 1.728 18.528 1.76 21.036 ;
  LAYER M3 ;
        RECT 1.792 18.528 1.824 21.036 ;
  LAYER M3 ;
        RECT 1.856 18.528 1.888 21.036 ;
  LAYER M3 ;
        RECT 1.92 18.528 1.952 21.036 ;
  LAYER M3 ;
        RECT 1.984 18.528 2.016 21.036 ;
  LAYER M3 ;
        RECT 2.048 18.528 2.08 21.036 ;
  LAYER M3 ;
        RECT 2.112 18.528 2.144 21.036 ;
  LAYER M3 ;
        RECT 2.176 18.528 2.208 21.036 ;
  LAYER M3 ;
        RECT 2.24 18.528 2.272 21.036 ;
  LAYER M3 ;
        RECT 2.304 18.528 2.336 21.036 ;
  LAYER M3 ;
        RECT 2.368 18.528 2.4 21.036 ;
  LAYER M3 ;
        RECT 2.464 18.528 2.496 21.036 ;
  LAYER M1 ;
        RECT 0.079 18.564 0.081 21 ;
  LAYER M1 ;
        RECT 0.159 18.564 0.161 21 ;
  LAYER M1 ;
        RECT 0.239 18.564 0.241 21 ;
  LAYER M1 ;
        RECT 0.319 18.564 0.321 21 ;
  LAYER M1 ;
        RECT 0.399 18.564 0.401 21 ;
  LAYER M1 ;
        RECT 0.479 18.564 0.481 21 ;
  LAYER M1 ;
        RECT 0.559 18.564 0.561 21 ;
  LAYER M1 ;
        RECT 0.639 18.564 0.641 21 ;
  LAYER M1 ;
        RECT 0.719 18.564 0.721 21 ;
  LAYER M1 ;
        RECT 0.799 18.564 0.801 21 ;
  LAYER M1 ;
        RECT 0.879 18.564 0.881 21 ;
  LAYER M1 ;
        RECT 0.959 18.564 0.961 21 ;
  LAYER M1 ;
        RECT 1.039 18.564 1.041 21 ;
  LAYER M1 ;
        RECT 1.119 18.564 1.121 21 ;
  LAYER M1 ;
        RECT 1.199 18.564 1.201 21 ;
  LAYER M1 ;
        RECT 1.279 18.564 1.281 21 ;
  LAYER M1 ;
        RECT 1.359 18.564 1.361 21 ;
  LAYER M1 ;
        RECT 1.439 18.564 1.441 21 ;
  LAYER M1 ;
        RECT 1.519 18.564 1.521 21 ;
  LAYER M1 ;
        RECT 1.599 18.564 1.601 21 ;
  LAYER M1 ;
        RECT 1.679 18.564 1.681 21 ;
  LAYER M1 ;
        RECT 1.759 18.564 1.761 21 ;
  LAYER M1 ;
        RECT 1.839 18.564 1.841 21 ;
  LAYER M1 ;
        RECT 1.919 18.564 1.921 21 ;
  LAYER M1 ;
        RECT 1.999 18.564 2.001 21 ;
  LAYER M1 ;
        RECT 2.079 18.564 2.081 21 ;
  LAYER M1 ;
        RECT 2.159 18.564 2.161 21 ;
  LAYER M1 ;
        RECT 2.239 18.564 2.241 21 ;
  LAYER M1 ;
        RECT 2.319 18.564 2.321 21 ;
  LAYER M1 ;
        RECT 2.399 18.564 2.401 21 ;
  LAYER M2 ;
        RECT 0.08 18.563 2.48 18.565 ;
  LAYER M2 ;
        RECT 0.08 18.647 2.48 18.649 ;
  LAYER M2 ;
        RECT 0.08 18.731 2.48 18.733 ;
  LAYER M2 ;
        RECT 0.08 18.815 2.48 18.817 ;
  LAYER M2 ;
        RECT 0.08 18.899 2.48 18.901 ;
  LAYER M2 ;
        RECT 0.08 18.983 2.48 18.985 ;
  LAYER M2 ;
        RECT 0.08 19.067 2.48 19.069 ;
  LAYER M2 ;
        RECT 0.08 19.151 2.48 19.153 ;
  LAYER M2 ;
        RECT 0.08 19.235 2.48 19.237 ;
  LAYER M2 ;
        RECT 0.08 19.319 2.48 19.321 ;
  LAYER M2 ;
        RECT 0.08 19.403 2.48 19.405 ;
  LAYER M2 ;
        RECT 0.08 19.487 2.48 19.489 ;
  LAYER M2 ;
        RECT 0.08 19.5705 2.48 19.5725 ;
  LAYER M2 ;
        RECT 0.08 19.655 2.48 19.657 ;
  LAYER M2 ;
        RECT 0.08 19.739 2.48 19.741 ;
  LAYER M2 ;
        RECT 0.08 19.823 2.48 19.825 ;
  LAYER M2 ;
        RECT 0.08 19.907 2.48 19.909 ;
  LAYER M2 ;
        RECT 0.08 19.991 2.48 19.993 ;
  LAYER M2 ;
        RECT 0.08 20.075 2.48 20.077 ;
  LAYER M2 ;
        RECT 0.08 20.159 2.48 20.161 ;
  LAYER M2 ;
        RECT 0.08 20.243 2.48 20.245 ;
  LAYER M2 ;
        RECT 0.08 20.327 2.48 20.329 ;
  LAYER M2 ;
        RECT 0.08 20.411 2.48 20.413 ;
  LAYER M2 ;
        RECT 0.08 20.495 2.48 20.497 ;
  LAYER M2 ;
        RECT 0.08 20.579 2.48 20.581 ;
  LAYER M2 ;
        RECT 0.08 20.663 2.48 20.665 ;
  LAYER M2 ;
        RECT 0.08 20.747 2.48 20.749 ;
  LAYER M2 ;
        RECT 0.08 20.831 2.48 20.833 ;
  LAYER M2 ;
        RECT 0.08 20.915 2.48 20.917 ;
  LAYER M1 ;
        RECT 3.264 0.888 3.296 3.396 ;
  LAYER M1 ;
        RECT 3.328 0.888 3.36 3.396 ;
  LAYER M1 ;
        RECT 3.392 0.888 3.424 3.396 ;
  LAYER M1 ;
        RECT 3.456 0.888 3.488 3.396 ;
  LAYER M1 ;
        RECT 3.52 0.888 3.552 3.396 ;
  LAYER M1 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M1 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M1 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M1 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M1 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M1 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M1 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M1 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M1 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M1 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M1 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M1 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M1 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M1 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M1 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M1 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M1 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M1 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M1 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M1 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M1 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M1 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M1 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M1 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M1 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M1 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M1 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M1 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M1 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M1 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M1 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M1 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M2 ;
        RECT 3.244 0.972 5.716 1.004 ;
  LAYER M2 ;
        RECT 3.244 1.036 5.716 1.068 ;
  LAYER M2 ;
        RECT 3.244 1.1 5.716 1.132 ;
  LAYER M2 ;
        RECT 3.244 1.164 5.716 1.196 ;
  LAYER M2 ;
        RECT 3.244 1.228 5.716 1.26 ;
  LAYER M2 ;
        RECT 3.244 1.292 5.716 1.324 ;
  LAYER M2 ;
        RECT 3.244 1.356 5.716 1.388 ;
  LAYER M2 ;
        RECT 3.244 1.42 5.716 1.452 ;
  LAYER M2 ;
        RECT 3.244 1.484 5.716 1.516 ;
  LAYER M2 ;
        RECT 3.244 1.548 5.716 1.58 ;
  LAYER M2 ;
        RECT 3.244 1.612 5.716 1.644 ;
  LAYER M2 ;
        RECT 3.244 1.676 5.716 1.708 ;
  LAYER M2 ;
        RECT 3.244 1.74 5.716 1.772 ;
  LAYER M2 ;
        RECT 3.244 1.804 5.716 1.836 ;
  LAYER M2 ;
        RECT 3.244 1.868 5.716 1.9 ;
  LAYER M2 ;
        RECT 3.244 1.932 5.716 1.964 ;
  LAYER M2 ;
        RECT 3.244 1.996 5.716 2.028 ;
  LAYER M2 ;
        RECT 3.244 2.06 5.716 2.092 ;
  LAYER M2 ;
        RECT 3.244 2.124 5.716 2.156 ;
  LAYER M2 ;
        RECT 3.244 2.188 5.716 2.22 ;
  LAYER M2 ;
        RECT 3.244 2.252 5.716 2.284 ;
  LAYER M2 ;
        RECT 3.244 2.316 5.716 2.348 ;
  LAYER M2 ;
        RECT 3.244 2.38 5.716 2.412 ;
  LAYER M2 ;
        RECT 3.244 2.444 5.716 2.476 ;
  LAYER M2 ;
        RECT 3.244 2.508 5.716 2.54 ;
  LAYER M2 ;
        RECT 3.244 2.572 5.716 2.604 ;
  LAYER M2 ;
        RECT 3.244 2.636 5.716 2.668 ;
  LAYER M2 ;
        RECT 3.244 2.7 5.716 2.732 ;
  LAYER M2 ;
        RECT 3.244 2.764 5.716 2.796 ;
  LAYER M2 ;
        RECT 3.244 2.828 5.716 2.86 ;
  LAYER M2 ;
        RECT 3.244 2.892 5.716 2.924 ;
  LAYER M2 ;
        RECT 3.244 2.956 5.716 2.988 ;
  LAYER M2 ;
        RECT 3.244 3.02 5.716 3.052 ;
  LAYER M2 ;
        RECT 3.244 3.084 5.716 3.116 ;
  LAYER M2 ;
        RECT 3.244 3.148 5.716 3.18 ;
  LAYER M2 ;
        RECT 3.244 3.212 5.716 3.244 ;
  LAYER M3 ;
        RECT 3.264 0.888 3.296 3.396 ;
  LAYER M3 ;
        RECT 3.328 0.888 3.36 3.396 ;
  LAYER M3 ;
        RECT 3.392 0.888 3.424 3.396 ;
  LAYER M3 ;
        RECT 3.456 0.888 3.488 3.396 ;
  LAYER M3 ;
        RECT 3.52 0.888 3.552 3.396 ;
  LAYER M3 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M3 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M3 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M3 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M3 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M3 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M3 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M3 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M3 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M3 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M3 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M3 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M3 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M3 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M3 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M3 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M3 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M3 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M3 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M3 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M3 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M3 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M3 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M3 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M3 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M3 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M3 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M3 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M3 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M3 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M3 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M3 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M3 ;
        RECT 5.664 0.888 5.696 3.396 ;
  LAYER M1 ;
        RECT 3.279 0.924 3.281 3.36 ;
  LAYER M1 ;
        RECT 3.359 0.924 3.361 3.36 ;
  LAYER M1 ;
        RECT 3.439 0.924 3.441 3.36 ;
  LAYER M1 ;
        RECT 3.519 0.924 3.521 3.36 ;
  LAYER M1 ;
        RECT 3.599 0.924 3.601 3.36 ;
  LAYER M1 ;
        RECT 3.679 0.924 3.681 3.36 ;
  LAYER M1 ;
        RECT 3.759 0.924 3.761 3.36 ;
  LAYER M1 ;
        RECT 3.839 0.924 3.841 3.36 ;
  LAYER M1 ;
        RECT 3.919 0.924 3.921 3.36 ;
  LAYER M1 ;
        RECT 3.999 0.924 4.001 3.36 ;
  LAYER M1 ;
        RECT 4.079 0.924 4.081 3.36 ;
  LAYER M1 ;
        RECT 4.159 0.924 4.161 3.36 ;
  LAYER M1 ;
        RECT 4.239 0.924 4.241 3.36 ;
  LAYER M1 ;
        RECT 4.319 0.924 4.321 3.36 ;
  LAYER M1 ;
        RECT 4.399 0.924 4.401 3.36 ;
  LAYER M1 ;
        RECT 4.479 0.924 4.481 3.36 ;
  LAYER M1 ;
        RECT 4.559 0.924 4.561 3.36 ;
  LAYER M1 ;
        RECT 4.639 0.924 4.641 3.36 ;
  LAYER M1 ;
        RECT 4.719 0.924 4.721 3.36 ;
  LAYER M1 ;
        RECT 4.799 0.924 4.801 3.36 ;
  LAYER M1 ;
        RECT 4.879 0.924 4.881 3.36 ;
  LAYER M1 ;
        RECT 4.959 0.924 4.961 3.36 ;
  LAYER M1 ;
        RECT 5.039 0.924 5.041 3.36 ;
  LAYER M1 ;
        RECT 5.119 0.924 5.121 3.36 ;
  LAYER M1 ;
        RECT 5.199 0.924 5.201 3.36 ;
  LAYER M1 ;
        RECT 5.279 0.924 5.281 3.36 ;
  LAYER M1 ;
        RECT 5.359 0.924 5.361 3.36 ;
  LAYER M1 ;
        RECT 5.439 0.924 5.441 3.36 ;
  LAYER M1 ;
        RECT 5.519 0.924 5.521 3.36 ;
  LAYER M1 ;
        RECT 5.599 0.924 5.601 3.36 ;
  LAYER M2 ;
        RECT 3.28 0.923 5.68 0.925 ;
  LAYER M2 ;
        RECT 3.28 1.007 5.68 1.009 ;
  LAYER M2 ;
        RECT 3.28 1.091 5.68 1.093 ;
  LAYER M2 ;
        RECT 3.28 1.175 5.68 1.177 ;
  LAYER M2 ;
        RECT 3.28 1.259 5.68 1.261 ;
  LAYER M2 ;
        RECT 3.28 1.343 5.68 1.345 ;
  LAYER M2 ;
        RECT 3.28 1.427 5.68 1.429 ;
  LAYER M2 ;
        RECT 3.28 1.511 5.68 1.513 ;
  LAYER M2 ;
        RECT 3.28 1.595 5.68 1.597 ;
  LAYER M2 ;
        RECT 3.28 1.679 5.68 1.681 ;
  LAYER M2 ;
        RECT 3.28 1.763 5.68 1.765 ;
  LAYER M2 ;
        RECT 3.28 1.847 5.68 1.849 ;
  LAYER M2 ;
        RECT 3.28 1.9305 5.68 1.9325 ;
  LAYER M2 ;
        RECT 3.28 2.015 5.68 2.017 ;
  LAYER M2 ;
        RECT 3.28 2.099 5.68 2.101 ;
  LAYER M2 ;
        RECT 3.28 2.183 5.68 2.185 ;
  LAYER M2 ;
        RECT 3.28 2.267 5.68 2.269 ;
  LAYER M2 ;
        RECT 3.28 2.351 5.68 2.353 ;
  LAYER M2 ;
        RECT 3.28 2.435 5.68 2.437 ;
  LAYER M2 ;
        RECT 3.28 2.519 5.68 2.521 ;
  LAYER M2 ;
        RECT 3.28 2.603 5.68 2.605 ;
  LAYER M2 ;
        RECT 3.28 2.687 5.68 2.689 ;
  LAYER M2 ;
        RECT 3.28 2.771 5.68 2.773 ;
  LAYER M2 ;
        RECT 3.28 2.855 5.68 2.857 ;
  LAYER M2 ;
        RECT 3.28 2.939 5.68 2.941 ;
  LAYER M2 ;
        RECT 3.28 3.023 5.68 3.025 ;
  LAYER M2 ;
        RECT 3.28 3.107 5.68 3.109 ;
  LAYER M2 ;
        RECT 3.28 3.191 5.68 3.193 ;
  LAYER M2 ;
        RECT 3.28 3.275 5.68 3.277 ;
  LAYER M1 ;
        RECT 3.264 3.828 3.296 6.336 ;
  LAYER M1 ;
        RECT 3.328 3.828 3.36 6.336 ;
  LAYER M1 ;
        RECT 3.392 3.828 3.424 6.336 ;
  LAYER M1 ;
        RECT 3.456 3.828 3.488 6.336 ;
  LAYER M1 ;
        RECT 3.52 3.828 3.552 6.336 ;
  LAYER M1 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M1 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M1 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M1 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M1 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M1 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M1 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M1 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M1 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M1 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M1 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M1 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M1 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M1 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M1 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M1 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M1 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M1 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M1 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M1 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M1 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M1 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M1 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M1 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M1 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M1 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M1 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M1 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M1 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M1 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M1 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M2 ;
        RECT 3.244 3.912 5.716 3.944 ;
  LAYER M2 ;
        RECT 3.244 3.976 5.716 4.008 ;
  LAYER M2 ;
        RECT 3.244 4.04 5.716 4.072 ;
  LAYER M2 ;
        RECT 3.244 4.104 5.716 4.136 ;
  LAYER M2 ;
        RECT 3.244 4.168 5.716 4.2 ;
  LAYER M2 ;
        RECT 3.244 4.232 5.716 4.264 ;
  LAYER M2 ;
        RECT 3.244 4.296 5.716 4.328 ;
  LAYER M2 ;
        RECT 3.244 4.36 5.716 4.392 ;
  LAYER M2 ;
        RECT 3.244 4.424 5.716 4.456 ;
  LAYER M2 ;
        RECT 3.244 4.488 5.716 4.52 ;
  LAYER M2 ;
        RECT 3.244 4.552 5.716 4.584 ;
  LAYER M2 ;
        RECT 3.244 4.616 5.716 4.648 ;
  LAYER M2 ;
        RECT 3.244 4.68 5.716 4.712 ;
  LAYER M2 ;
        RECT 3.244 4.744 5.716 4.776 ;
  LAYER M2 ;
        RECT 3.244 4.808 5.716 4.84 ;
  LAYER M2 ;
        RECT 3.244 4.872 5.716 4.904 ;
  LAYER M2 ;
        RECT 3.244 4.936 5.716 4.968 ;
  LAYER M2 ;
        RECT 3.244 5 5.716 5.032 ;
  LAYER M2 ;
        RECT 3.244 5.064 5.716 5.096 ;
  LAYER M2 ;
        RECT 3.244 5.128 5.716 5.16 ;
  LAYER M2 ;
        RECT 3.244 5.192 5.716 5.224 ;
  LAYER M2 ;
        RECT 3.244 5.256 5.716 5.288 ;
  LAYER M2 ;
        RECT 3.244 5.32 5.716 5.352 ;
  LAYER M2 ;
        RECT 3.244 5.384 5.716 5.416 ;
  LAYER M2 ;
        RECT 3.244 5.448 5.716 5.48 ;
  LAYER M2 ;
        RECT 3.244 5.512 5.716 5.544 ;
  LAYER M2 ;
        RECT 3.244 5.576 5.716 5.608 ;
  LAYER M2 ;
        RECT 3.244 5.64 5.716 5.672 ;
  LAYER M2 ;
        RECT 3.244 5.704 5.716 5.736 ;
  LAYER M2 ;
        RECT 3.244 5.768 5.716 5.8 ;
  LAYER M2 ;
        RECT 3.244 5.832 5.716 5.864 ;
  LAYER M2 ;
        RECT 3.244 5.896 5.716 5.928 ;
  LAYER M2 ;
        RECT 3.244 5.96 5.716 5.992 ;
  LAYER M2 ;
        RECT 3.244 6.024 5.716 6.056 ;
  LAYER M2 ;
        RECT 3.244 6.088 5.716 6.12 ;
  LAYER M2 ;
        RECT 3.244 6.152 5.716 6.184 ;
  LAYER M3 ;
        RECT 3.264 3.828 3.296 6.336 ;
  LAYER M3 ;
        RECT 3.328 3.828 3.36 6.336 ;
  LAYER M3 ;
        RECT 3.392 3.828 3.424 6.336 ;
  LAYER M3 ;
        RECT 3.456 3.828 3.488 6.336 ;
  LAYER M3 ;
        RECT 3.52 3.828 3.552 6.336 ;
  LAYER M3 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M3 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M3 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M3 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M3 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M3 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M3 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M3 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M3 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M3 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M3 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M3 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M3 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M3 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M3 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M3 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M3 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M3 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M3 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M3 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M3 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M3 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M3 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M3 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M3 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M3 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M3 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M3 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M3 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M3 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M3 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M3 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M3 ;
        RECT 5.664 3.828 5.696 6.336 ;
  LAYER M1 ;
        RECT 3.279 3.864 3.281 6.3 ;
  LAYER M1 ;
        RECT 3.359 3.864 3.361 6.3 ;
  LAYER M1 ;
        RECT 3.439 3.864 3.441 6.3 ;
  LAYER M1 ;
        RECT 3.519 3.864 3.521 6.3 ;
  LAYER M1 ;
        RECT 3.599 3.864 3.601 6.3 ;
  LAYER M1 ;
        RECT 3.679 3.864 3.681 6.3 ;
  LAYER M1 ;
        RECT 3.759 3.864 3.761 6.3 ;
  LAYER M1 ;
        RECT 3.839 3.864 3.841 6.3 ;
  LAYER M1 ;
        RECT 3.919 3.864 3.921 6.3 ;
  LAYER M1 ;
        RECT 3.999 3.864 4.001 6.3 ;
  LAYER M1 ;
        RECT 4.079 3.864 4.081 6.3 ;
  LAYER M1 ;
        RECT 4.159 3.864 4.161 6.3 ;
  LAYER M1 ;
        RECT 4.239 3.864 4.241 6.3 ;
  LAYER M1 ;
        RECT 4.319 3.864 4.321 6.3 ;
  LAYER M1 ;
        RECT 4.399 3.864 4.401 6.3 ;
  LAYER M1 ;
        RECT 4.479 3.864 4.481 6.3 ;
  LAYER M1 ;
        RECT 4.559 3.864 4.561 6.3 ;
  LAYER M1 ;
        RECT 4.639 3.864 4.641 6.3 ;
  LAYER M1 ;
        RECT 4.719 3.864 4.721 6.3 ;
  LAYER M1 ;
        RECT 4.799 3.864 4.801 6.3 ;
  LAYER M1 ;
        RECT 4.879 3.864 4.881 6.3 ;
  LAYER M1 ;
        RECT 4.959 3.864 4.961 6.3 ;
  LAYER M1 ;
        RECT 5.039 3.864 5.041 6.3 ;
  LAYER M1 ;
        RECT 5.119 3.864 5.121 6.3 ;
  LAYER M1 ;
        RECT 5.199 3.864 5.201 6.3 ;
  LAYER M1 ;
        RECT 5.279 3.864 5.281 6.3 ;
  LAYER M1 ;
        RECT 5.359 3.864 5.361 6.3 ;
  LAYER M1 ;
        RECT 5.439 3.864 5.441 6.3 ;
  LAYER M1 ;
        RECT 5.519 3.864 5.521 6.3 ;
  LAYER M1 ;
        RECT 5.599 3.864 5.601 6.3 ;
  LAYER M2 ;
        RECT 3.28 3.863 5.68 3.865 ;
  LAYER M2 ;
        RECT 3.28 3.947 5.68 3.949 ;
  LAYER M2 ;
        RECT 3.28 4.031 5.68 4.033 ;
  LAYER M2 ;
        RECT 3.28 4.115 5.68 4.117 ;
  LAYER M2 ;
        RECT 3.28 4.199 5.68 4.201 ;
  LAYER M2 ;
        RECT 3.28 4.283 5.68 4.285 ;
  LAYER M2 ;
        RECT 3.28 4.367 5.68 4.369 ;
  LAYER M2 ;
        RECT 3.28 4.451 5.68 4.453 ;
  LAYER M2 ;
        RECT 3.28 4.535 5.68 4.537 ;
  LAYER M2 ;
        RECT 3.28 4.619 5.68 4.621 ;
  LAYER M2 ;
        RECT 3.28 4.703 5.68 4.705 ;
  LAYER M2 ;
        RECT 3.28 4.787 5.68 4.789 ;
  LAYER M2 ;
        RECT 3.28 4.8705 5.68 4.8725 ;
  LAYER M2 ;
        RECT 3.28 4.955 5.68 4.957 ;
  LAYER M2 ;
        RECT 3.28 5.039 5.68 5.041 ;
  LAYER M2 ;
        RECT 3.28 5.123 5.68 5.125 ;
  LAYER M2 ;
        RECT 3.28 5.207 5.68 5.209 ;
  LAYER M2 ;
        RECT 3.28 5.291 5.68 5.293 ;
  LAYER M2 ;
        RECT 3.28 5.375 5.68 5.377 ;
  LAYER M2 ;
        RECT 3.28 5.459 5.68 5.461 ;
  LAYER M2 ;
        RECT 3.28 5.543 5.68 5.545 ;
  LAYER M2 ;
        RECT 3.28 5.627 5.68 5.629 ;
  LAYER M2 ;
        RECT 3.28 5.711 5.68 5.713 ;
  LAYER M2 ;
        RECT 3.28 5.795 5.68 5.797 ;
  LAYER M2 ;
        RECT 3.28 5.879 5.68 5.881 ;
  LAYER M2 ;
        RECT 3.28 5.963 5.68 5.965 ;
  LAYER M2 ;
        RECT 3.28 6.047 5.68 6.049 ;
  LAYER M2 ;
        RECT 3.28 6.131 5.68 6.133 ;
  LAYER M2 ;
        RECT 3.28 6.215 5.68 6.217 ;
  LAYER M1 ;
        RECT 3.264 6.768 3.296 9.276 ;
  LAYER M1 ;
        RECT 3.328 6.768 3.36 9.276 ;
  LAYER M1 ;
        RECT 3.392 6.768 3.424 9.276 ;
  LAYER M1 ;
        RECT 3.456 6.768 3.488 9.276 ;
  LAYER M1 ;
        RECT 3.52 6.768 3.552 9.276 ;
  LAYER M1 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M1 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M1 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M1 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M1 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M1 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M1 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M1 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M1 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M1 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M1 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M1 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M1 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M1 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M1 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M1 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M1 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M1 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M1 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M1 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M1 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M1 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M1 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M1 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M1 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M1 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M1 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M1 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M1 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M1 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M1 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M2 ;
        RECT 3.244 6.852 5.716 6.884 ;
  LAYER M2 ;
        RECT 3.244 6.916 5.716 6.948 ;
  LAYER M2 ;
        RECT 3.244 6.98 5.716 7.012 ;
  LAYER M2 ;
        RECT 3.244 7.044 5.716 7.076 ;
  LAYER M2 ;
        RECT 3.244 7.108 5.716 7.14 ;
  LAYER M2 ;
        RECT 3.244 7.172 5.716 7.204 ;
  LAYER M2 ;
        RECT 3.244 7.236 5.716 7.268 ;
  LAYER M2 ;
        RECT 3.244 7.3 5.716 7.332 ;
  LAYER M2 ;
        RECT 3.244 7.364 5.716 7.396 ;
  LAYER M2 ;
        RECT 3.244 7.428 5.716 7.46 ;
  LAYER M2 ;
        RECT 3.244 7.492 5.716 7.524 ;
  LAYER M2 ;
        RECT 3.244 7.556 5.716 7.588 ;
  LAYER M2 ;
        RECT 3.244 7.62 5.716 7.652 ;
  LAYER M2 ;
        RECT 3.244 7.684 5.716 7.716 ;
  LAYER M2 ;
        RECT 3.244 7.748 5.716 7.78 ;
  LAYER M2 ;
        RECT 3.244 7.812 5.716 7.844 ;
  LAYER M2 ;
        RECT 3.244 7.876 5.716 7.908 ;
  LAYER M2 ;
        RECT 3.244 7.94 5.716 7.972 ;
  LAYER M2 ;
        RECT 3.244 8.004 5.716 8.036 ;
  LAYER M2 ;
        RECT 3.244 8.068 5.716 8.1 ;
  LAYER M2 ;
        RECT 3.244 8.132 5.716 8.164 ;
  LAYER M2 ;
        RECT 3.244 8.196 5.716 8.228 ;
  LAYER M2 ;
        RECT 3.244 8.26 5.716 8.292 ;
  LAYER M2 ;
        RECT 3.244 8.324 5.716 8.356 ;
  LAYER M2 ;
        RECT 3.244 8.388 5.716 8.42 ;
  LAYER M2 ;
        RECT 3.244 8.452 5.716 8.484 ;
  LAYER M2 ;
        RECT 3.244 8.516 5.716 8.548 ;
  LAYER M2 ;
        RECT 3.244 8.58 5.716 8.612 ;
  LAYER M2 ;
        RECT 3.244 8.644 5.716 8.676 ;
  LAYER M2 ;
        RECT 3.244 8.708 5.716 8.74 ;
  LAYER M2 ;
        RECT 3.244 8.772 5.716 8.804 ;
  LAYER M2 ;
        RECT 3.244 8.836 5.716 8.868 ;
  LAYER M2 ;
        RECT 3.244 8.9 5.716 8.932 ;
  LAYER M2 ;
        RECT 3.244 8.964 5.716 8.996 ;
  LAYER M2 ;
        RECT 3.244 9.028 5.716 9.06 ;
  LAYER M2 ;
        RECT 3.244 9.092 5.716 9.124 ;
  LAYER M3 ;
        RECT 3.264 6.768 3.296 9.276 ;
  LAYER M3 ;
        RECT 3.328 6.768 3.36 9.276 ;
  LAYER M3 ;
        RECT 3.392 6.768 3.424 9.276 ;
  LAYER M3 ;
        RECT 3.456 6.768 3.488 9.276 ;
  LAYER M3 ;
        RECT 3.52 6.768 3.552 9.276 ;
  LAYER M3 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M3 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M3 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M3 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M3 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M3 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M3 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M3 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M3 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M3 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M3 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M3 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M3 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M3 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M3 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M3 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M3 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M3 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M3 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M3 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M3 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M3 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M3 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M3 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M3 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M3 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M3 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M3 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M3 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M3 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M3 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M3 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M3 ;
        RECT 5.664 6.768 5.696 9.276 ;
  LAYER M1 ;
        RECT 3.279 6.804 3.281 9.24 ;
  LAYER M1 ;
        RECT 3.359 6.804 3.361 9.24 ;
  LAYER M1 ;
        RECT 3.439 6.804 3.441 9.24 ;
  LAYER M1 ;
        RECT 3.519 6.804 3.521 9.24 ;
  LAYER M1 ;
        RECT 3.599 6.804 3.601 9.24 ;
  LAYER M1 ;
        RECT 3.679 6.804 3.681 9.24 ;
  LAYER M1 ;
        RECT 3.759 6.804 3.761 9.24 ;
  LAYER M1 ;
        RECT 3.839 6.804 3.841 9.24 ;
  LAYER M1 ;
        RECT 3.919 6.804 3.921 9.24 ;
  LAYER M1 ;
        RECT 3.999 6.804 4.001 9.24 ;
  LAYER M1 ;
        RECT 4.079 6.804 4.081 9.24 ;
  LAYER M1 ;
        RECT 4.159 6.804 4.161 9.24 ;
  LAYER M1 ;
        RECT 4.239 6.804 4.241 9.24 ;
  LAYER M1 ;
        RECT 4.319 6.804 4.321 9.24 ;
  LAYER M1 ;
        RECT 4.399 6.804 4.401 9.24 ;
  LAYER M1 ;
        RECT 4.479 6.804 4.481 9.24 ;
  LAYER M1 ;
        RECT 4.559 6.804 4.561 9.24 ;
  LAYER M1 ;
        RECT 4.639 6.804 4.641 9.24 ;
  LAYER M1 ;
        RECT 4.719 6.804 4.721 9.24 ;
  LAYER M1 ;
        RECT 4.799 6.804 4.801 9.24 ;
  LAYER M1 ;
        RECT 4.879 6.804 4.881 9.24 ;
  LAYER M1 ;
        RECT 4.959 6.804 4.961 9.24 ;
  LAYER M1 ;
        RECT 5.039 6.804 5.041 9.24 ;
  LAYER M1 ;
        RECT 5.119 6.804 5.121 9.24 ;
  LAYER M1 ;
        RECT 5.199 6.804 5.201 9.24 ;
  LAYER M1 ;
        RECT 5.279 6.804 5.281 9.24 ;
  LAYER M1 ;
        RECT 5.359 6.804 5.361 9.24 ;
  LAYER M1 ;
        RECT 5.439 6.804 5.441 9.24 ;
  LAYER M1 ;
        RECT 5.519 6.804 5.521 9.24 ;
  LAYER M1 ;
        RECT 5.599 6.804 5.601 9.24 ;
  LAYER M2 ;
        RECT 3.28 6.803 5.68 6.805 ;
  LAYER M2 ;
        RECT 3.28 6.887 5.68 6.889 ;
  LAYER M2 ;
        RECT 3.28 6.971 5.68 6.973 ;
  LAYER M2 ;
        RECT 3.28 7.055 5.68 7.057 ;
  LAYER M2 ;
        RECT 3.28 7.139 5.68 7.141 ;
  LAYER M2 ;
        RECT 3.28 7.223 5.68 7.225 ;
  LAYER M2 ;
        RECT 3.28 7.307 5.68 7.309 ;
  LAYER M2 ;
        RECT 3.28 7.391 5.68 7.393 ;
  LAYER M2 ;
        RECT 3.28 7.475 5.68 7.477 ;
  LAYER M2 ;
        RECT 3.28 7.559 5.68 7.561 ;
  LAYER M2 ;
        RECT 3.28 7.643 5.68 7.645 ;
  LAYER M2 ;
        RECT 3.28 7.727 5.68 7.729 ;
  LAYER M2 ;
        RECT 3.28 7.8105 5.68 7.8125 ;
  LAYER M2 ;
        RECT 3.28 7.895 5.68 7.897 ;
  LAYER M2 ;
        RECT 3.28 7.979 5.68 7.981 ;
  LAYER M2 ;
        RECT 3.28 8.063 5.68 8.065 ;
  LAYER M2 ;
        RECT 3.28 8.147 5.68 8.149 ;
  LAYER M2 ;
        RECT 3.28 8.231 5.68 8.233 ;
  LAYER M2 ;
        RECT 3.28 8.315 5.68 8.317 ;
  LAYER M2 ;
        RECT 3.28 8.399 5.68 8.401 ;
  LAYER M2 ;
        RECT 3.28 8.483 5.68 8.485 ;
  LAYER M2 ;
        RECT 3.28 8.567 5.68 8.569 ;
  LAYER M2 ;
        RECT 3.28 8.651 5.68 8.653 ;
  LAYER M2 ;
        RECT 3.28 8.735 5.68 8.737 ;
  LAYER M2 ;
        RECT 3.28 8.819 5.68 8.821 ;
  LAYER M2 ;
        RECT 3.28 8.903 5.68 8.905 ;
  LAYER M2 ;
        RECT 3.28 8.987 5.68 8.989 ;
  LAYER M2 ;
        RECT 3.28 9.071 5.68 9.073 ;
  LAYER M2 ;
        RECT 3.28 9.155 5.68 9.157 ;
  LAYER M1 ;
        RECT 3.264 9.708 3.296 12.216 ;
  LAYER M1 ;
        RECT 3.328 9.708 3.36 12.216 ;
  LAYER M1 ;
        RECT 3.392 9.708 3.424 12.216 ;
  LAYER M1 ;
        RECT 3.456 9.708 3.488 12.216 ;
  LAYER M1 ;
        RECT 3.52 9.708 3.552 12.216 ;
  LAYER M1 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M1 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M1 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M1 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M1 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M1 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M1 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M1 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M1 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M1 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M1 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M1 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M1 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M1 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M1 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M1 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M1 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M1 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M1 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M1 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M1 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M1 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M1 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M1 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M1 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M1 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M1 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M1 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M1 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M1 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M1 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M2 ;
        RECT 3.244 9.792 5.716 9.824 ;
  LAYER M2 ;
        RECT 3.244 9.856 5.716 9.888 ;
  LAYER M2 ;
        RECT 3.244 9.92 5.716 9.952 ;
  LAYER M2 ;
        RECT 3.244 9.984 5.716 10.016 ;
  LAYER M2 ;
        RECT 3.244 10.048 5.716 10.08 ;
  LAYER M2 ;
        RECT 3.244 10.112 5.716 10.144 ;
  LAYER M2 ;
        RECT 3.244 10.176 5.716 10.208 ;
  LAYER M2 ;
        RECT 3.244 10.24 5.716 10.272 ;
  LAYER M2 ;
        RECT 3.244 10.304 5.716 10.336 ;
  LAYER M2 ;
        RECT 3.244 10.368 5.716 10.4 ;
  LAYER M2 ;
        RECT 3.244 10.432 5.716 10.464 ;
  LAYER M2 ;
        RECT 3.244 10.496 5.716 10.528 ;
  LAYER M2 ;
        RECT 3.244 10.56 5.716 10.592 ;
  LAYER M2 ;
        RECT 3.244 10.624 5.716 10.656 ;
  LAYER M2 ;
        RECT 3.244 10.688 5.716 10.72 ;
  LAYER M2 ;
        RECT 3.244 10.752 5.716 10.784 ;
  LAYER M2 ;
        RECT 3.244 10.816 5.716 10.848 ;
  LAYER M2 ;
        RECT 3.244 10.88 5.716 10.912 ;
  LAYER M2 ;
        RECT 3.244 10.944 5.716 10.976 ;
  LAYER M2 ;
        RECT 3.244 11.008 5.716 11.04 ;
  LAYER M2 ;
        RECT 3.244 11.072 5.716 11.104 ;
  LAYER M2 ;
        RECT 3.244 11.136 5.716 11.168 ;
  LAYER M2 ;
        RECT 3.244 11.2 5.716 11.232 ;
  LAYER M2 ;
        RECT 3.244 11.264 5.716 11.296 ;
  LAYER M2 ;
        RECT 3.244 11.328 5.716 11.36 ;
  LAYER M2 ;
        RECT 3.244 11.392 5.716 11.424 ;
  LAYER M2 ;
        RECT 3.244 11.456 5.716 11.488 ;
  LAYER M2 ;
        RECT 3.244 11.52 5.716 11.552 ;
  LAYER M2 ;
        RECT 3.244 11.584 5.716 11.616 ;
  LAYER M2 ;
        RECT 3.244 11.648 5.716 11.68 ;
  LAYER M2 ;
        RECT 3.244 11.712 5.716 11.744 ;
  LAYER M2 ;
        RECT 3.244 11.776 5.716 11.808 ;
  LAYER M2 ;
        RECT 3.244 11.84 5.716 11.872 ;
  LAYER M2 ;
        RECT 3.244 11.904 5.716 11.936 ;
  LAYER M2 ;
        RECT 3.244 11.968 5.716 12 ;
  LAYER M2 ;
        RECT 3.244 12.032 5.716 12.064 ;
  LAYER M3 ;
        RECT 3.264 9.708 3.296 12.216 ;
  LAYER M3 ;
        RECT 3.328 9.708 3.36 12.216 ;
  LAYER M3 ;
        RECT 3.392 9.708 3.424 12.216 ;
  LAYER M3 ;
        RECT 3.456 9.708 3.488 12.216 ;
  LAYER M3 ;
        RECT 3.52 9.708 3.552 12.216 ;
  LAYER M3 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M3 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M3 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M3 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M3 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M3 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M3 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M3 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M3 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M3 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M3 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M3 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M3 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M3 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M3 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M3 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M3 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M3 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M3 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M3 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M3 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M3 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M3 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M3 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M3 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M3 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M3 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M3 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M3 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M3 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M3 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M3 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M3 ;
        RECT 5.664 9.708 5.696 12.216 ;
  LAYER M1 ;
        RECT 3.279 9.744 3.281 12.18 ;
  LAYER M1 ;
        RECT 3.359 9.744 3.361 12.18 ;
  LAYER M1 ;
        RECT 3.439 9.744 3.441 12.18 ;
  LAYER M1 ;
        RECT 3.519 9.744 3.521 12.18 ;
  LAYER M1 ;
        RECT 3.599 9.744 3.601 12.18 ;
  LAYER M1 ;
        RECT 3.679 9.744 3.681 12.18 ;
  LAYER M1 ;
        RECT 3.759 9.744 3.761 12.18 ;
  LAYER M1 ;
        RECT 3.839 9.744 3.841 12.18 ;
  LAYER M1 ;
        RECT 3.919 9.744 3.921 12.18 ;
  LAYER M1 ;
        RECT 3.999 9.744 4.001 12.18 ;
  LAYER M1 ;
        RECT 4.079 9.744 4.081 12.18 ;
  LAYER M1 ;
        RECT 4.159 9.744 4.161 12.18 ;
  LAYER M1 ;
        RECT 4.239 9.744 4.241 12.18 ;
  LAYER M1 ;
        RECT 4.319 9.744 4.321 12.18 ;
  LAYER M1 ;
        RECT 4.399 9.744 4.401 12.18 ;
  LAYER M1 ;
        RECT 4.479 9.744 4.481 12.18 ;
  LAYER M1 ;
        RECT 4.559 9.744 4.561 12.18 ;
  LAYER M1 ;
        RECT 4.639 9.744 4.641 12.18 ;
  LAYER M1 ;
        RECT 4.719 9.744 4.721 12.18 ;
  LAYER M1 ;
        RECT 4.799 9.744 4.801 12.18 ;
  LAYER M1 ;
        RECT 4.879 9.744 4.881 12.18 ;
  LAYER M1 ;
        RECT 4.959 9.744 4.961 12.18 ;
  LAYER M1 ;
        RECT 5.039 9.744 5.041 12.18 ;
  LAYER M1 ;
        RECT 5.119 9.744 5.121 12.18 ;
  LAYER M1 ;
        RECT 5.199 9.744 5.201 12.18 ;
  LAYER M1 ;
        RECT 5.279 9.744 5.281 12.18 ;
  LAYER M1 ;
        RECT 5.359 9.744 5.361 12.18 ;
  LAYER M1 ;
        RECT 5.439 9.744 5.441 12.18 ;
  LAYER M1 ;
        RECT 5.519 9.744 5.521 12.18 ;
  LAYER M1 ;
        RECT 5.599 9.744 5.601 12.18 ;
  LAYER M2 ;
        RECT 3.28 9.743 5.68 9.745 ;
  LAYER M2 ;
        RECT 3.28 9.827 5.68 9.829 ;
  LAYER M2 ;
        RECT 3.28 9.911 5.68 9.913 ;
  LAYER M2 ;
        RECT 3.28 9.995 5.68 9.997 ;
  LAYER M2 ;
        RECT 3.28 10.079 5.68 10.081 ;
  LAYER M2 ;
        RECT 3.28 10.163 5.68 10.165 ;
  LAYER M2 ;
        RECT 3.28 10.247 5.68 10.249 ;
  LAYER M2 ;
        RECT 3.28 10.331 5.68 10.333 ;
  LAYER M2 ;
        RECT 3.28 10.415 5.68 10.417 ;
  LAYER M2 ;
        RECT 3.28 10.499 5.68 10.501 ;
  LAYER M2 ;
        RECT 3.28 10.583 5.68 10.585 ;
  LAYER M2 ;
        RECT 3.28 10.667 5.68 10.669 ;
  LAYER M2 ;
        RECT 3.28 10.7505 5.68 10.7525 ;
  LAYER M2 ;
        RECT 3.28 10.835 5.68 10.837 ;
  LAYER M2 ;
        RECT 3.28 10.919 5.68 10.921 ;
  LAYER M2 ;
        RECT 3.28 11.003 5.68 11.005 ;
  LAYER M2 ;
        RECT 3.28 11.087 5.68 11.089 ;
  LAYER M2 ;
        RECT 3.28 11.171 5.68 11.173 ;
  LAYER M2 ;
        RECT 3.28 11.255 5.68 11.257 ;
  LAYER M2 ;
        RECT 3.28 11.339 5.68 11.341 ;
  LAYER M2 ;
        RECT 3.28 11.423 5.68 11.425 ;
  LAYER M2 ;
        RECT 3.28 11.507 5.68 11.509 ;
  LAYER M2 ;
        RECT 3.28 11.591 5.68 11.593 ;
  LAYER M2 ;
        RECT 3.28 11.675 5.68 11.677 ;
  LAYER M2 ;
        RECT 3.28 11.759 5.68 11.761 ;
  LAYER M2 ;
        RECT 3.28 11.843 5.68 11.845 ;
  LAYER M2 ;
        RECT 3.28 11.927 5.68 11.929 ;
  LAYER M2 ;
        RECT 3.28 12.011 5.68 12.013 ;
  LAYER M2 ;
        RECT 3.28 12.095 5.68 12.097 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 15.156 ;
  LAYER M1 ;
        RECT 3.328 12.648 3.36 15.156 ;
  LAYER M1 ;
        RECT 3.392 12.648 3.424 15.156 ;
  LAYER M1 ;
        RECT 3.456 12.648 3.488 15.156 ;
  LAYER M1 ;
        RECT 3.52 12.648 3.552 15.156 ;
  LAYER M1 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M1 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M1 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M1 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M1 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M1 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M1 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M1 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M1 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M1 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M1 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M1 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M1 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M1 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M1 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M1 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M1 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M1 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M1 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M1 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M1 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M1 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M1 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M1 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M1 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M1 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M1 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M1 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M1 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M1 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M1 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M1 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M2 ;
        RECT 3.244 12.732 5.716 12.764 ;
  LAYER M2 ;
        RECT 3.244 12.796 5.716 12.828 ;
  LAYER M2 ;
        RECT 3.244 12.86 5.716 12.892 ;
  LAYER M2 ;
        RECT 3.244 12.924 5.716 12.956 ;
  LAYER M2 ;
        RECT 3.244 12.988 5.716 13.02 ;
  LAYER M2 ;
        RECT 3.244 13.052 5.716 13.084 ;
  LAYER M2 ;
        RECT 3.244 13.116 5.716 13.148 ;
  LAYER M2 ;
        RECT 3.244 13.18 5.716 13.212 ;
  LAYER M2 ;
        RECT 3.244 13.244 5.716 13.276 ;
  LAYER M2 ;
        RECT 3.244 13.308 5.716 13.34 ;
  LAYER M2 ;
        RECT 3.244 13.372 5.716 13.404 ;
  LAYER M2 ;
        RECT 3.244 13.436 5.716 13.468 ;
  LAYER M2 ;
        RECT 3.244 13.5 5.716 13.532 ;
  LAYER M2 ;
        RECT 3.244 13.564 5.716 13.596 ;
  LAYER M2 ;
        RECT 3.244 13.628 5.716 13.66 ;
  LAYER M2 ;
        RECT 3.244 13.692 5.716 13.724 ;
  LAYER M2 ;
        RECT 3.244 13.756 5.716 13.788 ;
  LAYER M2 ;
        RECT 3.244 13.82 5.716 13.852 ;
  LAYER M2 ;
        RECT 3.244 13.884 5.716 13.916 ;
  LAYER M2 ;
        RECT 3.244 13.948 5.716 13.98 ;
  LAYER M2 ;
        RECT 3.244 14.012 5.716 14.044 ;
  LAYER M2 ;
        RECT 3.244 14.076 5.716 14.108 ;
  LAYER M2 ;
        RECT 3.244 14.14 5.716 14.172 ;
  LAYER M2 ;
        RECT 3.244 14.204 5.716 14.236 ;
  LAYER M2 ;
        RECT 3.244 14.268 5.716 14.3 ;
  LAYER M2 ;
        RECT 3.244 14.332 5.716 14.364 ;
  LAYER M2 ;
        RECT 3.244 14.396 5.716 14.428 ;
  LAYER M2 ;
        RECT 3.244 14.46 5.716 14.492 ;
  LAYER M2 ;
        RECT 3.244 14.524 5.716 14.556 ;
  LAYER M2 ;
        RECT 3.244 14.588 5.716 14.62 ;
  LAYER M2 ;
        RECT 3.244 14.652 5.716 14.684 ;
  LAYER M2 ;
        RECT 3.244 14.716 5.716 14.748 ;
  LAYER M2 ;
        RECT 3.244 14.78 5.716 14.812 ;
  LAYER M2 ;
        RECT 3.244 14.844 5.716 14.876 ;
  LAYER M2 ;
        RECT 3.244 14.908 5.716 14.94 ;
  LAYER M2 ;
        RECT 3.244 14.972 5.716 15.004 ;
  LAYER M3 ;
        RECT 3.264 12.648 3.296 15.156 ;
  LAYER M3 ;
        RECT 3.328 12.648 3.36 15.156 ;
  LAYER M3 ;
        RECT 3.392 12.648 3.424 15.156 ;
  LAYER M3 ;
        RECT 3.456 12.648 3.488 15.156 ;
  LAYER M3 ;
        RECT 3.52 12.648 3.552 15.156 ;
  LAYER M3 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M3 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M3 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M3 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M3 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M3 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M3 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M3 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M3 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M3 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M3 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M3 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M3 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M3 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M3 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M3 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M3 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M3 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M3 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M3 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M3 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M3 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M3 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M3 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M3 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M3 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M3 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M3 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M3 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M3 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M3 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M3 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M3 ;
        RECT 5.664 12.648 5.696 15.156 ;
  LAYER M1 ;
        RECT 3.279 12.684 3.281 15.12 ;
  LAYER M1 ;
        RECT 3.359 12.684 3.361 15.12 ;
  LAYER M1 ;
        RECT 3.439 12.684 3.441 15.12 ;
  LAYER M1 ;
        RECT 3.519 12.684 3.521 15.12 ;
  LAYER M1 ;
        RECT 3.599 12.684 3.601 15.12 ;
  LAYER M1 ;
        RECT 3.679 12.684 3.681 15.12 ;
  LAYER M1 ;
        RECT 3.759 12.684 3.761 15.12 ;
  LAYER M1 ;
        RECT 3.839 12.684 3.841 15.12 ;
  LAYER M1 ;
        RECT 3.919 12.684 3.921 15.12 ;
  LAYER M1 ;
        RECT 3.999 12.684 4.001 15.12 ;
  LAYER M1 ;
        RECT 4.079 12.684 4.081 15.12 ;
  LAYER M1 ;
        RECT 4.159 12.684 4.161 15.12 ;
  LAYER M1 ;
        RECT 4.239 12.684 4.241 15.12 ;
  LAYER M1 ;
        RECT 4.319 12.684 4.321 15.12 ;
  LAYER M1 ;
        RECT 4.399 12.684 4.401 15.12 ;
  LAYER M1 ;
        RECT 4.479 12.684 4.481 15.12 ;
  LAYER M1 ;
        RECT 4.559 12.684 4.561 15.12 ;
  LAYER M1 ;
        RECT 4.639 12.684 4.641 15.12 ;
  LAYER M1 ;
        RECT 4.719 12.684 4.721 15.12 ;
  LAYER M1 ;
        RECT 4.799 12.684 4.801 15.12 ;
  LAYER M1 ;
        RECT 4.879 12.684 4.881 15.12 ;
  LAYER M1 ;
        RECT 4.959 12.684 4.961 15.12 ;
  LAYER M1 ;
        RECT 5.039 12.684 5.041 15.12 ;
  LAYER M1 ;
        RECT 5.119 12.684 5.121 15.12 ;
  LAYER M1 ;
        RECT 5.199 12.684 5.201 15.12 ;
  LAYER M1 ;
        RECT 5.279 12.684 5.281 15.12 ;
  LAYER M1 ;
        RECT 5.359 12.684 5.361 15.12 ;
  LAYER M1 ;
        RECT 5.439 12.684 5.441 15.12 ;
  LAYER M1 ;
        RECT 5.519 12.684 5.521 15.12 ;
  LAYER M1 ;
        RECT 5.599 12.684 5.601 15.12 ;
  LAYER M2 ;
        RECT 3.28 12.683 5.68 12.685 ;
  LAYER M2 ;
        RECT 3.28 12.767 5.68 12.769 ;
  LAYER M2 ;
        RECT 3.28 12.851 5.68 12.853 ;
  LAYER M2 ;
        RECT 3.28 12.935 5.68 12.937 ;
  LAYER M2 ;
        RECT 3.28 13.019 5.68 13.021 ;
  LAYER M2 ;
        RECT 3.28 13.103 5.68 13.105 ;
  LAYER M2 ;
        RECT 3.28 13.187 5.68 13.189 ;
  LAYER M2 ;
        RECT 3.28 13.271 5.68 13.273 ;
  LAYER M2 ;
        RECT 3.28 13.355 5.68 13.357 ;
  LAYER M2 ;
        RECT 3.28 13.439 5.68 13.441 ;
  LAYER M2 ;
        RECT 3.28 13.523 5.68 13.525 ;
  LAYER M2 ;
        RECT 3.28 13.607 5.68 13.609 ;
  LAYER M2 ;
        RECT 3.28 13.6905 5.68 13.6925 ;
  LAYER M2 ;
        RECT 3.28 13.775 5.68 13.777 ;
  LAYER M2 ;
        RECT 3.28 13.859 5.68 13.861 ;
  LAYER M2 ;
        RECT 3.28 13.943 5.68 13.945 ;
  LAYER M2 ;
        RECT 3.28 14.027 5.68 14.029 ;
  LAYER M2 ;
        RECT 3.28 14.111 5.68 14.113 ;
  LAYER M2 ;
        RECT 3.28 14.195 5.68 14.197 ;
  LAYER M2 ;
        RECT 3.28 14.279 5.68 14.281 ;
  LAYER M2 ;
        RECT 3.28 14.363 5.68 14.365 ;
  LAYER M2 ;
        RECT 3.28 14.447 5.68 14.449 ;
  LAYER M2 ;
        RECT 3.28 14.531 5.68 14.533 ;
  LAYER M2 ;
        RECT 3.28 14.615 5.68 14.617 ;
  LAYER M2 ;
        RECT 3.28 14.699 5.68 14.701 ;
  LAYER M2 ;
        RECT 3.28 14.783 5.68 14.785 ;
  LAYER M2 ;
        RECT 3.28 14.867 5.68 14.869 ;
  LAYER M2 ;
        RECT 3.28 14.951 5.68 14.953 ;
  LAYER M2 ;
        RECT 3.28 15.035 5.68 15.037 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 18.096 ;
  LAYER M1 ;
        RECT 3.328 15.588 3.36 18.096 ;
  LAYER M1 ;
        RECT 3.392 15.588 3.424 18.096 ;
  LAYER M1 ;
        RECT 3.456 15.588 3.488 18.096 ;
  LAYER M1 ;
        RECT 3.52 15.588 3.552 18.096 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M1 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M1 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M1 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M1 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M1 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M1 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M1 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M1 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M1 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M1 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M1 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M1 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M1 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M1 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M1 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M1 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M1 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M1 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M1 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M1 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M1 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M1 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M1 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M1 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M1 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M1 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M1 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M1 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M1 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M1 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M2 ;
        RECT 3.244 15.672 5.716 15.704 ;
  LAYER M2 ;
        RECT 3.244 15.736 5.716 15.768 ;
  LAYER M2 ;
        RECT 3.244 15.8 5.716 15.832 ;
  LAYER M2 ;
        RECT 3.244 15.864 5.716 15.896 ;
  LAYER M2 ;
        RECT 3.244 15.928 5.716 15.96 ;
  LAYER M2 ;
        RECT 3.244 15.992 5.716 16.024 ;
  LAYER M2 ;
        RECT 3.244 16.056 5.716 16.088 ;
  LAYER M2 ;
        RECT 3.244 16.12 5.716 16.152 ;
  LAYER M2 ;
        RECT 3.244 16.184 5.716 16.216 ;
  LAYER M2 ;
        RECT 3.244 16.248 5.716 16.28 ;
  LAYER M2 ;
        RECT 3.244 16.312 5.716 16.344 ;
  LAYER M2 ;
        RECT 3.244 16.376 5.716 16.408 ;
  LAYER M2 ;
        RECT 3.244 16.44 5.716 16.472 ;
  LAYER M2 ;
        RECT 3.244 16.504 5.716 16.536 ;
  LAYER M2 ;
        RECT 3.244 16.568 5.716 16.6 ;
  LAYER M2 ;
        RECT 3.244 16.632 5.716 16.664 ;
  LAYER M2 ;
        RECT 3.244 16.696 5.716 16.728 ;
  LAYER M2 ;
        RECT 3.244 16.76 5.716 16.792 ;
  LAYER M2 ;
        RECT 3.244 16.824 5.716 16.856 ;
  LAYER M2 ;
        RECT 3.244 16.888 5.716 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.952 5.716 16.984 ;
  LAYER M2 ;
        RECT 3.244 17.016 5.716 17.048 ;
  LAYER M2 ;
        RECT 3.244 17.08 5.716 17.112 ;
  LAYER M2 ;
        RECT 3.244 17.144 5.716 17.176 ;
  LAYER M2 ;
        RECT 3.244 17.208 5.716 17.24 ;
  LAYER M2 ;
        RECT 3.244 17.272 5.716 17.304 ;
  LAYER M2 ;
        RECT 3.244 17.336 5.716 17.368 ;
  LAYER M2 ;
        RECT 3.244 17.4 5.716 17.432 ;
  LAYER M2 ;
        RECT 3.244 17.464 5.716 17.496 ;
  LAYER M2 ;
        RECT 3.244 17.528 5.716 17.56 ;
  LAYER M2 ;
        RECT 3.244 17.592 5.716 17.624 ;
  LAYER M2 ;
        RECT 3.244 17.656 5.716 17.688 ;
  LAYER M2 ;
        RECT 3.244 17.72 5.716 17.752 ;
  LAYER M2 ;
        RECT 3.244 17.784 5.716 17.816 ;
  LAYER M2 ;
        RECT 3.244 17.848 5.716 17.88 ;
  LAYER M2 ;
        RECT 3.244 17.912 5.716 17.944 ;
  LAYER M3 ;
        RECT 3.264 15.588 3.296 18.096 ;
  LAYER M3 ;
        RECT 3.328 15.588 3.36 18.096 ;
  LAYER M3 ;
        RECT 3.392 15.588 3.424 18.096 ;
  LAYER M3 ;
        RECT 3.456 15.588 3.488 18.096 ;
  LAYER M3 ;
        RECT 3.52 15.588 3.552 18.096 ;
  LAYER M3 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M3 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M3 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M3 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M3 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M3 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M3 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M3 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M3 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M3 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M3 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M3 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M3 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M3 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M3 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M3 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M3 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M3 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M3 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M3 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M3 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M3 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M3 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M3 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M3 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M3 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M3 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M3 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M3 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M3 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M3 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M3 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M3 ;
        RECT 5.664 15.588 5.696 18.096 ;
  LAYER M1 ;
        RECT 3.279 15.624 3.281 18.06 ;
  LAYER M1 ;
        RECT 3.359 15.624 3.361 18.06 ;
  LAYER M1 ;
        RECT 3.439 15.624 3.441 18.06 ;
  LAYER M1 ;
        RECT 3.519 15.624 3.521 18.06 ;
  LAYER M1 ;
        RECT 3.599 15.624 3.601 18.06 ;
  LAYER M1 ;
        RECT 3.679 15.624 3.681 18.06 ;
  LAYER M1 ;
        RECT 3.759 15.624 3.761 18.06 ;
  LAYER M1 ;
        RECT 3.839 15.624 3.841 18.06 ;
  LAYER M1 ;
        RECT 3.919 15.624 3.921 18.06 ;
  LAYER M1 ;
        RECT 3.999 15.624 4.001 18.06 ;
  LAYER M1 ;
        RECT 4.079 15.624 4.081 18.06 ;
  LAYER M1 ;
        RECT 4.159 15.624 4.161 18.06 ;
  LAYER M1 ;
        RECT 4.239 15.624 4.241 18.06 ;
  LAYER M1 ;
        RECT 4.319 15.624 4.321 18.06 ;
  LAYER M1 ;
        RECT 4.399 15.624 4.401 18.06 ;
  LAYER M1 ;
        RECT 4.479 15.624 4.481 18.06 ;
  LAYER M1 ;
        RECT 4.559 15.624 4.561 18.06 ;
  LAYER M1 ;
        RECT 4.639 15.624 4.641 18.06 ;
  LAYER M1 ;
        RECT 4.719 15.624 4.721 18.06 ;
  LAYER M1 ;
        RECT 4.799 15.624 4.801 18.06 ;
  LAYER M1 ;
        RECT 4.879 15.624 4.881 18.06 ;
  LAYER M1 ;
        RECT 4.959 15.624 4.961 18.06 ;
  LAYER M1 ;
        RECT 5.039 15.624 5.041 18.06 ;
  LAYER M1 ;
        RECT 5.119 15.624 5.121 18.06 ;
  LAYER M1 ;
        RECT 5.199 15.624 5.201 18.06 ;
  LAYER M1 ;
        RECT 5.279 15.624 5.281 18.06 ;
  LAYER M1 ;
        RECT 5.359 15.624 5.361 18.06 ;
  LAYER M1 ;
        RECT 5.439 15.624 5.441 18.06 ;
  LAYER M1 ;
        RECT 5.519 15.624 5.521 18.06 ;
  LAYER M1 ;
        RECT 5.599 15.624 5.601 18.06 ;
  LAYER M2 ;
        RECT 3.28 15.623 5.68 15.625 ;
  LAYER M2 ;
        RECT 3.28 15.707 5.68 15.709 ;
  LAYER M2 ;
        RECT 3.28 15.791 5.68 15.793 ;
  LAYER M2 ;
        RECT 3.28 15.875 5.68 15.877 ;
  LAYER M2 ;
        RECT 3.28 15.959 5.68 15.961 ;
  LAYER M2 ;
        RECT 3.28 16.043 5.68 16.045 ;
  LAYER M2 ;
        RECT 3.28 16.127 5.68 16.129 ;
  LAYER M2 ;
        RECT 3.28 16.211 5.68 16.213 ;
  LAYER M2 ;
        RECT 3.28 16.295 5.68 16.297 ;
  LAYER M2 ;
        RECT 3.28 16.379 5.68 16.381 ;
  LAYER M2 ;
        RECT 3.28 16.463 5.68 16.465 ;
  LAYER M2 ;
        RECT 3.28 16.547 5.68 16.549 ;
  LAYER M2 ;
        RECT 3.28 16.6305 5.68 16.6325 ;
  LAYER M2 ;
        RECT 3.28 16.715 5.68 16.717 ;
  LAYER M2 ;
        RECT 3.28 16.799 5.68 16.801 ;
  LAYER M2 ;
        RECT 3.28 16.883 5.68 16.885 ;
  LAYER M2 ;
        RECT 3.28 16.967 5.68 16.969 ;
  LAYER M2 ;
        RECT 3.28 17.051 5.68 17.053 ;
  LAYER M2 ;
        RECT 3.28 17.135 5.68 17.137 ;
  LAYER M2 ;
        RECT 3.28 17.219 5.68 17.221 ;
  LAYER M2 ;
        RECT 3.28 17.303 5.68 17.305 ;
  LAYER M2 ;
        RECT 3.28 17.387 5.68 17.389 ;
  LAYER M2 ;
        RECT 3.28 17.471 5.68 17.473 ;
  LAYER M2 ;
        RECT 3.28 17.555 5.68 17.557 ;
  LAYER M2 ;
        RECT 3.28 17.639 5.68 17.641 ;
  LAYER M2 ;
        RECT 3.28 17.723 5.68 17.725 ;
  LAYER M2 ;
        RECT 3.28 17.807 5.68 17.809 ;
  LAYER M2 ;
        RECT 3.28 17.891 5.68 17.893 ;
  LAYER M2 ;
        RECT 3.28 17.975 5.68 17.977 ;
  LAYER M1 ;
        RECT 3.264 18.528 3.296 21.036 ;
  LAYER M1 ;
        RECT 3.328 18.528 3.36 21.036 ;
  LAYER M1 ;
        RECT 3.392 18.528 3.424 21.036 ;
  LAYER M1 ;
        RECT 3.456 18.528 3.488 21.036 ;
  LAYER M1 ;
        RECT 3.52 18.528 3.552 21.036 ;
  LAYER M1 ;
        RECT 3.584 18.528 3.616 21.036 ;
  LAYER M1 ;
        RECT 3.648 18.528 3.68 21.036 ;
  LAYER M1 ;
        RECT 3.712 18.528 3.744 21.036 ;
  LAYER M1 ;
        RECT 3.776 18.528 3.808 21.036 ;
  LAYER M1 ;
        RECT 3.84 18.528 3.872 21.036 ;
  LAYER M1 ;
        RECT 3.904 18.528 3.936 21.036 ;
  LAYER M1 ;
        RECT 3.968 18.528 4 21.036 ;
  LAYER M1 ;
        RECT 4.032 18.528 4.064 21.036 ;
  LAYER M1 ;
        RECT 4.096 18.528 4.128 21.036 ;
  LAYER M1 ;
        RECT 4.16 18.528 4.192 21.036 ;
  LAYER M1 ;
        RECT 4.224 18.528 4.256 21.036 ;
  LAYER M1 ;
        RECT 4.288 18.528 4.32 21.036 ;
  LAYER M1 ;
        RECT 4.352 18.528 4.384 21.036 ;
  LAYER M1 ;
        RECT 4.416 18.528 4.448 21.036 ;
  LAYER M1 ;
        RECT 4.48 18.528 4.512 21.036 ;
  LAYER M1 ;
        RECT 4.544 18.528 4.576 21.036 ;
  LAYER M1 ;
        RECT 4.608 18.528 4.64 21.036 ;
  LAYER M1 ;
        RECT 4.672 18.528 4.704 21.036 ;
  LAYER M1 ;
        RECT 4.736 18.528 4.768 21.036 ;
  LAYER M1 ;
        RECT 4.8 18.528 4.832 21.036 ;
  LAYER M1 ;
        RECT 4.864 18.528 4.896 21.036 ;
  LAYER M1 ;
        RECT 4.928 18.528 4.96 21.036 ;
  LAYER M1 ;
        RECT 4.992 18.528 5.024 21.036 ;
  LAYER M1 ;
        RECT 5.056 18.528 5.088 21.036 ;
  LAYER M1 ;
        RECT 5.12 18.528 5.152 21.036 ;
  LAYER M1 ;
        RECT 5.184 18.528 5.216 21.036 ;
  LAYER M1 ;
        RECT 5.248 18.528 5.28 21.036 ;
  LAYER M1 ;
        RECT 5.312 18.528 5.344 21.036 ;
  LAYER M1 ;
        RECT 5.376 18.528 5.408 21.036 ;
  LAYER M1 ;
        RECT 5.44 18.528 5.472 21.036 ;
  LAYER M1 ;
        RECT 5.504 18.528 5.536 21.036 ;
  LAYER M1 ;
        RECT 5.568 18.528 5.6 21.036 ;
  LAYER M2 ;
        RECT 3.244 18.612 5.716 18.644 ;
  LAYER M2 ;
        RECT 3.244 18.676 5.716 18.708 ;
  LAYER M2 ;
        RECT 3.244 18.74 5.716 18.772 ;
  LAYER M2 ;
        RECT 3.244 18.804 5.716 18.836 ;
  LAYER M2 ;
        RECT 3.244 18.868 5.716 18.9 ;
  LAYER M2 ;
        RECT 3.244 18.932 5.716 18.964 ;
  LAYER M2 ;
        RECT 3.244 18.996 5.716 19.028 ;
  LAYER M2 ;
        RECT 3.244 19.06 5.716 19.092 ;
  LAYER M2 ;
        RECT 3.244 19.124 5.716 19.156 ;
  LAYER M2 ;
        RECT 3.244 19.188 5.716 19.22 ;
  LAYER M2 ;
        RECT 3.244 19.252 5.716 19.284 ;
  LAYER M2 ;
        RECT 3.244 19.316 5.716 19.348 ;
  LAYER M2 ;
        RECT 3.244 19.38 5.716 19.412 ;
  LAYER M2 ;
        RECT 3.244 19.444 5.716 19.476 ;
  LAYER M2 ;
        RECT 3.244 19.508 5.716 19.54 ;
  LAYER M2 ;
        RECT 3.244 19.572 5.716 19.604 ;
  LAYER M2 ;
        RECT 3.244 19.636 5.716 19.668 ;
  LAYER M2 ;
        RECT 3.244 19.7 5.716 19.732 ;
  LAYER M2 ;
        RECT 3.244 19.764 5.716 19.796 ;
  LAYER M2 ;
        RECT 3.244 19.828 5.716 19.86 ;
  LAYER M2 ;
        RECT 3.244 19.892 5.716 19.924 ;
  LAYER M2 ;
        RECT 3.244 19.956 5.716 19.988 ;
  LAYER M2 ;
        RECT 3.244 20.02 5.716 20.052 ;
  LAYER M2 ;
        RECT 3.244 20.084 5.716 20.116 ;
  LAYER M2 ;
        RECT 3.244 20.148 5.716 20.18 ;
  LAYER M2 ;
        RECT 3.244 20.212 5.716 20.244 ;
  LAYER M2 ;
        RECT 3.244 20.276 5.716 20.308 ;
  LAYER M2 ;
        RECT 3.244 20.34 5.716 20.372 ;
  LAYER M2 ;
        RECT 3.244 20.404 5.716 20.436 ;
  LAYER M2 ;
        RECT 3.244 20.468 5.716 20.5 ;
  LAYER M2 ;
        RECT 3.244 20.532 5.716 20.564 ;
  LAYER M2 ;
        RECT 3.244 20.596 5.716 20.628 ;
  LAYER M2 ;
        RECT 3.244 20.66 5.716 20.692 ;
  LAYER M2 ;
        RECT 3.244 20.724 5.716 20.756 ;
  LAYER M2 ;
        RECT 3.244 20.788 5.716 20.82 ;
  LAYER M2 ;
        RECT 3.244 20.852 5.716 20.884 ;
  LAYER M3 ;
        RECT 3.264 18.528 3.296 21.036 ;
  LAYER M3 ;
        RECT 3.328 18.528 3.36 21.036 ;
  LAYER M3 ;
        RECT 3.392 18.528 3.424 21.036 ;
  LAYER M3 ;
        RECT 3.456 18.528 3.488 21.036 ;
  LAYER M3 ;
        RECT 3.52 18.528 3.552 21.036 ;
  LAYER M3 ;
        RECT 3.584 18.528 3.616 21.036 ;
  LAYER M3 ;
        RECT 3.648 18.528 3.68 21.036 ;
  LAYER M3 ;
        RECT 3.712 18.528 3.744 21.036 ;
  LAYER M3 ;
        RECT 3.776 18.528 3.808 21.036 ;
  LAYER M3 ;
        RECT 3.84 18.528 3.872 21.036 ;
  LAYER M3 ;
        RECT 3.904 18.528 3.936 21.036 ;
  LAYER M3 ;
        RECT 3.968 18.528 4 21.036 ;
  LAYER M3 ;
        RECT 4.032 18.528 4.064 21.036 ;
  LAYER M3 ;
        RECT 4.096 18.528 4.128 21.036 ;
  LAYER M3 ;
        RECT 4.16 18.528 4.192 21.036 ;
  LAYER M3 ;
        RECT 4.224 18.528 4.256 21.036 ;
  LAYER M3 ;
        RECT 4.288 18.528 4.32 21.036 ;
  LAYER M3 ;
        RECT 4.352 18.528 4.384 21.036 ;
  LAYER M3 ;
        RECT 4.416 18.528 4.448 21.036 ;
  LAYER M3 ;
        RECT 4.48 18.528 4.512 21.036 ;
  LAYER M3 ;
        RECT 4.544 18.528 4.576 21.036 ;
  LAYER M3 ;
        RECT 4.608 18.528 4.64 21.036 ;
  LAYER M3 ;
        RECT 4.672 18.528 4.704 21.036 ;
  LAYER M3 ;
        RECT 4.736 18.528 4.768 21.036 ;
  LAYER M3 ;
        RECT 4.8 18.528 4.832 21.036 ;
  LAYER M3 ;
        RECT 4.864 18.528 4.896 21.036 ;
  LAYER M3 ;
        RECT 4.928 18.528 4.96 21.036 ;
  LAYER M3 ;
        RECT 4.992 18.528 5.024 21.036 ;
  LAYER M3 ;
        RECT 5.056 18.528 5.088 21.036 ;
  LAYER M3 ;
        RECT 5.12 18.528 5.152 21.036 ;
  LAYER M3 ;
        RECT 5.184 18.528 5.216 21.036 ;
  LAYER M3 ;
        RECT 5.248 18.528 5.28 21.036 ;
  LAYER M3 ;
        RECT 5.312 18.528 5.344 21.036 ;
  LAYER M3 ;
        RECT 5.376 18.528 5.408 21.036 ;
  LAYER M3 ;
        RECT 5.44 18.528 5.472 21.036 ;
  LAYER M3 ;
        RECT 5.504 18.528 5.536 21.036 ;
  LAYER M3 ;
        RECT 5.568 18.528 5.6 21.036 ;
  LAYER M3 ;
        RECT 5.664 18.528 5.696 21.036 ;
  LAYER M1 ;
        RECT 3.279 18.564 3.281 21 ;
  LAYER M1 ;
        RECT 3.359 18.564 3.361 21 ;
  LAYER M1 ;
        RECT 3.439 18.564 3.441 21 ;
  LAYER M1 ;
        RECT 3.519 18.564 3.521 21 ;
  LAYER M1 ;
        RECT 3.599 18.564 3.601 21 ;
  LAYER M1 ;
        RECT 3.679 18.564 3.681 21 ;
  LAYER M1 ;
        RECT 3.759 18.564 3.761 21 ;
  LAYER M1 ;
        RECT 3.839 18.564 3.841 21 ;
  LAYER M1 ;
        RECT 3.919 18.564 3.921 21 ;
  LAYER M1 ;
        RECT 3.999 18.564 4.001 21 ;
  LAYER M1 ;
        RECT 4.079 18.564 4.081 21 ;
  LAYER M1 ;
        RECT 4.159 18.564 4.161 21 ;
  LAYER M1 ;
        RECT 4.239 18.564 4.241 21 ;
  LAYER M1 ;
        RECT 4.319 18.564 4.321 21 ;
  LAYER M1 ;
        RECT 4.399 18.564 4.401 21 ;
  LAYER M1 ;
        RECT 4.479 18.564 4.481 21 ;
  LAYER M1 ;
        RECT 4.559 18.564 4.561 21 ;
  LAYER M1 ;
        RECT 4.639 18.564 4.641 21 ;
  LAYER M1 ;
        RECT 4.719 18.564 4.721 21 ;
  LAYER M1 ;
        RECT 4.799 18.564 4.801 21 ;
  LAYER M1 ;
        RECT 4.879 18.564 4.881 21 ;
  LAYER M1 ;
        RECT 4.959 18.564 4.961 21 ;
  LAYER M1 ;
        RECT 5.039 18.564 5.041 21 ;
  LAYER M1 ;
        RECT 5.119 18.564 5.121 21 ;
  LAYER M1 ;
        RECT 5.199 18.564 5.201 21 ;
  LAYER M1 ;
        RECT 5.279 18.564 5.281 21 ;
  LAYER M1 ;
        RECT 5.359 18.564 5.361 21 ;
  LAYER M1 ;
        RECT 5.439 18.564 5.441 21 ;
  LAYER M1 ;
        RECT 5.519 18.564 5.521 21 ;
  LAYER M1 ;
        RECT 5.599 18.564 5.601 21 ;
  LAYER M2 ;
        RECT 3.28 18.563 5.68 18.565 ;
  LAYER M2 ;
        RECT 3.28 18.647 5.68 18.649 ;
  LAYER M2 ;
        RECT 3.28 18.731 5.68 18.733 ;
  LAYER M2 ;
        RECT 3.28 18.815 5.68 18.817 ;
  LAYER M2 ;
        RECT 3.28 18.899 5.68 18.901 ;
  LAYER M2 ;
        RECT 3.28 18.983 5.68 18.985 ;
  LAYER M2 ;
        RECT 3.28 19.067 5.68 19.069 ;
  LAYER M2 ;
        RECT 3.28 19.151 5.68 19.153 ;
  LAYER M2 ;
        RECT 3.28 19.235 5.68 19.237 ;
  LAYER M2 ;
        RECT 3.28 19.319 5.68 19.321 ;
  LAYER M2 ;
        RECT 3.28 19.403 5.68 19.405 ;
  LAYER M2 ;
        RECT 3.28 19.487 5.68 19.489 ;
  LAYER M2 ;
        RECT 3.28 19.5705 5.68 19.5725 ;
  LAYER M2 ;
        RECT 3.28 19.655 5.68 19.657 ;
  LAYER M2 ;
        RECT 3.28 19.739 5.68 19.741 ;
  LAYER M2 ;
        RECT 3.28 19.823 5.68 19.825 ;
  LAYER M2 ;
        RECT 3.28 19.907 5.68 19.909 ;
  LAYER M2 ;
        RECT 3.28 19.991 5.68 19.993 ;
  LAYER M2 ;
        RECT 3.28 20.075 5.68 20.077 ;
  LAYER M2 ;
        RECT 3.28 20.159 5.68 20.161 ;
  LAYER M2 ;
        RECT 3.28 20.243 5.68 20.245 ;
  LAYER M2 ;
        RECT 3.28 20.327 5.68 20.329 ;
  LAYER M2 ;
        RECT 3.28 20.411 5.68 20.413 ;
  LAYER M2 ;
        RECT 3.28 20.495 5.68 20.497 ;
  LAYER M2 ;
        RECT 3.28 20.579 5.68 20.581 ;
  LAYER M2 ;
        RECT 3.28 20.663 5.68 20.665 ;
  LAYER M2 ;
        RECT 3.28 20.747 5.68 20.749 ;
  LAYER M2 ;
        RECT 3.28 20.831 5.68 20.833 ;
  LAYER M2 ;
        RECT 3.28 20.915 5.68 20.917 ;
  LAYER M1 ;
        RECT 6.464 0.888 6.496 3.396 ;
  LAYER M1 ;
        RECT 6.528 0.888 6.56 3.396 ;
  LAYER M1 ;
        RECT 6.592 0.888 6.624 3.396 ;
  LAYER M1 ;
        RECT 6.656 0.888 6.688 3.396 ;
  LAYER M1 ;
        RECT 6.72 0.888 6.752 3.396 ;
  LAYER M1 ;
        RECT 6.784 0.888 6.816 3.396 ;
  LAYER M1 ;
        RECT 6.848 0.888 6.88 3.396 ;
  LAYER M1 ;
        RECT 6.912 0.888 6.944 3.396 ;
  LAYER M1 ;
        RECT 6.976 0.888 7.008 3.396 ;
  LAYER M1 ;
        RECT 7.04 0.888 7.072 3.396 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M1 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M1 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M1 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M1 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M1 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M1 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M1 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M1 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M1 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M1 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M1 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M1 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M1 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M1 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M1 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M1 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M1 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M1 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M1 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M1 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M1 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M1 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M1 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M1 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M1 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M1 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M2 ;
        RECT 6.444 0.972 8.916 1.004 ;
  LAYER M2 ;
        RECT 6.444 1.036 8.916 1.068 ;
  LAYER M2 ;
        RECT 6.444 1.1 8.916 1.132 ;
  LAYER M2 ;
        RECT 6.444 1.164 8.916 1.196 ;
  LAYER M2 ;
        RECT 6.444 1.228 8.916 1.26 ;
  LAYER M2 ;
        RECT 6.444 1.292 8.916 1.324 ;
  LAYER M2 ;
        RECT 6.444 1.356 8.916 1.388 ;
  LAYER M2 ;
        RECT 6.444 1.42 8.916 1.452 ;
  LAYER M2 ;
        RECT 6.444 1.484 8.916 1.516 ;
  LAYER M2 ;
        RECT 6.444 1.548 8.916 1.58 ;
  LAYER M2 ;
        RECT 6.444 1.612 8.916 1.644 ;
  LAYER M2 ;
        RECT 6.444 1.676 8.916 1.708 ;
  LAYER M2 ;
        RECT 6.444 1.74 8.916 1.772 ;
  LAYER M2 ;
        RECT 6.444 1.804 8.916 1.836 ;
  LAYER M2 ;
        RECT 6.444 1.868 8.916 1.9 ;
  LAYER M2 ;
        RECT 6.444 1.932 8.916 1.964 ;
  LAYER M2 ;
        RECT 6.444 1.996 8.916 2.028 ;
  LAYER M2 ;
        RECT 6.444 2.06 8.916 2.092 ;
  LAYER M2 ;
        RECT 6.444 2.124 8.916 2.156 ;
  LAYER M2 ;
        RECT 6.444 2.188 8.916 2.22 ;
  LAYER M2 ;
        RECT 6.444 2.252 8.916 2.284 ;
  LAYER M2 ;
        RECT 6.444 2.316 8.916 2.348 ;
  LAYER M2 ;
        RECT 6.444 2.38 8.916 2.412 ;
  LAYER M2 ;
        RECT 6.444 2.444 8.916 2.476 ;
  LAYER M2 ;
        RECT 6.444 2.508 8.916 2.54 ;
  LAYER M2 ;
        RECT 6.444 2.572 8.916 2.604 ;
  LAYER M2 ;
        RECT 6.444 2.636 8.916 2.668 ;
  LAYER M2 ;
        RECT 6.444 2.7 8.916 2.732 ;
  LAYER M2 ;
        RECT 6.444 2.764 8.916 2.796 ;
  LAYER M2 ;
        RECT 6.444 2.828 8.916 2.86 ;
  LAYER M2 ;
        RECT 6.444 2.892 8.916 2.924 ;
  LAYER M2 ;
        RECT 6.444 2.956 8.916 2.988 ;
  LAYER M2 ;
        RECT 6.444 3.02 8.916 3.052 ;
  LAYER M2 ;
        RECT 6.444 3.084 8.916 3.116 ;
  LAYER M2 ;
        RECT 6.444 3.148 8.916 3.18 ;
  LAYER M2 ;
        RECT 6.444 3.212 8.916 3.244 ;
  LAYER M3 ;
        RECT 6.464 0.888 6.496 3.396 ;
  LAYER M3 ;
        RECT 6.528 0.888 6.56 3.396 ;
  LAYER M3 ;
        RECT 6.592 0.888 6.624 3.396 ;
  LAYER M3 ;
        RECT 6.656 0.888 6.688 3.396 ;
  LAYER M3 ;
        RECT 6.72 0.888 6.752 3.396 ;
  LAYER M3 ;
        RECT 6.784 0.888 6.816 3.396 ;
  LAYER M3 ;
        RECT 6.848 0.888 6.88 3.396 ;
  LAYER M3 ;
        RECT 6.912 0.888 6.944 3.396 ;
  LAYER M3 ;
        RECT 6.976 0.888 7.008 3.396 ;
  LAYER M3 ;
        RECT 7.04 0.888 7.072 3.396 ;
  LAYER M3 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M3 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M3 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M3 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M3 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M3 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M3 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M3 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M3 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M3 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M3 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M3 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M3 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M3 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M3 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M3 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M3 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M3 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M3 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M3 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M3 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M3 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M3 ;
        RECT 8.512 0.888 8.544 3.396 ;
  LAYER M3 ;
        RECT 8.576 0.888 8.608 3.396 ;
  LAYER M3 ;
        RECT 8.64 0.888 8.672 3.396 ;
  LAYER M3 ;
        RECT 8.704 0.888 8.736 3.396 ;
  LAYER M3 ;
        RECT 8.768 0.888 8.8 3.396 ;
  LAYER M3 ;
        RECT 8.864 0.888 8.896 3.396 ;
  LAYER M1 ;
        RECT 6.479 0.924 6.481 3.36 ;
  LAYER M1 ;
        RECT 6.559 0.924 6.561 3.36 ;
  LAYER M1 ;
        RECT 6.639 0.924 6.641 3.36 ;
  LAYER M1 ;
        RECT 6.719 0.924 6.721 3.36 ;
  LAYER M1 ;
        RECT 6.799 0.924 6.801 3.36 ;
  LAYER M1 ;
        RECT 6.879 0.924 6.881 3.36 ;
  LAYER M1 ;
        RECT 6.959 0.924 6.961 3.36 ;
  LAYER M1 ;
        RECT 7.039 0.924 7.041 3.36 ;
  LAYER M1 ;
        RECT 7.119 0.924 7.121 3.36 ;
  LAYER M1 ;
        RECT 7.199 0.924 7.201 3.36 ;
  LAYER M1 ;
        RECT 7.279 0.924 7.281 3.36 ;
  LAYER M1 ;
        RECT 7.359 0.924 7.361 3.36 ;
  LAYER M1 ;
        RECT 7.439 0.924 7.441 3.36 ;
  LAYER M1 ;
        RECT 7.519 0.924 7.521 3.36 ;
  LAYER M1 ;
        RECT 7.599 0.924 7.601 3.36 ;
  LAYER M1 ;
        RECT 7.679 0.924 7.681 3.36 ;
  LAYER M1 ;
        RECT 7.759 0.924 7.761 3.36 ;
  LAYER M1 ;
        RECT 7.839 0.924 7.841 3.36 ;
  LAYER M1 ;
        RECT 7.919 0.924 7.921 3.36 ;
  LAYER M1 ;
        RECT 7.999 0.924 8.001 3.36 ;
  LAYER M1 ;
        RECT 8.079 0.924 8.081 3.36 ;
  LAYER M1 ;
        RECT 8.159 0.924 8.161 3.36 ;
  LAYER M1 ;
        RECT 8.239 0.924 8.241 3.36 ;
  LAYER M1 ;
        RECT 8.319 0.924 8.321 3.36 ;
  LAYER M1 ;
        RECT 8.399 0.924 8.401 3.36 ;
  LAYER M1 ;
        RECT 8.479 0.924 8.481 3.36 ;
  LAYER M1 ;
        RECT 8.559 0.924 8.561 3.36 ;
  LAYER M1 ;
        RECT 8.639 0.924 8.641 3.36 ;
  LAYER M1 ;
        RECT 8.719 0.924 8.721 3.36 ;
  LAYER M1 ;
        RECT 8.799 0.924 8.801 3.36 ;
  LAYER M2 ;
        RECT 6.48 0.923 8.88 0.925 ;
  LAYER M2 ;
        RECT 6.48 1.007 8.88 1.009 ;
  LAYER M2 ;
        RECT 6.48 1.091 8.88 1.093 ;
  LAYER M2 ;
        RECT 6.48 1.175 8.88 1.177 ;
  LAYER M2 ;
        RECT 6.48 1.259 8.88 1.261 ;
  LAYER M2 ;
        RECT 6.48 1.343 8.88 1.345 ;
  LAYER M2 ;
        RECT 6.48 1.427 8.88 1.429 ;
  LAYER M2 ;
        RECT 6.48 1.511 8.88 1.513 ;
  LAYER M2 ;
        RECT 6.48 1.595 8.88 1.597 ;
  LAYER M2 ;
        RECT 6.48 1.679 8.88 1.681 ;
  LAYER M2 ;
        RECT 6.48 1.763 8.88 1.765 ;
  LAYER M2 ;
        RECT 6.48 1.847 8.88 1.849 ;
  LAYER M2 ;
        RECT 6.48 1.9305 8.88 1.9325 ;
  LAYER M2 ;
        RECT 6.48 2.015 8.88 2.017 ;
  LAYER M2 ;
        RECT 6.48 2.099 8.88 2.101 ;
  LAYER M2 ;
        RECT 6.48 2.183 8.88 2.185 ;
  LAYER M2 ;
        RECT 6.48 2.267 8.88 2.269 ;
  LAYER M2 ;
        RECT 6.48 2.351 8.88 2.353 ;
  LAYER M2 ;
        RECT 6.48 2.435 8.88 2.437 ;
  LAYER M2 ;
        RECT 6.48 2.519 8.88 2.521 ;
  LAYER M2 ;
        RECT 6.48 2.603 8.88 2.605 ;
  LAYER M2 ;
        RECT 6.48 2.687 8.88 2.689 ;
  LAYER M2 ;
        RECT 6.48 2.771 8.88 2.773 ;
  LAYER M2 ;
        RECT 6.48 2.855 8.88 2.857 ;
  LAYER M2 ;
        RECT 6.48 2.939 8.88 2.941 ;
  LAYER M2 ;
        RECT 6.48 3.023 8.88 3.025 ;
  LAYER M2 ;
        RECT 6.48 3.107 8.88 3.109 ;
  LAYER M2 ;
        RECT 6.48 3.191 8.88 3.193 ;
  LAYER M2 ;
        RECT 6.48 3.275 8.88 3.277 ;
  LAYER M1 ;
        RECT 6.464 3.828 6.496 6.336 ;
  LAYER M1 ;
        RECT 6.528 3.828 6.56 6.336 ;
  LAYER M1 ;
        RECT 6.592 3.828 6.624 6.336 ;
  LAYER M1 ;
        RECT 6.656 3.828 6.688 6.336 ;
  LAYER M1 ;
        RECT 6.72 3.828 6.752 6.336 ;
  LAYER M1 ;
        RECT 6.784 3.828 6.816 6.336 ;
  LAYER M1 ;
        RECT 6.848 3.828 6.88 6.336 ;
  LAYER M1 ;
        RECT 6.912 3.828 6.944 6.336 ;
  LAYER M1 ;
        RECT 6.976 3.828 7.008 6.336 ;
  LAYER M1 ;
        RECT 7.04 3.828 7.072 6.336 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M1 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M1 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M1 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M1 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M1 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M1 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M1 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M1 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M1 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M1 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M1 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M1 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M1 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M1 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M1 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M1 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M1 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M1 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M1 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M1 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M1 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M1 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M1 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M1 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M1 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M1 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M2 ;
        RECT 6.444 3.912 8.916 3.944 ;
  LAYER M2 ;
        RECT 6.444 3.976 8.916 4.008 ;
  LAYER M2 ;
        RECT 6.444 4.04 8.916 4.072 ;
  LAYER M2 ;
        RECT 6.444 4.104 8.916 4.136 ;
  LAYER M2 ;
        RECT 6.444 4.168 8.916 4.2 ;
  LAYER M2 ;
        RECT 6.444 4.232 8.916 4.264 ;
  LAYER M2 ;
        RECT 6.444 4.296 8.916 4.328 ;
  LAYER M2 ;
        RECT 6.444 4.36 8.916 4.392 ;
  LAYER M2 ;
        RECT 6.444 4.424 8.916 4.456 ;
  LAYER M2 ;
        RECT 6.444 4.488 8.916 4.52 ;
  LAYER M2 ;
        RECT 6.444 4.552 8.916 4.584 ;
  LAYER M2 ;
        RECT 6.444 4.616 8.916 4.648 ;
  LAYER M2 ;
        RECT 6.444 4.68 8.916 4.712 ;
  LAYER M2 ;
        RECT 6.444 4.744 8.916 4.776 ;
  LAYER M2 ;
        RECT 6.444 4.808 8.916 4.84 ;
  LAYER M2 ;
        RECT 6.444 4.872 8.916 4.904 ;
  LAYER M2 ;
        RECT 6.444 4.936 8.916 4.968 ;
  LAYER M2 ;
        RECT 6.444 5 8.916 5.032 ;
  LAYER M2 ;
        RECT 6.444 5.064 8.916 5.096 ;
  LAYER M2 ;
        RECT 6.444 5.128 8.916 5.16 ;
  LAYER M2 ;
        RECT 6.444 5.192 8.916 5.224 ;
  LAYER M2 ;
        RECT 6.444 5.256 8.916 5.288 ;
  LAYER M2 ;
        RECT 6.444 5.32 8.916 5.352 ;
  LAYER M2 ;
        RECT 6.444 5.384 8.916 5.416 ;
  LAYER M2 ;
        RECT 6.444 5.448 8.916 5.48 ;
  LAYER M2 ;
        RECT 6.444 5.512 8.916 5.544 ;
  LAYER M2 ;
        RECT 6.444 5.576 8.916 5.608 ;
  LAYER M2 ;
        RECT 6.444 5.64 8.916 5.672 ;
  LAYER M2 ;
        RECT 6.444 5.704 8.916 5.736 ;
  LAYER M2 ;
        RECT 6.444 5.768 8.916 5.8 ;
  LAYER M2 ;
        RECT 6.444 5.832 8.916 5.864 ;
  LAYER M2 ;
        RECT 6.444 5.896 8.916 5.928 ;
  LAYER M2 ;
        RECT 6.444 5.96 8.916 5.992 ;
  LAYER M2 ;
        RECT 6.444 6.024 8.916 6.056 ;
  LAYER M2 ;
        RECT 6.444 6.088 8.916 6.12 ;
  LAYER M2 ;
        RECT 6.444 6.152 8.916 6.184 ;
  LAYER M3 ;
        RECT 6.464 3.828 6.496 6.336 ;
  LAYER M3 ;
        RECT 6.528 3.828 6.56 6.336 ;
  LAYER M3 ;
        RECT 6.592 3.828 6.624 6.336 ;
  LAYER M3 ;
        RECT 6.656 3.828 6.688 6.336 ;
  LAYER M3 ;
        RECT 6.72 3.828 6.752 6.336 ;
  LAYER M3 ;
        RECT 6.784 3.828 6.816 6.336 ;
  LAYER M3 ;
        RECT 6.848 3.828 6.88 6.336 ;
  LAYER M3 ;
        RECT 6.912 3.828 6.944 6.336 ;
  LAYER M3 ;
        RECT 6.976 3.828 7.008 6.336 ;
  LAYER M3 ;
        RECT 7.04 3.828 7.072 6.336 ;
  LAYER M3 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M3 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M3 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M3 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M3 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M3 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M3 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M3 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M3 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M3 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M3 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M3 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M3 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M3 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M3 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M3 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M3 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M3 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M3 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M3 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M3 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M3 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M3 ;
        RECT 8.512 3.828 8.544 6.336 ;
  LAYER M3 ;
        RECT 8.576 3.828 8.608 6.336 ;
  LAYER M3 ;
        RECT 8.64 3.828 8.672 6.336 ;
  LAYER M3 ;
        RECT 8.704 3.828 8.736 6.336 ;
  LAYER M3 ;
        RECT 8.768 3.828 8.8 6.336 ;
  LAYER M3 ;
        RECT 8.864 3.828 8.896 6.336 ;
  LAYER M1 ;
        RECT 6.479 3.864 6.481 6.3 ;
  LAYER M1 ;
        RECT 6.559 3.864 6.561 6.3 ;
  LAYER M1 ;
        RECT 6.639 3.864 6.641 6.3 ;
  LAYER M1 ;
        RECT 6.719 3.864 6.721 6.3 ;
  LAYER M1 ;
        RECT 6.799 3.864 6.801 6.3 ;
  LAYER M1 ;
        RECT 6.879 3.864 6.881 6.3 ;
  LAYER M1 ;
        RECT 6.959 3.864 6.961 6.3 ;
  LAYER M1 ;
        RECT 7.039 3.864 7.041 6.3 ;
  LAYER M1 ;
        RECT 7.119 3.864 7.121 6.3 ;
  LAYER M1 ;
        RECT 7.199 3.864 7.201 6.3 ;
  LAYER M1 ;
        RECT 7.279 3.864 7.281 6.3 ;
  LAYER M1 ;
        RECT 7.359 3.864 7.361 6.3 ;
  LAYER M1 ;
        RECT 7.439 3.864 7.441 6.3 ;
  LAYER M1 ;
        RECT 7.519 3.864 7.521 6.3 ;
  LAYER M1 ;
        RECT 7.599 3.864 7.601 6.3 ;
  LAYER M1 ;
        RECT 7.679 3.864 7.681 6.3 ;
  LAYER M1 ;
        RECT 7.759 3.864 7.761 6.3 ;
  LAYER M1 ;
        RECT 7.839 3.864 7.841 6.3 ;
  LAYER M1 ;
        RECT 7.919 3.864 7.921 6.3 ;
  LAYER M1 ;
        RECT 7.999 3.864 8.001 6.3 ;
  LAYER M1 ;
        RECT 8.079 3.864 8.081 6.3 ;
  LAYER M1 ;
        RECT 8.159 3.864 8.161 6.3 ;
  LAYER M1 ;
        RECT 8.239 3.864 8.241 6.3 ;
  LAYER M1 ;
        RECT 8.319 3.864 8.321 6.3 ;
  LAYER M1 ;
        RECT 8.399 3.864 8.401 6.3 ;
  LAYER M1 ;
        RECT 8.479 3.864 8.481 6.3 ;
  LAYER M1 ;
        RECT 8.559 3.864 8.561 6.3 ;
  LAYER M1 ;
        RECT 8.639 3.864 8.641 6.3 ;
  LAYER M1 ;
        RECT 8.719 3.864 8.721 6.3 ;
  LAYER M1 ;
        RECT 8.799 3.864 8.801 6.3 ;
  LAYER M2 ;
        RECT 6.48 3.863 8.88 3.865 ;
  LAYER M2 ;
        RECT 6.48 3.947 8.88 3.949 ;
  LAYER M2 ;
        RECT 6.48 4.031 8.88 4.033 ;
  LAYER M2 ;
        RECT 6.48 4.115 8.88 4.117 ;
  LAYER M2 ;
        RECT 6.48 4.199 8.88 4.201 ;
  LAYER M2 ;
        RECT 6.48 4.283 8.88 4.285 ;
  LAYER M2 ;
        RECT 6.48 4.367 8.88 4.369 ;
  LAYER M2 ;
        RECT 6.48 4.451 8.88 4.453 ;
  LAYER M2 ;
        RECT 6.48 4.535 8.88 4.537 ;
  LAYER M2 ;
        RECT 6.48 4.619 8.88 4.621 ;
  LAYER M2 ;
        RECT 6.48 4.703 8.88 4.705 ;
  LAYER M2 ;
        RECT 6.48 4.787 8.88 4.789 ;
  LAYER M2 ;
        RECT 6.48 4.8705 8.88 4.8725 ;
  LAYER M2 ;
        RECT 6.48 4.955 8.88 4.957 ;
  LAYER M2 ;
        RECT 6.48 5.039 8.88 5.041 ;
  LAYER M2 ;
        RECT 6.48 5.123 8.88 5.125 ;
  LAYER M2 ;
        RECT 6.48 5.207 8.88 5.209 ;
  LAYER M2 ;
        RECT 6.48 5.291 8.88 5.293 ;
  LAYER M2 ;
        RECT 6.48 5.375 8.88 5.377 ;
  LAYER M2 ;
        RECT 6.48 5.459 8.88 5.461 ;
  LAYER M2 ;
        RECT 6.48 5.543 8.88 5.545 ;
  LAYER M2 ;
        RECT 6.48 5.627 8.88 5.629 ;
  LAYER M2 ;
        RECT 6.48 5.711 8.88 5.713 ;
  LAYER M2 ;
        RECT 6.48 5.795 8.88 5.797 ;
  LAYER M2 ;
        RECT 6.48 5.879 8.88 5.881 ;
  LAYER M2 ;
        RECT 6.48 5.963 8.88 5.965 ;
  LAYER M2 ;
        RECT 6.48 6.047 8.88 6.049 ;
  LAYER M2 ;
        RECT 6.48 6.131 8.88 6.133 ;
  LAYER M2 ;
        RECT 6.48 6.215 8.88 6.217 ;
  LAYER M1 ;
        RECT 6.464 6.768 6.496 9.276 ;
  LAYER M1 ;
        RECT 6.528 6.768 6.56 9.276 ;
  LAYER M1 ;
        RECT 6.592 6.768 6.624 9.276 ;
  LAYER M1 ;
        RECT 6.656 6.768 6.688 9.276 ;
  LAYER M1 ;
        RECT 6.72 6.768 6.752 9.276 ;
  LAYER M1 ;
        RECT 6.784 6.768 6.816 9.276 ;
  LAYER M1 ;
        RECT 6.848 6.768 6.88 9.276 ;
  LAYER M1 ;
        RECT 6.912 6.768 6.944 9.276 ;
  LAYER M1 ;
        RECT 6.976 6.768 7.008 9.276 ;
  LAYER M1 ;
        RECT 7.04 6.768 7.072 9.276 ;
  LAYER M1 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M1 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M1 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M1 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M1 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M1 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M1 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M1 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M1 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M1 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M1 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M1 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M1 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M1 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M1 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M1 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M1 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M1 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M1 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M1 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M1 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M1 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M1 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M1 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M1 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M1 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M1 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M2 ;
        RECT 6.444 6.852 8.916 6.884 ;
  LAYER M2 ;
        RECT 6.444 6.916 8.916 6.948 ;
  LAYER M2 ;
        RECT 6.444 6.98 8.916 7.012 ;
  LAYER M2 ;
        RECT 6.444 7.044 8.916 7.076 ;
  LAYER M2 ;
        RECT 6.444 7.108 8.916 7.14 ;
  LAYER M2 ;
        RECT 6.444 7.172 8.916 7.204 ;
  LAYER M2 ;
        RECT 6.444 7.236 8.916 7.268 ;
  LAYER M2 ;
        RECT 6.444 7.3 8.916 7.332 ;
  LAYER M2 ;
        RECT 6.444 7.364 8.916 7.396 ;
  LAYER M2 ;
        RECT 6.444 7.428 8.916 7.46 ;
  LAYER M2 ;
        RECT 6.444 7.492 8.916 7.524 ;
  LAYER M2 ;
        RECT 6.444 7.556 8.916 7.588 ;
  LAYER M2 ;
        RECT 6.444 7.62 8.916 7.652 ;
  LAYER M2 ;
        RECT 6.444 7.684 8.916 7.716 ;
  LAYER M2 ;
        RECT 6.444 7.748 8.916 7.78 ;
  LAYER M2 ;
        RECT 6.444 7.812 8.916 7.844 ;
  LAYER M2 ;
        RECT 6.444 7.876 8.916 7.908 ;
  LAYER M2 ;
        RECT 6.444 7.94 8.916 7.972 ;
  LAYER M2 ;
        RECT 6.444 8.004 8.916 8.036 ;
  LAYER M2 ;
        RECT 6.444 8.068 8.916 8.1 ;
  LAYER M2 ;
        RECT 6.444 8.132 8.916 8.164 ;
  LAYER M2 ;
        RECT 6.444 8.196 8.916 8.228 ;
  LAYER M2 ;
        RECT 6.444 8.26 8.916 8.292 ;
  LAYER M2 ;
        RECT 6.444 8.324 8.916 8.356 ;
  LAYER M2 ;
        RECT 6.444 8.388 8.916 8.42 ;
  LAYER M2 ;
        RECT 6.444 8.452 8.916 8.484 ;
  LAYER M2 ;
        RECT 6.444 8.516 8.916 8.548 ;
  LAYER M2 ;
        RECT 6.444 8.58 8.916 8.612 ;
  LAYER M2 ;
        RECT 6.444 8.644 8.916 8.676 ;
  LAYER M2 ;
        RECT 6.444 8.708 8.916 8.74 ;
  LAYER M2 ;
        RECT 6.444 8.772 8.916 8.804 ;
  LAYER M2 ;
        RECT 6.444 8.836 8.916 8.868 ;
  LAYER M2 ;
        RECT 6.444 8.9 8.916 8.932 ;
  LAYER M2 ;
        RECT 6.444 8.964 8.916 8.996 ;
  LAYER M2 ;
        RECT 6.444 9.028 8.916 9.06 ;
  LAYER M2 ;
        RECT 6.444 9.092 8.916 9.124 ;
  LAYER M3 ;
        RECT 6.464 6.768 6.496 9.276 ;
  LAYER M3 ;
        RECT 6.528 6.768 6.56 9.276 ;
  LAYER M3 ;
        RECT 6.592 6.768 6.624 9.276 ;
  LAYER M3 ;
        RECT 6.656 6.768 6.688 9.276 ;
  LAYER M3 ;
        RECT 6.72 6.768 6.752 9.276 ;
  LAYER M3 ;
        RECT 6.784 6.768 6.816 9.276 ;
  LAYER M3 ;
        RECT 6.848 6.768 6.88 9.276 ;
  LAYER M3 ;
        RECT 6.912 6.768 6.944 9.276 ;
  LAYER M3 ;
        RECT 6.976 6.768 7.008 9.276 ;
  LAYER M3 ;
        RECT 7.04 6.768 7.072 9.276 ;
  LAYER M3 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M3 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M3 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M3 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M3 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M3 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M3 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M3 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M3 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M3 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M3 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M3 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M3 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M3 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M3 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M3 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M3 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M3 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M3 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M3 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M3 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M3 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M3 ;
        RECT 8.512 6.768 8.544 9.276 ;
  LAYER M3 ;
        RECT 8.576 6.768 8.608 9.276 ;
  LAYER M3 ;
        RECT 8.64 6.768 8.672 9.276 ;
  LAYER M3 ;
        RECT 8.704 6.768 8.736 9.276 ;
  LAYER M3 ;
        RECT 8.768 6.768 8.8 9.276 ;
  LAYER M3 ;
        RECT 8.864 6.768 8.896 9.276 ;
  LAYER M1 ;
        RECT 6.479 6.804 6.481 9.24 ;
  LAYER M1 ;
        RECT 6.559 6.804 6.561 9.24 ;
  LAYER M1 ;
        RECT 6.639 6.804 6.641 9.24 ;
  LAYER M1 ;
        RECT 6.719 6.804 6.721 9.24 ;
  LAYER M1 ;
        RECT 6.799 6.804 6.801 9.24 ;
  LAYER M1 ;
        RECT 6.879 6.804 6.881 9.24 ;
  LAYER M1 ;
        RECT 6.959 6.804 6.961 9.24 ;
  LAYER M1 ;
        RECT 7.039 6.804 7.041 9.24 ;
  LAYER M1 ;
        RECT 7.119 6.804 7.121 9.24 ;
  LAYER M1 ;
        RECT 7.199 6.804 7.201 9.24 ;
  LAYER M1 ;
        RECT 7.279 6.804 7.281 9.24 ;
  LAYER M1 ;
        RECT 7.359 6.804 7.361 9.24 ;
  LAYER M1 ;
        RECT 7.439 6.804 7.441 9.24 ;
  LAYER M1 ;
        RECT 7.519 6.804 7.521 9.24 ;
  LAYER M1 ;
        RECT 7.599 6.804 7.601 9.24 ;
  LAYER M1 ;
        RECT 7.679 6.804 7.681 9.24 ;
  LAYER M1 ;
        RECT 7.759 6.804 7.761 9.24 ;
  LAYER M1 ;
        RECT 7.839 6.804 7.841 9.24 ;
  LAYER M1 ;
        RECT 7.919 6.804 7.921 9.24 ;
  LAYER M1 ;
        RECT 7.999 6.804 8.001 9.24 ;
  LAYER M1 ;
        RECT 8.079 6.804 8.081 9.24 ;
  LAYER M1 ;
        RECT 8.159 6.804 8.161 9.24 ;
  LAYER M1 ;
        RECT 8.239 6.804 8.241 9.24 ;
  LAYER M1 ;
        RECT 8.319 6.804 8.321 9.24 ;
  LAYER M1 ;
        RECT 8.399 6.804 8.401 9.24 ;
  LAYER M1 ;
        RECT 8.479 6.804 8.481 9.24 ;
  LAYER M1 ;
        RECT 8.559 6.804 8.561 9.24 ;
  LAYER M1 ;
        RECT 8.639 6.804 8.641 9.24 ;
  LAYER M1 ;
        RECT 8.719 6.804 8.721 9.24 ;
  LAYER M1 ;
        RECT 8.799 6.804 8.801 9.24 ;
  LAYER M2 ;
        RECT 6.48 6.803 8.88 6.805 ;
  LAYER M2 ;
        RECT 6.48 6.887 8.88 6.889 ;
  LAYER M2 ;
        RECT 6.48 6.971 8.88 6.973 ;
  LAYER M2 ;
        RECT 6.48 7.055 8.88 7.057 ;
  LAYER M2 ;
        RECT 6.48 7.139 8.88 7.141 ;
  LAYER M2 ;
        RECT 6.48 7.223 8.88 7.225 ;
  LAYER M2 ;
        RECT 6.48 7.307 8.88 7.309 ;
  LAYER M2 ;
        RECT 6.48 7.391 8.88 7.393 ;
  LAYER M2 ;
        RECT 6.48 7.475 8.88 7.477 ;
  LAYER M2 ;
        RECT 6.48 7.559 8.88 7.561 ;
  LAYER M2 ;
        RECT 6.48 7.643 8.88 7.645 ;
  LAYER M2 ;
        RECT 6.48 7.727 8.88 7.729 ;
  LAYER M2 ;
        RECT 6.48 7.8105 8.88 7.8125 ;
  LAYER M2 ;
        RECT 6.48 7.895 8.88 7.897 ;
  LAYER M2 ;
        RECT 6.48 7.979 8.88 7.981 ;
  LAYER M2 ;
        RECT 6.48 8.063 8.88 8.065 ;
  LAYER M2 ;
        RECT 6.48 8.147 8.88 8.149 ;
  LAYER M2 ;
        RECT 6.48 8.231 8.88 8.233 ;
  LAYER M2 ;
        RECT 6.48 8.315 8.88 8.317 ;
  LAYER M2 ;
        RECT 6.48 8.399 8.88 8.401 ;
  LAYER M2 ;
        RECT 6.48 8.483 8.88 8.485 ;
  LAYER M2 ;
        RECT 6.48 8.567 8.88 8.569 ;
  LAYER M2 ;
        RECT 6.48 8.651 8.88 8.653 ;
  LAYER M2 ;
        RECT 6.48 8.735 8.88 8.737 ;
  LAYER M2 ;
        RECT 6.48 8.819 8.88 8.821 ;
  LAYER M2 ;
        RECT 6.48 8.903 8.88 8.905 ;
  LAYER M2 ;
        RECT 6.48 8.987 8.88 8.989 ;
  LAYER M2 ;
        RECT 6.48 9.071 8.88 9.073 ;
  LAYER M2 ;
        RECT 6.48 9.155 8.88 9.157 ;
  LAYER M1 ;
        RECT 6.464 9.708 6.496 12.216 ;
  LAYER M1 ;
        RECT 6.528 9.708 6.56 12.216 ;
  LAYER M1 ;
        RECT 6.592 9.708 6.624 12.216 ;
  LAYER M1 ;
        RECT 6.656 9.708 6.688 12.216 ;
  LAYER M1 ;
        RECT 6.72 9.708 6.752 12.216 ;
  LAYER M1 ;
        RECT 6.784 9.708 6.816 12.216 ;
  LAYER M1 ;
        RECT 6.848 9.708 6.88 12.216 ;
  LAYER M1 ;
        RECT 6.912 9.708 6.944 12.216 ;
  LAYER M1 ;
        RECT 6.976 9.708 7.008 12.216 ;
  LAYER M1 ;
        RECT 7.04 9.708 7.072 12.216 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M1 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M1 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M1 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M1 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M1 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M1 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M1 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M1 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M1 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M1 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M1 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M1 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M1 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M1 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M1 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M1 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M1 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M1 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M1 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M1 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M1 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M1 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M1 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M1 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M1 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M1 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M2 ;
        RECT 6.444 9.792 8.916 9.824 ;
  LAYER M2 ;
        RECT 6.444 9.856 8.916 9.888 ;
  LAYER M2 ;
        RECT 6.444 9.92 8.916 9.952 ;
  LAYER M2 ;
        RECT 6.444 9.984 8.916 10.016 ;
  LAYER M2 ;
        RECT 6.444 10.048 8.916 10.08 ;
  LAYER M2 ;
        RECT 6.444 10.112 8.916 10.144 ;
  LAYER M2 ;
        RECT 6.444 10.176 8.916 10.208 ;
  LAYER M2 ;
        RECT 6.444 10.24 8.916 10.272 ;
  LAYER M2 ;
        RECT 6.444 10.304 8.916 10.336 ;
  LAYER M2 ;
        RECT 6.444 10.368 8.916 10.4 ;
  LAYER M2 ;
        RECT 6.444 10.432 8.916 10.464 ;
  LAYER M2 ;
        RECT 6.444 10.496 8.916 10.528 ;
  LAYER M2 ;
        RECT 6.444 10.56 8.916 10.592 ;
  LAYER M2 ;
        RECT 6.444 10.624 8.916 10.656 ;
  LAYER M2 ;
        RECT 6.444 10.688 8.916 10.72 ;
  LAYER M2 ;
        RECT 6.444 10.752 8.916 10.784 ;
  LAYER M2 ;
        RECT 6.444 10.816 8.916 10.848 ;
  LAYER M2 ;
        RECT 6.444 10.88 8.916 10.912 ;
  LAYER M2 ;
        RECT 6.444 10.944 8.916 10.976 ;
  LAYER M2 ;
        RECT 6.444 11.008 8.916 11.04 ;
  LAYER M2 ;
        RECT 6.444 11.072 8.916 11.104 ;
  LAYER M2 ;
        RECT 6.444 11.136 8.916 11.168 ;
  LAYER M2 ;
        RECT 6.444 11.2 8.916 11.232 ;
  LAYER M2 ;
        RECT 6.444 11.264 8.916 11.296 ;
  LAYER M2 ;
        RECT 6.444 11.328 8.916 11.36 ;
  LAYER M2 ;
        RECT 6.444 11.392 8.916 11.424 ;
  LAYER M2 ;
        RECT 6.444 11.456 8.916 11.488 ;
  LAYER M2 ;
        RECT 6.444 11.52 8.916 11.552 ;
  LAYER M2 ;
        RECT 6.444 11.584 8.916 11.616 ;
  LAYER M2 ;
        RECT 6.444 11.648 8.916 11.68 ;
  LAYER M2 ;
        RECT 6.444 11.712 8.916 11.744 ;
  LAYER M2 ;
        RECT 6.444 11.776 8.916 11.808 ;
  LAYER M2 ;
        RECT 6.444 11.84 8.916 11.872 ;
  LAYER M2 ;
        RECT 6.444 11.904 8.916 11.936 ;
  LAYER M2 ;
        RECT 6.444 11.968 8.916 12 ;
  LAYER M2 ;
        RECT 6.444 12.032 8.916 12.064 ;
  LAYER M3 ;
        RECT 6.464 9.708 6.496 12.216 ;
  LAYER M3 ;
        RECT 6.528 9.708 6.56 12.216 ;
  LAYER M3 ;
        RECT 6.592 9.708 6.624 12.216 ;
  LAYER M3 ;
        RECT 6.656 9.708 6.688 12.216 ;
  LAYER M3 ;
        RECT 6.72 9.708 6.752 12.216 ;
  LAYER M3 ;
        RECT 6.784 9.708 6.816 12.216 ;
  LAYER M3 ;
        RECT 6.848 9.708 6.88 12.216 ;
  LAYER M3 ;
        RECT 6.912 9.708 6.944 12.216 ;
  LAYER M3 ;
        RECT 6.976 9.708 7.008 12.216 ;
  LAYER M3 ;
        RECT 7.04 9.708 7.072 12.216 ;
  LAYER M3 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M3 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M3 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M3 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M3 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M3 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M3 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M3 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M3 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M3 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M3 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M3 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M3 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M3 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M3 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M3 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M3 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M3 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M3 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M3 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M3 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M3 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M3 ;
        RECT 8.512 9.708 8.544 12.216 ;
  LAYER M3 ;
        RECT 8.576 9.708 8.608 12.216 ;
  LAYER M3 ;
        RECT 8.64 9.708 8.672 12.216 ;
  LAYER M3 ;
        RECT 8.704 9.708 8.736 12.216 ;
  LAYER M3 ;
        RECT 8.768 9.708 8.8 12.216 ;
  LAYER M3 ;
        RECT 8.864 9.708 8.896 12.216 ;
  LAYER M1 ;
        RECT 6.479 9.744 6.481 12.18 ;
  LAYER M1 ;
        RECT 6.559 9.744 6.561 12.18 ;
  LAYER M1 ;
        RECT 6.639 9.744 6.641 12.18 ;
  LAYER M1 ;
        RECT 6.719 9.744 6.721 12.18 ;
  LAYER M1 ;
        RECT 6.799 9.744 6.801 12.18 ;
  LAYER M1 ;
        RECT 6.879 9.744 6.881 12.18 ;
  LAYER M1 ;
        RECT 6.959 9.744 6.961 12.18 ;
  LAYER M1 ;
        RECT 7.039 9.744 7.041 12.18 ;
  LAYER M1 ;
        RECT 7.119 9.744 7.121 12.18 ;
  LAYER M1 ;
        RECT 7.199 9.744 7.201 12.18 ;
  LAYER M1 ;
        RECT 7.279 9.744 7.281 12.18 ;
  LAYER M1 ;
        RECT 7.359 9.744 7.361 12.18 ;
  LAYER M1 ;
        RECT 7.439 9.744 7.441 12.18 ;
  LAYER M1 ;
        RECT 7.519 9.744 7.521 12.18 ;
  LAYER M1 ;
        RECT 7.599 9.744 7.601 12.18 ;
  LAYER M1 ;
        RECT 7.679 9.744 7.681 12.18 ;
  LAYER M1 ;
        RECT 7.759 9.744 7.761 12.18 ;
  LAYER M1 ;
        RECT 7.839 9.744 7.841 12.18 ;
  LAYER M1 ;
        RECT 7.919 9.744 7.921 12.18 ;
  LAYER M1 ;
        RECT 7.999 9.744 8.001 12.18 ;
  LAYER M1 ;
        RECT 8.079 9.744 8.081 12.18 ;
  LAYER M1 ;
        RECT 8.159 9.744 8.161 12.18 ;
  LAYER M1 ;
        RECT 8.239 9.744 8.241 12.18 ;
  LAYER M1 ;
        RECT 8.319 9.744 8.321 12.18 ;
  LAYER M1 ;
        RECT 8.399 9.744 8.401 12.18 ;
  LAYER M1 ;
        RECT 8.479 9.744 8.481 12.18 ;
  LAYER M1 ;
        RECT 8.559 9.744 8.561 12.18 ;
  LAYER M1 ;
        RECT 8.639 9.744 8.641 12.18 ;
  LAYER M1 ;
        RECT 8.719 9.744 8.721 12.18 ;
  LAYER M1 ;
        RECT 8.799 9.744 8.801 12.18 ;
  LAYER M2 ;
        RECT 6.48 9.743 8.88 9.745 ;
  LAYER M2 ;
        RECT 6.48 9.827 8.88 9.829 ;
  LAYER M2 ;
        RECT 6.48 9.911 8.88 9.913 ;
  LAYER M2 ;
        RECT 6.48 9.995 8.88 9.997 ;
  LAYER M2 ;
        RECT 6.48 10.079 8.88 10.081 ;
  LAYER M2 ;
        RECT 6.48 10.163 8.88 10.165 ;
  LAYER M2 ;
        RECT 6.48 10.247 8.88 10.249 ;
  LAYER M2 ;
        RECT 6.48 10.331 8.88 10.333 ;
  LAYER M2 ;
        RECT 6.48 10.415 8.88 10.417 ;
  LAYER M2 ;
        RECT 6.48 10.499 8.88 10.501 ;
  LAYER M2 ;
        RECT 6.48 10.583 8.88 10.585 ;
  LAYER M2 ;
        RECT 6.48 10.667 8.88 10.669 ;
  LAYER M2 ;
        RECT 6.48 10.7505 8.88 10.7525 ;
  LAYER M2 ;
        RECT 6.48 10.835 8.88 10.837 ;
  LAYER M2 ;
        RECT 6.48 10.919 8.88 10.921 ;
  LAYER M2 ;
        RECT 6.48 11.003 8.88 11.005 ;
  LAYER M2 ;
        RECT 6.48 11.087 8.88 11.089 ;
  LAYER M2 ;
        RECT 6.48 11.171 8.88 11.173 ;
  LAYER M2 ;
        RECT 6.48 11.255 8.88 11.257 ;
  LAYER M2 ;
        RECT 6.48 11.339 8.88 11.341 ;
  LAYER M2 ;
        RECT 6.48 11.423 8.88 11.425 ;
  LAYER M2 ;
        RECT 6.48 11.507 8.88 11.509 ;
  LAYER M2 ;
        RECT 6.48 11.591 8.88 11.593 ;
  LAYER M2 ;
        RECT 6.48 11.675 8.88 11.677 ;
  LAYER M2 ;
        RECT 6.48 11.759 8.88 11.761 ;
  LAYER M2 ;
        RECT 6.48 11.843 8.88 11.845 ;
  LAYER M2 ;
        RECT 6.48 11.927 8.88 11.929 ;
  LAYER M2 ;
        RECT 6.48 12.011 8.88 12.013 ;
  LAYER M2 ;
        RECT 6.48 12.095 8.88 12.097 ;
  LAYER M1 ;
        RECT 6.464 12.648 6.496 15.156 ;
  LAYER M1 ;
        RECT 6.528 12.648 6.56 15.156 ;
  LAYER M1 ;
        RECT 6.592 12.648 6.624 15.156 ;
  LAYER M1 ;
        RECT 6.656 12.648 6.688 15.156 ;
  LAYER M1 ;
        RECT 6.72 12.648 6.752 15.156 ;
  LAYER M1 ;
        RECT 6.784 12.648 6.816 15.156 ;
  LAYER M1 ;
        RECT 6.848 12.648 6.88 15.156 ;
  LAYER M1 ;
        RECT 6.912 12.648 6.944 15.156 ;
  LAYER M1 ;
        RECT 6.976 12.648 7.008 15.156 ;
  LAYER M1 ;
        RECT 7.04 12.648 7.072 15.156 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M1 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M1 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M1 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M1 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M1 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M1 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M1 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M1 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M1 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M1 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M1 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M1 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M1 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M1 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M1 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M1 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M1 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M1 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M1 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M1 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M1 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M1 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M1 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M1 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M1 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M1 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M2 ;
        RECT 6.444 12.732 8.916 12.764 ;
  LAYER M2 ;
        RECT 6.444 12.796 8.916 12.828 ;
  LAYER M2 ;
        RECT 6.444 12.86 8.916 12.892 ;
  LAYER M2 ;
        RECT 6.444 12.924 8.916 12.956 ;
  LAYER M2 ;
        RECT 6.444 12.988 8.916 13.02 ;
  LAYER M2 ;
        RECT 6.444 13.052 8.916 13.084 ;
  LAYER M2 ;
        RECT 6.444 13.116 8.916 13.148 ;
  LAYER M2 ;
        RECT 6.444 13.18 8.916 13.212 ;
  LAYER M2 ;
        RECT 6.444 13.244 8.916 13.276 ;
  LAYER M2 ;
        RECT 6.444 13.308 8.916 13.34 ;
  LAYER M2 ;
        RECT 6.444 13.372 8.916 13.404 ;
  LAYER M2 ;
        RECT 6.444 13.436 8.916 13.468 ;
  LAYER M2 ;
        RECT 6.444 13.5 8.916 13.532 ;
  LAYER M2 ;
        RECT 6.444 13.564 8.916 13.596 ;
  LAYER M2 ;
        RECT 6.444 13.628 8.916 13.66 ;
  LAYER M2 ;
        RECT 6.444 13.692 8.916 13.724 ;
  LAYER M2 ;
        RECT 6.444 13.756 8.916 13.788 ;
  LAYER M2 ;
        RECT 6.444 13.82 8.916 13.852 ;
  LAYER M2 ;
        RECT 6.444 13.884 8.916 13.916 ;
  LAYER M2 ;
        RECT 6.444 13.948 8.916 13.98 ;
  LAYER M2 ;
        RECT 6.444 14.012 8.916 14.044 ;
  LAYER M2 ;
        RECT 6.444 14.076 8.916 14.108 ;
  LAYER M2 ;
        RECT 6.444 14.14 8.916 14.172 ;
  LAYER M2 ;
        RECT 6.444 14.204 8.916 14.236 ;
  LAYER M2 ;
        RECT 6.444 14.268 8.916 14.3 ;
  LAYER M2 ;
        RECT 6.444 14.332 8.916 14.364 ;
  LAYER M2 ;
        RECT 6.444 14.396 8.916 14.428 ;
  LAYER M2 ;
        RECT 6.444 14.46 8.916 14.492 ;
  LAYER M2 ;
        RECT 6.444 14.524 8.916 14.556 ;
  LAYER M2 ;
        RECT 6.444 14.588 8.916 14.62 ;
  LAYER M2 ;
        RECT 6.444 14.652 8.916 14.684 ;
  LAYER M2 ;
        RECT 6.444 14.716 8.916 14.748 ;
  LAYER M2 ;
        RECT 6.444 14.78 8.916 14.812 ;
  LAYER M2 ;
        RECT 6.444 14.844 8.916 14.876 ;
  LAYER M2 ;
        RECT 6.444 14.908 8.916 14.94 ;
  LAYER M2 ;
        RECT 6.444 14.972 8.916 15.004 ;
  LAYER M3 ;
        RECT 6.464 12.648 6.496 15.156 ;
  LAYER M3 ;
        RECT 6.528 12.648 6.56 15.156 ;
  LAYER M3 ;
        RECT 6.592 12.648 6.624 15.156 ;
  LAYER M3 ;
        RECT 6.656 12.648 6.688 15.156 ;
  LAYER M3 ;
        RECT 6.72 12.648 6.752 15.156 ;
  LAYER M3 ;
        RECT 6.784 12.648 6.816 15.156 ;
  LAYER M3 ;
        RECT 6.848 12.648 6.88 15.156 ;
  LAYER M3 ;
        RECT 6.912 12.648 6.944 15.156 ;
  LAYER M3 ;
        RECT 6.976 12.648 7.008 15.156 ;
  LAYER M3 ;
        RECT 7.04 12.648 7.072 15.156 ;
  LAYER M3 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M3 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M3 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M3 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M3 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M3 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M3 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M3 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M3 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M3 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M3 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M3 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M3 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M3 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M3 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M3 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M3 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M3 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M3 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M3 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M3 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M3 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M3 ;
        RECT 8.512 12.648 8.544 15.156 ;
  LAYER M3 ;
        RECT 8.576 12.648 8.608 15.156 ;
  LAYER M3 ;
        RECT 8.64 12.648 8.672 15.156 ;
  LAYER M3 ;
        RECT 8.704 12.648 8.736 15.156 ;
  LAYER M3 ;
        RECT 8.768 12.648 8.8 15.156 ;
  LAYER M3 ;
        RECT 8.864 12.648 8.896 15.156 ;
  LAYER M1 ;
        RECT 6.479 12.684 6.481 15.12 ;
  LAYER M1 ;
        RECT 6.559 12.684 6.561 15.12 ;
  LAYER M1 ;
        RECT 6.639 12.684 6.641 15.12 ;
  LAYER M1 ;
        RECT 6.719 12.684 6.721 15.12 ;
  LAYER M1 ;
        RECT 6.799 12.684 6.801 15.12 ;
  LAYER M1 ;
        RECT 6.879 12.684 6.881 15.12 ;
  LAYER M1 ;
        RECT 6.959 12.684 6.961 15.12 ;
  LAYER M1 ;
        RECT 7.039 12.684 7.041 15.12 ;
  LAYER M1 ;
        RECT 7.119 12.684 7.121 15.12 ;
  LAYER M1 ;
        RECT 7.199 12.684 7.201 15.12 ;
  LAYER M1 ;
        RECT 7.279 12.684 7.281 15.12 ;
  LAYER M1 ;
        RECT 7.359 12.684 7.361 15.12 ;
  LAYER M1 ;
        RECT 7.439 12.684 7.441 15.12 ;
  LAYER M1 ;
        RECT 7.519 12.684 7.521 15.12 ;
  LAYER M1 ;
        RECT 7.599 12.684 7.601 15.12 ;
  LAYER M1 ;
        RECT 7.679 12.684 7.681 15.12 ;
  LAYER M1 ;
        RECT 7.759 12.684 7.761 15.12 ;
  LAYER M1 ;
        RECT 7.839 12.684 7.841 15.12 ;
  LAYER M1 ;
        RECT 7.919 12.684 7.921 15.12 ;
  LAYER M1 ;
        RECT 7.999 12.684 8.001 15.12 ;
  LAYER M1 ;
        RECT 8.079 12.684 8.081 15.12 ;
  LAYER M1 ;
        RECT 8.159 12.684 8.161 15.12 ;
  LAYER M1 ;
        RECT 8.239 12.684 8.241 15.12 ;
  LAYER M1 ;
        RECT 8.319 12.684 8.321 15.12 ;
  LAYER M1 ;
        RECT 8.399 12.684 8.401 15.12 ;
  LAYER M1 ;
        RECT 8.479 12.684 8.481 15.12 ;
  LAYER M1 ;
        RECT 8.559 12.684 8.561 15.12 ;
  LAYER M1 ;
        RECT 8.639 12.684 8.641 15.12 ;
  LAYER M1 ;
        RECT 8.719 12.684 8.721 15.12 ;
  LAYER M1 ;
        RECT 8.799 12.684 8.801 15.12 ;
  LAYER M2 ;
        RECT 6.48 12.683 8.88 12.685 ;
  LAYER M2 ;
        RECT 6.48 12.767 8.88 12.769 ;
  LAYER M2 ;
        RECT 6.48 12.851 8.88 12.853 ;
  LAYER M2 ;
        RECT 6.48 12.935 8.88 12.937 ;
  LAYER M2 ;
        RECT 6.48 13.019 8.88 13.021 ;
  LAYER M2 ;
        RECT 6.48 13.103 8.88 13.105 ;
  LAYER M2 ;
        RECT 6.48 13.187 8.88 13.189 ;
  LAYER M2 ;
        RECT 6.48 13.271 8.88 13.273 ;
  LAYER M2 ;
        RECT 6.48 13.355 8.88 13.357 ;
  LAYER M2 ;
        RECT 6.48 13.439 8.88 13.441 ;
  LAYER M2 ;
        RECT 6.48 13.523 8.88 13.525 ;
  LAYER M2 ;
        RECT 6.48 13.607 8.88 13.609 ;
  LAYER M2 ;
        RECT 6.48 13.6905 8.88 13.6925 ;
  LAYER M2 ;
        RECT 6.48 13.775 8.88 13.777 ;
  LAYER M2 ;
        RECT 6.48 13.859 8.88 13.861 ;
  LAYER M2 ;
        RECT 6.48 13.943 8.88 13.945 ;
  LAYER M2 ;
        RECT 6.48 14.027 8.88 14.029 ;
  LAYER M2 ;
        RECT 6.48 14.111 8.88 14.113 ;
  LAYER M2 ;
        RECT 6.48 14.195 8.88 14.197 ;
  LAYER M2 ;
        RECT 6.48 14.279 8.88 14.281 ;
  LAYER M2 ;
        RECT 6.48 14.363 8.88 14.365 ;
  LAYER M2 ;
        RECT 6.48 14.447 8.88 14.449 ;
  LAYER M2 ;
        RECT 6.48 14.531 8.88 14.533 ;
  LAYER M2 ;
        RECT 6.48 14.615 8.88 14.617 ;
  LAYER M2 ;
        RECT 6.48 14.699 8.88 14.701 ;
  LAYER M2 ;
        RECT 6.48 14.783 8.88 14.785 ;
  LAYER M2 ;
        RECT 6.48 14.867 8.88 14.869 ;
  LAYER M2 ;
        RECT 6.48 14.951 8.88 14.953 ;
  LAYER M2 ;
        RECT 6.48 15.035 8.88 15.037 ;
  LAYER M1 ;
        RECT 6.464 15.588 6.496 18.096 ;
  LAYER M1 ;
        RECT 6.528 15.588 6.56 18.096 ;
  LAYER M1 ;
        RECT 6.592 15.588 6.624 18.096 ;
  LAYER M1 ;
        RECT 6.656 15.588 6.688 18.096 ;
  LAYER M1 ;
        RECT 6.72 15.588 6.752 18.096 ;
  LAYER M1 ;
        RECT 6.784 15.588 6.816 18.096 ;
  LAYER M1 ;
        RECT 6.848 15.588 6.88 18.096 ;
  LAYER M1 ;
        RECT 6.912 15.588 6.944 18.096 ;
  LAYER M1 ;
        RECT 6.976 15.588 7.008 18.096 ;
  LAYER M1 ;
        RECT 7.04 15.588 7.072 18.096 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M1 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M1 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M1 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M1 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M1 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M1 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M1 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M1 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M1 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M1 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M1 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M1 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M1 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M1 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M1 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M1 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M1 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M1 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M1 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M1 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M1 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M1 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M1 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M1 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M1 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M1 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M2 ;
        RECT 6.444 15.672 8.916 15.704 ;
  LAYER M2 ;
        RECT 6.444 15.736 8.916 15.768 ;
  LAYER M2 ;
        RECT 6.444 15.8 8.916 15.832 ;
  LAYER M2 ;
        RECT 6.444 15.864 8.916 15.896 ;
  LAYER M2 ;
        RECT 6.444 15.928 8.916 15.96 ;
  LAYER M2 ;
        RECT 6.444 15.992 8.916 16.024 ;
  LAYER M2 ;
        RECT 6.444 16.056 8.916 16.088 ;
  LAYER M2 ;
        RECT 6.444 16.12 8.916 16.152 ;
  LAYER M2 ;
        RECT 6.444 16.184 8.916 16.216 ;
  LAYER M2 ;
        RECT 6.444 16.248 8.916 16.28 ;
  LAYER M2 ;
        RECT 6.444 16.312 8.916 16.344 ;
  LAYER M2 ;
        RECT 6.444 16.376 8.916 16.408 ;
  LAYER M2 ;
        RECT 6.444 16.44 8.916 16.472 ;
  LAYER M2 ;
        RECT 6.444 16.504 8.916 16.536 ;
  LAYER M2 ;
        RECT 6.444 16.568 8.916 16.6 ;
  LAYER M2 ;
        RECT 6.444 16.632 8.916 16.664 ;
  LAYER M2 ;
        RECT 6.444 16.696 8.916 16.728 ;
  LAYER M2 ;
        RECT 6.444 16.76 8.916 16.792 ;
  LAYER M2 ;
        RECT 6.444 16.824 8.916 16.856 ;
  LAYER M2 ;
        RECT 6.444 16.888 8.916 16.92 ;
  LAYER M2 ;
        RECT 6.444 16.952 8.916 16.984 ;
  LAYER M2 ;
        RECT 6.444 17.016 8.916 17.048 ;
  LAYER M2 ;
        RECT 6.444 17.08 8.916 17.112 ;
  LAYER M2 ;
        RECT 6.444 17.144 8.916 17.176 ;
  LAYER M2 ;
        RECT 6.444 17.208 8.916 17.24 ;
  LAYER M2 ;
        RECT 6.444 17.272 8.916 17.304 ;
  LAYER M2 ;
        RECT 6.444 17.336 8.916 17.368 ;
  LAYER M2 ;
        RECT 6.444 17.4 8.916 17.432 ;
  LAYER M2 ;
        RECT 6.444 17.464 8.916 17.496 ;
  LAYER M2 ;
        RECT 6.444 17.528 8.916 17.56 ;
  LAYER M2 ;
        RECT 6.444 17.592 8.916 17.624 ;
  LAYER M2 ;
        RECT 6.444 17.656 8.916 17.688 ;
  LAYER M2 ;
        RECT 6.444 17.72 8.916 17.752 ;
  LAYER M2 ;
        RECT 6.444 17.784 8.916 17.816 ;
  LAYER M2 ;
        RECT 6.444 17.848 8.916 17.88 ;
  LAYER M2 ;
        RECT 6.444 17.912 8.916 17.944 ;
  LAYER M3 ;
        RECT 6.464 15.588 6.496 18.096 ;
  LAYER M3 ;
        RECT 6.528 15.588 6.56 18.096 ;
  LAYER M3 ;
        RECT 6.592 15.588 6.624 18.096 ;
  LAYER M3 ;
        RECT 6.656 15.588 6.688 18.096 ;
  LAYER M3 ;
        RECT 6.72 15.588 6.752 18.096 ;
  LAYER M3 ;
        RECT 6.784 15.588 6.816 18.096 ;
  LAYER M3 ;
        RECT 6.848 15.588 6.88 18.096 ;
  LAYER M3 ;
        RECT 6.912 15.588 6.944 18.096 ;
  LAYER M3 ;
        RECT 6.976 15.588 7.008 18.096 ;
  LAYER M3 ;
        RECT 7.04 15.588 7.072 18.096 ;
  LAYER M3 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M3 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M3 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M3 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M3 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M3 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M3 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M3 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M3 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M3 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M3 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M3 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M3 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M3 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M3 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M3 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M3 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M3 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M3 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M3 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M3 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M3 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M3 ;
        RECT 8.512 15.588 8.544 18.096 ;
  LAYER M3 ;
        RECT 8.576 15.588 8.608 18.096 ;
  LAYER M3 ;
        RECT 8.64 15.588 8.672 18.096 ;
  LAYER M3 ;
        RECT 8.704 15.588 8.736 18.096 ;
  LAYER M3 ;
        RECT 8.768 15.588 8.8 18.096 ;
  LAYER M3 ;
        RECT 8.864 15.588 8.896 18.096 ;
  LAYER M1 ;
        RECT 6.479 15.624 6.481 18.06 ;
  LAYER M1 ;
        RECT 6.559 15.624 6.561 18.06 ;
  LAYER M1 ;
        RECT 6.639 15.624 6.641 18.06 ;
  LAYER M1 ;
        RECT 6.719 15.624 6.721 18.06 ;
  LAYER M1 ;
        RECT 6.799 15.624 6.801 18.06 ;
  LAYER M1 ;
        RECT 6.879 15.624 6.881 18.06 ;
  LAYER M1 ;
        RECT 6.959 15.624 6.961 18.06 ;
  LAYER M1 ;
        RECT 7.039 15.624 7.041 18.06 ;
  LAYER M1 ;
        RECT 7.119 15.624 7.121 18.06 ;
  LAYER M1 ;
        RECT 7.199 15.624 7.201 18.06 ;
  LAYER M1 ;
        RECT 7.279 15.624 7.281 18.06 ;
  LAYER M1 ;
        RECT 7.359 15.624 7.361 18.06 ;
  LAYER M1 ;
        RECT 7.439 15.624 7.441 18.06 ;
  LAYER M1 ;
        RECT 7.519 15.624 7.521 18.06 ;
  LAYER M1 ;
        RECT 7.599 15.624 7.601 18.06 ;
  LAYER M1 ;
        RECT 7.679 15.624 7.681 18.06 ;
  LAYER M1 ;
        RECT 7.759 15.624 7.761 18.06 ;
  LAYER M1 ;
        RECT 7.839 15.624 7.841 18.06 ;
  LAYER M1 ;
        RECT 7.919 15.624 7.921 18.06 ;
  LAYER M1 ;
        RECT 7.999 15.624 8.001 18.06 ;
  LAYER M1 ;
        RECT 8.079 15.624 8.081 18.06 ;
  LAYER M1 ;
        RECT 8.159 15.624 8.161 18.06 ;
  LAYER M1 ;
        RECT 8.239 15.624 8.241 18.06 ;
  LAYER M1 ;
        RECT 8.319 15.624 8.321 18.06 ;
  LAYER M1 ;
        RECT 8.399 15.624 8.401 18.06 ;
  LAYER M1 ;
        RECT 8.479 15.624 8.481 18.06 ;
  LAYER M1 ;
        RECT 8.559 15.624 8.561 18.06 ;
  LAYER M1 ;
        RECT 8.639 15.624 8.641 18.06 ;
  LAYER M1 ;
        RECT 8.719 15.624 8.721 18.06 ;
  LAYER M1 ;
        RECT 8.799 15.624 8.801 18.06 ;
  LAYER M2 ;
        RECT 6.48 15.623 8.88 15.625 ;
  LAYER M2 ;
        RECT 6.48 15.707 8.88 15.709 ;
  LAYER M2 ;
        RECT 6.48 15.791 8.88 15.793 ;
  LAYER M2 ;
        RECT 6.48 15.875 8.88 15.877 ;
  LAYER M2 ;
        RECT 6.48 15.959 8.88 15.961 ;
  LAYER M2 ;
        RECT 6.48 16.043 8.88 16.045 ;
  LAYER M2 ;
        RECT 6.48 16.127 8.88 16.129 ;
  LAYER M2 ;
        RECT 6.48 16.211 8.88 16.213 ;
  LAYER M2 ;
        RECT 6.48 16.295 8.88 16.297 ;
  LAYER M2 ;
        RECT 6.48 16.379 8.88 16.381 ;
  LAYER M2 ;
        RECT 6.48 16.463 8.88 16.465 ;
  LAYER M2 ;
        RECT 6.48 16.547 8.88 16.549 ;
  LAYER M2 ;
        RECT 6.48 16.6305 8.88 16.6325 ;
  LAYER M2 ;
        RECT 6.48 16.715 8.88 16.717 ;
  LAYER M2 ;
        RECT 6.48 16.799 8.88 16.801 ;
  LAYER M2 ;
        RECT 6.48 16.883 8.88 16.885 ;
  LAYER M2 ;
        RECT 6.48 16.967 8.88 16.969 ;
  LAYER M2 ;
        RECT 6.48 17.051 8.88 17.053 ;
  LAYER M2 ;
        RECT 6.48 17.135 8.88 17.137 ;
  LAYER M2 ;
        RECT 6.48 17.219 8.88 17.221 ;
  LAYER M2 ;
        RECT 6.48 17.303 8.88 17.305 ;
  LAYER M2 ;
        RECT 6.48 17.387 8.88 17.389 ;
  LAYER M2 ;
        RECT 6.48 17.471 8.88 17.473 ;
  LAYER M2 ;
        RECT 6.48 17.555 8.88 17.557 ;
  LAYER M2 ;
        RECT 6.48 17.639 8.88 17.641 ;
  LAYER M2 ;
        RECT 6.48 17.723 8.88 17.725 ;
  LAYER M2 ;
        RECT 6.48 17.807 8.88 17.809 ;
  LAYER M2 ;
        RECT 6.48 17.891 8.88 17.893 ;
  LAYER M2 ;
        RECT 6.48 17.975 8.88 17.977 ;
  LAYER M1 ;
        RECT 6.464 18.528 6.496 21.036 ;
  LAYER M1 ;
        RECT 6.528 18.528 6.56 21.036 ;
  LAYER M1 ;
        RECT 6.592 18.528 6.624 21.036 ;
  LAYER M1 ;
        RECT 6.656 18.528 6.688 21.036 ;
  LAYER M1 ;
        RECT 6.72 18.528 6.752 21.036 ;
  LAYER M1 ;
        RECT 6.784 18.528 6.816 21.036 ;
  LAYER M1 ;
        RECT 6.848 18.528 6.88 21.036 ;
  LAYER M1 ;
        RECT 6.912 18.528 6.944 21.036 ;
  LAYER M1 ;
        RECT 6.976 18.528 7.008 21.036 ;
  LAYER M1 ;
        RECT 7.04 18.528 7.072 21.036 ;
  LAYER M1 ;
        RECT 7.104 18.528 7.136 21.036 ;
  LAYER M1 ;
        RECT 7.168 18.528 7.2 21.036 ;
  LAYER M1 ;
        RECT 7.232 18.528 7.264 21.036 ;
  LAYER M1 ;
        RECT 7.296 18.528 7.328 21.036 ;
  LAYER M1 ;
        RECT 7.36 18.528 7.392 21.036 ;
  LAYER M1 ;
        RECT 7.424 18.528 7.456 21.036 ;
  LAYER M1 ;
        RECT 7.488 18.528 7.52 21.036 ;
  LAYER M1 ;
        RECT 7.552 18.528 7.584 21.036 ;
  LAYER M1 ;
        RECT 7.616 18.528 7.648 21.036 ;
  LAYER M1 ;
        RECT 7.68 18.528 7.712 21.036 ;
  LAYER M1 ;
        RECT 7.744 18.528 7.776 21.036 ;
  LAYER M1 ;
        RECT 7.808 18.528 7.84 21.036 ;
  LAYER M1 ;
        RECT 7.872 18.528 7.904 21.036 ;
  LAYER M1 ;
        RECT 7.936 18.528 7.968 21.036 ;
  LAYER M1 ;
        RECT 8 18.528 8.032 21.036 ;
  LAYER M1 ;
        RECT 8.064 18.528 8.096 21.036 ;
  LAYER M1 ;
        RECT 8.128 18.528 8.16 21.036 ;
  LAYER M1 ;
        RECT 8.192 18.528 8.224 21.036 ;
  LAYER M1 ;
        RECT 8.256 18.528 8.288 21.036 ;
  LAYER M1 ;
        RECT 8.32 18.528 8.352 21.036 ;
  LAYER M1 ;
        RECT 8.384 18.528 8.416 21.036 ;
  LAYER M1 ;
        RECT 8.448 18.528 8.48 21.036 ;
  LAYER M1 ;
        RECT 8.512 18.528 8.544 21.036 ;
  LAYER M1 ;
        RECT 8.576 18.528 8.608 21.036 ;
  LAYER M1 ;
        RECT 8.64 18.528 8.672 21.036 ;
  LAYER M1 ;
        RECT 8.704 18.528 8.736 21.036 ;
  LAYER M1 ;
        RECT 8.768 18.528 8.8 21.036 ;
  LAYER M2 ;
        RECT 6.444 18.612 8.916 18.644 ;
  LAYER M2 ;
        RECT 6.444 18.676 8.916 18.708 ;
  LAYER M2 ;
        RECT 6.444 18.74 8.916 18.772 ;
  LAYER M2 ;
        RECT 6.444 18.804 8.916 18.836 ;
  LAYER M2 ;
        RECT 6.444 18.868 8.916 18.9 ;
  LAYER M2 ;
        RECT 6.444 18.932 8.916 18.964 ;
  LAYER M2 ;
        RECT 6.444 18.996 8.916 19.028 ;
  LAYER M2 ;
        RECT 6.444 19.06 8.916 19.092 ;
  LAYER M2 ;
        RECT 6.444 19.124 8.916 19.156 ;
  LAYER M2 ;
        RECT 6.444 19.188 8.916 19.22 ;
  LAYER M2 ;
        RECT 6.444 19.252 8.916 19.284 ;
  LAYER M2 ;
        RECT 6.444 19.316 8.916 19.348 ;
  LAYER M2 ;
        RECT 6.444 19.38 8.916 19.412 ;
  LAYER M2 ;
        RECT 6.444 19.444 8.916 19.476 ;
  LAYER M2 ;
        RECT 6.444 19.508 8.916 19.54 ;
  LAYER M2 ;
        RECT 6.444 19.572 8.916 19.604 ;
  LAYER M2 ;
        RECT 6.444 19.636 8.916 19.668 ;
  LAYER M2 ;
        RECT 6.444 19.7 8.916 19.732 ;
  LAYER M2 ;
        RECT 6.444 19.764 8.916 19.796 ;
  LAYER M2 ;
        RECT 6.444 19.828 8.916 19.86 ;
  LAYER M2 ;
        RECT 6.444 19.892 8.916 19.924 ;
  LAYER M2 ;
        RECT 6.444 19.956 8.916 19.988 ;
  LAYER M2 ;
        RECT 6.444 20.02 8.916 20.052 ;
  LAYER M2 ;
        RECT 6.444 20.084 8.916 20.116 ;
  LAYER M2 ;
        RECT 6.444 20.148 8.916 20.18 ;
  LAYER M2 ;
        RECT 6.444 20.212 8.916 20.244 ;
  LAYER M2 ;
        RECT 6.444 20.276 8.916 20.308 ;
  LAYER M2 ;
        RECT 6.444 20.34 8.916 20.372 ;
  LAYER M2 ;
        RECT 6.444 20.404 8.916 20.436 ;
  LAYER M2 ;
        RECT 6.444 20.468 8.916 20.5 ;
  LAYER M2 ;
        RECT 6.444 20.532 8.916 20.564 ;
  LAYER M2 ;
        RECT 6.444 20.596 8.916 20.628 ;
  LAYER M2 ;
        RECT 6.444 20.66 8.916 20.692 ;
  LAYER M2 ;
        RECT 6.444 20.724 8.916 20.756 ;
  LAYER M2 ;
        RECT 6.444 20.788 8.916 20.82 ;
  LAYER M2 ;
        RECT 6.444 20.852 8.916 20.884 ;
  LAYER M3 ;
        RECT 6.464 18.528 6.496 21.036 ;
  LAYER M3 ;
        RECT 6.528 18.528 6.56 21.036 ;
  LAYER M3 ;
        RECT 6.592 18.528 6.624 21.036 ;
  LAYER M3 ;
        RECT 6.656 18.528 6.688 21.036 ;
  LAYER M3 ;
        RECT 6.72 18.528 6.752 21.036 ;
  LAYER M3 ;
        RECT 6.784 18.528 6.816 21.036 ;
  LAYER M3 ;
        RECT 6.848 18.528 6.88 21.036 ;
  LAYER M3 ;
        RECT 6.912 18.528 6.944 21.036 ;
  LAYER M3 ;
        RECT 6.976 18.528 7.008 21.036 ;
  LAYER M3 ;
        RECT 7.04 18.528 7.072 21.036 ;
  LAYER M3 ;
        RECT 7.104 18.528 7.136 21.036 ;
  LAYER M3 ;
        RECT 7.168 18.528 7.2 21.036 ;
  LAYER M3 ;
        RECT 7.232 18.528 7.264 21.036 ;
  LAYER M3 ;
        RECT 7.296 18.528 7.328 21.036 ;
  LAYER M3 ;
        RECT 7.36 18.528 7.392 21.036 ;
  LAYER M3 ;
        RECT 7.424 18.528 7.456 21.036 ;
  LAYER M3 ;
        RECT 7.488 18.528 7.52 21.036 ;
  LAYER M3 ;
        RECT 7.552 18.528 7.584 21.036 ;
  LAYER M3 ;
        RECT 7.616 18.528 7.648 21.036 ;
  LAYER M3 ;
        RECT 7.68 18.528 7.712 21.036 ;
  LAYER M3 ;
        RECT 7.744 18.528 7.776 21.036 ;
  LAYER M3 ;
        RECT 7.808 18.528 7.84 21.036 ;
  LAYER M3 ;
        RECT 7.872 18.528 7.904 21.036 ;
  LAYER M3 ;
        RECT 7.936 18.528 7.968 21.036 ;
  LAYER M3 ;
        RECT 8 18.528 8.032 21.036 ;
  LAYER M3 ;
        RECT 8.064 18.528 8.096 21.036 ;
  LAYER M3 ;
        RECT 8.128 18.528 8.16 21.036 ;
  LAYER M3 ;
        RECT 8.192 18.528 8.224 21.036 ;
  LAYER M3 ;
        RECT 8.256 18.528 8.288 21.036 ;
  LAYER M3 ;
        RECT 8.32 18.528 8.352 21.036 ;
  LAYER M3 ;
        RECT 8.384 18.528 8.416 21.036 ;
  LAYER M3 ;
        RECT 8.448 18.528 8.48 21.036 ;
  LAYER M3 ;
        RECT 8.512 18.528 8.544 21.036 ;
  LAYER M3 ;
        RECT 8.576 18.528 8.608 21.036 ;
  LAYER M3 ;
        RECT 8.64 18.528 8.672 21.036 ;
  LAYER M3 ;
        RECT 8.704 18.528 8.736 21.036 ;
  LAYER M3 ;
        RECT 8.768 18.528 8.8 21.036 ;
  LAYER M3 ;
        RECT 8.864 18.528 8.896 21.036 ;
  LAYER M1 ;
        RECT 6.479 18.564 6.481 21 ;
  LAYER M1 ;
        RECT 6.559 18.564 6.561 21 ;
  LAYER M1 ;
        RECT 6.639 18.564 6.641 21 ;
  LAYER M1 ;
        RECT 6.719 18.564 6.721 21 ;
  LAYER M1 ;
        RECT 6.799 18.564 6.801 21 ;
  LAYER M1 ;
        RECT 6.879 18.564 6.881 21 ;
  LAYER M1 ;
        RECT 6.959 18.564 6.961 21 ;
  LAYER M1 ;
        RECT 7.039 18.564 7.041 21 ;
  LAYER M1 ;
        RECT 7.119 18.564 7.121 21 ;
  LAYER M1 ;
        RECT 7.199 18.564 7.201 21 ;
  LAYER M1 ;
        RECT 7.279 18.564 7.281 21 ;
  LAYER M1 ;
        RECT 7.359 18.564 7.361 21 ;
  LAYER M1 ;
        RECT 7.439 18.564 7.441 21 ;
  LAYER M1 ;
        RECT 7.519 18.564 7.521 21 ;
  LAYER M1 ;
        RECT 7.599 18.564 7.601 21 ;
  LAYER M1 ;
        RECT 7.679 18.564 7.681 21 ;
  LAYER M1 ;
        RECT 7.759 18.564 7.761 21 ;
  LAYER M1 ;
        RECT 7.839 18.564 7.841 21 ;
  LAYER M1 ;
        RECT 7.919 18.564 7.921 21 ;
  LAYER M1 ;
        RECT 7.999 18.564 8.001 21 ;
  LAYER M1 ;
        RECT 8.079 18.564 8.081 21 ;
  LAYER M1 ;
        RECT 8.159 18.564 8.161 21 ;
  LAYER M1 ;
        RECT 8.239 18.564 8.241 21 ;
  LAYER M1 ;
        RECT 8.319 18.564 8.321 21 ;
  LAYER M1 ;
        RECT 8.399 18.564 8.401 21 ;
  LAYER M1 ;
        RECT 8.479 18.564 8.481 21 ;
  LAYER M1 ;
        RECT 8.559 18.564 8.561 21 ;
  LAYER M1 ;
        RECT 8.639 18.564 8.641 21 ;
  LAYER M1 ;
        RECT 8.719 18.564 8.721 21 ;
  LAYER M1 ;
        RECT 8.799 18.564 8.801 21 ;
  LAYER M2 ;
        RECT 6.48 18.563 8.88 18.565 ;
  LAYER M2 ;
        RECT 6.48 18.647 8.88 18.649 ;
  LAYER M2 ;
        RECT 6.48 18.731 8.88 18.733 ;
  LAYER M2 ;
        RECT 6.48 18.815 8.88 18.817 ;
  LAYER M2 ;
        RECT 6.48 18.899 8.88 18.901 ;
  LAYER M2 ;
        RECT 6.48 18.983 8.88 18.985 ;
  LAYER M2 ;
        RECT 6.48 19.067 8.88 19.069 ;
  LAYER M2 ;
        RECT 6.48 19.151 8.88 19.153 ;
  LAYER M2 ;
        RECT 6.48 19.235 8.88 19.237 ;
  LAYER M2 ;
        RECT 6.48 19.319 8.88 19.321 ;
  LAYER M2 ;
        RECT 6.48 19.403 8.88 19.405 ;
  LAYER M2 ;
        RECT 6.48 19.487 8.88 19.489 ;
  LAYER M2 ;
        RECT 6.48 19.5705 8.88 19.5725 ;
  LAYER M2 ;
        RECT 6.48 19.655 8.88 19.657 ;
  LAYER M2 ;
        RECT 6.48 19.739 8.88 19.741 ;
  LAYER M2 ;
        RECT 6.48 19.823 8.88 19.825 ;
  LAYER M2 ;
        RECT 6.48 19.907 8.88 19.909 ;
  LAYER M2 ;
        RECT 6.48 19.991 8.88 19.993 ;
  LAYER M2 ;
        RECT 6.48 20.075 8.88 20.077 ;
  LAYER M2 ;
        RECT 6.48 20.159 8.88 20.161 ;
  LAYER M2 ;
        RECT 6.48 20.243 8.88 20.245 ;
  LAYER M2 ;
        RECT 6.48 20.327 8.88 20.329 ;
  LAYER M2 ;
        RECT 6.48 20.411 8.88 20.413 ;
  LAYER M2 ;
        RECT 6.48 20.495 8.88 20.497 ;
  LAYER M2 ;
        RECT 6.48 20.579 8.88 20.581 ;
  LAYER M2 ;
        RECT 6.48 20.663 8.88 20.665 ;
  LAYER M2 ;
        RECT 6.48 20.747 8.88 20.749 ;
  LAYER M2 ;
        RECT 6.48 20.831 8.88 20.833 ;
  LAYER M2 ;
        RECT 6.48 20.915 8.88 20.917 ;
  LAYER M1 ;
        RECT 9.664 0.888 9.696 3.396 ;
  LAYER M1 ;
        RECT 9.728 0.888 9.76 3.396 ;
  LAYER M1 ;
        RECT 9.792 0.888 9.824 3.396 ;
  LAYER M1 ;
        RECT 9.856 0.888 9.888 3.396 ;
  LAYER M1 ;
        RECT 9.92 0.888 9.952 3.396 ;
  LAYER M1 ;
        RECT 9.984 0.888 10.016 3.396 ;
  LAYER M1 ;
        RECT 10.048 0.888 10.08 3.396 ;
  LAYER M1 ;
        RECT 10.112 0.888 10.144 3.396 ;
  LAYER M1 ;
        RECT 10.176 0.888 10.208 3.396 ;
  LAYER M1 ;
        RECT 10.24 0.888 10.272 3.396 ;
  LAYER M1 ;
        RECT 10.304 0.888 10.336 3.396 ;
  LAYER M1 ;
        RECT 10.368 0.888 10.4 3.396 ;
  LAYER M1 ;
        RECT 10.432 0.888 10.464 3.396 ;
  LAYER M1 ;
        RECT 10.496 0.888 10.528 3.396 ;
  LAYER M1 ;
        RECT 10.56 0.888 10.592 3.396 ;
  LAYER M1 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M1 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M1 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M1 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M1 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M1 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M1 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M1 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M1 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M1 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M1 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M1 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M1 ;
        RECT 11.392 0.888 11.424 3.396 ;
  LAYER M1 ;
        RECT 11.456 0.888 11.488 3.396 ;
  LAYER M1 ;
        RECT 11.52 0.888 11.552 3.396 ;
  LAYER M1 ;
        RECT 11.584 0.888 11.616 3.396 ;
  LAYER M1 ;
        RECT 11.648 0.888 11.68 3.396 ;
  LAYER M1 ;
        RECT 11.712 0.888 11.744 3.396 ;
  LAYER M1 ;
        RECT 11.776 0.888 11.808 3.396 ;
  LAYER M1 ;
        RECT 11.84 0.888 11.872 3.396 ;
  LAYER M1 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M1 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M2 ;
        RECT 9.644 0.972 12.116 1.004 ;
  LAYER M2 ;
        RECT 9.644 1.036 12.116 1.068 ;
  LAYER M2 ;
        RECT 9.644 1.1 12.116 1.132 ;
  LAYER M2 ;
        RECT 9.644 1.164 12.116 1.196 ;
  LAYER M2 ;
        RECT 9.644 1.228 12.116 1.26 ;
  LAYER M2 ;
        RECT 9.644 1.292 12.116 1.324 ;
  LAYER M2 ;
        RECT 9.644 1.356 12.116 1.388 ;
  LAYER M2 ;
        RECT 9.644 1.42 12.116 1.452 ;
  LAYER M2 ;
        RECT 9.644 1.484 12.116 1.516 ;
  LAYER M2 ;
        RECT 9.644 1.548 12.116 1.58 ;
  LAYER M2 ;
        RECT 9.644 1.612 12.116 1.644 ;
  LAYER M2 ;
        RECT 9.644 1.676 12.116 1.708 ;
  LAYER M2 ;
        RECT 9.644 1.74 12.116 1.772 ;
  LAYER M2 ;
        RECT 9.644 1.804 12.116 1.836 ;
  LAYER M2 ;
        RECT 9.644 1.868 12.116 1.9 ;
  LAYER M2 ;
        RECT 9.644 1.932 12.116 1.964 ;
  LAYER M2 ;
        RECT 9.644 1.996 12.116 2.028 ;
  LAYER M2 ;
        RECT 9.644 2.06 12.116 2.092 ;
  LAYER M2 ;
        RECT 9.644 2.124 12.116 2.156 ;
  LAYER M2 ;
        RECT 9.644 2.188 12.116 2.22 ;
  LAYER M2 ;
        RECT 9.644 2.252 12.116 2.284 ;
  LAYER M2 ;
        RECT 9.644 2.316 12.116 2.348 ;
  LAYER M2 ;
        RECT 9.644 2.38 12.116 2.412 ;
  LAYER M2 ;
        RECT 9.644 2.444 12.116 2.476 ;
  LAYER M2 ;
        RECT 9.644 2.508 12.116 2.54 ;
  LAYER M2 ;
        RECT 9.644 2.572 12.116 2.604 ;
  LAYER M2 ;
        RECT 9.644 2.636 12.116 2.668 ;
  LAYER M2 ;
        RECT 9.644 2.7 12.116 2.732 ;
  LAYER M2 ;
        RECT 9.644 2.764 12.116 2.796 ;
  LAYER M2 ;
        RECT 9.644 2.828 12.116 2.86 ;
  LAYER M2 ;
        RECT 9.644 2.892 12.116 2.924 ;
  LAYER M2 ;
        RECT 9.644 2.956 12.116 2.988 ;
  LAYER M2 ;
        RECT 9.644 3.02 12.116 3.052 ;
  LAYER M2 ;
        RECT 9.644 3.084 12.116 3.116 ;
  LAYER M2 ;
        RECT 9.644 3.148 12.116 3.18 ;
  LAYER M2 ;
        RECT 9.644 3.212 12.116 3.244 ;
  LAYER M3 ;
        RECT 9.664 0.888 9.696 3.396 ;
  LAYER M3 ;
        RECT 9.728 0.888 9.76 3.396 ;
  LAYER M3 ;
        RECT 9.792 0.888 9.824 3.396 ;
  LAYER M3 ;
        RECT 9.856 0.888 9.888 3.396 ;
  LAYER M3 ;
        RECT 9.92 0.888 9.952 3.396 ;
  LAYER M3 ;
        RECT 9.984 0.888 10.016 3.396 ;
  LAYER M3 ;
        RECT 10.048 0.888 10.08 3.396 ;
  LAYER M3 ;
        RECT 10.112 0.888 10.144 3.396 ;
  LAYER M3 ;
        RECT 10.176 0.888 10.208 3.396 ;
  LAYER M3 ;
        RECT 10.24 0.888 10.272 3.396 ;
  LAYER M3 ;
        RECT 10.304 0.888 10.336 3.396 ;
  LAYER M3 ;
        RECT 10.368 0.888 10.4 3.396 ;
  LAYER M3 ;
        RECT 10.432 0.888 10.464 3.396 ;
  LAYER M3 ;
        RECT 10.496 0.888 10.528 3.396 ;
  LAYER M3 ;
        RECT 10.56 0.888 10.592 3.396 ;
  LAYER M3 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M3 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M3 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M3 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M3 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M3 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M3 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M3 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M3 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M3 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M3 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M3 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M3 ;
        RECT 11.392 0.888 11.424 3.396 ;
  LAYER M3 ;
        RECT 11.456 0.888 11.488 3.396 ;
  LAYER M3 ;
        RECT 11.52 0.888 11.552 3.396 ;
  LAYER M3 ;
        RECT 11.584 0.888 11.616 3.396 ;
  LAYER M3 ;
        RECT 11.648 0.888 11.68 3.396 ;
  LAYER M3 ;
        RECT 11.712 0.888 11.744 3.396 ;
  LAYER M3 ;
        RECT 11.776 0.888 11.808 3.396 ;
  LAYER M3 ;
        RECT 11.84 0.888 11.872 3.396 ;
  LAYER M3 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M3 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M3 ;
        RECT 12.064 0.888 12.096 3.396 ;
  LAYER M1 ;
        RECT 9.679 0.924 9.681 3.36 ;
  LAYER M1 ;
        RECT 9.759 0.924 9.761 3.36 ;
  LAYER M1 ;
        RECT 9.839 0.924 9.841 3.36 ;
  LAYER M1 ;
        RECT 9.919 0.924 9.921 3.36 ;
  LAYER M1 ;
        RECT 9.999 0.924 10.001 3.36 ;
  LAYER M1 ;
        RECT 10.079 0.924 10.081 3.36 ;
  LAYER M1 ;
        RECT 10.159 0.924 10.161 3.36 ;
  LAYER M1 ;
        RECT 10.239 0.924 10.241 3.36 ;
  LAYER M1 ;
        RECT 10.319 0.924 10.321 3.36 ;
  LAYER M1 ;
        RECT 10.399 0.924 10.401 3.36 ;
  LAYER M1 ;
        RECT 10.479 0.924 10.481 3.36 ;
  LAYER M1 ;
        RECT 10.559 0.924 10.561 3.36 ;
  LAYER M1 ;
        RECT 10.639 0.924 10.641 3.36 ;
  LAYER M1 ;
        RECT 10.719 0.924 10.721 3.36 ;
  LAYER M1 ;
        RECT 10.799 0.924 10.801 3.36 ;
  LAYER M1 ;
        RECT 10.879 0.924 10.881 3.36 ;
  LAYER M1 ;
        RECT 10.959 0.924 10.961 3.36 ;
  LAYER M1 ;
        RECT 11.039 0.924 11.041 3.36 ;
  LAYER M1 ;
        RECT 11.119 0.924 11.121 3.36 ;
  LAYER M1 ;
        RECT 11.199 0.924 11.201 3.36 ;
  LAYER M1 ;
        RECT 11.279 0.924 11.281 3.36 ;
  LAYER M1 ;
        RECT 11.359 0.924 11.361 3.36 ;
  LAYER M1 ;
        RECT 11.439 0.924 11.441 3.36 ;
  LAYER M1 ;
        RECT 11.519 0.924 11.521 3.36 ;
  LAYER M1 ;
        RECT 11.599 0.924 11.601 3.36 ;
  LAYER M1 ;
        RECT 11.679 0.924 11.681 3.36 ;
  LAYER M1 ;
        RECT 11.759 0.924 11.761 3.36 ;
  LAYER M1 ;
        RECT 11.839 0.924 11.841 3.36 ;
  LAYER M1 ;
        RECT 11.919 0.924 11.921 3.36 ;
  LAYER M1 ;
        RECT 11.999 0.924 12.001 3.36 ;
  LAYER M2 ;
        RECT 9.68 0.923 12.08 0.925 ;
  LAYER M2 ;
        RECT 9.68 1.007 12.08 1.009 ;
  LAYER M2 ;
        RECT 9.68 1.091 12.08 1.093 ;
  LAYER M2 ;
        RECT 9.68 1.175 12.08 1.177 ;
  LAYER M2 ;
        RECT 9.68 1.259 12.08 1.261 ;
  LAYER M2 ;
        RECT 9.68 1.343 12.08 1.345 ;
  LAYER M2 ;
        RECT 9.68 1.427 12.08 1.429 ;
  LAYER M2 ;
        RECT 9.68 1.511 12.08 1.513 ;
  LAYER M2 ;
        RECT 9.68 1.595 12.08 1.597 ;
  LAYER M2 ;
        RECT 9.68 1.679 12.08 1.681 ;
  LAYER M2 ;
        RECT 9.68 1.763 12.08 1.765 ;
  LAYER M2 ;
        RECT 9.68 1.847 12.08 1.849 ;
  LAYER M2 ;
        RECT 9.68 1.9305 12.08 1.9325 ;
  LAYER M2 ;
        RECT 9.68 2.015 12.08 2.017 ;
  LAYER M2 ;
        RECT 9.68 2.099 12.08 2.101 ;
  LAYER M2 ;
        RECT 9.68 2.183 12.08 2.185 ;
  LAYER M2 ;
        RECT 9.68 2.267 12.08 2.269 ;
  LAYER M2 ;
        RECT 9.68 2.351 12.08 2.353 ;
  LAYER M2 ;
        RECT 9.68 2.435 12.08 2.437 ;
  LAYER M2 ;
        RECT 9.68 2.519 12.08 2.521 ;
  LAYER M2 ;
        RECT 9.68 2.603 12.08 2.605 ;
  LAYER M2 ;
        RECT 9.68 2.687 12.08 2.689 ;
  LAYER M2 ;
        RECT 9.68 2.771 12.08 2.773 ;
  LAYER M2 ;
        RECT 9.68 2.855 12.08 2.857 ;
  LAYER M2 ;
        RECT 9.68 2.939 12.08 2.941 ;
  LAYER M2 ;
        RECT 9.68 3.023 12.08 3.025 ;
  LAYER M2 ;
        RECT 9.68 3.107 12.08 3.109 ;
  LAYER M2 ;
        RECT 9.68 3.191 12.08 3.193 ;
  LAYER M2 ;
        RECT 9.68 3.275 12.08 3.277 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 6.336 ;
  LAYER M1 ;
        RECT 9.728 3.828 9.76 6.336 ;
  LAYER M1 ;
        RECT 9.792 3.828 9.824 6.336 ;
  LAYER M1 ;
        RECT 9.856 3.828 9.888 6.336 ;
  LAYER M1 ;
        RECT 9.92 3.828 9.952 6.336 ;
  LAYER M1 ;
        RECT 9.984 3.828 10.016 6.336 ;
  LAYER M1 ;
        RECT 10.048 3.828 10.08 6.336 ;
  LAYER M1 ;
        RECT 10.112 3.828 10.144 6.336 ;
  LAYER M1 ;
        RECT 10.176 3.828 10.208 6.336 ;
  LAYER M1 ;
        RECT 10.24 3.828 10.272 6.336 ;
  LAYER M1 ;
        RECT 10.304 3.828 10.336 6.336 ;
  LAYER M1 ;
        RECT 10.368 3.828 10.4 6.336 ;
  LAYER M1 ;
        RECT 10.432 3.828 10.464 6.336 ;
  LAYER M1 ;
        RECT 10.496 3.828 10.528 6.336 ;
  LAYER M1 ;
        RECT 10.56 3.828 10.592 6.336 ;
  LAYER M1 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M1 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M1 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M1 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M1 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M1 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M1 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M1 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M1 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M1 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M1 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M1 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M1 ;
        RECT 11.392 3.828 11.424 6.336 ;
  LAYER M1 ;
        RECT 11.456 3.828 11.488 6.336 ;
  LAYER M1 ;
        RECT 11.52 3.828 11.552 6.336 ;
  LAYER M1 ;
        RECT 11.584 3.828 11.616 6.336 ;
  LAYER M1 ;
        RECT 11.648 3.828 11.68 6.336 ;
  LAYER M1 ;
        RECT 11.712 3.828 11.744 6.336 ;
  LAYER M1 ;
        RECT 11.776 3.828 11.808 6.336 ;
  LAYER M1 ;
        RECT 11.84 3.828 11.872 6.336 ;
  LAYER M1 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M1 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M2 ;
        RECT 9.644 3.912 12.116 3.944 ;
  LAYER M2 ;
        RECT 9.644 3.976 12.116 4.008 ;
  LAYER M2 ;
        RECT 9.644 4.04 12.116 4.072 ;
  LAYER M2 ;
        RECT 9.644 4.104 12.116 4.136 ;
  LAYER M2 ;
        RECT 9.644 4.168 12.116 4.2 ;
  LAYER M2 ;
        RECT 9.644 4.232 12.116 4.264 ;
  LAYER M2 ;
        RECT 9.644 4.296 12.116 4.328 ;
  LAYER M2 ;
        RECT 9.644 4.36 12.116 4.392 ;
  LAYER M2 ;
        RECT 9.644 4.424 12.116 4.456 ;
  LAYER M2 ;
        RECT 9.644 4.488 12.116 4.52 ;
  LAYER M2 ;
        RECT 9.644 4.552 12.116 4.584 ;
  LAYER M2 ;
        RECT 9.644 4.616 12.116 4.648 ;
  LAYER M2 ;
        RECT 9.644 4.68 12.116 4.712 ;
  LAYER M2 ;
        RECT 9.644 4.744 12.116 4.776 ;
  LAYER M2 ;
        RECT 9.644 4.808 12.116 4.84 ;
  LAYER M2 ;
        RECT 9.644 4.872 12.116 4.904 ;
  LAYER M2 ;
        RECT 9.644 4.936 12.116 4.968 ;
  LAYER M2 ;
        RECT 9.644 5 12.116 5.032 ;
  LAYER M2 ;
        RECT 9.644 5.064 12.116 5.096 ;
  LAYER M2 ;
        RECT 9.644 5.128 12.116 5.16 ;
  LAYER M2 ;
        RECT 9.644 5.192 12.116 5.224 ;
  LAYER M2 ;
        RECT 9.644 5.256 12.116 5.288 ;
  LAYER M2 ;
        RECT 9.644 5.32 12.116 5.352 ;
  LAYER M2 ;
        RECT 9.644 5.384 12.116 5.416 ;
  LAYER M2 ;
        RECT 9.644 5.448 12.116 5.48 ;
  LAYER M2 ;
        RECT 9.644 5.512 12.116 5.544 ;
  LAYER M2 ;
        RECT 9.644 5.576 12.116 5.608 ;
  LAYER M2 ;
        RECT 9.644 5.64 12.116 5.672 ;
  LAYER M2 ;
        RECT 9.644 5.704 12.116 5.736 ;
  LAYER M2 ;
        RECT 9.644 5.768 12.116 5.8 ;
  LAYER M2 ;
        RECT 9.644 5.832 12.116 5.864 ;
  LAYER M2 ;
        RECT 9.644 5.896 12.116 5.928 ;
  LAYER M2 ;
        RECT 9.644 5.96 12.116 5.992 ;
  LAYER M2 ;
        RECT 9.644 6.024 12.116 6.056 ;
  LAYER M2 ;
        RECT 9.644 6.088 12.116 6.12 ;
  LAYER M2 ;
        RECT 9.644 6.152 12.116 6.184 ;
  LAYER M3 ;
        RECT 9.664 3.828 9.696 6.336 ;
  LAYER M3 ;
        RECT 9.728 3.828 9.76 6.336 ;
  LAYER M3 ;
        RECT 9.792 3.828 9.824 6.336 ;
  LAYER M3 ;
        RECT 9.856 3.828 9.888 6.336 ;
  LAYER M3 ;
        RECT 9.92 3.828 9.952 6.336 ;
  LAYER M3 ;
        RECT 9.984 3.828 10.016 6.336 ;
  LAYER M3 ;
        RECT 10.048 3.828 10.08 6.336 ;
  LAYER M3 ;
        RECT 10.112 3.828 10.144 6.336 ;
  LAYER M3 ;
        RECT 10.176 3.828 10.208 6.336 ;
  LAYER M3 ;
        RECT 10.24 3.828 10.272 6.336 ;
  LAYER M3 ;
        RECT 10.304 3.828 10.336 6.336 ;
  LAYER M3 ;
        RECT 10.368 3.828 10.4 6.336 ;
  LAYER M3 ;
        RECT 10.432 3.828 10.464 6.336 ;
  LAYER M3 ;
        RECT 10.496 3.828 10.528 6.336 ;
  LAYER M3 ;
        RECT 10.56 3.828 10.592 6.336 ;
  LAYER M3 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M3 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M3 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M3 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M3 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M3 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M3 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M3 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M3 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M3 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M3 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M3 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M3 ;
        RECT 11.392 3.828 11.424 6.336 ;
  LAYER M3 ;
        RECT 11.456 3.828 11.488 6.336 ;
  LAYER M3 ;
        RECT 11.52 3.828 11.552 6.336 ;
  LAYER M3 ;
        RECT 11.584 3.828 11.616 6.336 ;
  LAYER M3 ;
        RECT 11.648 3.828 11.68 6.336 ;
  LAYER M3 ;
        RECT 11.712 3.828 11.744 6.336 ;
  LAYER M3 ;
        RECT 11.776 3.828 11.808 6.336 ;
  LAYER M3 ;
        RECT 11.84 3.828 11.872 6.336 ;
  LAYER M3 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M3 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M3 ;
        RECT 12.064 3.828 12.096 6.336 ;
  LAYER M1 ;
        RECT 9.679 3.864 9.681 6.3 ;
  LAYER M1 ;
        RECT 9.759 3.864 9.761 6.3 ;
  LAYER M1 ;
        RECT 9.839 3.864 9.841 6.3 ;
  LAYER M1 ;
        RECT 9.919 3.864 9.921 6.3 ;
  LAYER M1 ;
        RECT 9.999 3.864 10.001 6.3 ;
  LAYER M1 ;
        RECT 10.079 3.864 10.081 6.3 ;
  LAYER M1 ;
        RECT 10.159 3.864 10.161 6.3 ;
  LAYER M1 ;
        RECT 10.239 3.864 10.241 6.3 ;
  LAYER M1 ;
        RECT 10.319 3.864 10.321 6.3 ;
  LAYER M1 ;
        RECT 10.399 3.864 10.401 6.3 ;
  LAYER M1 ;
        RECT 10.479 3.864 10.481 6.3 ;
  LAYER M1 ;
        RECT 10.559 3.864 10.561 6.3 ;
  LAYER M1 ;
        RECT 10.639 3.864 10.641 6.3 ;
  LAYER M1 ;
        RECT 10.719 3.864 10.721 6.3 ;
  LAYER M1 ;
        RECT 10.799 3.864 10.801 6.3 ;
  LAYER M1 ;
        RECT 10.879 3.864 10.881 6.3 ;
  LAYER M1 ;
        RECT 10.959 3.864 10.961 6.3 ;
  LAYER M1 ;
        RECT 11.039 3.864 11.041 6.3 ;
  LAYER M1 ;
        RECT 11.119 3.864 11.121 6.3 ;
  LAYER M1 ;
        RECT 11.199 3.864 11.201 6.3 ;
  LAYER M1 ;
        RECT 11.279 3.864 11.281 6.3 ;
  LAYER M1 ;
        RECT 11.359 3.864 11.361 6.3 ;
  LAYER M1 ;
        RECT 11.439 3.864 11.441 6.3 ;
  LAYER M1 ;
        RECT 11.519 3.864 11.521 6.3 ;
  LAYER M1 ;
        RECT 11.599 3.864 11.601 6.3 ;
  LAYER M1 ;
        RECT 11.679 3.864 11.681 6.3 ;
  LAYER M1 ;
        RECT 11.759 3.864 11.761 6.3 ;
  LAYER M1 ;
        RECT 11.839 3.864 11.841 6.3 ;
  LAYER M1 ;
        RECT 11.919 3.864 11.921 6.3 ;
  LAYER M1 ;
        RECT 11.999 3.864 12.001 6.3 ;
  LAYER M2 ;
        RECT 9.68 3.863 12.08 3.865 ;
  LAYER M2 ;
        RECT 9.68 3.947 12.08 3.949 ;
  LAYER M2 ;
        RECT 9.68 4.031 12.08 4.033 ;
  LAYER M2 ;
        RECT 9.68 4.115 12.08 4.117 ;
  LAYER M2 ;
        RECT 9.68 4.199 12.08 4.201 ;
  LAYER M2 ;
        RECT 9.68 4.283 12.08 4.285 ;
  LAYER M2 ;
        RECT 9.68 4.367 12.08 4.369 ;
  LAYER M2 ;
        RECT 9.68 4.451 12.08 4.453 ;
  LAYER M2 ;
        RECT 9.68 4.535 12.08 4.537 ;
  LAYER M2 ;
        RECT 9.68 4.619 12.08 4.621 ;
  LAYER M2 ;
        RECT 9.68 4.703 12.08 4.705 ;
  LAYER M2 ;
        RECT 9.68 4.787 12.08 4.789 ;
  LAYER M2 ;
        RECT 9.68 4.8705 12.08 4.8725 ;
  LAYER M2 ;
        RECT 9.68 4.955 12.08 4.957 ;
  LAYER M2 ;
        RECT 9.68 5.039 12.08 5.041 ;
  LAYER M2 ;
        RECT 9.68 5.123 12.08 5.125 ;
  LAYER M2 ;
        RECT 9.68 5.207 12.08 5.209 ;
  LAYER M2 ;
        RECT 9.68 5.291 12.08 5.293 ;
  LAYER M2 ;
        RECT 9.68 5.375 12.08 5.377 ;
  LAYER M2 ;
        RECT 9.68 5.459 12.08 5.461 ;
  LAYER M2 ;
        RECT 9.68 5.543 12.08 5.545 ;
  LAYER M2 ;
        RECT 9.68 5.627 12.08 5.629 ;
  LAYER M2 ;
        RECT 9.68 5.711 12.08 5.713 ;
  LAYER M2 ;
        RECT 9.68 5.795 12.08 5.797 ;
  LAYER M2 ;
        RECT 9.68 5.879 12.08 5.881 ;
  LAYER M2 ;
        RECT 9.68 5.963 12.08 5.965 ;
  LAYER M2 ;
        RECT 9.68 6.047 12.08 6.049 ;
  LAYER M2 ;
        RECT 9.68 6.131 12.08 6.133 ;
  LAYER M2 ;
        RECT 9.68 6.215 12.08 6.217 ;
  LAYER M1 ;
        RECT 9.664 6.768 9.696 9.276 ;
  LAYER M1 ;
        RECT 9.728 6.768 9.76 9.276 ;
  LAYER M1 ;
        RECT 9.792 6.768 9.824 9.276 ;
  LAYER M1 ;
        RECT 9.856 6.768 9.888 9.276 ;
  LAYER M1 ;
        RECT 9.92 6.768 9.952 9.276 ;
  LAYER M1 ;
        RECT 9.984 6.768 10.016 9.276 ;
  LAYER M1 ;
        RECT 10.048 6.768 10.08 9.276 ;
  LAYER M1 ;
        RECT 10.112 6.768 10.144 9.276 ;
  LAYER M1 ;
        RECT 10.176 6.768 10.208 9.276 ;
  LAYER M1 ;
        RECT 10.24 6.768 10.272 9.276 ;
  LAYER M1 ;
        RECT 10.304 6.768 10.336 9.276 ;
  LAYER M1 ;
        RECT 10.368 6.768 10.4 9.276 ;
  LAYER M1 ;
        RECT 10.432 6.768 10.464 9.276 ;
  LAYER M1 ;
        RECT 10.496 6.768 10.528 9.276 ;
  LAYER M1 ;
        RECT 10.56 6.768 10.592 9.276 ;
  LAYER M1 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M1 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M1 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M1 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M1 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M1 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M1 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M1 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M1 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M1 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M1 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M1 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M1 ;
        RECT 11.392 6.768 11.424 9.276 ;
  LAYER M1 ;
        RECT 11.456 6.768 11.488 9.276 ;
  LAYER M1 ;
        RECT 11.52 6.768 11.552 9.276 ;
  LAYER M1 ;
        RECT 11.584 6.768 11.616 9.276 ;
  LAYER M1 ;
        RECT 11.648 6.768 11.68 9.276 ;
  LAYER M1 ;
        RECT 11.712 6.768 11.744 9.276 ;
  LAYER M1 ;
        RECT 11.776 6.768 11.808 9.276 ;
  LAYER M1 ;
        RECT 11.84 6.768 11.872 9.276 ;
  LAYER M1 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M1 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M2 ;
        RECT 9.644 6.852 12.116 6.884 ;
  LAYER M2 ;
        RECT 9.644 6.916 12.116 6.948 ;
  LAYER M2 ;
        RECT 9.644 6.98 12.116 7.012 ;
  LAYER M2 ;
        RECT 9.644 7.044 12.116 7.076 ;
  LAYER M2 ;
        RECT 9.644 7.108 12.116 7.14 ;
  LAYER M2 ;
        RECT 9.644 7.172 12.116 7.204 ;
  LAYER M2 ;
        RECT 9.644 7.236 12.116 7.268 ;
  LAYER M2 ;
        RECT 9.644 7.3 12.116 7.332 ;
  LAYER M2 ;
        RECT 9.644 7.364 12.116 7.396 ;
  LAYER M2 ;
        RECT 9.644 7.428 12.116 7.46 ;
  LAYER M2 ;
        RECT 9.644 7.492 12.116 7.524 ;
  LAYER M2 ;
        RECT 9.644 7.556 12.116 7.588 ;
  LAYER M2 ;
        RECT 9.644 7.62 12.116 7.652 ;
  LAYER M2 ;
        RECT 9.644 7.684 12.116 7.716 ;
  LAYER M2 ;
        RECT 9.644 7.748 12.116 7.78 ;
  LAYER M2 ;
        RECT 9.644 7.812 12.116 7.844 ;
  LAYER M2 ;
        RECT 9.644 7.876 12.116 7.908 ;
  LAYER M2 ;
        RECT 9.644 7.94 12.116 7.972 ;
  LAYER M2 ;
        RECT 9.644 8.004 12.116 8.036 ;
  LAYER M2 ;
        RECT 9.644 8.068 12.116 8.1 ;
  LAYER M2 ;
        RECT 9.644 8.132 12.116 8.164 ;
  LAYER M2 ;
        RECT 9.644 8.196 12.116 8.228 ;
  LAYER M2 ;
        RECT 9.644 8.26 12.116 8.292 ;
  LAYER M2 ;
        RECT 9.644 8.324 12.116 8.356 ;
  LAYER M2 ;
        RECT 9.644 8.388 12.116 8.42 ;
  LAYER M2 ;
        RECT 9.644 8.452 12.116 8.484 ;
  LAYER M2 ;
        RECT 9.644 8.516 12.116 8.548 ;
  LAYER M2 ;
        RECT 9.644 8.58 12.116 8.612 ;
  LAYER M2 ;
        RECT 9.644 8.644 12.116 8.676 ;
  LAYER M2 ;
        RECT 9.644 8.708 12.116 8.74 ;
  LAYER M2 ;
        RECT 9.644 8.772 12.116 8.804 ;
  LAYER M2 ;
        RECT 9.644 8.836 12.116 8.868 ;
  LAYER M2 ;
        RECT 9.644 8.9 12.116 8.932 ;
  LAYER M2 ;
        RECT 9.644 8.964 12.116 8.996 ;
  LAYER M2 ;
        RECT 9.644 9.028 12.116 9.06 ;
  LAYER M2 ;
        RECT 9.644 9.092 12.116 9.124 ;
  LAYER M3 ;
        RECT 9.664 6.768 9.696 9.276 ;
  LAYER M3 ;
        RECT 9.728 6.768 9.76 9.276 ;
  LAYER M3 ;
        RECT 9.792 6.768 9.824 9.276 ;
  LAYER M3 ;
        RECT 9.856 6.768 9.888 9.276 ;
  LAYER M3 ;
        RECT 9.92 6.768 9.952 9.276 ;
  LAYER M3 ;
        RECT 9.984 6.768 10.016 9.276 ;
  LAYER M3 ;
        RECT 10.048 6.768 10.08 9.276 ;
  LAYER M3 ;
        RECT 10.112 6.768 10.144 9.276 ;
  LAYER M3 ;
        RECT 10.176 6.768 10.208 9.276 ;
  LAYER M3 ;
        RECT 10.24 6.768 10.272 9.276 ;
  LAYER M3 ;
        RECT 10.304 6.768 10.336 9.276 ;
  LAYER M3 ;
        RECT 10.368 6.768 10.4 9.276 ;
  LAYER M3 ;
        RECT 10.432 6.768 10.464 9.276 ;
  LAYER M3 ;
        RECT 10.496 6.768 10.528 9.276 ;
  LAYER M3 ;
        RECT 10.56 6.768 10.592 9.276 ;
  LAYER M3 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M3 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M3 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M3 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M3 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M3 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M3 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M3 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M3 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M3 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M3 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M3 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M3 ;
        RECT 11.392 6.768 11.424 9.276 ;
  LAYER M3 ;
        RECT 11.456 6.768 11.488 9.276 ;
  LAYER M3 ;
        RECT 11.52 6.768 11.552 9.276 ;
  LAYER M3 ;
        RECT 11.584 6.768 11.616 9.276 ;
  LAYER M3 ;
        RECT 11.648 6.768 11.68 9.276 ;
  LAYER M3 ;
        RECT 11.712 6.768 11.744 9.276 ;
  LAYER M3 ;
        RECT 11.776 6.768 11.808 9.276 ;
  LAYER M3 ;
        RECT 11.84 6.768 11.872 9.276 ;
  LAYER M3 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M3 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M3 ;
        RECT 12.064 6.768 12.096 9.276 ;
  LAYER M1 ;
        RECT 9.679 6.804 9.681 9.24 ;
  LAYER M1 ;
        RECT 9.759 6.804 9.761 9.24 ;
  LAYER M1 ;
        RECT 9.839 6.804 9.841 9.24 ;
  LAYER M1 ;
        RECT 9.919 6.804 9.921 9.24 ;
  LAYER M1 ;
        RECT 9.999 6.804 10.001 9.24 ;
  LAYER M1 ;
        RECT 10.079 6.804 10.081 9.24 ;
  LAYER M1 ;
        RECT 10.159 6.804 10.161 9.24 ;
  LAYER M1 ;
        RECT 10.239 6.804 10.241 9.24 ;
  LAYER M1 ;
        RECT 10.319 6.804 10.321 9.24 ;
  LAYER M1 ;
        RECT 10.399 6.804 10.401 9.24 ;
  LAYER M1 ;
        RECT 10.479 6.804 10.481 9.24 ;
  LAYER M1 ;
        RECT 10.559 6.804 10.561 9.24 ;
  LAYER M1 ;
        RECT 10.639 6.804 10.641 9.24 ;
  LAYER M1 ;
        RECT 10.719 6.804 10.721 9.24 ;
  LAYER M1 ;
        RECT 10.799 6.804 10.801 9.24 ;
  LAYER M1 ;
        RECT 10.879 6.804 10.881 9.24 ;
  LAYER M1 ;
        RECT 10.959 6.804 10.961 9.24 ;
  LAYER M1 ;
        RECT 11.039 6.804 11.041 9.24 ;
  LAYER M1 ;
        RECT 11.119 6.804 11.121 9.24 ;
  LAYER M1 ;
        RECT 11.199 6.804 11.201 9.24 ;
  LAYER M1 ;
        RECT 11.279 6.804 11.281 9.24 ;
  LAYER M1 ;
        RECT 11.359 6.804 11.361 9.24 ;
  LAYER M1 ;
        RECT 11.439 6.804 11.441 9.24 ;
  LAYER M1 ;
        RECT 11.519 6.804 11.521 9.24 ;
  LAYER M1 ;
        RECT 11.599 6.804 11.601 9.24 ;
  LAYER M1 ;
        RECT 11.679 6.804 11.681 9.24 ;
  LAYER M1 ;
        RECT 11.759 6.804 11.761 9.24 ;
  LAYER M1 ;
        RECT 11.839 6.804 11.841 9.24 ;
  LAYER M1 ;
        RECT 11.919 6.804 11.921 9.24 ;
  LAYER M1 ;
        RECT 11.999 6.804 12.001 9.24 ;
  LAYER M2 ;
        RECT 9.68 6.803 12.08 6.805 ;
  LAYER M2 ;
        RECT 9.68 6.887 12.08 6.889 ;
  LAYER M2 ;
        RECT 9.68 6.971 12.08 6.973 ;
  LAYER M2 ;
        RECT 9.68 7.055 12.08 7.057 ;
  LAYER M2 ;
        RECT 9.68 7.139 12.08 7.141 ;
  LAYER M2 ;
        RECT 9.68 7.223 12.08 7.225 ;
  LAYER M2 ;
        RECT 9.68 7.307 12.08 7.309 ;
  LAYER M2 ;
        RECT 9.68 7.391 12.08 7.393 ;
  LAYER M2 ;
        RECT 9.68 7.475 12.08 7.477 ;
  LAYER M2 ;
        RECT 9.68 7.559 12.08 7.561 ;
  LAYER M2 ;
        RECT 9.68 7.643 12.08 7.645 ;
  LAYER M2 ;
        RECT 9.68 7.727 12.08 7.729 ;
  LAYER M2 ;
        RECT 9.68 7.8105 12.08 7.8125 ;
  LAYER M2 ;
        RECT 9.68 7.895 12.08 7.897 ;
  LAYER M2 ;
        RECT 9.68 7.979 12.08 7.981 ;
  LAYER M2 ;
        RECT 9.68 8.063 12.08 8.065 ;
  LAYER M2 ;
        RECT 9.68 8.147 12.08 8.149 ;
  LAYER M2 ;
        RECT 9.68 8.231 12.08 8.233 ;
  LAYER M2 ;
        RECT 9.68 8.315 12.08 8.317 ;
  LAYER M2 ;
        RECT 9.68 8.399 12.08 8.401 ;
  LAYER M2 ;
        RECT 9.68 8.483 12.08 8.485 ;
  LAYER M2 ;
        RECT 9.68 8.567 12.08 8.569 ;
  LAYER M2 ;
        RECT 9.68 8.651 12.08 8.653 ;
  LAYER M2 ;
        RECT 9.68 8.735 12.08 8.737 ;
  LAYER M2 ;
        RECT 9.68 8.819 12.08 8.821 ;
  LAYER M2 ;
        RECT 9.68 8.903 12.08 8.905 ;
  LAYER M2 ;
        RECT 9.68 8.987 12.08 8.989 ;
  LAYER M2 ;
        RECT 9.68 9.071 12.08 9.073 ;
  LAYER M2 ;
        RECT 9.68 9.155 12.08 9.157 ;
  LAYER M1 ;
        RECT 9.664 9.708 9.696 12.216 ;
  LAYER M1 ;
        RECT 9.728 9.708 9.76 12.216 ;
  LAYER M1 ;
        RECT 9.792 9.708 9.824 12.216 ;
  LAYER M1 ;
        RECT 9.856 9.708 9.888 12.216 ;
  LAYER M1 ;
        RECT 9.92 9.708 9.952 12.216 ;
  LAYER M1 ;
        RECT 9.984 9.708 10.016 12.216 ;
  LAYER M1 ;
        RECT 10.048 9.708 10.08 12.216 ;
  LAYER M1 ;
        RECT 10.112 9.708 10.144 12.216 ;
  LAYER M1 ;
        RECT 10.176 9.708 10.208 12.216 ;
  LAYER M1 ;
        RECT 10.24 9.708 10.272 12.216 ;
  LAYER M1 ;
        RECT 10.304 9.708 10.336 12.216 ;
  LAYER M1 ;
        RECT 10.368 9.708 10.4 12.216 ;
  LAYER M1 ;
        RECT 10.432 9.708 10.464 12.216 ;
  LAYER M1 ;
        RECT 10.496 9.708 10.528 12.216 ;
  LAYER M1 ;
        RECT 10.56 9.708 10.592 12.216 ;
  LAYER M1 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M1 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M1 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M1 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M1 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M1 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M1 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M1 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M1 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M1 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M1 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M1 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M1 ;
        RECT 11.392 9.708 11.424 12.216 ;
  LAYER M1 ;
        RECT 11.456 9.708 11.488 12.216 ;
  LAYER M1 ;
        RECT 11.52 9.708 11.552 12.216 ;
  LAYER M1 ;
        RECT 11.584 9.708 11.616 12.216 ;
  LAYER M1 ;
        RECT 11.648 9.708 11.68 12.216 ;
  LAYER M1 ;
        RECT 11.712 9.708 11.744 12.216 ;
  LAYER M1 ;
        RECT 11.776 9.708 11.808 12.216 ;
  LAYER M1 ;
        RECT 11.84 9.708 11.872 12.216 ;
  LAYER M1 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M1 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M2 ;
        RECT 9.644 9.792 12.116 9.824 ;
  LAYER M2 ;
        RECT 9.644 9.856 12.116 9.888 ;
  LAYER M2 ;
        RECT 9.644 9.92 12.116 9.952 ;
  LAYER M2 ;
        RECT 9.644 9.984 12.116 10.016 ;
  LAYER M2 ;
        RECT 9.644 10.048 12.116 10.08 ;
  LAYER M2 ;
        RECT 9.644 10.112 12.116 10.144 ;
  LAYER M2 ;
        RECT 9.644 10.176 12.116 10.208 ;
  LAYER M2 ;
        RECT 9.644 10.24 12.116 10.272 ;
  LAYER M2 ;
        RECT 9.644 10.304 12.116 10.336 ;
  LAYER M2 ;
        RECT 9.644 10.368 12.116 10.4 ;
  LAYER M2 ;
        RECT 9.644 10.432 12.116 10.464 ;
  LAYER M2 ;
        RECT 9.644 10.496 12.116 10.528 ;
  LAYER M2 ;
        RECT 9.644 10.56 12.116 10.592 ;
  LAYER M2 ;
        RECT 9.644 10.624 12.116 10.656 ;
  LAYER M2 ;
        RECT 9.644 10.688 12.116 10.72 ;
  LAYER M2 ;
        RECT 9.644 10.752 12.116 10.784 ;
  LAYER M2 ;
        RECT 9.644 10.816 12.116 10.848 ;
  LAYER M2 ;
        RECT 9.644 10.88 12.116 10.912 ;
  LAYER M2 ;
        RECT 9.644 10.944 12.116 10.976 ;
  LAYER M2 ;
        RECT 9.644 11.008 12.116 11.04 ;
  LAYER M2 ;
        RECT 9.644 11.072 12.116 11.104 ;
  LAYER M2 ;
        RECT 9.644 11.136 12.116 11.168 ;
  LAYER M2 ;
        RECT 9.644 11.2 12.116 11.232 ;
  LAYER M2 ;
        RECT 9.644 11.264 12.116 11.296 ;
  LAYER M2 ;
        RECT 9.644 11.328 12.116 11.36 ;
  LAYER M2 ;
        RECT 9.644 11.392 12.116 11.424 ;
  LAYER M2 ;
        RECT 9.644 11.456 12.116 11.488 ;
  LAYER M2 ;
        RECT 9.644 11.52 12.116 11.552 ;
  LAYER M2 ;
        RECT 9.644 11.584 12.116 11.616 ;
  LAYER M2 ;
        RECT 9.644 11.648 12.116 11.68 ;
  LAYER M2 ;
        RECT 9.644 11.712 12.116 11.744 ;
  LAYER M2 ;
        RECT 9.644 11.776 12.116 11.808 ;
  LAYER M2 ;
        RECT 9.644 11.84 12.116 11.872 ;
  LAYER M2 ;
        RECT 9.644 11.904 12.116 11.936 ;
  LAYER M2 ;
        RECT 9.644 11.968 12.116 12 ;
  LAYER M2 ;
        RECT 9.644 12.032 12.116 12.064 ;
  LAYER M3 ;
        RECT 9.664 9.708 9.696 12.216 ;
  LAYER M3 ;
        RECT 9.728 9.708 9.76 12.216 ;
  LAYER M3 ;
        RECT 9.792 9.708 9.824 12.216 ;
  LAYER M3 ;
        RECT 9.856 9.708 9.888 12.216 ;
  LAYER M3 ;
        RECT 9.92 9.708 9.952 12.216 ;
  LAYER M3 ;
        RECT 9.984 9.708 10.016 12.216 ;
  LAYER M3 ;
        RECT 10.048 9.708 10.08 12.216 ;
  LAYER M3 ;
        RECT 10.112 9.708 10.144 12.216 ;
  LAYER M3 ;
        RECT 10.176 9.708 10.208 12.216 ;
  LAYER M3 ;
        RECT 10.24 9.708 10.272 12.216 ;
  LAYER M3 ;
        RECT 10.304 9.708 10.336 12.216 ;
  LAYER M3 ;
        RECT 10.368 9.708 10.4 12.216 ;
  LAYER M3 ;
        RECT 10.432 9.708 10.464 12.216 ;
  LAYER M3 ;
        RECT 10.496 9.708 10.528 12.216 ;
  LAYER M3 ;
        RECT 10.56 9.708 10.592 12.216 ;
  LAYER M3 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M3 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M3 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M3 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M3 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M3 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M3 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M3 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M3 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M3 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M3 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M3 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M3 ;
        RECT 11.392 9.708 11.424 12.216 ;
  LAYER M3 ;
        RECT 11.456 9.708 11.488 12.216 ;
  LAYER M3 ;
        RECT 11.52 9.708 11.552 12.216 ;
  LAYER M3 ;
        RECT 11.584 9.708 11.616 12.216 ;
  LAYER M3 ;
        RECT 11.648 9.708 11.68 12.216 ;
  LAYER M3 ;
        RECT 11.712 9.708 11.744 12.216 ;
  LAYER M3 ;
        RECT 11.776 9.708 11.808 12.216 ;
  LAYER M3 ;
        RECT 11.84 9.708 11.872 12.216 ;
  LAYER M3 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M3 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M3 ;
        RECT 12.064 9.708 12.096 12.216 ;
  LAYER M1 ;
        RECT 9.679 9.744 9.681 12.18 ;
  LAYER M1 ;
        RECT 9.759 9.744 9.761 12.18 ;
  LAYER M1 ;
        RECT 9.839 9.744 9.841 12.18 ;
  LAYER M1 ;
        RECT 9.919 9.744 9.921 12.18 ;
  LAYER M1 ;
        RECT 9.999 9.744 10.001 12.18 ;
  LAYER M1 ;
        RECT 10.079 9.744 10.081 12.18 ;
  LAYER M1 ;
        RECT 10.159 9.744 10.161 12.18 ;
  LAYER M1 ;
        RECT 10.239 9.744 10.241 12.18 ;
  LAYER M1 ;
        RECT 10.319 9.744 10.321 12.18 ;
  LAYER M1 ;
        RECT 10.399 9.744 10.401 12.18 ;
  LAYER M1 ;
        RECT 10.479 9.744 10.481 12.18 ;
  LAYER M1 ;
        RECT 10.559 9.744 10.561 12.18 ;
  LAYER M1 ;
        RECT 10.639 9.744 10.641 12.18 ;
  LAYER M1 ;
        RECT 10.719 9.744 10.721 12.18 ;
  LAYER M1 ;
        RECT 10.799 9.744 10.801 12.18 ;
  LAYER M1 ;
        RECT 10.879 9.744 10.881 12.18 ;
  LAYER M1 ;
        RECT 10.959 9.744 10.961 12.18 ;
  LAYER M1 ;
        RECT 11.039 9.744 11.041 12.18 ;
  LAYER M1 ;
        RECT 11.119 9.744 11.121 12.18 ;
  LAYER M1 ;
        RECT 11.199 9.744 11.201 12.18 ;
  LAYER M1 ;
        RECT 11.279 9.744 11.281 12.18 ;
  LAYER M1 ;
        RECT 11.359 9.744 11.361 12.18 ;
  LAYER M1 ;
        RECT 11.439 9.744 11.441 12.18 ;
  LAYER M1 ;
        RECT 11.519 9.744 11.521 12.18 ;
  LAYER M1 ;
        RECT 11.599 9.744 11.601 12.18 ;
  LAYER M1 ;
        RECT 11.679 9.744 11.681 12.18 ;
  LAYER M1 ;
        RECT 11.759 9.744 11.761 12.18 ;
  LAYER M1 ;
        RECT 11.839 9.744 11.841 12.18 ;
  LAYER M1 ;
        RECT 11.919 9.744 11.921 12.18 ;
  LAYER M1 ;
        RECT 11.999 9.744 12.001 12.18 ;
  LAYER M2 ;
        RECT 9.68 9.743 12.08 9.745 ;
  LAYER M2 ;
        RECT 9.68 9.827 12.08 9.829 ;
  LAYER M2 ;
        RECT 9.68 9.911 12.08 9.913 ;
  LAYER M2 ;
        RECT 9.68 9.995 12.08 9.997 ;
  LAYER M2 ;
        RECT 9.68 10.079 12.08 10.081 ;
  LAYER M2 ;
        RECT 9.68 10.163 12.08 10.165 ;
  LAYER M2 ;
        RECT 9.68 10.247 12.08 10.249 ;
  LAYER M2 ;
        RECT 9.68 10.331 12.08 10.333 ;
  LAYER M2 ;
        RECT 9.68 10.415 12.08 10.417 ;
  LAYER M2 ;
        RECT 9.68 10.499 12.08 10.501 ;
  LAYER M2 ;
        RECT 9.68 10.583 12.08 10.585 ;
  LAYER M2 ;
        RECT 9.68 10.667 12.08 10.669 ;
  LAYER M2 ;
        RECT 9.68 10.7505 12.08 10.7525 ;
  LAYER M2 ;
        RECT 9.68 10.835 12.08 10.837 ;
  LAYER M2 ;
        RECT 9.68 10.919 12.08 10.921 ;
  LAYER M2 ;
        RECT 9.68 11.003 12.08 11.005 ;
  LAYER M2 ;
        RECT 9.68 11.087 12.08 11.089 ;
  LAYER M2 ;
        RECT 9.68 11.171 12.08 11.173 ;
  LAYER M2 ;
        RECT 9.68 11.255 12.08 11.257 ;
  LAYER M2 ;
        RECT 9.68 11.339 12.08 11.341 ;
  LAYER M2 ;
        RECT 9.68 11.423 12.08 11.425 ;
  LAYER M2 ;
        RECT 9.68 11.507 12.08 11.509 ;
  LAYER M2 ;
        RECT 9.68 11.591 12.08 11.593 ;
  LAYER M2 ;
        RECT 9.68 11.675 12.08 11.677 ;
  LAYER M2 ;
        RECT 9.68 11.759 12.08 11.761 ;
  LAYER M2 ;
        RECT 9.68 11.843 12.08 11.845 ;
  LAYER M2 ;
        RECT 9.68 11.927 12.08 11.929 ;
  LAYER M2 ;
        RECT 9.68 12.011 12.08 12.013 ;
  LAYER M2 ;
        RECT 9.68 12.095 12.08 12.097 ;
  LAYER M1 ;
        RECT 9.664 12.648 9.696 15.156 ;
  LAYER M1 ;
        RECT 9.728 12.648 9.76 15.156 ;
  LAYER M1 ;
        RECT 9.792 12.648 9.824 15.156 ;
  LAYER M1 ;
        RECT 9.856 12.648 9.888 15.156 ;
  LAYER M1 ;
        RECT 9.92 12.648 9.952 15.156 ;
  LAYER M1 ;
        RECT 9.984 12.648 10.016 15.156 ;
  LAYER M1 ;
        RECT 10.048 12.648 10.08 15.156 ;
  LAYER M1 ;
        RECT 10.112 12.648 10.144 15.156 ;
  LAYER M1 ;
        RECT 10.176 12.648 10.208 15.156 ;
  LAYER M1 ;
        RECT 10.24 12.648 10.272 15.156 ;
  LAYER M1 ;
        RECT 10.304 12.648 10.336 15.156 ;
  LAYER M1 ;
        RECT 10.368 12.648 10.4 15.156 ;
  LAYER M1 ;
        RECT 10.432 12.648 10.464 15.156 ;
  LAYER M1 ;
        RECT 10.496 12.648 10.528 15.156 ;
  LAYER M1 ;
        RECT 10.56 12.648 10.592 15.156 ;
  LAYER M1 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M1 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M1 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M1 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M1 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M1 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M1 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M1 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M1 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M1 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M1 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M1 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M1 ;
        RECT 11.392 12.648 11.424 15.156 ;
  LAYER M1 ;
        RECT 11.456 12.648 11.488 15.156 ;
  LAYER M1 ;
        RECT 11.52 12.648 11.552 15.156 ;
  LAYER M1 ;
        RECT 11.584 12.648 11.616 15.156 ;
  LAYER M1 ;
        RECT 11.648 12.648 11.68 15.156 ;
  LAYER M1 ;
        RECT 11.712 12.648 11.744 15.156 ;
  LAYER M1 ;
        RECT 11.776 12.648 11.808 15.156 ;
  LAYER M1 ;
        RECT 11.84 12.648 11.872 15.156 ;
  LAYER M1 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M1 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M2 ;
        RECT 9.644 12.732 12.116 12.764 ;
  LAYER M2 ;
        RECT 9.644 12.796 12.116 12.828 ;
  LAYER M2 ;
        RECT 9.644 12.86 12.116 12.892 ;
  LAYER M2 ;
        RECT 9.644 12.924 12.116 12.956 ;
  LAYER M2 ;
        RECT 9.644 12.988 12.116 13.02 ;
  LAYER M2 ;
        RECT 9.644 13.052 12.116 13.084 ;
  LAYER M2 ;
        RECT 9.644 13.116 12.116 13.148 ;
  LAYER M2 ;
        RECT 9.644 13.18 12.116 13.212 ;
  LAYER M2 ;
        RECT 9.644 13.244 12.116 13.276 ;
  LAYER M2 ;
        RECT 9.644 13.308 12.116 13.34 ;
  LAYER M2 ;
        RECT 9.644 13.372 12.116 13.404 ;
  LAYER M2 ;
        RECT 9.644 13.436 12.116 13.468 ;
  LAYER M2 ;
        RECT 9.644 13.5 12.116 13.532 ;
  LAYER M2 ;
        RECT 9.644 13.564 12.116 13.596 ;
  LAYER M2 ;
        RECT 9.644 13.628 12.116 13.66 ;
  LAYER M2 ;
        RECT 9.644 13.692 12.116 13.724 ;
  LAYER M2 ;
        RECT 9.644 13.756 12.116 13.788 ;
  LAYER M2 ;
        RECT 9.644 13.82 12.116 13.852 ;
  LAYER M2 ;
        RECT 9.644 13.884 12.116 13.916 ;
  LAYER M2 ;
        RECT 9.644 13.948 12.116 13.98 ;
  LAYER M2 ;
        RECT 9.644 14.012 12.116 14.044 ;
  LAYER M2 ;
        RECT 9.644 14.076 12.116 14.108 ;
  LAYER M2 ;
        RECT 9.644 14.14 12.116 14.172 ;
  LAYER M2 ;
        RECT 9.644 14.204 12.116 14.236 ;
  LAYER M2 ;
        RECT 9.644 14.268 12.116 14.3 ;
  LAYER M2 ;
        RECT 9.644 14.332 12.116 14.364 ;
  LAYER M2 ;
        RECT 9.644 14.396 12.116 14.428 ;
  LAYER M2 ;
        RECT 9.644 14.46 12.116 14.492 ;
  LAYER M2 ;
        RECT 9.644 14.524 12.116 14.556 ;
  LAYER M2 ;
        RECT 9.644 14.588 12.116 14.62 ;
  LAYER M2 ;
        RECT 9.644 14.652 12.116 14.684 ;
  LAYER M2 ;
        RECT 9.644 14.716 12.116 14.748 ;
  LAYER M2 ;
        RECT 9.644 14.78 12.116 14.812 ;
  LAYER M2 ;
        RECT 9.644 14.844 12.116 14.876 ;
  LAYER M2 ;
        RECT 9.644 14.908 12.116 14.94 ;
  LAYER M2 ;
        RECT 9.644 14.972 12.116 15.004 ;
  LAYER M3 ;
        RECT 9.664 12.648 9.696 15.156 ;
  LAYER M3 ;
        RECT 9.728 12.648 9.76 15.156 ;
  LAYER M3 ;
        RECT 9.792 12.648 9.824 15.156 ;
  LAYER M3 ;
        RECT 9.856 12.648 9.888 15.156 ;
  LAYER M3 ;
        RECT 9.92 12.648 9.952 15.156 ;
  LAYER M3 ;
        RECT 9.984 12.648 10.016 15.156 ;
  LAYER M3 ;
        RECT 10.048 12.648 10.08 15.156 ;
  LAYER M3 ;
        RECT 10.112 12.648 10.144 15.156 ;
  LAYER M3 ;
        RECT 10.176 12.648 10.208 15.156 ;
  LAYER M3 ;
        RECT 10.24 12.648 10.272 15.156 ;
  LAYER M3 ;
        RECT 10.304 12.648 10.336 15.156 ;
  LAYER M3 ;
        RECT 10.368 12.648 10.4 15.156 ;
  LAYER M3 ;
        RECT 10.432 12.648 10.464 15.156 ;
  LAYER M3 ;
        RECT 10.496 12.648 10.528 15.156 ;
  LAYER M3 ;
        RECT 10.56 12.648 10.592 15.156 ;
  LAYER M3 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M3 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M3 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M3 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M3 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M3 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M3 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M3 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M3 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M3 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M3 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M3 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M3 ;
        RECT 11.392 12.648 11.424 15.156 ;
  LAYER M3 ;
        RECT 11.456 12.648 11.488 15.156 ;
  LAYER M3 ;
        RECT 11.52 12.648 11.552 15.156 ;
  LAYER M3 ;
        RECT 11.584 12.648 11.616 15.156 ;
  LAYER M3 ;
        RECT 11.648 12.648 11.68 15.156 ;
  LAYER M3 ;
        RECT 11.712 12.648 11.744 15.156 ;
  LAYER M3 ;
        RECT 11.776 12.648 11.808 15.156 ;
  LAYER M3 ;
        RECT 11.84 12.648 11.872 15.156 ;
  LAYER M3 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M3 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M3 ;
        RECT 12.064 12.648 12.096 15.156 ;
  LAYER M1 ;
        RECT 9.679 12.684 9.681 15.12 ;
  LAYER M1 ;
        RECT 9.759 12.684 9.761 15.12 ;
  LAYER M1 ;
        RECT 9.839 12.684 9.841 15.12 ;
  LAYER M1 ;
        RECT 9.919 12.684 9.921 15.12 ;
  LAYER M1 ;
        RECT 9.999 12.684 10.001 15.12 ;
  LAYER M1 ;
        RECT 10.079 12.684 10.081 15.12 ;
  LAYER M1 ;
        RECT 10.159 12.684 10.161 15.12 ;
  LAYER M1 ;
        RECT 10.239 12.684 10.241 15.12 ;
  LAYER M1 ;
        RECT 10.319 12.684 10.321 15.12 ;
  LAYER M1 ;
        RECT 10.399 12.684 10.401 15.12 ;
  LAYER M1 ;
        RECT 10.479 12.684 10.481 15.12 ;
  LAYER M1 ;
        RECT 10.559 12.684 10.561 15.12 ;
  LAYER M1 ;
        RECT 10.639 12.684 10.641 15.12 ;
  LAYER M1 ;
        RECT 10.719 12.684 10.721 15.12 ;
  LAYER M1 ;
        RECT 10.799 12.684 10.801 15.12 ;
  LAYER M1 ;
        RECT 10.879 12.684 10.881 15.12 ;
  LAYER M1 ;
        RECT 10.959 12.684 10.961 15.12 ;
  LAYER M1 ;
        RECT 11.039 12.684 11.041 15.12 ;
  LAYER M1 ;
        RECT 11.119 12.684 11.121 15.12 ;
  LAYER M1 ;
        RECT 11.199 12.684 11.201 15.12 ;
  LAYER M1 ;
        RECT 11.279 12.684 11.281 15.12 ;
  LAYER M1 ;
        RECT 11.359 12.684 11.361 15.12 ;
  LAYER M1 ;
        RECT 11.439 12.684 11.441 15.12 ;
  LAYER M1 ;
        RECT 11.519 12.684 11.521 15.12 ;
  LAYER M1 ;
        RECT 11.599 12.684 11.601 15.12 ;
  LAYER M1 ;
        RECT 11.679 12.684 11.681 15.12 ;
  LAYER M1 ;
        RECT 11.759 12.684 11.761 15.12 ;
  LAYER M1 ;
        RECT 11.839 12.684 11.841 15.12 ;
  LAYER M1 ;
        RECT 11.919 12.684 11.921 15.12 ;
  LAYER M1 ;
        RECT 11.999 12.684 12.001 15.12 ;
  LAYER M2 ;
        RECT 9.68 12.683 12.08 12.685 ;
  LAYER M2 ;
        RECT 9.68 12.767 12.08 12.769 ;
  LAYER M2 ;
        RECT 9.68 12.851 12.08 12.853 ;
  LAYER M2 ;
        RECT 9.68 12.935 12.08 12.937 ;
  LAYER M2 ;
        RECT 9.68 13.019 12.08 13.021 ;
  LAYER M2 ;
        RECT 9.68 13.103 12.08 13.105 ;
  LAYER M2 ;
        RECT 9.68 13.187 12.08 13.189 ;
  LAYER M2 ;
        RECT 9.68 13.271 12.08 13.273 ;
  LAYER M2 ;
        RECT 9.68 13.355 12.08 13.357 ;
  LAYER M2 ;
        RECT 9.68 13.439 12.08 13.441 ;
  LAYER M2 ;
        RECT 9.68 13.523 12.08 13.525 ;
  LAYER M2 ;
        RECT 9.68 13.607 12.08 13.609 ;
  LAYER M2 ;
        RECT 9.68 13.6905 12.08 13.6925 ;
  LAYER M2 ;
        RECT 9.68 13.775 12.08 13.777 ;
  LAYER M2 ;
        RECT 9.68 13.859 12.08 13.861 ;
  LAYER M2 ;
        RECT 9.68 13.943 12.08 13.945 ;
  LAYER M2 ;
        RECT 9.68 14.027 12.08 14.029 ;
  LAYER M2 ;
        RECT 9.68 14.111 12.08 14.113 ;
  LAYER M2 ;
        RECT 9.68 14.195 12.08 14.197 ;
  LAYER M2 ;
        RECT 9.68 14.279 12.08 14.281 ;
  LAYER M2 ;
        RECT 9.68 14.363 12.08 14.365 ;
  LAYER M2 ;
        RECT 9.68 14.447 12.08 14.449 ;
  LAYER M2 ;
        RECT 9.68 14.531 12.08 14.533 ;
  LAYER M2 ;
        RECT 9.68 14.615 12.08 14.617 ;
  LAYER M2 ;
        RECT 9.68 14.699 12.08 14.701 ;
  LAYER M2 ;
        RECT 9.68 14.783 12.08 14.785 ;
  LAYER M2 ;
        RECT 9.68 14.867 12.08 14.869 ;
  LAYER M2 ;
        RECT 9.68 14.951 12.08 14.953 ;
  LAYER M2 ;
        RECT 9.68 15.035 12.08 15.037 ;
  LAYER M1 ;
        RECT 9.664 15.588 9.696 18.096 ;
  LAYER M1 ;
        RECT 9.728 15.588 9.76 18.096 ;
  LAYER M1 ;
        RECT 9.792 15.588 9.824 18.096 ;
  LAYER M1 ;
        RECT 9.856 15.588 9.888 18.096 ;
  LAYER M1 ;
        RECT 9.92 15.588 9.952 18.096 ;
  LAYER M1 ;
        RECT 9.984 15.588 10.016 18.096 ;
  LAYER M1 ;
        RECT 10.048 15.588 10.08 18.096 ;
  LAYER M1 ;
        RECT 10.112 15.588 10.144 18.096 ;
  LAYER M1 ;
        RECT 10.176 15.588 10.208 18.096 ;
  LAYER M1 ;
        RECT 10.24 15.588 10.272 18.096 ;
  LAYER M1 ;
        RECT 10.304 15.588 10.336 18.096 ;
  LAYER M1 ;
        RECT 10.368 15.588 10.4 18.096 ;
  LAYER M1 ;
        RECT 10.432 15.588 10.464 18.096 ;
  LAYER M1 ;
        RECT 10.496 15.588 10.528 18.096 ;
  LAYER M1 ;
        RECT 10.56 15.588 10.592 18.096 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M1 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M1 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M1 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M1 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M1 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M1 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M1 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M1 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M1 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M1 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M1 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M1 ;
        RECT 11.392 15.588 11.424 18.096 ;
  LAYER M1 ;
        RECT 11.456 15.588 11.488 18.096 ;
  LAYER M1 ;
        RECT 11.52 15.588 11.552 18.096 ;
  LAYER M1 ;
        RECT 11.584 15.588 11.616 18.096 ;
  LAYER M1 ;
        RECT 11.648 15.588 11.68 18.096 ;
  LAYER M1 ;
        RECT 11.712 15.588 11.744 18.096 ;
  LAYER M1 ;
        RECT 11.776 15.588 11.808 18.096 ;
  LAYER M1 ;
        RECT 11.84 15.588 11.872 18.096 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M1 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M2 ;
        RECT 9.644 15.672 12.116 15.704 ;
  LAYER M2 ;
        RECT 9.644 15.736 12.116 15.768 ;
  LAYER M2 ;
        RECT 9.644 15.8 12.116 15.832 ;
  LAYER M2 ;
        RECT 9.644 15.864 12.116 15.896 ;
  LAYER M2 ;
        RECT 9.644 15.928 12.116 15.96 ;
  LAYER M2 ;
        RECT 9.644 15.992 12.116 16.024 ;
  LAYER M2 ;
        RECT 9.644 16.056 12.116 16.088 ;
  LAYER M2 ;
        RECT 9.644 16.12 12.116 16.152 ;
  LAYER M2 ;
        RECT 9.644 16.184 12.116 16.216 ;
  LAYER M2 ;
        RECT 9.644 16.248 12.116 16.28 ;
  LAYER M2 ;
        RECT 9.644 16.312 12.116 16.344 ;
  LAYER M2 ;
        RECT 9.644 16.376 12.116 16.408 ;
  LAYER M2 ;
        RECT 9.644 16.44 12.116 16.472 ;
  LAYER M2 ;
        RECT 9.644 16.504 12.116 16.536 ;
  LAYER M2 ;
        RECT 9.644 16.568 12.116 16.6 ;
  LAYER M2 ;
        RECT 9.644 16.632 12.116 16.664 ;
  LAYER M2 ;
        RECT 9.644 16.696 12.116 16.728 ;
  LAYER M2 ;
        RECT 9.644 16.76 12.116 16.792 ;
  LAYER M2 ;
        RECT 9.644 16.824 12.116 16.856 ;
  LAYER M2 ;
        RECT 9.644 16.888 12.116 16.92 ;
  LAYER M2 ;
        RECT 9.644 16.952 12.116 16.984 ;
  LAYER M2 ;
        RECT 9.644 17.016 12.116 17.048 ;
  LAYER M2 ;
        RECT 9.644 17.08 12.116 17.112 ;
  LAYER M2 ;
        RECT 9.644 17.144 12.116 17.176 ;
  LAYER M2 ;
        RECT 9.644 17.208 12.116 17.24 ;
  LAYER M2 ;
        RECT 9.644 17.272 12.116 17.304 ;
  LAYER M2 ;
        RECT 9.644 17.336 12.116 17.368 ;
  LAYER M2 ;
        RECT 9.644 17.4 12.116 17.432 ;
  LAYER M2 ;
        RECT 9.644 17.464 12.116 17.496 ;
  LAYER M2 ;
        RECT 9.644 17.528 12.116 17.56 ;
  LAYER M2 ;
        RECT 9.644 17.592 12.116 17.624 ;
  LAYER M2 ;
        RECT 9.644 17.656 12.116 17.688 ;
  LAYER M2 ;
        RECT 9.644 17.72 12.116 17.752 ;
  LAYER M2 ;
        RECT 9.644 17.784 12.116 17.816 ;
  LAYER M2 ;
        RECT 9.644 17.848 12.116 17.88 ;
  LAYER M2 ;
        RECT 9.644 17.912 12.116 17.944 ;
  LAYER M3 ;
        RECT 9.664 15.588 9.696 18.096 ;
  LAYER M3 ;
        RECT 9.728 15.588 9.76 18.096 ;
  LAYER M3 ;
        RECT 9.792 15.588 9.824 18.096 ;
  LAYER M3 ;
        RECT 9.856 15.588 9.888 18.096 ;
  LAYER M3 ;
        RECT 9.92 15.588 9.952 18.096 ;
  LAYER M3 ;
        RECT 9.984 15.588 10.016 18.096 ;
  LAYER M3 ;
        RECT 10.048 15.588 10.08 18.096 ;
  LAYER M3 ;
        RECT 10.112 15.588 10.144 18.096 ;
  LAYER M3 ;
        RECT 10.176 15.588 10.208 18.096 ;
  LAYER M3 ;
        RECT 10.24 15.588 10.272 18.096 ;
  LAYER M3 ;
        RECT 10.304 15.588 10.336 18.096 ;
  LAYER M3 ;
        RECT 10.368 15.588 10.4 18.096 ;
  LAYER M3 ;
        RECT 10.432 15.588 10.464 18.096 ;
  LAYER M3 ;
        RECT 10.496 15.588 10.528 18.096 ;
  LAYER M3 ;
        RECT 10.56 15.588 10.592 18.096 ;
  LAYER M3 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M3 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M3 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M3 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M3 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M3 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M3 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M3 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M3 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M3 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M3 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M3 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M3 ;
        RECT 11.392 15.588 11.424 18.096 ;
  LAYER M3 ;
        RECT 11.456 15.588 11.488 18.096 ;
  LAYER M3 ;
        RECT 11.52 15.588 11.552 18.096 ;
  LAYER M3 ;
        RECT 11.584 15.588 11.616 18.096 ;
  LAYER M3 ;
        RECT 11.648 15.588 11.68 18.096 ;
  LAYER M3 ;
        RECT 11.712 15.588 11.744 18.096 ;
  LAYER M3 ;
        RECT 11.776 15.588 11.808 18.096 ;
  LAYER M3 ;
        RECT 11.84 15.588 11.872 18.096 ;
  LAYER M3 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M3 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M3 ;
        RECT 12.064 15.588 12.096 18.096 ;
  LAYER M1 ;
        RECT 9.679 15.624 9.681 18.06 ;
  LAYER M1 ;
        RECT 9.759 15.624 9.761 18.06 ;
  LAYER M1 ;
        RECT 9.839 15.624 9.841 18.06 ;
  LAYER M1 ;
        RECT 9.919 15.624 9.921 18.06 ;
  LAYER M1 ;
        RECT 9.999 15.624 10.001 18.06 ;
  LAYER M1 ;
        RECT 10.079 15.624 10.081 18.06 ;
  LAYER M1 ;
        RECT 10.159 15.624 10.161 18.06 ;
  LAYER M1 ;
        RECT 10.239 15.624 10.241 18.06 ;
  LAYER M1 ;
        RECT 10.319 15.624 10.321 18.06 ;
  LAYER M1 ;
        RECT 10.399 15.624 10.401 18.06 ;
  LAYER M1 ;
        RECT 10.479 15.624 10.481 18.06 ;
  LAYER M1 ;
        RECT 10.559 15.624 10.561 18.06 ;
  LAYER M1 ;
        RECT 10.639 15.624 10.641 18.06 ;
  LAYER M1 ;
        RECT 10.719 15.624 10.721 18.06 ;
  LAYER M1 ;
        RECT 10.799 15.624 10.801 18.06 ;
  LAYER M1 ;
        RECT 10.879 15.624 10.881 18.06 ;
  LAYER M1 ;
        RECT 10.959 15.624 10.961 18.06 ;
  LAYER M1 ;
        RECT 11.039 15.624 11.041 18.06 ;
  LAYER M1 ;
        RECT 11.119 15.624 11.121 18.06 ;
  LAYER M1 ;
        RECT 11.199 15.624 11.201 18.06 ;
  LAYER M1 ;
        RECT 11.279 15.624 11.281 18.06 ;
  LAYER M1 ;
        RECT 11.359 15.624 11.361 18.06 ;
  LAYER M1 ;
        RECT 11.439 15.624 11.441 18.06 ;
  LAYER M1 ;
        RECT 11.519 15.624 11.521 18.06 ;
  LAYER M1 ;
        RECT 11.599 15.624 11.601 18.06 ;
  LAYER M1 ;
        RECT 11.679 15.624 11.681 18.06 ;
  LAYER M1 ;
        RECT 11.759 15.624 11.761 18.06 ;
  LAYER M1 ;
        RECT 11.839 15.624 11.841 18.06 ;
  LAYER M1 ;
        RECT 11.919 15.624 11.921 18.06 ;
  LAYER M1 ;
        RECT 11.999 15.624 12.001 18.06 ;
  LAYER M2 ;
        RECT 9.68 15.623 12.08 15.625 ;
  LAYER M2 ;
        RECT 9.68 15.707 12.08 15.709 ;
  LAYER M2 ;
        RECT 9.68 15.791 12.08 15.793 ;
  LAYER M2 ;
        RECT 9.68 15.875 12.08 15.877 ;
  LAYER M2 ;
        RECT 9.68 15.959 12.08 15.961 ;
  LAYER M2 ;
        RECT 9.68 16.043 12.08 16.045 ;
  LAYER M2 ;
        RECT 9.68 16.127 12.08 16.129 ;
  LAYER M2 ;
        RECT 9.68 16.211 12.08 16.213 ;
  LAYER M2 ;
        RECT 9.68 16.295 12.08 16.297 ;
  LAYER M2 ;
        RECT 9.68 16.379 12.08 16.381 ;
  LAYER M2 ;
        RECT 9.68 16.463 12.08 16.465 ;
  LAYER M2 ;
        RECT 9.68 16.547 12.08 16.549 ;
  LAYER M2 ;
        RECT 9.68 16.6305 12.08 16.6325 ;
  LAYER M2 ;
        RECT 9.68 16.715 12.08 16.717 ;
  LAYER M2 ;
        RECT 9.68 16.799 12.08 16.801 ;
  LAYER M2 ;
        RECT 9.68 16.883 12.08 16.885 ;
  LAYER M2 ;
        RECT 9.68 16.967 12.08 16.969 ;
  LAYER M2 ;
        RECT 9.68 17.051 12.08 17.053 ;
  LAYER M2 ;
        RECT 9.68 17.135 12.08 17.137 ;
  LAYER M2 ;
        RECT 9.68 17.219 12.08 17.221 ;
  LAYER M2 ;
        RECT 9.68 17.303 12.08 17.305 ;
  LAYER M2 ;
        RECT 9.68 17.387 12.08 17.389 ;
  LAYER M2 ;
        RECT 9.68 17.471 12.08 17.473 ;
  LAYER M2 ;
        RECT 9.68 17.555 12.08 17.557 ;
  LAYER M2 ;
        RECT 9.68 17.639 12.08 17.641 ;
  LAYER M2 ;
        RECT 9.68 17.723 12.08 17.725 ;
  LAYER M2 ;
        RECT 9.68 17.807 12.08 17.809 ;
  LAYER M2 ;
        RECT 9.68 17.891 12.08 17.893 ;
  LAYER M2 ;
        RECT 9.68 17.975 12.08 17.977 ;
  LAYER M1 ;
        RECT 9.664 18.528 9.696 21.036 ;
  LAYER M1 ;
        RECT 9.728 18.528 9.76 21.036 ;
  LAYER M1 ;
        RECT 9.792 18.528 9.824 21.036 ;
  LAYER M1 ;
        RECT 9.856 18.528 9.888 21.036 ;
  LAYER M1 ;
        RECT 9.92 18.528 9.952 21.036 ;
  LAYER M1 ;
        RECT 9.984 18.528 10.016 21.036 ;
  LAYER M1 ;
        RECT 10.048 18.528 10.08 21.036 ;
  LAYER M1 ;
        RECT 10.112 18.528 10.144 21.036 ;
  LAYER M1 ;
        RECT 10.176 18.528 10.208 21.036 ;
  LAYER M1 ;
        RECT 10.24 18.528 10.272 21.036 ;
  LAYER M1 ;
        RECT 10.304 18.528 10.336 21.036 ;
  LAYER M1 ;
        RECT 10.368 18.528 10.4 21.036 ;
  LAYER M1 ;
        RECT 10.432 18.528 10.464 21.036 ;
  LAYER M1 ;
        RECT 10.496 18.528 10.528 21.036 ;
  LAYER M1 ;
        RECT 10.56 18.528 10.592 21.036 ;
  LAYER M1 ;
        RECT 10.624 18.528 10.656 21.036 ;
  LAYER M1 ;
        RECT 10.688 18.528 10.72 21.036 ;
  LAYER M1 ;
        RECT 10.752 18.528 10.784 21.036 ;
  LAYER M1 ;
        RECT 10.816 18.528 10.848 21.036 ;
  LAYER M1 ;
        RECT 10.88 18.528 10.912 21.036 ;
  LAYER M1 ;
        RECT 10.944 18.528 10.976 21.036 ;
  LAYER M1 ;
        RECT 11.008 18.528 11.04 21.036 ;
  LAYER M1 ;
        RECT 11.072 18.528 11.104 21.036 ;
  LAYER M1 ;
        RECT 11.136 18.528 11.168 21.036 ;
  LAYER M1 ;
        RECT 11.2 18.528 11.232 21.036 ;
  LAYER M1 ;
        RECT 11.264 18.528 11.296 21.036 ;
  LAYER M1 ;
        RECT 11.328 18.528 11.36 21.036 ;
  LAYER M1 ;
        RECT 11.392 18.528 11.424 21.036 ;
  LAYER M1 ;
        RECT 11.456 18.528 11.488 21.036 ;
  LAYER M1 ;
        RECT 11.52 18.528 11.552 21.036 ;
  LAYER M1 ;
        RECT 11.584 18.528 11.616 21.036 ;
  LAYER M1 ;
        RECT 11.648 18.528 11.68 21.036 ;
  LAYER M1 ;
        RECT 11.712 18.528 11.744 21.036 ;
  LAYER M1 ;
        RECT 11.776 18.528 11.808 21.036 ;
  LAYER M1 ;
        RECT 11.84 18.528 11.872 21.036 ;
  LAYER M1 ;
        RECT 11.904 18.528 11.936 21.036 ;
  LAYER M1 ;
        RECT 11.968 18.528 12 21.036 ;
  LAYER M2 ;
        RECT 9.644 18.612 12.116 18.644 ;
  LAYER M2 ;
        RECT 9.644 18.676 12.116 18.708 ;
  LAYER M2 ;
        RECT 9.644 18.74 12.116 18.772 ;
  LAYER M2 ;
        RECT 9.644 18.804 12.116 18.836 ;
  LAYER M2 ;
        RECT 9.644 18.868 12.116 18.9 ;
  LAYER M2 ;
        RECT 9.644 18.932 12.116 18.964 ;
  LAYER M2 ;
        RECT 9.644 18.996 12.116 19.028 ;
  LAYER M2 ;
        RECT 9.644 19.06 12.116 19.092 ;
  LAYER M2 ;
        RECT 9.644 19.124 12.116 19.156 ;
  LAYER M2 ;
        RECT 9.644 19.188 12.116 19.22 ;
  LAYER M2 ;
        RECT 9.644 19.252 12.116 19.284 ;
  LAYER M2 ;
        RECT 9.644 19.316 12.116 19.348 ;
  LAYER M2 ;
        RECT 9.644 19.38 12.116 19.412 ;
  LAYER M2 ;
        RECT 9.644 19.444 12.116 19.476 ;
  LAYER M2 ;
        RECT 9.644 19.508 12.116 19.54 ;
  LAYER M2 ;
        RECT 9.644 19.572 12.116 19.604 ;
  LAYER M2 ;
        RECT 9.644 19.636 12.116 19.668 ;
  LAYER M2 ;
        RECT 9.644 19.7 12.116 19.732 ;
  LAYER M2 ;
        RECT 9.644 19.764 12.116 19.796 ;
  LAYER M2 ;
        RECT 9.644 19.828 12.116 19.86 ;
  LAYER M2 ;
        RECT 9.644 19.892 12.116 19.924 ;
  LAYER M2 ;
        RECT 9.644 19.956 12.116 19.988 ;
  LAYER M2 ;
        RECT 9.644 20.02 12.116 20.052 ;
  LAYER M2 ;
        RECT 9.644 20.084 12.116 20.116 ;
  LAYER M2 ;
        RECT 9.644 20.148 12.116 20.18 ;
  LAYER M2 ;
        RECT 9.644 20.212 12.116 20.244 ;
  LAYER M2 ;
        RECT 9.644 20.276 12.116 20.308 ;
  LAYER M2 ;
        RECT 9.644 20.34 12.116 20.372 ;
  LAYER M2 ;
        RECT 9.644 20.404 12.116 20.436 ;
  LAYER M2 ;
        RECT 9.644 20.468 12.116 20.5 ;
  LAYER M2 ;
        RECT 9.644 20.532 12.116 20.564 ;
  LAYER M2 ;
        RECT 9.644 20.596 12.116 20.628 ;
  LAYER M2 ;
        RECT 9.644 20.66 12.116 20.692 ;
  LAYER M2 ;
        RECT 9.644 20.724 12.116 20.756 ;
  LAYER M2 ;
        RECT 9.644 20.788 12.116 20.82 ;
  LAYER M2 ;
        RECT 9.644 20.852 12.116 20.884 ;
  LAYER M3 ;
        RECT 9.664 18.528 9.696 21.036 ;
  LAYER M3 ;
        RECT 9.728 18.528 9.76 21.036 ;
  LAYER M3 ;
        RECT 9.792 18.528 9.824 21.036 ;
  LAYER M3 ;
        RECT 9.856 18.528 9.888 21.036 ;
  LAYER M3 ;
        RECT 9.92 18.528 9.952 21.036 ;
  LAYER M3 ;
        RECT 9.984 18.528 10.016 21.036 ;
  LAYER M3 ;
        RECT 10.048 18.528 10.08 21.036 ;
  LAYER M3 ;
        RECT 10.112 18.528 10.144 21.036 ;
  LAYER M3 ;
        RECT 10.176 18.528 10.208 21.036 ;
  LAYER M3 ;
        RECT 10.24 18.528 10.272 21.036 ;
  LAYER M3 ;
        RECT 10.304 18.528 10.336 21.036 ;
  LAYER M3 ;
        RECT 10.368 18.528 10.4 21.036 ;
  LAYER M3 ;
        RECT 10.432 18.528 10.464 21.036 ;
  LAYER M3 ;
        RECT 10.496 18.528 10.528 21.036 ;
  LAYER M3 ;
        RECT 10.56 18.528 10.592 21.036 ;
  LAYER M3 ;
        RECT 10.624 18.528 10.656 21.036 ;
  LAYER M3 ;
        RECT 10.688 18.528 10.72 21.036 ;
  LAYER M3 ;
        RECT 10.752 18.528 10.784 21.036 ;
  LAYER M3 ;
        RECT 10.816 18.528 10.848 21.036 ;
  LAYER M3 ;
        RECT 10.88 18.528 10.912 21.036 ;
  LAYER M3 ;
        RECT 10.944 18.528 10.976 21.036 ;
  LAYER M3 ;
        RECT 11.008 18.528 11.04 21.036 ;
  LAYER M3 ;
        RECT 11.072 18.528 11.104 21.036 ;
  LAYER M3 ;
        RECT 11.136 18.528 11.168 21.036 ;
  LAYER M3 ;
        RECT 11.2 18.528 11.232 21.036 ;
  LAYER M3 ;
        RECT 11.264 18.528 11.296 21.036 ;
  LAYER M3 ;
        RECT 11.328 18.528 11.36 21.036 ;
  LAYER M3 ;
        RECT 11.392 18.528 11.424 21.036 ;
  LAYER M3 ;
        RECT 11.456 18.528 11.488 21.036 ;
  LAYER M3 ;
        RECT 11.52 18.528 11.552 21.036 ;
  LAYER M3 ;
        RECT 11.584 18.528 11.616 21.036 ;
  LAYER M3 ;
        RECT 11.648 18.528 11.68 21.036 ;
  LAYER M3 ;
        RECT 11.712 18.528 11.744 21.036 ;
  LAYER M3 ;
        RECT 11.776 18.528 11.808 21.036 ;
  LAYER M3 ;
        RECT 11.84 18.528 11.872 21.036 ;
  LAYER M3 ;
        RECT 11.904 18.528 11.936 21.036 ;
  LAYER M3 ;
        RECT 11.968 18.528 12 21.036 ;
  LAYER M3 ;
        RECT 12.064 18.528 12.096 21.036 ;
  LAYER M1 ;
        RECT 9.679 18.564 9.681 21 ;
  LAYER M1 ;
        RECT 9.759 18.564 9.761 21 ;
  LAYER M1 ;
        RECT 9.839 18.564 9.841 21 ;
  LAYER M1 ;
        RECT 9.919 18.564 9.921 21 ;
  LAYER M1 ;
        RECT 9.999 18.564 10.001 21 ;
  LAYER M1 ;
        RECT 10.079 18.564 10.081 21 ;
  LAYER M1 ;
        RECT 10.159 18.564 10.161 21 ;
  LAYER M1 ;
        RECT 10.239 18.564 10.241 21 ;
  LAYER M1 ;
        RECT 10.319 18.564 10.321 21 ;
  LAYER M1 ;
        RECT 10.399 18.564 10.401 21 ;
  LAYER M1 ;
        RECT 10.479 18.564 10.481 21 ;
  LAYER M1 ;
        RECT 10.559 18.564 10.561 21 ;
  LAYER M1 ;
        RECT 10.639 18.564 10.641 21 ;
  LAYER M1 ;
        RECT 10.719 18.564 10.721 21 ;
  LAYER M1 ;
        RECT 10.799 18.564 10.801 21 ;
  LAYER M1 ;
        RECT 10.879 18.564 10.881 21 ;
  LAYER M1 ;
        RECT 10.959 18.564 10.961 21 ;
  LAYER M1 ;
        RECT 11.039 18.564 11.041 21 ;
  LAYER M1 ;
        RECT 11.119 18.564 11.121 21 ;
  LAYER M1 ;
        RECT 11.199 18.564 11.201 21 ;
  LAYER M1 ;
        RECT 11.279 18.564 11.281 21 ;
  LAYER M1 ;
        RECT 11.359 18.564 11.361 21 ;
  LAYER M1 ;
        RECT 11.439 18.564 11.441 21 ;
  LAYER M1 ;
        RECT 11.519 18.564 11.521 21 ;
  LAYER M1 ;
        RECT 11.599 18.564 11.601 21 ;
  LAYER M1 ;
        RECT 11.679 18.564 11.681 21 ;
  LAYER M1 ;
        RECT 11.759 18.564 11.761 21 ;
  LAYER M1 ;
        RECT 11.839 18.564 11.841 21 ;
  LAYER M1 ;
        RECT 11.919 18.564 11.921 21 ;
  LAYER M1 ;
        RECT 11.999 18.564 12.001 21 ;
  LAYER M2 ;
        RECT 9.68 18.563 12.08 18.565 ;
  LAYER M2 ;
        RECT 9.68 18.647 12.08 18.649 ;
  LAYER M2 ;
        RECT 9.68 18.731 12.08 18.733 ;
  LAYER M2 ;
        RECT 9.68 18.815 12.08 18.817 ;
  LAYER M2 ;
        RECT 9.68 18.899 12.08 18.901 ;
  LAYER M2 ;
        RECT 9.68 18.983 12.08 18.985 ;
  LAYER M2 ;
        RECT 9.68 19.067 12.08 19.069 ;
  LAYER M2 ;
        RECT 9.68 19.151 12.08 19.153 ;
  LAYER M2 ;
        RECT 9.68 19.235 12.08 19.237 ;
  LAYER M2 ;
        RECT 9.68 19.319 12.08 19.321 ;
  LAYER M2 ;
        RECT 9.68 19.403 12.08 19.405 ;
  LAYER M2 ;
        RECT 9.68 19.487 12.08 19.489 ;
  LAYER M2 ;
        RECT 9.68 19.5705 12.08 19.5725 ;
  LAYER M2 ;
        RECT 9.68 19.655 12.08 19.657 ;
  LAYER M2 ;
        RECT 9.68 19.739 12.08 19.741 ;
  LAYER M2 ;
        RECT 9.68 19.823 12.08 19.825 ;
  LAYER M2 ;
        RECT 9.68 19.907 12.08 19.909 ;
  LAYER M2 ;
        RECT 9.68 19.991 12.08 19.993 ;
  LAYER M2 ;
        RECT 9.68 20.075 12.08 20.077 ;
  LAYER M2 ;
        RECT 9.68 20.159 12.08 20.161 ;
  LAYER M2 ;
        RECT 9.68 20.243 12.08 20.245 ;
  LAYER M2 ;
        RECT 9.68 20.327 12.08 20.329 ;
  LAYER M2 ;
        RECT 9.68 20.411 12.08 20.413 ;
  LAYER M2 ;
        RECT 9.68 20.495 12.08 20.497 ;
  LAYER M2 ;
        RECT 9.68 20.579 12.08 20.581 ;
  LAYER M2 ;
        RECT 9.68 20.663 12.08 20.665 ;
  LAYER M2 ;
        RECT 9.68 20.747 12.08 20.749 ;
  LAYER M2 ;
        RECT 9.68 20.831 12.08 20.833 ;
  LAYER M2 ;
        RECT 9.68 20.915 12.08 20.917 ;
  LAYER M1 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M1 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M1 ;
        RECT 12.992 0.888 13.024 3.396 ;
  LAYER M1 ;
        RECT 13.056 0.888 13.088 3.396 ;
  LAYER M1 ;
        RECT 13.12 0.888 13.152 3.396 ;
  LAYER M1 ;
        RECT 13.184 0.888 13.216 3.396 ;
  LAYER M1 ;
        RECT 13.248 0.888 13.28 3.396 ;
  LAYER M1 ;
        RECT 13.312 0.888 13.344 3.396 ;
  LAYER M1 ;
        RECT 13.376 0.888 13.408 3.396 ;
  LAYER M1 ;
        RECT 13.44 0.888 13.472 3.396 ;
  LAYER M1 ;
        RECT 13.504 0.888 13.536 3.396 ;
  LAYER M1 ;
        RECT 13.568 0.888 13.6 3.396 ;
  LAYER M1 ;
        RECT 13.632 0.888 13.664 3.396 ;
  LAYER M1 ;
        RECT 13.696 0.888 13.728 3.396 ;
  LAYER M1 ;
        RECT 13.76 0.888 13.792 3.396 ;
  LAYER M1 ;
        RECT 13.824 0.888 13.856 3.396 ;
  LAYER M1 ;
        RECT 13.888 0.888 13.92 3.396 ;
  LAYER M1 ;
        RECT 13.952 0.888 13.984 3.396 ;
  LAYER M1 ;
        RECT 14.016 0.888 14.048 3.396 ;
  LAYER M1 ;
        RECT 14.08 0.888 14.112 3.396 ;
  LAYER M1 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M1 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M1 ;
        RECT 14.272 0.888 14.304 3.396 ;
  LAYER M1 ;
        RECT 14.336 0.888 14.368 3.396 ;
  LAYER M1 ;
        RECT 14.4 0.888 14.432 3.396 ;
  LAYER M1 ;
        RECT 14.464 0.888 14.496 3.396 ;
  LAYER M1 ;
        RECT 14.528 0.888 14.56 3.396 ;
  LAYER M1 ;
        RECT 14.592 0.888 14.624 3.396 ;
  LAYER M1 ;
        RECT 14.656 0.888 14.688 3.396 ;
  LAYER M1 ;
        RECT 14.72 0.888 14.752 3.396 ;
  LAYER M1 ;
        RECT 14.784 0.888 14.816 3.396 ;
  LAYER M1 ;
        RECT 14.848 0.888 14.88 3.396 ;
  LAYER M1 ;
        RECT 14.912 0.888 14.944 3.396 ;
  LAYER M1 ;
        RECT 14.976 0.888 15.008 3.396 ;
  LAYER M1 ;
        RECT 15.04 0.888 15.072 3.396 ;
  LAYER M1 ;
        RECT 15.104 0.888 15.136 3.396 ;
  LAYER M1 ;
        RECT 15.168 0.888 15.2 3.396 ;
  LAYER M2 ;
        RECT 12.844 0.972 15.316 1.004 ;
  LAYER M2 ;
        RECT 12.844 1.036 15.316 1.068 ;
  LAYER M2 ;
        RECT 12.844 1.1 15.316 1.132 ;
  LAYER M2 ;
        RECT 12.844 1.164 15.316 1.196 ;
  LAYER M2 ;
        RECT 12.844 1.228 15.316 1.26 ;
  LAYER M2 ;
        RECT 12.844 1.292 15.316 1.324 ;
  LAYER M2 ;
        RECT 12.844 1.356 15.316 1.388 ;
  LAYER M2 ;
        RECT 12.844 1.42 15.316 1.452 ;
  LAYER M2 ;
        RECT 12.844 1.484 15.316 1.516 ;
  LAYER M2 ;
        RECT 12.844 1.548 15.316 1.58 ;
  LAYER M2 ;
        RECT 12.844 1.612 15.316 1.644 ;
  LAYER M2 ;
        RECT 12.844 1.676 15.316 1.708 ;
  LAYER M2 ;
        RECT 12.844 1.74 15.316 1.772 ;
  LAYER M2 ;
        RECT 12.844 1.804 15.316 1.836 ;
  LAYER M2 ;
        RECT 12.844 1.868 15.316 1.9 ;
  LAYER M2 ;
        RECT 12.844 1.932 15.316 1.964 ;
  LAYER M2 ;
        RECT 12.844 1.996 15.316 2.028 ;
  LAYER M2 ;
        RECT 12.844 2.06 15.316 2.092 ;
  LAYER M2 ;
        RECT 12.844 2.124 15.316 2.156 ;
  LAYER M2 ;
        RECT 12.844 2.188 15.316 2.22 ;
  LAYER M2 ;
        RECT 12.844 2.252 15.316 2.284 ;
  LAYER M2 ;
        RECT 12.844 2.316 15.316 2.348 ;
  LAYER M2 ;
        RECT 12.844 2.38 15.316 2.412 ;
  LAYER M2 ;
        RECT 12.844 2.444 15.316 2.476 ;
  LAYER M2 ;
        RECT 12.844 2.508 15.316 2.54 ;
  LAYER M2 ;
        RECT 12.844 2.572 15.316 2.604 ;
  LAYER M2 ;
        RECT 12.844 2.636 15.316 2.668 ;
  LAYER M2 ;
        RECT 12.844 2.7 15.316 2.732 ;
  LAYER M2 ;
        RECT 12.844 2.764 15.316 2.796 ;
  LAYER M2 ;
        RECT 12.844 2.828 15.316 2.86 ;
  LAYER M2 ;
        RECT 12.844 2.892 15.316 2.924 ;
  LAYER M2 ;
        RECT 12.844 2.956 15.316 2.988 ;
  LAYER M2 ;
        RECT 12.844 3.02 15.316 3.052 ;
  LAYER M2 ;
        RECT 12.844 3.084 15.316 3.116 ;
  LAYER M2 ;
        RECT 12.844 3.148 15.316 3.18 ;
  LAYER M2 ;
        RECT 12.844 3.212 15.316 3.244 ;
  LAYER M3 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M3 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M3 ;
        RECT 12.992 0.888 13.024 3.396 ;
  LAYER M3 ;
        RECT 13.056 0.888 13.088 3.396 ;
  LAYER M3 ;
        RECT 13.12 0.888 13.152 3.396 ;
  LAYER M3 ;
        RECT 13.184 0.888 13.216 3.396 ;
  LAYER M3 ;
        RECT 13.248 0.888 13.28 3.396 ;
  LAYER M3 ;
        RECT 13.312 0.888 13.344 3.396 ;
  LAYER M3 ;
        RECT 13.376 0.888 13.408 3.396 ;
  LAYER M3 ;
        RECT 13.44 0.888 13.472 3.396 ;
  LAYER M3 ;
        RECT 13.504 0.888 13.536 3.396 ;
  LAYER M3 ;
        RECT 13.568 0.888 13.6 3.396 ;
  LAYER M3 ;
        RECT 13.632 0.888 13.664 3.396 ;
  LAYER M3 ;
        RECT 13.696 0.888 13.728 3.396 ;
  LAYER M3 ;
        RECT 13.76 0.888 13.792 3.396 ;
  LAYER M3 ;
        RECT 13.824 0.888 13.856 3.396 ;
  LAYER M3 ;
        RECT 13.888 0.888 13.92 3.396 ;
  LAYER M3 ;
        RECT 13.952 0.888 13.984 3.396 ;
  LAYER M3 ;
        RECT 14.016 0.888 14.048 3.396 ;
  LAYER M3 ;
        RECT 14.08 0.888 14.112 3.396 ;
  LAYER M3 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M3 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M3 ;
        RECT 14.272 0.888 14.304 3.396 ;
  LAYER M3 ;
        RECT 14.336 0.888 14.368 3.396 ;
  LAYER M3 ;
        RECT 14.4 0.888 14.432 3.396 ;
  LAYER M3 ;
        RECT 14.464 0.888 14.496 3.396 ;
  LAYER M3 ;
        RECT 14.528 0.888 14.56 3.396 ;
  LAYER M3 ;
        RECT 14.592 0.888 14.624 3.396 ;
  LAYER M3 ;
        RECT 14.656 0.888 14.688 3.396 ;
  LAYER M3 ;
        RECT 14.72 0.888 14.752 3.396 ;
  LAYER M3 ;
        RECT 14.784 0.888 14.816 3.396 ;
  LAYER M3 ;
        RECT 14.848 0.888 14.88 3.396 ;
  LAYER M3 ;
        RECT 14.912 0.888 14.944 3.396 ;
  LAYER M3 ;
        RECT 14.976 0.888 15.008 3.396 ;
  LAYER M3 ;
        RECT 15.04 0.888 15.072 3.396 ;
  LAYER M3 ;
        RECT 15.104 0.888 15.136 3.396 ;
  LAYER M3 ;
        RECT 15.168 0.888 15.2 3.396 ;
  LAYER M3 ;
        RECT 15.264 0.888 15.296 3.396 ;
  LAYER M1 ;
        RECT 12.879 0.924 12.881 3.36 ;
  LAYER M1 ;
        RECT 12.959 0.924 12.961 3.36 ;
  LAYER M1 ;
        RECT 13.039 0.924 13.041 3.36 ;
  LAYER M1 ;
        RECT 13.119 0.924 13.121 3.36 ;
  LAYER M1 ;
        RECT 13.199 0.924 13.201 3.36 ;
  LAYER M1 ;
        RECT 13.279 0.924 13.281 3.36 ;
  LAYER M1 ;
        RECT 13.359 0.924 13.361 3.36 ;
  LAYER M1 ;
        RECT 13.439 0.924 13.441 3.36 ;
  LAYER M1 ;
        RECT 13.519 0.924 13.521 3.36 ;
  LAYER M1 ;
        RECT 13.599 0.924 13.601 3.36 ;
  LAYER M1 ;
        RECT 13.679 0.924 13.681 3.36 ;
  LAYER M1 ;
        RECT 13.759 0.924 13.761 3.36 ;
  LAYER M1 ;
        RECT 13.839 0.924 13.841 3.36 ;
  LAYER M1 ;
        RECT 13.919 0.924 13.921 3.36 ;
  LAYER M1 ;
        RECT 13.999 0.924 14.001 3.36 ;
  LAYER M1 ;
        RECT 14.079 0.924 14.081 3.36 ;
  LAYER M1 ;
        RECT 14.159 0.924 14.161 3.36 ;
  LAYER M1 ;
        RECT 14.239 0.924 14.241 3.36 ;
  LAYER M1 ;
        RECT 14.319 0.924 14.321 3.36 ;
  LAYER M1 ;
        RECT 14.399 0.924 14.401 3.36 ;
  LAYER M1 ;
        RECT 14.479 0.924 14.481 3.36 ;
  LAYER M1 ;
        RECT 14.559 0.924 14.561 3.36 ;
  LAYER M1 ;
        RECT 14.639 0.924 14.641 3.36 ;
  LAYER M1 ;
        RECT 14.719 0.924 14.721 3.36 ;
  LAYER M1 ;
        RECT 14.799 0.924 14.801 3.36 ;
  LAYER M1 ;
        RECT 14.879 0.924 14.881 3.36 ;
  LAYER M1 ;
        RECT 14.959 0.924 14.961 3.36 ;
  LAYER M1 ;
        RECT 15.039 0.924 15.041 3.36 ;
  LAYER M1 ;
        RECT 15.119 0.924 15.121 3.36 ;
  LAYER M1 ;
        RECT 15.199 0.924 15.201 3.36 ;
  LAYER M2 ;
        RECT 12.88 0.923 15.28 0.925 ;
  LAYER M2 ;
        RECT 12.88 1.007 15.28 1.009 ;
  LAYER M2 ;
        RECT 12.88 1.091 15.28 1.093 ;
  LAYER M2 ;
        RECT 12.88 1.175 15.28 1.177 ;
  LAYER M2 ;
        RECT 12.88 1.259 15.28 1.261 ;
  LAYER M2 ;
        RECT 12.88 1.343 15.28 1.345 ;
  LAYER M2 ;
        RECT 12.88 1.427 15.28 1.429 ;
  LAYER M2 ;
        RECT 12.88 1.511 15.28 1.513 ;
  LAYER M2 ;
        RECT 12.88 1.595 15.28 1.597 ;
  LAYER M2 ;
        RECT 12.88 1.679 15.28 1.681 ;
  LAYER M2 ;
        RECT 12.88 1.763 15.28 1.765 ;
  LAYER M2 ;
        RECT 12.88 1.847 15.28 1.849 ;
  LAYER M2 ;
        RECT 12.88 1.9305 15.28 1.9325 ;
  LAYER M2 ;
        RECT 12.88 2.015 15.28 2.017 ;
  LAYER M2 ;
        RECT 12.88 2.099 15.28 2.101 ;
  LAYER M2 ;
        RECT 12.88 2.183 15.28 2.185 ;
  LAYER M2 ;
        RECT 12.88 2.267 15.28 2.269 ;
  LAYER M2 ;
        RECT 12.88 2.351 15.28 2.353 ;
  LAYER M2 ;
        RECT 12.88 2.435 15.28 2.437 ;
  LAYER M2 ;
        RECT 12.88 2.519 15.28 2.521 ;
  LAYER M2 ;
        RECT 12.88 2.603 15.28 2.605 ;
  LAYER M2 ;
        RECT 12.88 2.687 15.28 2.689 ;
  LAYER M2 ;
        RECT 12.88 2.771 15.28 2.773 ;
  LAYER M2 ;
        RECT 12.88 2.855 15.28 2.857 ;
  LAYER M2 ;
        RECT 12.88 2.939 15.28 2.941 ;
  LAYER M2 ;
        RECT 12.88 3.023 15.28 3.025 ;
  LAYER M2 ;
        RECT 12.88 3.107 15.28 3.109 ;
  LAYER M2 ;
        RECT 12.88 3.191 15.28 3.193 ;
  LAYER M2 ;
        RECT 12.88 3.275 15.28 3.277 ;
  LAYER M1 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M1 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M1 ;
        RECT 12.992 3.828 13.024 6.336 ;
  LAYER M1 ;
        RECT 13.056 3.828 13.088 6.336 ;
  LAYER M1 ;
        RECT 13.12 3.828 13.152 6.336 ;
  LAYER M1 ;
        RECT 13.184 3.828 13.216 6.336 ;
  LAYER M1 ;
        RECT 13.248 3.828 13.28 6.336 ;
  LAYER M1 ;
        RECT 13.312 3.828 13.344 6.336 ;
  LAYER M1 ;
        RECT 13.376 3.828 13.408 6.336 ;
  LAYER M1 ;
        RECT 13.44 3.828 13.472 6.336 ;
  LAYER M1 ;
        RECT 13.504 3.828 13.536 6.336 ;
  LAYER M1 ;
        RECT 13.568 3.828 13.6 6.336 ;
  LAYER M1 ;
        RECT 13.632 3.828 13.664 6.336 ;
  LAYER M1 ;
        RECT 13.696 3.828 13.728 6.336 ;
  LAYER M1 ;
        RECT 13.76 3.828 13.792 6.336 ;
  LAYER M1 ;
        RECT 13.824 3.828 13.856 6.336 ;
  LAYER M1 ;
        RECT 13.888 3.828 13.92 6.336 ;
  LAYER M1 ;
        RECT 13.952 3.828 13.984 6.336 ;
  LAYER M1 ;
        RECT 14.016 3.828 14.048 6.336 ;
  LAYER M1 ;
        RECT 14.08 3.828 14.112 6.336 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M1 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M1 ;
        RECT 14.272 3.828 14.304 6.336 ;
  LAYER M1 ;
        RECT 14.336 3.828 14.368 6.336 ;
  LAYER M1 ;
        RECT 14.4 3.828 14.432 6.336 ;
  LAYER M1 ;
        RECT 14.464 3.828 14.496 6.336 ;
  LAYER M1 ;
        RECT 14.528 3.828 14.56 6.336 ;
  LAYER M1 ;
        RECT 14.592 3.828 14.624 6.336 ;
  LAYER M1 ;
        RECT 14.656 3.828 14.688 6.336 ;
  LAYER M1 ;
        RECT 14.72 3.828 14.752 6.336 ;
  LAYER M1 ;
        RECT 14.784 3.828 14.816 6.336 ;
  LAYER M1 ;
        RECT 14.848 3.828 14.88 6.336 ;
  LAYER M1 ;
        RECT 14.912 3.828 14.944 6.336 ;
  LAYER M1 ;
        RECT 14.976 3.828 15.008 6.336 ;
  LAYER M1 ;
        RECT 15.04 3.828 15.072 6.336 ;
  LAYER M1 ;
        RECT 15.104 3.828 15.136 6.336 ;
  LAYER M1 ;
        RECT 15.168 3.828 15.2 6.336 ;
  LAYER M2 ;
        RECT 12.844 3.912 15.316 3.944 ;
  LAYER M2 ;
        RECT 12.844 3.976 15.316 4.008 ;
  LAYER M2 ;
        RECT 12.844 4.04 15.316 4.072 ;
  LAYER M2 ;
        RECT 12.844 4.104 15.316 4.136 ;
  LAYER M2 ;
        RECT 12.844 4.168 15.316 4.2 ;
  LAYER M2 ;
        RECT 12.844 4.232 15.316 4.264 ;
  LAYER M2 ;
        RECT 12.844 4.296 15.316 4.328 ;
  LAYER M2 ;
        RECT 12.844 4.36 15.316 4.392 ;
  LAYER M2 ;
        RECT 12.844 4.424 15.316 4.456 ;
  LAYER M2 ;
        RECT 12.844 4.488 15.316 4.52 ;
  LAYER M2 ;
        RECT 12.844 4.552 15.316 4.584 ;
  LAYER M2 ;
        RECT 12.844 4.616 15.316 4.648 ;
  LAYER M2 ;
        RECT 12.844 4.68 15.316 4.712 ;
  LAYER M2 ;
        RECT 12.844 4.744 15.316 4.776 ;
  LAYER M2 ;
        RECT 12.844 4.808 15.316 4.84 ;
  LAYER M2 ;
        RECT 12.844 4.872 15.316 4.904 ;
  LAYER M2 ;
        RECT 12.844 4.936 15.316 4.968 ;
  LAYER M2 ;
        RECT 12.844 5 15.316 5.032 ;
  LAYER M2 ;
        RECT 12.844 5.064 15.316 5.096 ;
  LAYER M2 ;
        RECT 12.844 5.128 15.316 5.16 ;
  LAYER M2 ;
        RECT 12.844 5.192 15.316 5.224 ;
  LAYER M2 ;
        RECT 12.844 5.256 15.316 5.288 ;
  LAYER M2 ;
        RECT 12.844 5.32 15.316 5.352 ;
  LAYER M2 ;
        RECT 12.844 5.384 15.316 5.416 ;
  LAYER M2 ;
        RECT 12.844 5.448 15.316 5.48 ;
  LAYER M2 ;
        RECT 12.844 5.512 15.316 5.544 ;
  LAYER M2 ;
        RECT 12.844 5.576 15.316 5.608 ;
  LAYER M2 ;
        RECT 12.844 5.64 15.316 5.672 ;
  LAYER M2 ;
        RECT 12.844 5.704 15.316 5.736 ;
  LAYER M2 ;
        RECT 12.844 5.768 15.316 5.8 ;
  LAYER M2 ;
        RECT 12.844 5.832 15.316 5.864 ;
  LAYER M2 ;
        RECT 12.844 5.896 15.316 5.928 ;
  LAYER M2 ;
        RECT 12.844 5.96 15.316 5.992 ;
  LAYER M2 ;
        RECT 12.844 6.024 15.316 6.056 ;
  LAYER M2 ;
        RECT 12.844 6.088 15.316 6.12 ;
  LAYER M2 ;
        RECT 12.844 6.152 15.316 6.184 ;
  LAYER M3 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M3 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M3 ;
        RECT 12.992 3.828 13.024 6.336 ;
  LAYER M3 ;
        RECT 13.056 3.828 13.088 6.336 ;
  LAYER M3 ;
        RECT 13.12 3.828 13.152 6.336 ;
  LAYER M3 ;
        RECT 13.184 3.828 13.216 6.336 ;
  LAYER M3 ;
        RECT 13.248 3.828 13.28 6.336 ;
  LAYER M3 ;
        RECT 13.312 3.828 13.344 6.336 ;
  LAYER M3 ;
        RECT 13.376 3.828 13.408 6.336 ;
  LAYER M3 ;
        RECT 13.44 3.828 13.472 6.336 ;
  LAYER M3 ;
        RECT 13.504 3.828 13.536 6.336 ;
  LAYER M3 ;
        RECT 13.568 3.828 13.6 6.336 ;
  LAYER M3 ;
        RECT 13.632 3.828 13.664 6.336 ;
  LAYER M3 ;
        RECT 13.696 3.828 13.728 6.336 ;
  LAYER M3 ;
        RECT 13.76 3.828 13.792 6.336 ;
  LAYER M3 ;
        RECT 13.824 3.828 13.856 6.336 ;
  LAYER M3 ;
        RECT 13.888 3.828 13.92 6.336 ;
  LAYER M3 ;
        RECT 13.952 3.828 13.984 6.336 ;
  LAYER M3 ;
        RECT 14.016 3.828 14.048 6.336 ;
  LAYER M3 ;
        RECT 14.08 3.828 14.112 6.336 ;
  LAYER M3 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M3 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M3 ;
        RECT 14.272 3.828 14.304 6.336 ;
  LAYER M3 ;
        RECT 14.336 3.828 14.368 6.336 ;
  LAYER M3 ;
        RECT 14.4 3.828 14.432 6.336 ;
  LAYER M3 ;
        RECT 14.464 3.828 14.496 6.336 ;
  LAYER M3 ;
        RECT 14.528 3.828 14.56 6.336 ;
  LAYER M3 ;
        RECT 14.592 3.828 14.624 6.336 ;
  LAYER M3 ;
        RECT 14.656 3.828 14.688 6.336 ;
  LAYER M3 ;
        RECT 14.72 3.828 14.752 6.336 ;
  LAYER M3 ;
        RECT 14.784 3.828 14.816 6.336 ;
  LAYER M3 ;
        RECT 14.848 3.828 14.88 6.336 ;
  LAYER M3 ;
        RECT 14.912 3.828 14.944 6.336 ;
  LAYER M3 ;
        RECT 14.976 3.828 15.008 6.336 ;
  LAYER M3 ;
        RECT 15.04 3.828 15.072 6.336 ;
  LAYER M3 ;
        RECT 15.104 3.828 15.136 6.336 ;
  LAYER M3 ;
        RECT 15.168 3.828 15.2 6.336 ;
  LAYER M3 ;
        RECT 15.264 3.828 15.296 6.336 ;
  LAYER M1 ;
        RECT 12.879 3.864 12.881 6.3 ;
  LAYER M1 ;
        RECT 12.959 3.864 12.961 6.3 ;
  LAYER M1 ;
        RECT 13.039 3.864 13.041 6.3 ;
  LAYER M1 ;
        RECT 13.119 3.864 13.121 6.3 ;
  LAYER M1 ;
        RECT 13.199 3.864 13.201 6.3 ;
  LAYER M1 ;
        RECT 13.279 3.864 13.281 6.3 ;
  LAYER M1 ;
        RECT 13.359 3.864 13.361 6.3 ;
  LAYER M1 ;
        RECT 13.439 3.864 13.441 6.3 ;
  LAYER M1 ;
        RECT 13.519 3.864 13.521 6.3 ;
  LAYER M1 ;
        RECT 13.599 3.864 13.601 6.3 ;
  LAYER M1 ;
        RECT 13.679 3.864 13.681 6.3 ;
  LAYER M1 ;
        RECT 13.759 3.864 13.761 6.3 ;
  LAYER M1 ;
        RECT 13.839 3.864 13.841 6.3 ;
  LAYER M1 ;
        RECT 13.919 3.864 13.921 6.3 ;
  LAYER M1 ;
        RECT 13.999 3.864 14.001 6.3 ;
  LAYER M1 ;
        RECT 14.079 3.864 14.081 6.3 ;
  LAYER M1 ;
        RECT 14.159 3.864 14.161 6.3 ;
  LAYER M1 ;
        RECT 14.239 3.864 14.241 6.3 ;
  LAYER M1 ;
        RECT 14.319 3.864 14.321 6.3 ;
  LAYER M1 ;
        RECT 14.399 3.864 14.401 6.3 ;
  LAYER M1 ;
        RECT 14.479 3.864 14.481 6.3 ;
  LAYER M1 ;
        RECT 14.559 3.864 14.561 6.3 ;
  LAYER M1 ;
        RECT 14.639 3.864 14.641 6.3 ;
  LAYER M1 ;
        RECT 14.719 3.864 14.721 6.3 ;
  LAYER M1 ;
        RECT 14.799 3.864 14.801 6.3 ;
  LAYER M1 ;
        RECT 14.879 3.864 14.881 6.3 ;
  LAYER M1 ;
        RECT 14.959 3.864 14.961 6.3 ;
  LAYER M1 ;
        RECT 15.039 3.864 15.041 6.3 ;
  LAYER M1 ;
        RECT 15.119 3.864 15.121 6.3 ;
  LAYER M1 ;
        RECT 15.199 3.864 15.201 6.3 ;
  LAYER M2 ;
        RECT 12.88 3.863 15.28 3.865 ;
  LAYER M2 ;
        RECT 12.88 3.947 15.28 3.949 ;
  LAYER M2 ;
        RECT 12.88 4.031 15.28 4.033 ;
  LAYER M2 ;
        RECT 12.88 4.115 15.28 4.117 ;
  LAYER M2 ;
        RECT 12.88 4.199 15.28 4.201 ;
  LAYER M2 ;
        RECT 12.88 4.283 15.28 4.285 ;
  LAYER M2 ;
        RECT 12.88 4.367 15.28 4.369 ;
  LAYER M2 ;
        RECT 12.88 4.451 15.28 4.453 ;
  LAYER M2 ;
        RECT 12.88 4.535 15.28 4.537 ;
  LAYER M2 ;
        RECT 12.88 4.619 15.28 4.621 ;
  LAYER M2 ;
        RECT 12.88 4.703 15.28 4.705 ;
  LAYER M2 ;
        RECT 12.88 4.787 15.28 4.789 ;
  LAYER M2 ;
        RECT 12.88 4.8705 15.28 4.8725 ;
  LAYER M2 ;
        RECT 12.88 4.955 15.28 4.957 ;
  LAYER M2 ;
        RECT 12.88 5.039 15.28 5.041 ;
  LAYER M2 ;
        RECT 12.88 5.123 15.28 5.125 ;
  LAYER M2 ;
        RECT 12.88 5.207 15.28 5.209 ;
  LAYER M2 ;
        RECT 12.88 5.291 15.28 5.293 ;
  LAYER M2 ;
        RECT 12.88 5.375 15.28 5.377 ;
  LAYER M2 ;
        RECT 12.88 5.459 15.28 5.461 ;
  LAYER M2 ;
        RECT 12.88 5.543 15.28 5.545 ;
  LAYER M2 ;
        RECT 12.88 5.627 15.28 5.629 ;
  LAYER M2 ;
        RECT 12.88 5.711 15.28 5.713 ;
  LAYER M2 ;
        RECT 12.88 5.795 15.28 5.797 ;
  LAYER M2 ;
        RECT 12.88 5.879 15.28 5.881 ;
  LAYER M2 ;
        RECT 12.88 5.963 15.28 5.965 ;
  LAYER M2 ;
        RECT 12.88 6.047 15.28 6.049 ;
  LAYER M2 ;
        RECT 12.88 6.131 15.28 6.133 ;
  LAYER M2 ;
        RECT 12.88 6.215 15.28 6.217 ;
  LAYER M1 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M1 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M1 ;
        RECT 12.992 6.768 13.024 9.276 ;
  LAYER M1 ;
        RECT 13.056 6.768 13.088 9.276 ;
  LAYER M1 ;
        RECT 13.12 6.768 13.152 9.276 ;
  LAYER M1 ;
        RECT 13.184 6.768 13.216 9.276 ;
  LAYER M1 ;
        RECT 13.248 6.768 13.28 9.276 ;
  LAYER M1 ;
        RECT 13.312 6.768 13.344 9.276 ;
  LAYER M1 ;
        RECT 13.376 6.768 13.408 9.276 ;
  LAYER M1 ;
        RECT 13.44 6.768 13.472 9.276 ;
  LAYER M1 ;
        RECT 13.504 6.768 13.536 9.276 ;
  LAYER M1 ;
        RECT 13.568 6.768 13.6 9.276 ;
  LAYER M1 ;
        RECT 13.632 6.768 13.664 9.276 ;
  LAYER M1 ;
        RECT 13.696 6.768 13.728 9.276 ;
  LAYER M1 ;
        RECT 13.76 6.768 13.792 9.276 ;
  LAYER M1 ;
        RECT 13.824 6.768 13.856 9.276 ;
  LAYER M1 ;
        RECT 13.888 6.768 13.92 9.276 ;
  LAYER M1 ;
        RECT 13.952 6.768 13.984 9.276 ;
  LAYER M1 ;
        RECT 14.016 6.768 14.048 9.276 ;
  LAYER M1 ;
        RECT 14.08 6.768 14.112 9.276 ;
  LAYER M1 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M1 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M1 ;
        RECT 14.272 6.768 14.304 9.276 ;
  LAYER M1 ;
        RECT 14.336 6.768 14.368 9.276 ;
  LAYER M1 ;
        RECT 14.4 6.768 14.432 9.276 ;
  LAYER M1 ;
        RECT 14.464 6.768 14.496 9.276 ;
  LAYER M1 ;
        RECT 14.528 6.768 14.56 9.276 ;
  LAYER M1 ;
        RECT 14.592 6.768 14.624 9.276 ;
  LAYER M1 ;
        RECT 14.656 6.768 14.688 9.276 ;
  LAYER M1 ;
        RECT 14.72 6.768 14.752 9.276 ;
  LAYER M1 ;
        RECT 14.784 6.768 14.816 9.276 ;
  LAYER M1 ;
        RECT 14.848 6.768 14.88 9.276 ;
  LAYER M1 ;
        RECT 14.912 6.768 14.944 9.276 ;
  LAYER M1 ;
        RECT 14.976 6.768 15.008 9.276 ;
  LAYER M1 ;
        RECT 15.04 6.768 15.072 9.276 ;
  LAYER M1 ;
        RECT 15.104 6.768 15.136 9.276 ;
  LAYER M1 ;
        RECT 15.168 6.768 15.2 9.276 ;
  LAYER M2 ;
        RECT 12.844 6.852 15.316 6.884 ;
  LAYER M2 ;
        RECT 12.844 6.916 15.316 6.948 ;
  LAYER M2 ;
        RECT 12.844 6.98 15.316 7.012 ;
  LAYER M2 ;
        RECT 12.844 7.044 15.316 7.076 ;
  LAYER M2 ;
        RECT 12.844 7.108 15.316 7.14 ;
  LAYER M2 ;
        RECT 12.844 7.172 15.316 7.204 ;
  LAYER M2 ;
        RECT 12.844 7.236 15.316 7.268 ;
  LAYER M2 ;
        RECT 12.844 7.3 15.316 7.332 ;
  LAYER M2 ;
        RECT 12.844 7.364 15.316 7.396 ;
  LAYER M2 ;
        RECT 12.844 7.428 15.316 7.46 ;
  LAYER M2 ;
        RECT 12.844 7.492 15.316 7.524 ;
  LAYER M2 ;
        RECT 12.844 7.556 15.316 7.588 ;
  LAYER M2 ;
        RECT 12.844 7.62 15.316 7.652 ;
  LAYER M2 ;
        RECT 12.844 7.684 15.316 7.716 ;
  LAYER M2 ;
        RECT 12.844 7.748 15.316 7.78 ;
  LAYER M2 ;
        RECT 12.844 7.812 15.316 7.844 ;
  LAYER M2 ;
        RECT 12.844 7.876 15.316 7.908 ;
  LAYER M2 ;
        RECT 12.844 7.94 15.316 7.972 ;
  LAYER M2 ;
        RECT 12.844 8.004 15.316 8.036 ;
  LAYER M2 ;
        RECT 12.844 8.068 15.316 8.1 ;
  LAYER M2 ;
        RECT 12.844 8.132 15.316 8.164 ;
  LAYER M2 ;
        RECT 12.844 8.196 15.316 8.228 ;
  LAYER M2 ;
        RECT 12.844 8.26 15.316 8.292 ;
  LAYER M2 ;
        RECT 12.844 8.324 15.316 8.356 ;
  LAYER M2 ;
        RECT 12.844 8.388 15.316 8.42 ;
  LAYER M2 ;
        RECT 12.844 8.452 15.316 8.484 ;
  LAYER M2 ;
        RECT 12.844 8.516 15.316 8.548 ;
  LAYER M2 ;
        RECT 12.844 8.58 15.316 8.612 ;
  LAYER M2 ;
        RECT 12.844 8.644 15.316 8.676 ;
  LAYER M2 ;
        RECT 12.844 8.708 15.316 8.74 ;
  LAYER M2 ;
        RECT 12.844 8.772 15.316 8.804 ;
  LAYER M2 ;
        RECT 12.844 8.836 15.316 8.868 ;
  LAYER M2 ;
        RECT 12.844 8.9 15.316 8.932 ;
  LAYER M2 ;
        RECT 12.844 8.964 15.316 8.996 ;
  LAYER M2 ;
        RECT 12.844 9.028 15.316 9.06 ;
  LAYER M2 ;
        RECT 12.844 9.092 15.316 9.124 ;
  LAYER M3 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M3 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M3 ;
        RECT 12.992 6.768 13.024 9.276 ;
  LAYER M3 ;
        RECT 13.056 6.768 13.088 9.276 ;
  LAYER M3 ;
        RECT 13.12 6.768 13.152 9.276 ;
  LAYER M3 ;
        RECT 13.184 6.768 13.216 9.276 ;
  LAYER M3 ;
        RECT 13.248 6.768 13.28 9.276 ;
  LAYER M3 ;
        RECT 13.312 6.768 13.344 9.276 ;
  LAYER M3 ;
        RECT 13.376 6.768 13.408 9.276 ;
  LAYER M3 ;
        RECT 13.44 6.768 13.472 9.276 ;
  LAYER M3 ;
        RECT 13.504 6.768 13.536 9.276 ;
  LAYER M3 ;
        RECT 13.568 6.768 13.6 9.276 ;
  LAYER M3 ;
        RECT 13.632 6.768 13.664 9.276 ;
  LAYER M3 ;
        RECT 13.696 6.768 13.728 9.276 ;
  LAYER M3 ;
        RECT 13.76 6.768 13.792 9.276 ;
  LAYER M3 ;
        RECT 13.824 6.768 13.856 9.276 ;
  LAYER M3 ;
        RECT 13.888 6.768 13.92 9.276 ;
  LAYER M3 ;
        RECT 13.952 6.768 13.984 9.276 ;
  LAYER M3 ;
        RECT 14.016 6.768 14.048 9.276 ;
  LAYER M3 ;
        RECT 14.08 6.768 14.112 9.276 ;
  LAYER M3 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M3 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M3 ;
        RECT 14.272 6.768 14.304 9.276 ;
  LAYER M3 ;
        RECT 14.336 6.768 14.368 9.276 ;
  LAYER M3 ;
        RECT 14.4 6.768 14.432 9.276 ;
  LAYER M3 ;
        RECT 14.464 6.768 14.496 9.276 ;
  LAYER M3 ;
        RECT 14.528 6.768 14.56 9.276 ;
  LAYER M3 ;
        RECT 14.592 6.768 14.624 9.276 ;
  LAYER M3 ;
        RECT 14.656 6.768 14.688 9.276 ;
  LAYER M3 ;
        RECT 14.72 6.768 14.752 9.276 ;
  LAYER M3 ;
        RECT 14.784 6.768 14.816 9.276 ;
  LAYER M3 ;
        RECT 14.848 6.768 14.88 9.276 ;
  LAYER M3 ;
        RECT 14.912 6.768 14.944 9.276 ;
  LAYER M3 ;
        RECT 14.976 6.768 15.008 9.276 ;
  LAYER M3 ;
        RECT 15.04 6.768 15.072 9.276 ;
  LAYER M3 ;
        RECT 15.104 6.768 15.136 9.276 ;
  LAYER M3 ;
        RECT 15.168 6.768 15.2 9.276 ;
  LAYER M3 ;
        RECT 15.264 6.768 15.296 9.276 ;
  LAYER M1 ;
        RECT 12.879 6.804 12.881 9.24 ;
  LAYER M1 ;
        RECT 12.959 6.804 12.961 9.24 ;
  LAYER M1 ;
        RECT 13.039 6.804 13.041 9.24 ;
  LAYER M1 ;
        RECT 13.119 6.804 13.121 9.24 ;
  LAYER M1 ;
        RECT 13.199 6.804 13.201 9.24 ;
  LAYER M1 ;
        RECT 13.279 6.804 13.281 9.24 ;
  LAYER M1 ;
        RECT 13.359 6.804 13.361 9.24 ;
  LAYER M1 ;
        RECT 13.439 6.804 13.441 9.24 ;
  LAYER M1 ;
        RECT 13.519 6.804 13.521 9.24 ;
  LAYER M1 ;
        RECT 13.599 6.804 13.601 9.24 ;
  LAYER M1 ;
        RECT 13.679 6.804 13.681 9.24 ;
  LAYER M1 ;
        RECT 13.759 6.804 13.761 9.24 ;
  LAYER M1 ;
        RECT 13.839 6.804 13.841 9.24 ;
  LAYER M1 ;
        RECT 13.919 6.804 13.921 9.24 ;
  LAYER M1 ;
        RECT 13.999 6.804 14.001 9.24 ;
  LAYER M1 ;
        RECT 14.079 6.804 14.081 9.24 ;
  LAYER M1 ;
        RECT 14.159 6.804 14.161 9.24 ;
  LAYER M1 ;
        RECT 14.239 6.804 14.241 9.24 ;
  LAYER M1 ;
        RECT 14.319 6.804 14.321 9.24 ;
  LAYER M1 ;
        RECT 14.399 6.804 14.401 9.24 ;
  LAYER M1 ;
        RECT 14.479 6.804 14.481 9.24 ;
  LAYER M1 ;
        RECT 14.559 6.804 14.561 9.24 ;
  LAYER M1 ;
        RECT 14.639 6.804 14.641 9.24 ;
  LAYER M1 ;
        RECT 14.719 6.804 14.721 9.24 ;
  LAYER M1 ;
        RECT 14.799 6.804 14.801 9.24 ;
  LAYER M1 ;
        RECT 14.879 6.804 14.881 9.24 ;
  LAYER M1 ;
        RECT 14.959 6.804 14.961 9.24 ;
  LAYER M1 ;
        RECT 15.039 6.804 15.041 9.24 ;
  LAYER M1 ;
        RECT 15.119 6.804 15.121 9.24 ;
  LAYER M1 ;
        RECT 15.199 6.804 15.201 9.24 ;
  LAYER M2 ;
        RECT 12.88 6.803 15.28 6.805 ;
  LAYER M2 ;
        RECT 12.88 6.887 15.28 6.889 ;
  LAYER M2 ;
        RECT 12.88 6.971 15.28 6.973 ;
  LAYER M2 ;
        RECT 12.88 7.055 15.28 7.057 ;
  LAYER M2 ;
        RECT 12.88 7.139 15.28 7.141 ;
  LAYER M2 ;
        RECT 12.88 7.223 15.28 7.225 ;
  LAYER M2 ;
        RECT 12.88 7.307 15.28 7.309 ;
  LAYER M2 ;
        RECT 12.88 7.391 15.28 7.393 ;
  LAYER M2 ;
        RECT 12.88 7.475 15.28 7.477 ;
  LAYER M2 ;
        RECT 12.88 7.559 15.28 7.561 ;
  LAYER M2 ;
        RECT 12.88 7.643 15.28 7.645 ;
  LAYER M2 ;
        RECT 12.88 7.727 15.28 7.729 ;
  LAYER M2 ;
        RECT 12.88 7.8105 15.28 7.8125 ;
  LAYER M2 ;
        RECT 12.88 7.895 15.28 7.897 ;
  LAYER M2 ;
        RECT 12.88 7.979 15.28 7.981 ;
  LAYER M2 ;
        RECT 12.88 8.063 15.28 8.065 ;
  LAYER M2 ;
        RECT 12.88 8.147 15.28 8.149 ;
  LAYER M2 ;
        RECT 12.88 8.231 15.28 8.233 ;
  LAYER M2 ;
        RECT 12.88 8.315 15.28 8.317 ;
  LAYER M2 ;
        RECT 12.88 8.399 15.28 8.401 ;
  LAYER M2 ;
        RECT 12.88 8.483 15.28 8.485 ;
  LAYER M2 ;
        RECT 12.88 8.567 15.28 8.569 ;
  LAYER M2 ;
        RECT 12.88 8.651 15.28 8.653 ;
  LAYER M2 ;
        RECT 12.88 8.735 15.28 8.737 ;
  LAYER M2 ;
        RECT 12.88 8.819 15.28 8.821 ;
  LAYER M2 ;
        RECT 12.88 8.903 15.28 8.905 ;
  LAYER M2 ;
        RECT 12.88 8.987 15.28 8.989 ;
  LAYER M2 ;
        RECT 12.88 9.071 15.28 9.073 ;
  LAYER M2 ;
        RECT 12.88 9.155 15.28 9.157 ;
  LAYER M1 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M1 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M1 ;
        RECT 12.992 9.708 13.024 12.216 ;
  LAYER M1 ;
        RECT 13.056 9.708 13.088 12.216 ;
  LAYER M1 ;
        RECT 13.12 9.708 13.152 12.216 ;
  LAYER M1 ;
        RECT 13.184 9.708 13.216 12.216 ;
  LAYER M1 ;
        RECT 13.248 9.708 13.28 12.216 ;
  LAYER M1 ;
        RECT 13.312 9.708 13.344 12.216 ;
  LAYER M1 ;
        RECT 13.376 9.708 13.408 12.216 ;
  LAYER M1 ;
        RECT 13.44 9.708 13.472 12.216 ;
  LAYER M1 ;
        RECT 13.504 9.708 13.536 12.216 ;
  LAYER M1 ;
        RECT 13.568 9.708 13.6 12.216 ;
  LAYER M1 ;
        RECT 13.632 9.708 13.664 12.216 ;
  LAYER M1 ;
        RECT 13.696 9.708 13.728 12.216 ;
  LAYER M1 ;
        RECT 13.76 9.708 13.792 12.216 ;
  LAYER M1 ;
        RECT 13.824 9.708 13.856 12.216 ;
  LAYER M1 ;
        RECT 13.888 9.708 13.92 12.216 ;
  LAYER M1 ;
        RECT 13.952 9.708 13.984 12.216 ;
  LAYER M1 ;
        RECT 14.016 9.708 14.048 12.216 ;
  LAYER M1 ;
        RECT 14.08 9.708 14.112 12.216 ;
  LAYER M1 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M1 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M1 ;
        RECT 14.272 9.708 14.304 12.216 ;
  LAYER M1 ;
        RECT 14.336 9.708 14.368 12.216 ;
  LAYER M1 ;
        RECT 14.4 9.708 14.432 12.216 ;
  LAYER M1 ;
        RECT 14.464 9.708 14.496 12.216 ;
  LAYER M1 ;
        RECT 14.528 9.708 14.56 12.216 ;
  LAYER M1 ;
        RECT 14.592 9.708 14.624 12.216 ;
  LAYER M1 ;
        RECT 14.656 9.708 14.688 12.216 ;
  LAYER M1 ;
        RECT 14.72 9.708 14.752 12.216 ;
  LAYER M1 ;
        RECT 14.784 9.708 14.816 12.216 ;
  LAYER M1 ;
        RECT 14.848 9.708 14.88 12.216 ;
  LAYER M1 ;
        RECT 14.912 9.708 14.944 12.216 ;
  LAYER M1 ;
        RECT 14.976 9.708 15.008 12.216 ;
  LAYER M1 ;
        RECT 15.04 9.708 15.072 12.216 ;
  LAYER M1 ;
        RECT 15.104 9.708 15.136 12.216 ;
  LAYER M1 ;
        RECT 15.168 9.708 15.2 12.216 ;
  LAYER M2 ;
        RECT 12.844 9.792 15.316 9.824 ;
  LAYER M2 ;
        RECT 12.844 9.856 15.316 9.888 ;
  LAYER M2 ;
        RECT 12.844 9.92 15.316 9.952 ;
  LAYER M2 ;
        RECT 12.844 9.984 15.316 10.016 ;
  LAYER M2 ;
        RECT 12.844 10.048 15.316 10.08 ;
  LAYER M2 ;
        RECT 12.844 10.112 15.316 10.144 ;
  LAYER M2 ;
        RECT 12.844 10.176 15.316 10.208 ;
  LAYER M2 ;
        RECT 12.844 10.24 15.316 10.272 ;
  LAYER M2 ;
        RECT 12.844 10.304 15.316 10.336 ;
  LAYER M2 ;
        RECT 12.844 10.368 15.316 10.4 ;
  LAYER M2 ;
        RECT 12.844 10.432 15.316 10.464 ;
  LAYER M2 ;
        RECT 12.844 10.496 15.316 10.528 ;
  LAYER M2 ;
        RECT 12.844 10.56 15.316 10.592 ;
  LAYER M2 ;
        RECT 12.844 10.624 15.316 10.656 ;
  LAYER M2 ;
        RECT 12.844 10.688 15.316 10.72 ;
  LAYER M2 ;
        RECT 12.844 10.752 15.316 10.784 ;
  LAYER M2 ;
        RECT 12.844 10.816 15.316 10.848 ;
  LAYER M2 ;
        RECT 12.844 10.88 15.316 10.912 ;
  LAYER M2 ;
        RECT 12.844 10.944 15.316 10.976 ;
  LAYER M2 ;
        RECT 12.844 11.008 15.316 11.04 ;
  LAYER M2 ;
        RECT 12.844 11.072 15.316 11.104 ;
  LAYER M2 ;
        RECT 12.844 11.136 15.316 11.168 ;
  LAYER M2 ;
        RECT 12.844 11.2 15.316 11.232 ;
  LAYER M2 ;
        RECT 12.844 11.264 15.316 11.296 ;
  LAYER M2 ;
        RECT 12.844 11.328 15.316 11.36 ;
  LAYER M2 ;
        RECT 12.844 11.392 15.316 11.424 ;
  LAYER M2 ;
        RECT 12.844 11.456 15.316 11.488 ;
  LAYER M2 ;
        RECT 12.844 11.52 15.316 11.552 ;
  LAYER M2 ;
        RECT 12.844 11.584 15.316 11.616 ;
  LAYER M2 ;
        RECT 12.844 11.648 15.316 11.68 ;
  LAYER M2 ;
        RECT 12.844 11.712 15.316 11.744 ;
  LAYER M2 ;
        RECT 12.844 11.776 15.316 11.808 ;
  LAYER M2 ;
        RECT 12.844 11.84 15.316 11.872 ;
  LAYER M2 ;
        RECT 12.844 11.904 15.316 11.936 ;
  LAYER M2 ;
        RECT 12.844 11.968 15.316 12 ;
  LAYER M2 ;
        RECT 12.844 12.032 15.316 12.064 ;
  LAYER M3 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M3 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M3 ;
        RECT 12.992 9.708 13.024 12.216 ;
  LAYER M3 ;
        RECT 13.056 9.708 13.088 12.216 ;
  LAYER M3 ;
        RECT 13.12 9.708 13.152 12.216 ;
  LAYER M3 ;
        RECT 13.184 9.708 13.216 12.216 ;
  LAYER M3 ;
        RECT 13.248 9.708 13.28 12.216 ;
  LAYER M3 ;
        RECT 13.312 9.708 13.344 12.216 ;
  LAYER M3 ;
        RECT 13.376 9.708 13.408 12.216 ;
  LAYER M3 ;
        RECT 13.44 9.708 13.472 12.216 ;
  LAYER M3 ;
        RECT 13.504 9.708 13.536 12.216 ;
  LAYER M3 ;
        RECT 13.568 9.708 13.6 12.216 ;
  LAYER M3 ;
        RECT 13.632 9.708 13.664 12.216 ;
  LAYER M3 ;
        RECT 13.696 9.708 13.728 12.216 ;
  LAYER M3 ;
        RECT 13.76 9.708 13.792 12.216 ;
  LAYER M3 ;
        RECT 13.824 9.708 13.856 12.216 ;
  LAYER M3 ;
        RECT 13.888 9.708 13.92 12.216 ;
  LAYER M3 ;
        RECT 13.952 9.708 13.984 12.216 ;
  LAYER M3 ;
        RECT 14.016 9.708 14.048 12.216 ;
  LAYER M3 ;
        RECT 14.08 9.708 14.112 12.216 ;
  LAYER M3 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M3 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M3 ;
        RECT 14.272 9.708 14.304 12.216 ;
  LAYER M3 ;
        RECT 14.336 9.708 14.368 12.216 ;
  LAYER M3 ;
        RECT 14.4 9.708 14.432 12.216 ;
  LAYER M3 ;
        RECT 14.464 9.708 14.496 12.216 ;
  LAYER M3 ;
        RECT 14.528 9.708 14.56 12.216 ;
  LAYER M3 ;
        RECT 14.592 9.708 14.624 12.216 ;
  LAYER M3 ;
        RECT 14.656 9.708 14.688 12.216 ;
  LAYER M3 ;
        RECT 14.72 9.708 14.752 12.216 ;
  LAYER M3 ;
        RECT 14.784 9.708 14.816 12.216 ;
  LAYER M3 ;
        RECT 14.848 9.708 14.88 12.216 ;
  LAYER M3 ;
        RECT 14.912 9.708 14.944 12.216 ;
  LAYER M3 ;
        RECT 14.976 9.708 15.008 12.216 ;
  LAYER M3 ;
        RECT 15.04 9.708 15.072 12.216 ;
  LAYER M3 ;
        RECT 15.104 9.708 15.136 12.216 ;
  LAYER M3 ;
        RECT 15.168 9.708 15.2 12.216 ;
  LAYER M3 ;
        RECT 15.264 9.708 15.296 12.216 ;
  LAYER M1 ;
        RECT 12.879 9.744 12.881 12.18 ;
  LAYER M1 ;
        RECT 12.959 9.744 12.961 12.18 ;
  LAYER M1 ;
        RECT 13.039 9.744 13.041 12.18 ;
  LAYER M1 ;
        RECT 13.119 9.744 13.121 12.18 ;
  LAYER M1 ;
        RECT 13.199 9.744 13.201 12.18 ;
  LAYER M1 ;
        RECT 13.279 9.744 13.281 12.18 ;
  LAYER M1 ;
        RECT 13.359 9.744 13.361 12.18 ;
  LAYER M1 ;
        RECT 13.439 9.744 13.441 12.18 ;
  LAYER M1 ;
        RECT 13.519 9.744 13.521 12.18 ;
  LAYER M1 ;
        RECT 13.599 9.744 13.601 12.18 ;
  LAYER M1 ;
        RECT 13.679 9.744 13.681 12.18 ;
  LAYER M1 ;
        RECT 13.759 9.744 13.761 12.18 ;
  LAYER M1 ;
        RECT 13.839 9.744 13.841 12.18 ;
  LAYER M1 ;
        RECT 13.919 9.744 13.921 12.18 ;
  LAYER M1 ;
        RECT 13.999 9.744 14.001 12.18 ;
  LAYER M1 ;
        RECT 14.079 9.744 14.081 12.18 ;
  LAYER M1 ;
        RECT 14.159 9.744 14.161 12.18 ;
  LAYER M1 ;
        RECT 14.239 9.744 14.241 12.18 ;
  LAYER M1 ;
        RECT 14.319 9.744 14.321 12.18 ;
  LAYER M1 ;
        RECT 14.399 9.744 14.401 12.18 ;
  LAYER M1 ;
        RECT 14.479 9.744 14.481 12.18 ;
  LAYER M1 ;
        RECT 14.559 9.744 14.561 12.18 ;
  LAYER M1 ;
        RECT 14.639 9.744 14.641 12.18 ;
  LAYER M1 ;
        RECT 14.719 9.744 14.721 12.18 ;
  LAYER M1 ;
        RECT 14.799 9.744 14.801 12.18 ;
  LAYER M1 ;
        RECT 14.879 9.744 14.881 12.18 ;
  LAYER M1 ;
        RECT 14.959 9.744 14.961 12.18 ;
  LAYER M1 ;
        RECT 15.039 9.744 15.041 12.18 ;
  LAYER M1 ;
        RECT 15.119 9.744 15.121 12.18 ;
  LAYER M1 ;
        RECT 15.199 9.744 15.201 12.18 ;
  LAYER M2 ;
        RECT 12.88 9.743 15.28 9.745 ;
  LAYER M2 ;
        RECT 12.88 9.827 15.28 9.829 ;
  LAYER M2 ;
        RECT 12.88 9.911 15.28 9.913 ;
  LAYER M2 ;
        RECT 12.88 9.995 15.28 9.997 ;
  LAYER M2 ;
        RECT 12.88 10.079 15.28 10.081 ;
  LAYER M2 ;
        RECT 12.88 10.163 15.28 10.165 ;
  LAYER M2 ;
        RECT 12.88 10.247 15.28 10.249 ;
  LAYER M2 ;
        RECT 12.88 10.331 15.28 10.333 ;
  LAYER M2 ;
        RECT 12.88 10.415 15.28 10.417 ;
  LAYER M2 ;
        RECT 12.88 10.499 15.28 10.501 ;
  LAYER M2 ;
        RECT 12.88 10.583 15.28 10.585 ;
  LAYER M2 ;
        RECT 12.88 10.667 15.28 10.669 ;
  LAYER M2 ;
        RECT 12.88 10.7505 15.28 10.7525 ;
  LAYER M2 ;
        RECT 12.88 10.835 15.28 10.837 ;
  LAYER M2 ;
        RECT 12.88 10.919 15.28 10.921 ;
  LAYER M2 ;
        RECT 12.88 11.003 15.28 11.005 ;
  LAYER M2 ;
        RECT 12.88 11.087 15.28 11.089 ;
  LAYER M2 ;
        RECT 12.88 11.171 15.28 11.173 ;
  LAYER M2 ;
        RECT 12.88 11.255 15.28 11.257 ;
  LAYER M2 ;
        RECT 12.88 11.339 15.28 11.341 ;
  LAYER M2 ;
        RECT 12.88 11.423 15.28 11.425 ;
  LAYER M2 ;
        RECT 12.88 11.507 15.28 11.509 ;
  LAYER M2 ;
        RECT 12.88 11.591 15.28 11.593 ;
  LAYER M2 ;
        RECT 12.88 11.675 15.28 11.677 ;
  LAYER M2 ;
        RECT 12.88 11.759 15.28 11.761 ;
  LAYER M2 ;
        RECT 12.88 11.843 15.28 11.845 ;
  LAYER M2 ;
        RECT 12.88 11.927 15.28 11.929 ;
  LAYER M2 ;
        RECT 12.88 12.011 15.28 12.013 ;
  LAYER M2 ;
        RECT 12.88 12.095 15.28 12.097 ;
  LAYER M1 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M1 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M1 ;
        RECT 12.992 12.648 13.024 15.156 ;
  LAYER M1 ;
        RECT 13.056 12.648 13.088 15.156 ;
  LAYER M1 ;
        RECT 13.12 12.648 13.152 15.156 ;
  LAYER M1 ;
        RECT 13.184 12.648 13.216 15.156 ;
  LAYER M1 ;
        RECT 13.248 12.648 13.28 15.156 ;
  LAYER M1 ;
        RECT 13.312 12.648 13.344 15.156 ;
  LAYER M1 ;
        RECT 13.376 12.648 13.408 15.156 ;
  LAYER M1 ;
        RECT 13.44 12.648 13.472 15.156 ;
  LAYER M1 ;
        RECT 13.504 12.648 13.536 15.156 ;
  LAYER M1 ;
        RECT 13.568 12.648 13.6 15.156 ;
  LAYER M1 ;
        RECT 13.632 12.648 13.664 15.156 ;
  LAYER M1 ;
        RECT 13.696 12.648 13.728 15.156 ;
  LAYER M1 ;
        RECT 13.76 12.648 13.792 15.156 ;
  LAYER M1 ;
        RECT 13.824 12.648 13.856 15.156 ;
  LAYER M1 ;
        RECT 13.888 12.648 13.92 15.156 ;
  LAYER M1 ;
        RECT 13.952 12.648 13.984 15.156 ;
  LAYER M1 ;
        RECT 14.016 12.648 14.048 15.156 ;
  LAYER M1 ;
        RECT 14.08 12.648 14.112 15.156 ;
  LAYER M1 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M1 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M1 ;
        RECT 14.272 12.648 14.304 15.156 ;
  LAYER M1 ;
        RECT 14.336 12.648 14.368 15.156 ;
  LAYER M1 ;
        RECT 14.4 12.648 14.432 15.156 ;
  LAYER M1 ;
        RECT 14.464 12.648 14.496 15.156 ;
  LAYER M1 ;
        RECT 14.528 12.648 14.56 15.156 ;
  LAYER M1 ;
        RECT 14.592 12.648 14.624 15.156 ;
  LAYER M1 ;
        RECT 14.656 12.648 14.688 15.156 ;
  LAYER M1 ;
        RECT 14.72 12.648 14.752 15.156 ;
  LAYER M1 ;
        RECT 14.784 12.648 14.816 15.156 ;
  LAYER M1 ;
        RECT 14.848 12.648 14.88 15.156 ;
  LAYER M1 ;
        RECT 14.912 12.648 14.944 15.156 ;
  LAYER M1 ;
        RECT 14.976 12.648 15.008 15.156 ;
  LAYER M1 ;
        RECT 15.04 12.648 15.072 15.156 ;
  LAYER M1 ;
        RECT 15.104 12.648 15.136 15.156 ;
  LAYER M1 ;
        RECT 15.168 12.648 15.2 15.156 ;
  LAYER M2 ;
        RECT 12.844 12.732 15.316 12.764 ;
  LAYER M2 ;
        RECT 12.844 12.796 15.316 12.828 ;
  LAYER M2 ;
        RECT 12.844 12.86 15.316 12.892 ;
  LAYER M2 ;
        RECT 12.844 12.924 15.316 12.956 ;
  LAYER M2 ;
        RECT 12.844 12.988 15.316 13.02 ;
  LAYER M2 ;
        RECT 12.844 13.052 15.316 13.084 ;
  LAYER M2 ;
        RECT 12.844 13.116 15.316 13.148 ;
  LAYER M2 ;
        RECT 12.844 13.18 15.316 13.212 ;
  LAYER M2 ;
        RECT 12.844 13.244 15.316 13.276 ;
  LAYER M2 ;
        RECT 12.844 13.308 15.316 13.34 ;
  LAYER M2 ;
        RECT 12.844 13.372 15.316 13.404 ;
  LAYER M2 ;
        RECT 12.844 13.436 15.316 13.468 ;
  LAYER M2 ;
        RECT 12.844 13.5 15.316 13.532 ;
  LAYER M2 ;
        RECT 12.844 13.564 15.316 13.596 ;
  LAYER M2 ;
        RECT 12.844 13.628 15.316 13.66 ;
  LAYER M2 ;
        RECT 12.844 13.692 15.316 13.724 ;
  LAYER M2 ;
        RECT 12.844 13.756 15.316 13.788 ;
  LAYER M2 ;
        RECT 12.844 13.82 15.316 13.852 ;
  LAYER M2 ;
        RECT 12.844 13.884 15.316 13.916 ;
  LAYER M2 ;
        RECT 12.844 13.948 15.316 13.98 ;
  LAYER M2 ;
        RECT 12.844 14.012 15.316 14.044 ;
  LAYER M2 ;
        RECT 12.844 14.076 15.316 14.108 ;
  LAYER M2 ;
        RECT 12.844 14.14 15.316 14.172 ;
  LAYER M2 ;
        RECT 12.844 14.204 15.316 14.236 ;
  LAYER M2 ;
        RECT 12.844 14.268 15.316 14.3 ;
  LAYER M2 ;
        RECT 12.844 14.332 15.316 14.364 ;
  LAYER M2 ;
        RECT 12.844 14.396 15.316 14.428 ;
  LAYER M2 ;
        RECT 12.844 14.46 15.316 14.492 ;
  LAYER M2 ;
        RECT 12.844 14.524 15.316 14.556 ;
  LAYER M2 ;
        RECT 12.844 14.588 15.316 14.62 ;
  LAYER M2 ;
        RECT 12.844 14.652 15.316 14.684 ;
  LAYER M2 ;
        RECT 12.844 14.716 15.316 14.748 ;
  LAYER M2 ;
        RECT 12.844 14.78 15.316 14.812 ;
  LAYER M2 ;
        RECT 12.844 14.844 15.316 14.876 ;
  LAYER M2 ;
        RECT 12.844 14.908 15.316 14.94 ;
  LAYER M2 ;
        RECT 12.844 14.972 15.316 15.004 ;
  LAYER M3 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M3 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M3 ;
        RECT 12.992 12.648 13.024 15.156 ;
  LAYER M3 ;
        RECT 13.056 12.648 13.088 15.156 ;
  LAYER M3 ;
        RECT 13.12 12.648 13.152 15.156 ;
  LAYER M3 ;
        RECT 13.184 12.648 13.216 15.156 ;
  LAYER M3 ;
        RECT 13.248 12.648 13.28 15.156 ;
  LAYER M3 ;
        RECT 13.312 12.648 13.344 15.156 ;
  LAYER M3 ;
        RECT 13.376 12.648 13.408 15.156 ;
  LAYER M3 ;
        RECT 13.44 12.648 13.472 15.156 ;
  LAYER M3 ;
        RECT 13.504 12.648 13.536 15.156 ;
  LAYER M3 ;
        RECT 13.568 12.648 13.6 15.156 ;
  LAYER M3 ;
        RECT 13.632 12.648 13.664 15.156 ;
  LAYER M3 ;
        RECT 13.696 12.648 13.728 15.156 ;
  LAYER M3 ;
        RECT 13.76 12.648 13.792 15.156 ;
  LAYER M3 ;
        RECT 13.824 12.648 13.856 15.156 ;
  LAYER M3 ;
        RECT 13.888 12.648 13.92 15.156 ;
  LAYER M3 ;
        RECT 13.952 12.648 13.984 15.156 ;
  LAYER M3 ;
        RECT 14.016 12.648 14.048 15.156 ;
  LAYER M3 ;
        RECT 14.08 12.648 14.112 15.156 ;
  LAYER M3 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M3 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M3 ;
        RECT 14.272 12.648 14.304 15.156 ;
  LAYER M3 ;
        RECT 14.336 12.648 14.368 15.156 ;
  LAYER M3 ;
        RECT 14.4 12.648 14.432 15.156 ;
  LAYER M3 ;
        RECT 14.464 12.648 14.496 15.156 ;
  LAYER M3 ;
        RECT 14.528 12.648 14.56 15.156 ;
  LAYER M3 ;
        RECT 14.592 12.648 14.624 15.156 ;
  LAYER M3 ;
        RECT 14.656 12.648 14.688 15.156 ;
  LAYER M3 ;
        RECT 14.72 12.648 14.752 15.156 ;
  LAYER M3 ;
        RECT 14.784 12.648 14.816 15.156 ;
  LAYER M3 ;
        RECT 14.848 12.648 14.88 15.156 ;
  LAYER M3 ;
        RECT 14.912 12.648 14.944 15.156 ;
  LAYER M3 ;
        RECT 14.976 12.648 15.008 15.156 ;
  LAYER M3 ;
        RECT 15.04 12.648 15.072 15.156 ;
  LAYER M3 ;
        RECT 15.104 12.648 15.136 15.156 ;
  LAYER M3 ;
        RECT 15.168 12.648 15.2 15.156 ;
  LAYER M3 ;
        RECT 15.264 12.648 15.296 15.156 ;
  LAYER M1 ;
        RECT 12.879 12.684 12.881 15.12 ;
  LAYER M1 ;
        RECT 12.959 12.684 12.961 15.12 ;
  LAYER M1 ;
        RECT 13.039 12.684 13.041 15.12 ;
  LAYER M1 ;
        RECT 13.119 12.684 13.121 15.12 ;
  LAYER M1 ;
        RECT 13.199 12.684 13.201 15.12 ;
  LAYER M1 ;
        RECT 13.279 12.684 13.281 15.12 ;
  LAYER M1 ;
        RECT 13.359 12.684 13.361 15.12 ;
  LAYER M1 ;
        RECT 13.439 12.684 13.441 15.12 ;
  LAYER M1 ;
        RECT 13.519 12.684 13.521 15.12 ;
  LAYER M1 ;
        RECT 13.599 12.684 13.601 15.12 ;
  LAYER M1 ;
        RECT 13.679 12.684 13.681 15.12 ;
  LAYER M1 ;
        RECT 13.759 12.684 13.761 15.12 ;
  LAYER M1 ;
        RECT 13.839 12.684 13.841 15.12 ;
  LAYER M1 ;
        RECT 13.919 12.684 13.921 15.12 ;
  LAYER M1 ;
        RECT 13.999 12.684 14.001 15.12 ;
  LAYER M1 ;
        RECT 14.079 12.684 14.081 15.12 ;
  LAYER M1 ;
        RECT 14.159 12.684 14.161 15.12 ;
  LAYER M1 ;
        RECT 14.239 12.684 14.241 15.12 ;
  LAYER M1 ;
        RECT 14.319 12.684 14.321 15.12 ;
  LAYER M1 ;
        RECT 14.399 12.684 14.401 15.12 ;
  LAYER M1 ;
        RECT 14.479 12.684 14.481 15.12 ;
  LAYER M1 ;
        RECT 14.559 12.684 14.561 15.12 ;
  LAYER M1 ;
        RECT 14.639 12.684 14.641 15.12 ;
  LAYER M1 ;
        RECT 14.719 12.684 14.721 15.12 ;
  LAYER M1 ;
        RECT 14.799 12.684 14.801 15.12 ;
  LAYER M1 ;
        RECT 14.879 12.684 14.881 15.12 ;
  LAYER M1 ;
        RECT 14.959 12.684 14.961 15.12 ;
  LAYER M1 ;
        RECT 15.039 12.684 15.041 15.12 ;
  LAYER M1 ;
        RECT 15.119 12.684 15.121 15.12 ;
  LAYER M1 ;
        RECT 15.199 12.684 15.201 15.12 ;
  LAYER M2 ;
        RECT 12.88 12.683 15.28 12.685 ;
  LAYER M2 ;
        RECT 12.88 12.767 15.28 12.769 ;
  LAYER M2 ;
        RECT 12.88 12.851 15.28 12.853 ;
  LAYER M2 ;
        RECT 12.88 12.935 15.28 12.937 ;
  LAYER M2 ;
        RECT 12.88 13.019 15.28 13.021 ;
  LAYER M2 ;
        RECT 12.88 13.103 15.28 13.105 ;
  LAYER M2 ;
        RECT 12.88 13.187 15.28 13.189 ;
  LAYER M2 ;
        RECT 12.88 13.271 15.28 13.273 ;
  LAYER M2 ;
        RECT 12.88 13.355 15.28 13.357 ;
  LAYER M2 ;
        RECT 12.88 13.439 15.28 13.441 ;
  LAYER M2 ;
        RECT 12.88 13.523 15.28 13.525 ;
  LAYER M2 ;
        RECT 12.88 13.607 15.28 13.609 ;
  LAYER M2 ;
        RECT 12.88 13.6905 15.28 13.6925 ;
  LAYER M2 ;
        RECT 12.88 13.775 15.28 13.777 ;
  LAYER M2 ;
        RECT 12.88 13.859 15.28 13.861 ;
  LAYER M2 ;
        RECT 12.88 13.943 15.28 13.945 ;
  LAYER M2 ;
        RECT 12.88 14.027 15.28 14.029 ;
  LAYER M2 ;
        RECT 12.88 14.111 15.28 14.113 ;
  LAYER M2 ;
        RECT 12.88 14.195 15.28 14.197 ;
  LAYER M2 ;
        RECT 12.88 14.279 15.28 14.281 ;
  LAYER M2 ;
        RECT 12.88 14.363 15.28 14.365 ;
  LAYER M2 ;
        RECT 12.88 14.447 15.28 14.449 ;
  LAYER M2 ;
        RECT 12.88 14.531 15.28 14.533 ;
  LAYER M2 ;
        RECT 12.88 14.615 15.28 14.617 ;
  LAYER M2 ;
        RECT 12.88 14.699 15.28 14.701 ;
  LAYER M2 ;
        RECT 12.88 14.783 15.28 14.785 ;
  LAYER M2 ;
        RECT 12.88 14.867 15.28 14.869 ;
  LAYER M2 ;
        RECT 12.88 14.951 15.28 14.953 ;
  LAYER M2 ;
        RECT 12.88 15.035 15.28 15.037 ;
  LAYER M1 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M1 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M1 ;
        RECT 12.992 15.588 13.024 18.096 ;
  LAYER M1 ;
        RECT 13.056 15.588 13.088 18.096 ;
  LAYER M1 ;
        RECT 13.12 15.588 13.152 18.096 ;
  LAYER M1 ;
        RECT 13.184 15.588 13.216 18.096 ;
  LAYER M1 ;
        RECT 13.248 15.588 13.28 18.096 ;
  LAYER M1 ;
        RECT 13.312 15.588 13.344 18.096 ;
  LAYER M1 ;
        RECT 13.376 15.588 13.408 18.096 ;
  LAYER M1 ;
        RECT 13.44 15.588 13.472 18.096 ;
  LAYER M1 ;
        RECT 13.504 15.588 13.536 18.096 ;
  LAYER M1 ;
        RECT 13.568 15.588 13.6 18.096 ;
  LAYER M1 ;
        RECT 13.632 15.588 13.664 18.096 ;
  LAYER M1 ;
        RECT 13.696 15.588 13.728 18.096 ;
  LAYER M1 ;
        RECT 13.76 15.588 13.792 18.096 ;
  LAYER M1 ;
        RECT 13.824 15.588 13.856 18.096 ;
  LAYER M1 ;
        RECT 13.888 15.588 13.92 18.096 ;
  LAYER M1 ;
        RECT 13.952 15.588 13.984 18.096 ;
  LAYER M1 ;
        RECT 14.016 15.588 14.048 18.096 ;
  LAYER M1 ;
        RECT 14.08 15.588 14.112 18.096 ;
  LAYER M1 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M1 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M1 ;
        RECT 14.272 15.588 14.304 18.096 ;
  LAYER M1 ;
        RECT 14.336 15.588 14.368 18.096 ;
  LAYER M1 ;
        RECT 14.4 15.588 14.432 18.096 ;
  LAYER M1 ;
        RECT 14.464 15.588 14.496 18.096 ;
  LAYER M1 ;
        RECT 14.528 15.588 14.56 18.096 ;
  LAYER M1 ;
        RECT 14.592 15.588 14.624 18.096 ;
  LAYER M1 ;
        RECT 14.656 15.588 14.688 18.096 ;
  LAYER M1 ;
        RECT 14.72 15.588 14.752 18.096 ;
  LAYER M1 ;
        RECT 14.784 15.588 14.816 18.096 ;
  LAYER M1 ;
        RECT 14.848 15.588 14.88 18.096 ;
  LAYER M1 ;
        RECT 14.912 15.588 14.944 18.096 ;
  LAYER M1 ;
        RECT 14.976 15.588 15.008 18.096 ;
  LAYER M1 ;
        RECT 15.04 15.588 15.072 18.096 ;
  LAYER M1 ;
        RECT 15.104 15.588 15.136 18.096 ;
  LAYER M1 ;
        RECT 15.168 15.588 15.2 18.096 ;
  LAYER M2 ;
        RECT 12.844 15.672 15.316 15.704 ;
  LAYER M2 ;
        RECT 12.844 15.736 15.316 15.768 ;
  LAYER M2 ;
        RECT 12.844 15.8 15.316 15.832 ;
  LAYER M2 ;
        RECT 12.844 15.864 15.316 15.896 ;
  LAYER M2 ;
        RECT 12.844 15.928 15.316 15.96 ;
  LAYER M2 ;
        RECT 12.844 15.992 15.316 16.024 ;
  LAYER M2 ;
        RECT 12.844 16.056 15.316 16.088 ;
  LAYER M2 ;
        RECT 12.844 16.12 15.316 16.152 ;
  LAYER M2 ;
        RECT 12.844 16.184 15.316 16.216 ;
  LAYER M2 ;
        RECT 12.844 16.248 15.316 16.28 ;
  LAYER M2 ;
        RECT 12.844 16.312 15.316 16.344 ;
  LAYER M2 ;
        RECT 12.844 16.376 15.316 16.408 ;
  LAYER M2 ;
        RECT 12.844 16.44 15.316 16.472 ;
  LAYER M2 ;
        RECT 12.844 16.504 15.316 16.536 ;
  LAYER M2 ;
        RECT 12.844 16.568 15.316 16.6 ;
  LAYER M2 ;
        RECT 12.844 16.632 15.316 16.664 ;
  LAYER M2 ;
        RECT 12.844 16.696 15.316 16.728 ;
  LAYER M2 ;
        RECT 12.844 16.76 15.316 16.792 ;
  LAYER M2 ;
        RECT 12.844 16.824 15.316 16.856 ;
  LAYER M2 ;
        RECT 12.844 16.888 15.316 16.92 ;
  LAYER M2 ;
        RECT 12.844 16.952 15.316 16.984 ;
  LAYER M2 ;
        RECT 12.844 17.016 15.316 17.048 ;
  LAYER M2 ;
        RECT 12.844 17.08 15.316 17.112 ;
  LAYER M2 ;
        RECT 12.844 17.144 15.316 17.176 ;
  LAYER M2 ;
        RECT 12.844 17.208 15.316 17.24 ;
  LAYER M2 ;
        RECT 12.844 17.272 15.316 17.304 ;
  LAYER M2 ;
        RECT 12.844 17.336 15.316 17.368 ;
  LAYER M2 ;
        RECT 12.844 17.4 15.316 17.432 ;
  LAYER M2 ;
        RECT 12.844 17.464 15.316 17.496 ;
  LAYER M2 ;
        RECT 12.844 17.528 15.316 17.56 ;
  LAYER M2 ;
        RECT 12.844 17.592 15.316 17.624 ;
  LAYER M2 ;
        RECT 12.844 17.656 15.316 17.688 ;
  LAYER M2 ;
        RECT 12.844 17.72 15.316 17.752 ;
  LAYER M2 ;
        RECT 12.844 17.784 15.316 17.816 ;
  LAYER M2 ;
        RECT 12.844 17.848 15.316 17.88 ;
  LAYER M2 ;
        RECT 12.844 17.912 15.316 17.944 ;
  LAYER M3 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M3 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M3 ;
        RECT 12.992 15.588 13.024 18.096 ;
  LAYER M3 ;
        RECT 13.056 15.588 13.088 18.096 ;
  LAYER M3 ;
        RECT 13.12 15.588 13.152 18.096 ;
  LAYER M3 ;
        RECT 13.184 15.588 13.216 18.096 ;
  LAYER M3 ;
        RECT 13.248 15.588 13.28 18.096 ;
  LAYER M3 ;
        RECT 13.312 15.588 13.344 18.096 ;
  LAYER M3 ;
        RECT 13.376 15.588 13.408 18.096 ;
  LAYER M3 ;
        RECT 13.44 15.588 13.472 18.096 ;
  LAYER M3 ;
        RECT 13.504 15.588 13.536 18.096 ;
  LAYER M3 ;
        RECT 13.568 15.588 13.6 18.096 ;
  LAYER M3 ;
        RECT 13.632 15.588 13.664 18.096 ;
  LAYER M3 ;
        RECT 13.696 15.588 13.728 18.096 ;
  LAYER M3 ;
        RECT 13.76 15.588 13.792 18.096 ;
  LAYER M3 ;
        RECT 13.824 15.588 13.856 18.096 ;
  LAYER M3 ;
        RECT 13.888 15.588 13.92 18.096 ;
  LAYER M3 ;
        RECT 13.952 15.588 13.984 18.096 ;
  LAYER M3 ;
        RECT 14.016 15.588 14.048 18.096 ;
  LAYER M3 ;
        RECT 14.08 15.588 14.112 18.096 ;
  LAYER M3 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M3 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M3 ;
        RECT 14.272 15.588 14.304 18.096 ;
  LAYER M3 ;
        RECT 14.336 15.588 14.368 18.096 ;
  LAYER M3 ;
        RECT 14.4 15.588 14.432 18.096 ;
  LAYER M3 ;
        RECT 14.464 15.588 14.496 18.096 ;
  LAYER M3 ;
        RECT 14.528 15.588 14.56 18.096 ;
  LAYER M3 ;
        RECT 14.592 15.588 14.624 18.096 ;
  LAYER M3 ;
        RECT 14.656 15.588 14.688 18.096 ;
  LAYER M3 ;
        RECT 14.72 15.588 14.752 18.096 ;
  LAYER M3 ;
        RECT 14.784 15.588 14.816 18.096 ;
  LAYER M3 ;
        RECT 14.848 15.588 14.88 18.096 ;
  LAYER M3 ;
        RECT 14.912 15.588 14.944 18.096 ;
  LAYER M3 ;
        RECT 14.976 15.588 15.008 18.096 ;
  LAYER M3 ;
        RECT 15.04 15.588 15.072 18.096 ;
  LAYER M3 ;
        RECT 15.104 15.588 15.136 18.096 ;
  LAYER M3 ;
        RECT 15.168 15.588 15.2 18.096 ;
  LAYER M3 ;
        RECT 15.264 15.588 15.296 18.096 ;
  LAYER M1 ;
        RECT 12.879 15.624 12.881 18.06 ;
  LAYER M1 ;
        RECT 12.959 15.624 12.961 18.06 ;
  LAYER M1 ;
        RECT 13.039 15.624 13.041 18.06 ;
  LAYER M1 ;
        RECT 13.119 15.624 13.121 18.06 ;
  LAYER M1 ;
        RECT 13.199 15.624 13.201 18.06 ;
  LAYER M1 ;
        RECT 13.279 15.624 13.281 18.06 ;
  LAYER M1 ;
        RECT 13.359 15.624 13.361 18.06 ;
  LAYER M1 ;
        RECT 13.439 15.624 13.441 18.06 ;
  LAYER M1 ;
        RECT 13.519 15.624 13.521 18.06 ;
  LAYER M1 ;
        RECT 13.599 15.624 13.601 18.06 ;
  LAYER M1 ;
        RECT 13.679 15.624 13.681 18.06 ;
  LAYER M1 ;
        RECT 13.759 15.624 13.761 18.06 ;
  LAYER M1 ;
        RECT 13.839 15.624 13.841 18.06 ;
  LAYER M1 ;
        RECT 13.919 15.624 13.921 18.06 ;
  LAYER M1 ;
        RECT 13.999 15.624 14.001 18.06 ;
  LAYER M1 ;
        RECT 14.079 15.624 14.081 18.06 ;
  LAYER M1 ;
        RECT 14.159 15.624 14.161 18.06 ;
  LAYER M1 ;
        RECT 14.239 15.624 14.241 18.06 ;
  LAYER M1 ;
        RECT 14.319 15.624 14.321 18.06 ;
  LAYER M1 ;
        RECT 14.399 15.624 14.401 18.06 ;
  LAYER M1 ;
        RECT 14.479 15.624 14.481 18.06 ;
  LAYER M1 ;
        RECT 14.559 15.624 14.561 18.06 ;
  LAYER M1 ;
        RECT 14.639 15.624 14.641 18.06 ;
  LAYER M1 ;
        RECT 14.719 15.624 14.721 18.06 ;
  LAYER M1 ;
        RECT 14.799 15.624 14.801 18.06 ;
  LAYER M1 ;
        RECT 14.879 15.624 14.881 18.06 ;
  LAYER M1 ;
        RECT 14.959 15.624 14.961 18.06 ;
  LAYER M1 ;
        RECT 15.039 15.624 15.041 18.06 ;
  LAYER M1 ;
        RECT 15.119 15.624 15.121 18.06 ;
  LAYER M1 ;
        RECT 15.199 15.624 15.201 18.06 ;
  LAYER M2 ;
        RECT 12.88 15.623 15.28 15.625 ;
  LAYER M2 ;
        RECT 12.88 15.707 15.28 15.709 ;
  LAYER M2 ;
        RECT 12.88 15.791 15.28 15.793 ;
  LAYER M2 ;
        RECT 12.88 15.875 15.28 15.877 ;
  LAYER M2 ;
        RECT 12.88 15.959 15.28 15.961 ;
  LAYER M2 ;
        RECT 12.88 16.043 15.28 16.045 ;
  LAYER M2 ;
        RECT 12.88 16.127 15.28 16.129 ;
  LAYER M2 ;
        RECT 12.88 16.211 15.28 16.213 ;
  LAYER M2 ;
        RECT 12.88 16.295 15.28 16.297 ;
  LAYER M2 ;
        RECT 12.88 16.379 15.28 16.381 ;
  LAYER M2 ;
        RECT 12.88 16.463 15.28 16.465 ;
  LAYER M2 ;
        RECT 12.88 16.547 15.28 16.549 ;
  LAYER M2 ;
        RECT 12.88 16.6305 15.28 16.6325 ;
  LAYER M2 ;
        RECT 12.88 16.715 15.28 16.717 ;
  LAYER M2 ;
        RECT 12.88 16.799 15.28 16.801 ;
  LAYER M2 ;
        RECT 12.88 16.883 15.28 16.885 ;
  LAYER M2 ;
        RECT 12.88 16.967 15.28 16.969 ;
  LAYER M2 ;
        RECT 12.88 17.051 15.28 17.053 ;
  LAYER M2 ;
        RECT 12.88 17.135 15.28 17.137 ;
  LAYER M2 ;
        RECT 12.88 17.219 15.28 17.221 ;
  LAYER M2 ;
        RECT 12.88 17.303 15.28 17.305 ;
  LAYER M2 ;
        RECT 12.88 17.387 15.28 17.389 ;
  LAYER M2 ;
        RECT 12.88 17.471 15.28 17.473 ;
  LAYER M2 ;
        RECT 12.88 17.555 15.28 17.557 ;
  LAYER M2 ;
        RECT 12.88 17.639 15.28 17.641 ;
  LAYER M2 ;
        RECT 12.88 17.723 15.28 17.725 ;
  LAYER M2 ;
        RECT 12.88 17.807 15.28 17.809 ;
  LAYER M2 ;
        RECT 12.88 17.891 15.28 17.893 ;
  LAYER M2 ;
        RECT 12.88 17.975 15.28 17.977 ;
  LAYER M1 ;
        RECT 12.864 18.528 12.896 21.036 ;
  LAYER M1 ;
        RECT 12.928 18.528 12.96 21.036 ;
  LAYER M1 ;
        RECT 12.992 18.528 13.024 21.036 ;
  LAYER M1 ;
        RECT 13.056 18.528 13.088 21.036 ;
  LAYER M1 ;
        RECT 13.12 18.528 13.152 21.036 ;
  LAYER M1 ;
        RECT 13.184 18.528 13.216 21.036 ;
  LAYER M1 ;
        RECT 13.248 18.528 13.28 21.036 ;
  LAYER M1 ;
        RECT 13.312 18.528 13.344 21.036 ;
  LAYER M1 ;
        RECT 13.376 18.528 13.408 21.036 ;
  LAYER M1 ;
        RECT 13.44 18.528 13.472 21.036 ;
  LAYER M1 ;
        RECT 13.504 18.528 13.536 21.036 ;
  LAYER M1 ;
        RECT 13.568 18.528 13.6 21.036 ;
  LAYER M1 ;
        RECT 13.632 18.528 13.664 21.036 ;
  LAYER M1 ;
        RECT 13.696 18.528 13.728 21.036 ;
  LAYER M1 ;
        RECT 13.76 18.528 13.792 21.036 ;
  LAYER M1 ;
        RECT 13.824 18.528 13.856 21.036 ;
  LAYER M1 ;
        RECT 13.888 18.528 13.92 21.036 ;
  LAYER M1 ;
        RECT 13.952 18.528 13.984 21.036 ;
  LAYER M1 ;
        RECT 14.016 18.528 14.048 21.036 ;
  LAYER M1 ;
        RECT 14.08 18.528 14.112 21.036 ;
  LAYER M1 ;
        RECT 14.144 18.528 14.176 21.036 ;
  LAYER M1 ;
        RECT 14.208 18.528 14.24 21.036 ;
  LAYER M1 ;
        RECT 14.272 18.528 14.304 21.036 ;
  LAYER M1 ;
        RECT 14.336 18.528 14.368 21.036 ;
  LAYER M1 ;
        RECT 14.4 18.528 14.432 21.036 ;
  LAYER M1 ;
        RECT 14.464 18.528 14.496 21.036 ;
  LAYER M1 ;
        RECT 14.528 18.528 14.56 21.036 ;
  LAYER M1 ;
        RECT 14.592 18.528 14.624 21.036 ;
  LAYER M1 ;
        RECT 14.656 18.528 14.688 21.036 ;
  LAYER M1 ;
        RECT 14.72 18.528 14.752 21.036 ;
  LAYER M1 ;
        RECT 14.784 18.528 14.816 21.036 ;
  LAYER M1 ;
        RECT 14.848 18.528 14.88 21.036 ;
  LAYER M1 ;
        RECT 14.912 18.528 14.944 21.036 ;
  LAYER M1 ;
        RECT 14.976 18.528 15.008 21.036 ;
  LAYER M1 ;
        RECT 15.04 18.528 15.072 21.036 ;
  LAYER M1 ;
        RECT 15.104 18.528 15.136 21.036 ;
  LAYER M1 ;
        RECT 15.168 18.528 15.2 21.036 ;
  LAYER M2 ;
        RECT 12.844 18.612 15.316 18.644 ;
  LAYER M2 ;
        RECT 12.844 18.676 15.316 18.708 ;
  LAYER M2 ;
        RECT 12.844 18.74 15.316 18.772 ;
  LAYER M2 ;
        RECT 12.844 18.804 15.316 18.836 ;
  LAYER M2 ;
        RECT 12.844 18.868 15.316 18.9 ;
  LAYER M2 ;
        RECT 12.844 18.932 15.316 18.964 ;
  LAYER M2 ;
        RECT 12.844 18.996 15.316 19.028 ;
  LAYER M2 ;
        RECT 12.844 19.06 15.316 19.092 ;
  LAYER M2 ;
        RECT 12.844 19.124 15.316 19.156 ;
  LAYER M2 ;
        RECT 12.844 19.188 15.316 19.22 ;
  LAYER M2 ;
        RECT 12.844 19.252 15.316 19.284 ;
  LAYER M2 ;
        RECT 12.844 19.316 15.316 19.348 ;
  LAYER M2 ;
        RECT 12.844 19.38 15.316 19.412 ;
  LAYER M2 ;
        RECT 12.844 19.444 15.316 19.476 ;
  LAYER M2 ;
        RECT 12.844 19.508 15.316 19.54 ;
  LAYER M2 ;
        RECT 12.844 19.572 15.316 19.604 ;
  LAYER M2 ;
        RECT 12.844 19.636 15.316 19.668 ;
  LAYER M2 ;
        RECT 12.844 19.7 15.316 19.732 ;
  LAYER M2 ;
        RECT 12.844 19.764 15.316 19.796 ;
  LAYER M2 ;
        RECT 12.844 19.828 15.316 19.86 ;
  LAYER M2 ;
        RECT 12.844 19.892 15.316 19.924 ;
  LAYER M2 ;
        RECT 12.844 19.956 15.316 19.988 ;
  LAYER M2 ;
        RECT 12.844 20.02 15.316 20.052 ;
  LAYER M2 ;
        RECT 12.844 20.084 15.316 20.116 ;
  LAYER M2 ;
        RECT 12.844 20.148 15.316 20.18 ;
  LAYER M2 ;
        RECT 12.844 20.212 15.316 20.244 ;
  LAYER M2 ;
        RECT 12.844 20.276 15.316 20.308 ;
  LAYER M2 ;
        RECT 12.844 20.34 15.316 20.372 ;
  LAYER M2 ;
        RECT 12.844 20.404 15.316 20.436 ;
  LAYER M2 ;
        RECT 12.844 20.468 15.316 20.5 ;
  LAYER M2 ;
        RECT 12.844 20.532 15.316 20.564 ;
  LAYER M2 ;
        RECT 12.844 20.596 15.316 20.628 ;
  LAYER M2 ;
        RECT 12.844 20.66 15.316 20.692 ;
  LAYER M2 ;
        RECT 12.844 20.724 15.316 20.756 ;
  LAYER M2 ;
        RECT 12.844 20.788 15.316 20.82 ;
  LAYER M2 ;
        RECT 12.844 20.852 15.316 20.884 ;
  LAYER M3 ;
        RECT 12.864 18.528 12.896 21.036 ;
  LAYER M3 ;
        RECT 12.928 18.528 12.96 21.036 ;
  LAYER M3 ;
        RECT 12.992 18.528 13.024 21.036 ;
  LAYER M3 ;
        RECT 13.056 18.528 13.088 21.036 ;
  LAYER M3 ;
        RECT 13.12 18.528 13.152 21.036 ;
  LAYER M3 ;
        RECT 13.184 18.528 13.216 21.036 ;
  LAYER M3 ;
        RECT 13.248 18.528 13.28 21.036 ;
  LAYER M3 ;
        RECT 13.312 18.528 13.344 21.036 ;
  LAYER M3 ;
        RECT 13.376 18.528 13.408 21.036 ;
  LAYER M3 ;
        RECT 13.44 18.528 13.472 21.036 ;
  LAYER M3 ;
        RECT 13.504 18.528 13.536 21.036 ;
  LAYER M3 ;
        RECT 13.568 18.528 13.6 21.036 ;
  LAYER M3 ;
        RECT 13.632 18.528 13.664 21.036 ;
  LAYER M3 ;
        RECT 13.696 18.528 13.728 21.036 ;
  LAYER M3 ;
        RECT 13.76 18.528 13.792 21.036 ;
  LAYER M3 ;
        RECT 13.824 18.528 13.856 21.036 ;
  LAYER M3 ;
        RECT 13.888 18.528 13.92 21.036 ;
  LAYER M3 ;
        RECT 13.952 18.528 13.984 21.036 ;
  LAYER M3 ;
        RECT 14.016 18.528 14.048 21.036 ;
  LAYER M3 ;
        RECT 14.08 18.528 14.112 21.036 ;
  LAYER M3 ;
        RECT 14.144 18.528 14.176 21.036 ;
  LAYER M3 ;
        RECT 14.208 18.528 14.24 21.036 ;
  LAYER M3 ;
        RECT 14.272 18.528 14.304 21.036 ;
  LAYER M3 ;
        RECT 14.336 18.528 14.368 21.036 ;
  LAYER M3 ;
        RECT 14.4 18.528 14.432 21.036 ;
  LAYER M3 ;
        RECT 14.464 18.528 14.496 21.036 ;
  LAYER M3 ;
        RECT 14.528 18.528 14.56 21.036 ;
  LAYER M3 ;
        RECT 14.592 18.528 14.624 21.036 ;
  LAYER M3 ;
        RECT 14.656 18.528 14.688 21.036 ;
  LAYER M3 ;
        RECT 14.72 18.528 14.752 21.036 ;
  LAYER M3 ;
        RECT 14.784 18.528 14.816 21.036 ;
  LAYER M3 ;
        RECT 14.848 18.528 14.88 21.036 ;
  LAYER M3 ;
        RECT 14.912 18.528 14.944 21.036 ;
  LAYER M3 ;
        RECT 14.976 18.528 15.008 21.036 ;
  LAYER M3 ;
        RECT 15.04 18.528 15.072 21.036 ;
  LAYER M3 ;
        RECT 15.104 18.528 15.136 21.036 ;
  LAYER M3 ;
        RECT 15.168 18.528 15.2 21.036 ;
  LAYER M3 ;
        RECT 15.264 18.528 15.296 21.036 ;
  LAYER M1 ;
        RECT 12.879 18.564 12.881 21 ;
  LAYER M1 ;
        RECT 12.959 18.564 12.961 21 ;
  LAYER M1 ;
        RECT 13.039 18.564 13.041 21 ;
  LAYER M1 ;
        RECT 13.119 18.564 13.121 21 ;
  LAYER M1 ;
        RECT 13.199 18.564 13.201 21 ;
  LAYER M1 ;
        RECT 13.279 18.564 13.281 21 ;
  LAYER M1 ;
        RECT 13.359 18.564 13.361 21 ;
  LAYER M1 ;
        RECT 13.439 18.564 13.441 21 ;
  LAYER M1 ;
        RECT 13.519 18.564 13.521 21 ;
  LAYER M1 ;
        RECT 13.599 18.564 13.601 21 ;
  LAYER M1 ;
        RECT 13.679 18.564 13.681 21 ;
  LAYER M1 ;
        RECT 13.759 18.564 13.761 21 ;
  LAYER M1 ;
        RECT 13.839 18.564 13.841 21 ;
  LAYER M1 ;
        RECT 13.919 18.564 13.921 21 ;
  LAYER M1 ;
        RECT 13.999 18.564 14.001 21 ;
  LAYER M1 ;
        RECT 14.079 18.564 14.081 21 ;
  LAYER M1 ;
        RECT 14.159 18.564 14.161 21 ;
  LAYER M1 ;
        RECT 14.239 18.564 14.241 21 ;
  LAYER M1 ;
        RECT 14.319 18.564 14.321 21 ;
  LAYER M1 ;
        RECT 14.399 18.564 14.401 21 ;
  LAYER M1 ;
        RECT 14.479 18.564 14.481 21 ;
  LAYER M1 ;
        RECT 14.559 18.564 14.561 21 ;
  LAYER M1 ;
        RECT 14.639 18.564 14.641 21 ;
  LAYER M1 ;
        RECT 14.719 18.564 14.721 21 ;
  LAYER M1 ;
        RECT 14.799 18.564 14.801 21 ;
  LAYER M1 ;
        RECT 14.879 18.564 14.881 21 ;
  LAYER M1 ;
        RECT 14.959 18.564 14.961 21 ;
  LAYER M1 ;
        RECT 15.039 18.564 15.041 21 ;
  LAYER M1 ;
        RECT 15.119 18.564 15.121 21 ;
  LAYER M1 ;
        RECT 15.199 18.564 15.201 21 ;
  LAYER M2 ;
        RECT 12.88 18.563 15.28 18.565 ;
  LAYER M2 ;
        RECT 12.88 18.647 15.28 18.649 ;
  LAYER M2 ;
        RECT 12.88 18.731 15.28 18.733 ;
  LAYER M2 ;
        RECT 12.88 18.815 15.28 18.817 ;
  LAYER M2 ;
        RECT 12.88 18.899 15.28 18.901 ;
  LAYER M2 ;
        RECT 12.88 18.983 15.28 18.985 ;
  LAYER M2 ;
        RECT 12.88 19.067 15.28 19.069 ;
  LAYER M2 ;
        RECT 12.88 19.151 15.28 19.153 ;
  LAYER M2 ;
        RECT 12.88 19.235 15.28 19.237 ;
  LAYER M2 ;
        RECT 12.88 19.319 15.28 19.321 ;
  LAYER M2 ;
        RECT 12.88 19.403 15.28 19.405 ;
  LAYER M2 ;
        RECT 12.88 19.487 15.28 19.489 ;
  LAYER M2 ;
        RECT 12.88 19.5705 15.28 19.5725 ;
  LAYER M2 ;
        RECT 12.88 19.655 15.28 19.657 ;
  LAYER M2 ;
        RECT 12.88 19.739 15.28 19.741 ;
  LAYER M2 ;
        RECT 12.88 19.823 15.28 19.825 ;
  LAYER M2 ;
        RECT 12.88 19.907 15.28 19.909 ;
  LAYER M2 ;
        RECT 12.88 19.991 15.28 19.993 ;
  LAYER M2 ;
        RECT 12.88 20.075 15.28 20.077 ;
  LAYER M2 ;
        RECT 12.88 20.159 15.28 20.161 ;
  LAYER M2 ;
        RECT 12.88 20.243 15.28 20.245 ;
  LAYER M2 ;
        RECT 12.88 20.327 15.28 20.329 ;
  LAYER M2 ;
        RECT 12.88 20.411 15.28 20.413 ;
  LAYER M2 ;
        RECT 12.88 20.495 15.28 20.497 ;
  LAYER M2 ;
        RECT 12.88 20.579 15.28 20.581 ;
  LAYER M2 ;
        RECT 12.88 20.663 15.28 20.665 ;
  LAYER M2 ;
        RECT 12.88 20.747 15.28 20.749 ;
  LAYER M2 ;
        RECT 12.88 20.831 15.28 20.833 ;
  LAYER M2 ;
        RECT 12.88 20.915 15.28 20.917 ;
  END 
END Cap_60fF_Cap_60fF
