MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 17.04 BY 19.992 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.78 19.536 6.812 19.608 ;
      LAYER M2 ;
        RECT 6.76 19.556 6.832 19.588 ;
      LAYER M1 ;
        RECT 10.396 19.536 10.428 19.608 ;
      LAYER M2 ;
        RECT 10.376 19.556 10.448 19.588 ;
      LAYER M2 ;
        RECT 6.796 19.556 10.412 19.588 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.3 0.384 6.332 0.456 ;
      LAYER M2 ;
        RECT 6.28 0.404 6.352 0.436 ;
      LAYER M1 ;
        RECT 9.916 0.384 9.948 0.456 ;
      LAYER M2 ;
        RECT 9.896 0.404 9.968 0.436 ;
      LAYER M2 ;
        RECT 6.316 0.404 9.932 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.94 19.704 6.972 19.776 ;
      LAYER M2 ;
        RECT 6.92 19.724 6.992 19.756 ;
      LAYER M1 ;
        RECT 10.556 19.704 10.588 19.776 ;
      LAYER M2 ;
        RECT 10.536 19.724 10.608 19.756 ;
      LAYER M2 ;
        RECT 6.956 19.724 10.572 19.756 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.46 0.216 6.492 0.288 ;
      LAYER M2 ;
        RECT 6.44 0.236 6.512 0.268 ;
      LAYER M1 ;
        RECT 10.076 0.216 10.108 0.288 ;
      LAYER M2 ;
        RECT 10.056 0.236 10.128 0.268 ;
      LAYER M2 ;
        RECT 6.476 0.236 10.092 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 9.692 7.188 9.724 7.26 ;
  LAYER M2 ;
        RECT 9.672 7.208 9.744 7.24 ;
  LAYER M2 ;
        RECT 6.316 7.208 9.708 7.24 ;
  LAYER M1 ;
        RECT 6.3 7.188 6.332 7.26 ;
  LAYER M2 ;
        RECT 6.28 7.208 6.352 7.24 ;
  LAYER M1 ;
        RECT 6.076 13.404 6.108 13.476 ;
  LAYER M2 ;
        RECT 6.056 13.424 6.128 13.456 ;
  LAYER M1 ;
        RECT 6.076 13.272 6.108 13.44 ;
  LAYER M1 ;
        RECT 6.076 13.236 6.108 13.308 ;
  LAYER M2 ;
        RECT 6.056 13.256 6.128 13.288 ;
  LAYER M2 ;
        RECT 6.092 13.256 6.316 13.288 ;
  LAYER M1 ;
        RECT 6.3 13.236 6.332 13.308 ;
  LAYER M2 ;
        RECT 6.28 13.256 6.352 13.288 ;
  LAYER M1 ;
        RECT 6.3 0.384 6.332 0.456 ;
  LAYER M2 ;
        RECT 6.28 0.404 6.352 0.436 ;
  LAYER M1 ;
        RECT 6.3 0.42 6.332 0.672 ;
  LAYER M1 ;
        RECT 6.3 0.672 6.332 13.272 ;
  LAYER M1 ;
        RECT 13.308 4.08 13.34 4.152 ;
  LAYER M2 ;
        RECT 13.288 4.1 13.36 4.132 ;
  LAYER M2 ;
        RECT 9.932 4.1 13.324 4.132 ;
  LAYER M1 ;
        RECT 9.916 4.08 9.948 4.152 ;
  LAYER M2 ;
        RECT 9.896 4.1 9.968 4.132 ;
  LAYER M1 ;
        RECT 9.916 0.384 9.948 0.456 ;
  LAYER M2 ;
        RECT 9.896 0.404 9.968 0.436 ;
  LAYER M1 ;
        RECT 9.916 0.42 9.948 0.672 ;
  LAYER M1 ;
        RECT 9.916 0.672 9.948 4.116 ;
  LAYER M2 ;
        RECT 6.316 0.404 9.932 0.436 ;
  LAYER M1 ;
        RECT 6.076 7.188 6.108 7.26 ;
  LAYER M2 ;
        RECT 6.056 7.208 6.128 7.24 ;
  LAYER M1 ;
        RECT 6.076 7.056 6.108 7.224 ;
  LAYER M1 ;
        RECT 6.076 7.02 6.108 7.092 ;
  LAYER M2 ;
        RECT 6.056 7.04 6.128 7.072 ;
  LAYER M2 ;
        RECT 6.092 7.04 6.476 7.072 ;
  LAYER M1 ;
        RECT 6.46 7.02 6.492 7.092 ;
  LAYER M2 ;
        RECT 6.44 7.04 6.512 7.072 ;
  LAYER M1 ;
        RECT 6.076 10.296 6.108 10.368 ;
  LAYER M2 ;
        RECT 6.056 10.316 6.128 10.348 ;
  LAYER M1 ;
        RECT 6.076 10.164 6.108 10.332 ;
  LAYER M1 ;
        RECT 6.076 10.128 6.108 10.2 ;
  LAYER M2 ;
        RECT 6.056 10.148 6.128 10.18 ;
  LAYER M2 ;
        RECT 6.092 10.148 6.476 10.18 ;
  LAYER M1 ;
        RECT 6.46 10.128 6.492 10.2 ;
  LAYER M2 ;
        RECT 6.44 10.148 6.512 10.18 ;
  LAYER M1 ;
        RECT 9.692 4.08 9.724 4.152 ;
  LAYER M2 ;
        RECT 9.672 4.1 9.744 4.132 ;
  LAYER M2 ;
        RECT 6.476 4.1 9.708 4.132 ;
  LAYER M1 ;
        RECT 6.46 4.08 6.492 4.152 ;
  LAYER M2 ;
        RECT 6.44 4.1 6.512 4.132 ;
  LAYER M1 ;
        RECT 9.692 13.404 9.724 13.476 ;
  LAYER M2 ;
        RECT 9.672 13.424 9.744 13.456 ;
  LAYER M2 ;
        RECT 6.476 13.424 9.708 13.456 ;
  LAYER M1 ;
        RECT 6.46 13.404 6.492 13.476 ;
  LAYER M2 ;
        RECT 6.44 13.424 6.512 13.456 ;
  LAYER M1 ;
        RECT 6.46 0.216 6.492 0.288 ;
  LAYER M2 ;
        RECT 6.44 0.236 6.512 0.268 ;
  LAYER M1 ;
        RECT 6.46 0.252 6.492 0.672 ;
  LAYER M1 ;
        RECT 6.46 0.672 6.492 13.44 ;
  LAYER M1 ;
        RECT 13.308 10.296 13.34 10.368 ;
  LAYER M2 ;
        RECT 13.288 10.316 13.36 10.348 ;
  LAYER M2 ;
        RECT 10.092 10.316 13.324 10.348 ;
  LAYER M1 ;
        RECT 10.076 10.296 10.108 10.368 ;
  LAYER M2 ;
        RECT 10.056 10.316 10.128 10.348 ;
  LAYER M1 ;
        RECT 13.308 7.188 13.34 7.26 ;
  LAYER M2 ;
        RECT 13.288 7.208 13.36 7.24 ;
  LAYER M2 ;
        RECT 10.092 7.208 13.324 7.24 ;
  LAYER M1 ;
        RECT 10.076 7.188 10.108 7.26 ;
  LAYER M2 ;
        RECT 10.056 7.208 10.128 7.24 ;
  LAYER M1 ;
        RECT 10.076 0.216 10.108 0.288 ;
  LAYER M2 ;
        RECT 10.056 0.236 10.128 0.268 ;
  LAYER M1 ;
        RECT 10.076 0.252 10.108 0.672 ;
  LAYER M1 ;
        RECT 10.076 0.672 10.108 10.332 ;
  LAYER M2 ;
        RECT 6.476 0.236 10.092 0.268 ;
  LAYER M1 ;
        RECT 6.076 0.972 6.108 1.044 ;
  LAYER M2 ;
        RECT 6.056 0.992 6.128 1.024 ;
  LAYER M1 ;
        RECT 6.076 0.84 6.108 1.008 ;
  LAYER M1 ;
        RECT 6.076 0.804 6.108 0.876 ;
  LAYER M2 ;
        RECT 6.056 0.824 6.128 0.856 ;
  LAYER M2 ;
        RECT 6.092 0.824 6.636 0.856 ;
  LAYER M1 ;
        RECT 6.62 0.804 6.652 0.876 ;
  LAYER M2 ;
        RECT 6.6 0.824 6.672 0.856 ;
  LAYER M1 ;
        RECT 6.076 4.08 6.108 4.152 ;
  LAYER M2 ;
        RECT 6.056 4.1 6.128 4.132 ;
  LAYER M1 ;
        RECT 6.076 3.948 6.108 4.116 ;
  LAYER M1 ;
        RECT 6.076 3.912 6.108 3.984 ;
  LAYER M2 ;
        RECT 6.056 3.932 6.128 3.964 ;
  LAYER M2 ;
        RECT 6.092 3.932 6.636 3.964 ;
  LAYER M1 ;
        RECT 6.62 3.912 6.652 3.984 ;
  LAYER M2 ;
        RECT 6.6 3.932 6.672 3.964 ;
  LAYER M1 ;
        RECT 6.076 16.512 6.108 16.584 ;
  LAYER M2 ;
        RECT 6.056 16.532 6.128 16.564 ;
  LAYER M1 ;
        RECT 6.076 16.38 6.108 16.548 ;
  LAYER M1 ;
        RECT 6.076 16.344 6.108 16.416 ;
  LAYER M2 ;
        RECT 6.056 16.364 6.128 16.396 ;
  LAYER M2 ;
        RECT 6.092 16.364 6.636 16.396 ;
  LAYER M1 ;
        RECT 6.62 16.344 6.652 16.416 ;
  LAYER M2 ;
        RECT 6.6 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 9.692 0.972 9.724 1.044 ;
  LAYER M2 ;
        RECT 9.672 0.992 9.744 1.024 ;
  LAYER M2 ;
        RECT 6.636 0.992 9.708 1.024 ;
  LAYER M1 ;
        RECT 6.62 0.972 6.652 1.044 ;
  LAYER M2 ;
        RECT 6.6 0.992 6.672 1.024 ;
  LAYER M1 ;
        RECT 9.692 10.296 9.724 10.368 ;
  LAYER M2 ;
        RECT 9.672 10.316 9.744 10.348 ;
  LAYER M2 ;
        RECT 6.636 10.316 9.708 10.348 ;
  LAYER M1 ;
        RECT 6.62 10.296 6.652 10.368 ;
  LAYER M2 ;
        RECT 6.6 10.316 6.672 10.348 ;
  LAYER M1 ;
        RECT 9.692 16.512 9.724 16.584 ;
  LAYER M2 ;
        RECT 9.672 16.532 9.744 16.564 ;
  LAYER M2 ;
        RECT 6.636 16.532 9.708 16.564 ;
  LAYER M1 ;
        RECT 6.62 16.512 6.652 16.584 ;
  LAYER M2 ;
        RECT 6.6 16.532 6.672 16.564 ;
  LAYER M1 ;
        RECT 6.62 0.048 6.652 0.12 ;
  LAYER M2 ;
        RECT 6.6 0.068 6.672 0.1 ;
  LAYER M1 ;
        RECT 6.62 0.084 6.652 0.672 ;
  LAYER M1 ;
        RECT 6.62 0.672 6.652 16.548 ;
  LAYER M1 ;
        RECT 13.308 0.972 13.34 1.044 ;
  LAYER M2 ;
        RECT 13.288 0.992 13.36 1.024 ;
  LAYER M2 ;
        RECT 10.252 0.992 13.324 1.024 ;
  LAYER M1 ;
        RECT 10.236 0.972 10.268 1.044 ;
  LAYER M2 ;
        RECT 10.216 0.992 10.288 1.024 ;
  LAYER M1 ;
        RECT 13.308 13.404 13.34 13.476 ;
  LAYER M2 ;
        RECT 13.288 13.424 13.36 13.456 ;
  LAYER M2 ;
        RECT 10.252 13.424 13.324 13.456 ;
  LAYER M1 ;
        RECT 10.236 13.404 10.268 13.476 ;
  LAYER M2 ;
        RECT 10.216 13.424 10.288 13.456 ;
  LAYER M1 ;
        RECT 13.308 16.512 13.34 16.584 ;
  LAYER M2 ;
        RECT 13.288 16.532 13.36 16.564 ;
  LAYER M2 ;
        RECT 10.252 16.532 13.324 16.564 ;
  LAYER M1 ;
        RECT 10.236 16.512 10.268 16.584 ;
  LAYER M2 ;
        RECT 10.216 16.532 10.288 16.564 ;
  LAYER M1 ;
        RECT 10.236 0.048 10.268 0.12 ;
  LAYER M2 ;
        RECT 10.216 0.068 10.288 0.1 ;
  LAYER M1 ;
        RECT 10.236 0.084 10.268 0.672 ;
  LAYER M1 ;
        RECT 10.236 0.672 10.268 16.548 ;
  LAYER M2 ;
        RECT 6.636 0.068 10.252 0.1 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M2 ;
        RECT 2.476 16.532 6.092 16.564 ;
  LAYER M1 ;
        RECT 6.076 16.512 6.108 16.584 ;
  LAYER M2 ;
        RECT 6.056 16.532 6.128 16.564 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 13.44 2.492 16.548 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 16.584 ;
  LAYER M2 ;
        RECT 2.44 16.532 2.512 16.564 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 10.332 2.492 13.44 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 13.476 ;
  LAYER M2 ;
        RECT 2.44 13.424 2.512 13.456 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 7.224 2.492 10.332 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 10.368 ;
  LAYER M2 ;
        RECT 2.44 10.316 2.512 10.348 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 2.46 4.116 2.492 7.224 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 7.26 ;
  LAYER M2 ;
        RECT 2.44 7.208 2.512 7.24 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 1.044 ;
  LAYER M2 ;
        RECT 2.44 0.992 2.512 1.024 ;
  LAYER M1 ;
        RECT 2.46 1.008 2.492 4.116 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 4.152 ;
  LAYER M2 ;
        RECT 2.44 4.1 2.512 4.132 ;
  LAYER M1 ;
        RECT 16.924 16.512 16.956 16.584 ;
  LAYER M2 ;
        RECT 16.904 16.532 16.976 16.564 ;
  LAYER M2 ;
        RECT 13.324 16.532 16.94 16.564 ;
  LAYER M1 ;
        RECT 13.308 16.512 13.34 16.584 ;
  LAYER M2 ;
        RECT 13.288 16.532 13.36 16.564 ;
  LAYER M1 ;
        RECT 16.924 13.404 16.956 13.476 ;
  LAYER M2 ;
        RECT 16.904 13.424 16.976 13.456 ;
  LAYER M2 ;
        RECT 13.324 13.424 16.94 13.456 ;
  LAYER M1 ;
        RECT 13.308 13.404 13.34 13.476 ;
  LAYER M2 ;
        RECT 13.288 13.424 13.36 13.456 ;
  LAYER M1 ;
        RECT 16.924 10.296 16.956 10.368 ;
  LAYER M2 ;
        RECT 16.904 10.316 16.976 10.348 ;
  LAYER M1 ;
        RECT 16.924 10.332 16.956 13.44 ;
  LAYER M1 ;
        RECT 16.924 13.404 16.956 13.476 ;
  LAYER M2 ;
        RECT 16.904 13.424 16.976 13.456 ;
  LAYER M1 ;
        RECT 16.924 7.188 16.956 7.26 ;
  LAYER M2 ;
        RECT 16.904 7.208 16.976 7.24 ;
  LAYER M1 ;
        RECT 16.924 7.224 16.956 10.332 ;
  LAYER M1 ;
        RECT 16.924 10.296 16.956 10.368 ;
  LAYER M2 ;
        RECT 16.904 10.316 16.976 10.348 ;
  LAYER M1 ;
        RECT 16.924 4.08 16.956 4.152 ;
  LAYER M2 ;
        RECT 16.904 4.1 16.976 4.132 ;
  LAYER M1 ;
        RECT 16.924 4.116 16.956 7.224 ;
  LAYER M1 ;
        RECT 16.924 7.188 16.956 7.26 ;
  LAYER M2 ;
        RECT 16.904 7.208 16.976 7.24 ;
  LAYER M1 ;
        RECT 16.924 0.972 16.956 1.044 ;
  LAYER M2 ;
        RECT 16.904 0.992 16.976 1.024 ;
  LAYER M1 ;
        RECT 16.924 1.008 16.956 4.116 ;
  LAYER M1 ;
        RECT 16.924 4.08 16.956 4.152 ;
  LAYER M2 ;
        RECT 16.904 4.1 16.976 4.132 ;
  LAYER M1 ;
        RECT 7.324 9.624 7.356 9.696 ;
  LAYER M2 ;
        RECT 7.304 9.644 7.376 9.676 ;
  LAYER M2 ;
        RECT 6.796 9.644 7.34 9.676 ;
  LAYER M1 ;
        RECT 6.78 9.624 6.812 9.696 ;
  LAYER M2 ;
        RECT 6.76 9.644 6.832 9.676 ;
  LAYER M1 ;
        RECT 3.708 15.84 3.74 15.912 ;
  LAYER M2 ;
        RECT 3.688 15.86 3.76 15.892 ;
  LAYER M1 ;
        RECT 3.708 15.876 3.74 16.044 ;
  LAYER M1 ;
        RECT 3.708 16.008 3.74 16.08 ;
  LAYER M2 ;
        RECT 3.688 16.028 3.76 16.06 ;
  LAYER M2 ;
        RECT 3.724 16.028 6.796 16.06 ;
  LAYER M1 ;
        RECT 6.78 16.008 6.812 16.08 ;
  LAYER M2 ;
        RECT 6.76 16.028 6.832 16.06 ;
  LAYER M1 ;
        RECT 6.78 19.536 6.812 19.608 ;
  LAYER M2 ;
        RECT 6.76 19.556 6.832 19.588 ;
  LAYER M1 ;
        RECT 6.78 19.32 6.812 19.572 ;
  LAYER M1 ;
        RECT 6.78 9.66 6.812 19.32 ;
  LAYER M1 ;
        RECT 10.94 6.516 10.972 6.588 ;
  LAYER M2 ;
        RECT 10.92 6.536 10.992 6.568 ;
  LAYER M2 ;
        RECT 10.412 6.536 10.956 6.568 ;
  LAYER M1 ;
        RECT 10.396 6.516 10.428 6.588 ;
  LAYER M2 ;
        RECT 10.376 6.536 10.448 6.568 ;
  LAYER M1 ;
        RECT 10.396 19.536 10.428 19.608 ;
  LAYER M2 ;
        RECT 10.376 19.556 10.448 19.588 ;
  LAYER M1 ;
        RECT 10.396 19.32 10.428 19.572 ;
  LAYER M1 ;
        RECT 10.396 6.552 10.428 19.32 ;
  LAYER M2 ;
        RECT 6.796 19.556 10.412 19.588 ;
  LAYER M1 ;
        RECT 3.708 9.624 3.74 9.696 ;
  LAYER M2 ;
        RECT 3.688 9.644 3.76 9.676 ;
  LAYER M1 ;
        RECT 3.708 9.66 3.74 9.828 ;
  LAYER M1 ;
        RECT 3.708 9.792 3.74 9.864 ;
  LAYER M2 ;
        RECT 3.688 9.812 3.76 9.844 ;
  LAYER M2 ;
        RECT 3.724 9.812 6.956 9.844 ;
  LAYER M1 ;
        RECT 6.94 9.792 6.972 9.864 ;
  LAYER M2 ;
        RECT 6.92 9.812 6.992 9.844 ;
  LAYER M1 ;
        RECT 3.708 12.732 3.74 12.804 ;
  LAYER M2 ;
        RECT 3.688 12.752 3.76 12.784 ;
  LAYER M1 ;
        RECT 3.708 12.768 3.74 12.936 ;
  LAYER M1 ;
        RECT 3.708 12.9 3.74 12.972 ;
  LAYER M2 ;
        RECT 3.688 12.92 3.76 12.952 ;
  LAYER M2 ;
        RECT 3.724 12.92 6.956 12.952 ;
  LAYER M1 ;
        RECT 6.94 12.9 6.972 12.972 ;
  LAYER M2 ;
        RECT 6.92 12.92 6.992 12.952 ;
  LAYER M1 ;
        RECT 7.324 6.516 7.356 6.588 ;
  LAYER M2 ;
        RECT 7.304 6.536 7.376 6.568 ;
  LAYER M2 ;
        RECT 6.956 6.536 7.34 6.568 ;
  LAYER M1 ;
        RECT 6.94 6.516 6.972 6.588 ;
  LAYER M2 ;
        RECT 6.92 6.536 6.992 6.568 ;
  LAYER M1 ;
        RECT 7.324 15.84 7.356 15.912 ;
  LAYER M2 ;
        RECT 7.304 15.86 7.376 15.892 ;
  LAYER M2 ;
        RECT 6.956 15.86 7.34 15.892 ;
  LAYER M1 ;
        RECT 6.94 15.84 6.972 15.912 ;
  LAYER M2 ;
        RECT 6.92 15.86 6.992 15.892 ;
  LAYER M1 ;
        RECT 6.94 19.704 6.972 19.776 ;
  LAYER M2 ;
        RECT 6.92 19.724 6.992 19.756 ;
  LAYER M1 ;
        RECT 6.94 19.32 6.972 19.74 ;
  LAYER M1 ;
        RECT 6.94 6.552 6.972 19.32 ;
  LAYER M1 ;
        RECT 10.94 12.732 10.972 12.804 ;
  LAYER M2 ;
        RECT 10.92 12.752 10.992 12.784 ;
  LAYER M2 ;
        RECT 10.572 12.752 10.956 12.784 ;
  LAYER M1 ;
        RECT 10.556 12.732 10.588 12.804 ;
  LAYER M2 ;
        RECT 10.536 12.752 10.608 12.784 ;
  LAYER M1 ;
        RECT 10.94 9.624 10.972 9.696 ;
  LAYER M2 ;
        RECT 10.92 9.644 10.992 9.676 ;
  LAYER M2 ;
        RECT 10.572 9.644 10.956 9.676 ;
  LAYER M1 ;
        RECT 10.556 9.624 10.588 9.696 ;
  LAYER M2 ;
        RECT 10.536 9.644 10.608 9.676 ;
  LAYER M1 ;
        RECT 10.556 19.704 10.588 19.776 ;
  LAYER M2 ;
        RECT 10.536 19.724 10.608 19.756 ;
  LAYER M1 ;
        RECT 10.556 19.32 10.588 19.74 ;
  LAYER M1 ;
        RECT 10.556 9.66 10.588 19.32 ;
  LAYER M2 ;
        RECT 6.956 19.724 10.572 19.756 ;
  LAYER M1 ;
        RECT 3.708 3.408 3.74 3.48 ;
  LAYER M2 ;
        RECT 3.688 3.428 3.76 3.46 ;
  LAYER M1 ;
        RECT 3.708 3.444 3.74 3.612 ;
  LAYER M1 ;
        RECT 3.708 3.576 3.74 3.648 ;
  LAYER M2 ;
        RECT 3.688 3.596 3.76 3.628 ;
  LAYER M2 ;
        RECT 3.724 3.596 7.116 3.628 ;
  LAYER M1 ;
        RECT 7.1 3.576 7.132 3.648 ;
  LAYER M2 ;
        RECT 7.08 3.596 7.152 3.628 ;
  LAYER M1 ;
        RECT 3.708 6.516 3.74 6.588 ;
  LAYER M2 ;
        RECT 3.688 6.536 3.76 6.568 ;
  LAYER M1 ;
        RECT 3.708 6.552 3.74 6.72 ;
  LAYER M1 ;
        RECT 3.708 6.684 3.74 6.756 ;
  LAYER M2 ;
        RECT 3.688 6.704 3.76 6.736 ;
  LAYER M2 ;
        RECT 3.724 6.704 7.116 6.736 ;
  LAYER M1 ;
        RECT 7.1 6.684 7.132 6.756 ;
  LAYER M2 ;
        RECT 7.08 6.704 7.152 6.736 ;
  LAYER M1 ;
        RECT 3.708 18.948 3.74 19.02 ;
  LAYER M2 ;
        RECT 3.688 18.968 3.76 19 ;
  LAYER M1 ;
        RECT 3.708 18.984 3.74 19.152 ;
  LAYER M1 ;
        RECT 3.708 19.116 3.74 19.188 ;
  LAYER M2 ;
        RECT 3.688 19.136 3.76 19.168 ;
  LAYER M2 ;
        RECT 3.724 19.136 7.116 19.168 ;
  LAYER M1 ;
        RECT 7.1 19.116 7.132 19.188 ;
  LAYER M2 ;
        RECT 7.08 19.136 7.152 19.168 ;
  LAYER M1 ;
        RECT 7.324 3.408 7.356 3.48 ;
  LAYER M2 ;
        RECT 7.304 3.428 7.376 3.46 ;
  LAYER M2 ;
        RECT 7.116 3.428 7.34 3.46 ;
  LAYER M1 ;
        RECT 7.1 3.408 7.132 3.48 ;
  LAYER M2 ;
        RECT 7.08 3.428 7.152 3.46 ;
  LAYER M1 ;
        RECT 7.324 12.732 7.356 12.804 ;
  LAYER M2 ;
        RECT 7.304 12.752 7.376 12.784 ;
  LAYER M2 ;
        RECT 7.116 12.752 7.34 12.784 ;
  LAYER M1 ;
        RECT 7.1 12.732 7.132 12.804 ;
  LAYER M2 ;
        RECT 7.08 12.752 7.152 12.784 ;
  LAYER M1 ;
        RECT 7.324 18.948 7.356 19.02 ;
  LAYER M2 ;
        RECT 7.304 18.968 7.376 19 ;
  LAYER M2 ;
        RECT 7.116 18.968 7.34 19 ;
  LAYER M1 ;
        RECT 7.1 18.948 7.132 19.02 ;
  LAYER M2 ;
        RECT 7.08 18.968 7.152 19 ;
  LAYER M1 ;
        RECT 7.1 19.872 7.132 19.944 ;
  LAYER M2 ;
        RECT 7.08 19.892 7.152 19.924 ;
  LAYER M1 ;
        RECT 7.1 19.32 7.132 19.908 ;
  LAYER M1 ;
        RECT 7.1 3.444 7.132 19.32 ;
  LAYER M1 ;
        RECT 10.94 3.408 10.972 3.48 ;
  LAYER M2 ;
        RECT 10.92 3.428 10.992 3.46 ;
  LAYER M2 ;
        RECT 10.732 3.428 10.956 3.46 ;
  LAYER M1 ;
        RECT 10.716 3.408 10.748 3.48 ;
  LAYER M2 ;
        RECT 10.696 3.428 10.768 3.46 ;
  LAYER M1 ;
        RECT 10.94 15.84 10.972 15.912 ;
  LAYER M2 ;
        RECT 10.92 15.86 10.992 15.892 ;
  LAYER M2 ;
        RECT 10.732 15.86 10.956 15.892 ;
  LAYER M1 ;
        RECT 10.716 15.84 10.748 15.912 ;
  LAYER M2 ;
        RECT 10.696 15.86 10.768 15.892 ;
  LAYER M1 ;
        RECT 10.94 18.948 10.972 19.02 ;
  LAYER M2 ;
        RECT 10.92 18.968 10.992 19 ;
  LAYER M2 ;
        RECT 10.732 18.968 10.956 19 ;
  LAYER M1 ;
        RECT 10.716 18.948 10.748 19.02 ;
  LAYER M2 ;
        RECT 10.696 18.968 10.768 19 ;
  LAYER M1 ;
        RECT 10.716 19.872 10.748 19.944 ;
  LAYER M2 ;
        RECT 10.696 19.892 10.768 19.924 ;
  LAYER M1 ;
        RECT 10.716 19.32 10.748 19.908 ;
  LAYER M1 ;
        RECT 10.716 3.444 10.748 19.32 ;
  LAYER M2 ;
        RECT 7.116 19.892 10.732 19.924 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M2 ;
        RECT 0.108 18.968 3.724 19 ;
  LAYER M1 ;
        RECT 3.708 18.948 3.74 19.02 ;
  LAYER M2 ;
        RECT 3.688 18.968 3.76 19 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 15.876 0.124 18.984 ;
  LAYER M1 ;
        RECT 0.092 18.948 0.124 19.02 ;
  LAYER M2 ;
        RECT 0.072 18.968 0.144 19 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 12.768 0.124 15.876 ;
  LAYER M1 ;
        RECT 0.092 15.84 0.124 15.912 ;
  LAYER M2 ;
        RECT 0.072 15.86 0.144 15.892 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 9.66 0.124 12.768 ;
  LAYER M1 ;
        RECT 0.092 12.732 0.124 12.804 ;
  LAYER M2 ;
        RECT 0.072 12.752 0.144 12.784 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 0.092 6.552 0.124 9.66 ;
  LAYER M1 ;
        RECT 0.092 9.624 0.124 9.696 ;
  LAYER M2 ;
        RECT 0.072 9.644 0.144 9.676 ;
  LAYER M1 ;
        RECT 0.092 3.408 0.124 3.48 ;
  LAYER M2 ;
        RECT 0.072 3.428 0.144 3.46 ;
  LAYER M1 ;
        RECT 0.092 3.444 0.124 6.552 ;
  LAYER M1 ;
        RECT 0.092 6.516 0.124 6.588 ;
  LAYER M2 ;
        RECT 0.072 6.536 0.144 6.568 ;
  LAYER M1 ;
        RECT 14.556 18.948 14.588 19.02 ;
  LAYER M2 ;
        RECT 14.536 18.968 14.608 19 ;
  LAYER M2 ;
        RECT 10.956 18.968 14.572 19 ;
  LAYER M1 ;
        RECT 10.94 18.948 10.972 19.02 ;
  LAYER M2 ;
        RECT 10.92 18.968 10.992 19 ;
  LAYER M1 ;
        RECT 14.556 15.84 14.588 15.912 ;
  LAYER M2 ;
        RECT 14.536 15.86 14.608 15.892 ;
  LAYER M2 ;
        RECT 10.956 15.86 14.572 15.892 ;
  LAYER M1 ;
        RECT 10.94 15.84 10.972 15.912 ;
  LAYER M2 ;
        RECT 10.92 15.86 10.992 15.892 ;
  LAYER M1 ;
        RECT 14.556 12.732 14.588 12.804 ;
  LAYER M2 ;
        RECT 14.536 12.752 14.608 12.784 ;
  LAYER M1 ;
        RECT 14.556 12.768 14.588 15.876 ;
  LAYER M1 ;
        RECT 14.556 15.84 14.588 15.912 ;
  LAYER M2 ;
        RECT 14.536 15.86 14.608 15.892 ;
  LAYER M1 ;
        RECT 14.556 9.624 14.588 9.696 ;
  LAYER M2 ;
        RECT 14.536 9.644 14.608 9.676 ;
  LAYER M1 ;
        RECT 14.556 9.66 14.588 12.768 ;
  LAYER M1 ;
        RECT 14.556 12.732 14.588 12.804 ;
  LAYER M2 ;
        RECT 14.536 12.752 14.608 12.784 ;
  LAYER M1 ;
        RECT 14.556 6.516 14.588 6.588 ;
  LAYER M2 ;
        RECT 14.536 6.536 14.608 6.568 ;
  LAYER M1 ;
        RECT 14.556 6.552 14.588 9.66 ;
  LAYER M1 ;
        RECT 14.556 9.624 14.588 9.696 ;
  LAYER M2 ;
        RECT 14.536 9.644 14.608 9.676 ;
  LAYER M1 ;
        RECT 14.556 3.408 14.588 3.48 ;
  LAYER M2 ;
        RECT 14.536 3.428 14.608 3.46 ;
  LAYER M1 ;
        RECT 14.556 3.444 14.588 6.552 ;
  LAYER M1 ;
        RECT 14.556 6.516 14.588 6.588 ;
  LAYER M2 ;
        RECT 14.536 6.536 14.608 6.568 ;
  LAYER M1 ;
        RECT 0.092 0.972 0.124 3.48 ;
  LAYER M3 ;
        RECT 0.092 3.428 0.124 3.46 ;
  LAYER M1 ;
        RECT 0.156 0.972 0.188 3.48 ;
  LAYER M3 ;
        RECT 0.156 0.992 0.188 1.024 ;
  LAYER M1 ;
        RECT 0.22 0.972 0.252 3.48 ;
  LAYER M3 ;
        RECT 0.22 3.428 0.252 3.46 ;
  LAYER M1 ;
        RECT 0.284 0.972 0.316 3.48 ;
  LAYER M3 ;
        RECT 0.284 0.992 0.316 1.024 ;
  LAYER M1 ;
        RECT 0.348 0.972 0.38 3.48 ;
  LAYER M3 ;
        RECT 0.348 3.428 0.38 3.46 ;
  LAYER M1 ;
        RECT 0.412 0.972 0.444 3.48 ;
  LAYER M3 ;
        RECT 0.412 0.992 0.444 1.024 ;
  LAYER M1 ;
        RECT 0.476 0.972 0.508 3.48 ;
  LAYER M3 ;
        RECT 0.476 3.428 0.508 3.46 ;
  LAYER M1 ;
        RECT 0.54 0.972 0.572 3.48 ;
  LAYER M3 ;
        RECT 0.54 0.992 0.572 1.024 ;
  LAYER M1 ;
        RECT 0.604 0.972 0.636 3.48 ;
  LAYER M3 ;
        RECT 0.604 3.428 0.636 3.46 ;
  LAYER M1 ;
        RECT 0.668 0.972 0.7 3.48 ;
  LAYER M3 ;
        RECT 0.668 0.992 0.7 1.024 ;
  LAYER M1 ;
        RECT 0.732 0.972 0.764 3.48 ;
  LAYER M3 ;
        RECT 0.732 3.428 0.764 3.46 ;
  LAYER M1 ;
        RECT 0.796 0.972 0.828 3.48 ;
  LAYER M3 ;
        RECT 0.796 0.992 0.828 1.024 ;
  LAYER M1 ;
        RECT 0.86 0.972 0.892 3.48 ;
  LAYER M3 ;
        RECT 0.86 3.428 0.892 3.46 ;
  LAYER M1 ;
        RECT 0.924 0.972 0.956 3.48 ;
  LAYER M3 ;
        RECT 0.924 0.992 0.956 1.024 ;
  LAYER M1 ;
        RECT 0.988 0.972 1.02 3.48 ;
  LAYER M3 ;
        RECT 0.988 3.428 1.02 3.46 ;
  LAYER M1 ;
        RECT 1.052 0.972 1.084 3.48 ;
  LAYER M3 ;
        RECT 1.052 0.992 1.084 1.024 ;
  LAYER M1 ;
        RECT 1.116 0.972 1.148 3.48 ;
  LAYER M3 ;
        RECT 1.116 3.428 1.148 3.46 ;
  LAYER M1 ;
        RECT 1.18 0.972 1.212 3.48 ;
  LAYER M3 ;
        RECT 1.18 0.992 1.212 1.024 ;
  LAYER M1 ;
        RECT 1.244 0.972 1.276 3.48 ;
  LAYER M3 ;
        RECT 1.244 3.428 1.276 3.46 ;
  LAYER M1 ;
        RECT 1.308 0.972 1.34 3.48 ;
  LAYER M3 ;
        RECT 1.308 0.992 1.34 1.024 ;
  LAYER M1 ;
        RECT 1.372 0.972 1.404 3.48 ;
  LAYER M3 ;
        RECT 1.372 3.428 1.404 3.46 ;
  LAYER M1 ;
        RECT 1.436 0.972 1.468 3.48 ;
  LAYER M3 ;
        RECT 1.436 0.992 1.468 1.024 ;
  LAYER M1 ;
        RECT 1.5 0.972 1.532 3.48 ;
  LAYER M3 ;
        RECT 1.5 3.428 1.532 3.46 ;
  LAYER M1 ;
        RECT 1.564 0.972 1.596 3.48 ;
  LAYER M3 ;
        RECT 1.564 0.992 1.596 1.024 ;
  LAYER M1 ;
        RECT 1.628 0.972 1.66 3.48 ;
  LAYER M3 ;
        RECT 1.628 3.428 1.66 3.46 ;
  LAYER M1 ;
        RECT 1.692 0.972 1.724 3.48 ;
  LAYER M3 ;
        RECT 1.692 0.992 1.724 1.024 ;
  LAYER M1 ;
        RECT 1.756 0.972 1.788 3.48 ;
  LAYER M3 ;
        RECT 1.756 3.428 1.788 3.46 ;
  LAYER M1 ;
        RECT 1.82 0.972 1.852 3.48 ;
  LAYER M3 ;
        RECT 1.82 0.992 1.852 1.024 ;
  LAYER M1 ;
        RECT 1.884 0.972 1.916 3.48 ;
  LAYER M3 ;
        RECT 1.884 3.428 1.916 3.46 ;
  LAYER M1 ;
        RECT 1.948 0.972 1.98 3.48 ;
  LAYER M3 ;
        RECT 1.948 0.992 1.98 1.024 ;
  LAYER M1 ;
        RECT 2.012 0.972 2.044 3.48 ;
  LAYER M3 ;
        RECT 2.012 3.428 2.044 3.46 ;
  LAYER M1 ;
        RECT 2.076 0.972 2.108 3.48 ;
  LAYER M3 ;
        RECT 2.076 0.992 2.108 1.024 ;
  LAYER M1 ;
        RECT 2.14 0.972 2.172 3.48 ;
  LAYER M3 ;
        RECT 2.14 3.428 2.172 3.46 ;
  LAYER M1 ;
        RECT 2.204 0.972 2.236 3.48 ;
  LAYER M3 ;
        RECT 2.204 0.992 2.236 1.024 ;
  LAYER M1 ;
        RECT 2.268 0.972 2.3 3.48 ;
  LAYER M3 ;
        RECT 2.268 3.428 2.3 3.46 ;
  LAYER M1 ;
        RECT 2.332 0.972 2.364 3.48 ;
  LAYER M3 ;
        RECT 2.332 0.992 2.364 1.024 ;
  LAYER M1 ;
        RECT 2.396 0.972 2.428 3.48 ;
  LAYER M3 ;
        RECT 2.396 3.428 2.428 3.46 ;
  LAYER M1 ;
        RECT 2.46 0.972 2.492 3.48 ;
  LAYER M3 ;
        RECT 0.092 1.056 0.124 1.088 ;
  LAYER M2 ;
        RECT 2.46 1.12 2.492 1.152 ;
  LAYER M2 ;
        RECT 0.092 1.184 0.124 1.216 ;
  LAYER M2 ;
        RECT 2.46 1.248 2.492 1.28 ;
  LAYER M2 ;
        RECT 0.092 1.312 0.124 1.344 ;
  LAYER M2 ;
        RECT 2.46 1.376 2.492 1.408 ;
  LAYER M2 ;
        RECT 0.092 1.44 0.124 1.472 ;
  LAYER M2 ;
        RECT 2.46 1.504 2.492 1.536 ;
  LAYER M2 ;
        RECT 0.092 1.568 0.124 1.6 ;
  LAYER M2 ;
        RECT 2.46 1.632 2.492 1.664 ;
  LAYER M2 ;
        RECT 0.092 1.696 0.124 1.728 ;
  LAYER M2 ;
        RECT 2.46 1.76 2.492 1.792 ;
  LAYER M2 ;
        RECT 0.092 1.824 0.124 1.856 ;
  LAYER M2 ;
        RECT 2.46 1.888 2.492 1.92 ;
  LAYER M2 ;
        RECT 0.092 1.952 0.124 1.984 ;
  LAYER M2 ;
        RECT 2.46 2.016 2.492 2.048 ;
  LAYER M2 ;
        RECT 0.092 2.08 0.124 2.112 ;
  LAYER M2 ;
        RECT 2.46 2.144 2.492 2.176 ;
  LAYER M2 ;
        RECT 0.092 2.208 0.124 2.24 ;
  LAYER M2 ;
        RECT 2.46 2.272 2.492 2.304 ;
  LAYER M2 ;
        RECT 0.092 2.336 0.124 2.368 ;
  LAYER M2 ;
        RECT 2.46 2.4 2.492 2.432 ;
  LAYER M2 ;
        RECT 0.092 2.464 0.124 2.496 ;
  LAYER M2 ;
        RECT 2.46 2.528 2.492 2.56 ;
  LAYER M2 ;
        RECT 0.092 2.592 0.124 2.624 ;
  LAYER M2 ;
        RECT 2.46 2.656 2.492 2.688 ;
  LAYER M2 ;
        RECT 0.092 2.72 0.124 2.752 ;
  LAYER M2 ;
        RECT 2.46 2.784 2.492 2.816 ;
  LAYER M2 ;
        RECT 0.092 2.848 0.124 2.88 ;
  LAYER M2 ;
        RECT 2.46 2.912 2.492 2.944 ;
  LAYER M2 ;
        RECT 0.092 2.976 0.124 3.008 ;
  LAYER M2 ;
        RECT 2.46 3.04 2.492 3.072 ;
  LAYER M2 ;
        RECT 0.092 3.104 0.124 3.136 ;
  LAYER M2 ;
        RECT 2.46 3.168 2.492 3.2 ;
  LAYER M2 ;
        RECT 0.092 3.232 0.124 3.264 ;
  LAYER M2 ;
        RECT 2.46 3.296 2.492 3.328 ;
  LAYER M2 ;
        RECT 0.044 0.924 2.54 3.528 ;
  LAYER M1 ;
        RECT 0.092 4.08 0.124 6.588 ;
  LAYER M3 ;
        RECT 0.092 6.536 0.124 6.568 ;
  LAYER M1 ;
        RECT 0.156 4.08 0.188 6.588 ;
  LAYER M3 ;
        RECT 0.156 4.1 0.188 4.132 ;
  LAYER M1 ;
        RECT 0.22 4.08 0.252 6.588 ;
  LAYER M3 ;
        RECT 0.22 6.536 0.252 6.568 ;
  LAYER M1 ;
        RECT 0.284 4.08 0.316 6.588 ;
  LAYER M3 ;
        RECT 0.284 4.1 0.316 4.132 ;
  LAYER M1 ;
        RECT 0.348 4.08 0.38 6.588 ;
  LAYER M3 ;
        RECT 0.348 6.536 0.38 6.568 ;
  LAYER M1 ;
        RECT 0.412 4.08 0.444 6.588 ;
  LAYER M3 ;
        RECT 0.412 4.1 0.444 4.132 ;
  LAYER M1 ;
        RECT 0.476 4.08 0.508 6.588 ;
  LAYER M3 ;
        RECT 0.476 6.536 0.508 6.568 ;
  LAYER M1 ;
        RECT 0.54 4.08 0.572 6.588 ;
  LAYER M3 ;
        RECT 0.54 4.1 0.572 4.132 ;
  LAYER M1 ;
        RECT 0.604 4.08 0.636 6.588 ;
  LAYER M3 ;
        RECT 0.604 6.536 0.636 6.568 ;
  LAYER M1 ;
        RECT 0.668 4.08 0.7 6.588 ;
  LAYER M3 ;
        RECT 0.668 4.1 0.7 4.132 ;
  LAYER M1 ;
        RECT 0.732 4.08 0.764 6.588 ;
  LAYER M3 ;
        RECT 0.732 6.536 0.764 6.568 ;
  LAYER M1 ;
        RECT 0.796 4.08 0.828 6.588 ;
  LAYER M3 ;
        RECT 0.796 4.1 0.828 4.132 ;
  LAYER M1 ;
        RECT 0.86 4.08 0.892 6.588 ;
  LAYER M3 ;
        RECT 0.86 6.536 0.892 6.568 ;
  LAYER M1 ;
        RECT 0.924 4.08 0.956 6.588 ;
  LAYER M3 ;
        RECT 0.924 4.1 0.956 4.132 ;
  LAYER M1 ;
        RECT 0.988 4.08 1.02 6.588 ;
  LAYER M3 ;
        RECT 0.988 6.536 1.02 6.568 ;
  LAYER M1 ;
        RECT 1.052 4.08 1.084 6.588 ;
  LAYER M3 ;
        RECT 1.052 4.1 1.084 4.132 ;
  LAYER M1 ;
        RECT 1.116 4.08 1.148 6.588 ;
  LAYER M3 ;
        RECT 1.116 6.536 1.148 6.568 ;
  LAYER M1 ;
        RECT 1.18 4.08 1.212 6.588 ;
  LAYER M3 ;
        RECT 1.18 4.1 1.212 4.132 ;
  LAYER M1 ;
        RECT 1.244 4.08 1.276 6.588 ;
  LAYER M3 ;
        RECT 1.244 6.536 1.276 6.568 ;
  LAYER M1 ;
        RECT 1.308 4.08 1.34 6.588 ;
  LAYER M3 ;
        RECT 1.308 4.1 1.34 4.132 ;
  LAYER M1 ;
        RECT 1.372 4.08 1.404 6.588 ;
  LAYER M3 ;
        RECT 1.372 6.536 1.404 6.568 ;
  LAYER M1 ;
        RECT 1.436 4.08 1.468 6.588 ;
  LAYER M3 ;
        RECT 1.436 4.1 1.468 4.132 ;
  LAYER M1 ;
        RECT 1.5 4.08 1.532 6.588 ;
  LAYER M3 ;
        RECT 1.5 6.536 1.532 6.568 ;
  LAYER M1 ;
        RECT 1.564 4.08 1.596 6.588 ;
  LAYER M3 ;
        RECT 1.564 4.1 1.596 4.132 ;
  LAYER M1 ;
        RECT 1.628 4.08 1.66 6.588 ;
  LAYER M3 ;
        RECT 1.628 6.536 1.66 6.568 ;
  LAYER M1 ;
        RECT 1.692 4.08 1.724 6.588 ;
  LAYER M3 ;
        RECT 1.692 4.1 1.724 4.132 ;
  LAYER M1 ;
        RECT 1.756 4.08 1.788 6.588 ;
  LAYER M3 ;
        RECT 1.756 6.536 1.788 6.568 ;
  LAYER M1 ;
        RECT 1.82 4.08 1.852 6.588 ;
  LAYER M3 ;
        RECT 1.82 4.1 1.852 4.132 ;
  LAYER M1 ;
        RECT 1.884 4.08 1.916 6.588 ;
  LAYER M3 ;
        RECT 1.884 6.536 1.916 6.568 ;
  LAYER M1 ;
        RECT 1.948 4.08 1.98 6.588 ;
  LAYER M3 ;
        RECT 1.948 4.1 1.98 4.132 ;
  LAYER M1 ;
        RECT 2.012 4.08 2.044 6.588 ;
  LAYER M3 ;
        RECT 2.012 6.536 2.044 6.568 ;
  LAYER M1 ;
        RECT 2.076 4.08 2.108 6.588 ;
  LAYER M3 ;
        RECT 2.076 4.1 2.108 4.132 ;
  LAYER M1 ;
        RECT 2.14 4.08 2.172 6.588 ;
  LAYER M3 ;
        RECT 2.14 6.536 2.172 6.568 ;
  LAYER M1 ;
        RECT 2.204 4.08 2.236 6.588 ;
  LAYER M3 ;
        RECT 2.204 4.1 2.236 4.132 ;
  LAYER M1 ;
        RECT 2.268 4.08 2.3 6.588 ;
  LAYER M3 ;
        RECT 2.268 6.536 2.3 6.568 ;
  LAYER M1 ;
        RECT 2.332 4.08 2.364 6.588 ;
  LAYER M3 ;
        RECT 2.332 4.1 2.364 4.132 ;
  LAYER M1 ;
        RECT 2.396 4.08 2.428 6.588 ;
  LAYER M3 ;
        RECT 2.396 6.536 2.428 6.568 ;
  LAYER M1 ;
        RECT 2.46 4.08 2.492 6.588 ;
  LAYER M3 ;
        RECT 0.092 4.164 0.124 4.196 ;
  LAYER M2 ;
        RECT 2.46 4.228 2.492 4.26 ;
  LAYER M2 ;
        RECT 0.092 4.292 0.124 4.324 ;
  LAYER M2 ;
        RECT 2.46 4.356 2.492 4.388 ;
  LAYER M2 ;
        RECT 0.092 4.42 0.124 4.452 ;
  LAYER M2 ;
        RECT 2.46 4.484 2.492 4.516 ;
  LAYER M2 ;
        RECT 0.092 4.548 0.124 4.58 ;
  LAYER M2 ;
        RECT 2.46 4.612 2.492 4.644 ;
  LAYER M2 ;
        RECT 0.092 4.676 0.124 4.708 ;
  LAYER M2 ;
        RECT 2.46 4.74 2.492 4.772 ;
  LAYER M2 ;
        RECT 0.092 4.804 0.124 4.836 ;
  LAYER M2 ;
        RECT 2.46 4.868 2.492 4.9 ;
  LAYER M2 ;
        RECT 0.092 4.932 0.124 4.964 ;
  LAYER M2 ;
        RECT 2.46 4.996 2.492 5.028 ;
  LAYER M2 ;
        RECT 0.092 5.06 0.124 5.092 ;
  LAYER M2 ;
        RECT 2.46 5.124 2.492 5.156 ;
  LAYER M2 ;
        RECT 0.092 5.188 0.124 5.22 ;
  LAYER M2 ;
        RECT 2.46 5.252 2.492 5.284 ;
  LAYER M2 ;
        RECT 0.092 5.316 0.124 5.348 ;
  LAYER M2 ;
        RECT 2.46 5.38 2.492 5.412 ;
  LAYER M2 ;
        RECT 0.092 5.444 0.124 5.476 ;
  LAYER M2 ;
        RECT 2.46 5.508 2.492 5.54 ;
  LAYER M2 ;
        RECT 0.092 5.572 0.124 5.604 ;
  LAYER M2 ;
        RECT 2.46 5.636 2.492 5.668 ;
  LAYER M2 ;
        RECT 0.092 5.7 0.124 5.732 ;
  LAYER M2 ;
        RECT 2.46 5.764 2.492 5.796 ;
  LAYER M2 ;
        RECT 0.092 5.828 0.124 5.86 ;
  LAYER M2 ;
        RECT 2.46 5.892 2.492 5.924 ;
  LAYER M2 ;
        RECT 0.092 5.956 0.124 5.988 ;
  LAYER M2 ;
        RECT 2.46 6.02 2.492 6.052 ;
  LAYER M2 ;
        RECT 0.092 6.084 0.124 6.116 ;
  LAYER M2 ;
        RECT 2.46 6.148 2.492 6.18 ;
  LAYER M2 ;
        RECT 0.092 6.212 0.124 6.244 ;
  LAYER M2 ;
        RECT 2.46 6.276 2.492 6.308 ;
  LAYER M2 ;
        RECT 0.092 6.34 0.124 6.372 ;
  LAYER M2 ;
        RECT 2.46 6.404 2.492 6.436 ;
  LAYER M2 ;
        RECT 0.044 4.032 2.54 6.636 ;
  LAYER M1 ;
        RECT 0.092 7.188 0.124 9.696 ;
  LAYER M3 ;
        RECT 0.092 9.644 0.124 9.676 ;
  LAYER M1 ;
        RECT 0.156 7.188 0.188 9.696 ;
  LAYER M3 ;
        RECT 0.156 7.208 0.188 7.24 ;
  LAYER M1 ;
        RECT 0.22 7.188 0.252 9.696 ;
  LAYER M3 ;
        RECT 0.22 9.644 0.252 9.676 ;
  LAYER M1 ;
        RECT 0.284 7.188 0.316 9.696 ;
  LAYER M3 ;
        RECT 0.284 7.208 0.316 7.24 ;
  LAYER M1 ;
        RECT 0.348 7.188 0.38 9.696 ;
  LAYER M3 ;
        RECT 0.348 9.644 0.38 9.676 ;
  LAYER M1 ;
        RECT 0.412 7.188 0.444 9.696 ;
  LAYER M3 ;
        RECT 0.412 7.208 0.444 7.24 ;
  LAYER M1 ;
        RECT 0.476 7.188 0.508 9.696 ;
  LAYER M3 ;
        RECT 0.476 9.644 0.508 9.676 ;
  LAYER M1 ;
        RECT 0.54 7.188 0.572 9.696 ;
  LAYER M3 ;
        RECT 0.54 7.208 0.572 7.24 ;
  LAYER M1 ;
        RECT 0.604 7.188 0.636 9.696 ;
  LAYER M3 ;
        RECT 0.604 9.644 0.636 9.676 ;
  LAYER M1 ;
        RECT 0.668 7.188 0.7 9.696 ;
  LAYER M3 ;
        RECT 0.668 7.208 0.7 7.24 ;
  LAYER M1 ;
        RECT 0.732 7.188 0.764 9.696 ;
  LAYER M3 ;
        RECT 0.732 9.644 0.764 9.676 ;
  LAYER M1 ;
        RECT 0.796 7.188 0.828 9.696 ;
  LAYER M3 ;
        RECT 0.796 7.208 0.828 7.24 ;
  LAYER M1 ;
        RECT 0.86 7.188 0.892 9.696 ;
  LAYER M3 ;
        RECT 0.86 9.644 0.892 9.676 ;
  LAYER M1 ;
        RECT 0.924 7.188 0.956 9.696 ;
  LAYER M3 ;
        RECT 0.924 7.208 0.956 7.24 ;
  LAYER M1 ;
        RECT 0.988 7.188 1.02 9.696 ;
  LAYER M3 ;
        RECT 0.988 9.644 1.02 9.676 ;
  LAYER M1 ;
        RECT 1.052 7.188 1.084 9.696 ;
  LAYER M3 ;
        RECT 1.052 7.208 1.084 7.24 ;
  LAYER M1 ;
        RECT 1.116 7.188 1.148 9.696 ;
  LAYER M3 ;
        RECT 1.116 9.644 1.148 9.676 ;
  LAYER M1 ;
        RECT 1.18 7.188 1.212 9.696 ;
  LAYER M3 ;
        RECT 1.18 7.208 1.212 7.24 ;
  LAYER M1 ;
        RECT 1.244 7.188 1.276 9.696 ;
  LAYER M3 ;
        RECT 1.244 9.644 1.276 9.676 ;
  LAYER M1 ;
        RECT 1.308 7.188 1.34 9.696 ;
  LAYER M3 ;
        RECT 1.308 7.208 1.34 7.24 ;
  LAYER M1 ;
        RECT 1.372 7.188 1.404 9.696 ;
  LAYER M3 ;
        RECT 1.372 9.644 1.404 9.676 ;
  LAYER M1 ;
        RECT 1.436 7.188 1.468 9.696 ;
  LAYER M3 ;
        RECT 1.436 7.208 1.468 7.24 ;
  LAYER M1 ;
        RECT 1.5 7.188 1.532 9.696 ;
  LAYER M3 ;
        RECT 1.5 9.644 1.532 9.676 ;
  LAYER M1 ;
        RECT 1.564 7.188 1.596 9.696 ;
  LAYER M3 ;
        RECT 1.564 7.208 1.596 7.24 ;
  LAYER M1 ;
        RECT 1.628 7.188 1.66 9.696 ;
  LAYER M3 ;
        RECT 1.628 9.644 1.66 9.676 ;
  LAYER M1 ;
        RECT 1.692 7.188 1.724 9.696 ;
  LAYER M3 ;
        RECT 1.692 7.208 1.724 7.24 ;
  LAYER M1 ;
        RECT 1.756 7.188 1.788 9.696 ;
  LAYER M3 ;
        RECT 1.756 9.644 1.788 9.676 ;
  LAYER M1 ;
        RECT 1.82 7.188 1.852 9.696 ;
  LAYER M3 ;
        RECT 1.82 7.208 1.852 7.24 ;
  LAYER M1 ;
        RECT 1.884 7.188 1.916 9.696 ;
  LAYER M3 ;
        RECT 1.884 9.644 1.916 9.676 ;
  LAYER M1 ;
        RECT 1.948 7.188 1.98 9.696 ;
  LAYER M3 ;
        RECT 1.948 7.208 1.98 7.24 ;
  LAYER M1 ;
        RECT 2.012 7.188 2.044 9.696 ;
  LAYER M3 ;
        RECT 2.012 9.644 2.044 9.676 ;
  LAYER M1 ;
        RECT 2.076 7.188 2.108 9.696 ;
  LAYER M3 ;
        RECT 2.076 7.208 2.108 7.24 ;
  LAYER M1 ;
        RECT 2.14 7.188 2.172 9.696 ;
  LAYER M3 ;
        RECT 2.14 9.644 2.172 9.676 ;
  LAYER M1 ;
        RECT 2.204 7.188 2.236 9.696 ;
  LAYER M3 ;
        RECT 2.204 7.208 2.236 7.24 ;
  LAYER M1 ;
        RECT 2.268 7.188 2.3 9.696 ;
  LAYER M3 ;
        RECT 2.268 9.644 2.3 9.676 ;
  LAYER M1 ;
        RECT 2.332 7.188 2.364 9.696 ;
  LAYER M3 ;
        RECT 2.332 7.208 2.364 7.24 ;
  LAYER M1 ;
        RECT 2.396 7.188 2.428 9.696 ;
  LAYER M3 ;
        RECT 2.396 9.644 2.428 9.676 ;
  LAYER M1 ;
        RECT 2.46 7.188 2.492 9.696 ;
  LAYER M3 ;
        RECT 0.092 7.272 0.124 7.304 ;
  LAYER M2 ;
        RECT 2.46 7.336 2.492 7.368 ;
  LAYER M2 ;
        RECT 0.092 7.4 0.124 7.432 ;
  LAYER M2 ;
        RECT 2.46 7.464 2.492 7.496 ;
  LAYER M2 ;
        RECT 0.092 7.528 0.124 7.56 ;
  LAYER M2 ;
        RECT 2.46 7.592 2.492 7.624 ;
  LAYER M2 ;
        RECT 0.092 7.656 0.124 7.688 ;
  LAYER M2 ;
        RECT 2.46 7.72 2.492 7.752 ;
  LAYER M2 ;
        RECT 0.092 7.784 0.124 7.816 ;
  LAYER M2 ;
        RECT 2.46 7.848 2.492 7.88 ;
  LAYER M2 ;
        RECT 0.092 7.912 0.124 7.944 ;
  LAYER M2 ;
        RECT 2.46 7.976 2.492 8.008 ;
  LAYER M2 ;
        RECT 0.092 8.04 0.124 8.072 ;
  LAYER M2 ;
        RECT 2.46 8.104 2.492 8.136 ;
  LAYER M2 ;
        RECT 0.092 8.168 0.124 8.2 ;
  LAYER M2 ;
        RECT 2.46 8.232 2.492 8.264 ;
  LAYER M2 ;
        RECT 0.092 8.296 0.124 8.328 ;
  LAYER M2 ;
        RECT 2.46 8.36 2.492 8.392 ;
  LAYER M2 ;
        RECT 0.092 8.424 0.124 8.456 ;
  LAYER M2 ;
        RECT 2.46 8.488 2.492 8.52 ;
  LAYER M2 ;
        RECT 0.092 8.552 0.124 8.584 ;
  LAYER M2 ;
        RECT 2.46 8.616 2.492 8.648 ;
  LAYER M2 ;
        RECT 0.092 8.68 0.124 8.712 ;
  LAYER M2 ;
        RECT 2.46 8.744 2.492 8.776 ;
  LAYER M2 ;
        RECT 0.092 8.808 0.124 8.84 ;
  LAYER M2 ;
        RECT 2.46 8.872 2.492 8.904 ;
  LAYER M2 ;
        RECT 0.092 8.936 0.124 8.968 ;
  LAYER M2 ;
        RECT 2.46 9 2.492 9.032 ;
  LAYER M2 ;
        RECT 0.092 9.064 0.124 9.096 ;
  LAYER M2 ;
        RECT 2.46 9.128 2.492 9.16 ;
  LAYER M2 ;
        RECT 0.092 9.192 0.124 9.224 ;
  LAYER M2 ;
        RECT 2.46 9.256 2.492 9.288 ;
  LAYER M2 ;
        RECT 0.092 9.32 0.124 9.352 ;
  LAYER M2 ;
        RECT 2.46 9.384 2.492 9.416 ;
  LAYER M2 ;
        RECT 0.092 9.448 0.124 9.48 ;
  LAYER M2 ;
        RECT 2.46 9.512 2.492 9.544 ;
  LAYER M2 ;
        RECT 0.044 7.14 2.54 9.744 ;
  LAYER M1 ;
        RECT 0.092 10.296 0.124 12.804 ;
  LAYER M3 ;
        RECT 0.092 12.752 0.124 12.784 ;
  LAYER M1 ;
        RECT 0.156 10.296 0.188 12.804 ;
  LAYER M3 ;
        RECT 0.156 10.316 0.188 10.348 ;
  LAYER M1 ;
        RECT 0.22 10.296 0.252 12.804 ;
  LAYER M3 ;
        RECT 0.22 12.752 0.252 12.784 ;
  LAYER M1 ;
        RECT 0.284 10.296 0.316 12.804 ;
  LAYER M3 ;
        RECT 0.284 10.316 0.316 10.348 ;
  LAYER M1 ;
        RECT 0.348 10.296 0.38 12.804 ;
  LAYER M3 ;
        RECT 0.348 12.752 0.38 12.784 ;
  LAYER M1 ;
        RECT 0.412 10.296 0.444 12.804 ;
  LAYER M3 ;
        RECT 0.412 10.316 0.444 10.348 ;
  LAYER M1 ;
        RECT 0.476 10.296 0.508 12.804 ;
  LAYER M3 ;
        RECT 0.476 12.752 0.508 12.784 ;
  LAYER M1 ;
        RECT 0.54 10.296 0.572 12.804 ;
  LAYER M3 ;
        RECT 0.54 10.316 0.572 10.348 ;
  LAYER M1 ;
        RECT 0.604 10.296 0.636 12.804 ;
  LAYER M3 ;
        RECT 0.604 12.752 0.636 12.784 ;
  LAYER M1 ;
        RECT 0.668 10.296 0.7 12.804 ;
  LAYER M3 ;
        RECT 0.668 10.316 0.7 10.348 ;
  LAYER M1 ;
        RECT 0.732 10.296 0.764 12.804 ;
  LAYER M3 ;
        RECT 0.732 12.752 0.764 12.784 ;
  LAYER M1 ;
        RECT 0.796 10.296 0.828 12.804 ;
  LAYER M3 ;
        RECT 0.796 10.316 0.828 10.348 ;
  LAYER M1 ;
        RECT 0.86 10.296 0.892 12.804 ;
  LAYER M3 ;
        RECT 0.86 12.752 0.892 12.784 ;
  LAYER M1 ;
        RECT 0.924 10.296 0.956 12.804 ;
  LAYER M3 ;
        RECT 0.924 10.316 0.956 10.348 ;
  LAYER M1 ;
        RECT 0.988 10.296 1.02 12.804 ;
  LAYER M3 ;
        RECT 0.988 12.752 1.02 12.784 ;
  LAYER M1 ;
        RECT 1.052 10.296 1.084 12.804 ;
  LAYER M3 ;
        RECT 1.052 10.316 1.084 10.348 ;
  LAYER M1 ;
        RECT 1.116 10.296 1.148 12.804 ;
  LAYER M3 ;
        RECT 1.116 12.752 1.148 12.784 ;
  LAYER M1 ;
        RECT 1.18 10.296 1.212 12.804 ;
  LAYER M3 ;
        RECT 1.18 10.316 1.212 10.348 ;
  LAYER M1 ;
        RECT 1.244 10.296 1.276 12.804 ;
  LAYER M3 ;
        RECT 1.244 12.752 1.276 12.784 ;
  LAYER M1 ;
        RECT 1.308 10.296 1.34 12.804 ;
  LAYER M3 ;
        RECT 1.308 10.316 1.34 10.348 ;
  LAYER M1 ;
        RECT 1.372 10.296 1.404 12.804 ;
  LAYER M3 ;
        RECT 1.372 12.752 1.404 12.784 ;
  LAYER M1 ;
        RECT 1.436 10.296 1.468 12.804 ;
  LAYER M3 ;
        RECT 1.436 10.316 1.468 10.348 ;
  LAYER M1 ;
        RECT 1.5 10.296 1.532 12.804 ;
  LAYER M3 ;
        RECT 1.5 12.752 1.532 12.784 ;
  LAYER M1 ;
        RECT 1.564 10.296 1.596 12.804 ;
  LAYER M3 ;
        RECT 1.564 10.316 1.596 10.348 ;
  LAYER M1 ;
        RECT 1.628 10.296 1.66 12.804 ;
  LAYER M3 ;
        RECT 1.628 12.752 1.66 12.784 ;
  LAYER M1 ;
        RECT 1.692 10.296 1.724 12.804 ;
  LAYER M3 ;
        RECT 1.692 10.316 1.724 10.348 ;
  LAYER M1 ;
        RECT 1.756 10.296 1.788 12.804 ;
  LAYER M3 ;
        RECT 1.756 12.752 1.788 12.784 ;
  LAYER M1 ;
        RECT 1.82 10.296 1.852 12.804 ;
  LAYER M3 ;
        RECT 1.82 10.316 1.852 10.348 ;
  LAYER M1 ;
        RECT 1.884 10.296 1.916 12.804 ;
  LAYER M3 ;
        RECT 1.884 12.752 1.916 12.784 ;
  LAYER M1 ;
        RECT 1.948 10.296 1.98 12.804 ;
  LAYER M3 ;
        RECT 1.948 10.316 1.98 10.348 ;
  LAYER M1 ;
        RECT 2.012 10.296 2.044 12.804 ;
  LAYER M3 ;
        RECT 2.012 12.752 2.044 12.784 ;
  LAYER M1 ;
        RECT 2.076 10.296 2.108 12.804 ;
  LAYER M3 ;
        RECT 2.076 10.316 2.108 10.348 ;
  LAYER M1 ;
        RECT 2.14 10.296 2.172 12.804 ;
  LAYER M3 ;
        RECT 2.14 12.752 2.172 12.784 ;
  LAYER M1 ;
        RECT 2.204 10.296 2.236 12.804 ;
  LAYER M3 ;
        RECT 2.204 10.316 2.236 10.348 ;
  LAYER M1 ;
        RECT 2.268 10.296 2.3 12.804 ;
  LAYER M3 ;
        RECT 2.268 12.752 2.3 12.784 ;
  LAYER M1 ;
        RECT 2.332 10.296 2.364 12.804 ;
  LAYER M3 ;
        RECT 2.332 10.316 2.364 10.348 ;
  LAYER M1 ;
        RECT 2.396 10.296 2.428 12.804 ;
  LAYER M3 ;
        RECT 2.396 12.752 2.428 12.784 ;
  LAYER M1 ;
        RECT 2.46 10.296 2.492 12.804 ;
  LAYER M3 ;
        RECT 0.092 10.38 0.124 10.412 ;
  LAYER M2 ;
        RECT 2.46 10.444 2.492 10.476 ;
  LAYER M2 ;
        RECT 0.092 10.508 0.124 10.54 ;
  LAYER M2 ;
        RECT 2.46 10.572 2.492 10.604 ;
  LAYER M2 ;
        RECT 0.092 10.636 0.124 10.668 ;
  LAYER M2 ;
        RECT 2.46 10.7 2.492 10.732 ;
  LAYER M2 ;
        RECT 0.092 10.764 0.124 10.796 ;
  LAYER M2 ;
        RECT 2.46 10.828 2.492 10.86 ;
  LAYER M2 ;
        RECT 0.092 10.892 0.124 10.924 ;
  LAYER M2 ;
        RECT 2.46 10.956 2.492 10.988 ;
  LAYER M2 ;
        RECT 0.092 11.02 0.124 11.052 ;
  LAYER M2 ;
        RECT 2.46 11.084 2.492 11.116 ;
  LAYER M2 ;
        RECT 0.092 11.148 0.124 11.18 ;
  LAYER M2 ;
        RECT 2.46 11.212 2.492 11.244 ;
  LAYER M2 ;
        RECT 0.092 11.276 0.124 11.308 ;
  LAYER M2 ;
        RECT 2.46 11.34 2.492 11.372 ;
  LAYER M2 ;
        RECT 0.092 11.404 0.124 11.436 ;
  LAYER M2 ;
        RECT 2.46 11.468 2.492 11.5 ;
  LAYER M2 ;
        RECT 0.092 11.532 0.124 11.564 ;
  LAYER M2 ;
        RECT 2.46 11.596 2.492 11.628 ;
  LAYER M2 ;
        RECT 0.092 11.66 0.124 11.692 ;
  LAYER M2 ;
        RECT 2.46 11.724 2.492 11.756 ;
  LAYER M2 ;
        RECT 0.092 11.788 0.124 11.82 ;
  LAYER M2 ;
        RECT 2.46 11.852 2.492 11.884 ;
  LAYER M2 ;
        RECT 0.092 11.916 0.124 11.948 ;
  LAYER M2 ;
        RECT 2.46 11.98 2.492 12.012 ;
  LAYER M2 ;
        RECT 0.092 12.044 0.124 12.076 ;
  LAYER M2 ;
        RECT 2.46 12.108 2.492 12.14 ;
  LAYER M2 ;
        RECT 0.092 12.172 0.124 12.204 ;
  LAYER M2 ;
        RECT 2.46 12.236 2.492 12.268 ;
  LAYER M2 ;
        RECT 0.092 12.3 0.124 12.332 ;
  LAYER M2 ;
        RECT 2.46 12.364 2.492 12.396 ;
  LAYER M2 ;
        RECT 0.092 12.428 0.124 12.46 ;
  LAYER M2 ;
        RECT 2.46 12.492 2.492 12.524 ;
  LAYER M2 ;
        RECT 0.092 12.556 0.124 12.588 ;
  LAYER M2 ;
        RECT 2.46 12.62 2.492 12.652 ;
  LAYER M2 ;
        RECT 0.044 10.248 2.54 12.852 ;
  LAYER M1 ;
        RECT 0.092 13.404 0.124 15.912 ;
  LAYER M3 ;
        RECT 0.092 15.86 0.124 15.892 ;
  LAYER M1 ;
        RECT 0.156 13.404 0.188 15.912 ;
  LAYER M3 ;
        RECT 0.156 13.424 0.188 13.456 ;
  LAYER M1 ;
        RECT 0.22 13.404 0.252 15.912 ;
  LAYER M3 ;
        RECT 0.22 15.86 0.252 15.892 ;
  LAYER M1 ;
        RECT 0.284 13.404 0.316 15.912 ;
  LAYER M3 ;
        RECT 0.284 13.424 0.316 13.456 ;
  LAYER M1 ;
        RECT 0.348 13.404 0.38 15.912 ;
  LAYER M3 ;
        RECT 0.348 15.86 0.38 15.892 ;
  LAYER M1 ;
        RECT 0.412 13.404 0.444 15.912 ;
  LAYER M3 ;
        RECT 0.412 13.424 0.444 13.456 ;
  LAYER M1 ;
        RECT 0.476 13.404 0.508 15.912 ;
  LAYER M3 ;
        RECT 0.476 15.86 0.508 15.892 ;
  LAYER M1 ;
        RECT 0.54 13.404 0.572 15.912 ;
  LAYER M3 ;
        RECT 0.54 13.424 0.572 13.456 ;
  LAYER M1 ;
        RECT 0.604 13.404 0.636 15.912 ;
  LAYER M3 ;
        RECT 0.604 15.86 0.636 15.892 ;
  LAYER M1 ;
        RECT 0.668 13.404 0.7 15.912 ;
  LAYER M3 ;
        RECT 0.668 13.424 0.7 13.456 ;
  LAYER M1 ;
        RECT 0.732 13.404 0.764 15.912 ;
  LAYER M3 ;
        RECT 0.732 15.86 0.764 15.892 ;
  LAYER M1 ;
        RECT 0.796 13.404 0.828 15.912 ;
  LAYER M3 ;
        RECT 0.796 13.424 0.828 13.456 ;
  LAYER M1 ;
        RECT 0.86 13.404 0.892 15.912 ;
  LAYER M3 ;
        RECT 0.86 15.86 0.892 15.892 ;
  LAYER M1 ;
        RECT 0.924 13.404 0.956 15.912 ;
  LAYER M3 ;
        RECT 0.924 13.424 0.956 13.456 ;
  LAYER M1 ;
        RECT 0.988 13.404 1.02 15.912 ;
  LAYER M3 ;
        RECT 0.988 15.86 1.02 15.892 ;
  LAYER M1 ;
        RECT 1.052 13.404 1.084 15.912 ;
  LAYER M3 ;
        RECT 1.052 13.424 1.084 13.456 ;
  LAYER M1 ;
        RECT 1.116 13.404 1.148 15.912 ;
  LAYER M3 ;
        RECT 1.116 15.86 1.148 15.892 ;
  LAYER M1 ;
        RECT 1.18 13.404 1.212 15.912 ;
  LAYER M3 ;
        RECT 1.18 13.424 1.212 13.456 ;
  LAYER M1 ;
        RECT 1.244 13.404 1.276 15.912 ;
  LAYER M3 ;
        RECT 1.244 15.86 1.276 15.892 ;
  LAYER M1 ;
        RECT 1.308 13.404 1.34 15.912 ;
  LAYER M3 ;
        RECT 1.308 13.424 1.34 13.456 ;
  LAYER M1 ;
        RECT 1.372 13.404 1.404 15.912 ;
  LAYER M3 ;
        RECT 1.372 15.86 1.404 15.892 ;
  LAYER M1 ;
        RECT 1.436 13.404 1.468 15.912 ;
  LAYER M3 ;
        RECT 1.436 13.424 1.468 13.456 ;
  LAYER M1 ;
        RECT 1.5 13.404 1.532 15.912 ;
  LAYER M3 ;
        RECT 1.5 15.86 1.532 15.892 ;
  LAYER M1 ;
        RECT 1.564 13.404 1.596 15.912 ;
  LAYER M3 ;
        RECT 1.564 13.424 1.596 13.456 ;
  LAYER M1 ;
        RECT 1.628 13.404 1.66 15.912 ;
  LAYER M3 ;
        RECT 1.628 15.86 1.66 15.892 ;
  LAYER M1 ;
        RECT 1.692 13.404 1.724 15.912 ;
  LAYER M3 ;
        RECT 1.692 13.424 1.724 13.456 ;
  LAYER M1 ;
        RECT 1.756 13.404 1.788 15.912 ;
  LAYER M3 ;
        RECT 1.756 15.86 1.788 15.892 ;
  LAYER M1 ;
        RECT 1.82 13.404 1.852 15.912 ;
  LAYER M3 ;
        RECT 1.82 13.424 1.852 13.456 ;
  LAYER M1 ;
        RECT 1.884 13.404 1.916 15.912 ;
  LAYER M3 ;
        RECT 1.884 15.86 1.916 15.892 ;
  LAYER M1 ;
        RECT 1.948 13.404 1.98 15.912 ;
  LAYER M3 ;
        RECT 1.948 13.424 1.98 13.456 ;
  LAYER M1 ;
        RECT 2.012 13.404 2.044 15.912 ;
  LAYER M3 ;
        RECT 2.012 15.86 2.044 15.892 ;
  LAYER M1 ;
        RECT 2.076 13.404 2.108 15.912 ;
  LAYER M3 ;
        RECT 2.076 13.424 2.108 13.456 ;
  LAYER M1 ;
        RECT 2.14 13.404 2.172 15.912 ;
  LAYER M3 ;
        RECT 2.14 15.86 2.172 15.892 ;
  LAYER M1 ;
        RECT 2.204 13.404 2.236 15.912 ;
  LAYER M3 ;
        RECT 2.204 13.424 2.236 13.456 ;
  LAYER M1 ;
        RECT 2.268 13.404 2.3 15.912 ;
  LAYER M3 ;
        RECT 2.268 15.86 2.3 15.892 ;
  LAYER M1 ;
        RECT 2.332 13.404 2.364 15.912 ;
  LAYER M3 ;
        RECT 2.332 13.424 2.364 13.456 ;
  LAYER M1 ;
        RECT 2.396 13.404 2.428 15.912 ;
  LAYER M3 ;
        RECT 2.396 15.86 2.428 15.892 ;
  LAYER M1 ;
        RECT 2.46 13.404 2.492 15.912 ;
  LAYER M3 ;
        RECT 0.092 13.488 0.124 13.52 ;
  LAYER M2 ;
        RECT 2.46 13.552 2.492 13.584 ;
  LAYER M2 ;
        RECT 0.092 13.616 0.124 13.648 ;
  LAYER M2 ;
        RECT 2.46 13.68 2.492 13.712 ;
  LAYER M2 ;
        RECT 0.092 13.744 0.124 13.776 ;
  LAYER M2 ;
        RECT 2.46 13.808 2.492 13.84 ;
  LAYER M2 ;
        RECT 0.092 13.872 0.124 13.904 ;
  LAYER M2 ;
        RECT 2.46 13.936 2.492 13.968 ;
  LAYER M2 ;
        RECT 0.092 14 0.124 14.032 ;
  LAYER M2 ;
        RECT 2.46 14.064 2.492 14.096 ;
  LAYER M2 ;
        RECT 0.092 14.128 0.124 14.16 ;
  LAYER M2 ;
        RECT 2.46 14.192 2.492 14.224 ;
  LAYER M2 ;
        RECT 0.092 14.256 0.124 14.288 ;
  LAYER M2 ;
        RECT 2.46 14.32 2.492 14.352 ;
  LAYER M2 ;
        RECT 0.092 14.384 0.124 14.416 ;
  LAYER M2 ;
        RECT 2.46 14.448 2.492 14.48 ;
  LAYER M2 ;
        RECT 0.092 14.512 0.124 14.544 ;
  LAYER M2 ;
        RECT 2.46 14.576 2.492 14.608 ;
  LAYER M2 ;
        RECT 0.092 14.64 0.124 14.672 ;
  LAYER M2 ;
        RECT 2.46 14.704 2.492 14.736 ;
  LAYER M2 ;
        RECT 0.092 14.768 0.124 14.8 ;
  LAYER M2 ;
        RECT 2.46 14.832 2.492 14.864 ;
  LAYER M2 ;
        RECT 0.092 14.896 0.124 14.928 ;
  LAYER M2 ;
        RECT 2.46 14.96 2.492 14.992 ;
  LAYER M2 ;
        RECT 0.092 15.024 0.124 15.056 ;
  LAYER M2 ;
        RECT 2.46 15.088 2.492 15.12 ;
  LAYER M2 ;
        RECT 0.092 15.152 0.124 15.184 ;
  LAYER M2 ;
        RECT 2.46 15.216 2.492 15.248 ;
  LAYER M2 ;
        RECT 0.092 15.28 0.124 15.312 ;
  LAYER M2 ;
        RECT 2.46 15.344 2.492 15.376 ;
  LAYER M2 ;
        RECT 0.092 15.408 0.124 15.44 ;
  LAYER M2 ;
        RECT 2.46 15.472 2.492 15.504 ;
  LAYER M2 ;
        RECT 0.092 15.536 0.124 15.568 ;
  LAYER M2 ;
        RECT 2.46 15.6 2.492 15.632 ;
  LAYER M2 ;
        RECT 0.092 15.664 0.124 15.696 ;
  LAYER M2 ;
        RECT 2.46 15.728 2.492 15.76 ;
  LAYER M2 ;
        RECT 0.044 13.356 2.54 15.96 ;
  LAYER M1 ;
        RECT 0.092 16.512 0.124 19.02 ;
  LAYER M3 ;
        RECT 0.092 18.968 0.124 19 ;
  LAYER M1 ;
        RECT 0.156 16.512 0.188 19.02 ;
  LAYER M3 ;
        RECT 0.156 16.532 0.188 16.564 ;
  LAYER M1 ;
        RECT 0.22 16.512 0.252 19.02 ;
  LAYER M3 ;
        RECT 0.22 18.968 0.252 19 ;
  LAYER M1 ;
        RECT 0.284 16.512 0.316 19.02 ;
  LAYER M3 ;
        RECT 0.284 16.532 0.316 16.564 ;
  LAYER M1 ;
        RECT 0.348 16.512 0.38 19.02 ;
  LAYER M3 ;
        RECT 0.348 18.968 0.38 19 ;
  LAYER M1 ;
        RECT 0.412 16.512 0.444 19.02 ;
  LAYER M3 ;
        RECT 0.412 16.532 0.444 16.564 ;
  LAYER M1 ;
        RECT 0.476 16.512 0.508 19.02 ;
  LAYER M3 ;
        RECT 0.476 18.968 0.508 19 ;
  LAYER M1 ;
        RECT 0.54 16.512 0.572 19.02 ;
  LAYER M3 ;
        RECT 0.54 16.532 0.572 16.564 ;
  LAYER M1 ;
        RECT 0.604 16.512 0.636 19.02 ;
  LAYER M3 ;
        RECT 0.604 18.968 0.636 19 ;
  LAYER M1 ;
        RECT 0.668 16.512 0.7 19.02 ;
  LAYER M3 ;
        RECT 0.668 16.532 0.7 16.564 ;
  LAYER M1 ;
        RECT 0.732 16.512 0.764 19.02 ;
  LAYER M3 ;
        RECT 0.732 18.968 0.764 19 ;
  LAYER M1 ;
        RECT 0.796 16.512 0.828 19.02 ;
  LAYER M3 ;
        RECT 0.796 16.532 0.828 16.564 ;
  LAYER M1 ;
        RECT 0.86 16.512 0.892 19.02 ;
  LAYER M3 ;
        RECT 0.86 18.968 0.892 19 ;
  LAYER M1 ;
        RECT 0.924 16.512 0.956 19.02 ;
  LAYER M3 ;
        RECT 0.924 16.532 0.956 16.564 ;
  LAYER M1 ;
        RECT 0.988 16.512 1.02 19.02 ;
  LAYER M3 ;
        RECT 0.988 18.968 1.02 19 ;
  LAYER M1 ;
        RECT 1.052 16.512 1.084 19.02 ;
  LAYER M3 ;
        RECT 1.052 16.532 1.084 16.564 ;
  LAYER M1 ;
        RECT 1.116 16.512 1.148 19.02 ;
  LAYER M3 ;
        RECT 1.116 18.968 1.148 19 ;
  LAYER M1 ;
        RECT 1.18 16.512 1.212 19.02 ;
  LAYER M3 ;
        RECT 1.18 16.532 1.212 16.564 ;
  LAYER M1 ;
        RECT 1.244 16.512 1.276 19.02 ;
  LAYER M3 ;
        RECT 1.244 18.968 1.276 19 ;
  LAYER M1 ;
        RECT 1.308 16.512 1.34 19.02 ;
  LAYER M3 ;
        RECT 1.308 16.532 1.34 16.564 ;
  LAYER M1 ;
        RECT 1.372 16.512 1.404 19.02 ;
  LAYER M3 ;
        RECT 1.372 18.968 1.404 19 ;
  LAYER M1 ;
        RECT 1.436 16.512 1.468 19.02 ;
  LAYER M3 ;
        RECT 1.436 16.532 1.468 16.564 ;
  LAYER M1 ;
        RECT 1.5 16.512 1.532 19.02 ;
  LAYER M3 ;
        RECT 1.5 18.968 1.532 19 ;
  LAYER M1 ;
        RECT 1.564 16.512 1.596 19.02 ;
  LAYER M3 ;
        RECT 1.564 16.532 1.596 16.564 ;
  LAYER M1 ;
        RECT 1.628 16.512 1.66 19.02 ;
  LAYER M3 ;
        RECT 1.628 18.968 1.66 19 ;
  LAYER M1 ;
        RECT 1.692 16.512 1.724 19.02 ;
  LAYER M3 ;
        RECT 1.692 16.532 1.724 16.564 ;
  LAYER M1 ;
        RECT 1.756 16.512 1.788 19.02 ;
  LAYER M3 ;
        RECT 1.756 18.968 1.788 19 ;
  LAYER M1 ;
        RECT 1.82 16.512 1.852 19.02 ;
  LAYER M3 ;
        RECT 1.82 16.532 1.852 16.564 ;
  LAYER M1 ;
        RECT 1.884 16.512 1.916 19.02 ;
  LAYER M3 ;
        RECT 1.884 18.968 1.916 19 ;
  LAYER M1 ;
        RECT 1.948 16.512 1.98 19.02 ;
  LAYER M3 ;
        RECT 1.948 16.532 1.98 16.564 ;
  LAYER M1 ;
        RECT 2.012 16.512 2.044 19.02 ;
  LAYER M3 ;
        RECT 2.012 18.968 2.044 19 ;
  LAYER M1 ;
        RECT 2.076 16.512 2.108 19.02 ;
  LAYER M3 ;
        RECT 2.076 16.532 2.108 16.564 ;
  LAYER M1 ;
        RECT 2.14 16.512 2.172 19.02 ;
  LAYER M3 ;
        RECT 2.14 18.968 2.172 19 ;
  LAYER M1 ;
        RECT 2.204 16.512 2.236 19.02 ;
  LAYER M3 ;
        RECT 2.204 16.532 2.236 16.564 ;
  LAYER M1 ;
        RECT 2.268 16.512 2.3 19.02 ;
  LAYER M3 ;
        RECT 2.268 18.968 2.3 19 ;
  LAYER M1 ;
        RECT 2.332 16.512 2.364 19.02 ;
  LAYER M3 ;
        RECT 2.332 16.532 2.364 16.564 ;
  LAYER M1 ;
        RECT 2.396 16.512 2.428 19.02 ;
  LAYER M3 ;
        RECT 2.396 18.968 2.428 19 ;
  LAYER M1 ;
        RECT 2.46 16.512 2.492 19.02 ;
  LAYER M3 ;
        RECT 0.092 16.596 0.124 16.628 ;
  LAYER M2 ;
        RECT 2.46 16.66 2.492 16.692 ;
  LAYER M2 ;
        RECT 0.092 16.724 0.124 16.756 ;
  LAYER M2 ;
        RECT 2.46 16.788 2.492 16.82 ;
  LAYER M2 ;
        RECT 0.092 16.852 0.124 16.884 ;
  LAYER M2 ;
        RECT 2.46 16.916 2.492 16.948 ;
  LAYER M2 ;
        RECT 0.092 16.98 0.124 17.012 ;
  LAYER M2 ;
        RECT 2.46 17.044 2.492 17.076 ;
  LAYER M2 ;
        RECT 0.092 17.108 0.124 17.14 ;
  LAYER M2 ;
        RECT 2.46 17.172 2.492 17.204 ;
  LAYER M2 ;
        RECT 0.092 17.236 0.124 17.268 ;
  LAYER M2 ;
        RECT 2.46 17.3 2.492 17.332 ;
  LAYER M2 ;
        RECT 0.092 17.364 0.124 17.396 ;
  LAYER M2 ;
        RECT 2.46 17.428 2.492 17.46 ;
  LAYER M2 ;
        RECT 0.092 17.492 0.124 17.524 ;
  LAYER M2 ;
        RECT 2.46 17.556 2.492 17.588 ;
  LAYER M2 ;
        RECT 0.092 17.62 0.124 17.652 ;
  LAYER M2 ;
        RECT 2.46 17.684 2.492 17.716 ;
  LAYER M2 ;
        RECT 0.092 17.748 0.124 17.78 ;
  LAYER M2 ;
        RECT 2.46 17.812 2.492 17.844 ;
  LAYER M2 ;
        RECT 0.092 17.876 0.124 17.908 ;
  LAYER M2 ;
        RECT 2.46 17.94 2.492 17.972 ;
  LAYER M2 ;
        RECT 0.092 18.004 0.124 18.036 ;
  LAYER M2 ;
        RECT 2.46 18.068 2.492 18.1 ;
  LAYER M2 ;
        RECT 0.092 18.132 0.124 18.164 ;
  LAYER M2 ;
        RECT 2.46 18.196 2.492 18.228 ;
  LAYER M2 ;
        RECT 0.092 18.26 0.124 18.292 ;
  LAYER M2 ;
        RECT 2.46 18.324 2.492 18.356 ;
  LAYER M2 ;
        RECT 0.092 18.388 0.124 18.42 ;
  LAYER M2 ;
        RECT 2.46 18.452 2.492 18.484 ;
  LAYER M2 ;
        RECT 0.092 18.516 0.124 18.548 ;
  LAYER M2 ;
        RECT 2.46 18.58 2.492 18.612 ;
  LAYER M2 ;
        RECT 0.092 18.644 0.124 18.676 ;
  LAYER M2 ;
        RECT 2.46 18.708 2.492 18.74 ;
  LAYER M2 ;
        RECT 0.092 18.772 0.124 18.804 ;
  LAYER M2 ;
        RECT 2.46 18.836 2.492 18.868 ;
  LAYER M2 ;
        RECT 0.044 16.464 2.54 19.068 ;
  LAYER M1 ;
        RECT 3.708 0.972 3.74 3.48 ;
  LAYER M3 ;
        RECT 3.708 3.428 3.74 3.46 ;
  LAYER M1 ;
        RECT 3.772 0.972 3.804 3.48 ;
  LAYER M3 ;
        RECT 3.772 0.992 3.804 1.024 ;
  LAYER M1 ;
        RECT 3.836 0.972 3.868 3.48 ;
  LAYER M3 ;
        RECT 3.836 3.428 3.868 3.46 ;
  LAYER M1 ;
        RECT 3.9 0.972 3.932 3.48 ;
  LAYER M3 ;
        RECT 3.9 0.992 3.932 1.024 ;
  LAYER M1 ;
        RECT 3.964 0.972 3.996 3.48 ;
  LAYER M3 ;
        RECT 3.964 3.428 3.996 3.46 ;
  LAYER M1 ;
        RECT 4.028 0.972 4.06 3.48 ;
  LAYER M3 ;
        RECT 4.028 0.992 4.06 1.024 ;
  LAYER M1 ;
        RECT 4.092 0.972 4.124 3.48 ;
  LAYER M3 ;
        RECT 4.092 3.428 4.124 3.46 ;
  LAYER M1 ;
        RECT 4.156 0.972 4.188 3.48 ;
  LAYER M3 ;
        RECT 4.156 0.992 4.188 1.024 ;
  LAYER M1 ;
        RECT 4.22 0.972 4.252 3.48 ;
  LAYER M3 ;
        RECT 4.22 3.428 4.252 3.46 ;
  LAYER M1 ;
        RECT 4.284 0.972 4.316 3.48 ;
  LAYER M3 ;
        RECT 4.284 0.992 4.316 1.024 ;
  LAYER M1 ;
        RECT 4.348 0.972 4.38 3.48 ;
  LAYER M3 ;
        RECT 4.348 3.428 4.38 3.46 ;
  LAYER M1 ;
        RECT 4.412 0.972 4.444 3.48 ;
  LAYER M3 ;
        RECT 4.412 0.992 4.444 1.024 ;
  LAYER M1 ;
        RECT 4.476 0.972 4.508 3.48 ;
  LAYER M3 ;
        RECT 4.476 3.428 4.508 3.46 ;
  LAYER M1 ;
        RECT 4.54 0.972 4.572 3.48 ;
  LAYER M3 ;
        RECT 4.54 0.992 4.572 1.024 ;
  LAYER M1 ;
        RECT 4.604 0.972 4.636 3.48 ;
  LAYER M3 ;
        RECT 4.604 3.428 4.636 3.46 ;
  LAYER M1 ;
        RECT 4.668 0.972 4.7 3.48 ;
  LAYER M3 ;
        RECT 4.668 0.992 4.7 1.024 ;
  LAYER M1 ;
        RECT 4.732 0.972 4.764 3.48 ;
  LAYER M3 ;
        RECT 4.732 3.428 4.764 3.46 ;
  LAYER M1 ;
        RECT 4.796 0.972 4.828 3.48 ;
  LAYER M3 ;
        RECT 4.796 0.992 4.828 1.024 ;
  LAYER M1 ;
        RECT 4.86 0.972 4.892 3.48 ;
  LAYER M3 ;
        RECT 4.86 3.428 4.892 3.46 ;
  LAYER M1 ;
        RECT 4.924 0.972 4.956 3.48 ;
  LAYER M3 ;
        RECT 4.924 0.992 4.956 1.024 ;
  LAYER M1 ;
        RECT 4.988 0.972 5.02 3.48 ;
  LAYER M3 ;
        RECT 4.988 3.428 5.02 3.46 ;
  LAYER M1 ;
        RECT 5.052 0.972 5.084 3.48 ;
  LAYER M3 ;
        RECT 5.052 0.992 5.084 1.024 ;
  LAYER M1 ;
        RECT 5.116 0.972 5.148 3.48 ;
  LAYER M3 ;
        RECT 5.116 3.428 5.148 3.46 ;
  LAYER M1 ;
        RECT 5.18 0.972 5.212 3.48 ;
  LAYER M3 ;
        RECT 5.18 0.992 5.212 1.024 ;
  LAYER M1 ;
        RECT 5.244 0.972 5.276 3.48 ;
  LAYER M3 ;
        RECT 5.244 3.428 5.276 3.46 ;
  LAYER M1 ;
        RECT 5.308 0.972 5.34 3.48 ;
  LAYER M3 ;
        RECT 5.308 0.992 5.34 1.024 ;
  LAYER M1 ;
        RECT 5.372 0.972 5.404 3.48 ;
  LAYER M3 ;
        RECT 5.372 3.428 5.404 3.46 ;
  LAYER M1 ;
        RECT 5.436 0.972 5.468 3.48 ;
  LAYER M3 ;
        RECT 5.436 0.992 5.468 1.024 ;
  LAYER M1 ;
        RECT 5.5 0.972 5.532 3.48 ;
  LAYER M3 ;
        RECT 5.5 3.428 5.532 3.46 ;
  LAYER M1 ;
        RECT 5.564 0.972 5.596 3.48 ;
  LAYER M3 ;
        RECT 5.564 0.992 5.596 1.024 ;
  LAYER M1 ;
        RECT 5.628 0.972 5.66 3.48 ;
  LAYER M3 ;
        RECT 5.628 3.428 5.66 3.46 ;
  LAYER M1 ;
        RECT 5.692 0.972 5.724 3.48 ;
  LAYER M3 ;
        RECT 5.692 0.992 5.724 1.024 ;
  LAYER M1 ;
        RECT 5.756 0.972 5.788 3.48 ;
  LAYER M3 ;
        RECT 5.756 3.428 5.788 3.46 ;
  LAYER M1 ;
        RECT 5.82 0.972 5.852 3.48 ;
  LAYER M3 ;
        RECT 5.82 0.992 5.852 1.024 ;
  LAYER M1 ;
        RECT 5.884 0.972 5.916 3.48 ;
  LAYER M3 ;
        RECT 5.884 3.428 5.916 3.46 ;
  LAYER M1 ;
        RECT 5.948 0.972 5.98 3.48 ;
  LAYER M3 ;
        RECT 5.948 0.992 5.98 1.024 ;
  LAYER M1 ;
        RECT 6.012 0.972 6.044 3.48 ;
  LAYER M3 ;
        RECT 6.012 3.428 6.044 3.46 ;
  LAYER M1 ;
        RECT 6.076 0.972 6.108 3.48 ;
  LAYER M3 ;
        RECT 3.708 1.056 3.74 1.088 ;
  LAYER M2 ;
        RECT 6.076 1.12 6.108 1.152 ;
  LAYER M2 ;
        RECT 3.708 1.184 3.74 1.216 ;
  LAYER M2 ;
        RECT 6.076 1.248 6.108 1.28 ;
  LAYER M2 ;
        RECT 3.708 1.312 3.74 1.344 ;
  LAYER M2 ;
        RECT 6.076 1.376 6.108 1.408 ;
  LAYER M2 ;
        RECT 3.708 1.44 3.74 1.472 ;
  LAYER M2 ;
        RECT 6.076 1.504 6.108 1.536 ;
  LAYER M2 ;
        RECT 3.708 1.568 3.74 1.6 ;
  LAYER M2 ;
        RECT 6.076 1.632 6.108 1.664 ;
  LAYER M2 ;
        RECT 3.708 1.696 3.74 1.728 ;
  LAYER M2 ;
        RECT 6.076 1.76 6.108 1.792 ;
  LAYER M2 ;
        RECT 3.708 1.824 3.74 1.856 ;
  LAYER M2 ;
        RECT 6.076 1.888 6.108 1.92 ;
  LAYER M2 ;
        RECT 3.708 1.952 3.74 1.984 ;
  LAYER M2 ;
        RECT 6.076 2.016 6.108 2.048 ;
  LAYER M2 ;
        RECT 3.708 2.08 3.74 2.112 ;
  LAYER M2 ;
        RECT 6.076 2.144 6.108 2.176 ;
  LAYER M2 ;
        RECT 3.708 2.208 3.74 2.24 ;
  LAYER M2 ;
        RECT 6.076 2.272 6.108 2.304 ;
  LAYER M2 ;
        RECT 3.708 2.336 3.74 2.368 ;
  LAYER M2 ;
        RECT 6.076 2.4 6.108 2.432 ;
  LAYER M2 ;
        RECT 3.708 2.464 3.74 2.496 ;
  LAYER M2 ;
        RECT 6.076 2.528 6.108 2.56 ;
  LAYER M2 ;
        RECT 3.708 2.592 3.74 2.624 ;
  LAYER M2 ;
        RECT 6.076 2.656 6.108 2.688 ;
  LAYER M2 ;
        RECT 3.708 2.72 3.74 2.752 ;
  LAYER M2 ;
        RECT 6.076 2.784 6.108 2.816 ;
  LAYER M2 ;
        RECT 3.708 2.848 3.74 2.88 ;
  LAYER M2 ;
        RECT 6.076 2.912 6.108 2.944 ;
  LAYER M2 ;
        RECT 3.708 2.976 3.74 3.008 ;
  LAYER M2 ;
        RECT 6.076 3.04 6.108 3.072 ;
  LAYER M2 ;
        RECT 3.708 3.104 3.74 3.136 ;
  LAYER M2 ;
        RECT 6.076 3.168 6.108 3.2 ;
  LAYER M2 ;
        RECT 3.708 3.232 3.74 3.264 ;
  LAYER M2 ;
        RECT 6.076 3.296 6.108 3.328 ;
  LAYER M2 ;
        RECT 3.66 0.924 6.156 3.528 ;
  LAYER M1 ;
        RECT 3.708 4.08 3.74 6.588 ;
  LAYER M3 ;
        RECT 3.708 6.536 3.74 6.568 ;
  LAYER M1 ;
        RECT 3.772 4.08 3.804 6.588 ;
  LAYER M3 ;
        RECT 3.772 4.1 3.804 4.132 ;
  LAYER M1 ;
        RECT 3.836 4.08 3.868 6.588 ;
  LAYER M3 ;
        RECT 3.836 6.536 3.868 6.568 ;
  LAYER M1 ;
        RECT 3.9 4.08 3.932 6.588 ;
  LAYER M3 ;
        RECT 3.9 4.1 3.932 4.132 ;
  LAYER M1 ;
        RECT 3.964 4.08 3.996 6.588 ;
  LAYER M3 ;
        RECT 3.964 6.536 3.996 6.568 ;
  LAYER M1 ;
        RECT 4.028 4.08 4.06 6.588 ;
  LAYER M3 ;
        RECT 4.028 4.1 4.06 4.132 ;
  LAYER M1 ;
        RECT 4.092 4.08 4.124 6.588 ;
  LAYER M3 ;
        RECT 4.092 6.536 4.124 6.568 ;
  LAYER M1 ;
        RECT 4.156 4.08 4.188 6.588 ;
  LAYER M3 ;
        RECT 4.156 4.1 4.188 4.132 ;
  LAYER M1 ;
        RECT 4.22 4.08 4.252 6.588 ;
  LAYER M3 ;
        RECT 4.22 6.536 4.252 6.568 ;
  LAYER M1 ;
        RECT 4.284 4.08 4.316 6.588 ;
  LAYER M3 ;
        RECT 4.284 4.1 4.316 4.132 ;
  LAYER M1 ;
        RECT 4.348 4.08 4.38 6.588 ;
  LAYER M3 ;
        RECT 4.348 6.536 4.38 6.568 ;
  LAYER M1 ;
        RECT 4.412 4.08 4.444 6.588 ;
  LAYER M3 ;
        RECT 4.412 4.1 4.444 4.132 ;
  LAYER M1 ;
        RECT 4.476 4.08 4.508 6.588 ;
  LAYER M3 ;
        RECT 4.476 6.536 4.508 6.568 ;
  LAYER M1 ;
        RECT 4.54 4.08 4.572 6.588 ;
  LAYER M3 ;
        RECT 4.54 4.1 4.572 4.132 ;
  LAYER M1 ;
        RECT 4.604 4.08 4.636 6.588 ;
  LAYER M3 ;
        RECT 4.604 6.536 4.636 6.568 ;
  LAYER M1 ;
        RECT 4.668 4.08 4.7 6.588 ;
  LAYER M3 ;
        RECT 4.668 4.1 4.7 4.132 ;
  LAYER M1 ;
        RECT 4.732 4.08 4.764 6.588 ;
  LAYER M3 ;
        RECT 4.732 6.536 4.764 6.568 ;
  LAYER M1 ;
        RECT 4.796 4.08 4.828 6.588 ;
  LAYER M3 ;
        RECT 4.796 4.1 4.828 4.132 ;
  LAYER M1 ;
        RECT 4.86 4.08 4.892 6.588 ;
  LAYER M3 ;
        RECT 4.86 6.536 4.892 6.568 ;
  LAYER M1 ;
        RECT 4.924 4.08 4.956 6.588 ;
  LAYER M3 ;
        RECT 4.924 4.1 4.956 4.132 ;
  LAYER M1 ;
        RECT 4.988 4.08 5.02 6.588 ;
  LAYER M3 ;
        RECT 4.988 6.536 5.02 6.568 ;
  LAYER M1 ;
        RECT 5.052 4.08 5.084 6.588 ;
  LAYER M3 ;
        RECT 5.052 4.1 5.084 4.132 ;
  LAYER M1 ;
        RECT 5.116 4.08 5.148 6.588 ;
  LAYER M3 ;
        RECT 5.116 6.536 5.148 6.568 ;
  LAYER M1 ;
        RECT 5.18 4.08 5.212 6.588 ;
  LAYER M3 ;
        RECT 5.18 4.1 5.212 4.132 ;
  LAYER M1 ;
        RECT 5.244 4.08 5.276 6.588 ;
  LAYER M3 ;
        RECT 5.244 6.536 5.276 6.568 ;
  LAYER M1 ;
        RECT 5.308 4.08 5.34 6.588 ;
  LAYER M3 ;
        RECT 5.308 4.1 5.34 4.132 ;
  LAYER M1 ;
        RECT 5.372 4.08 5.404 6.588 ;
  LAYER M3 ;
        RECT 5.372 6.536 5.404 6.568 ;
  LAYER M1 ;
        RECT 5.436 4.08 5.468 6.588 ;
  LAYER M3 ;
        RECT 5.436 4.1 5.468 4.132 ;
  LAYER M1 ;
        RECT 5.5 4.08 5.532 6.588 ;
  LAYER M3 ;
        RECT 5.5 6.536 5.532 6.568 ;
  LAYER M1 ;
        RECT 5.564 4.08 5.596 6.588 ;
  LAYER M3 ;
        RECT 5.564 4.1 5.596 4.132 ;
  LAYER M1 ;
        RECT 5.628 4.08 5.66 6.588 ;
  LAYER M3 ;
        RECT 5.628 6.536 5.66 6.568 ;
  LAYER M1 ;
        RECT 5.692 4.08 5.724 6.588 ;
  LAYER M3 ;
        RECT 5.692 4.1 5.724 4.132 ;
  LAYER M1 ;
        RECT 5.756 4.08 5.788 6.588 ;
  LAYER M3 ;
        RECT 5.756 6.536 5.788 6.568 ;
  LAYER M1 ;
        RECT 5.82 4.08 5.852 6.588 ;
  LAYER M3 ;
        RECT 5.82 4.1 5.852 4.132 ;
  LAYER M1 ;
        RECT 5.884 4.08 5.916 6.588 ;
  LAYER M3 ;
        RECT 5.884 6.536 5.916 6.568 ;
  LAYER M1 ;
        RECT 5.948 4.08 5.98 6.588 ;
  LAYER M3 ;
        RECT 5.948 4.1 5.98 4.132 ;
  LAYER M1 ;
        RECT 6.012 4.08 6.044 6.588 ;
  LAYER M3 ;
        RECT 6.012 6.536 6.044 6.568 ;
  LAYER M1 ;
        RECT 6.076 4.08 6.108 6.588 ;
  LAYER M3 ;
        RECT 3.708 4.164 3.74 4.196 ;
  LAYER M2 ;
        RECT 6.076 4.228 6.108 4.26 ;
  LAYER M2 ;
        RECT 3.708 4.292 3.74 4.324 ;
  LAYER M2 ;
        RECT 6.076 4.356 6.108 4.388 ;
  LAYER M2 ;
        RECT 3.708 4.42 3.74 4.452 ;
  LAYER M2 ;
        RECT 6.076 4.484 6.108 4.516 ;
  LAYER M2 ;
        RECT 3.708 4.548 3.74 4.58 ;
  LAYER M2 ;
        RECT 6.076 4.612 6.108 4.644 ;
  LAYER M2 ;
        RECT 3.708 4.676 3.74 4.708 ;
  LAYER M2 ;
        RECT 6.076 4.74 6.108 4.772 ;
  LAYER M2 ;
        RECT 3.708 4.804 3.74 4.836 ;
  LAYER M2 ;
        RECT 6.076 4.868 6.108 4.9 ;
  LAYER M2 ;
        RECT 3.708 4.932 3.74 4.964 ;
  LAYER M2 ;
        RECT 6.076 4.996 6.108 5.028 ;
  LAYER M2 ;
        RECT 3.708 5.06 3.74 5.092 ;
  LAYER M2 ;
        RECT 6.076 5.124 6.108 5.156 ;
  LAYER M2 ;
        RECT 3.708 5.188 3.74 5.22 ;
  LAYER M2 ;
        RECT 6.076 5.252 6.108 5.284 ;
  LAYER M2 ;
        RECT 3.708 5.316 3.74 5.348 ;
  LAYER M2 ;
        RECT 6.076 5.38 6.108 5.412 ;
  LAYER M2 ;
        RECT 3.708 5.444 3.74 5.476 ;
  LAYER M2 ;
        RECT 6.076 5.508 6.108 5.54 ;
  LAYER M2 ;
        RECT 3.708 5.572 3.74 5.604 ;
  LAYER M2 ;
        RECT 6.076 5.636 6.108 5.668 ;
  LAYER M2 ;
        RECT 3.708 5.7 3.74 5.732 ;
  LAYER M2 ;
        RECT 6.076 5.764 6.108 5.796 ;
  LAYER M2 ;
        RECT 3.708 5.828 3.74 5.86 ;
  LAYER M2 ;
        RECT 6.076 5.892 6.108 5.924 ;
  LAYER M2 ;
        RECT 3.708 5.956 3.74 5.988 ;
  LAYER M2 ;
        RECT 6.076 6.02 6.108 6.052 ;
  LAYER M2 ;
        RECT 3.708 6.084 3.74 6.116 ;
  LAYER M2 ;
        RECT 6.076 6.148 6.108 6.18 ;
  LAYER M2 ;
        RECT 3.708 6.212 3.74 6.244 ;
  LAYER M2 ;
        RECT 6.076 6.276 6.108 6.308 ;
  LAYER M2 ;
        RECT 3.708 6.34 3.74 6.372 ;
  LAYER M2 ;
        RECT 6.076 6.404 6.108 6.436 ;
  LAYER M2 ;
        RECT 3.66 4.032 6.156 6.636 ;
  LAYER M1 ;
        RECT 3.708 7.188 3.74 9.696 ;
  LAYER M3 ;
        RECT 3.708 9.644 3.74 9.676 ;
  LAYER M1 ;
        RECT 3.772 7.188 3.804 9.696 ;
  LAYER M3 ;
        RECT 3.772 7.208 3.804 7.24 ;
  LAYER M1 ;
        RECT 3.836 7.188 3.868 9.696 ;
  LAYER M3 ;
        RECT 3.836 9.644 3.868 9.676 ;
  LAYER M1 ;
        RECT 3.9 7.188 3.932 9.696 ;
  LAYER M3 ;
        RECT 3.9 7.208 3.932 7.24 ;
  LAYER M1 ;
        RECT 3.964 7.188 3.996 9.696 ;
  LAYER M3 ;
        RECT 3.964 9.644 3.996 9.676 ;
  LAYER M1 ;
        RECT 4.028 7.188 4.06 9.696 ;
  LAYER M3 ;
        RECT 4.028 7.208 4.06 7.24 ;
  LAYER M1 ;
        RECT 4.092 7.188 4.124 9.696 ;
  LAYER M3 ;
        RECT 4.092 9.644 4.124 9.676 ;
  LAYER M1 ;
        RECT 4.156 7.188 4.188 9.696 ;
  LAYER M3 ;
        RECT 4.156 7.208 4.188 7.24 ;
  LAYER M1 ;
        RECT 4.22 7.188 4.252 9.696 ;
  LAYER M3 ;
        RECT 4.22 9.644 4.252 9.676 ;
  LAYER M1 ;
        RECT 4.284 7.188 4.316 9.696 ;
  LAYER M3 ;
        RECT 4.284 7.208 4.316 7.24 ;
  LAYER M1 ;
        RECT 4.348 7.188 4.38 9.696 ;
  LAYER M3 ;
        RECT 4.348 9.644 4.38 9.676 ;
  LAYER M1 ;
        RECT 4.412 7.188 4.444 9.696 ;
  LAYER M3 ;
        RECT 4.412 7.208 4.444 7.24 ;
  LAYER M1 ;
        RECT 4.476 7.188 4.508 9.696 ;
  LAYER M3 ;
        RECT 4.476 9.644 4.508 9.676 ;
  LAYER M1 ;
        RECT 4.54 7.188 4.572 9.696 ;
  LAYER M3 ;
        RECT 4.54 7.208 4.572 7.24 ;
  LAYER M1 ;
        RECT 4.604 7.188 4.636 9.696 ;
  LAYER M3 ;
        RECT 4.604 9.644 4.636 9.676 ;
  LAYER M1 ;
        RECT 4.668 7.188 4.7 9.696 ;
  LAYER M3 ;
        RECT 4.668 7.208 4.7 7.24 ;
  LAYER M1 ;
        RECT 4.732 7.188 4.764 9.696 ;
  LAYER M3 ;
        RECT 4.732 9.644 4.764 9.676 ;
  LAYER M1 ;
        RECT 4.796 7.188 4.828 9.696 ;
  LAYER M3 ;
        RECT 4.796 7.208 4.828 7.24 ;
  LAYER M1 ;
        RECT 4.86 7.188 4.892 9.696 ;
  LAYER M3 ;
        RECT 4.86 9.644 4.892 9.676 ;
  LAYER M1 ;
        RECT 4.924 7.188 4.956 9.696 ;
  LAYER M3 ;
        RECT 4.924 7.208 4.956 7.24 ;
  LAYER M1 ;
        RECT 4.988 7.188 5.02 9.696 ;
  LAYER M3 ;
        RECT 4.988 9.644 5.02 9.676 ;
  LAYER M1 ;
        RECT 5.052 7.188 5.084 9.696 ;
  LAYER M3 ;
        RECT 5.052 7.208 5.084 7.24 ;
  LAYER M1 ;
        RECT 5.116 7.188 5.148 9.696 ;
  LAYER M3 ;
        RECT 5.116 9.644 5.148 9.676 ;
  LAYER M1 ;
        RECT 5.18 7.188 5.212 9.696 ;
  LAYER M3 ;
        RECT 5.18 7.208 5.212 7.24 ;
  LAYER M1 ;
        RECT 5.244 7.188 5.276 9.696 ;
  LAYER M3 ;
        RECT 5.244 9.644 5.276 9.676 ;
  LAYER M1 ;
        RECT 5.308 7.188 5.34 9.696 ;
  LAYER M3 ;
        RECT 5.308 7.208 5.34 7.24 ;
  LAYER M1 ;
        RECT 5.372 7.188 5.404 9.696 ;
  LAYER M3 ;
        RECT 5.372 9.644 5.404 9.676 ;
  LAYER M1 ;
        RECT 5.436 7.188 5.468 9.696 ;
  LAYER M3 ;
        RECT 5.436 7.208 5.468 7.24 ;
  LAYER M1 ;
        RECT 5.5 7.188 5.532 9.696 ;
  LAYER M3 ;
        RECT 5.5 9.644 5.532 9.676 ;
  LAYER M1 ;
        RECT 5.564 7.188 5.596 9.696 ;
  LAYER M3 ;
        RECT 5.564 7.208 5.596 7.24 ;
  LAYER M1 ;
        RECT 5.628 7.188 5.66 9.696 ;
  LAYER M3 ;
        RECT 5.628 9.644 5.66 9.676 ;
  LAYER M1 ;
        RECT 5.692 7.188 5.724 9.696 ;
  LAYER M3 ;
        RECT 5.692 7.208 5.724 7.24 ;
  LAYER M1 ;
        RECT 5.756 7.188 5.788 9.696 ;
  LAYER M3 ;
        RECT 5.756 9.644 5.788 9.676 ;
  LAYER M1 ;
        RECT 5.82 7.188 5.852 9.696 ;
  LAYER M3 ;
        RECT 5.82 7.208 5.852 7.24 ;
  LAYER M1 ;
        RECT 5.884 7.188 5.916 9.696 ;
  LAYER M3 ;
        RECT 5.884 9.644 5.916 9.676 ;
  LAYER M1 ;
        RECT 5.948 7.188 5.98 9.696 ;
  LAYER M3 ;
        RECT 5.948 7.208 5.98 7.24 ;
  LAYER M1 ;
        RECT 6.012 7.188 6.044 9.696 ;
  LAYER M3 ;
        RECT 6.012 9.644 6.044 9.676 ;
  LAYER M1 ;
        RECT 6.076 7.188 6.108 9.696 ;
  LAYER M3 ;
        RECT 3.708 7.272 3.74 7.304 ;
  LAYER M2 ;
        RECT 6.076 7.336 6.108 7.368 ;
  LAYER M2 ;
        RECT 3.708 7.4 3.74 7.432 ;
  LAYER M2 ;
        RECT 6.076 7.464 6.108 7.496 ;
  LAYER M2 ;
        RECT 3.708 7.528 3.74 7.56 ;
  LAYER M2 ;
        RECT 6.076 7.592 6.108 7.624 ;
  LAYER M2 ;
        RECT 3.708 7.656 3.74 7.688 ;
  LAYER M2 ;
        RECT 6.076 7.72 6.108 7.752 ;
  LAYER M2 ;
        RECT 3.708 7.784 3.74 7.816 ;
  LAYER M2 ;
        RECT 6.076 7.848 6.108 7.88 ;
  LAYER M2 ;
        RECT 3.708 7.912 3.74 7.944 ;
  LAYER M2 ;
        RECT 6.076 7.976 6.108 8.008 ;
  LAYER M2 ;
        RECT 3.708 8.04 3.74 8.072 ;
  LAYER M2 ;
        RECT 6.076 8.104 6.108 8.136 ;
  LAYER M2 ;
        RECT 3.708 8.168 3.74 8.2 ;
  LAYER M2 ;
        RECT 6.076 8.232 6.108 8.264 ;
  LAYER M2 ;
        RECT 3.708 8.296 3.74 8.328 ;
  LAYER M2 ;
        RECT 6.076 8.36 6.108 8.392 ;
  LAYER M2 ;
        RECT 3.708 8.424 3.74 8.456 ;
  LAYER M2 ;
        RECT 6.076 8.488 6.108 8.52 ;
  LAYER M2 ;
        RECT 3.708 8.552 3.74 8.584 ;
  LAYER M2 ;
        RECT 6.076 8.616 6.108 8.648 ;
  LAYER M2 ;
        RECT 3.708 8.68 3.74 8.712 ;
  LAYER M2 ;
        RECT 6.076 8.744 6.108 8.776 ;
  LAYER M2 ;
        RECT 3.708 8.808 3.74 8.84 ;
  LAYER M2 ;
        RECT 6.076 8.872 6.108 8.904 ;
  LAYER M2 ;
        RECT 3.708 8.936 3.74 8.968 ;
  LAYER M2 ;
        RECT 6.076 9 6.108 9.032 ;
  LAYER M2 ;
        RECT 3.708 9.064 3.74 9.096 ;
  LAYER M2 ;
        RECT 6.076 9.128 6.108 9.16 ;
  LAYER M2 ;
        RECT 3.708 9.192 3.74 9.224 ;
  LAYER M2 ;
        RECT 6.076 9.256 6.108 9.288 ;
  LAYER M2 ;
        RECT 3.708 9.32 3.74 9.352 ;
  LAYER M2 ;
        RECT 6.076 9.384 6.108 9.416 ;
  LAYER M2 ;
        RECT 3.708 9.448 3.74 9.48 ;
  LAYER M2 ;
        RECT 6.076 9.512 6.108 9.544 ;
  LAYER M2 ;
        RECT 3.66 7.14 6.156 9.744 ;
  LAYER M1 ;
        RECT 3.708 10.296 3.74 12.804 ;
  LAYER M3 ;
        RECT 3.708 12.752 3.74 12.784 ;
  LAYER M1 ;
        RECT 3.772 10.296 3.804 12.804 ;
  LAYER M3 ;
        RECT 3.772 10.316 3.804 10.348 ;
  LAYER M1 ;
        RECT 3.836 10.296 3.868 12.804 ;
  LAYER M3 ;
        RECT 3.836 12.752 3.868 12.784 ;
  LAYER M1 ;
        RECT 3.9 10.296 3.932 12.804 ;
  LAYER M3 ;
        RECT 3.9 10.316 3.932 10.348 ;
  LAYER M1 ;
        RECT 3.964 10.296 3.996 12.804 ;
  LAYER M3 ;
        RECT 3.964 12.752 3.996 12.784 ;
  LAYER M1 ;
        RECT 4.028 10.296 4.06 12.804 ;
  LAYER M3 ;
        RECT 4.028 10.316 4.06 10.348 ;
  LAYER M1 ;
        RECT 4.092 10.296 4.124 12.804 ;
  LAYER M3 ;
        RECT 4.092 12.752 4.124 12.784 ;
  LAYER M1 ;
        RECT 4.156 10.296 4.188 12.804 ;
  LAYER M3 ;
        RECT 4.156 10.316 4.188 10.348 ;
  LAYER M1 ;
        RECT 4.22 10.296 4.252 12.804 ;
  LAYER M3 ;
        RECT 4.22 12.752 4.252 12.784 ;
  LAYER M1 ;
        RECT 4.284 10.296 4.316 12.804 ;
  LAYER M3 ;
        RECT 4.284 10.316 4.316 10.348 ;
  LAYER M1 ;
        RECT 4.348 10.296 4.38 12.804 ;
  LAYER M3 ;
        RECT 4.348 12.752 4.38 12.784 ;
  LAYER M1 ;
        RECT 4.412 10.296 4.444 12.804 ;
  LAYER M3 ;
        RECT 4.412 10.316 4.444 10.348 ;
  LAYER M1 ;
        RECT 4.476 10.296 4.508 12.804 ;
  LAYER M3 ;
        RECT 4.476 12.752 4.508 12.784 ;
  LAYER M1 ;
        RECT 4.54 10.296 4.572 12.804 ;
  LAYER M3 ;
        RECT 4.54 10.316 4.572 10.348 ;
  LAYER M1 ;
        RECT 4.604 10.296 4.636 12.804 ;
  LAYER M3 ;
        RECT 4.604 12.752 4.636 12.784 ;
  LAYER M1 ;
        RECT 4.668 10.296 4.7 12.804 ;
  LAYER M3 ;
        RECT 4.668 10.316 4.7 10.348 ;
  LAYER M1 ;
        RECT 4.732 10.296 4.764 12.804 ;
  LAYER M3 ;
        RECT 4.732 12.752 4.764 12.784 ;
  LAYER M1 ;
        RECT 4.796 10.296 4.828 12.804 ;
  LAYER M3 ;
        RECT 4.796 10.316 4.828 10.348 ;
  LAYER M1 ;
        RECT 4.86 10.296 4.892 12.804 ;
  LAYER M3 ;
        RECT 4.86 12.752 4.892 12.784 ;
  LAYER M1 ;
        RECT 4.924 10.296 4.956 12.804 ;
  LAYER M3 ;
        RECT 4.924 10.316 4.956 10.348 ;
  LAYER M1 ;
        RECT 4.988 10.296 5.02 12.804 ;
  LAYER M3 ;
        RECT 4.988 12.752 5.02 12.784 ;
  LAYER M1 ;
        RECT 5.052 10.296 5.084 12.804 ;
  LAYER M3 ;
        RECT 5.052 10.316 5.084 10.348 ;
  LAYER M1 ;
        RECT 5.116 10.296 5.148 12.804 ;
  LAYER M3 ;
        RECT 5.116 12.752 5.148 12.784 ;
  LAYER M1 ;
        RECT 5.18 10.296 5.212 12.804 ;
  LAYER M3 ;
        RECT 5.18 10.316 5.212 10.348 ;
  LAYER M1 ;
        RECT 5.244 10.296 5.276 12.804 ;
  LAYER M3 ;
        RECT 5.244 12.752 5.276 12.784 ;
  LAYER M1 ;
        RECT 5.308 10.296 5.34 12.804 ;
  LAYER M3 ;
        RECT 5.308 10.316 5.34 10.348 ;
  LAYER M1 ;
        RECT 5.372 10.296 5.404 12.804 ;
  LAYER M3 ;
        RECT 5.372 12.752 5.404 12.784 ;
  LAYER M1 ;
        RECT 5.436 10.296 5.468 12.804 ;
  LAYER M3 ;
        RECT 5.436 10.316 5.468 10.348 ;
  LAYER M1 ;
        RECT 5.5 10.296 5.532 12.804 ;
  LAYER M3 ;
        RECT 5.5 12.752 5.532 12.784 ;
  LAYER M1 ;
        RECT 5.564 10.296 5.596 12.804 ;
  LAYER M3 ;
        RECT 5.564 10.316 5.596 10.348 ;
  LAYER M1 ;
        RECT 5.628 10.296 5.66 12.804 ;
  LAYER M3 ;
        RECT 5.628 12.752 5.66 12.784 ;
  LAYER M1 ;
        RECT 5.692 10.296 5.724 12.804 ;
  LAYER M3 ;
        RECT 5.692 10.316 5.724 10.348 ;
  LAYER M1 ;
        RECT 5.756 10.296 5.788 12.804 ;
  LAYER M3 ;
        RECT 5.756 12.752 5.788 12.784 ;
  LAYER M1 ;
        RECT 5.82 10.296 5.852 12.804 ;
  LAYER M3 ;
        RECT 5.82 10.316 5.852 10.348 ;
  LAYER M1 ;
        RECT 5.884 10.296 5.916 12.804 ;
  LAYER M3 ;
        RECT 5.884 12.752 5.916 12.784 ;
  LAYER M1 ;
        RECT 5.948 10.296 5.98 12.804 ;
  LAYER M3 ;
        RECT 5.948 10.316 5.98 10.348 ;
  LAYER M1 ;
        RECT 6.012 10.296 6.044 12.804 ;
  LAYER M3 ;
        RECT 6.012 12.752 6.044 12.784 ;
  LAYER M1 ;
        RECT 6.076 10.296 6.108 12.804 ;
  LAYER M3 ;
        RECT 3.708 10.38 3.74 10.412 ;
  LAYER M2 ;
        RECT 6.076 10.444 6.108 10.476 ;
  LAYER M2 ;
        RECT 3.708 10.508 3.74 10.54 ;
  LAYER M2 ;
        RECT 6.076 10.572 6.108 10.604 ;
  LAYER M2 ;
        RECT 3.708 10.636 3.74 10.668 ;
  LAYER M2 ;
        RECT 6.076 10.7 6.108 10.732 ;
  LAYER M2 ;
        RECT 3.708 10.764 3.74 10.796 ;
  LAYER M2 ;
        RECT 6.076 10.828 6.108 10.86 ;
  LAYER M2 ;
        RECT 3.708 10.892 3.74 10.924 ;
  LAYER M2 ;
        RECT 6.076 10.956 6.108 10.988 ;
  LAYER M2 ;
        RECT 3.708 11.02 3.74 11.052 ;
  LAYER M2 ;
        RECT 6.076 11.084 6.108 11.116 ;
  LAYER M2 ;
        RECT 3.708 11.148 3.74 11.18 ;
  LAYER M2 ;
        RECT 6.076 11.212 6.108 11.244 ;
  LAYER M2 ;
        RECT 3.708 11.276 3.74 11.308 ;
  LAYER M2 ;
        RECT 6.076 11.34 6.108 11.372 ;
  LAYER M2 ;
        RECT 3.708 11.404 3.74 11.436 ;
  LAYER M2 ;
        RECT 6.076 11.468 6.108 11.5 ;
  LAYER M2 ;
        RECT 3.708 11.532 3.74 11.564 ;
  LAYER M2 ;
        RECT 6.076 11.596 6.108 11.628 ;
  LAYER M2 ;
        RECT 3.708 11.66 3.74 11.692 ;
  LAYER M2 ;
        RECT 6.076 11.724 6.108 11.756 ;
  LAYER M2 ;
        RECT 3.708 11.788 3.74 11.82 ;
  LAYER M2 ;
        RECT 6.076 11.852 6.108 11.884 ;
  LAYER M2 ;
        RECT 3.708 11.916 3.74 11.948 ;
  LAYER M2 ;
        RECT 6.076 11.98 6.108 12.012 ;
  LAYER M2 ;
        RECT 3.708 12.044 3.74 12.076 ;
  LAYER M2 ;
        RECT 6.076 12.108 6.108 12.14 ;
  LAYER M2 ;
        RECT 3.708 12.172 3.74 12.204 ;
  LAYER M2 ;
        RECT 6.076 12.236 6.108 12.268 ;
  LAYER M2 ;
        RECT 3.708 12.3 3.74 12.332 ;
  LAYER M2 ;
        RECT 6.076 12.364 6.108 12.396 ;
  LAYER M2 ;
        RECT 3.708 12.428 3.74 12.46 ;
  LAYER M2 ;
        RECT 6.076 12.492 6.108 12.524 ;
  LAYER M2 ;
        RECT 3.708 12.556 3.74 12.588 ;
  LAYER M2 ;
        RECT 6.076 12.62 6.108 12.652 ;
  LAYER M2 ;
        RECT 3.66 10.248 6.156 12.852 ;
  LAYER M1 ;
        RECT 3.708 13.404 3.74 15.912 ;
  LAYER M3 ;
        RECT 3.708 15.86 3.74 15.892 ;
  LAYER M1 ;
        RECT 3.772 13.404 3.804 15.912 ;
  LAYER M3 ;
        RECT 3.772 13.424 3.804 13.456 ;
  LAYER M1 ;
        RECT 3.836 13.404 3.868 15.912 ;
  LAYER M3 ;
        RECT 3.836 15.86 3.868 15.892 ;
  LAYER M1 ;
        RECT 3.9 13.404 3.932 15.912 ;
  LAYER M3 ;
        RECT 3.9 13.424 3.932 13.456 ;
  LAYER M1 ;
        RECT 3.964 13.404 3.996 15.912 ;
  LAYER M3 ;
        RECT 3.964 15.86 3.996 15.892 ;
  LAYER M1 ;
        RECT 4.028 13.404 4.06 15.912 ;
  LAYER M3 ;
        RECT 4.028 13.424 4.06 13.456 ;
  LAYER M1 ;
        RECT 4.092 13.404 4.124 15.912 ;
  LAYER M3 ;
        RECT 4.092 15.86 4.124 15.892 ;
  LAYER M1 ;
        RECT 4.156 13.404 4.188 15.912 ;
  LAYER M3 ;
        RECT 4.156 13.424 4.188 13.456 ;
  LAYER M1 ;
        RECT 4.22 13.404 4.252 15.912 ;
  LAYER M3 ;
        RECT 4.22 15.86 4.252 15.892 ;
  LAYER M1 ;
        RECT 4.284 13.404 4.316 15.912 ;
  LAYER M3 ;
        RECT 4.284 13.424 4.316 13.456 ;
  LAYER M1 ;
        RECT 4.348 13.404 4.38 15.912 ;
  LAYER M3 ;
        RECT 4.348 15.86 4.38 15.892 ;
  LAYER M1 ;
        RECT 4.412 13.404 4.444 15.912 ;
  LAYER M3 ;
        RECT 4.412 13.424 4.444 13.456 ;
  LAYER M1 ;
        RECT 4.476 13.404 4.508 15.912 ;
  LAYER M3 ;
        RECT 4.476 15.86 4.508 15.892 ;
  LAYER M1 ;
        RECT 4.54 13.404 4.572 15.912 ;
  LAYER M3 ;
        RECT 4.54 13.424 4.572 13.456 ;
  LAYER M1 ;
        RECT 4.604 13.404 4.636 15.912 ;
  LAYER M3 ;
        RECT 4.604 15.86 4.636 15.892 ;
  LAYER M1 ;
        RECT 4.668 13.404 4.7 15.912 ;
  LAYER M3 ;
        RECT 4.668 13.424 4.7 13.456 ;
  LAYER M1 ;
        RECT 4.732 13.404 4.764 15.912 ;
  LAYER M3 ;
        RECT 4.732 15.86 4.764 15.892 ;
  LAYER M1 ;
        RECT 4.796 13.404 4.828 15.912 ;
  LAYER M3 ;
        RECT 4.796 13.424 4.828 13.456 ;
  LAYER M1 ;
        RECT 4.86 13.404 4.892 15.912 ;
  LAYER M3 ;
        RECT 4.86 15.86 4.892 15.892 ;
  LAYER M1 ;
        RECT 4.924 13.404 4.956 15.912 ;
  LAYER M3 ;
        RECT 4.924 13.424 4.956 13.456 ;
  LAYER M1 ;
        RECT 4.988 13.404 5.02 15.912 ;
  LAYER M3 ;
        RECT 4.988 15.86 5.02 15.892 ;
  LAYER M1 ;
        RECT 5.052 13.404 5.084 15.912 ;
  LAYER M3 ;
        RECT 5.052 13.424 5.084 13.456 ;
  LAYER M1 ;
        RECT 5.116 13.404 5.148 15.912 ;
  LAYER M3 ;
        RECT 5.116 15.86 5.148 15.892 ;
  LAYER M1 ;
        RECT 5.18 13.404 5.212 15.912 ;
  LAYER M3 ;
        RECT 5.18 13.424 5.212 13.456 ;
  LAYER M1 ;
        RECT 5.244 13.404 5.276 15.912 ;
  LAYER M3 ;
        RECT 5.244 15.86 5.276 15.892 ;
  LAYER M1 ;
        RECT 5.308 13.404 5.34 15.912 ;
  LAYER M3 ;
        RECT 5.308 13.424 5.34 13.456 ;
  LAYER M1 ;
        RECT 5.372 13.404 5.404 15.912 ;
  LAYER M3 ;
        RECT 5.372 15.86 5.404 15.892 ;
  LAYER M1 ;
        RECT 5.436 13.404 5.468 15.912 ;
  LAYER M3 ;
        RECT 5.436 13.424 5.468 13.456 ;
  LAYER M1 ;
        RECT 5.5 13.404 5.532 15.912 ;
  LAYER M3 ;
        RECT 5.5 15.86 5.532 15.892 ;
  LAYER M1 ;
        RECT 5.564 13.404 5.596 15.912 ;
  LAYER M3 ;
        RECT 5.564 13.424 5.596 13.456 ;
  LAYER M1 ;
        RECT 5.628 13.404 5.66 15.912 ;
  LAYER M3 ;
        RECT 5.628 15.86 5.66 15.892 ;
  LAYER M1 ;
        RECT 5.692 13.404 5.724 15.912 ;
  LAYER M3 ;
        RECT 5.692 13.424 5.724 13.456 ;
  LAYER M1 ;
        RECT 5.756 13.404 5.788 15.912 ;
  LAYER M3 ;
        RECT 5.756 15.86 5.788 15.892 ;
  LAYER M1 ;
        RECT 5.82 13.404 5.852 15.912 ;
  LAYER M3 ;
        RECT 5.82 13.424 5.852 13.456 ;
  LAYER M1 ;
        RECT 5.884 13.404 5.916 15.912 ;
  LAYER M3 ;
        RECT 5.884 15.86 5.916 15.892 ;
  LAYER M1 ;
        RECT 5.948 13.404 5.98 15.912 ;
  LAYER M3 ;
        RECT 5.948 13.424 5.98 13.456 ;
  LAYER M1 ;
        RECT 6.012 13.404 6.044 15.912 ;
  LAYER M3 ;
        RECT 6.012 15.86 6.044 15.892 ;
  LAYER M1 ;
        RECT 6.076 13.404 6.108 15.912 ;
  LAYER M3 ;
        RECT 3.708 13.488 3.74 13.52 ;
  LAYER M2 ;
        RECT 6.076 13.552 6.108 13.584 ;
  LAYER M2 ;
        RECT 3.708 13.616 3.74 13.648 ;
  LAYER M2 ;
        RECT 6.076 13.68 6.108 13.712 ;
  LAYER M2 ;
        RECT 3.708 13.744 3.74 13.776 ;
  LAYER M2 ;
        RECT 6.076 13.808 6.108 13.84 ;
  LAYER M2 ;
        RECT 3.708 13.872 3.74 13.904 ;
  LAYER M2 ;
        RECT 6.076 13.936 6.108 13.968 ;
  LAYER M2 ;
        RECT 3.708 14 3.74 14.032 ;
  LAYER M2 ;
        RECT 6.076 14.064 6.108 14.096 ;
  LAYER M2 ;
        RECT 3.708 14.128 3.74 14.16 ;
  LAYER M2 ;
        RECT 6.076 14.192 6.108 14.224 ;
  LAYER M2 ;
        RECT 3.708 14.256 3.74 14.288 ;
  LAYER M2 ;
        RECT 6.076 14.32 6.108 14.352 ;
  LAYER M2 ;
        RECT 3.708 14.384 3.74 14.416 ;
  LAYER M2 ;
        RECT 6.076 14.448 6.108 14.48 ;
  LAYER M2 ;
        RECT 3.708 14.512 3.74 14.544 ;
  LAYER M2 ;
        RECT 6.076 14.576 6.108 14.608 ;
  LAYER M2 ;
        RECT 3.708 14.64 3.74 14.672 ;
  LAYER M2 ;
        RECT 6.076 14.704 6.108 14.736 ;
  LAYER M2 ;
        RECT 3.708 14.768 3.74 14.8 ;
  LAYER M2 ;
        RECT 6.076 14.832 6.108 14.864 ;
  LAYER M2 ;
        RECT 3.708 14.896 3.74 14.928 ;
  LAYER M2 ;
        RECT 6.076 14.96 6.108 14.992 ;
  LAYER M2 ;
        RECT 3.708 15.024 3.74 15.056 ;
  LAYER M2 ;
        RECT 6.076 15.088 6.108 15.12 ;
  LAYER M2 ;
        RECT 3.708 15.152 3.74 15.184 ;
  LAYER M2 ;
        RECT 6.076 15.216 6.108 15.248 ;
  LAYER M2 ;
        RECT 3.708 15.28 3.74 15.312 ;
  LAYER M2 ;
        RECT 6.076 15.344 6.108 15.376 ;
  LAYER M2 ;
        RECT 3.708 15.408 3.74 15.44 ;
  LAYER M2 ;
        RECT 6.076 15.472 6.108 15.504 ;
  LAYER M2 ;
        RECT 3.708 15.536 3.74 15.568 ;
  LAYER M2 ;
        RECT 6.076 15.6 6.108 15.632 ;
  LAYER M2 ;
        RECT 3.708 15.664 3.74 15.696 ;
  LAYER M2 ;
        RECT 6.076 15.728 6.108 15.76 ;
  LAYER M2 ;
        RECT 3.66 13.356 6.156 15.96 ;
  LAYER M1 ;
        RECT 3.708 16.512 3.74 19.02 ;
  LAYER M3 ;
        RECT 3.708 18.968 3.74 19 ;
  LAYER M1 ;
        RECT 3.772 16.512 3.804 19.02 ;
  LAYER M3 ;
        RECT 3.772 16.532 3.804 16.564 ;
  LAYER M1 ;
        RECT 3.836 16.512 3.868 19.02 ;
  LAYER M3 ;
        RECT 3.836 18.968 3.868 19 ;
  LAYER M1 ;
        RECT 3.9 16.512 3.932 19.02 ;
  LAYER M3 ;
        RECT 3.9 16.532 3.932 16.564 ;
  LAYER M1 ;
        RECT 3.964 16.512 3.996 19.02 ;
  LAYER M3 ;
        RECT 3.964 18.968 3.996 19 ;
  LAYER M1 ;
        RECT 4.028 16.512 4.06 19.02 ;
  LAYER M3 ;
        RECT 4.028 16.532 4.06 16.564 ;
  LAYER M1 ;
        RECT 4.092 16.512 4.124 19.02 ;
  LAYER M3 ;
        RECT 4.092 18.968 4.124 19 ;
  LAYER M1 ;
        RECT 4.156 16.512 4.188 19.02 ;
  LAYER M3 ;
        RECT 4.156 16.532 4.188 16.564 ;
  LAYER M1 ;
        RECT 4.22 16.512 4.252 19.02 ;
  LAYER M3 ;
        RECT 4.22 18.968 4.252 19 ;
  LAYER M1 ;
        RECT 4.284 16.512 4.316 19.02 ;
  LAYER M3 ;
        RECT 4.284 16.532 4.316 16.564 ;
  LAYER M1 ;
        RECT 4.348 16.512 4.38 19.02 ;
  LAYER M3 ;
        RECT 4.348 18.968 4.38 19 ;
  LAYER M1 ;
        RECT 4.412 16.512 4.444 19.02 ;
  LAYER M3 ;
        RECT 4.412 16.532 4.444 16.564 ;
  LAYER M1 ;
        RECT 4.476 16.512 4.508 19.02 ;
  LAYER M3 ;
        RECT 4.476 18.968 4.508 19 ;
  LAYER M1 ;
        RECT 4.54 16.512 4.572 19.02 ;
  LAYER M3 ;
        RECT 4.54 16.532 4.572 16.564 ;
  LAYER M1 ;
        RECT 4.604 16.512 4.636 19.02 ;
  LAYER M3 ;
        RECT 4.604 18.968 4.636 19 ;
  LAYER M1 ;
        RECT 4.668 16.512 4.7 19.02 ;
  LAYER M3 ;
        RECT 4.668 16.532 4.7 16.564 ;
  LAYER M1 ;
        RECT 4.732 16.512 4.764 19.02 ;
  LAYER M3 ;
        RECT 4.732 18.968 4.764 19 ;
  LAYER M1 ;
        RECT 4.796 16.512 4.828 19.02 ;
  LAYER M3 ;
        RECT 4.796 16.532 4.828 16.564 ;
  LAYER M1 ;
        RECT 4.86 16.512 4.892 19.02 ;
  LAYER M3 ;
        RECT 4.86 18.968 4.892 19 ;
  LAYER M1 ;
        RECT 4.924 16.512 4.956 19.02 ;
  LAYER M3 ;
        RECT 4.924 16.532 4.956 16.564 ;
  LAYER M1 ;
        RECT 4.988 16.512 5.02 19.02 ;
  LAYER M3 ;
        RECT 4.988 18.968 5.02 19 ;
  LAYER M1 ;
        RECT 5.052 16.512 5.084 19.02 ;
  LAYER M3 ;
        RECT 5.052 16.532 5.084 16.564 ;
  LAYER M1 ;
        RECT 5.116 16.512 5.148 19.02 ;
  LAYER M3 ;
        RECT 5.116 18.968 5.148 19 ;
  LAYER M1 ;
        RECT 5.18 16.512 5.212 19.02 ;
  LAYER M3 ;
        RECT 5.18 16.532 5.212 16.564 ;
  LAYER M1 ;
        RECT 5.244 16.512 5.276 19.02 ;
  LAYER M3 ;
        RECT 5.244 18.968 5.276 19 ;
  LAYER M1 ;
        RECT 5.308 16.512 5.34 19.02 ;
  LAYER M3 ;
        RECT 5.308 16.532 5.34 16.564 ;
  LAYER M1 ;
        RECT 5.372 16.512 5.404 19.02 ;
  LAYER M3 ;
        RECT 5.372 18.968 5.404 19 ;
  LAYER M1 ;
        RECT 5.436 16.512 5.468 19.02 ;
  LAYER M3 ;
        RECT 5.436 16.532 5.468 16.564 ;
  LAYER M1 ;
        RECT 5.5 16.512 5.532 19.02 ;
  LAYER M3 ;
        RECT 5.5 18.968 5.532 19 ;
  LAYER M1 ;
        RECT 5.564 16.512 5.596 19.02 ;
  LAYER M3 ;
        RECT 5.564 16.532 5.596 16.564 ;
  LAYER M1 ;
        RECT 5.628 16.512 5.66 19.02 ;
  LAYER M3 ;
        RECT 5.628 18.968 5.66 19 ;
  LAYER M1 ;
        RECT 5.692 16.512 5.724 19.02 ;
  LAYER M3 ;
        RECT 5.692 16.532 5.724 16.564 ;
  LAYER M1 ;
        RECT 5.756 16.512 5.788 19.02 ;
  LAYER M3 ;
        RECT 5.756 18.968 5.788 19 ;
  LAYER M1 ;
        RECT 5.82 16.512 5.852 19.02 ;
  LAYER M3 ;
        RECT 5.82 16.532 5.852 16.564 ;
  LAYER M1 ;
        RECT 5.884 16.512 5.916 19.02 ;
  LAYER M3 ;
        RECT 5.884 18.968 5.916 19 ;
  LAYER M1 ;
        RECT 5.948 16.512 5.98 19.02 ;
  LAYER M3 ;
        RECT 5.948 16.532 5.98 16.564 ;
  LAYER M1 ;
        RECT 6.012 16.512 6.044 19.02 ;
  LAYER M3 ;
        RECT 6.012 18.968 6.044 19 ;
  LAYER M1 ;
        RECT 6.076 16.512 6.108 19.02 ;
  LAYER M3 ;
        RECT 3.708 16.596 3.74 16.628 ;
  LAYER M2 ;
        RECT 6.076 16.66 6.108 16.692 ;
  LAYER M2 ;
        RECT 3.708 16.724 3.74 16.756 ;
  LAYER M2 ;
        RECT 6.076 16.788 6.108 16.82 ;
  LAYER M2 ;
        RECT 3.708 16.852 3.74 16.884 ;
  LAYER M2 ;
        RECT 6.076 16.916 6.108 16.948 ;
  LAYER M2 ;
        RECT 3.708 16.98 3.74 17.012 ;
  LAYER M2 ;
        RECT 6.076 17.044 6.108 17.076 ;
  LAYER M2 ;
        RECT 3.708 17.108 3.74 17.14 ;
  LAYER M2 ;
        RECT 6.076 17.172 6.108 17.204 ;
  LAYER M2 ;
        RECT 3.708 17.236 3.74 17.268 ;
  LAYER M2 ;
        RECT 6.076 17.3 6.108 17.332 ;
  LAYER M2 ;
        RECT 3.708 17.364 3.74 17.396 ;
  LAYER M2 ;
        RECT 6.076 17.428 6.108 17.46 ;
  LAYER M2 ;
        RECT 3.708 17.492 3.74 17.524 ;
  LAYER M2 ;
        RECT 6.076 17.556 6.108 17.588 ;
  LAYER M2 ;
        RECT 3.708 17.62 3.74 17.652 ;
  LAYER M2 ;
        RECT 6.076 17.684 6.108 17.716 ;
  LAYER M2 ;
        RECT 3.708 17.748 3.74 17.78 ;
  LAYER M2 ;
        RECT 6.076 17.812 6.108 17.844 ;
  LAYER M2 ;
        RECT 3.708 17.876 3.74 17.908 ;
  LAYER M2 ;
        RECT 6.076 17.94 6.108 17.972 ;
  LAYER M2 ;
        RECT 3.708 18.004 3.74 18.036 ;
  LAYER M2 ;
        RECT 6.076 18.068 6.108 18.1 ;
  LAYER M2 ;
        RECT 3.708 18.132 3.74 18.164 ;
  LAYER M2 ;
        RECT 6.076 18.196 6.108 18.228 ;
  LAYER M2 ;
        RECT 3.708 18.26 3.74 18.292 ;
  LAYER M2 ;
        RECT 6.076 18.324 6.108 18.356 ;
  LAYER M2 ;
        RECT 3.708 18.388 3.74 18.42 ;
  LAYER M2 ;
        RECT 6.076 18.452 6.108 18.484 ;
  LAYER M2 ;
        RECT 3.708 18.516 3.74 18.548 ;
  LAYER M2 ;
        RECT 6.076 18.58 6.108 18.612 ;
  LAYER M2 ;
        RECT 3.708 18.644 3.74 18.676 ;
  LAYER M2 ;
        RECT 6.076 18.708 6.108 18.74 ;
  LAYER M2 ;
        RECT 3.708 18.772 3.74 18.804 ;
  LAYER M2 ;
        RECT 6.076 18.836 6.108 18.868 ;
  LAYER M2 ;
        RECT 3.66 16.464 6.156 19.068 ;
  LAYER M1 ;
        RECT 7.324 0.972 7.356 3.48 ;
  LAYER M3 ;
        RECT 7.324 3.428 7.356 3.46 ;
  LAYER M1 ;
        RECT 7.388 0.972 7.42 3.48 ;
  LAYER M3 ;
        RECT 7.388 0.992 7.42 1.024 ;
  LAYER M1 ;
        RECT 7.452 0.972 7.484 3.48 ;
  LAYER M3 ;
        RECT 7.452 3.428 7.484 3.46 ;
  LAYER M1 ;
        RECT 7.516 0.972 7.548 3.48 ;
  LAYER M3 ;
        RECT 7.516 0.992 7.548 1.024 ;
  LAYER M1 ;
        RECT 7.58 0.972 7.612 3.48 ;
  LAYER M3 ;
        RECT 7.58 3.428 7.612 3.46 ;
  LAYER M1 ;
        RECT 7.644 0.972 7.676 3.48 ;
  LAYER M3 ;
        RECT 7.644 0.992 7.676 1.024 ;
  LAYER M1 ;
        RECT 7.708 0.972 7.74 3.48 ;
  LAYER M3 ;
        RECT 7.708 3.428 7.74 3.46 ;
  LAYER M1 ;
        RECT 7.772 0.972 7.804 3.48 ;
  LAYER M3 ;
        RECT 7.772 0.992 7.804 1.024 ;
  LAYER M1 ;
        RECT 7.836 0.972 7.868 3.48 ;
  LAYER M3 ;
        RECT 7.836 3.428 7.868 3.46 ;
  LAYER M1 ;
        RECT 7.9 0.972 7.932 3.48 ;
  LAYER M3 ;
        RECT 7.9 0.992 7.932 1.024 ;
  LAYER M1 ;
        RECT 7.964 0.972 7.996 3.48 ;
  LAYER M3 ;
        RECT 7.964 3.428 7.996 3.46 ;
  LAYER M1 ;
        RECT 8.028 0.972 8.06 3.48 ;
  LAYER M3 ;
        RECT 8.028 0.992 8.06 1.024 ;
  LAYER M1 ;
        RECT 8.092 0.972 8.124 3.48 ;
  LAYER M3 ;
        RECT 8.092 3.428 8.124 3.46 ;
  LAYER M1 ;
        RECT 8.156 0.972 8.188 3.48 ;
  LAYER M3 ;
        RECT 8.156 0.992 8.188 1.024 ;
  LAYER M1 ;
        RECT 8.22 0.972 8.252 3.48 ;
  LAYER M3 ;
        RECT 8.22 3.428 8.252 3.46 ;
  LAYER M1 ;
        RECT 8.284 0.972 8.316 3.48 ;
  LAYER M3 ;
        RECT 8.284 0.992 8.316 1.024 ;
  LAYER M1 ;
        RECT 8.348 0.972 8.38 3.48 ;
  LAYER M3 ;
        RECT 8.348 3.428 8.38 3.46 ;
  LAYER M1 ;
        RECT 8.412 0.972 8.444 3.48 ;
  LAYER M3 ;
        RECT 8.412 0.992 8.444 1.024 ;
  LAYER M1 ;
        RECT 8.476 0.972 8.508 3.48 ;
  LAYER M3 ;
        RECT 8.476 3.428 8.508 3.46 ;
  LAYER M1 ;
        RECT 8.54 0.972 8.572 3.48 ;
  LAYER M3 ;
        RECT 8.54 0.992 8.572 1.024 ;
  LAYER M1 ;
        RECT 8.604 0.972 8.636 3.48 ;
  LAYER M3 ;
        RECT 8.604 3.428 8.636 3.46 ;
  LAYER M1 ;
        RECT 8.668 0.972 8.7 3.48 ;
  LAYER M3 ;
        RECT 8.668 0.992 8.7 1.024 ;
  LAYER M1 ;
        RECT 8.732 0.972 8.764 3.48 ;
  LAYER M3 ;
        RECT 8.732 3.428 8.764 3.46 ;
  LAYER M1 ;
        RECT 8.796 0.972 8.828 3.48 ;
  LAYER M3 ;
        RECT 8.796 0.992 8.828 1.024 ;
  LAYER M1 ;
        RECT 8.86 0.972 8.892 3.48 ;
  LAYER M3 ;
        RECT 8.86 3.428 8.892 3.46 ;
  LAYER M1 ;
        RECT 8.924 0.972 8.956 3.48 ;
  LAYER M3 ;
        RECT 8.924 0.992 8.956 1.024 ;
  LAYER M1 ;
        RECT 8.988 0.972 9.02 3.48 ;
  LAYER M3 ;
        RECT 8.988 3.428 9.02 3.46 ;
  LAYER M1 ;
        RECT 9.052 0.972 9.084 3.48 ;
  LAYER M3 ;
        RECT 9.052 0.992 9.084 1.024 ;
  LAYER M1 ;
        RECT 9.116 0.972 9.148 3.48 ;
  LAYER M3 ;
        RECT 9.116 3.428 9.148 3.46 ;
  LAYER M1 ;
        RECT 9.18 0.972 9.212 3.48 ;
  LAYER M3 ;
        RECT 9.18 0.992 9.212 1.024 ;
  LAYER M1 ;
        RECT 9.244 0.972 9.276 3.48 ;
  LAYER M3 ;
        RECT 9.244 3.428 9.276 3.46 ;
  LAYER M1 ;
        RECT 9.308 0.972 9.34 3.48 ;
  LAYER M3 ;
        RECT 9.308 0.992 9.34 1.024 ;
  LAYER M1 ;
        RECT 9.372 0.972 9.404 3.48 ;
  LAYER M3 ;
        RECT 9.372 3.428 9.404 3.46 ;
  LAYER M1 ;
        RECT 9.436 0.972 9.468 3.48 ;
  LAYER M3 ;
        RECT 9.436 0.992 9.468 1.024 ;
  LAYER M1 ;
        RECT 9.5 0.972 9.532 3.48 ;
  LAYER M3 ;
        RECT 9.5 3.428 9.532 3.46 ;
  LAYER M1 ;
        RECT 9.564 0.972 9.596 3.48 ;
  LAYER M3 ;
        RECT 9.564 0.992 9.596 1.024 ;
  LAYER M1 ;
        RECT 9.628 0.972 9.66 3.48 ;
  LAYER M3 ;
        RECT 9.628 3.428 9.66 3.46 ;
  LAYER M1 ;
        RECT 9.692 0.972 9.724 3.48 ;
  LAYER M3 ;
        RECT 7.324 1.056 7.356 1.088 ;
  LAYER M2 ;
        RECT 9.692 1.12 9.724 1.152 ;
  LAYER M2 ;
        RECT 7.324 1.184 7.356 1.216 ;
  LAYER M2 ;
        RECT 9.692 1.248 9.724 1.28 ;
  LAYER M2 ;
        RECT 7.324 1.312 7.356 1.344 ;
  LAYER M2 ;
        RECT 9.692 1.376 9.724 1.408 ;
  LAYER M2 ;
        RECT 7.324 1.44 7.356 1.472 ;
  LAYER M2 ;
        RECT 9.692 1.504 9.724 1.536 ;
  LAYER M2 ;
        RECT 7.324 1.568 7.356 1.6 ;
  LAYER M2 ;
        RECT 9.692 1.632 9.724 1.664 ;
  LAYER M2 ;
        RECT 7.324 1.696 7.356 1.728 ;
  LAYER M2 ;
        RECT 9.692 1.76 9.724 1.792 ;
  LAYER M2 ;
        RECT 7.324 1.824 7.356 1.856 ;
  LAYER M2 ;
        RECT 9.692 1.888 9.724 1.92 ;
  LAYER M2 ;
        RECT 7.324 1.952 7.356 1.984 ;
  LAYER M2 ;
        RECT 9.692 2.016 9.724 2.048 ;
  LAYER M2 ;
        RECT 7.324 2.08 7.356 2.112 ;
  LAYER M2 ;
        RECT 9.692 2.144 9.724 2.176 ;
  LAYER M2 ;
        RECT 7.324 2.208 7.356 2.24 ;
  LAYER M2 ;
        RECT 9.692 2.272 9.724 2.304 ;
  LAYER M2 ;
        RECT 7.324 2.336 7.356 2.368 ;
  LAYER M2 ;
        RECT 9.692 2.4 9.724 2.432 ;
  LAYER M2 ;
        RECT 7.324 2.464 7.356 2.496 ;
  LAYER M2 ;
        RECT 9.692 2.528 9.724 2.56 ;
  LAYER M2 ;
        RECT 7.324 2.592 7.356 2.624 ;
  LAYER M2 ;
        RECT 9.692 2.656 9.724 2.688 ;
  LAYER M2 ;
        RECT 7.324 2.72 7.356 2.752 ;
  LAYER M2 ;
        RECT 9.692 2.784 9.724 2.816 ;
  LAYER M2 ;
        RECT 7.324 2.848 7.356 2.88 ;
  LAYER M2 ;
        RECT 9.692 2.912 9.724 2.944 ;
  LAYER M2 ;
        RECT 7.324 2.976 7.356 3.008 ;
  LAYER M2 ;
        RECT 9.692 3.04 9.724 3.072 ;
  LAYER M2 ;
        RECT 7.324 3.104 7.356 3.136 ;
  LAYER M2 ;
        RECT 9.692 3.168 9.724 3.2 ;
  LAYER M2 ;
        RECT 7.324 3.232 7.356 3.264 ;
  LAYER M2 ;
        RECT 9.692 3.296 9.724 3.328 ;
  LAYER M2 ;
        RECT 7.276 0.924 9.772 3.528 ;
  LAYER M1 ;
        RECT 7.324 4.08 7.356 6.588 ;
  LAYER M3 ;
        RECT 7.324 6.536 7.356 6.568 ;
  LAYER M1 ;
        RECT 7.388 4.08 7.42 6.588 ;
  LAYER M3 ;
        RECT 7.388 4.1 7.42 4.132 ;
  LAYER M1 ;
        RECT 7.452 4.08 7.484 6.588 ;
  LAYER M3 ;
        RECT 7.452 6.536 7.484 6.568 ;
  LAYER M1 ;
        RECT 7.516 4.08 7.548 6.588 ;
  LAYER M3 ;
        RECT 7.516 4.1 7.548 4.132 ;
  LAYER M1 ;
        RECT 7.58 4.08 7.612 6.588 ;
  LAYER M3 ;
        RECT 7.58 6.536 7.612 6.568 ;
  LAYER M1 ;
        RECT 7.644 4.08 7.676 6.588 ;
  LAYER M3 ;
        RECT 7.644 4.1 7.676 4.132 ;
  LAYER M1 ;
        RECT 7.708 4.08 7.74 6.588 ;
  LAYER M3 ;
        RECT 7.708 6.536 7.74 6.568 ;
  LAYER M1 ;
        RECT 7.772 4.08 7.804 6.588 ;
  LAYER M3 ;
        RECT 7.772 4.1 7.804 4.132 ;
  LAYER M1 ;
        RECT 7.836 4.08 7.868 6.588 ;
  LAYER M3 ;
        RECT 7.836 6.536 7.868 6.568 ;
  LAYER M1 ;
        RECT 7.9 4.08 7.932 6.588 ;
  LAYER M3 ;
        RECT 7.9 4.1 7.932 4.132 ;
  LAYER M1 ;
        RECT 7.964 4.08 7.996 6.588 ;
  LAYER M3 ;
        RECT 7.964 6.536 7.996 6.568 ;
  LAYER M1 ;
        RECT 8.028 4.08 8.06 6.588 ;
  LAYER M3 ;
        RECT 8.028 4.1 8.06 4.132 ;
  LAYER M1 ;
        RECT 8.092 4.08 8.124 6.588 ;
  LAYER M3 ;
        RECT 8.092 6.536 8.124 6.568 ;
  LAYER M1 ;
        RECT 8.156 4.08 8.188 6.588 ;
  LAYER M3 ;
        RECT 8.156 4.1 8.188 4.132 ;
  LAYER M1 ;
        RECT 8.22 4.08 8.252 6.588 ;
  LAYER M3 ;
        RECT 8.22 6.536 8.252 6.568 ;
  LAYER M1 ;
        RECT 8.284 4.08 8.316 6.588 ;
  LAYER M3 ;
        RECT 8.284 4.1 8.316 4.132 ;
  LAYER M1 ;
        RECT 8.348 4.08 8.38 6.588 ;
  LAYER M3 ;
        RECT 8.348 6.536 8.38 6.568 ;
  LAYER M1 ;
        RECT 8.412 4.08 8.444 6.588 ;
  LAYER M3 ;
        RECT 8.412 4.1 8.444 4.132 ;
  LAYER M1 ;
        RECT 8.476 4.08 8.508 6.588 ;
  LAYER M3 ;
        RECT 8.476 6.536 8.508 6.568 ;
  LAYER M1 ;
        RECT 8.54 4.08 8.572 6.588 ;
  LAYER M3 ;
        RECT 8.54 4.1 8.572 4.132 ;
  LAYER M1 ;
        RECT 8.604 4.08 8.636 6.588 ;
  LAYER M3 ;
        RECT 8.604 6.536 8.636 6.568 ;
  LAYER M1 ;
        RECT 8.668 4.08 8.7 6.588 ;
  LAYER M3 ;
        RECT 8.668 4.1 8.7 4.132 ;
  LAYER M1 ;
        RECT 8.732 4.08 8.764 6.588 ;
  LAYER M3 ;
        RECT 8.732 6.536 8.764 6.568 ;
  LAYER M1 ;
        RECT 8.796 4.08 8.828 6.588 ;
  LAYER M3 ;
        RECT 8.796 4.1 8.828 4.132 ;
  LAYER M1 ;
        RECT 8.86 4.08 8.892 6.588 ;
  LAYER M3 ;
        RECT 8.86 6.536 8.892 6.568 ;
  LAYER M1 ;
        RECT 8.924 4.08 8.956 6.588 ;
  LAYER M3 ;
        RECT 8.924 4.1 8.956 4.132 ;
  LAYER M1 ;
        RECT 8.988 4.08 9.02 6.588 ;
  LAYER M3 ;
        RECT 8.988 6.536 9.02 6.568 ;
  LAYER M1 ;
        RECT 9.052 4.08 9.084 6.588 ;
  LAYER M3 ;
        RECT 9.052 4.1 9.084 4.132 ;
  LAYER M1 ;
        RECT 9.116 4.08 9.148 6.588 ;
  LAYER M3 ;
        RECT 9.116 6.536 9.148 6.568 ;
  LAYER M1 ;
        RECT 9.18 4.08 9.212 6.588 ;
  LAYER M3 ;
        RECT 9.18 4.1 9.212 4.132 ;
  LAYER M1 ;
        RECT 9.244 4.08 9.276 6.588 ;
  LAYER M3 ;
        RECT 9.244 6.536 9.276 6.568 ;
  LAYER M1 ;
        RECT 9.308 4.08 9.34 6.588 ;
  LAYER M3 ;
        RECT 9.308 4.1 9.34 4.132 ;
  LAYER M1 ;
        RECT 9.372 4.08 9.404 6.588 ;
  LAYER M3 ;
        RECT 9.372 6.536 9.404 6.568 ;
  LAYER M1 ;
        RECT 9.436 4.08 9.468 6.588 ;
  LAYER M3 ;
        RECT 9.436 4.1 9.468 4.132 ;
  LAYER M1 ;
        RECT 9.5 4.08 9.532 6.588 ;
  LAYER M3 ;
        RECT 9.5 6.536 9.532 6.568 ;
  LAYER M1 ;
        RECT 9.564 4.08 9.596 6.588 ;
  LAYER M3 ;
        RECT 9.564 4.1 9.596 4.132 ;
  LAYER M1 ;
        RECT 9.628 4.08 9.66 6.588 ;
  LAYER M3 ;
        RECT 9.628 6.536 9.66 6.568 ;
  LAYER M1 ;
        RECT 9.692 4.08 9.724 6.588 ;
  LAYER M3 ;
        RECT 7.324 4.164 7.356 4.196 ;
  LAYER M2 ;
        RECT 9.692 4.228 9.724 4.26 ;
  LAYER M2 ;
        RECT 7.324 4.292 7.356 4.324 ;
  LAYER M2 ;
        RECT 9.692 4.356 9.724 4.388 ;
  LAYER M2 ;
        RECT 7.324 4.42 7.356 4.452 ;
  LAYER M2 ;
        RECT 9.692 4.484 9.724 4.516 ;
  LAYER M2 ;
        RECT 7.324 4.548 7.356 4.58 ;
  LAYER M2 ;
        RECT 9.692 4.612 9.724 4.644 ;
  LAYER M2 ;
        RECT 7.324 4.676 7.356 4.708 ;
  LAYER M2 ;
        RECT 9.692 4.74 9.724 4.772 ;
  LAYER M2 ;
        RECT 7.324 4.804 7.356 4.836 ;
  LAYER M2 ;
        RECT 9.692 4.868 9.724 4.9 ;
  LAYER M2 ;
        RECT 7.324 4.932 7.356 4.964 ;
  LAYER M2 ;
        RECT 9.692 4.996 9.724 5.028 ;
  LAYER M2 ;
        RECT 7.324 5.06 7.356 5.092 ;
  LAYER M2 ;
        RECT 9.692 5.124 9.724 5.156 ;
  LAYER M2 ;
        RECT 7.324 5.188 7.356 5.22 ;
  LAYER M2 ;
        RECT 9.692 5.252 9.724 5.284 ;
  LAYER M2 ;
        RECT 7.324 5.316 7.356 5.348 ;
  LAYER M2 ;
        RECT 9.692 5.38 9.724 5.412 ;
  LAYER M2 ;
        RECT 7.324 5.444 7.356 5.476 ;
  LAYER M2 ;
        RECT 9.692 5.508 9.724 5.54 ;
  LAYER M2 ;
        RECT 7.324 5.572 7.356 5.604 ;
  LAYER M2 ;
        RECT 9.692 5.636 9.724 5.668 ;
  LAYER M2 ;
        RECT 7.324 5.7 7.356 5.732 ;
  LAYER M2 ;
        RECT 9.692 5.764 9.724 5.796 ;
  LAYER M2 ;
        RECT 7.324 5.828 7.356 5.86 ;
  LAYER M2 ;
        RECT 9.692 5.892 9.724 5.924 ;
  LAYER M2 ;
        RECT 7.324 5.956 7.356 5.988 ;
  LAYER M2 ;
        RECT 9.692 6.02 9.724 6.052 ;
  LAYER M2 ;
        RECT 7.324 6.084 7.356 6.116 ;
  LAYER M2 ;
        RECT 9.692 6.148 9.724 6.18 ;
  LAYER M2 ;
        RECT 7.324 6.212 7.356 6.244 ;
  LAYER M2 ;
        RECT 9.692 6.276 9.724 6.308 ;
  LAYER M2 ;
        RECT 7.324 6.34 7.356 6.372 ;
  LAYER M2 ;
        RECT 9.692 6.404 9.724 6.436 ;
  LAYER M2 ;
        RECT 7.276 4.032 9.772 6.636 ;
  LAYER M1 ;
        RECT 7.324 7.188 7.356 9.696 ;
  LAYER M3 ;
        RECT 7.324 9.644 7.356 9.676 ;
  LAYER M1 ;
        RECT 7.388 7.188 7.42 9.696 ;
  LAYER M3 ;
        RECT 7.388 7.208 7.42 7.24 ;
  LAYER M1 ;
        RECT 7.452 7.188 7.484 9.696 ;
  LAYER M3 ;
        RECT 7.452 9.644 7.484 9.676 ;
  LAYER M1 ;
        RECT 7.516 7.188 7.548 9.696 ;
  LAYER M3 ;
        RECT 7.516 7.208 7.548 7.24 ;
  LAYER M1 ;
        RECT 7.58 7.188 7.612 9.696 ;
  LAYER M3 ;
        RECT 7.58 9.644 7.612 9.676 ;
  LAYER M1 ;
        RECT 7.644 7.188 7.676 9.696 ;
  LAYER M3 ;
        RECT 7.644 7.208 7.676 7.24 ;
  LAYER M1 ;
        RECT 7.708 7.188 7.74 9.696 ;
  LAYER M3 ;
        RECT 7.708 9.644 7.74 9.676 ;
  LAYER M1 ;
        RECT 7.772 7.188 7.804 9.696 ;
  LAYER M3 ;
        RECT 7.772 7.208 7.804 7.24 ;
  LAYER M1 ;
        RECT 7.836 7.188 7.868 9.696 ;
  LAYER M3 ;
        RECT 7.836 9.644 7.868 9.676 ;
  LAYER M1 ;
        RECT 7.9 7.188 7.932 9.696 ;
  LAYER M3 ;
        RECT 7.9 7.208 7.932 7.24 ;
  LAYER M1 ;
        RECT 7.964 7.188 7.996 9.696 ;
  LAYER M3 ;
        RECT 7.964 9.644 7.996 9.676 ;
  LAYER M1 ;
        RECT 8.028 7.188 8.06 9.696 ;
  LAYER M3 ;
        RECT 8.028 7.208 8.06 7.24 ;
  LAYER M1 ;
        RECT 8.092 7.188 8.124 9.696 ;
  LAYER M3 ;
        RECT 8.092 9.644 8.124 9.676 ;
  LAYER M1 ;
        RECT 8.156 7.188 8.188 9.696 ;
  LAYER M3 ;
        RECT 8.156 7.208 8.188 7.24 ;
  LAYER M1 ;
        RECT 8.22 7.188 8.252 9.696 ;
  LAYER M3 ;
        RECT 8.22 9.644 8.252 9.676 ;
  LAYER M1 ;
        RECT 8.284 7.188 8.316 9.696 ;
  LAYER M3 ;
        RECT 8.284 7.208 8.316 7.24 ;
  LAYER M1 ;
        RECT 8.348 7.188 8.38 9.696 ;
  LAYER M3 ;
        RECT 8.348 9.644 8.38 9.676 ;
  LAYER M1 ;
        RECT 8.412 7.188 8.444 9.696 ;
  LAYER M3 ;
        RECT 8.412 7.208 8.444 7.24 ;
  LAYER M1 ;
        RECT 8.476 7.188 8.508 9.696 ;
  LAYER M3 ;
        RECT 8.476 9.644 8.508 9.676 ;
  LAYER M1 ;
        RECT 8.54 7.188 8.572 9.696 ;
  LAYER M3 ;
        RECT 8.54 7.208 8.572 7.24 ;
  LAYER M1 ;
        RECT 8.604 7.188 8.636 9.696 ;
  LAYER M3 ;
        RECT 8.604 9.644 8.636 9.676 ;
  LAYER M1 ;
        RECT 8.668 7.188 8.7 9.696 ;
  LAYER M3 ;
        RECT 8.668 7.208 8.7 7.24 ;
  LAYER M1 ;
        RECT 8.732 7.188 8.764 9.696 ;
  LAYER M3 ;
        RECT 8.732 9.644 8.764 9.676 ;
  LAYER M1 ;
        RECT 8.796 7.188 8.828 9.696 ;
  LAYER M3 ;
        RECT 8.796 7.208 8.828 7.24 ;
  LAYER M1 ;
        RECT 8.86 7.188 8.892 9.696 ;
  LAYER M3 ;
        RECT 8.86 9.644 8.892 9.676 ;
  LAYER M1 ;
        RECT 8.924 7.188 8.956 9.696 ;
  LAYER M3 ;
        RECT 8.924 7.208 8.956 7.24 ;
  LAYER M1 ;
        RECT 8.988 7.188 9.02 9.696 ;
  LAYER M3 ;
        RECT 8.988 9.644 9.02 9.676 ;
  LAYER M1 ;
        RECT 9.052 7.188 9.084 9.696 ;
  LAYER M3 ;
        RECT 9.052 7.208 9.084 7.24 ;
  LAYER M1 ;
        RECT 9.116 7.188 9.148 9.696 ;
  LAYER M3 ;
        RECT 9.116 9.644 9.148 9.676 ;
  LAYER M1 ;
        RECT 9.18 7.188 9.212 9.696 ;
  LAYER M3 ;
        RECT 9.18 7.208 9.212 7.24 ;
  LAYER M1 ;
        RECT 9.244 7.188 9.276 9.696 ;
  LAYER M3 ;
        RECT 9.244 9.644 9.276 9.676 ;
  LAYER M1 ;
        RECT 9.308 7.188 9.34 9.696 ;
  LAYER M3 ;
        RECT 9.308 7.208 9.34 7.24 ;
  LAYER M1 ;
        RECT 9.372 7.188 9.404 9.696 ;
  LAYER M3 ;
        RECT 9.372 9.644 9.404 9.676 ;
  LAYER M1 ;
        RECT 9.436 7.188 9.468 9.696 ;
  LAYER M3 ;
        RECT 9.436 7.208 9.468 7.24 ;
  LAYER M1 ;
        RECT 9.5 7.188 9.532 9.696 ;
  LAYER M3 ;
        RECT 9.5 9.644 9.532 9.676 ;
  LAYER M1 ;
        RECT 9.564 7.188 9.596 9.696 ;
  LAYER M3 ;
        RECT 9.564 7.208 9.596 7.24 ;
  LAYER M1 ;
        RECT 9.628 7.188 9.66 9.696 ;
  LAYER M3 ;
        RECT 9.628 9.644 9.66 9.676 ;
  LAYER M1 ;
        RECT 9.692 7.188 9.724 9.696 ;
  LAYER M3 ;
        RECT 7.324 7.272 7.356 7.304 ;
  LAYER M2 ;
        RECT 9.692 7.336 9.724 7.368 ;
  LAYER M2 ;
        RECT 7.324 7.4 7.356 7.432 ;
  LAYER M2 ;
        RECT 9.692 7.464 9.724 7.496 ;
  LAYER M2 ;
        RECT 7.324 7.528 7.356 7.56 ;
  LAYER M2 ;
        RECT 9.692 7.592 9.724 7.624 ;
  LAYER M2 ;
        RECT 7.324 7.656 7.356 7.688 ;
  LAYER M2 ;
        RECT 9.692 7.72 9.724 7.752 ;
  LAYER M2 ;
        RECT 7.324 7.784 7.356 7.816 ;
  LAYER M2 ;
        RECT 9.692 7.848 9.724 7.88 ;
  LAYER M2 ;
        RECT 7.324 7.912 7.356 7.944 ;
  LAYER M2 ;
        RECT 9.692 7.976 9.724 8.008 ;
  LAYER M2 ;
        RECT 7.324 8.04 7.356 8.072 ;
  LAYER M2 ;
        RECT 9.692 8.104 9.724 8.136 ;
  LAYER M2 ;
        RECT 7.324 8.168 7.356 8.2 ;
  LAYER M2 ;
        RECT 9.692 8.232 9.724 8.264 ;
  LAYER M2 ;
        RECT 7.324 8.296 7.356 8.328 ;
  LAYER M2 ;
        RECT 9.692 8.36 9.724 8.392 ;
  LAYER M2 ;
        RECT 7.324 8.424 7.356 8.456 ;
  LAYER M2 ;
        RECT 9.692 8.488 9.724 8.52 ;
  LAYER M2 ;
        RECT 7.324 8.552 7.356 8.584 ;
  LAYER M2 ;
        RECT 9.692 8.616 9.724 8.648 ;
  LAYER M2 ;
        RECT 7.324 8.68 7.356 8.712 ;
  LAYER M2 ;
        RECT 9.692 8.744 9.724 8.776 ;
  LAYER M2 ;
        RECT 7.324 8.808 7.356 8.84 ;
  LAYER M2 ;
        RECT 9.692 8.872 9.724 8.904 ;
  LAYER M2 ;
        RECT 7.324 8.936 7.356 8.968 ;
  LAYER M2 ;
        RECT 9.692 9 9.724 9.032 ;
  LAYER M2 ;
        RECT 7.324 9.064 7.356 9.096 ;
  LAYER M2 ;
        RECT 9.692 9.128 9.724 9.16 ;
  LAYER M2 ;
        RECT 7.324 9.192 7.356 9.224 ;
  LAYER M2 ;
        RECT 9.692 9.256 9.724 9.288 ;
  LAYER M2 ;
        RECT 7.324 9.32 7.356 9.352 ;
  LAYER M2 ;
        RECT 9.692 9.384 9.724 9.416 ;
  LAYER M2 ;
        RECT 7.324 9.448 7.356 9.48 ;
  LAYER M2 ;
        RECT 9.692 9.512 9.724 9.544 ;
  LAYER M2 ;
        RECT 7.276 7.14 9.772 9.744 ;
  LAYER M1 ;
        RECT 7.324 10.296 7.356 12.804 ;
  LAYER M3 ;
        RECT 7.324 12.752 7.356 12.784 ;
  LAYER M1 ;
        RECT 7.388 10.296 7.42 12.804 ;
  LAYER M3 ;
        RECT 7.388 10.316 7.42 10.348 ;
  LAYER M1 ;
        RECT 7.452 10.296 7.484 12.804 ;
  LAYER M3 ;
        RECT 7.452 12.752 7.484 12.784 ;
  LAYER M1 ;
        RECT 7.516 10.296 7.548 12.804 ;
  LAYER M3 ;
        RECT 7.516 10.316 7.548 10.348 ;
  LAYER M1 ;
        RECT 7.58 10.296 7.612 12.804 ;
  LAYER M3 ;
        RECT 7.58 12.752 7.612 12.784 ;
  LAYER M1 ;
        RECT 7.644 10.296 7.676 12.804 ;
  LAYER M3 ;
        RECT 7.644 10.316 7.676 10.348 ;
  LAYER M1 ;
        RECT 7.708 10.296 7.74 12.804 ;
  LAYER M3 ;
        RECT 7.708 12.752 7.74 12.784 ;
  LAYER M1 ;
        RECT 7.772 10.296 7.804 12.804 ;
  LAYER M3 ;
        RECT 7.772 10.316 7.804 10.348 ;
  LAYER M1 ;
        RECT 7.836 10.296 7.868 12.804 ;
  LAYER M3 ;
        RECT 7.836 12.752 7.868 12.784 ;
  LAYER M1 ;
        RECT 7.9 10.296 7.932 12.804 ;
  LAYER M3 ;
        RECT 7.9 10.316 7.932 10.348 ;
  LAYER M1 ;
        RECT 7.964 10.296 7.996 12.804 ;
  LAYER M3 ;
        RECT 7.964 12.752 7.996 12.784 ;
  LAYER M1 ;
        RECT 8.028 10.296 8.06 12.804 ;
  LAYER M3 ;
        RECT 8.028 10.316 8.06 10.348 ;
  LAYER M1 ;
        RECT 8.092 10.296 8.124 12.804 ;
  LAYER M3 ;
        RECT 8.092 12.752 8.124 12.784 ;
  LAYER M1 ;
        RECT 8.156 10.296 8.188 12.804 ;
  LAYER M3 ;
        RECT 8.156 10.316 8.188 10.348 ;
  LAYER M1 ;
        RECT 8.22 10.296 8.252 12.804 ;
  LAYER M3 ;
        RECT 8.22 12.752 8.252 12.784 ;
  LAYER M1 ;
        RECT 8.284 10.296 8.316 12.804 ;
  LAYER M3 ;
        RECT 8.284 10.316 8.316 10.348 ;
  LAYER M1 ;
        RECT 8.348 10.296 8.38 12.804 ;
  LAYER M3 ;
        RECT 8.348 12.752 8.38 12.784 ;
  LAYER M1 ;
        RECT 8.412 10.296 8.444 12.804 ;
  LAYER M3 ;
        RECT 8.412 10.316 8.444 10.348 ;
  LAYER M1 ;
        RECT 8.476 10.296 8.508 12.804 ;
  LAYER M3 ;
        RECT 8.476 12.752 8.508 12.784 ;
  LAYER M1 ;
        RECT 8.54 10.296 8.572 12.804 ;
  LAYER M3 ;
        RECT 8.54 10.316 8.572 10.348 ;
  LAYER M1 ;
        RECT 8.604 10.296 8.636 12.804 ;
  LAYER M3 ;
        RECT 8.604 12.752 8.636 12.784 ;
  LAYER M1 ;
        RECT 8.668 10.296 8.7 12.804 ;
  LAYER M3 ;
        RECT 8.668 10.316 8.7 10.348 ;
  LAYER M1 ;
        RECT 8.732 10.296 8.764 12.804 ;
  LAYER M3 ;
        RECT 8.732 12.752 8.764 12.784 ;
  LAYER M1 ;
        RECT 8.796 10.296 8.828 12.804 ;
  LAYER M3 ;
        RECT 8.796 10.316 8.828 10.348 ;
  LAYER M1 ;
        RECT 8.86 10.296 8.892 12.804 ;
  LAYER M3 ;
        RECT 8.86 12.752 8.892 12.784 ;
  LAYER M1 ;
        RECT 8.924 10.296 8.956 12.804 ;
  LAYER M3 ;
        RECT 8.924 10.316 8.956 10.348 ;
  LAYER M1 ;
        RECT 8.988 10.296 9.02 12.804 ;
  LAYER M3 ;
        RECT 8.988 12.752 9.02 12.784 ;
  LAYER M1 ;
        RECT 9.052 10.296 9.084 12.804 ;
  LAYER M3 ;
        RECT 9.052 10.316 9.084 10.348 ;
  LAYER M1 ;
        RECT 9.116 10.296 9.148 12.804 ;
  LAYER M3 ;
        RECT 9.116 12.752 9.148 12.784 ;
  LAYER M1 ;
        RECT 9.18 10.296 9.212 12.804 ;
  LAYER M3 ;
        RECT 9.18 10.316 9.212 10.348 ;
  LAYER M1 ;
        RECT 9.244 10.296 9.276 12.804 ;
  LAYER M3 ;
        RECT 9.244 12.752 9.276 12.784 ;
  LAYER M1 ;
        RECT 9.308 10.296 9.34 12.804 ;
  LAYER M3 ;
        RECT 9.308 10.316 9.34 10.348 ;
  LAYER M1 ;
        RECT 9.372 10.296 9.404 12.804 ;
  LAYER M3 ;
        RECT 9.372 12.752 9.404 12.784 ;
  LAYER M1 ;
        RECT 9.436 10.296 9.468 12.804 ;
  LAYER M3 ;
        RECT 9.436 10.316 9.468 10.348 ;
  LAYER M1 ;
        RECT 9.5 10.296 9.532 12.804 ;
  LAYER M3 ;
        RECT 9.5 12.752 9.532 12.784 ;
  LAYER M1 ;
        RECT 9.564 10.296 9.596 12.804 ;
  LAYER M3 ;
        RECT 9.564 10.316 9.596 10.348 ;
  LAYER M1 ;
        RECT 9.628 10.296 9.66 12.804 ;
  LAYER M3 ;
        RECT 9.628 12.752 9.66 12.784 ;
  LAYER M1 ;
        RECT 9.692 10.296 9.724 12.804 ;
  LAYER M3 ;
        RECT 7.324 10.38 7.356 10.412 ;
  LAYER M2 ;
        RECT 9.692 10.444 9.724 10.476 ;
  LAYER M2 ;
        RECT 7.324 10.508 7.356 10.54 ;
  LAYER M2 ;
        RECT 9.692 10.572 9.724 10.604 ;
  LAYER M2 ;
        RECT 7.324 10.636 7.356 10.668 ;
  LAYER M2 ;
        RECT 9.692 10.7 9.724 10.732 ;
  LAYER M2 ;
        RECT 7.324 10.764 7.356 10.796 ;
  LAYER M2 ;
        RECT 9.692 10.828 9.724 10.86 ;
  LAYER M2 ;
        RECT 7.324 10.892 7.356 10.924 ;
  LAYER M2 ;
        RECT 9.692 10.956 9.724 10.988 ;
  LAYER M2 ;
        RECT 7.324 11.02 7.356 11.052 ;
  LAYER M2 ;
        RECT 9.692 11.084 9.724 11.116 ;
  LAYER M2 ;
        RECT 7.324 11.148 7.356 11.18 ;
  LAYER M2 ;
        RECT 9.692 11.212 9.724 11.244 ;
  LAYER M2 ;
        RECT 7.324 11.276 7.356 11.308 ;
  LAYER M2 ;
        RECT 9.692 11.34 9.724 11.372 ;
  LAYER M2 ;
        RECT 7.324 11.404 7.356 11.436 ;
  LAYER M2 ;
        RECT 9.692 11.468 9.724 11.5 ;
  LAYER M2 ;
        RECT 7.324 11.532 7.356 11.564 ;
  LAYER M2 ;
        RECT 9.692 11.596 9.724 11.628 ;
  LAYER M2 ;
        RECT 7.324 11.66 7.356 11.692 ;
  LAYER M2 ;
        RECT 9.692 11.724 9.724 11.756 ;
  LAYER M2 ;
        RECT 7.324 11.788 7.356 11.82 ;
  LAYER M2 ;
        RECT 9.692 11.852 9.724 11.884 ;
  LAYER M2 ;
        RECT 7.324 11.916 7.356 11.948 ;
  LAYER M2 ;
        RECT 9.692 11.98 9.724 12.012 ;
  LAYER M2 ;
        RECT 7.324 12.044 7.356 12.076 ;
  LAYER M2 ;
        RECT 9.692 12.108 9.724 12.14 ;
  LAYER M2 ;
        RECT 7.324 12.172 7.356 12.204 ;
  LAYER M2 ;
        RECT 9.692 12.236 9.724 12.268 ;
  LAYER M2 ;
        RECT 7.324 12.3 7.356 12.332 ;
  LAYER M2 ;
        RECT 9.692 12.364 9.724 12.396 ;
  LAYER M2 ;
        RECT 7.324 12.428 7.356 12.46 ;
  LAYER M2 ;
        RECT 9.692 12.492 9.724 12.524 ;
  LAYER M2 ;
        RECT 7.324 12.556 7.356 12.588 ;
  LAYER M2 ;
        RECT 9.692 12.62 9.724 12.652 ;
  LAYER M2 ;
        RECT 7.276 10.248 9.772 12.852 ;
  LAYER M1 ;
        RECT 7.324 13.404 7.356 15.912 ;
  LAYER M3 ;
        RECT 7.324 15.86 7.356 15.892 ;
  LAYER M1 ;
        RECT 7.388 13.404 7.42 15.912 ;
  LAYER M3 ;
        RECT 7.388 13.424 7.42 13.456 ;
  LAYER M1 ;
        RECT 7.452 13.404 7.484 15.912 ;
  LAYER M3 ;
        RECT 7.452 15.86 7.484 15.892 ;
  LAYER M1 ;
        RECT 7.516 13.404 7.548 15.912 ;
  LAYER M3 ;
        RECT 7.516 13.424 7.548 13.456 ;
  LAYER M1 ;
        RECT 7.58 13.404 7.612 15.912 ;
  LAYER M3 ;
        RECT 7.58 15.86 7.612 15.892 ;
  LAYER M1 ;
        RECT 7.644 13.404 7.676 15.912 ;
  LAYER M3 ;
        RECT 7.644 13.424 7.676 13.456 ;
  LAYER M1 ;
        RECT 7.708 13.404 7.74 15.912 ;
  LAYER M3 ;
        RECT 7.708 15.86 7.74 15.892 ;
  LAYER M1 ;
        RECT 7.772 13.404 7.804 15.912 ;
  LAYER M3 ;
        RECT 7.772 13.424 7.804 13.456 ;
  LAYER M1 ;
        RECT 7.836 13.404 7.868 15.912 ;
  LAYER M3 ;
        RECT 7.836 15.86 7.868 15.892 ;
  LAYER M1 ;
        RECT 7.9 13.404 7.932 15.912 ;
  LAYER M3 ;
        RECT 7.9 13.424 7.932 13.456 ;
  LAYER M1 ;
        RECT 7.964 13.404 7.996 15.912 ;
  LAYER M3 ;
        RECT 7.964 15.86 7.996 15.892 ;
  LAYER M1 ;
        RECT 8.028 13.404 8.06 15.912 ;
  LAYER M3 ;
        RECT 8.028 13.424 8.06 13.456 ;
  LAYER M1 ;
        RECT 8.092 13.404 8.124 15.912 ;
  LAYER M3 ;
        RECT 8.092 15.86 8.124 15.892 ;
  LAYER M1 ;
        RECT 8.156 13.404 8.188 15.912 ;
  LAYER M3 ;
        RECT 8.156 13.424 8.188 13.456 ;
  LAYER M1 ;
        RECT 8.22 13.404 8.252 15.912 ;
  LAYER M3 ;
        RECT 8.22 15.86 8.252 15.892 ;
  LAYER M1 ;
        RECT 8.284 13.404 8.316 15.912 ;
  LAYER M3 ;
        RECT 8.284 13.424 8.316 13.456 ;
  LAYER M1 ;
        RECT 8.348 13.404 8.38 15.912 ;
  LAYER M3 ;
        RECT 8.348 15.86 8.38 15.892 ;
  LAYER M1 ;
        RECT 8.412 13.404 8.444 15.912 ;
  LAYER M3 ;
        RECT 8.412 13.424 8.444 13.456 ;
  LAYER M1 ;
        RECT 8.476 13.404 8.508 15.912 ;
  LAYER M3 ;
        RECT 8.476 15.86 8.508 15.892 ;
  LAYER M1 ;
        RECT 8.54 13.404 8.572 15.912 ;
  LAYER M3 ;
        RECT 8.54 13.424 8.572 13.456 ;
  LAYER M1 ;
        RECT 8.604 13.404 8.636 15.912 ;
  LAYER M3 ;
        RECT 8.604 15.86 8.636 15.892 ;
  LAYER M1 ;
        RECT 8.668 13.404 8.7 15.912 ;
  LAYER M3 ;
        RECT 8.668 13.424 8.7 13.456 ;
  LAYER M1 ;
        RECT 8.732 13.404 8.764 15.912 ;
  LAYER M3 ;
        RECT 8.732 15.86 8.764 15.892 ;
  LAYER M1 ;
        RECT 8.796 13.404 8.828 15.912 ;
  LAYER M3 ;
        RECT 8.796 13.424 8.828 13.456 ;
  LAYER M1 ;
        RECT 8.86 13.404 8.892 15.912 ;
  LAYER M3 ;
        RECT 8.86 15.86 8.892 15.892 ;
  LAYER M1 ;
        RECT 8.924 13.404 8.956 15.912 ;
  LAYER M3 ;
        RECT 8.924 13.424 8.956 13.456 ;
  LAYER M1 ;
        RECT 8.988 13.404 9.02 15.912 ;
  LAYER M3 ;
        RECT 8.988 15.86 9.02 15.892 ;
  LAYER M1 ;
        RECT 9.052 13.404 9.084 15.912 ;
  LAYER M3 ;
        RECT 9.052 13.424 9.084 13.456 ;
  LAYER M1 ;
        RECT 9.116 13.404 9.148 15.912 ;
  LAYER M3 ;
        RECT 9.116 15.86 9.148 15.892 ;
  LAYER M1 ;
        RECT 9.18 13.404 9.212 15.912 ;
  LAYER M3 ;
        RECT 9.18 13.424 9.212 13.456 ;
  LAYER M1 ;
        RECT 9.244 13.404 9.276 15.912 ;
  LAYER M3 ;
        RECT 9.244 15.86 9.276 15.892 ;
  LAYER M1 ;
        RECT 9.308 13.404 9.34 15.912 ;
  LAYER M3 ;
        RECT 9.308 13.424 9.34 13.456 ;
  LAYER M1 ;
        RECT 9.372 13.404 9.404 15.912 ;
  LAYER M3 ;
        RECT 9.372 15.86 9.404 15.892 ;
  LAYER M1 ;
        RECT 9.436 13.404 9.468 15.912 ;
  LAYER M3 ;
        RECT 9.436 13.424 9.468 13.456 ;
  LAYER M1 ;
        RECT 9.5 13.404 9.532 15.912 ;
  LAYER M3 ;
        RECT 9.5 15.86 9.532 15.892 ;
  LAYER M1 ;
        RECT 9.564 13.404 9.596 15.912 ;
  LAYER M3 ;
        RECT 9.564 13.424 9.596 13.456 ;
  LAYER M1 ;
        RECT 9.628 13.404 9.66 15.912 ;
  LAYER M3 ;
        RECT 9.628 15.86 9.66 15.892 ;
  LAYER M1 ;
        RECT 9.692 13.404 9.724 15.912 ;
  LAYER M3 ;
        RECT 7.324 13.488 7.356 13.52 ;
  LAYER M2 ;
        RECT 9.692 13.552 9.724 13.584 ;
  LAYER M2 ;
        RECT 7.324 13.616 7.356 13.648 ;
  LAYER M2 ;
        RECT 9.692 13.68 9.724 13.712 ;
  LAYER M2 ;
        RECT 7.324 13.744 7.356 13.776 ;
  LAYER M2 ;
        RECT 9.692 13.808 9.724 13.84 ;
  LAYER M2 ;
        RECT 7.324 13.872 7.356 13.904 ;
  LAYER M2 ;
        RECT 9.692 13.936 9.724 13.968 ;
  LAYER M2 ;
        RECT 7.324 14 7.356 14.032 ;
  LAYER M2 ;
        RECT 9.692 14.064 9.724 14.096 ;
  LAYER M2 ;
        RECT 7.324 14.128 7.356 14.16 ;
  LAYER M2 ;
        RECT 9.692 14.192 9.724 14.224 ;
  LAYER M2 ;
        RECT 7.324 14.256 7.356 14.288 ;
  LAYER M2 ;
        RECT 9.692 14.32 9.724 14.352 ;
  LAYER M2 ;
        RECT 7.324 14.384 7.356 14.416 ;
  LAYER M2 ;
        RECT 9.692 14.448 9.724 14.48 ;
  LAYER M2 ;
        RECT 7.324 14.512 7.356 14.544 ;
  LAYER M2 ;
        RECT 9.692 14.576 9.724 14.608 ;
  LAYER M2 ;
        RECT 7.324 14.64 7.356 14.672 ;
  LAYER M2 ;
        RECT 9.692 14.704 9.724 14.736 ;
  LAYER M2 ;
        RECT 7.324 14.768 7.356 14.8 ;
  LAYER M2 ;
        RECT 9.692 14.832 9.724 14.864 ;
  LAYER M2 ;
        RECT 7.324 14.896 7.356 14.928 ;
  LAYER M2 ;
        RECT 9.692 14.96 9.724 14.992 ;
  LAYER M2 ;
        RECT 7.324 15.024 7.356 15.056 ;
  LAYER M2 ;
        RECT 9.692 15.088 9.724 15.12 ;
  LAYER M2 ;
        RECT 7.324 15.152 7.356 15.184 ;
  LAYER M2 ;
        RECT 9.692 15.216 9.724 15.248 ;
  LAYER M2 ;
        RECT 7.324 15.28 7.356 15.312 ;
  LAYER M2 ;
        RECT 9.692 15.344 9.724 15.376 ;
  LAYER M2 ;
        RECT 7.324 15.408 7.356 15.44 ;
  LAYER M2 ;
        RECT 9.692 15.472 9.724 15.504 ;
  LAYER M2 ;
        RECT 7.324 15.536 7.356 15.568 ;
  LAYER M2 ;
        RECT 9.692 15.6 9.724 15.632 ;
  LAYER M2 ;
        RECT 7.324 15.664 7.356 15.696 ;
  LAYER M2 ;
        RECT 9.692 15.728 9.724 15.76 ;
  LAYER M2 ;
        RECT 7.276 13.356 9.772 15.96 ;
  LAYER M1 ;
        RECT 7.324 16.512 7.356 19.02 ;
  LAYER M3 ;
        RECT 7.324 18.968 7.356 19 ;
  LAYER M1 ;
        RECT 7.388 16.512 7.42 19.02 ;
  LAYER M3 ;
        RECT 7.388 16.532 7.42 16.564 ;
  LAYER M1 ;
        RECT 7.452 16.512 7.484 19.02 ;
  LAYER M3 ;
        RECT 7.452 18.968 7.484 19 ;
  LAYER M1 ;
        RECT 7.516 16.512 7.548 19.02 ;
  LAYER M3 ;
        RECT 7.516 16.532 7.548 16.564 ;
  LAYER M1 ;
        RECT 7.58 16.512 7.612 19.02 ;
  LAYER M3 ;
        RECT 7.58 18.968 7.612 19 ;
  LAYER M1 ;
        RECT 7.644 16.512 7.676 19.02 ;
  LAYER M3 ;
        RECT 7.644 16.532 7.676 16.564 ;
  LAYER M1 ;
        RECT 7.708 16.512 7.74 19.02 ;
  LAYER M3 ;
        RECT 7.708 18.968 7.74 19 ;
  LAYER M1 ;
        RECT 7.772 16.512 7.804 19.02 ;
  LAYER M3 ;
        RECT 7.772 16.532 7.804 16.564 ;
  LAYER M1 ;
        RECT 7.836 16.512 7.868 19.02 ;
  LAYER M3 ;
        RECT 7.836 18.968 7.868 19 ;
  LAYER M1 ;
        RECT 7.9 16.512 7.932 19.02 ;
  LAYER M3 ;
        RECT 7.9 16.532 7.932 16.564 ;
  LAYER M1 ;
        RECT 7.964 16.512 7.996 19.02 ;
  LAYER M3 ;
        RECT 7.964 18.968 7.996 19 ;
  LAYER M1 ;
        RECT 8.028 16.512 8.06 19.02 ;
  LAYER M3 ;
        RECT 8.028 16.532 8.06 16.564 ;
  LAYER M1 ;
        RECT 8.092 16.512 8.124 19.02 ;
  LAYER M3 ;
        RECT 8.092 18.968 8.124 19 ;
  LAYER M1 ;
        RECT 8.156 16.512 8.188 19.02 ;
  LAYER M3 ;
        RECT 8.156 16.532 8.188 16.564 ;
  LAYER M1 ;
        RECT 8.22 16.512 8.252 19.02 ;
  LAYER M3 ;
        RECT 8.22 18.968 8.252 19 ;
  LAYER M1 ;
        RECT 8.284 16.512 8.316 19.02 ;
  LAYER M3 ;
        RECT 8.284 16.532 8.316 16.564 ;
  LAYER M1 ;
        RECT 8.348 16.512 8.38 19.02 ;
  LAYER M3 ;
        RECT 8.348 18.968 8.38 19 ;
  LAYER M1 ;
        RECT 8.412 16.512 8.444 19.02 ;
  LAYER M3 ;
        RECT 8.412 16.532 8.444 16.564 ;
  LAYER M1 ;
        RECT 8.476 16.512 8.508 19.02 ;
  LAYER M3 ;
        RECT 8.476 18.968 8.508 19 ;
  LAYER M1 ;
        RECT 8.54 16.512 8.572 19.02 ;
  LAYER M3 ;
        RECT 8.54 16.532 8.572 16.564 ;
  LAYER M1 ;
        RECT 8.604 16.512 8.636 19.02 ;
  LAYER M3 ;
        RECT 8.604 18.968 8.636 19 ;
  LAYER M1 ;
        RECT 8.668 16.512 8.7 19.02 ;
  LAYER M3 ;
        RECT 8.668 16.532 8.7 16.564 ;
  LAYER M1 ;
        RECT 8.732 16.512 8.764 19.02 ;
  LAYER M3 ;
        RECT 8.732 18.968 8.764 19 ;
  LAYER M1 ;
        RECT 8.796 16.512 8.828 19.02 ;
  LAYER M3 ;
        RECT 8.796 16.532 8.828 16.564 ;
  LAYER M1 ;
        RECT 8.86 16.512 8.892 19.02 ;
  LAYER M3 ;
        RECT 8.86 18.968 8.892 19 ;
  LAYER M1 ;
        RECT 8.924 16.512 8.956 19.02 ;
  LAYER M3 ;
        RECT 8.924 16.532 8.956 16.564 ;
  LAYER M1 ;
        RECT 8.988 16.512 9.02 19.02 ;
  LAYER M3 ;
        RECT 8.988 18.968 9.02 19 ;
  LAYER M1 ;
        RECT 9.052 16.512 9.084 19.02 ;
  LAYER M3 ;
        RECT 9.052 16.532 9.084 16.564 ;
  LAYER M1 ;
        RECT 9.116 16.512 9.148 19.02 ;
  LAYER M3 ;
        RECT 9.116 18.968 9.148 19 ;
  LAYER M1 ;
        RECT 9.18 16.512 9.212 19.02 ;
  LAYER M3 ;
        RECT 9.18 16.532 9.212 16.564 ;
  LAYER M1 ;
        RECT 9.244 16.512 9.276 19.02 ;
  LAYER M3 ;
        RECT 9.244 18.968 9.276 19 ;
  LAYER M1 ;
        RECT 9.308 16.512 9.34 19.02 ;
  LAYER M3 ;
        RECT 9.308 16.532 9.34 16.564 ;
  LAYER M1 ;
        RECT 9.372 16.512 9.404 19.02 ;
  LAYER M3 ;
        RECT 9.372 18.968 9.404 19 ;
  LAYER M1 ;
        RECT 9.436 16.512 9.468 19.02 ;
  LAYER M3 ;
        RECT 9.436 16.532 9.468 16.564 ;
  LAYER M1 ;
        RECT 9.5 16.512 9.532 19.02 ;
  LAYER M3 ;
        RECT 9.5 18.968 9.532 19 ;
  LAYER M1 ;
        RECT 9.564 16.512 9.596 19.02 ;
  LAYER M3 ;
        RECT 9.564 16.532 9.596 16.564 ;
  LAYER M1 ;
        RECT 9.628 16.512 9.66 19.02 ;
  LAYER M3 ;
        RECT 9.628 18.968 9.66 19 ;
  LAYER M1 ;
        RECT 9.692 16.512 9.724 19.02 ;
  LAYER M3 ;
        RECT 7.324 16.596 7.356 16.628 ;
  LAYER M2 ;
        RECT 9.692 16.66 9.724 16.692 ;
  LAYER M2 ;
        RECT 7.324 16.724 7.356 16.756 ;
  LAYER M2 ;
        RECT 9.692 16.788 9.724 16.82 ;
  LAYER M2 ;
        RECT 7.324 16.852 7.356 16.884 ;
  LAYER M2 ;
        RECT 9.692 16.916 9.724 16.948 ;
  LAYER M2 ;
        RECT 7.324 16.98 7.356 17.012 ;
  LAYER M2 ;
        RECT 9.692 17.044 9.724 17.076 ;
  LAYER M2 ;
        RECT 7.324 17.108 7.356 17.14 ;
  LAYER M2 ;
        RECT 9.692 17.172 9.724 17.204 ;
  LAYER M2 ;
        RECT 7.324 17.236 7.356 17.268 ;
  LAYER M2 ;
        RECT 9.692 17.3 9.724 17.332 ;
  LAYER M2 ;
        RECT 7.324 17.364 7.356 17.396 ;
  LAYER M2 ;
        RECT 9.692 17.428 9.724 17.46 ;
  LAYER M2 ;
        RECT 7.324 17.492 7.356 17.524 ;
  LAYER M2 ;
        RECT 9.692 17.556 9.724 17.588 ;
  LAYER M2 ;
        RECT 7.324 17.62 7.356 17.652 ;
  LAYER M2 ;
        RECT 9.692 17.684 9.724 17.716 ;
  LAYER M2 ;
        RECT 7.324 17.748 7.356 17.78 ;
  LAYER M2 ;
        RECT 9.692 17.812 9.724 17.844 ;
  LAYER M2 ;
        RECT 7.324 17.876 7.356 17.908 ;
  LAYER M2 ;
        RECT 9.692 17.94 9.724 17.972 ;
  LAYER M2 ;
        RECT 7.324 18.004 7.356 18.036 ;
  LAYER M2 ;
        RECT 9.692 18.068 9.724 18.1 ;
  LAYER M2 ;
        RECT 7.324 18.132 7.356 18.164 ;
  LAYER M2 ;
        RECT 9.692 18.196 9.724 18.228 ;
  LAYER M2 ;
        RECT 7.324 18.26 7.356 18.292 ;
  LAYER M2 ;
        RECT 9.692 18.324 9.724 18.356 ;
  LAYER M2 ;
        RECT 7.324 18.388 7.356 18.42 ;
  LAYER M2 ;
        RECT 9.692 18.452 9.724 18.484 ;
  LAYER M2 ;
        RECT 7.324 18.516 7.356 18.548 ;
  LAYER M2 ;
        RECT 9.692 18.58 9.724 18.612 ;
  LAYER M2 ;
        RECT 7.324 18.644 7.356 18.676 ;
  LAYER M2 ;
        RECT 9.692 18.708 9.724 18.74 ;
  LAYER M2 ;
        RECT 7.324 18.772 7.356 18.804 ;
  LAYER M2 ;
        RECT 9.692 18.836 9.724 18.868 ;
  LAYER M2 ;
        RECT 7.276 16.464 9.772 19.068 ;
  LAYER M1 ;
        RECT 10.94 0.972 10.972 3.48 ;
  LAYER M3 ;
        RECT 10.94 3.428 10.972 3.46 ;
  LAYER M1 ;
        RECT 11.004 0.972 11.036 3.48 ;
  LAYER M3 ;
        RECT 11.004 0.992 11.036 1.024 ;
  LAYER M1 ;
        RECT 11.068 0.972 11.1 3.48 ;
  LAYER M3 ;
        RECT 11.068 3.428 11.1 3.46 ;
  LAYER M1 ;
        RECT 11.132 0.972 11.164 3.48 ;
  LAYER M3 ;
        RECT 11.132 0.992 11.164 1.024 ;
  LAYER M1 ;
        RECT 11.196 0.972 11.228 3.48 ;
  LAYER M3 ;
        RECT 11.196 3.428 11.228 3.46 ;
  LAYER M1 ;
        RECT 11.26 0.972 11.292 3.48 ;
  LAYER M3 ;
        RECT 11.26 0.992 11.292 1.024 ;
  LAYER M1 ;
        RECT 11.324 0.972 11.356 3.48 ;
  LAYER M3 ;
        RECT 11.324 3.428 11.356 3.46 ;
  LAYER M1 ;
        RECT 11.388 0.972 11.42 3.48 ;
  LAYER M3 ;
        RECT 11.388 0.992 11.42 1.024 ;
  LAYER M1 ;
        RECT 11.452 0.972 11.484 3.48 ;
  LAYER M3 ;
        RECT 11.452 3.428 11.484 3.46 ;
  LAYER M1 ;
        RECT 11.516 0.972 11.548 3.48 ;
  LAYER M3 ;
        RECT 11.516 0.992 11.548 1.024 ;
  LAYER M1 ;
        RECT 11.58 0.972 11.612 3.48 ;
  LAYER M3 ;
        RECT 11.58 3.428 11.612 3.46 ;
  LAYER M1 ;
        RECT 11.644 0.972 11.676 3.48 ;
  LAYER M3 ;
        RECT 11.644 0.992 11.676 1.024 ;
  LAYER M1 ;
        RECT 11.708 0.972 11.74 3.48 ;
  LAYER M3 ;
        RECT 11.708 3.428 11.74 3.46 ;
  LAYER M1 ;
        RECT 11.772 0.972 11.804 3.48 ;
  LAYER M3 ;
        RECT 11.772 0.992 11.804 1.024 ;
  LAYER M1 ;
        RECT 11.836 0.972 11.868 3.48 ;
  LAYER M3 ;
        RECT 11.836 3.428 11.868 3.46 ;
  LAYER M1 ;
        RECT 11.9 0.972 11.932 3.48 ;
  LAYER M3 ;
        RECT 11.9 0.992 11.932 1.024 ;
  LAYER M1 ;
        RECT 11.964 0.972 11.996 3.48 ;
  LAYER M3 ;
        RECT 11.964 3.428 11.996 3.46 ;
  LAYER M1 ;
        RECT 12.028 0.972 12.06 3.48 ;
  LAYER M3 ;
        RECT 12.028 0.992 12.06 1.024 ;
  LAYER M1 ;
        RECT 12.092 0.972 12.124 3.48 ;
  LAYER M3 ;
        RECT 12.092 3.428 12.124 3.46 ;
  LAYER M1 ;
        RECT 12.156 0.972 12.188 3.48 ;
  LAYER M3 ;
        RECT 12.156 0.992 12.188 1.024 ;
  LAYER M1 ;
        RECT 12.22 0.972 12.252 3.48 ;
  LAYER M3 ;
        RECT 12.22 3.428 12.252 3.46 ;
  LAYER M1 ;
        RECT 12.284 0.972 12.316 3.48 ;
  LAYER M3 ;
        RECT 12.284 0.992 12.316 1.024 ;
  LAYER M1 ;
        RECT 12.348 0.972 12.38 3.48 ;
  LAYER M3 ;
        RECT 12.348 3.428 12.38 3.46 ;
  LAYER M1 ;
        RECT 12.412 0.972 12.444 3.48 ;
  LAYER M3 ;
        RECT 12.412 0.992 12.444 1.024 ;
  LAYER M1 ;
        RECT 12.476 0.972 12.508 3.48 ;
  LAYER M3 ;
        RECT 12.476 3.428 12.508 3.46 ;
  LAYER M1 ;
        RECT 12.54 0.972 12.572 3.48 ;
  LAYER M3 ;
        RECT 12.54 0.992 12.572 1.024 ;
  LAYER M1 ;
        RECT 12.604 0.972 12.636 3.48 ;
  LAYER M3 ;
        RECT 12.604 3.428 12.636 3.46 ;
  LAYER M1 ;
        RECT 12.668 0.972 12.7 3.48 ;
  LAYER M3 ;
        RECT 12.668 0.992 12.7 1.024 ;
  LAYER M1 ;
        RECT 12.732 0.972 12.764 3.48 ;
  LAYER M3 ;
        RECT 12.732 3.428 12.764 3.46 ;
  LAYER M1 ;
        RECT 12.796 0.972 12.828 3.48 ;
  LAYER M3 ;
        RECT 12.796 0.992 12.828 1.024 ;
  LAYER M1 ;
        RECT 12.86 0.972 12.892 3.48 ;
  LAYER M3 ;
        RECT 12.86 3.428 12.892 3.46 ;
  LAYER M1 ;
        RECT 12.924 0.972 12.956 3.48 ;
  LAYER M3 ;
        RECT 12.924 0.992 12.956 1.024 ;
  LAYER M1 ;
        RECT 12.988 0.972 13.02 3.48 ;
  LAYER M3 ;
        RECT 12.988 3.428 13.02 3.46 ;
  LAYER M1 ;
        RECT 13.052 0.972 13.084 3.48 ;
  LAYER M3 ;
        RECT 13.052 0.992 13.084 1.024 ;
  LAYER M1 ;
        RECT 13.116 0.972 13.148 3.48 ;
  LAYER M3 ;
        RECT 13.116 3.428 13.148 3.46 ;
  LAYER M1 ;
        RECT 13.18 0.972 13.212 3.48 ;
  LAYER M3 ;
        RECT 13.18 0.992 13.212 1.024 ;
  LAYER M1 ;
        RECT 13.244 0.972 13.276 3.48 ;
  LAYER M3 ;
        RECT 13.244 3.428 13.276 3.46 ;
  LAYER M1 ;
        RECT 13.308 0.972 13.34 3.48 ;
  LAYER M3 ;
        RECT 10.94 1.056 10.972 1.088 ;
  LAYER M2 ;
        RECT 13.308 1.12 13.34 1.152 ;
  LAYER M2 ;
        RECT 10.94 1.184 10.972 1.216 ;
  LAYER M2 ;
        RECT 13.308 1.248 13.34 1.28 ;
  LAYER M2 ;
        RECT 10.94 1.312 10.972 1.344 ;
  LAYER M2 ;
        RECT 13.308 1.376 13.34 1.408 ;
  LAYER M2 ;
        RECT 10.94 1.44 10.972 1.472 ;
  LAYER M2 ;
        RECT 13.308 1.504 13.34 1.536 ;
  LAYER M2 ;
        RECT 10.94 1.568 10.972 1.6 ;
  LAYER M2 ;
        RECT 13.308 1.632 13.34 1.664 ;
  LAYER M2 ;
        RECT 10.94 1.696 10.972 1.728 ;
  LAYER M2 ;
        RECT 13.308 1.76 13.34 1.792 ;
  LAYER M2 ;
        RECT 10.94 1.824 10.972 1.856 ;
  LAYER M2 ;
        RECT 13.308 1.888 13.34 1.92 ;
  LAYER M2 ;
        RECT 10.94 1.952 10.972 1.984 ;
  LAYER M2 ;
        RECT 13.308 2.016 13.34 2.048 ;
  LAYER M2 ;
        RECT 10.94 2.08 10.972 2.112 ;
  LAYER M2 ;
        RECT 13.308 2.144 13.34 2.176 ;
  LAYER M2 ;
        RECT 10.94 2.208 10.972 2.24 ;
  LAYER M2 ;
        RECT 13.308 2.272 13.34 2.304 ;
  LAYER M2 ;
        RECT 10.94 2.336 10.972 2.368 ;
  LAYER M2 ;
        RECT 13.308 2.4 13.34 2.432 ;
  LAYER M2 ;
        RECT 10.94 2.464 10.972 2.496 ;
  LAYER M2 ;
        RECT 13.308 2.528 13.34 2.56 ;
  LAYER M2 ;
        RECT 10.94 2.592 10.972 2.624 ;
  LAYER M2 ;
        RECT 13.308 2.656 13.34 2.688 ;
  LAYER M2 ;
        RECT 10.94 2.72 10.972 2.752 ;
  LAYER M2 ;
        RECT 13.308 2.784 13.34 2.816 ;
  LAYER M2 ;
        RECT 10.94 2.848 10.972 2.88 ;
  LAYER M2 ;
        RECT 13.308 2.912 13.34 2.944 ;
  LAYER M2 ;
        RECT 10.94 2.976 10.972 3.008 ;
  LAYER M2 ;
        RECT 13.308 3.04 13.34 3.072 ;
  LAYER M2 ;
        RECT 10.94 3.104 10.972 3.136 ;
  LAYER M2 ;
        RECT 13.308 3.168 13.34 3.2 ;
  LAYER M2 ;
        RECT 10.94 3.232 10.972 3.264 ;
  LAYER M2 ;
        RECT 13.308 3.296 13.34 3.328 ;
  LAYER M2 ;
        RECT 10.892 0.924 13.388 3.528 ;
  LAYER M1 ;
        RECT 10.94 4.08 10.972 6.588 ;
  LAYER M3 ;
        RECT 10.94 6.536 10.972 6.568 ;
  LAYER M1 ;
        RECT 11.004 4.08 11.036 6.588 ;
  LAYER M3 ;
        RECT 11.004 4.1 11.036 4.132 ;
  LAYER M1 ;
        RECT 11.068 4.08 11.1 6.588 ;
  LAYER M3 ;
        RECT 11.068 6.536 11.1 6.568 ;
  LAYER M1 ;
        RECT 11.132 4.08 11.164 6.588 ;
  LAYER M3 ;
        RECT 11.132 4.1 11.164 4.132 ;
  LAYER M1 ;
        RECT 11.196 4.08 11.228 6.588 ;
  LAYER M3 ;
        RECT 11.196 6.536 11.228 6.568 ;
  LAYER M1 ;
        RECT 11.26 4.08 11.292 6.588 ;
  LAYER M3 ;
        RECT 11.26 4.1 11.292 4.132 ;
  LAYER M1 ;
        RECT 11.324 4.08 11.356 6.588 ;
  LAYER M3 ;
        RECT 11.324 6.536 11.356 6.568 ;
  LAYER M1 ;
        RECT 11.388 4.08 11.42 6.588 ;
  LAYER M3 ;
        RECT 11.388 4.1 11.42 4.132 ;
  LAYER M1 ;
        RECT 11.452 4.08 11.484 6.588 ;
  LAYER M3 ;
        RECT 11.452 6.536 11.484 6.568 ;
  LAYER M1 ;
        RECT 11.516 4.08 11.548 6.588 ;
  LAYER M3 ;
        RECT 11.516 4.1 11.548 4.132 ;
  LAYER M1 ;
        RECT 11.58 4.08 11.612 6.588 ;
  LAYER M3 ;
        RECT 11.58 6.536 11.612 6.568 ;
  LAYER M1 ;
        RECT 11.644 4.08 11.676 6.588 ;
  LAYER M3 ;
        RECT 11.644 4.1 11.676 4.132 ;
  LAYER M1 ;
        RECT 11.708 4.08 11.74 6.588 ;
  LAYER M3 ;
        RECT 11.708 6.536 11.74 6.568 ;
  LAYER M1 ;
        RECT 11.772 4.08 11.804 6.588 ;
  LAYER M3 ;
        RECT 11.772 4.1 11.804 4.132 ;
  LAYER M1 ;
        RECT 11.836 4.08 11.868 6.588 ;
  LAYER M3 ;
        RECT 11.836 6.536 11.868 6.568 ;
  LAYER M1 ;
        RECT 11.9 4.08 11.932 6.588 ;
  LAYER M3 ;
        RECT 11.9 4.1 11.932 4.132 ;
  LAYER M1 ;
        RECT 11.964 4.08 11.996 6.588 ;
  LAYER M3 ;
        RECT 11.964 6.536 11.996 6.568 ;
  LAYER M1 ;
        RECT 12.028 4.08 12.06 6.588 ;
  LAYER M3 ;
        RECT 12.028 4.1 12.06 4.132 ;
  LAYER M1 ;
        RECT 12.092 4.08 12.124 6.588 ;
  LAYER M3 ;
        RECT 12.092 6.536 12.124 6.568 ;
  LAYER M1 ;
        RECT 12.156 4.08 12.188 6.588 ;
  LAYER M3 ;
        RECT 12.156 4.1 12.188 4.132 ;
  LAYER M1 ;
        RECT 12.22 4.08 12.252 6.588 ;
  LAYER M3 ;
        RECT 12.22 6.536 12.252 6.568 ;
  LAYER M1 ;
        RECT 12.284 4.08 12.316 6.588 ;
  LAYER M3 ;
        RECT 12.284 4.1 12.316 4.132 ;
  LAYER M1 ;
        RECT 12.348 4.08 12.38 6.588 ;
  LAYER M3 ;
        RECT 12.348 6.536 12.38 6.568 ;
  LAYER M1 ;
        RECT 12.412 4.08 12.444 6.588 ;
  LAYER M3 ;
        RECT 12.412 4.1 12.444 4.132 ;
  LAYER M1 ;
        RECT 12.476 4.08 12.508 6.588 ;
  LAYER M3 ;
        RECT 12.476 6.536 12.508 6.568 ;
  LAYER M1 ;
        RECT 12.54 4.08 12.572 6.588 ;
  LAYER M3 ;
        RECT 12.54 4.1 12.572 4.132 ;
  LAYER M1 ;
        RECT 12.604 4.08 12.636 6.588 ;
  LAYER M3 ;
        RECT 12.604 6.536 12.636 6.568 ;
  LAYER M1 ;
        RECT 12.668 4.08 12.7 6.588 ;
  LAYER M3 ;
        RECT 12.668 4.1 12.7 4.132 ;
  LAYER M1 ;
        RECT 12.732 4.08 12.764 6.588 ;
  LAYER M3 ;
        RECT 12.732 6.536 12.764 6.568 ;
  LAYER M1 ;
        RECT 12.796 4.08 12.828 6.588 ;
  LAYER M3 ;
        RECT 12.796 4.1 12.828 4.132 ;
  LAYER M1 ;
        RECT 12.86 4.08 12.892 6.588 ;
  LAYER M3 ;
        RECT 12.86 6.536 12.892 6.568 ;
  LAYER M1 ;
        RECT 12.924 4.08 12.956 6.588 ;
  LAYER M3 ;
        RECT 12.924 4.1 12.956 4.132 ;
  LAYER M1 ;
        RECT 12.988 4.08 13.02 6.588 ;
  LAYER M3 ;
        RECT 12.988 6.536 13.02 6.568 ;
  LAYER M1 ;
        RECT 13.052 4.08 13.084 6.588 ;
  LAYER M3 ;
        RECT 13.052 4.1 13.084 4.132 ;
  LAYER M1 ;
        RECT 13.116 4.08 13.148 6.588 ;
  LAYER M3 ;
        RECT 13.116 6.536 13.148 6.568 ;
  LAYER M1 ;
        RECT 13.18 4.08 13.212 6.588 ;
  LAYER M3 ;
        RECT 13.18 4.1 13.212 4.132 ;
  LAYER M1 ;
        RECT 13.244 4.08 13.276 6.588 ;
  LAYER M3 ;
        RECT 13.244 6.536 13.276 6.568 ;
  LAYER M1 ;
        RECT 13.308 4.08 13.34 6.588 ;
  LAYER M3 ;
        RECT 10.94 4.164 10.972 4.196 ;
  LAYER M2 ;
        RECT 13.308 4.228 13.34 4.26 ;
  LAYER M2 ;
        RECT 10.94 4.292 10.972 4.324 ;
  LAYER M2 ;
        RECT 13.308 4.356 13.34 4.388 ;
  LAYER M2 ;
        RECT 10.94 4.42 10.972 4.452 ;
  LAYER M2 ;
        RECT 13.308 4.484 13.34 4.516 ;
  LAYER M2 ;
        RECT 10.94 4.548 10.972 4.58 ;
  LAYER M2 ;
        RECT 13.308 4.612 13.34 4.644 ;
  LAYER M2 ;
        RECT 10.94 4.676 10.972 4.708 ;
  LAYER M2 ;
        RECT 13.308 4.74 13.34 4.772 ;
  LAYER M2 ;
        RECT 10.94 4.804 10.972 4.836 ;
  LAYER M2 ;
        RECT 13.308 4.868 13.34 4.9 ;
  LAYER M2 ;
        RECT 10.94 4.932 10.972 4.964 ;
  LAYER M2 ;
        RECT 13.308 4.996 13.34 5.028 ;
  LAYER M2 ;
        RECT 10.94 5.06 10.972 5.092 ;
  LAYER M2 ;
        RECT 13.308 5.124 13.34 5.156 ;
  LAYER M2 ;
        RECT 10.94 5.188 10.972 5.22 ;
  LAYER M2 ;
        RECT 13.308 5.252 13.34 5.284 ;
  LAYER M2 ;
        RECT 10.94 5.316 10.972 5.348 ;
  LAYER M2 ;
        RECT 13.308 5.38 13.34 5.412 ;
  LAYER M2 ;
        RECT 10.94 5.444 10.972 5.476 ;
  LAYER M2 ;
        RECT 13.308 5.508 13.34 5.54 ;
  LAYER M2 ;
        RECT 10.94 5.572 10.972 5.604 ;
  LAYER M2 ;
        RECT 13.308 5.636 13.34 5.668 ;
  LAYER M2 ;
        RECT 10.94 5.7 10.972 5.732 ;
  LAYER M2 ;
        RECT 13.308 5.764 13.34 5.796 ;
  LAYER M2 ;
        RECT 10.94 5.828 10.972 5.86 ;
  LAYER M2 ;
        RECT 13.308 5.892 13.34 5.924 ;
  LAYER M2 ;
        RECT 10.94 5.956 10.972 5.988 ;
  LAYER M2 ;
        RECT 13.308 6.02 13.34 6.052 ;
  LAYER M2 ;
        RECT 10.94 6.084 10.972 6.116 ;
  LAYER M2 ;
        RECT 13.308 6.148 13.34 6.18 ;
  LAYER M2 ;
        RECT 10.94 6.212 10.972 6.244 ;
  LAYER M2 ;
        RECT 13.308 6.276 13.34 6.308 ;
  LAYER M2 ;
        RECT 10.94 6.34 10.972 6.372 ;
  LAYER M2 ;
        RECT 13.308 6.404 13.34 6.436 ;
  LAYER M2 ;
        RECT 10.892 4.032 13.388 6.636 ;
  LAYER M1 ;
        RECT 10.94 7.188 10.972 9.696 ;
  LAYER M3 ;
        RECT 10.94 9.644 10.972 9.676 ;
  LAYER M1 ;
        RECT 11.004 7.188 11.036 9.696 ;
  LAYER M3 ;
        RECT 11.004 7.208 11.036 7.24 ;
  LAYER M1 ;
        RECT 11.068 7.188 11.1 9.696 ;
  LAYER M3 ;
        RECT 11.068 9.644 11.1 9.676 ;
  LAYER M1 ;
        RECT 11.132 7.188 11.164 9.696 ;
  LAYER M3 ;
        RECT 11.132 7.208 11.164 7.24 ;
  LAYER M1 ;
        RECT 11.196 7.188 11.228 9.696 ;
  LAYER M3 ;
        RECT 11.196 9.644 11.228 9.676 ;
  LAYER M1 ;
        RECT 11.26 7.188 11.292 9.696 ;
  LAYER M3 ;
        RECT 11.26 7.208 11.292 7.24 ;
  LAYER M1 ;
        RECT 11.324 7.188 11.356 9.696 ;
  LAYER M3 ;
        RECT 11.324 9.644 11.356 9.676 ;
  LAYER M1 ;
        RECT 11.388 7.188 11.42 9.696 ;
  LAYER M3 ;
        RECT 11.388 7.208 11.42 7.24 ;
  LAYER M1 ;
        RECT 11.452 7.188 11.484 9.696 ;
  LAYER M3 ;
        RECT 11.452 9.644 11.484 9.676 ;
  LAYER M1 ;
        RECT 11.516 7.188 11.548 9.696 ;
  LAYER M3 ;
        RECT 11.516 7.208 11.548 7.24 ;
  LAYER M1 ;
        RECT 11.58 7.188 11.612 9.696 ;
  LAYER M3 ;
        RECT 11.58 9.644 11.612 9.676 ;
  LAYER M1 ;
        RECT 11.644 7.188 11.676 9.696 ;
  LAYER M3 ;
        RECT 11.644 7.208 11.676 7.24 ;
  LAYER M1 ;
        RECT 11.708 7.188 11.74 9.696 ;
  LAYER M3 ;
        RECT 11.708 9.644 11.74 9.676 ;
  LAYER M1 ;
        RECT 11.772 7.188 11.804 9.696 ;
  LAYER M3 ;
        RECT 11.772 7.208 11.804 7.24 ;
  LAYER M1 ;
        RECT 11.836 7.188 11.868 9.696 ;
  LAYER M3 ;
        RECT 11.836 9.644 11.868 9.676 ;
  LAYER M1 ;
        RECT 11.9 7.188 11.932 9.696 ;
  LAYER M3 ;
        RECT 11.9 7.208 11.932 7.24 ;
  LAYER M1 ;
        RECT 11.964 7.188 11.996 9.696 ;
  LAYER M3 ;
        RECT 11.964 9.644 11.996 9.676 ;
  LAYER M1 ;
        RECT 12.028 7.188 12.06 9.696 ;
  LAYER M3 ;
        RECT 12.028 7.208 12.06 7.24 ;
  LAYER M1 ;
        RECT 12.092 7.188 12.124 9.696 ;
  LAYER M3 ;
        RECT 12.092 9.644 12.124 9.676 ;
  LAYER M1 ;
        RECT 12.156 7.188 12.188 9.696 ;
  LAYER M3 ;
        RECT 12.156 7.208 12.188 7.24 ;
  LAYER M1 ;
        RECT 12.22 7.188 12.252 9.696 ;
  LAYER M3 ;
        RECT 12.22 9.644 12.252 9.676 ;
  LAYER M1 ;
        RECT 12.284 7.188 12.316 9.696 ;
  LAYER M3 ;
        RECT 12.284 7.208 12.316 7.24 ;
  LAYER M1 ;
        RECT 12.348 7.188 12.38 9.696 ;
  LAYER M3 ;
        RECT 12.348 9.644 12.38 9.676 ;
  LAYER M1 ;
        RECT 12.412 7.188 12.444 9.696 ;
  LAYER M3 ;
        RECT 12.412 7.208 12.444 7.24 ;
  LAYER M1 ;
        RECT 12.476 7.188 12.508 9.696 ;
  LAYER M3 ;
        RECT 12.476 9.644 12.508 9.676 ;
  LAYER M1 ;
        RECT 12.54 7.188 12.572 9.696 ;
  LAYER M3 ;
        RECT 12.54 7.208 12.572 7.24 ;
  LAYER M1 ;
        RECT 12.604 7.188 12.636 9.696 ;
  LAYER M3 ;
        RECT 12.604 9.644 12.636 9.676 ;
  LAYER M1 ;
        RECT 12.668 7.188 12.7 9.696 ;
  LAYER M3 ;
        RECT 12.668 7.208 12.7 7.24 ;
  LAYER M1 ;
        RECT 12.732 7.188 12.764 9.696 ;
  LAYER M3 ;
        RECT 12.732 9.644 12.764 9.676 ;
  LAYER M1 ;
        RECT 12.796 7.188 12.828 9.696 ;
  LAYER M3 ;
        RECT 12.796 7.208 12.828 7.24 ;
  LAYER M1 ;
        RECT 12.86 7.188 12.892 9.696 ;
  LAYER M3 ;
        RECT 12.86 9.644 12.892 9.676 ;
  LAYER M1 ;
        RECT 12.924 7.188 12.956 9.696 ;
  LAYER M3 ;
        RECT 12.924 7.208 12.956 7.24 ;
  LAYER M1 ;
        RECT 12.988 7.188 13.02 9.696 ;
  LAYER M3 ;
        RECT 12.988 9.644 13.02 9.676 ;
  LAYER M1 ;
        RECT 13.052 7.188 13.084 9.696 ;
  LAYER M3 ;
        RECT 13.052 7.208 13.084 7.24 ;
  LAYER M1 ;
        RECT 13.116 7.188 13.148 9.696 ;
  LAYER M3 ;
        RECT 13.116 9.644 13.148 9.676 ;
  LAYER M1 ;
        RECT 13.18 7.188 13.212 9.696 ;
  LAYER M3 ;
        RECT 13.18 7.208 13.212 7.24 ;
  LAYER M1 ;
        RECT 13.244 7.188 13.276 9.696 ;
  LAYER M3 ;
        RECT 13.244 9.644 13.276 9.676 ;
  LAYER M1 ;
        RECT 13.308 7.188 13.34 9.696 ;
  LAYER M3 ;
        RECT 10.94 7.272 10.972 7.304 ;
  LAYER M2 ;
        RECT 13.308 7.336 13.34 7.368 ;
  LAYER M2 ;
        RECT 10.94 7.4 10.972 7.432 ;
  LAYER M2 ;
        RECT 13.308 7.464 13.34 7.496 ;
  LAYER M2 ;
        RECT 10.94 7.528 10.972 7.56 ;
  LAYER M2 ;
        RECT 13.308 7.592 13.34 7.624 ;
  LAYER M2 ;
        RECT 10.94 7.656 10.972 7.688 ;
  LAYER M2 ;
        RECT 13.308 7.72 13.34 7.752 ;
  LAYER M2 ;
        RECT 10.94 7.784 10.972 7.816 ;
  LAYER M2 ;
        RECT 13.308 7.848 13.34 7.88 ;
  LAYER M2 ;
        RECT 10.94 7.912 10.972 7.944 ;
  LAYER M2 ;
        RECT 13.308 7.976 13.34 8.008 ;
  LAYER M2 ;
        RECT 10.94 8.04 10.972 8.072 ;
  LAYER M2 ;
        RECT 13.308 8.104 13.34 8.136 ;
  LAYER M2 ;
        RECT 10.94 8.168 10.972 8.2 ;
  LAYER M2 ;
        RECT 13.308 8.232 13.34 8.264 ;
  LAYER M2 ;
        RECT 10.94 8.296 10.972 8.328 ;
  LAYER M2 ;
        RECT 13.308 8.36 13.34 8.392 ;
  LAYER M2 ;
        RECT 10.94 8.424 10.972 8.456 ;
  LAYER M2 ;
        RECT 13.308 8.488 13.34 8.52 ;
  LAYER M2 ;
        RECT 10.94 8.552 10.972 8.584 ;
  LAYER M2 ;
        RECT 13.308 8.616 13.34 8.648 ;
  LAYER M2 ;
        RECT 10.94 8.68 10.972 8.712 ;
  LAYER M2 ;
        RECT 13.308 8.744 13.34 8.776 ;
  LAYER M2 ;
        RECT 10.94 8.808 10.972 8.84 ;
  LAYER M2 ;
        RECT 13.308 8.872 13.34 8.904 ;
  LAYER M2 ;
        RECT 10.94 8.936 10.972 8.968 ;
  LAYER M2 ;
        RECT 13.308 9 13.34 9.032 ;
  LAYER M2 ;
        RECT 10.94 9.064 10.972 9.096 ;
  LAYER M2 ;
        RECT 13.308 9.128 13.34 9.16 ;
  LAYER M2 ;
        RECT 10.94 9.192 10.972 9.224 ;
  LAYER M2 ;
        RECT 13.308 9.256 13.34 9.288 ;
  LAYER M2 ;
        RECT 10.94 9.32 10.972 9.352 ;
  LAYER M2 ;
        RECT 13.308 9.384 13.34 9.416 ;
  LAYER M2 ;
        RECT 10.94 9.448 10.972 9.48 ;
  LAYER M2 ;
        RECT 13.308 9.512 13.34 9.544 ;
  LAYER M2 ;
        RECT 10.892 7.14 13.388 9.744 ;
  LAYER M1 ;
        RECT 10.94 10.296 10.972 12.804 ;
  LAYER M3 ;
        RECT 10.94 12.752 10.972 12.784 ;
  LAYER M1 ;
        RECT 11.004 10.296 11.036 12.804 ;
  LAYER M3 ;
        RECT 11.004 10.316 11.036 10.348 ;
  LAYER M1 ;
        RECT 11.068 10.296 11.1 12.804 ;
  LAYER M3 ;
        RECT 11.068 12.752 11.1 12.784 ;
  LAYER M1 ;
        RECT 11.132 10.296 11.164 12.804 ;
  LAYER M3 ;
        RECT 11.132 10.316 11.164 10.348 ;
  LAYER M1 ;
        RECT 11.196 10.296 11.228 12.804 ;
  LAYER M3 ;
        RECT 11.196 12.752 11.228 12.784 ;
  LAYER M1 ;
        RECT 11.26 10.296 11.292 12.804 ;
  LAYER M3 ;
        RECT 11.26 10.316 11.292 10.348 ;
  LAYER M1 ;
        RECT 11.324 10.296 11.356 12.804 ;
  LAYER M3 ;
        RECT 11.324 12.752 11.356 12.784 ;
  LAYER M1 ;
        RECT 11.388 10.296 11.42 12.804 ;
  LAYER M3 ;
        RECT 11.388 10.316 11.42 10.348 ;
  LAYER M1 ;
        RECT 11.452 10.296 11.484 12.804 ;
  LAYER M3 ;
        RECT 11.452 12.752 11.484 12.784 ;
  LAYER M1 ;
        RECT 11.516 10.296 11.548 12.804 ;
  LAYER M3 ;
        RECT 11.516 10.316 11.548 10.348 ;
  LAYER M1 ;
        RECT 11.58 10.296 11.612 12.804 ;
  LAYER M3 ;
        RECT 11.58 12.752 11.612 12.784 ;
  LAYER M1 ;
        RECT 11.644 10.296 11.676 12.804 ;
  LAYER M3 ;
        RECT 11.644 10.316 11.676 10.348 ;
  LAYER M1 ;
        RECT 11.708 10.296 11.74 12.804 ;
  LAYER M3 ;
        RECT 11.708 12.752 11.74 12.784 ;
  LAYER M1 ;
        RECT 11.772 10.296 11.804 12.804 ;
  LAYER M3 ;
        RECT 11.772 10.316 11.804 10.348 ;
  LAYER M1 ;
        RECT 11.836 10.296 11.868 12.804 ;
  LAYER M3 ;
        RECT 11.836 12.752 11.868 12.784 ;
  LAYER M1 ;
        RECT 11.9 10.296 11.932 12.804 ;
  LAYER M3 ;
        RECT 11.9 10.316 11.932 10.348 ;
  LAYER M1 ;
        RECT 11.964 10.296 11.996 12.804 ;
  LAYER M3 ;
        RECT 11.964 12.752 11.996 12.784 ;
  LAYER M1 ;
        RECT 12.028 10.296 12.06 12.804 ;
  LAYER M3 ;
        RECT 12.028 10.316 12.06 10.348 ;
  LAYER M1 ;
        RECT 12.092 10.296 12.124 12.804 ;
  LAYER M3 ;
        RECT 12.092 12.752 12.124 12.784 ;
  LAYER M1 ;
        RECT 12.156 10.296 12.188 12.804 ;
  LAYER M3 ;
        RECT 12.156 10.316 12.188 10.348 ;
  LAYER M1 ;
        RECT 12.22 10.296 12.252 12.804 ;
  LAYER M3 ;
        RECT 12.22 12.752 12.252 12.784 ;
  LAYER M1 ;
        RECT 12.284 10.296 12.316 12.804 ;
  LAYER M3 ;
        RECT 12.284 10.316 12.316 10.348 ;
  LAYER M1 ;
        RECT 12.348 10.296 12.38 12.804 ;
  LAYER M3 ;
        RECT 12.348 12.752 12.38 12.784 ;
  LAYER M1 ;
        RECT 12.412 10.296 12.444 12.804 ;
  LAYER M3 ;
        RECT 12.412 10.316 12.444 10.348 ;
  LAYER M1 ;
        RECT 12.476 10.296 12.508 12.804 ;
  LAYER M3 ;
        RECT 12.476 12.752 12.508 12.784 ;
  LAYER M1 ;
        RECT 12.54 10.296 12.572 12.804 ;
  LAYER M3 ;
        RECT 12.54 10.316 12.572 10.348 ;
  LAYER M1 ;
        RECT 12.604 10.296 12.636 12.804 ;
  LAYER M3 ;
        RECT 12.604 12.752 12.636 12.784 ;
  LAYER M1 ;
        RECT 12.668 10.296 12.7 12.804 ;
  LAYER M3 ;
        RECT 12.668 10.316 12.7 10.348 ;
  LAYER M1 ;
        RECT 12.732 10.296 12.764 12.804 ;
  LAYER M3 ;
        RECT 12.732 12.752 12.764 12.784 ;
  LAYER M1 ;
        RECT 12.796 10.296 12.828 12.804 ;
  LAYER M3 ;
        RECT 12.796 10.316 12.828 10.348 ;
  LAYER M1 ;
        RECT 12.86 10.296 12.892 12.804 ;
  LAYER M3 ;
        RECT 12.86 12.752 12.892 12.784 ;
  LAYER M1 ;
        RECT 12.924 10.296 12.956 12.804 ;
  LAYER M3 ;
        RECT 12.924 10.316 12.956 10.348 ;
  LAYER M1 ;
        RECT 12.988 10.296 13.02 12.804 ;
  LAYER M3 ;
        RECT 12.988 12.752 13.02 12.784 ;
  LAYER M1 ;
        RECT 13.052 10.296 13.084 12.804 ;
  LAYER M3 ;
        RECT 13.052 10.316 13.084 10.348 ;
  LAYER M1 ;
        RECT 13.116 10.296 13.148 12.804 ;
  LAYER M3 ;
        RECT 13.116 12.752 13.148 12.784 ;
  LAYER M1 ;
        RECT 13.18 10.296 13.212 12.804 ;
  LAYER M3 ;
        RECT 13.18 10.316 13.212 10.348 ;
  LAYER M1 ;
        RECT 13.244 10.296 13.276 12.804 ;
  LAYER M3 ;
        RECT 13.244 12.752 13.276 12.784 ;
  LAYER M1 ;
        RECT 13.308 10.296 13.34 12.804 ;
  LAYER M3 ;
        RECT 10.94 10.38 10.972 10.412 ;
  LAYER M2 ;
        RECT 13.308 10.444 13.34 10.476 ;
  LAYER M2 ;
        RECT 10.94 10.508 10.972 10.54 ;
  LAYER M2 ;
        RECT 13.308 10.572 13.34 10.604 ;
  LAYER M2 ;
        RECT 10.94 10.636 10.972 10.668 ;
  LAYER M2 ;
        RECT 13.308 10.7 13.34 10.732 ;
  LAYER M2 ;
        RECT 10.94 10.764 10.972 10.796 ;
  LAYER M2 ;
        RECT 13.308 10.828 13.34 10.86 ;
  LAYER M2 ;
        RECT 10.94 10.892 10.972 10.924 ;
  LAYER M2 ;
        RECT 13.308 10.956 13.34 10.988 ;
  LAYER M2 ;
        RECT 10.94 11.02 10.972 11.052 ;
  LAYER M2 ;
        RECT 13.308 11.084 13.34 11.116 ;
  LAYER M2 ;
        RECT 10.94 11.148 10.972 11.18 ;
  LAYER M2 ;
        RECT 13.308 11.212 13.34 11.244 ;
  LAYER M2 ;
        RECT 10.94 11.276 10.972 11.308 ;
  LAYER M2 ;
        RECT 13.308 11.34 13.34 11.372 ;
  LAYER M2 ;
        RECT 10.94 11.404 10.972 11.436 ;
  LAYER M2 ;
        RECT 13.308 11.468 13.34 11.5 ;
  LAYER M2 ;
        RECT 10.94 11.532 10.972 11.564 ;
  LAYER M2 ;
        RECT 13.308 11.596 13.34 11.628 ;
  LAYER M2 ;
        RECT 10.94 11.66 10.972 11.692 ;
  LAYER M2 ;
        RECT 13.308 11.724 13.34 11.756 ;
  LAYER M2 ;
        RECT 10.94 11.788 10.972 11.82 ;
  LAYER M2 ;
        RECT 13.308 11.852 13.34 11.884 ;
  LAYER M2 ;
        RECT 10.94 11.916 10.972 11.948 ;
  LAYER M2 ;
        RECT 13.308 11.98 13.34 12.012 ;
  LAYER M2 ;
        RECT 10.94 12.044 10.972 12.076 ;
  LAYER M2 ;
        RECT 13.308 12.108 13.34 12.14 ;
  LAYER M2 ;
        RECT 10.94 12.172 10.972 12.204 ;
  LAYER M2 ;
        RECT 13.308 12.236 13.34 12.268 ;
  LAYER M2 ;
        RECT 10.94 12.3 10.972 12.332 ;
  LAYER M2 ;
        RECT 13.308 12.364 13.34 12.396 ;
  LAYER M2 ;
        RECT 10.94 12.428 10.972 12.46 ;
  LAYER M2 ;
        RECT 13.308 12.492 13.34 12.524 ;
  LAYER M2 ;
        RECT 10.94 12.556 10.972 12.588 ;
  LAYER M2 ;
        RECT 13.308 12.62 13.34 12.652 ;
  LAYER M2 ;
        RECT 10.892 10.248 13.388 12.852 ;
  LAYER M1 ;
        RECT 10.94 13.404 10.972 15.912 ;
  LAYER M3 ;
        RECT 10.94 15.86 10.972 15.892 ;
  LAYER M1 ;
        RECT 11.004 13.404 11.036 15.912 ;
  LAYER M3 ;
        RECT 11.004 13.424 11.036 13.456 ;
  LAYER M1 ;
        RECT 11.068 13.404 11.1 15.912 ;
  LAYER M3 ;
        RECT 11.068 15.86 11.1 15.892 ;
  LAYER M1 ;
        RECT 11.132 13.404 11.164 15.912 ;
  LAYER M3 ;
        RECT 11.132 13.424 11.164 13.456 ;
  LAYER M1 ;
        RECT 11.196 13.404 11.228 15.912 ;
  LAYER M3 ;
        RECT 11.196 15.86 11.228 15.892 ;
  LAYER M1 ;
        RECT 11.26 13.404 11.292 15.912 ;
  LAYER M3 ;
        RECT 11.26 13.424 11.292 13.456 ;
  LAYER M1 ;
        RECT 11.324 13.404 11.356 15.912 ;
  LAYER M3 ;
        RECT 11.324 15.86 11.356 15.892 ;
  LAYER M1 ;
        RECT 11.388 13.404 11.42 15.912 ;
  LAYER M3 ;
        RECT 11.388 13.424 11.42 13.456 ;
  LAYER M1 ;
        RECT 11.452 13.404 11.484 15.912 ;
  LAYER M3 ;
        RECT 11.452 15.86 11.484 15.892 ;
  LAYER M1 ;
        RECT 11.516 13.404 11.548 15.912 ;
  LAYER M3 ;
        RECT 11.516 13.424 11.548 13.456 ;
  LAYER M1 ;
        RECT 11.58 13.404 11.612 15.912 ;
  LAYER M3 ;
        RECT 11.58 15.86 11.612 15.892 ;
  LAYER M1 ;
        RECT 11.644 13.404 11.676 15.912 ;
  LAYER M3 ;
        RECT 11.644 13.424 11.676 13.456 ;
  LAYER M1 ;
        RECT 11.708 13.404 11.74 15.912 ;
  LAYER M3 ;
        RECT 11.708 15.86 11.74 15.892 ;
  LAYER M1 ;
        RECT 11.772 13.404 11.804 15.912 ;
  LAYER M3 ;
        RECT 11.772 13.424 11.804 13.456 ;
  LAYER M1 ;
        RECT 11.836 13.404 11.868 15.912 ;
  LAYER M3 ;
        RECT 11.836 15.86 11.868 15.892 ;
  LAYER M1 ;
        RECT 11.9 13.404 11.932 15.912 ;
  LAYER M3 ;
        RECT 11.9 13.424 11.932 13.456 ;
  LAYER M1 ;
        RECT 11.964 13.404 11.996 15.912 ;
  LAYER M3 ;
        RECT 11.964 15.86 11.996 15.892 ;
  LAYER M1 ;
        RECT 12.028 13.404 12.06 15.912 ;
  LAYER M3 ;
        RECT 12.028 13.424 12.06 13.456 ;
  LAYER M1 ;
        RECT 12.092 13.404 12.124 15.912 ;
  LAYER M3 ;
        RECT 12.092 15.86 12.124 15.892 ;
  LAYER M1 ;
        RECT 12.156 13.404 12.188 15.912 ;
  LAYER M3 ;
        RECT 12.156 13.424 12.188 13.456 ;
  LAYER M1 ;
        RECT 12.22 13.404 12.252 15.912 ;
  LAYER M3 ;
        RECT 12.22 15.86 12.252 15.892 ;
  LAYER M1 ;
        RECT 12.284 13.404 12.316 15.912 ;
  LAYER M3 ;
        RECT 12.284 13.424 12.316 13.456 ;
  LAYER M1 ;
        RECT 12.348 13.404 12.38 15.912 ;
  LAYER M3 ;
        RECT 12.348 15.86 12.38 15.892 ;
  LAYER M1 ;
        RECT 12.412 13.404 12.444 15.912 ;
  LAYER M3 ;
        RECT 12.412 13.424 12.444 13.456 ;
  LAYER M1 ;
        RECT 12.476 13.404 12.508 15.912 ;
  LAYER M3 ;
        RECT 12.476 15.86 12.508 15.892 ;
  LAYER M1 ;
        RECT 12.54 13.404 12.572 15.912 ;
  LAYER M3 ;
        RECT 12.54 13.424 12.572 13.456 ;
  LAYER M1 ;
        RECT 12.604 13.404 12.636 15.912 ;
  LAYER M3 ;
        RECT 12.604 15.86 12.636 15.892 ;
  LAYER M1 ;
        RECT 12.668 13.404 12.7 15.912 ;
  LAYER M3 ;
        RECT 12.668 13.424 12.7 13.456 ;
  LAYER M1 ;
        RECT 12.732 13.404 12.764 15.912 ;
  LAYER M3 ;
        RECT 12.732 15.86 12.764 15.892 ;
  LAYER M1 ;
        RECT 12.796 13.404 12.828 15.912 ;
  LAYER M3 ;
        RECT 12.796 13.424 12.828 13.456 ;
  LAYER M1 ;
        RECT 12.86 13.404 12.892 15.912 ;
  LAYER M3 ;
        RECT 12.86 15.86 12.892 15.892 ;
  LAYER M1 ;
        RECT 12.924 13.404 12.956 15.912 ;
  LAYER M3 ;
        RECT 12.924 13.424 12.956 13.456 ;
  LAYER M1 ;
        RECT 12.988 13.404 13.02 15.912 ;
  LAYER M3 ;
        RECT 12.988 15.86 13.02 15.892 ;
  LAYER M1 ;
        RECT 13.052 13.404 13.084 15.912 ;
  LAYER M3 ;
        RECT 13.052 13.424 13.084 13.456 ;
  LAYER M1 ;
        RECT 13.116 13.404 13.148 15.912 ;
  LAYER M3 ;
        RECT 13.116 15.86 13.148 15.892 ;
  LAYER M1 ;
        RECT 13.18 13.404 13.212 15.912 ;
  LAYER M3 ;
        RECT 13.18 13.424 13.212 13.456 ;
  LAYER M1 ;
        RECT 13.244 13.404 13.276 15.912 ;
  LAYER M3 ;
        RECT 13.244 15.86 13.276 15.892 ;
  LAYER M1 ;
        RECT 13.308 13.404 13.34 15.912 ;
  LAYER M3 ;
        RECT 10.94 13.488 10.972 13.52 ;
  LAYER M2 ;
        RECT 13.308 13.552 13.34 13.584 ;
  LAYER M2 ;
        RECT 10.94 13.616 10.972 13.648 ;
  LAYER M2 ;
        RECT 13.308 13.68 13.34 13.712 ;
  LAYER M2 ;
        RECT 10.94 13.744 10.972 13.776 ;
  LAYER M2 ;
        RECT 13.308 13.808 13.34 13.84 ;
  LAYER M2 ;
        RECT 10.94 13.872 10.972 13.904 ;
  LAYER M2 ;
        RECT 13.308 13.936 13.34 13.968 ;
  LAYER M2 ;
        RECT 10.94 14 10.972 14.032 ;
  LAYER M2 ;
        RECT 13.308 14.064 13.34 14.096 ;
  LAYER M2 ;
        RECT 10.94 14.128 10.972 14.16 ;
  LAYER M2 ;
        RECT 13.308 14.192 13.34 14.224 ;
  LAYER M2 ;
        RECT 10.94 14.256 10.972 14.288 ;
  LAYER M2 ;
        RECT 13.308 14.32 13.34 14.352 ;
  LAYER M2 ;
        RECT 10.94 14.384 10.972 14.416 ;
  LAYER M2 ;
        RECT 13.308 14.448 13.34 14.48 ;
  LAYER M2 ;
        RECT 10.94 14.512 10.972 14.544 ;
  LAYER M2 ;
        RECT 13.308 14.576 13.34 14.608 ;
  LAYER M2 ;
        RECT 10.94 14.64 10.972 14.672 ;
  LAYER M2 ;
        RECT 13.308 14.704 13.34 14.736 ;
  LAYER M2 ;
        RECT 10.94 14.768 10.972 14.8 ;
  LAYER M2 ;
        RECT 13.308 14.832 13.34 14.864 ;
  LAYER M2 ;
        RECT 10.94 14.896 10.972 14.928 ;
  LAYER M2 ;
        RECT 13.308 14.96 13.34 14.992 ;
  LAYER M2 ;
        RECT 10.94 15.024 10.972 15.056 ;
  LAYER M2 ;
        RECT 13.308 15.088 13.34 15.12 ;
  LAYER M2 ;
        RECT 10.94 15.152 10.972 15.184 ;
  LAYER M2 ;
        RECT 13.308 15.216 13.34 15.248 ;
  LAYER M2 ;
        RECT 10.94 15.28 10.972 15.312 ;
  LAYER M2 ;
        RECT 13.308 15.344 13.34 15.376 ;
  LAYER M2 ;
        RECT 10.94 15.408 10.972 15.44 ;
  LAYER M2 ;
        RECT 13.308 15.472 13.34 15.504 ;
  LAYER M2 ;
        RECT 10.94 15.536 10.972 15.568 ;
  LAYER M2 ;
        RECT 13.308 15.6 13.34 15.632 ;
  LAYER M2 ;
        RECT 10.94 15.664 10.972 15.696 ;
  LAYER M2 ;
        RECT 13.308 15.728 13.34 15.76 ;
  LAYER M2 ;
        RECT 10.892 13.356 13.388 15.96 ;
  LAYER M1 ;
        RECT 10.94 16.512 10.972 19.02 ;
  LAYER M3 ;
        RECT 10.94 18.968 10.972 19 ;
  LAYER M1 ;
        RECT 11.004 16.512 11.036 19.02 ;
  LAYER M3 ;
        RECT 11.004 16.532 11.036 16.564 ;
  LAYER M1 ;
        RECT 11.068 16.512 11.1 19.02 ;
  LAYER M3 ;
        RECT 11.068 18.968 11.1 19 ;
  LAYER M1 ;
        RECT 11.132 16.512 11.164 19.02 ;
  LAYER M3 ;
        RECT 11.132 16.532 11.164 16.564 ;
  LAYER M1 ;
        RECT 11.196 16.512 11.228 19.02 ;
  LAYER M3 ;
        RECT 11.196 18.968 11.228 19 ;
  LAYER M1 ;
        RECT 11.26 16.512 11.292 19.02 ;
  LAYER M3 ;
        RECT 11.26 16.532 11.292 16.564 ;
  LAYER M1 ;
        RECT 11.324 16.512 11.356 19.02 ;
  LAYER M3 ;
        RECT 11.324 18.968 11.356 19 ;
  LAYER M1 ;
        RECT 11.388 16.512 11.42 19.02 ;
  LAYER M3 ;
        RECT 11.388 16.532 11.42 16.564 ;
  LAYER M1 ;
        RECT 11.452 16.512 11.484 19.02 ;
  LAYER M3 ;
        RECT 11.452 18.968 11.484 19 ;
  LAYER M1 ;
        RECT 11.516 16.512 11.548 19.02 ;
  LAYER M3 ;
        RECT 11.516 16.532 11.548 16.564 ;
  LAYER M1 ;
        RECT 11.58 16.512 11.612 19.02 ;
  LAYER M3 ;
        RECT 11.58 18.968 11.612 19 ;
  LAYER M1 ;
        RECT 11.644 16.512 11.676 19.02 ;
  LAYER M3 ;
        RECT 11.644 16.532 11.676 16.564 ;
  LAYER M1 ;
        RECT 11.708 16.512 11.74 19.02 ;
  LAYER M3 ;
        RECT 11.708 18.968 11.74 19 ;
  LAYER M1 ;
        RECT 11.772 16.512 11.804 19.02 ;
  LAYER M3 ;
        RECT 11.772 16.532 11.804 16.564 ;
  LAYER M1 ;
        RECT 11.836 16.512 11.868 19.02 ;
  LAYER M3 ;
        RECT 11.836 18.968 11.868 19 ;
  LAYER M1 ;
        RECT 11.9 16.512 11.932 19.02 ;
  LAYER M3 ;
        RECT 11.9 16.532 11.932 16.564 ;
  LAYER M1 ;
        RECT 11.964 16.512 11.996 19.02 ;
  LAYER M3 ;
        RECT 11.964 18.968 11.996 19 ;
  LAYER M1 ;
        RECT 12.028 16.512 12.06 19.02 ;
  LAYER M3 ;
        RECT 12.028 16.532 12.06 16.564 ;
  LAYER M1 ;
        RECT 12.092 16.512 12.124 19.02 ;
  LAYER M3 ;
        RECT 12.092 18.968 12.124 19 ;
  LAYER M1 ;
        RECT 12.156 16.512 12.188 19.02 ;
  LAYER M3 ;
        RECT 12.156 16.532 12.188 16.564 ;
  LAYER M1 ;
        RECT 12.22 16.512 12.252 19.02 ;
  LAYER M3 ;
        RECT 12.22 18.968 12.252 19 ;
  LAYER M1 ;
        RECT 12.284 16.512 12.316 19.02 ;
  LAYER M3 ;
        RECT 12.284 16.532 12.316 16.564 ;
  LAYER M1 ;
        RECT 12.348 16.512 12.38 19.02 ;
  LAYER M3 ;
        RECT 12.348 18.968 12.38 19 ;
  LAYER M1 ;
        RECT 12.412 16.512 12.444 19.02 ;
  LAYER M3 ;
        RECT 12.412 16.532 12.444 16.564 ;
  LAYER M1 ;
        RECT 12.476 16.512 12.508 19.02 ;
  LAYER M3 ;
        RECT 12.476 18.968 12.508 19 ;
  LAYER M1 ;
        RECT 12.54 16.512 12.572 19.02 ;
  LAYER M3 ;
        RECT 12.54 16.532 12.572 16.564 ;
  LAYER M1 ;
        RECT 12.604 16.512 12.636 19.02 ;
  LAYER M3 ;
        RECT 12.604 18.968 12.636 19 ;
  LAYER M1 ;
        RECT 12.668 16.512 12.7 19.02 ;
  LAYER M3 ;
        RECT 12.668 16.532 12.7 16.564 ;
  LAYER M1 ;
        RECT 12.732 16.512 12.764 19.02 ;
  LAYER M3 ;
        RECT 12.732 18.968 12.764 19 ;
  LAYER M1 ;
        RECT 12.796 16.512 12.828 19.02 ;
  LAYER M3 ;
        RECT 12.796 16.532 12.828 16.564 ;
  LAYER M1 ;
        RECT 12.86 16.512 12.892 19.02 ;
  LAYER M3 ;
        RECT 12.86 18.968 12.892 19 ;
  LAYER M1 ;
        RECT 12.924 16.512 12.956 19.02 ;
  LAYER M3 ;
        RECT 12.924 16.532 12.956 16.564 ;
  LAYER M1 ;
        RECT 12.988 16.512 13.02 19.02 ;
  LAYER M3 ;
        RECT 12.988 18.968 13.02 19 ;
  LAYER M1 ;
        RECT 13.052 16.512 13.084 19.02 ;
  LAYER M3 ;
        RECT 13.052 16.532 13.084 16.564 ;
  LAYER M1 ;
        RECT 13.116 16.512 13.148 19.02 ;
  LAYER M3 ;
        RECT 13.116 18.968 13.148 19 ;
  LAYER M1 ;
        RECT 13.18 16.512 13.212 19.02 ;
  LAYER M3 ;
        RECT 13.18 16.532 13.212 16.564 ;
  LAYER M1 ;
        RECT 13.244 16.512 13.276 19.02 ;
  LAYER M3 ;
        RECT 13.244 18.968 13.276 19 ;
  LAYER M1 ;
        RECT 13.308 16.512 13.34 19.02 ;
  LAYER M3 ;
        RECT 10.94 16.596 10.972 16.628 ;
  LAYER M2 ;
        RECT 13.308 16.66 13.34 16.692 ;
  LAYER M2 ;
        RECT 10.94 16.724 10.972 16.756 ;
  LAYER M2 ;
        RECT 13.308 16.788 13.34 16.82 ;
  LAYER M2 ;
        RECT 10.94 16.852 10.972 16.884 ;
  LAYER M2 ;
        RECT 13.308 16.916 13.34 16.948 ;
  LAYER M2 ;
        RECT 10.94 16.98 10.972 17.012 ;
  LAYER M2 ;
        RECT 13.308 17.044 13.34 17.076 ;
  LAYER M2 ;
        RECT 10.94 17.108 10.972 17.14 ;
  LAYER M2 ;
        RECT 13.308 17.172 13.34 17.204 ;
  LAYER M2 ;
        RECT 10.94 17.236 10.972 17.268 ;
  LAYER M2 ;
        RECT 13.308 17.3 13.34 17.332 ;
  LAYER M2 ;
        RECT 10.94 17.364 10.972 17.396 ;
  LAYER M2 ;
        RECT 13.308 17.428 13.34 17.46 ;
  LAYER M2 ;
        RECT 10.94 17.492 10.972 17.524 ;
  LAYER M2 ;
        RECT 13.308 17.556 13.34 17.588 ;
  LAYER M2 ;
        RECT 10.94 17.62 10.972 17.652 ;
  LAYER M2 ;
        RECT 13.308 17.684 13.34 17.716 ;
  LAYER M2 ;
        RECT 10.94 17.748 10.972 17.78 ;
  LAYER M2 ;
        RECT 13.308 17.812 13.34 17.844 ;
  LAYER M2 ;
        RECT 10.94 17.876 10.972 17.908 ;
  LAYER M2 ;
        RECT 13.308 17.94 13.34 17.972 ;
  LAYER M2 ;
        RECT 10.94 18.004 10.972 18.036 ;
  LAYER M2 ;
        RECT 13.308 18.068 13.34 18.1 ;
  LAYER M2 ;
        RECT 10.94 18.132 10.972 18.164 ;
  LAYER M2 ;
        RECT 13.308 18.196 13.34 18.228 ;
  LAYER M2 ;
        RECT 10.94 18.26 10.972 18.292 ;
  LAYER M2 ;
        RECT 13.308 18.324 13.34 18.356 ;
  LAYER M2 ;
        RECT 10.94 18.388 10.972 18.42 ;
  LAYER M2 ;
        RECT 13.308 18.452 13.34 18.484 ;
  LAYER M2 ;
        RECT 10.94 18.516 10.972 18.548 ;
  LAYER M2 ;
        RECT 13.308 18.58 13.34 18.612 ;
  LAYER M2 ;
        RECT 10.94 18.644 10.972 18.676 ;
  LAYER M2 ;
        RECT 13.308 18.708 13.34 18.74 ;
  LAYER M2 ;
        RECT 10.94 18.772 10.972 18.804 ;
  LAYER M2 ;
        RECT 13.308 18.836 13.34 18.868 ;
  LAYER M2 ;
        RECT 10.892 16.464 13.388 19.068 ;
  LAYER M1 ;
        RECT 14.556 0.972 14.588 3.48 ;
  LAYER M3 ;
        RECT 14.556 3.428 14.588 3.46 ;
  LAYER M1 ;
        RECT 14.62 0.972 14.652 3.48 ;
  LAYER M3 ;
        RECT 14.62 0.992 14.652 1.024 ;
  LAYER M1 ;
        RECT 14.684 0.972 14.716 3.48 ;
  LAYER M3 ;
        RECT 14.684 3.428 14.716 3.46 ;
  LAYER M1 ;
        RECT 14.748 0.972 14.78 3.48 ;
  LAYER M3 ;
        RECT 14.748 0.992 14.78 1.024 ;
  LAYER M1 ;
        RECT 14.812 0.972 14.844 3.48 ;
  LAYER M3 ;
        RECT 14.812 3.428 14.844 3.46 ;
  LAYER M1 ;
        RECT 14.876 0.972 14.908 3.48 ;
  LAYER M3 ;
        RECT 14.876 0.992 14.908 1.024 ;
  LAYER M1 ;
        RECT 14.94 0.972 14.972 3.48 ;
  LAYER M3 ;
        RECT 14.94 3.428 14.972 3.46 ;
  LAYER M1 ;
        RECT 15.004 0.972 15.036 3.48 ;
  LAYER M3 ;
        RECT 15.004 0.992 15.036 1.024 ;
  LAYER M1 ;
        RECT 15.068 0.972 15.1 3.48 ;
  LAYER M3 ;
        RECT 15.068 3.428 15.1 3.46 ;
  LAYER M1 ;
        RECT 15.132 0.972 15.164 3.48 ;
  LAYER M3 ;
        RECT 15.132 0.992 15.164 1.024 ;
  LAYER M1 ;
        RECT 15.196 0.972 15.228 3.48 ;
  LAYER M3 ;
        RECT 15.196 3.428 15.228 3.46 ;
  LAYER M1 ;
        RECT 15.26 0.972 15.292 3.48 ;
  LAYER M3 ;
        RECT 15.26 0.992 15.292 1.024 ;
  LAYER M1 ;
        RECT 15.324 0.972 15.356 3.48 ;
  LAYER M3 ;
        RECT 15.324 3.428 15.356 3.46 ;
  LAYER M1 ;
        RECT 15.388 0.972 15.42 3.48 ;
  LAYER M3 ;
        RECT 15.388 0.992 15.42 1.024 ;
  LAYER M1 ;
        RECT 15.452 0.972 15.484 3.48 ;
  LAYER M3 ;
        RECT 15.452 3.428 15.484 3.46 ;
  LAYER M1 ;
        RECT 15.516 0.972 15.548 3.48 ;
  LAYER M3 ;
        RECT 15.516 0.992 15.548 1.024 ;
  LAYER M1 ;
        RECT 15.58 0.972 15.612 3.48 ;
  LAYER M3 ;
        RECT 15.58 3.428 15.612 3.46 ;
  LAYER M1 ;
        RECT 15.644 0.972 15.676 3.48 ;
  LAYER M3 ;
        RECT 15.644 0.992 15.676 1.024 ;
  LAYER M1 ;
        RECT 15.708 0.972 15.74 3.48 ;
  LAYER M3 ;
        RECT 15.708 3.428 15.74 3.46 ;
  LAYER M1 ;
        RECT 15.772 0.972 15.804 3.48 ;
  LAYER M3 ;
        RECT 15.772 0.992 15.804 1.024 ;
  LAYER M1 ;
        RECT 15.836 0.972 15.868 3.48 ;
  LAYER M3 ;
        RECT 15.836 3.428 15.868 3.46 ;
  LAYER M1 ;
        RECT 15.9 0.972 15.932 3.48 ;
  LAYER M3 ;
        RECT 15.9 0.992 15.932 1.024 ;
  LAYER M1 ;
        RECT 15.964 0.972 15.996 3.48 ;
  LAYER M3 ;
        RECT 15.964 3.428 15.996 3.46 ;
  LAYER M1 ;
        RECT 16.028 0.972 16.06 3.48 ;
  LAYER M3 ;
        RECT 16.028 0.992 16.06 1.024 ;
  LAYER M1 ;
        RECT 16.092 0.972 16.124 3.48 ;
  LAYER M3 ;
        RECT 16.092 3.428 16.124 3.46 ;
  LAYER M1 ;
        RECT 16.156 0.972 16.188 3.48 ;
  LAYER M3 ;
        RECT 16.156 0.992 16.188 1.024 ;
  LAYER M1 ;
        RECT 16.22 0.972 16.252 3.48 ;
  LAYER M3 ;
        RECT 16.22 3.428 16.252 3.46 ;
  LAYER M1 ;
        RECT 16.284 0.972 16.316 3.48 ;
  LAYER M3 ;
        RECT 16.284 0.992 16.316 1.024 ;
  LAYER M1 ;
        RECT 16.348 0.972 16.38 3.48 ;
  LAYER M3 ;
        RECT 16.348 3.428 16.38 3.46 ;
  LAYER M1 ;
        RECT 16.412 0.972 16.444 3.48 ;
  LAYER M3 ;
        RECT 16.412 0.992 16.444 1.024 ;
  LAYER M1 ;
        RECT 16.476 0.972 16.508 3.48 ;
  LAYER M3 ;
        RECT 16.476 3.428 16.508 3.46 ;
  LAYER M1 ;
        RECT 16.54 0.972 16.572 3.48 ;
  LAYER M3 ;
        RECT 16.54 0.992 16.572 1.024 ;
  LAYER M1 ;
        RECT 16.604 0.972 16.636 3.48 ;
  LAYER M3 ;
        RECT 16.604 3.428 16.636 3.46 ;
  LAYER M1 ;
        RECT 16.668 0.972 16.7 3.48 ;
  LAYER M3 ;
        RECT 16.668 0.992 16.7 1.024 ;
  LAYER M1 ;
        RECT 16.732 0.972 16.764 3.48 ;
  LAYER M3 ;
        RECT 16.732 3.428 16.764 3.46 ;
  LAYER M1 ;
        RECT 16.796 0.972 16.828 3.48 ;
  LAYER M3 ;
        RECT 16.796 0.992 16.828 1.024 ;
  LAYER M1 ;
        RECT 16.86 0.972 16.892 3.48 ;
  LAYER M3 ;
        RECT 16.86 3.428 16.892 3.46 ;
  LAYER M1 ;
        RECT 16.924 0.972 16.956 3.48 ;
  LAYER M3 ;
        RECT 14.556 1.056 14.588 1.088 ;
  LAYER M2 ;
        RECT 16.924 1.12 16.956 1.152 ;
  LAYER M2 ;
        RECT 14.556 1.184 14.588 1.216 ;
  LAYER M2 ;
        RECT 16.924 1.248 16.956 1.28 ;
  LAYER M2 ;
        RECT 14.556 1.312 14.588 1.344 ;
  LAYER M2 ;
        RECT 16.924 1.376 16.956 1.408 ;
  LAYER M2 ;
        RECT 14.556 1.44 14.588 1.472 ;
  LAYER M2 ;
        RECT 16.924 1.504 16.956 1.536 ;
  LAYER M2 ;
        RECT 14.556 1.568 14.588 1.6 ;
  LAYER M2 ;
        RECT 16.924 1.632 16.956 1.664 ;
  LAYER M2 ;
        RECT 14.556 1.696 14.588 1.728 ;
  LAYER M2 ;
        RECT 16.924 1.76 16.956 1.792 ;
  LAYER M2 ;
        RECT 14.556 1.824 14.588 1.856 ;
  LAYER M2 ;
        RECT 16.924 1.888 16.956 1.92 ;
  LAYER M2 ;
        RECT 14.556 1.952 14.588 1.984 ;
  LAYER M2 ;
        RECT 16.924 2.016 16.956 2.048 ;
  LAYER M2 ;
        RECT 14.556 2.08 14.588 2.112 ;
  LAYER M2 ;
        RECT 16.924 2.144 16.956 2.176 ;
  LAYER M2 ;
        RECT 14.556 2.208 14.588 2.24 ;
  LAYER M2 ;
        RECT 16.924 2.272 16.956 2.304 ;
  LAYER M2 ;
        RECT 14.556 2.336 14.588 2.368 ;
  LAYER M2 ;
        RECT 16.924 2.4 16.956 2.432 ;
  LAYER M2 ;
        RECT 14.556 2.464 14.588 2.496 ;
  LAYER M2 ;
        RECT 16.924 2.528 16.956 2.56 ;
  LAYER M2 ;
        RECT 14.556 2.592 14.588 2.624 ;
  LAYER M2 ;
        RECT 16.924 2.656 16.956 2.688 ;
  LAYER M2 ;
        RECT 14.556 2.72 14.588 2.752 ;
  LAYER M2 ;
        RECT 16.924 2.784 16.956 2.816 ;
  LAYER M2 ;
        RECT 14.556 2.848 14.588 2.88 ;
  LAYER M2 ;
        RECT 16.924 2.912 16.956 2.944 ;
  LAYER M2 ;
        RECT 14.556 2.976 14.588 3.008 ;
  LAYER M2 ;
        RECT 16.924 3.04 16.956 3.072 ;
  LAYER M2 ;
        RECT 14.556 3.104 14.588 3.136 ;
  LAYER M2 ;
        RECT 16.924 3.168 16.956 3.2 ;
  LAYER M2 ;
        RECT 14.556 3.232 14.588 3.264 ;
  LAYER M2 ;
        RECT 16.924 3.296 16.956 3.328 ;
  LAYER M2 ;
        RECT 14.508 0.924 17.004 3.528 ;
  LAYER M1 ;
        RECT 14.556 4.08 14.588 6.588 ;
  LAYER M3 ;
        RECT 14.556 6.536 14.588 6.568 ;
  LAYER M1 ;
        RECT 14.62 4.08 14.652 6.588 ;
  LAYER M3 ;
        RECT 14.62 4.1 14.652 4.132 ;
  LAYER M1 ;
        RECT 14.684 4.08 14.716 6.588 ;
  LAYER M3 ;
        RECT 14.684 6.536 14.716 6.568 ;
  LAYER M1 ;
        RECT 14.748 4.08 14.78 6.588 ;
  LAYER M3 ;
        RECT 14.748 4.1 14.78 4.132 ;
  LAYER M1 ;
        RECT 14.812 4.08 14.844 6.588 ;
  LAYER M3 ;
        RECT 14.812 6.536 14.844 6.568 ;
  LAYER M1 ;
        RECT 14.876 4.08 14.908 6.588 ;
  LAYER M3 ;
        RECT 14.876 4.1 14.908 4.132 ;
  LAYER M1 ;
        RECT 14.94 4.08 14.972 6.588 ;
  LAYER M3 ;
        RECT 14.94 6.536 14.972 6.568 ;
  LAYER M1 ;
        RECT 15.004 4.08 15.036 6.588 ;
  LAYER M3 ;
        RECT 15.004 4.1 15.036 4.132 ;
  LAYER M1 ;
        RECT 15.068 4.08 15.1 6.588 ;
  LAYER M3 ;
        RECT 15.068 6.536 15.1 6.568 ;
  LAYER M1 ;
        RECT 15.132 4.08 15.164 6.588 ;
  LAYER M3 ;
        RECT 15.132 4.1 15.164 4.132 ;
  LAYER M1 ;
        RECT 15.196 4.08 15.228 6.588 ;
  LAYER M3 ;
        RECT 15.196 6.536 15.228 6.568 ;
  LAYER M1 ;
        RECT 15.26 4.08 15.292 6.588 ;
  LAYER M3 ;
        RECT 15.26 4.1 15.292 4.132 ;
  LAYER M1 ;
        RECT 15.324 4.08 15.356 6.588 ;
  LAYER M3 ;
        RECT 15.324 6.536 15.356 6.568 ;
  LAYER M1 ;
        RECT 15.388 4.08 15.42 6.588 ;
  LAYER M3 ;
        RECT 15.388 4.1 15.42 4.132 ;
  LAYER M1 ;
        RECT 15.452 4.08 15.484 6.588 ;
  LAYER M3 ;
        RECT 15.452 6.536 15.484 6.568 ;
  LAYER M1 ;
        RECT 15.516 4.08 15.548 6.588 ;
  LAYER M3 ;
        RECT 15.516 4.1 15.548 4.132 ;
  LAYER M1 ;
        RECT 15.58 4.08 15.612 6.588 ;
  LAYER M3 ;
        RECT 15.58 6.536 15.612 6.568 ;
  LAYER M1 ;
        RECT 15.644 4.08 15.676 6.588 ;
  LAYER M3 ;
        RECT 15.644 4.1 15.676 4.132 ;
  LAYER M1 ;
        RECT 15.708 4.08 15.74 6.588 ;
  LAYER M3 ;
        RECT 15.708 6.536 15.74 6.568 ;
  LAYER M1 ;
        RECT 15.772 4.08 15.804 6.588 ;
  LAYER M3 ;
        RECT 15.772 4.1 15.804 4.132 ;
  LAYER M1 ;
        RECT 15.836 4.08 15.868 6.588 ;
  LAYER M3 ;
        RECT 15.836 6.536 15.868 6.568 ;
  LAYER M1 ;
        RECT 15.9 4.08 15.932 6.588 ;
  LAYER M3 ;
        RECT 15.9 4.1 15.932 4.132 ;
  LAYER M1 ;
        RECT 15.964 4.08 15.996 6.588 ;
  LAYER M3 ;
        RECT 15.964 6.536 15.996 6.568 ;
  LAYER M1 ;
        RECT 16.028 4.08 16.06 6.588 ;
  LAYER M3 ;
        RECT 16.028 4.1 16.06 4.132 ;
  LAYER M1 ;
        RECT 16.092 4.08 16.124 6.588 ;
  LAYER M3 ;
        RECT 16.092 6.536 16.124 6.568 ;
  LAYER M1 ;
        RECT 16.156 4.08 16.188 6.588 ;
  LAYER M3 ;
        RECT 16.156 4.1 16.188 4.132 ;
  LAYER M1 ;
        RECT 16.22 4.08 16.252 6.588 ;
  LAYER M3 ;
        RECT 16.22 6.536 16.252 6.568 ;
  LAYER M1 ;
        RECT 16.284 4.08 16.316 6.588 ;
  LAYER M3 ;
        RECT 16.284 4.1 16.316 4.132 ;
  LAYER M1 ;
        RECT 16.348 4.08 16.38 6.588 ;
  LAYER M3 ;
        RECT 16.348 6.536 16.38 6.568 ;
  LAYER M1 ;
        RECT 16.412 4.08 16.444 6.588 ;
  LAYER M3 ;
        RECT 16.412 4.1 16.444 4.132 ;
  LAYER M1 ;
        RECT 16.476 4.08 16.508 6.588 ;
  LAYER M3 ;
        RECT 16.476 6.536 16.508 6.568 ;
  LAYER M1 ;
        RECT 16.54 4.08 16.572 6.588 ;
  LAYER M3 ;
        RECT 16.54 4.1 16.572 4.132 ;
  LAYER M1 ;
        RECT 16.604 4.08 16.636 6.588 ;
  LAYER M3 ;
        RECT 16.604 6.536 16.636 6.568 ;
  LAYER M1 ;
        RECT 16.668 4.08 16.7 6.588 ;
  LAYER M3 ;
        RECT 16.668 4.1 16.7 4.132 ;
  LAYER M1 ;
        RECT 16.732 4.08 16.764 6.588 ;
  LAYER M3 ;
        RECT 16.732 6.536 16.764 6.568 ;
  LAYER M1 ;
        RECT 16.796 4.08 16.828 6.588 ;
  LAYER M3 ;
        RECT 16.796 4.1 16.828 4.132 ;
  LAYER M1 ;
        RECT 16.86 4.08 16.892 6.588 ;
  LAYER M3 ;
        RECT 16.86 6.536 16.892 6.568 ;
  LAYER M1 ;
        RECT 16.924 4.08 16.956 6.588 ;
  LAYER M3 ;
        RECT 14.556 4.164 14.588 4.196 ;
  LAYER M2 ;
        RECT 16.924 4.228 16.956 4.26 ;
  LAYER M2 ;
        RECT 14.556 4.292 14.588 4.324 ;
  LAYER M2 ;
        RECT 16.924 4.356 16.956 4.388 ;
  LAYER M2 ;
        RECT 14.556 4.42 14.588 4.452 ;
  LAYER M2 ;
        RECT 16.924 4.484 16.956 4.516 ;
  LAYER M2 ;
        RECT 14.556 4.548 14.588 4.58 ;
  LAYER M2 ;
        RECT 16.924 4.612 16.956 4.644 ;
  LAYER M2 ;
        RECT 14.556 4.676 14.588 4.708 ;
  LAYER M2 ;
        RECT 16.924 4.74 16.956 4.772 ;
  LAYER M2 ;
        RECT 14.556 4.804 14.588 4.836 ;
  LAYER M2 ;
        RECT 16.924 4.868 16.956 4.9 ;
  LAYER M2 ;
        RECT 14.556 4.932 14.588 4.964 ;
  LAYER M2 ;
        RECT 16.924 4.996 16.956 5.028 ;
  LAYER M2 ;
        RECT 14.556 5.06 14.588 5.092 ;
  LAYER M2 ;
        RECT 16.924 5.124 16.956 5.156 ;
  LAYER M2 ;
        RECT 14.556 5.188 14.588 5.22 ;
  LAYER M2 ;
        RECT 16.924 5.252 16.956 5.284 ;
  LAYER M2 ;
        RECT 14.556 5.316 14.588 5.348 ;
  LAYER M2 ;
        RECT 16.924 5.38 16.956 5.412 ;
  LAYER M2 ;
        RECT 14.556 5.444 14.588 5.476 ;
  LAYER M2 ;
        RECT 16.924 5.508 16.956 5.54 ;
  LAYER M2 ;
        RECT 14.556 5.572 14.588 5.604 ;
  LAYER M2 ;
        RECT 16.924 5.636 16.956 5.668 ;
  LAYER M2 ;
        RECT 14.556 5.7 14.588 5.732 ;
  LAYER M2 ;
        RECT 16.924 5.764 16.956 5.796 ;
  LAYER M2 ;
        RECT 14.556 5.828 14.588 5.86 ;
  LAYER M2 ;
        RECT 16.924 5.892 16.956 5.924 ;
  LAYER M2 ;
        RECT 14.556 5.956 14.588 5.988 ;
  LAYER M2 ;
        RECT 16.924 6.02 16.956 6.052 ;
  LAYER M2 ;
        RECT 14.556 6.084 14.588 6.116 ;
  LAYER M2 ;
        RECT 16.924 6.148 16.956 6.18 ;
  LAYER M2 ;
        RECT 14.556 6.212 14.588 6.244 ;
  LAYER M2 ;
        RECT 16.924 6.276 16.956 6.308 ;
  LAYER M2 ;
        RECT 14.556 6.34 14.588 6.372 ;
  LAYER M2 ;
        RECT 16.924 6.404 16.956 6.436 ;
  LAYER M2 ;
        RECT 14.508 4.032 17.004 6.636 ;
  LAYER M1 ;
        RECT 14.556 7.188 14.588 9.696 ;
  LAYER M3 ;
        RECT 14.556 9.644 14.588 9.676 ;
  LAYER M1 ;
        RECT 14.62 7.188 14.652 9.696 ;
  LAYER M3 ;
        RECT 14.62 7.208 14.652 7.24 ;
  LAYER M1 ;
        RECT 14.684 7.188 14.716 9.696 ;
  LAYER M3 ;
        RECT 14.684 9.644 14.716 9.676 ;
  LAYER M1 ;
        RECT 14.748 7.188 14.78 9.696 ;
  LAYER M3 ;
        RECT 14.748 7.208 14.78 7.24 ;
  LAYER M1 ;
        RECT 14.812 7.188 14.844 9.696 ;
  LAYER M3 ;
        RECT 14.812 9.644 14.844 9.676 ;
  LAYER M1 ;
        RECT 14.876 7.188 14.908 9.696 ;
  LAYER M3 ;
        RECT 14.876 7.208 14.908 7.24 ;
  LAYER M1 ;
        RECT 14.94 7.188 14.972 9.696 ;
  LAYER M3 ;
        RECT 14.94 9.644 14.972 9.676 ;
  LAYER M1 ;
        RECT 15.004 7.188 15.036 9.696 ;
  LAYER M3 ;
        RECT 15.004 7.208 15.036 7.24 ;
  LAYER M1 ;
        RECT 15.068 7.188 15.1 9.696 ;
  LAYER M3 ;
        RECT 15.068 9.644 15.1 9.676 ;
  LAYER M1 ;
        RECT 15.132 7.188 15.164 9.696 ;
  LAYER M3 ;
        RECT 15.132 7.208 15.164 7.24 ;
  LAYER M1 ;
        RECT 15.196 7.188 15.228 9.696 ;
  LAYER M3 ;
        RECT 15.196 9.644 15.228 9.676 ;
  LAYER M1 ;
        RECT 15.26 7.188 15.292 9.696 ;
  LAYER M3 ;
        RECT 15.26 7.208 15.292 7.24 ;
  LAYER M1 ;
        RECT 15.324 7.188 15.356 9.696 ;
  LAYER M3 ;
        RECT 15.324 9.644 15.356 9.676 ;
  LAYER M1 ;
        RECT 15.388 7.188 15.42 9.696 ;
  LAYER M3 ;
        RECT 15.388 7.208 15.42 7.24 ;
  LAYER M1 ;
        RECT 15.452 7.188 15.484 9.696 ;
  LAYER M3 ;
        RECT 15.452 9.644 15.484 9.676 ;
  LAYER M1 ;
        RECT 15.516 7.188 15.548 9.696 ;
  LAYER M3 ;
        RECT 15.516 7.208 15.548 7.24 ;
  LAYER M1 ;
        RECT 15.58 7.188 15.612 9.696 ;
  LAYER M3 ;
        RECT 15.58 9.644 15.612 9.676 ;
  LAYER M1 ;
        RECT 15.644 7.188 15.676 9.696 ;
  LAYER M3 ;
        RECT 15.644 7.208 15.676 7.24 ;
  LAYER M1 ;
        RECT 15.708 7.188 15.74 9.696 ;
  LAYER M3 ;
        RECT 15.708 9.644 15.74 9.676 ;
  LAYER M1 ;
        RECT 15.772 7.188 15.804 9.696 ;
  LAYER M3 ;
        RECT 15.772 7.208 15.804 7.24 ;
  LAYER M1 ;
        RECT 15.836 7.188 15.868 9.696 ;
  LAYER M3 ;
        RECT 15.836 9.644 15.868 9.676 ;
  LAYER M1 ;
        RECT 15.9 7.188 15.932 9.696 ;
  LAYER M3 ;
        RECT 15.9 7.208 15.932 7.24 ;
  LAYER M1 ;
        RECT 15.964 7.188 15.996 9.696 ;
  LAYER M3 ;
        RECT 15.964 9.644 15.996 9.676 ;
  LAYER M1 ;
        RECT 16.028 7.188 16.06 9.696 ;
  LAYER M3 ;
        RECT 16.028 7.208 16.06 7.24 ;
  LAYER M1 ;
        RECT 16.092 7.188 16.124 9.696 ;
  LAYER M3 ;
        RECT 16.092 9.644 16.124 9.676 ;
  LAYER M1 ;
        RECT 16.156 7.188 16.188 9.696 ;
  LAYER M3 ;
        RECT 16.156 7.208 16.188 7.24 ;
  LAYER M1 ;
        RECT 16.22 7.188 16.252 9.696 ;
  LAYER M3 ;
        RECT 16.22 9.644 16.252 9.676 ;
  LAYER M1 ;
        RECT 16.284 7.188 16.316 9.696 ;
  LAYER M3 ;
        RECT 16.284 7.208 16.316 7.24 ;
  LAYER M1 ;
        RECT 16.348 7.188 16.38 9.696 ;
  LAYER M3 ;
        RECT 16.348 9.644 16.38 9.676 ;
  LAYER M1 ;
        RECT 16.412 7.188 16.444 9.696 ;
  LAYER M3 ;
        RECT 16.412 7.208 16.444 7.24 ;
  LAYER M1 ;
        RECT 16.476 7.188 16.508 9.696 ;
  LAYER M3 ;
        RECT 16.476 9.644 16.508 9.676 ;
  LAYER M1 ;
        RECT 16.54 7.188 16.572 9.696 ;
  LAYER M3 ;
        RECT 16.54 7.208 16.572 7.24 ;
  LAYER M1 ;
        RECT 16.604 7.188 16.636 9.696 ;
  LAYER M3 ;
        RECT 16.604 9.644 16.636 9.676 ;
  LAYER M1 ;
        RECT 16.668 7.188 16.7 9.696 ;
  LAYER M3 ;
        RECT 16.668 7.208 16.7 7.24 ;
  LAYER M1 ;
        RECT 16.732 7.188 16.764 9.696 ;
  LAYER M3 ;
        RECT 16.732 9.644 16.764 9.676 ;
  LAYER M1 ;
        RECT 16.796 7.188 16.828 9.696 ;
  LAYER M3 ;
        RECT 16.796 7.208 16.828 7.24 ;
  LAYER M1 ;
        RECT 16.86 7.188 16.892 9.696 ;
  LAYER M3 ;
        RECT 16.86 9.644 16.892 9.676 ;
  LAYER M1 ;
        RECT 16.924 7.188 16.956 9.696 ;
  LAYER M3 ;
        RECT 14.556 7.272 14.588 7.304 ;
  LAYER M2 ;
        RECT 16.924 7.336 16.956 7.368 ;
  LAYER M2 ;
        RECT 14.556 7.4 14.588 7.432 ;
  LAYER M2 ;
        RECT 16.924 7.464 16.956 7.496 ;
  LAYER M2 ;
        RECT 14.556 7.528 14.588 7.56 ;
  LAYER M2 ;
        RECT 16.924 7.592 16.956 7.624 ;
  LAYER M2 ;
        RECT 14.556 7.656 14.588 7.688 ;
  LAYER M2 ;
        RECT 16.924 7.72 16.956 7.752 ;
  LAYER M2 ;
        RECT 14.556 7.784 14.588 7.816 ;
  LAYER M2 ;
        RECT 16.924 7.848 16.956 7.88 ;
  LAYER M2 ;
        RECT 14.556 7.912 14.588 7.944 ;
  LAYER M2 ;
        RECT 16.924 7.976 16.956 8.008 ;
  LAYER M2 ;
        RECT 14.556 8.04 14.588 8.072 ;
  LAYER M2 ;
        RECT 16.924 8.104 16.956 8.136 ;
  LAYER M2 ;
        RECT 14.556 8.168 14.588 8.2 ;
  LAYER M2 ;
        RECT 16.924 8.232 16.956 8.264 ;
  LAYER M2 ;
        RECT 14.556 8.296 14.588 8.328 ;
  LAYER M2 ;
        RECT 16.924 8.36 16.956 8.392 ;
  LAYER M2 ;
        RECT 14.556 8.424 14.588 8.456 ;
  LAYER M2 ;
        RECT 16.924 8.488 16.956 8.52 ;
  LAYER M2 ;
        RECT 14.556 8.552 14.588 8.584 ;
  LAYER M2 ;
        RECT 16.924 8.616 16.956 8.648 ;
  LAYER M2 ;
        RECT 14.556 8.68 14.588 8.712 ;
  LAYER M2 ;
        RECT 16.924 8.744 16.956 8.776 ;
  LAYER M2 ;
        RECT 14.556 8.808 14.588 8.84 ;
  LAYER M2 ;
        RECT 16.924 8.872 16.956 8.904 ;
  LAYER M2 ;
        RECT 14.556 8.936 14.588 8.968 ;
  LAYER M2 ;
        RECT 16.924 9 16.956 9.032 ;
  LAYER M2 ;
        RECT 14.556 9.064 14.588 9.096 ;
  LAYER M2 ;
        RECT 16.924 9.128 16.956 9.16 ;
  LAYER M2 ;
        RECT 14.556 9.192 14.588 9.224 ;
  LAYER M2 ;
        RECT 16.924 9.256 16.956 9.288 ;
  LAYER M2 ;
        RECT 14.556 9.32 14.588 9.352 ;
  LAYER M2 ;
        RECT 16.924 9.384 16.956 9.416 ;
  LAYER M2 ;
        RECT 14.556 9.448 14.588 9.48 ;
  LAYER M2 ;
        RECT 16.924 9.512 16.956 9.544 ;
  LAYER M2 ;
        RECT 14.508 7.14 17.004 9.744 ;
  LAYER M1 ;
        RECT 14.556 10.296 14.588 12.804 ;
  LAYER M3 ;
        RECT 14.556 12.752 14.588 12.784 ;
  LAYER M1 ;
        RECT 14.62 10.296 14.652 12.804 ;
  LAYER M3 ;
        RECT 14.62 10.316 14.652 10.348 ;
  LAYER M1 ;
        RECT 14.684 10.296 14.716 12.804 ;
  LAYER M3 ;
        RECT 14.684 12.752 14.716 12.784 ;
  LAYER M1 ;
        RECT 14.748 10.296 14.78 12.804 ;
  LAYER M3 ;
        RECT 14.748 10.316 14.78 10.348 ;
  LAYER M1 ;
        RECT 14.812 10.296 14.844 12.804 ;
  LAYER M3 ;
        RECT 14.812 12.752 14.844 12.784 ;
  LAYER M1 ;
        RECT 14.876 10.296 14.908 12.804 ;
  LAYER M3 ;
        RECT 14.876 10.316 14.908 10.348 ;
  LAYER M1 ;
        RECT 14.94 10.296 14.972 12.804 ;
  LAYER M3 ;
        RECT 14.94 12.752 14.972 12.784 ;
  LAYER M1 ;
        RECT 15.004 10.296 15.036 12.804 ;
  LAYER M3 ;
        RECT 15.004 10.316 15.036 10.348 ;
  LAYER M1 ;
        RECT 15.068 10.296 15.1 12.804 ;
  LAYER M3 ;
        RECT 15.068 12.752 15.1 12.784 ;
  LAYER M1 ;
        RECT 15.132 10.296 15.164 12.804 ;
  LAYER M3 ;
        RECT 15.132 10.316 15.164 10.348 ;
  LAYER M1 ;
        RECT 15.196 10.296 15.228 12.804 ;
  LAYER M3 ;
        RECT 15.196 12.752 15.228 12.784 ;
  LAYER M1 ;
        RECT 15.26 10.296 15.292 12.804 ;
  LAYER M3 ;
        RECT 15.26 10.316 15.292 10.348 ;
  LAYER M1 ;
        RECT 15.324 10.296 15.356 12.804 ;
  LAYER M3 ;
        RECT 15.324 12.752 15.356 12.784 ;
  LAYER M1 ;
        RECT 15.388 10.296 15.42 12.804 ;
  LAYER M3 ;
        RECT 15.388 10.316 15.42 10.348 ;
  LAYER M1 ;
        RECT 15.452 10.296 15.484 12.804 ;
  LAYER M3 ;
        RECT 15.452 12.752 15.484 12.784 ;
  LAYER M1 ;
        RECT 15.516 10.296 15.548 12.804 ;
  LAYER M3 ;
        RECT 15.516 10.316 15.548 10.348 ;
  LAYER M1 ;
        RECT 15.58 10.296 15.612 12.804 ;
  LAYER M3 ;
        RECT 15.58 12.752 15.612 12.784 ;
  LAYER M1 ;
        RECT 15.644 10.296 15.676 12.804 ;
  LAYER M3 ;
        RECT 15.644 10.316 15.676 10.348 ;
  LAYER M1 ;
        RECT 15.708 10.296 15.74 12.804 ;
  LAYER M3 ;
        RECT 15.708 12.752 15.74 12.784 ;
  LAYER M1 ;
        RECT 15.772 10.296 15.804 12.804 ;
  LAYER M3 ;
        RECT 15.772 10.316 15.804 10.348 ;
  LAYER M1 ;
        RECT 15.836 10.296 15.868 12.804 ;
  LAYER M3 ;
        RECT 15.836 12.752 15.868 12.784 ;
  LAYER M1 ;
        RECT 15.9 10.296 15.932 12.804 ;
  LAYER M3 ;
        RECT 15.9 10.316 15.932 10.348 ;
  LAYER M1 ;
        RECT 15.964 10.296 15.996 12.804 ;
  LAYER M3 ;
        RECT 15.964 12.752 15.996 12.784 ;
  LAYER M1 ;
        RECT 16.028 10.296 16.06 12.804 ;
  LAYER M3 ;
        RECT 16.028 10.316 16.06 10.348 ;
  LAYER M1 ;
        RECT 16.092 10.296 16.124 12.804 ;
  LAYER M3 ;
        RECT 16.092 12.752 16.124 12.784 ;
  LAYER M1 ;
        RECT 16.156 10.296 16.188 12.804 ;
  LAYER M3 ;
        RECT 16.156 10.316 16.188 10.348 ;
  LAYER M1 ;
        RECT 16.22 10.296 16.252 12.804 ;
  LAYER M3 ;
        RECT 16.22 12.752 16.252 12.784 ;
  LAYER M1 ;
        RECT 16.284 10.296 16.316 12.804 ;
  LAYER M3 ;
        RECT 16.284 10.316 16.316 10.348 ;
  LAYER M1 ;
        RECT 16.348 10.296 16.38 12.804 ;
  LAYER M3 ;
        RECT 16.348 12.752 16.38 12.784 ;
  LAYER M1 ;
        RECT 16.412 10.296 16.444 12.804 ;
  LAYER M3 ;
        RECT 16.412 10.316 16.444 10.348 ;
  LAYER M1 ;
        RECT 16.476 10.296 16.508 12.804 ;
  LAYER M3 ;
        RECT 16.476 12.752 16.508 12.784 ;
  LAYER M1 ;
        RECT 16.54 10.296 16.572 12.804 ;
  LAYER M3 ;
        RECT 16.54 10.316 16.572 10.348 ;
  LAYER M1 ;
        RECT 16.604 10.296 16.636 12.804 ;
  LAYER M3 ;
        RECT 16.604 12.752 16.636 12.784 ;
  LAYER M1 ;
        RECT 16.668 10.296 16.7 12.804 ;
  LAYER M3 ;
        RECT 16.668 10.316 16.7 10.348 ;
  LAYER M1 ;
        RECT 16.732 10.296 16.764 12.804 ;
  LAYER M3 ;
        RECT 16.732 12.752 16.764 12.784 ;
  LAYER M1 ;
        RECT 16.796 10.296 16.828 12.804 ;
  LAYER M3 ;
        RECT 16.796 10.316 16.828 10.348 ;
  LAYER M1 ;
        RECT 16.86 10.296 16.892 12.804 ;
  LAYER M3 ;
        RECT 16.86 12.752 16.892 12.784 ;
  LAYER M1 ;
        RECT 16.924 10.296 16.956 12.804 ;
  LAYER M3 ;
        RECT 14.556 10.38 14.588 10.412 ;
  LAYER M2 ;
        RECT 16.924 10.444 16.956 10.476 ;
  LAYER M2 ;
        RECT 14.556 10.508 14.588 10.54 ;
  LAYER M2 ;
        RECT 16.924 10.572 16.956 10.604 ;
  LAYER M2 ;
        RECT 14.556 10.636 14.588 10.668 ;
  LAYER M2 ;
        RECT 16.924 10.7 16.956 10.732 ;
  LAYER M2 ;
        RECT 14.556 10.764 14.588 10.796 ;
  LAYER M2 ;
        RECT 16.924 10.828 16.956 10.86 ;
  LAYER M2 ;
        RECT 14.556 10.892 14.588 10.924 ;
  LAYER M2 ;
        RECT 16.924 10.956 16.956 10.988 ;
  LAYER M2 ;
        RECT 14.556 11.02 14.588 11.052 ;
  LAYER M2 ;
        RECT 16.924 11.084 16.956 11.116 ;
  LAYER M2 ;
        RECT 14.556 11.148 14.588 11.18 ;
  LAYER M2 ;
        RECT 16.924 11.212 16.956 11.244 ;
  LAYER M2 ;
        RECT 14.556 11.276 14.588 11.308 ;
  LAYER M2 ;
        RECT 16.924 11.34 16.956 11.372 ;
  LAYER M2 ;
        RECT 14.556 11.404 14.588 11.436 ;
  LAYER M2 ;
        RECT 16.924 11.468 16.956 11.5 ;
  LAYER M2 ;
        RECT 14.556 11.532 14.588 11.564 ;
  LAYER M2 ;
        RECT 16.924 11.596 16.956 11.628 ;
  LAYER M2 ;
        RECT 14.556 11.66 14.588 11.692 ;
  LAYER M2 ;
        RECT 16.924 11.724 16.956 11.756 ;
  LAYER M2 ;
        RECT 14.556 11.788 14.588 11.82 ;
  LAYER M2 ;
        RECT 16.924 11.852 16.956 11.884 ;
  LAYER M2 ;
        RECT 14.556 11.916 14.588 11.948 ;
  LAYER M2 ;
        RECT 16.924 11.98 16.956 12.012 ;
  LAYER M2 ;
        RECT 14.556 12.044 14.588 12.076 ;
  LAYER M2 ;
        RECT 16.924 12.108 16.956 12.14 ;
  LAYER M2 ;
        RECT 14.556 12.172 14.588 12.204 ;
  LAYER M2 ;
        RECT 16.924 12.236 16.956 12.268 ;
  LAYER M2 ;
        RECT 14.556 12.3 14.588 12.332 ;
  LAYER M2 ;
        RECT 16.924 12.364 16.956 12.396 ;
  LAYER M2 ;
        RECT 14.556 12.428 14.588 12.46 ;
  LAYER M2 ;
        RECT 16.924 12.492 16.956 12.524 ;
  LAYER M2 ;
        RECT 14.556 12.556 14.588 12.588 ;
  LAYER M2 ;
        RECT 16.924 12.62 16.956 12.652 ;
  LAYER M2 ;
        RECT 14.508 10.248 17.004 12.852 ;
  LAYER M1 ;
        RECT 14.556 13.404 14.588 15.912 ;
  LAYER M3 ;
        RECT 14.556 15.86 14.588 15.892 ;
  LAYER M1 ;
        RECT 14.62 13.404 14.652 15.912 ;
  LAYER M3 ;
        RECT 14.62 13.424 14.652 13.456 ;
  LAYER M1 ;
        RECT 14.684 13.404 14.716 15.912 ;
  LAYER M3 ;
        RECT 14.684 15.86 14.716 15.892 ;
  LAYER M1 ;
        RECT 14.748 13.404 14.78 15.912 ;
  LAYER M3 ;
        RECT 14.748 13.424 14.78 13.456 ;
  LAYER M1 ;
        RECT 14.812 13.404 14.844 15.912 ;
  LAYER M3 ;
        RECT 14.812 15.86 14.844 15.892 ;
  LAYER M1 ;
        RECT 14.876 13.404 14.908 15.912 ;
  LAYER M3 ;
        RECT 14.876 13.424 14.908 13.456 ;
  LAYER M1 ;
        RECT 14.94 13.404 14.972 15.912 ;
  LAYER M3 ;
        RECT 14.94 15.86 14.972 15.892 ;
  LAYER M1 ;
        RECT 15.004 13.404 15.036 15.912 ;
  LAYER M3 ;
        RECT 15.004 13.424 15.036 13.456 ;
  LAYER M1 ;
        RECT 15.068 13.404 15.1 15.912 ;
  LAYER M3 ;
        RECT 15.068 15.86 15.1 15.892 ;
  LAYER M1 ;
        RECT 15.132 13.404 15.164 15.912 ;
  LAYER M3 ;
        RECT 15.132 13.424 15.164 13.456 ;
  LAYER M1 ;
        RECT 15.196 13.404 15.228 15.912 ;
  LAYER M3 ;
        RECT 15.196 15.86 15.228 15.892 ;
  LAYER M1 ;
        RECT 15.26 13.404 15.292 15.912 ;
  LAYER M3 ;
        RECT 15.26 13.424 15.292 13.456 ;
  LAYER M1 ;
        RECT 15.324 13.404 15.356 15.912 ;
  LAYER M3 ;
        RECT 15.324 15.86 15.356 15.892 ;
  LAYER M1 ;
        RECT 15.388 13.404 15.42 15.912 ;
  LAYER M3 ;
        RECT 15.388 13.424 15.42 13.456 ;
  LAYER M1 ;
        RECT 15.452 13.404 15.484 15.912 ;
  LAYER M3 ;
        RECT 15.452 15.86 15.484 15.892 ;
  LAYER M1 ;
        RECT 15.516 13.404 15.548 15.912 ;
  LAYER M3 ;
        RECT 15.516 13.424 15.548 13.456 ;
  LAYER M1 ;
        RECT 15.58 13.404 15.612 15.912 ;
  LAYER M3 ;
        RECT 15.58 15.86 15.612 15.892 ;
  LAYER M1 ;
        RECT 15.644 13.404 15.676 15.912 ;
  LAYER M3 ;
        RECT 15.644 13.424 15.676 13.456 ;
  LAYER M1 ;
        RECT 15.708 13.404 15.74 15.912 ;
  LAYER M3 ;
        RECT 15.708 15.86 15.74 15.892 ;
  LAYER M1 ;
        RECT 15.772 13.404 15.804 15.912 ;
  LAYER M3 ;
        RECT 15.772 13.424 15.804 13.456 ;
  LAYER M1 ;
        RECT 15.836 13.404 15.868 15.912 ;
  LAYER M3 ;
        RECT 15.836 15.86 15.868 15.892 ;
  LAYER M1 ;
        RECT 15.9 13.404 15.932 15.912 ;
  LAYER M3 ;
        RECT 15.9 13.424 15.932 13.456 ;
  LAYER M1 ;
        RECT 15.964 13.404 15.996 15.912 ;
  LAYER M3 ;
        RECT 15.964 15.86 15.996 15.892 ;
  LAYER M1 ;
        RECT 16.028 13.404 16.06 15.912 ;
  LAYER M3 ;
        RECT 16.028 13.424 16.06 13.456 ;
  LAYER M1 ;
        RECT 16.092 13.404 16.124 15.912 ;
  LAYER M3 ;
        RECT 16.092 15.86 16.124 15.892 ;
  LAYER M1 ;
        RECT 16.156 13.404 16.188 15.912 ;
  LAYER M3 ;
        RECT 16.156 13.424 16.188 13.456 ;
  LAYER M1 ;
        RECT 16.22 13.404 16.252 15.912 ;
  LAYER M3 ;
        RECT 16.22 15.86 16.252 15.892 ;
  LAYER M1 ;
        RECT 16.284 13.404 16.316 15.912 ;
  LAYER M3 ;
        RECT 16.284 13.424 16.316 13.456 ;
  LAYER M1 ;
        RECT 16.348 13.404 16.38 15.912 ;
  LAYER M3 ;
        RECT 16.348 15.86 16.38 15.892 ;
  LAYER M1 ;
        RECT 16.412 13.404 16.444 15.912 ;
  LAYER M3 ;
        RECT 16.412 13.424 16.444 13.456 ;
  LAYER M1 ;
        RECT 16.476 13.404 16.508 15.912 ;
  LAYER M3 ;
        RECT 16.476 15.86 16.508 15.892 ;
  LAYER M1 ;
        RECT 16.54 13.404 16.572 15.912 ;
  LAYER M3 ;
        RECT 16.54 13.424 16.572 13.456 ;
  LAYER M1 ;
        RECT 16.604 13.404 16.636 15.912 ;
  LAYER M3 ;
        RECT 16.604 15.86 16.636 15.892 ;
  LAYER M1 ;
        RECT 16.668 13.404 16.7 15.912 ;
  LAYER M3 ;
        RECT 16.668 13.424 16.7 13.456 ;
  LAYER M1 ;
        RECT 16.732 13.404 16.764 15.912 ;
  LAYER M3 ;
        RECT 16.732 15.86 16.764 15.892 ;
  LAYER M1 ;
        RECT 16.796 13.404 16.828 15.912 ;
  LAYER M3 ;
        RECT 16.796 13.424 16.828 13.456 ;
  LAYER M1 ;
        RECT 16.86 13.404 16.892 15.912 ;
  LAYER M3 ;
        RECT 16.86 15.86 16.892 15.892 ;
  LAYER M1 ;
        RECT 16.924 13.404 16.956 15.912 ;
  LAYER M3 ;
        RECT 14.556 13.488 14.588 13.52 ;
  LAYER M2 ;
        RECT 16.924 13.552 16.956 13.584 ;
  LAYER M2 ;
        RECT 14.556 13.616 14.588 13.648 ;
  LAYER M2 ;
        RECT 16.924 13.68 16.956 13.712 ;
  LAYER M2 ;
        RECT 14.556 13.744 14.588 13.776 ;
  LAYER M2 ;
        RECT 16.924 13.808 16.956 13.84 ;
  LAYER M2 ;
        RECT 14.556 13.872 14.588 13.904 ;
  LAYER M2 ;
        RECT 16.924 13.936 16.956 13.968 ;
  LAYER M2 ;
        RECT 14.556 14 14.588 14.032 ;
  LAYER M2 ;
        RECT 16.924 14.064 16.956 14.096 ;
  LAYER M2 ;
        RECT 14.556 14.128 14.588 14.16 ;
  LAYER M2 ;
        RECT 16.924 14.192 16.956 14.224 ;
  LAYER M2 ;
        RECT 14.556 14.256 14.588 14.288 ;
  LAYER M2 ;
        RECT 16.924 14.32 16.956 14.352 ;
  LAYER M2 ;
        RECT 14.556 14.384 14.588 14.416 ;
  LAYER M2 ;
        RECT 16.924 14.448 16.956 14.48 ;
  LAYER M2 ;
        RECT 14.556 14.512 14.588 14.544 ;
  LAYER M2 ;
        RECT 16.924 14.576 16.956 14.608 ;
  LAYER M2 ;
        RECT 14.556 14.64 14.588 14.672 ;
  LAYER M2 ;
        RECT 16.924 14.704 16.956 14.736 ;
  LAYER M2 ;
        RECT 14.556 14.768 14.588 14.8 ;
  LAYER M2 ;
        RECT 16.924 14.832 16.956 14.864 ;
  LAYER M2 ;
        RECT 14.556 14.896 14.588 14.928 ;
  LAYER M2 ;
        RECT 16.924 14.96 16.956 14.992 ;
  LAYER M2 ;
        RECT 14.556 15.024 14.588 15.056 ;
  LAYER M2 ;
        RECT 16.924 15.088 16.956 15.12 ;
  LAYER M2 ;
        RECT 14.556 15.152 14.588 15.184 ;
  LAYER M2 ;
        RECT 16.924 15.216 16.956 15.248 ;
  LAYER M2 ;
        RECT 14.556 15.28 14.588 15.312 ;
  LAYER M2 ;
        RECT 16.924 15.344 16.956 15.376 ;
  LAYER M2 ;
        RECT 14.556 15.408 14.588 15.44 ;
  LAYER M2 ;
        RECT 16.924 15.472 16.956 15.504 ;
  LAYER M2 ;
        RECT 14.556 15.536 14.588 15.568 ;
  LAYER M2 ;
        RECT 16.924 15.6 16.956 15.632 ;
  LAYER M2 ;
        RECT 14.556 15.664 14.588 15.696 ;
  LAYER M2 ;
        RECT 16.924 15.728 16.956 15.76 ;
  LAYER M2 ;
        RECT 14.508 13.356 17.004 15.96 ;
  LAYER M1 ;
        RECT 14.556 16.512 14.588 19.02 ;
  LAYER M3 ;
        RECT 14.556 18.968 14.588 19 ;
  LAYER M1 ;
        RECT 14.62 16.512 14.652 19.02 ;
  LAYER M3 ;
        RECT 14.62 16.532 14.652 16.564 ;
  LAYER M1 ;
        RECT 14.684 16.512 14.716 19.02 ;
  LAYER M3 ;
        RECT 14.684 18.968 14.716 19 ;
  LAYER M1 ;
        RECT 14.748 16.512 14.78 19.02 ;
  LAYER M3 ;
        RECT 14.748 16.532 14.78 16.564 ;
  LAYER M1 ;
        RECT 14.812 16.512 14.844 19.02 ;
  LAYER M3 ;
        RECT 14.812 18.968 14.844 19 ;
  LAYER M1 ;
        RECT 14.876 16.512 14.908 19.02 ;
  LAYER M3 ;
        RECT 14.876 16.532 14.908 16.564 ;
  LAYER M1 ;
        RECT 14.94 16.512 14.972 19.02 ;
  LAYER M3 ;
        RECT 14.94 18.968 14.972 19 ;
  LAYER M1 ;
        RECT 15.004 16.512 15.036 19.02 ;
  LAYER M3 ;
        RECT 15.004 16.532 15.036 16.564 ;
  LAYER M1 ;
        RECT 15.068 16.512 15.1 19.02 ;
  LAYER M3 ;
        RECT 15.068 18.968 15.1 19 ;
  LAYER M1 ;
        RECT 15.132 16.512 15.164 19.02 ;
  LAYER M3 ;
        RECT 15.132 16.532 15.164 16.564 ;
  LAYER M1 ;
        RECT 15.196 16.512 15.228 19.02 ;
  LAYER M3 ;
        RECT 15.196 18.968 15.228 19 ;
  LAYER M1 ;
        RECT 15.26 16.512 15.292 19.02 ;
  LAYER M3 ;
        RECT 15.26 16.532 15.292 16.564 ;
  LAYER M1 ;
        RECT 15.324 16.512 15.356 19.02 ;
  LAYER M3 ;
        RECT 15.324 18.968 15.356 19 ;
  LAYER M1 ;
        RECT 15.388 16.512 15.42 19.02 ;
  LAYER M3 ;
        RECT 15.388 16.532 15.42 16.564 ;
  LAYER M1 ;
        RECT 15.452 16.512 15.484 19.02 ;
  LAYER M3 ;
        RECT 15.452 18.968 15.484 19 ;
  LAYER M1 ;
        RECT 15.516 16.512 15.548 19.02 ;
  LAYER M3 ;
        RECT 15.516 16.532 15.548 16.564 ;
  LAYER M1 ;
        RECT 15.58 16.512 15.612 19.02 ;
  LAYER M3 ;
        RECT 15.58 18.968 15.612 19 ;
  LAYER M1 ;
        RECT 15.644 16.512 15.676 19.02 ;
  LAYER M3 ;
        RECT 15.644 16.532 15.676 16.564 ;
  LAYER M1 ;
        RECT 15.708 16.512 15.74 19.02 ;
  LAYER M3 ;
        RECT 15.708 18.968 15.74 19 ;
  LAYER M1 ;
        RECT 15.772 16.512 15.804 19.02 ;
  LAYER M3 ;
        RECT 15.772 16.532 15.804 16.564 ;
  LAYER M1 ;
        RECT 15.836 16.512 15.868 19.02 ;
  LAYER M3 ;
        RECT 15.836 18.968 15.868 19 ;
  LAYER M1 ;
        RECT 15.9 16.512 15.932 19.02 ;
  LAYER M3 ;
        RECT 15.9 16.532 15.932 16.564 ;
  LAYER M1 ;
        RECT 15.964 16.512 15.996 19.02 ;
  LAYER M3 ;
        RECT 15.964 18.968 15.996 19 ;
  LAYER M1 ;
        RECT 16.028 16.512 16.06 19.02 ;
  LAYER M3 ;
        RECT 16.028 16.532 16.06 16.564 ;
  LAYER M1 ;
        RECT 16.092 16.512 16.124 19.02 ;
  LAYER M3 ;
        RECT 16.092 18.968 16.124 19 ;
  LAYER M1 ;
        RECT 16.156 16.512 16.188 19.02 ;
  LAYER M3 ;
        RECT 16.156 16.532 16.188 16.564 ;
  LAYER M1 ;
        RECT 16.22 16.512 16.252 19.02 ;
  LAYER M3 ;
        RECT 16.22 18.968 16.252 19 ;
  LAYER M1 ;
        RECT 16.284 16.512 16.316 19.02 ;
  LAYER M3 ;
        RECT 16.284 16.532 16.316 16.564 ;
  LAYER M1 ;
        RECT 16.348 16.512 16.38 19.02 ;
  LAYER M3 ;
        RECT 16.348 18.968 16.38 19 ;
  LAYER M1 ;
        RECT 16.412 16.512 16.444 19.02 ;
  LAYER M3 ;
        RECT 16.412 16.532 16.444 16.564 ;
  LAYER M1 ;
        RECT 16.476 16.512 16.508 19.02 ;
  LAYER M3 ;
        RECT 16.476 18.968 16.508 19 ;
  LAYER M1 ;
        RECT 16.54 16.512 16.572 19.02 ;
  LAYER M3 ;
        RECT 16.54 16.532 16.572 16.564 ;
  LAYER M1 ;
        RECT 16.604 16.512 16.636 19.02 ;
  LAYER M3 ;
        RECT 16.604 18.968 16.636 19 ;
  LAYER M1 ;
        RECT 16.668 16.512 16.7 19.02 ;
  LAYER M3 ;
        RECT 16.668 16.532 16.7 16.564 ;
  LAYER M1 ;
        RECT 16.732 16.512 16.764 19.02 ;
  LAYER M3 ;
        RECT 16.732 18.968 16.764 19 ;
  LAYER M1 ;
        RECT 16.796 16.512 16.828 19.02 ;
  LAYER M3 ;
        RECT 16.796 16.532 16.828 16.564 ;
  LAYER M1 ;
        RECT 16.86 16.512 16.892 19.02 ;
  LAYER M3 ;
        RECT 16.86 18.968 16.892 19 ;
  LAYER M1 ;
        RECT 16.924 16.512 16.956 19.02 ;
  LAYER M3 ;
        RECT 14.556 16.596 14.588 16.628 ;
  LAYER M2 ;
        RECT 16.924 16.66 16.956 16.692 ;
  LAYER M2 ;
        RECT 14.556 16.724 14.588 16.756 ;
  LAYER M2 ;
        RECT 16.924 16.788 16.956 16.82 ;
  LAYER M2 ;
        RECT 14.556 16.852 14.588 16.884 ;
  LAYER M2 ;
        RECT 16.924 16.916 16.956 16.948 ;
  LAYER M2 ;
        RECT 14.556 16.98 14.588 17.012 ;
  LAYER M2 ;
        RECT 16.924 17.044 16.956 17.076 ;
  LAYER M2 ;
        RECT 14.556 17.108 14.588 17.14 ;
  LAYER M2 ;
        RECT 16.924 17.172 16.956 17.204 ;
  LAYER M2 ;
        RECT 14.556 17.236 14.588 17.268 ;
  LAYER M2 ;
        RECT 16.924 17.3 16.956 17.332 ;
  LAYER M2 ;
        RECT 14.556 17.364 14.588 17.396 ;
  LAYER M2 ;
        RECT 16.924 17.428 16.956 17.46 ;
  LAYER M2 ;
        RECT 14.556 17.492 14.588 17.524 ;
  LAYER M2 ;
        RECT 16.924 17.556 16.956 17.588 ;
  LAYER M2 ;
        RECT 14.556 17.62 14.588 17.652 ;
  LAYER M2 ;
        RECT 16.924 17.684 16.956 17.716 ;
  LAYER M2 ;
        RECT 14.556 17.748 14.588 17.78 ;
  LAYER M2 ;
        RECT 16.924 17.812 16.956 17.844 ;
  LAYER M2 ;
        RECT 14.556 17.876 14.588 17.908 ;
  LAYER M2 ;
        RECT 16.924 17.94 16.956 17.972 ;
  LAYER M2 ;
        RECT 14.556 18.004 14.588 18.036 ;
  LAYER M2 ;
        RECT 16.924 18.068 16.956 18.1 ;
  LAYER M2 ;
        RECT 14.556 18.132 14.588 18.164 ;
  LAYER M2 ;
        RECT 16.924 18.196 16.956 18.228 ;
  LAYER M2 ;
        RECT 14.556 18.26 14.588 18.292 ;
  LAYER M2 ;
        RECT 16.924 18.324 16.956 18.356 ;
  LAYER M2 ;
        RECT 14.556 18.388 14.588 18.42 ;
  LAYER M2 ;
        RECT 16.924 18.452 16.956 18.484 ;
  LAYER M2 ;
        RECT 14.556 18.516 14.588 18.548 ;
  LAYER M2 ;
        RECT 16.924 18.58 16.956 18.612 ;
  LAYER M2 ;
        RECT 14.556 18.644 14.588 18.676 ;
  LAYER M2 ;
        RECT 16.924 18.708 16.956 18.74 ;
  LAYER M2 ;
        RECT 14.556 18.772 14.588 18.804 ;
  LAYER M2 ;
        RECT 16.924 18.836 16.956 18.868 ;
  LAYER M2 ;
        RECT 14.508 16.464 17.004 19.068 ;
  END 
END Cap_30fF_Cap_60fF
