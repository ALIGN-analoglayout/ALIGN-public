VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Cap_10f_1x1
  ORIGIN 0 0 ;
  FOREIGN Cap_10f_1x1 0 0 ;
  SIZE 2.214 BY 2.214 ;
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 2.196 2.214 2.214 ;
    END
  END PLUS
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0 2.214 0.018 ;
    END
  END MINUS
  OBS
      LAYER M1 ;
        RECT 0 0 2.214 2.214 ;
      END
  OBS
      LAYER M2 ;
        RECT 0.018 0.018 2.196 2.196 ;
      END
  OBS
      LAYER M3 ;
        RECT 0 0 2.214 2.214 ;
      END
END Cap_10f_1x1

MACRO Switch_NMOS_10_1x1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_10_1x1 0 0 ;
  SIZE 0.432 BY 0.402 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.064 0.284 0.082 ;
    END
  END S
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.148 0.192 0.392 0.21 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.128 0.338 0.146 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 0.384 0.432 0.402 ;
    END
  END VDD

END Switch_NMOS_10_1x1


END LIBRARY
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

VIA M2_M1_0
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0.005 0.005 0 ;
  ROWCOL 1 1 ;
END M2_M1_0

VIA M2_M1_1
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0.005 0.005 0 ;
  ROWCOL 1 1 ;
END M2_M1_1


END LIBRARY
