MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 14.72 BY 18.984 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.984 18.528 6.016 18.6 ;
      LAYER M2 ;
        RECT 5.964 18.548 6.036 18.58 ;
      LAYER M1 ;
        RECT 8.864 18.528 8.896 18.6 ;
      LAYER M2 ;
        RECT 8.844 18.548 8.916 18.58 ;
      LAYER M2 ;
        RECT 6 18.548 8.88 18.58 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
      LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
      LAYER M1 ;
        RECT 8.704 0.384 8.736 0.456 ;
      LAYER M2 ;
        RECT 8.684 0.404 8.756 0.436 ;
      LAYER M2 ;
        RECT 5.84 0.404 8.72 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 18.696 3.136 18.768 ;
      LAYER M2 ;
        RECT 3.084 18.716 3.156 18.748 ;
      LAYER M1 ;
        RECT 11.744 18.696 11.776 18.768 ;
      LAYER M2 ;
        RECT 11.724 18.716 11.796 18.748 ;
      LAYER M2 ;
        RECT 3.12 18.716 11.76 18.748 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
      LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
      LAYER M1 ;
        RECT 11.584 0.216 11.616 0.288 ;
      LAYER M2 ;
        RECT 11.564 0.236 11.636 0.268 ;
      LAYER M2 ;
        RECT 2.96 0.236 11.6 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.144 6.768 6.176 6.84 ;
  LAYER M2 ;
        RECT 6.124 6.788 6.196 6.82 ;
  LAYER M2 ;
        RECT 5.84 6.788 6.16 6.82 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 6.84 ;
  LAYER M2 ;
        RECT 5.804 6.788 5.876 6.82 ;
  LAYER M1 ;
        RECT 6.144 9.708 6.176 9.78 ;
  LAYER M2 ;
        RECT 6.124 9.728 6.196 9.76 ;
  LAYER M2 ;
        RECT 5.84 9.728 6.16 9.76 ;
  LAYER M1 ;
        RECT 5.824 9.708 5.856 9.78 ;
  LAYER M2 ;
        RECT 5.804 9.728 5.876 9.76 ;
  LAYER M1 ;
        RECT 3.264 6.768 3.296 6.84 ;
  LAYER M2 ;
        RECT 3.244 6.788 3.316 6.82 ;
  LAYER M1 ;
        RECT 3.264 6.636 3.296 6.804 ;
  LAYER M1 ;
        RECT 3.264 6.6 3.296 6.672 ;
  LAYER M2 ;
        RECT 3.244 6.62 3.316 6.652 ;
  LAYER M2 ;
        RECT 3.28 6.62 5.84 6.652 ;
  LAYER M1 ;
        RECT 5.824 6.6 5.856 6.672 ;
  LAYER M2 ;
        RECT 5.804 6.62 5.876 6.652 ;
  LAYER M1 ;
        RECT 3.264 9.708 3.296 9.78 ;
  LAYER M2 ;
        RECT 3.244 9.728 3.316 9.76 ;
  LAYER M1 ;
        RECT 3.264 9.576 3.296 9.744 ;
  LAYER M1 ;
        RECT 3.264 9.54 3.296 9.612 ;
  LAYER M2 ;
        RECT 3.244 9.56 3.316 9.592 ;
  LAYER M2 ;
        RECT 3.28 9.56 5.84 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
  LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 0.588 ;
  LAYER M1 ;
        RECT 5.824 0.588 5.856 9.744 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 9.78 ;
  LAYER M2 ;
        RECT 9.004 9.728 9.076 9.76 ;
  LAYER M2 ;
        RECT 8.72 9.728 9.04 9.76 ;
  LAYER M1 ;
        RECT 8.704 9.708 8.736 9.78 ;
  LAYER M2 ;
        RECT 8.684 9.728 8.756 9.76 ;
  LAYER M1 ;
        RECT 9.024 6.768 9.056 6.84 ;
  LAYER M2 ;
        RECT 9.004 6.788 9.076 6.82 ;
  LAYER M2 ;
        RECT 8.72 6.788 9.04 6.82 ;
  LAYER M1 ;
        RECT 8.704 6.768 8.736 6.84 ;
  LAYER M2 ;
        RECT 8.684 6.788 8.756 6.82 ;
  LAYER M1 ;
        RECT 8.704 0.384 8.736 0.456 ;
  LAYER M2 ;
        RECT 8.684 0.404 8.756 0.436 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 0.588 ;
  LAYER M1 ;
        RECT 8.704 0.588 8.736 9.744 ;
  LAYER M2 ;
        RECT 5.84 0.404 8.72 0.436 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 12.72 ;
  LAYER M2 ;
        RECT 3.244 12.668 3.316 12.7 ;
  LAYER M2 ;
        RECT 2.96 12.668 3.28 12.7 ;
  LAYER M1 ;
        RECT 2.944 12.648 2.976 12.72 ;
  LAYER M2 ;
        RECT 2.924 12.668 2.996 12.7 ;
  LAYER M1 ;
        RECT 3.264 3.828 3.296 3.9 ;
  LAYER M2 ;
        RECT 3.244 3.848 3.316 3.88 ;
  LAYER M2 ;
        RECT 2.96 3.848 3.28 3.88 ;
  LAYER M1 ;
        RECT 2.944 3.828 2.976 3.9 ;
  LAYER M2 ;
        RECT 2.924 3.848 2.996 3.88 ;
  LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
  LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
  LAYER M1 ;
        RECT 2.944 0.252 2.976 0.588 ;
  LAYER M1 ;
        RECT 2.944 0.588 2.976 12.684 ;
  LAYER M1 ;
        RECT 9.024 3.828 9.056 3.9 ;
  LAYER M2 ;
        RECT 9.004 3.848 9.076 3.88 ;
  LAYER M1 ;
        RECT 9.024 3.696 9.056 3.864 ;
  LAYER M1 ;
        RECT 9.024 3.66 9.056 3.732 ;
  LAYER M2 ;
        RECT 9.004 3.68 9.076 3.712 ;
  LAYER M2 ;
        RECT 9.04 3.68 11.6 3.712 ;
  LAYER M1 ;
        RECT 11.584 3.66 11.616 3.732 ;
  LAYER M2 ;
        RECT 11.564 3.68 11.636 3.712 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 12.72 ;
  LAYER M2 ;
        RECT 9.004 12.668 9.076 12.7 ;
  LAYER M1 ;
        RECT 9.024 12.516 9.056 12.684 ;
  LAYER M1 ;
        RECT 9.024 12.48 9.056 12.552 ;
  LAYER M2 ;
        RECT 9.004 12.5 9.076 12.532 ;
  LAYER M2 ;
        RECT 9.04 12.5 11.6 12.532 ;
  LAYER M1 ;
        RECT 11.584 12.48 11.616 12.552 ;
  LAYER M2 ;
        RECT 11.564 12.5 11.636 12.532 ;
  LAYER M1 ;
        RECT 11.584 0.216 11.616 0.288 ;
  LAYER M2 ;
        RECT 11.564 0.236 11.636 0.268 ;
  LAYER M1 ;
        RECT 11.584 0.252 11.616 0.588 ;
  LAYER M1 ;
        RECT 11.584 0.588 11.616 12.516 ;
  LAYER M2 ;
        RECT 2.96 0.236 11.6 0.268 ;
  LAYER M1 ;
        RECT 6.144 3.828 6.176 3.9 ;
  LAYER M2 ;
        RECT 6.124 3.848 6.196 3.88 ;
  LAYER M2 ;
        RECT 6.16 3.848 9.04 3.88 ;
  LAYER M1 ;
        RECT 9.024 3.828 9.056 3.9 ;
  LAYER M2 ;
        RECT 9.004 3.848 9.076 3.88 ;
  LAYER M1 ;
        RECT 6.144 12.648 6.176 12.72 ;
  LAYER M2 ;
        RECT 6.124 12.668 6.196 12.7 ;
  LAYER M2 ;
        RECT 3.28 12.668 6.16 12.7 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 12.72 ;
  LAYER M2 ;
        RECT 3.244 12.668 3.316 12.7 ;
  LAYER M1 ;
        RECT 0.384 0.888 0.416 0.96 ;
  LAYER M2 ;
        RECT 0.364 0.908 0.436 0.94 ;
  LAYER M2 ;
        RECT 0.08 0.908 0.4 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 0.384 3.828 0.416 3.9 ;
  LAYER M2 ;
        RECT 0.364 3.848 0.436 3.88 ;
  LAYER M2 ;
        RECT 0.08 3.848 0.4 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 0.384 6.768 0.416 6.84 ;
  LAYER M2 ;
        RECT 0.364 6.788 0.436 6.82 ;
  LAYER M2 ;
        RECT 0.08 6.788 0.4 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 0.384 9.708 0.416 9.78 ;
  LAYER M2 ;
        RECT 0.364 9.728 0.436 9.76 ;
  LAYER M2 ;
        RECT 0.08 9.728 0.4 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 0.384 12.648 0.416 12.72 ;
  LAYER M2 ;
        RECT 0.364 12.668 0.436 12.7 ;
  LAYER M2 ;
        RECT 0.08 12.668 0.4 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 0.384 15.588 0.416 15.66 ;
  LAYER M2 ;
        RECT 0.364 15.608 0.436 15.64 ;
  LAYER M2 ;
        RECT 0.08 15.608 0.4 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.588 ;
  LAYER M1 ;
        RECT 0.064 0.588 0.096 15.624 ;
  LAYER M1 ;
        RECT 11.904 0.888 11.936 0.96 ;
  LAYER M2 ;
        RECT 11.884 0.908 11.956 0.94 ;
  LAYER M1 ;
        RECT 11.904 0.756 11.936 0.924 ;
  LAYER M1 ;
        RECT 11.904 0.72 11.936 0.792 ;
  LAYER M2 ;
        RECT 11.884 0.74 11.956 0.772 ;
  LAYER M2 ;
        RECT 11.92 0.74 14.48 0.772 ;
  LAYER M1 ;
        RECT 14.464 0.72 14.496 0.792 ;
  LAYER M2 ;
        RECT 14.444 0.74 14.516 0.772 ;
  LAYER M1 ;
        RECT 11.904 3.828 11.936 3.9 ;
  LAYER M2 ;
        RECT 11.884 3.848 11.956 3.88 ;
  LAYER M1 ;
        RECT 11.904 3.696 11.936 3.864 ;
  LAYER M1 ;
        RECT 11.904 3.66 11.936 3.732 ;
  LAYER M2 ;
        RECT 11.884 3.68 11.956 3.712 ;
  LAYER M2 ;
        RECT 11.92 3.68 14.48 3.712 ;
  LAYER M1 ;
        RECT 14.464 3.66 14.496 3.732 ;
  LAYER M2 ;
        RECT 14.444 3.68 14.516 3.712 ;
  LAYER M1 ;
        RECT 11.904 6.768 11.936 6.84 ;
  LAYER M2 ;
        RECT 11.884 6.788 11.956 6.82 ;
  LAYER M1 ;
        RECT 11.904 6.636 11.936 6.804 ;
  LAYER M1 ;
        RECT 11.904 6.6 11.936 6.672 ;
  LAYER M2 ;
        RECT 11.884 6.62 11.956 6.652 ;
  LAYER M2 ;
        RECT 11.92 6.62 14.48 6.652 ;
  LAYER M1 ;
        RECT 14.464 6.6 14.496 6.672 ;
  LAYER M2 ;
        RECT 14.444 6.62 14.516 6.652 ;
  LAYER M1 ;
        RECT 11.904 9.708 11.936 9.78 ;
  LAYER M2 ;
        RECT 11.884 9.728 11.956 9.76 ;
  LAYER M1 ;
        RECT 11.904 9.576 11.936 9.744 ;
  LAYER M1 ;
        RECT 11.904 9.54 11.936 9.612 ;
  LAYER M2 ;
        RECT 11.884 9.56 11.956 9.592 ;
  LAYER M2 ;
        RECT 11.92 9.56 14.48 9.592 ;
  LAYER M1 ;
        RECT 14.464 9.54 14.496 9.612 ;
  LAYER M2 ;
        RECT 14.444 9.56 14.516 9.592 ;
  LAYER M1 ;
        RECT 11.904 12.648 11.936 12.72 ;
  LAYER M2 ;
        RECT 11.884 12.668 11.956 12.7 ;
  LAYER M1 ;
        RECT 11.904 12.516 11.936 12.684 ;
  LAYER M1 ;
        RECT 11.904 12.48 11.936 12.552 ;
  LAYER M2 ;
        RECT 11.884 12.5 11.956 12.532 ;
  LAYER M2 ;
        RECT 11.92 12.5 14.48 12.532 ;
  LAYER M1 ;
        RECT 14.464 12.48 14.496 12.552 ;
  LAYER M2 ;
        RECT 14.444 12.5 14.516 12.532 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 15.66 ;
  LAYER M2 ;
        RECT 11.884 15.608 11.956 15.64 ;
  LAYER M1 ;
        RECT 11.904 15.456 11.936 15.624 ;
  LAYER M1 ;
        RECT 11.904 15.42 11.936 15.492 ;
  LAYER M2 ;
        RECT 11.884 15.44 11.956 15.472 ;
  LAYER M2 ;
        RECT 11.92 15.44 14.48 15.472 ;
  LAYER M1 ;
        RECT 14.464 15.42 14.496 15.492 ;
  LAYER M2 ;
        RECT 14.444 15.44 14.516 15.472 ;
  LAYER M1 ;
        RECT 14.464 0.048 14.496 0.12 ;
  LAYER M2 ;
        RECT 14.444 0.068 14.516 0.1 ;
  LAYER M1 ;
        RECT 14.464 0.084 14.496 0.588 ;
  LAYER M1 ;
        RECT 14.464 0.588 14.496 15.456 ;
  LAYER M2 ;
        RECT 0.08 0.068 14.48 0.1 ;
  LAYER M1 ;
        RECT 3.264 0.888 3.296 0.96 ;
  LAYER M2 ;
        RECT 3.244 0.908 3.316 0.94 ;
  LAYER M2 ;
        RECT 0.4 0.908 3.28 0.94 ;
  LAYER M1 ;
        RECT 0.384 0.888 0.416 0.96 ;
  LAYER M2 ;
        RECT 0.364 0.908 0.436 0.94 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M2 ;
        RECT 0.4 15.608 3.28 15.64 ;
  LAYER M1 ;
        RECT 0.384 15.588 0.416 15.66 ;
  LAYER M2 ;
        RECT 0.364 15.608 0.436 15.64 ;
  LAYER M1 ;
        RECT 6.144 15.588 6.176 15.66 ;
  LAYER M2 ;
        RECT 6.124 15.608 6.196 15.64 ;
  LAYER M2 ;
        RECT 3.28 15.608 6.16 15.64 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 15.66 ;
  LAYER M2 ;
        RECT 3.244 15.608 3.316 15.64 ;
  LAYER M1 ;
        RECT 9.024 15.588 9.056 15.66 ;
  LAYER M2 ;
        RECT 9.004 15.608 9.076 15.64 ;
  LAYER M2 ;
        RECT 6.16 15.608 9.04 15.64 ;
  LAYER M1 ;
        RECT 6.144 15.588 6.176 15.66 ;
  LAYER M2 ;
        RECT 6.124 15.608 6.196 15.64 ;
  LAYER M1 ;
        RECT 9.024 0.888 9.056 0.96 ;
  LAYER M2 ;
        RECT 9.004 0.908 9.076 0.94 ;
  LAYER M2 ;
        RECT 9.04 0.908 11.92 0.94 ;
  LAYER M1 ;
        RECT 11.904 0.888 11.936 0.96 ;
  LAYER M2 ;
        RECT 11.884 0.908 11.956 0.94 ;
  LAYER M1 ;
        RECT 6.144 0.888 6.176 0.96 ;
  LAYER M2 ;
        RECT 6.124 0.908 6.196 0.94 ;
  LAYER M2 ;
        RECT 6.16 0.908 9.04 0.94 ;
  LAYER M1 ;
        RECT 9.024 0.888 9.056 0.96 ;
  LAYER M2 ;
        RECT 9.004 0.908 9.076 0.94 ;
  LAYER M1 ;
        RECT 8.544 9.204 8.576 9.276 ;
  LAYER M2 ;
        RECT 8.524 9.224 8.596 9.256 ;
  LAYER M2 ;
        RECT 6 9.224 8.56 9.256 ;
  LAYER M1 ;
        RECT 5.984 9.204 6.016 9.276 ;
  LAYER M2 ;
        RECT 5.964 9.224 6.036 9.256 ;
  LAYER M1 ;
        RECT 8.544 12.144 8.576 12.216 ;
  LAYER M2 ;
        RECT 8.524 12.164 8.596 12.196 ;
  LAYER M2 ;
        RECT 6 12.164 8.56 12.196 ;
  LAYER M1 ;
        RECT 5.984 12.144 6.016 12.216 ;
  LAYER M2 ;
        RECT 5.964 12.164 6.036 12.196 ;
  LAYER M1 ;
        RECT 5.664 9.204 5.696 9.276 ;
  LAYER M2 ;
        RECT 5.644 9.224 5.716 9.256 ;
  LAYER M1 ;
        RECT 5.664 9.24 5.696 9.408 ;
  LAYER M1 ;
        RECT 5.664 9.372 5.696 9.444 ;
  LAYER M2 ;
        RECT 5.644 9.392 5.716 9.424 ;
  LAYER M2 ;
        RECT 5.68 9.392 6 9.424 ;
  LAYER M1 ;
        RECT 5.984 9.372 6.016 9.444 ;
  LAYER M2 ;
        RECT 5.964 9.392 6.036 9.424 ;
  LAYER M1 ;
        RECT 5.664 12.144 5.696 12.216 ;
  LAYER M2 ;
        RECT 5.644 12.164 5.716 12.196 ;
  LAYER M1 ;
        RECT 5.664 12.18 5.696 12.348 ;
  LAYER M1 ;
        RECT 5.664 12.312 5.696 12.384 ;
  LAYER M2 ;
        RECT 5.644 12.332 5.716 12.364 ;
  LAYER M2 ;
        RECT 5.68 12.332 6 12.364 ;
  LAYER M1 ;
        RECT 5.984 12.312 6.016 12.384 ;
  LAYER M2 ;
        RECT 5.964 12.332 6.036 12.364 ;
  LAYER M1 ;
        RECT 5.984 18.528 6.016 18.6 ;
  LAYER M2 ;
        RECT 5.964 18.548 6.036 18.58 ;
  LAYER M1 ;
        RECT 5.984 18.396 6.016 18.564 ;
  LAYER M1 ;
        RECT 5.984 9.24 6.016 18.396 ;
  LAYER M1 ;
        RECT 11.424 12.144 11.456 12.216 ;
  LAYER M2 ;
        RECT 11.404 12.164 11.476 12.196 ;
  LAYER M2 ;
        RECT 8.88 12.164 11.44 12.196 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M1 ;
        RECT 11.424 9.204 11.456 9.276 ;
  LAYER M2 ;
        RECT 11.404 9.224 11.476 9.256 ;
  LAYER M2 ;
        RECT 8.88 9.224 11.44 9.256 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M1 ;
        RECT 8.864 18.528 8.896 18.6 ;
  LAYER M2 ;
        RECT 8.844 18.548 8.916 18.58 ;
  LAYER M1 ;
        RECT 8.864 18.396 8.896 18.564 ;
  LAYER M1 ;
        RECT 8.864 9.24 8.896 18.396 ;
  LAYER M2 ;
        RECT 6 18.548 8.88 18.58 ;
  LAYER M1 ;
        RECT 5.664 15.084 5.696 15.156 ;
  LAYER M2 ;
        RECT 5.644 15.104 5.716 15.136 ;
  LAYER M2 ;
        RECT 3.12 15.104 5.68 15.136 ;
  LAYER M1 ;
        RECT 3.104 15.084 3.136 15.156 ;
  LAYER M2 ;
        RECT 3.084 15.104 3.156 15.136 ;
  LAYER M1 ;
        RECT 5.664 6.264 5.696 6.336 ;
  LAYER M2 ;
        RECT 5.644 6.284 5.716 6.316 ;
  LAYER M2 ;
        RECT 3.12 6.284 5.68 6.316 ;
  LAYER M1 ;
        RECT 3.104 6.264 3.136 6.336 ;
  LAYER M2 ;
        RECT 3.084 6.284 3.156 6.316 ;
  LAYER M1 ;
        RECT 3.104 18.696 3.136 18.768 ;
  LAYER M2 ;
        RECT 3.084 18.716 3.156 18.748 ;
  LAYER M1 ;
        RECT 3.104 18.396 3.136 18.732 ;
  LAYER M1 ;
        RECT 3.104 6.3 3.136 18.396 ;
  LAYER M1 ;
        RECT 11.424 6.264 11.456 6.336 ;
  LAYER M2 ;
        RECT 11.404 6.284 11.476 6.316 ;
  LAYER M1 ;
        RECT 11.424 6.3 11.456 6.468 ;
  LAYER M1 ;
        RECT 11.424 6.432 11.456 6.504 ;
  LAYER M2 ;
        RECT 11.404 6.452 11.476 6.484 ;
  LAYER M2 ;
        RECT 11.44 6.452 11.76 6.484 ;
  LAYER M1 ;
        RECT 11.744 6.432 11.776 6.504 ;
  LAYER M2 ;
        RECT 11.724 6.452 11.796 6.484 ;
  LAYER M1 ;
        RECT 11.424 15.084 11.456 15.156 ;
  LAYER M2 ;
        RECT 11.404 15.104 11.476 15.136 ;
  LAYER M1 ;
        RECT 11.424 15.12 11.456 15.288 ;
  LAYER M1 ;
        RECT 11.424 15.252 11.456 15.324 ;
  LAYER M2 ;
        RECT 11.404 15.272 11.476 15.304 ;
  LAYER M2 ;
        RECT 11.44 15.272 11.76 15.304 ;
  LAYER M1 ;
        RECT 11.744 15.252 11.776 15.324 ;
  LAYER M2 ;
        RECT 11.724 15.272 11.796 15.304 ;
  LAYER M1 ;
        RECT 11.744 18.696 11.776 18.768 ;
  LAYER M2 ;
        RECT 11.724 18.716 11.796 18.748 ;
  LAYER M1 ;
        RECT 11.744 18.396 11.776 18.732 ;
  LAYER M1 ;
        RECT 11.744 6.468 11.776 18.396 ;
  LAYER M2 ;
        RECT 3.12 18.716 11.76 18.748 ;
  LAYER M1 ;
        RECT 8.544 6.264 8.576 6.336 ;
  LAYER M2 ;
        RECT 8.524 6.284 8.596 6.316 ;
  LAYER M2 ;
        RECT 8.56 6.284 11.44 6.316 ;
  LAYER M1 ;
        RECT 11.424 6.264 11.456 6.336 ;
  LAYER M2 ;
        RECT 11.404 6.284 11.476 6.316 ;
  LAYER M1 ;
        RECT 8.544 15.084 8.576 15.156 ;
  LAYER M2 ;
        RECT 8.524 15.104 8.596 15.136 ;
  LAYER M2 ;
        RECT 5.68 15.104 8.56 15.136 ;
  LAYER M1 ;
        RECT 5.664 15.084 5.696 15.156 ;
  LAYER M2 ;
        RECT 5.644 15.104 5.716 15.136 ;
  LAYER M1 ;
        RECT 2.784 3.324 2.816 3.396 ;
  LAYER M2 ;
        RECT 2.764 3.344 2.836 3.376 ;
  LAYER M2 ;
        RECT 0.24 3.344 2.8 3.376 ;
  LAYER M1 ;
        RECT 0.224 3.324 0.256 3.396 ;
  LAYER M2 ;
        RECT 0.204 3.344 0.276 3.376 ;
  LAYER M1 ;
        RECT 2.784 6.264 2.816 6.336 ;
  LAYER M2 ;
        RECT 2.764 6.284 2.836 6.316 ;
  LAYER M2 ;
        RECT 0.24 6.284 2.8 6.316 ;
  LAYER M1 ;
        RECT 0.224 6.264 0.256 6.336 ;
  LAYER M2 ;
        RECT 0.204 6.284 0.276 6.316 ;
  LAYER M1 ;
        RECT 2.784 9.204 2.816 9.276 ;
  LAYER M2 ;
        RECT 2.764 9.224 2.836 9.256 ;
  LAYER M2 ;
        RECT 0.24 9.224 2.8 9.256 ;
  LAYER M1 ;
        RECT 0.224 9.204 0.256 9.276 ;
  LAYER M2 ;
        RECT 0.204 9.224 0.276 9.256 ;
  LAYER M1 ;
        RECT 2.784 12.144 2.816 12.216 ;
  LAYER M2 ;
        RECT 2.764 12.164 2.836 12.196 ;
  LAYER M2 ;
        RECT 0.24 12.164 2.8 12.196 ;
  LAYER M1 ;
        RECT 0.224 12.144 0.256 12.216 ;
  LAYER M2 ;
        RECT 0.204 12.164 0.276 12.196 ;
  LAYER M1 ;
        RECT 2.784 15.084 2.816 15.156 ;
  LAYER M2 ;
        RECT 2.764 15.104 2.836 15.136 ;
  LAYER M2 ;
        RECT 0.24 15.104 2.8 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.084 0.256 15.156 ;
  LAYER M2 ;
        RECT 0.204 15.104 0.276 15.136 ;
  LAYER M1 ;
        RECT 2.784 18.024 2.816 18.096 ;
  LAYER M2 ;
        RECT 2.764 18.044 2.836 18.076 ;
  LAYER M2 ;
        RECT 0.24 18.044 2.8 18.076 ;
  LAYER M1 ;
        RECT 0.224 18.024 0.256 18.096 ;
  LAYER M2 ;
        RECT 0.204 18.044 0.276 18.076 ;
  LAYER M1 ;
        RECT 0.224 18.864 0.256 18.936 ;
  LAYER M2 ;
        RECT 0.204 18.884 0.276 18.916 ;
  LAYER M1 ;
        RECT 0.224 18.396 0.256 18.9 ;
  LAYER M1 ;
        RECT 0.224 3.36 0.256 18.396 ;
  LAYER M1 ;
        RECT 14.304 3.324 14.336 3.396 ;
  LAYER M2 ;
        RECT 14.284 3.344 14.356 3.376 ;
  LAYER M1 ;
        RECT 14.304 3.36 14.336 3.528 ;
  LAYER M1 ;
        RECT 14.304 3.492 14.336 3.564 ;
  LAYER M2 ;
        RECT 14.284 3.512 14.356 3.544 ;
  LAYER M2 ;
        RECT 14.32 3.512 14.64 3.544 ;
  LAYER M1 ;
        RECT 14.624 3.492 14.656 3.564 ;
  LAYER M2 ;
        RECT 14.604 3.512 14.676 3.544 ;
  LAYER M1 ;
        RECT 14.304 6.264 14.336 6.336 ;
  LAYER M2 ;
        RECT 14.284 6.284 14.356 6.316 ;
  LAYER M1 ;
        RECT 14.304 6.3 14.336 6.468 ;
  LAYER M1 ;
        RECT 14.304 6.432 14.336 6.504 ;
  LAYER M2 ;
        RECT 14.284 6.452 14.356 6.484 ;
  LAYER M2 ;
        RECT 14.32 6.452 14.64 6.484 ;
  LAYER M1 ;
        RECT 14.624 6.432 14.656 6.504 ;
  LAYER M2 ;
        RECT 14.604 6.452 14.676 6.484 ;
  LAYER M1 ;
        RECT 14.304 9.204 14.336 9.276 ;
  LAYER M2 ;
        RECT 14.284 9.224 14.356 9.256 ;
  LAYER M1 ;
        RECT 14.304 9.24 14.336 9.408 ;
  LAYER M1 ;
        RECT 14.304 9.372 14.336 9.444 ;
  LAYER M2 ;
        RECT 14.284 9.392 14.356 9.424 ;
  LAYER M2 ;
        RECT 14.32 9.392 14.64 9.424 ;
  LAYER M1 ;
        RECT 14.624 9.372 14.656 9.444 ;
  LAYER M2 ;
        RECT 14.604 9.392 14.676 9.424 ;
  LAYER M1 ;
        RECT 14.304 12.144 14.336 12.216 ;
  LAYER M2 ;
        RECT 14.284 12.164 14.356 12.196 ;
  LAYER M1 ;
        RECT 14.304 12.18 14.336 12.348 ;
  LAYER M1 ;
        RECT 14.304 12.312 14.336 12.384 ;
  LAYER M2 ;
        RECT 14.284 12.332 14.356 12.364 ;
  LAYER M2 ;
        RECT 14.32 12.332 14.64 12.364 ;
  LAYER M1 ;
        RECT 14.624 12.312 14.656 12.384 ;
  LAYER M2 ;
        RECT 14.604 12.332 14.676 12.364 ;
  LAYER M1 ;
        RECT 14.304 15.084 14.336 15.156 ;
  LAYER M2 ;
        RECT 14.284 15.104 14.356 15.136 ;
  LAYER M1 ;
        RECT 14.304 15.12 14.336 15.288 ;
  LAYER M1 ;
        RECT 14.304 15.252 14.336 15.324 ;
  LAYER M2 ;
        RECT 14.284 15.272 14.356 15.304 ;
  LAYER M2 ;
        RECT 14.32 15.272 14.64 15.304 ;
  LAYER M1 ;
        RECT 14.624 15.252 14.656 15.324 ;
  LAYER M2 ;
        RECT 14.604 15.272 14.676 15.304 ;
  LAYER M1 ;
        RECT 14.304 18.024 14.336 18.096 ;
  LAYER M2 ;
        RECT 14.284 18.044 14.356 18.076 ;
  LAYER M1 ;
        RECT 14.304 18.06 14.336 18.228 ;
  LAYER M1 ;
        RECT 14.304 18.192 14.336 18.264 ;
  LAYER M2 ;
        RECT 14.284 18.212 14.356 18.244 ;
  LAYER M2 ;
        RECT 14.32 18.212 14.64 18.244 ;
  LAYER M1 ;
        RECT 14.624 18.192 14.656 18.264 ;
  LAYER M2 ;
        RECT 14.604 18.212 14.676 18.244 ;
  LAYER M1 ;
        RECT 14.624 18.864 14.656 18.936 ;
  LAYER M2 ;
        RECT 14.604 18.884 14.676 18.916 ;
  LAYER M1 ;
        RECT 14.624 18.396 14.656 18.9 ;
  LAYER M1 ;
        RECT 14.624 3.528 14.656 18.396 ;
  LAYER M2 ;
        RECT 0.24 18.884 14.64 18.916 ;
  LAYER M1 ;
        RECT 5.664 3.324 5.696 3.396 ;
  LAYER M2 ;
        RECT 5.644 3.344 5.716 3.376 ;
  LAYER M2 ;
        RECT 2.8 3.344 5.68 3.376 ;
  LAYER M1 ;
        RECT 2.784 3.324 2.816 3.396 ;
  LAYER M2 ;
        RECT 2.764 3.344 2.836 3.376 ;
  LAYER M1 ;
        RECT 5.664 18.024 5.696 18.096 ;
  LAYER M2 ;
        RECT 5.644 18.044 5.716 18.076 ;
  LAYER M2 ;
        RECT 2.8 18.044 5.68 18.076 ;
  LAYER M1 ;
        RECT 2.784 18.024 2.816 18.096 ;
  LAYER M2 ;
        RECT 2.764 18.044 2.836 18.076 ;
  LAYER M1 ;
        RECT 8.544 18.024 8.576 18.096 ;
  LAYER M2 ;
        RECT 8.524 18.044 8.596 18.076 ;
  LAYER M2 ;
        RECT 5.68 18.044 8.56 18.076 ;
  LAYER M1 ;
        RECT 5.664 18.024 5.696 18.096 ;
  LAYER M2 ;
        RECT 5.644 18.044 5.716 18.076 ;
  LAYER M1 ;
        RECT 11.424 18.024 11.456 18.096 ;
  LAYER M2 ;
        RECT 11.404 18.044 11.476 18.076 ;
  LAYER M2 ;
        RECT 8.56 18.044 11.44 18.076 ;
  LAYER M1 ;
        RECT 8.544 18.024 8.576 18.096 ;
  LAYER M2 ;
        RECT 8.524 18.044 8.596 18.076 ;
  LAYER M1 ;
        RECT 11.424 3.324 11.456 3.396 ;
  LAYER M2 ;
        RECT 11.404 3.344 11.476 3.376 ;
  LAYER M2 ;
        RECT 11.44 3.344 14.32 3.376 ;
  LAYER M1 ;
        RECT 14.304 3.324 14.336 3.396 ;
  LAYER M2 ;
        RECT 14.284 3.344 14.356 3.376 ;
  LAYER M1 ;
        RECT 8.544 3.324 8.576 3.396 ;
  LAYER M2 ;
        RECT 8.524 3.344 8.596 3.376 ;
  LAYER M2 ;
        RECT 8.56 3.344 11.44 3.376 ;
  LAYER M1 ;
        RECT 11.424 3.324 11.456 3.396 ;
  LAYER M2 ;
        RECT 11.404 3.344 11.476 3.376 ;
  LAYER M1 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M1 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M1 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M1 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M1 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M1 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M1 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M1 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M1 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M1 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M1 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M1 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M1 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M1 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M1 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M1 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M1 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M1 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M1 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M1 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M1 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M1 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M1 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M1 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M1 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M1 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M1 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M1 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M1 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M1 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M1 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M1 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M1 ;
        RECT 2.432 0.888 2.464 3.396 ;
  LAYER M1 ;
        RECT 2.496 0.888 2.528 3.396 ;
  LAYER M1 ;
        RECT 2.56 0.888 2.592 3.396 ;
  LAYER M1 ;
        RECT 2.624 0.888 2.656 3.396 ;
  LAYER M1 ;
        RECT 2.688 0.888 2.72 3.396 ;
  LAYER M2 ;
        RECT 0.364 0.972 2.836 1.004 ;
  LAYER M2 ;
        RECT 0.364 1.036 2.836 1.068 ;
  LAYER M2 ;
        RECT 0.364 1.1 2.836 1.132 ;
  LAYER M2 ;
        RECT 0.364 1.164 2.836 1.196 ;
  LAYER M2 ;
        RECT 0.364 1.228 2.836 1.26 ;
  LAYER M2 ;
        RECT 0.364 1.292 2.836 1.324 ;
  LAYER M2 ;
        RECT 0.364 1.356 2.836 1.388 ;
  LAYER M2 ;
        RECT 0.364 1.42 2.836 1.452 ;
  LAYER M2 ;
        RECT 0.364 1.484 2.836 1.516 ;
  LAYER M2 ;
        RECT 0.364 1.548 2.836 1.58 ;
  LAYER M2 ;
        RECT 0.364 1.612 2.836 1.644 ;
  LAYER M2 ;
        RECT 0.364 1.676 2.836 1.708 ;
  LAYER M2 ;
        RECT 0.364 1.74 2.836 1.772 ;
  LAYER M2 ;
        RECT 0.364 1.804 2.836 1.836 ;
  LAYER M2 ;
        RECT 0.364 1.868 2.836 1.9 ;
  LAYER M2 ;
        RECT 0.364 1.932 2.836 1.964 ;
  LAYER M2 ;
        RECT 0.364 1.996 2.836 2.028 ;
  LAYER M2 ;
        RECT 0.364 2.06 2.836 2.092 ;
  LAYER M2 ;
        RECT 0.364 2.124 2.836 2.156 ;
  LAYER M2 ;
        RECT 0.364 2.188 2.836 2.22 ;
  LAYER M2 ;
        RECT 0.364 2.252 2.836 2.284 ;
  LAYER M2 ;
        RECT 0.364 2.316 2.836 2.348 ;
  LAYER M2 ;
        RECT 0.364 2.38 2.836 2.412 ;
  LAYER M2 ;
        RECT 0.364 2.444 2.836 2.476 ;
  LAYER M2 ;
        RECT 0.364 2.508 2.836 2.54 ;
  LAYER M2 ;
        RECT 0.364 2.572 2.836 2.604 ;
  LAYER M2 ;
        RECT 0.364 2.636 2.836 2.668 ;
  LAYER M2 ;
        RECT 0.364 2.7 2.836 2.732 ;
  LAYER M2 ;
        RECT 0.364 2.764 2.836 2.796 ;
  LAYER M2 ;
        RECT 0.364 2.828 2.836 2.86 ;
  LAYER M2 ;
        RECT 0.364 2.892 2.836 2.924 ;
  LAYER M2 ;
        RECT 0.364 2.956 2.836 2.988 ;
  LAYER M2 ;
        RECT 0.364 3.02 2.836 3.052 ;
  LAYER M2 ;
        RECT 0.364 3.084 2.836 3.116 ;
  LAYER M2 ;
        RECT 0.364 3.148 2.836 3.18 ;
  LAYER M2 ;
        RECT 0.364 3.212 2.836 3.244 ;
  LAYER M3 ;
        RECT 0.384 0.888 0.416 3.396 ;
  LAYER M3 ;
        RECT 0.448 0.888 0.48 3.396 ;
  LAYER M3 ;
        RECT 0.512 0.888 0.544 3.396 ;
  LAYER M3 ;
        RECT 0.576 0.888 0.608 3.396 ;
  LAYER M3 ;
        RECT 0.64 0.888 0.672 3.396 ;
  LAYER M3 ;
        RECT 0.704 0.888 0.736 3.396 ;
  LAYER M3 ;
        RECT 0.768 0.888 0.8 3.396 ;
  LAYER M3 ;
        RECT 0.832 0.888 0.864 3.396 ;
  LAYER M3 ;
        RECT 0.896 0.888 0.928 3.396 ;
  LAYER M3 ;
        RECT 0.96 0.888 0.992 3.396 ;
  LAYER M3 ;
        RECT 1.024 0.888 1.056 3.396 ;
  LAYER M3 ;
        RECT 1.088 0.888 1.12 3.396 ;
  LAYER M3 ;
        RECT 1.152 0.888 1.184 3.396 ;
  LAYER M3 ;
        RECT 1.216 0.888 1.248 3.396 ;
  LAYER M3 ;
        RECT 1.28 0.888 1.312 3.396 ;
  LAYER M3 ;
        RECT 1.344 0.888 1.376 3.396 ;
  LAYER M3 ;
        RECT 1.408 0.888 1.44 3.396 ;
  LAYER M3 ;
        RECT 1.472 0.888 1.504 3.396 ;
  LAYER M3 ;
        RECT 1.536 0.888 1.568 3.396 ;
  LAYER M3 ;
        RECT 1.6 0.888 1.632 3.396 ;
  LAYER M3 ;
        RECT 1.664 0.888 1.696 3.396 ;
  LAYER M3 ;
        RECT 1.728 0.888 1.76 3.396 ;
  LAYER M3 ;
        RECT 1.792 0.888 1.824 3.396 ;
  LAYER M3 ;
        RECT 1.856 0.888 1.888 3.396 ;
  LAYER M3 ;
        RECT 1.92 0.888 1.952 3.396 ;
  LAYER M3 ;
        RECT 1.984 0.888 2.016 3.396 ;
  LAYER M3 ;
        RECT 2.048 0.888 2.08 3.396 ;
  LAYER M3 ;
        RECT 2.112 0.888 2.144 3.396 ;
  LAYER M3 ;
        RECT 2.176 0.888 2.208 3.396 ;
  LAYER M3 ;
        RECT 2.24 0.888 2.272 3.396 ;
  LAYER M3 ;
        RECT 2.304 0.888 2.336 3.396 ;
  LAYER M3 ;
        RECT 2.368 0.888 2.4 3.396 ;
  LAYER M3 ;
        RECT 2.432 0.888 2.464 3.396 ;
  LAYER M3 ;
        RECT 2.496 0.888 2.528 3.396 ;
  LAYER M3 ;
        RECT 2.56 0.888 2.592 3.396 ;
  LAYER M3 ;
        RECT 2.624 0.888 2.656 3.396 ;
  LAYER M3 ;
        RECT 2.688 0.888 2.72 3.396 ;
  LAYER M3 ;
        RECT 2.784 0.888 2.816 3.396 ;
  LAYER M1 ;
        RECT 0.399 0.924 0.401 3.36 ;
  LAYER M1 ;
        RECT 0.479 0.924 0.481 3.36 ;
  LAYER M1 ;
        RECT 0.559 0.924 0.561 3.36 ;
  LAYER M1 ;
        RECT 0.639 0.924 0.641 3.36 ;
  LAYER M1 ;
        RECT 0.719 0.924 0.721 3.36 ;
  LAYER M1 ;
        RECT 0.799 0.924 0.801 3.36 ;
  LAYER M1 ;
        RECT 0.879 0.924 0.881 3.36 ;
  LAYER M1 ;
        RECT 0.959 0.924 0.961 3.36 ;
  LAYER M1 ;
        RECT 1.039 0.924 1.041 3.36 ;
  LAYER M1 ;
        RECT 1.119 0.924 1.121 3.36 ;
  LAYER M1 ;
        RECT 1.199 0.924 1.201 3.36 ;
  LAYER M1 ;
        RECT 1.279 0.924 1.281 3.36 ;
  LAYER M1 ;
        RECT 1.359 0.924 1.361 3.36 ;
  LAYER M1 ;
        RECT 1.439 0.924 1.441 3.36 ;
  LAYER M1 ;
        RECT 1.519 0.924 1.521 3.36 ;
  LAYER M1 ;
        RECT 1.599 0.924 1.601 3.36 ;
  LAYER M1 ;
        RECT 1.679 0.924 1.681 3.36 ;
  LAYER M1 ;
        RECT 1.759 0.924 1.761 3.36 ;
  LAYER M1 ;
        RECT 1.839 0.924 1.841 3.36 ;
  LAYER M1 ;
        RECT 1.919 0.924 1.921 3.36 ;
  LAYER M1 ;
        RECT 1.999 0.924 2.001 3.36 ;
  LAYER M1 ;
        RECT 2.079 0.924 2.081 3.36 ;
  LAYER M1 ;
        RECT 2.159 0.924 2.161 3.36 ;
  LAYER M1 ;
        RECT 2.239 0.924 2.241 3.36 ;
  LAYER M1 ;
        RECT 2.319 0.924 2.321 3.36 ;
  LAYER M1 ;
        RECT 2.399 0.924 2.401 3.36 ;
  LAYER M1 ;
        RECT 2.479 0.924 2.481 3.36 ;
  LAYER M1 ;
        RECT 2.559 0.924 2.561 3.36 ;
  LAYER M1 ;
        RECT 2.639 0.924 2.641 3.36 ;
  LAYER M1 ;
        RECT 2.719 0.924 2.721 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.923 2.8 0.925 ;
  LAYER M2 ;
        RECT 0.4 1.007 2.8 1.009 ;
  LAYER M2 ;
        RECT 0.4 1.091 2.8 1.093 ;
  LAYER M2 ;
        RECT 0.4 1.175 2.8 1.177 ;
  LAYER M2 ;
        RECT 0.4 1.259 2.8 1.261 ;
  LAYER M2 ;
        RECT 0.4 1.343 2.8 1.345 ;
  LAYER M2 ;
        RECT 0.4 1.427 2.8 1.429 ;
  LAYER M2 ;
        RECT 0.4 1.511 2.8 1.513 ;
  LAYER M2 ;
        RECT 0.4 1.595 2.8 1.597 ;
  LAYER M2 ;
        RECT 0.4 1.679 2.8 1.681 ;
  LAYER M2 ;
        RECT 0.4 1.763 2.8 1.765 ;
  LAYER M2 ;
        RECT 0.4 1.847 2.8 1.849 ;
  LAYER M2 ;
        RECT 0.4 1.9305 2.8 1.9325 ;
  LAYER M2 ;
        RECT 0.4 2.015 2.8 2.017 ;
  LAYER M2 ;
        RECT 0.4 2.099 2.8 2.101 ;
  LAYER M2 ;
        RECT 0.4 2.183 2.8 2.185 ;
  LAYER M2 ;
        RECT 0.4 2.267 2.8 2.269 ;
  LAYER M2 ;
        RECT 0.4 2.351 2.8 2.353 ;
  LAYER M2 ;
        RECT 0.4 2.435 2.8 2.437 ;
  LAYER M2 ;
        RECT 0.4 2.519 2.8 2.521 ;
  LAYER M2 ;
        RECT 0.4 2.603 2.8 2.605 ;
  LAYER M2 ;
        RECT 0.4 2.687 2.8 2.689 ;
  LAYER M2 ;
        RECT 0.4 2.771 2.8 2.773 ;
  LAYER M2 ;
        RECT 0.4 2.855 2.8 2.857 ;
  LAYER M2 ;
        RECT 0.4 2.939 2.8 2.941 ;
  LAYER M2 ;
        RECT 0.4 3.023 2.8 3.025 ;
  LAYER M2 ;
        RECT 0.4 3.107 2.8 3.109 ;
  LAYER M2 ;
        RECT 0.4 3.191 2.8 3.193 ;
  LAYER M2 ;
        RECT 0.4 3.275 2.8 3.277 ;
  LAYER M1 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M1 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M1 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M1 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M1 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M1 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M1 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M1 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M1 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M1 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M1 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M1 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M1 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M1 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M1 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M1 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M1 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M1 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M1 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M1 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M1 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M1 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M1 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M1 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M1 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M1 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M1 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M1 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M1 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M1 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M1 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M1 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M1 ;
        RECT 2.432 3.828 2.464 6.336 ;
  LAYER M1 ;
        RECT 2.496 3.828 2.528 6.336 ;
  LAYER M1 ;
        RECT 2.56 3.828 2.592 6.336 ;
  LAYER M1 ;
        RECT 2.624 3.828 2.656 6.336 ;
  LAYER M1 ;
        RECT 2.688 3.828 2.72 6.336 ;
  LAYER M2 ;
        RECT 0.364 3.912 2.836 3.944 ;
  LAYER M2 ;
        RECT 0.364 3.976 2.836 4.008 ;
  LAYER M2 ;
        RECT 0.364 4.04 2.836 4.072 ;
  LAYER M2 ;
        RECT 0.364 4.104 2.836 4.136 ;
  LAYER M2 ;
        RECT 0.364 4.168 2.836 4.2 ;
  LAYER M2 ;
        RECT 0.364 4.232 2.836 4.264 ;
  LAYER M2 ;
        RECT 0.364 4.296 2.836 4.328 ;
  LAYER M2 ;
        RECT 0.364 4.36 2.836 4.392 ;
  LAYER M2 ;
        RECT 0.364 4.424 2.836 4.456 ;
  LAYER M2 ;
        RECT 0.364 4.488 2.836 4.52 ;
  LAYER M2 ;
        RECT 0.364 4.552 2.836 4.584 ;
  LAYER M2 ;
        RECT 0.364 4.616 2.836 4.648 ;
  LAYER M2 ;
        RECT 0.364 4.68 2.836 4.712 ;
  LAYER M2 ;
        RECT 0.364 4.744 2.836 4.776 ;
  LAYER M2 ;
        RECT 0.364 4.808 2.836 4.84 ;
  LAYER M2 ;
        RECT 0.364 4.872 2.836 4.904 ;
  LAYER M2 ;
        RECT 0.364 4.936 2.836 4.968 ;
  LAYER M2 ;
        RECT 0.364 5 2.836 5.032 ;
  LAYER M2 ;
        RECT 0.364 5.064 2.836 5.096 ;
  LAYER M2 ;
        RECT 0.364 5.128 2.836 5.16 ;
  LAYER M2 ;
        RECT 0.364 5.192 2.836 5.224 ;
  LAYER M2 ;
        RECT 0.364 5.256 2.836 5.288 ;
  LAYER M2 ;
        RECT 0.364 5.32 2.836 5.352 ;
  LAYER M2 ;
        RECT 0.364 5.384 2.836 5.416 ;
  LAYER M2 ;
        RECT 0.364 5.448 2.836 5.48 ;
  LAYER M2 ;
        RECT 0.364 5.512 2.836 5.544 ;
  LAYER M2 ;
        RECT 0.364 5.576 2.836 5.608 ;
  LAYER M2 ;
        RECT 0.364 5.64 2.836 5.672 ;
  LAYER M2 ;
        RECT 0.364 5.704 2.836 5.736 ;
  LAYER M2 ;
        RECT 0.364 5.768 2.836 5.8 ;
  LAYER M2 ;
        RECT 0.364 5.832 2.836 5.864 ;
  LAYER M2 ;
        RECT 0.364 5.896 2.836 5.928 ;
  LAYER M2 ;
        RECT 0.364 5.96 2.836 5.992 ;
  LAYER M2 ;
        RECT 0.364 6.024 2.836 6.056 ;
  LAYER M2 ;
        RECT 0.364 6.088 2.836 6.12 ;
  LAYER M2 ;
        RECT 0.364 6.152 2.836 6.184 ;
  LAYER M3 ;
        RECT 0.384 3.828 0.416 6.336 ;
  LAYER M3 ;
        RECT 0.448 3.828 0.48 6.336 ;
  LAYER M3 ;
        RECT 0.512 3.828 0.544 6.336 ;
  LAYER M3 ;
        RECT 0.576 3.828 0.608 6.336 ;
  LAYER M3 ;
        RECT 0.64 3.828 0.672 6.336 ;
  LAYER M3 ;
        RECT 0.704 3.828 0.736 6.336 ;
  LAYER M3 ;
        RECT 0.768 3.828 0.8 6.336 ;
  LAYER M3 ;
        RECT 0.832 3.828 0.864 6.336 ;
  LAYER M3 ;
        RECT 0.896 3.828 0.928 6.336 ;
  LAYER M3 ;
        RECT 0.96 3.828 0.992 6.336 ;
  LAYER M3 ;
        RECT 1.024 3.828 1.056 6.336 ;
  LAYER M3 ;
        RECT 1.088 3.828 1.12 6.336 ;
  LAYER M3 ;
        RECT 1.152 3.828 1.184 6.336 ;
  LAYER M3 ;
        RECT 1.216 3.828 1.248 6.336 ;
  LAYER M3 ;
        RECT 1.28 3.828 1.312 6.336 ;
  LAYER M3 ;
        RECT 1.344 3.828 1.376 6.336 ;
  LAYER M3 ;
        RECT 1.408 3.828 1.44 6.336 ;
  LAYER M3 ;
        RECT 1.472 3.828 1.504 6.336 ;
  LAYER M3 ;
        RECT 1.536 3.828 1.568 6.336 ;
  LAYER M3 ;
        RECT 1.6 3.828 1.632 6.336 ;
  LAYER M3 ;
        RECT 1.664 3.828 1.696 6.336 ;
  LAYER M3 ;
        RECT 1.728 3.828 1.76 6.336 ;
  LAYER M3 ;
        RECT 1.792 3.828 1.824 6.336 ;
  LAYER M3 ;
        RECT 1.856 3.828 1.888 6.336 ;
  LAYER M3 ;
        RECT 1.92 3.828 1.952 6.336 ;
  LAYER M3 ;
        RECT 1.984 3.828 2.016 6.336 ;
  LAYER M3 ;
        RECT 2.048 3.828 2.08 6.336 ;
  LAYER M3 ;
        RECT 2.112 3.828 2.144 6.336 ;
  LAYER M3 ;
        RECT 2.176 3.828 2.208 6.336 ;
  LAYER M3 ;
        RECT 2.24 3.828 2.272 6.336 ;
  LAYER M3 ;
        RECT 2.304 3.828 2.336 6.336 ;
  LAYER M3 ;
        RECT 2.368 3.828 2.4 6.336 ;
  LAYER M3 ;
        RECT 2.432 3.828 2.464 6.336 ;
  LAYER M3 ;
        RECT 2.496 3.828 2.528 6.336 ;
  LAYER M3 ;
        RECT 2.56 3.828 2.592 6.336 ;
  LAYER M3 ;
        RECT 2.624 3.828 2.656 6.336 ;
  LAYER M3 ;
        RECT 2.688 3.828 2.72 6.336 ;
  LAYER M3 ;
        RECT 2.784 3.828 2.816 6.336 ;
  LAYER M1 ;
        RECT 0.399 3.864 0.401 6.3 ;
  LAYER M1 ;
        RECT 0.479 3.864 0.481 6.3 ;
  LAYER M1 ;
        RECT 0.559 3.864 0.561 6.3 ;
  LAYER M1 ;
        RECT 0.639 3.864 0.641 6.3 ;
  LAYER M1 ;
        RECT 0.719 3.864 0.721 6.3 ;
  LAYER M1 ;
        RECT 0.799 3.864 0.801 6.3 ;
  LAYER M1 ;
        RECT 0.879 3.864 0.881 6.3 ;
  LAYER M1 ;
        RECT 0.959 3.864 0.961 6.3 ;
  LAYER M1 ;
        RECT 1.039 3.864 1.041 6.3 ;
  LAYER M1 ;
        RECT 1.119 3.864 1.121 6.3 ;
  LAYER M1 ;
        RECT 1.199 3.864 1.201 6.3 ;
  LAYER M1 ;
        RECT 1.279 3.864 1.281 6.3 ;
  LAYER M1 ;
        RECT 1.359 3.864 1.361 6.3 ;
  LAYER M1 ;
        RECT 1.439 3.864 1.441 6.3 ;
  LAYER M1 ;
        RECT 1.519 3.864 1.521 6.3 ;
  LAYER M1 ;
        RECT 1.599 3.864 1.601 6.3 ;
  LAYER M1 ;
        RECT 1.679 3.864 1.681 6.3 ;
  LAYER M1 ;
        RECT 1.759 3.864 1.761 6.3 ;
  LAYER M1 ;
        RECT 1.839 3.864 1.841 6.3 ;
  LAYER M1 ;
        RECT 1.919 3.864 1.921 6.3 ;
  LAYER M1 ;
        RECT 1.999 3.864 2.001 6.3 ;
  LAYER M1 ;
        RECT 2.079 3.864 2.081 6.3 ;
  LAYER M1 ;
        RECT 2.159 3.864 2.161 6.3 ;
  LAYER M1 ;
        RECT 2.239 3.864 2.241 6.3 ;
  LAYER M1 ;
        RECT 2.319 3.864 2.321 6.3 ;
  LAYER M1 ;
        RECT 2.399 3.864 2.401 6.3 ;
  LAYER M1 ;
        RECT 2.479 3.864 2.481 6.3 ;
  LAYER M1 ;
        RECT 2.559 3.864 2.561 6.3 ;
  LAYER M1 ;
        RECT 2.639 3.864 2.641 6.3 ;
  LAYER M1 ;
        RECT 2.719 3.864 2.721 6.3 ;
  LAYER M2 ;
        RECT 0.4 3.863 2.8 3.865 ;
  LAYER M2 ;
        RECT 0.4 3.947 2.8 3.949 ;
  LAYER M2 ;
        RECT 0.4 4.031 2.8 4.033 ;
  LAYER M2 ;
        RECT 0.4 4.115 2.8 4.117 ;
  LAYER M2 ;
        RECT 0.4 4.199 2.8 4.201 ;
  LAYER M2 ;
        RECT 0.4 4.283 2.8 4.285 ;
  LAYER M2 ;
        RECT 0.4 4.367 2.8 4.369 ;
  LAYER M2 ;
        RECT 0.4 4.451 2.8 4.453 ;
  LAYER M2 ;
        RECT 0.4 4.535 2.8 4.537 ;
  LAYER M2 ;
        RECT 0.4 4.619 2.8 4.621 ;
  LAYER M2 ;
        RECT 0.4 4.703 2.8 4.705 ;
  LAYER M2 ;
        RECT 0.4 4.787 2.8 4.789 ;
  LAYER M2 ;
        RECT 0.4 4.8705 2.8 4.8725 ;
  LAYER M2 ;
        RECT 0.4 4.955 2.8 4.957 ;
  LAYER M2 ;
        RECT 0.4 5.039 2.8 5.041 ;
  LAYER M2 ;
        RECT 0.4 5.123 2.8 5.125 ;
  LAYER M2 ;
        RECT 0.4 5.207 2.8 5.209 ;
  LAYER M2 ;
        RECT 0.4 5.291 2.8 5.293 ;
  LAYER M2 ;
        RECT 0.4 5.375 2.8 5.377 ;
  LAYER M2 ;
        RECT 0.4 5.459 2.8 5.461 ;
  LAYER M2 ;
        RECT 0.4 5.543 2.8 5.545 ;
  LAYER M2 ;
        RECT 0.4 5.627 2.8 5.629 ;
  LAYER M2 ;
        RECT 0.4 5.711 2.8 5.713 ;
  LAYER M2 ;
        RECT 0.4 5.795 2.8 5.797 ;
  LAYER M2 ;
        RECT 0.4 5.879 2.8 5.881 ;
  LAYER M2 ;
        RECT 0.4 5.963 2.8 5.965 ;
  LAYER M2 ;
        RECT 0.4 6.047 2.8 6.049 ;
  LAYER M2 ;
        RECT 0.4 6.131 2.8 6.133 ;
  LAYER M2 ;
        RECT 0.4 6.215 2.8 6.217 ;
  LAYER M1 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M1 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M1 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M1 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M1 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M1 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M1 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M1 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M1 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M1 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M1 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M1 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M1 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M1 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M1 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M1 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M1 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M1 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M1 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M1 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M1 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M1 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M1 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M1 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M1 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M1 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M1 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M1 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M1 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M1 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M1 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M1 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M1 ;
        RECT 2.432 6.768 2.464 9.276 ;
  LAYER M1 ;
        RECT 2.496 6.768 2.528 9.276 ;
  LAYER M1 ;
        RECT 2.56 6.768 2.592 9.276 ;
  LAYER M1 ;
        RECT 2.624 6.768 2.656 9.276 ;
  LAYER M1 ;
        RECT 2.688 6.768 2.72 9.276 ;
  LAYER M2 ;
        RECT 0.364 6.852 2.836 6.884 ;
  LAYER M2 ;
        RECT 0.364 6.916 2.836 6.948 ;
  LAYER M2 ;
        RECT 0.364 6.98 2.836 7.012 ;
  LAYER M2 ;
        RECT 0.364 7.044 2.836 7.076 ;
  LAYER M2 ;
        RECT 0.364 7.108 2.836 7.14 ;
  LAYER M2 ;
        RECT 0.364 7.172 2.836 7.204 ;
  LAYER M2 ;
        RECT 0.364 7.236 2.836 7.268 ;
  LAYER M2 ;
        RECT 0.364 7.3 2.836 7.332 ;
  LAYER M2 ;
        RECT 0.364 7.364 2.836 7.396 ;
  LAYER M2 ;
        RECT 0.364 7.428 2.836 7.46 ;
  LAYER M2 ;
        RECT 0.364 7.492 2.836 7.524 ;
  LAYER M2 ;
        RECT 0.364 7.556 2.836 7.588 ;
  LAYER M2 ;
        RECT 0.364 7.62 2.836 7.652 ;
  LAYER M2 ;
        RECT 0.364 7.684 2.836 7.716 ;
  LAYER M2 ;
        RECT 0.364 7.748 2.836 7.78 ;
  LAYER M2 ;
        RECT 0.364 7.812 2.836 7.844 ;
  LAYER M2 ;
        RECT 0.364 7.876 2.836 7.908 ;
  LAYER M2 ;
        RECT 0.364 7.94 2.836 7.972 ;
  LAYER M2 ;
        RECT 0.364 8.004 2.836 8.036 ;
  LAYER M2 ;
        RECT 0.364 8.068 2.836 8.1 ;
  LAYER M2 ;
        RECT 0.364 8.132 2.836 8.164 ;
  LAYER M2 ;
        RECT 0.364 8.196 2.836 8.228 ;
  LAYER M2 ;
        RECT 0.364 8.26 2.836 8.292 ;
  LAYER M2 ;
        RECT 0.364 8.324 2.836 8.356 ;
  LAYER M2 ;
        RECT 0.364 8.388 2.836 8.42 ;
  LAYER M2 ;
        RECT 0.364 8.452 2.836 8.484 ;
  LAYER M2 ;
        RECT 0.364 8.516 2.836 8.548 ;
  LAYER M2 ;
        RECT 0.364 8.58 2.836 8.612 ;
  LAYER M2 ;
        RECT 0.364 8.644 2.836 8.676 ;
  LAYER M2 ;
        RECT 0.364 8.708 2.836 8.74 ;
  LAYER M2 ;
        RECT 0.364 8.772 2.836 8.804 ;
  LAYER M2 ;
        RECT 0.364 8.836 2.836 8.868 ;
  LAYER M2 ;
        RECT 0.364 8.9 2.836 8.932 ;
  LAYER M2 ;
        RECT 0.364 8.964 2.836 8.996 ;
  LAYER M2 ;
        RECT 0.364 9.028 2.836 9.06 ;
  LAYER M2 ;
        RECT 0.364 9.092 2.836 9.124 ;
  LAYER M3 ;
        RECT 0.384 6.768 0.416 9.276 ;
  LAYER M3 ;
        RECT 0.448 6.768 0.48 9.276 ;
  LAYER M3 ;
        RECT 0.512 6.768 0.544 9.276 ;
  LAYER M3 ;
        RECT 0.576 6.768 0.608 9.276 ;
  LAYER M3 ;
        RECT 0.64 6.768 0.672 9.276 ;
  LAYER M3 ;
        RECT 0.704 6.768 0.736 9.276 ;
  LAYER M3 ;
        RECT 0.768 6.768 0.8 9.276 ;
  LAYER M3 ;
        RECT 0.832 6.768 0.864 9.276 ;
  LAYER M3 ;
        RECT 0.896 6.768 0.928 9.276 ;
  LAYER M3 ;
        RECT 0.96 6.768 0.992 9.276 ;
  LAYER M3 ;
        RECT 1.024 6.768 1.056 9.276 ;
  LAYER M3 ;
        RECT 1.088 6.768 1.12 9.276 ;
  LAYER M3 ;
        RECT 1.152 6.768 1.184 9.276 ;
  LAYER M3 ;
        RECT 1.216 6.768 1.248 9.276 ;
  LAYER M3 ;
        RECT 1.28 6.768 1.312 9.276 ;
  LAYER M3 ;
        RECT 1.344 6.768 1.376 9.276 ;
  LAYER M3 ;
        RECT 1.408 6.768 1.44 9.276 ;
  LAYER M3 ;
        RECT 1.472 6.768 1.504 9.276 ;
  LAYER M3 ;
        RECT 1.536 6.768 1.568 9.276 ;
  LAYER M3 ;
        RECT 1.6 6.768 1.632 9.276 ;
  LAYER M3 ;
        RECT 1.664 6.768 1.696 9.276 ;
  LAYER M3 ;
        RECT 1.728 6.768 1.76 9.276 ;
  LAYER M3 ;
        RECT 1.792 6.768 1.824 9.276 ;
  LAYER M3 ;
        RECT 1.856 6.768 1.888 9.276 ;
  LAYER M3 ;
        RECT 1.92 6.768 1.952 9.276 ;
  LAYER M3 ;
        RECT 1.984 6.768 2.016 9.276 ;
  LAYER M3 ;
        RECT 2.048 6.768 2.08 9.276 ;
  LAYER M3 ;
        RECT 2.112 6.768 2.144 9.276 ;
  LAYER M3 ;
        RECT 2.176 6.768 2.208 9.276 ;
  LAYER M3 ;
        RECT 2.24 6.768 2.272 9.276 ;
  LAYER M3 ;
        RECT 2.304 6.768 2.336 9.276 ;
  LAYER M3 ;
        RECT 2.368 6.768 2.4 9.276 ;
  LAYER M3 ;
        RECT 2.432 6.768 2.464 9.276 ;
  LAYER M3 ;
        RECT 2.496 6.768 2.528 9.276 ;
  LAYER M3 ;
        RECT 2.56 6.768 2.592 9.276 ;
  LAYER M3 ;
        RECT 2.624 6.768 2.656 9.276 ;
  LAYER M3 ;
        RECT 2.688 6.768 2.72 9.276 ;
  LAYER M3 ;
        RECT 2.784 6.768 2.816 9.276 ;
  LAYER M1 ;
        RECT 0.399 6.804 0.401 9.24 ;
  LAYER M1 ;
        RECT 0.479 6.804 0.481 9.24 ;
  LAYER M1 ;
        RECT 0.559 6.804 0.561 9.24 ;
  LAYER M1 ;
        RECT 0.639 6.804 0.641 9.24 ;
  LAYER M1 ;
        RECT 0.719 6.804 0.721 9.24 ;
  LAYER M1 ;
        RECT 0.799 6.804 0.801 9.24 ;
  LAYER M1 ;
        RECT 0.879 6.804 0.881 9.24 ;
  LAYER M1 ;
        RECT 0.959 6.804 0.961 9.24 ;
  LAYER M1 ;
        RECT 1.039 6.804 1.041 9.24 ;
  LAYER M1 ;
        RECT 1.119 6.804 1.121 9.24 ;
  LAYER M1 ;
        RECT 1.199 6.804 1.201 9.24 ;
  LAYER M1 ;
        RECT 1.279 6.804 1.281 9.24 ;
  LAYER M1 ;
        RECT 1.359 6.804 1.361 9.24 ;
  LAYER M1 ;
        RECT 1.439 6.804 1.441 9.24 ;
  LAYER M1 ;
        RECT 1.519 6.804 1.521 9.24 ;
  LAYER M1 ;
        RECT 1.599 6.804 1.601 9.24 ;
  LAYER M1 ;
        RECT 1.679 6.804 1.681 9.24 ;
  LAYER M1 ;
        RECT 1.759 6.804 1.761 9.24 ;
  LAYER M1 ;
        RECT 1.839 6.804 1.841 9.24 ;
  LAYER M1 ;
        RECT 1.919 6.804 1.921 9.24 ;
  LAYER M1 ;
        RECT 1.999 6.804 2.001 9.24 ;
  LAYER M1 ;
        RECT 2.079 6.804 2.081 9.24 ;
  LAYER M1 ;
        RECT 2.159 6.804 2.161 9.24 ;
  LAYER M1 ;
        RECT 2.239 6.804 2.241 9.24 ;
  LAYER M1 ;
        RECT 2.319 6.804 2.321 9.24 ;
  LAYER M1 ;
        RECT 2.399 6.804 2.401 9.24 ;
  LAYER M1 ;
        RECT 2.479 6.804 2.481 9.24 ;
  LAYER M1 ;
        RECT 2.559 6.804 2.561 9.24 ;
  LAYER M1 ;
        RECT 2.639 6.804 2.641 9.24 ;
  LAYER M1 ;
        RECT 2.719 6.804 2.721 9.24 ;
  LAYER M2 ;
        RECT 0.4 6.803 2.8 6.805 ;
  LAYER M2 ;
        RECT 0.4 6.887 2.8 6.889 ;
  LAYER M2 ;
        RECT 0.4 6.971 2.8 6.973 ;
  LAYER M2 ;
        RECT 0.4 7.055 2.8 7.057 ;
  LAYER M2 ;
        RECT 0.4 7.139 2.8 7.141 ;
  LAYER M2 ;
        RECT 0.4 7.223 2.8 7.225 ;
  LAYER M2 ;
        RECT 0.4 7.307 2.8 7.309 ;
  LAYER M2 ;
        RECT 0.4 7.391 2.8 7.393 ;
  LAYER M2 ;
        RECT 0.4 7.475 2.8 7.477 ;
  LAYER M2 ;
        RECT 0.4 7.559 2.8 7.561 ;
  LAYER M2 ;
        RECT 0.4 7.643 2.8 7.645 ;
  LAYER M2 ;
        RECT 0.4 7.727 2.8 7.729 ;
  LAYER M2 ;
        RECT 0.4 7.8105 2.8 7.8125 ;
  LAYER M2 ;
        RECT 0.4 7.895 2.8 7.897 ;
  LAYER M2 ;
        RECT 0.4 7.979 2.8 7.981 ;
  LAYER M2 ;
        RECT 0.4 8.063 2.8 8.065 ;
  LAYER M2 ;
        RECT 0.4 8.147 2.8 8.149 ;
  LAYER M2 ;
        RECT 0.4 8.231 2.8 8.233 ;
  LAYER M2 ;
        RECT 0.4 8.315 2.8 8.317 ;
  LAYER M2 ;
        RECT 0.4 8.399 2.8 8.401 ;
  LAYER M2 ;
        RECT 0.4 8.483 2.8 8.485 ;
  LAYER M2 ;
        RECT 0.4 8.567 2.8 8.569 ;
  LAYER M2 ;
        RECT 0.4 8.651 2.8 8.653 ;
  LAYER M2 ;
        RECT 0.4 8.735 2.8 8.737 ;
  LAYER M2 ;
        RECT 0.4 8.819 2.8 8.821 ;
  LAYER M2 ;
        RECT 0.4 8.903 2.8 8.905 ;
  LAYER M2 ;
        RECT 0.4 8.987 2.8 8.989 ;
  LAYER M2 ;
        RECT 0.4 9.071 2.8 9.073 ;
  LAYER M2 ;
        RECT 0.4 9.155 2.8 9.157 ;
  LAYER M1 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M1 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M1 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M1 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M1 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M1 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M1 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M1 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M1 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M1 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M1 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M1 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M1 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M1 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M1 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M1 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M1 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M1 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M1 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M1 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M1 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M1 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M1 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M1 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M1 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M1 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M1 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M1 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M1 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M1 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M1 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M1 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M1 ;
        RECT 2.432 9.708 2.464 12.216 ;
  LAYER M1 ;
        RECT 2.496 9.708 2.528 12.216 ;
  LAYER M1 ;
        RECT 2.56 9.708 2.592 12.216 ;
  LAYER M1 ;
        RECT 2.624 9.708 2.656 12.216 ;
  LAYER M1 ;
        RECT 2.688 9.708 2.72 12.216 ;
  LAYER M2 ;
        RECT 0.364 9.792 2.836 9.824 ;
  LAYER M2 ;
        RECT 0.364 9.856 2.836 9.888 ;
  LAYER M2 ;
        RECT 0.364 9.92 2.836 9.952 ;
  LAYER M2 ;
        RECT 0.364 9.984 2.836 10.016 ;
  LAYER M2 ;
        RECT 0.364 10.048 2.836 10.08 ;
  LAYER M2 ;
        RECT 0.364 10.112 2.836 10.144 ;
  LAYER M2 ;
        RECT 0.364 10.176 2.836 10.208 ;
  LAYER M2 ;
        RECT 0.364 10.24 2.836 10.272 ;
  LAYER M2 ;
        RECT 0.364 10.304 2.836 10.336 ;
  LAYER M2 ;
        RECT 0.364 10.368 2.836 10.4 ;
  LAYER M2 ;
        RECT 0.364 10.432 2.836 10.464 ;
  LAYER M2 ;
        RECT 0.364 10.496 2.836 10.528 ;
  LAYER M2 ;
        RECT 0.364 10.56 2.836 10.592 ;
  LAYER M2 ;
        RECT 0.364 10.624 2.836 10.656 ;
  LAYER M2 ;
        RECT 0.364 10.688 2.836 10.72 ;
  LAYER M2 ;
        RECT 0.364 10.752 2.836 10.784 ;
  LAYER M2 ;
        RECT 0.364 10.816 2.836 10.848 ;
  LAYER M2 ;
        RECT 0.364 10.88 2.836 10.912 ;
  LAYER M2 ;
        RECT 0.364 10.944 2.836 10.976 ;
  LAYER M2 ;
        RECT 0.364 11.008 2.836 11.04 ;
  LAYER M2 ;
        RECT 0.364 11.072 2.836 11.104 ;
  LAYER M2 ;
        RECT 0.364 11.136 2.836 11.168 ;
  LAYER M2 ;
        RECT 0.364 11.2 2.836 11.232 ;
  LAYER M2 ;
        RECT 0.364 11.264 2.836 11.296 ;
  LAYER M2 ;
        RECT 0.364 11.328 2.836 11.36 ;
  LAYER M2 ;
        RECT 0.364 11.392 2.836 11.424 ;
  LAYER M2 ;
        RECT 0.364 11.456 2.836 11.488 ;
  LAYER M2 ;
        RECT 0.364 11.52 2.836 11.552 ;
  LAYER M2 ;
        RECT 0.364 11.584 2.836 11.616 ;
  LAYER M2 ;
        RECT 0.364 11.648 2.836 11.68 ;
  LAYER M2 ;
        RECT 0.364 11.712 2.836 11.744 ;
  LAYER M2 ;
        RECT 0.364 11.776 2.836 11.808 ;
  LAYER M2 ;
        RECT 0.364 11.84 2.836 11.872 ;
  LAYER M2 ;
        RECT 0.364 11.904 2.836 11.936 ;
  LAYER M2 ;
        RECT 0.364 11.968 2.836 12 ;
  LAYER M2 ;
        RECT 0.364 12.032 2.836 12.064 ;
  LAYER M3 ;
        RECT 0.384 9.708 0.416 12.216 ;
  LAYER M3 ;
        RECT 0.448 9.708 0.48 12.216 ;
  LAYER M3 ;
        RECT 0.512 9.708 0.544 12.216 ;
  LAYER M3 ;
        RECT 0.576 9.708 0.608 12.216 ;
  LAYER M3 ;
        RECT 0.64 9.708 0.672 12.216 ;
  LAYER M3 ;
        RECT 0.704 9.708 0.736 12.216 ;
  LAYER M3 ;
        RECT 0.768 9.708 0.8 12.216 ;
  LAYER M3 ;
        RECT 0.832 9.708 0.864 12.216 ;
  LAYER M3 ;
        RECT 0.896 9.708 0.928 12.216 ;
  LAYER M3 ;
        RECT 0.96 9.708 0.992 12.216 ;
  LAYER M3 ;
        RECT 1.024 9.708 1.056 12.216 ;
  LAYER M3 ;
        RECT 1.088 9.708 1.12 12.216 ;
  LAYER M3 ;
        RECT 1.152 9.708 1.184 12.216 ;
  LAYER M3 ;
        RECT 1.216 9.708 1.248 12.216 ;
  LAYER M3 ;
        RECT 1.28 9.708 1.312 12.216 ;
  LAYER M3 ;
        RECT 1.344 9.708 1.376 12.216 ;
  LAYER M3 ;
        RECT 1.408 9.708 1.44 12.216 ;
  LAYER M3 ;
        RECT 1.472 9.708 1.504 12.216 ;
  LAYER M3 ;
        RECT 1.536 9.708 1.568 12.216 ;
  LAYER M3 ;
        RECT 1.6 9.708 1.632 12.216 ;
  LAYER M3 ;
        RECT 1.664 9.708 1.696 12.216 ;
  LAYER M3 ;
        RECT 1.728 9.708 1.76 12.216 ;
  LAYER M3 ;
        RECT 1.792 9.708 1.824 12.216 ;
  LAYER M3 ;
        RECT 1.856 9.708 1.888 12.216 ;
  LAYER M3 ;
        RECT 1.92 9.708 1.952 12.216 ;
  LAYER M3 ;
        RECT 1.984 9.708 2.016 12.216 ;
  LAYER M3 ;
        RECT 2.048 9.708 2.08 12.216 ;
  LAYER M3 ;
        RECT 2.112 9.708 2.144 12.216 ;
  LAYER M3 ;
        RECT 2.176 9.708 2.208 12.216 ;
  LAYER M3 ;
        RECT 2.24 9.708 2.272 12.216 ;
  LAYER M3 ;
        RECT 2.304 9.708 2.336 12.216 ;
  LAYER M3 ;
        RECT 2.368 9.708 2.4 12.216 ;
  LAYER M3 ;
        RECT 2.432 9.708 2.464 12.216 ;
  LAYER M3 ;
        RECT 2.496 9.708 2.528 12.216 ;
  LAYER M3 ;
        RECT 2.56 9.708 2.592 12.216 ;
  LAYER M3 ;
        RECT 2.624 9.708 2.656 12.216 ;
  LAYER M3 ;
        RECT 2.688 9.708 2.72 12.216 ;
  LAYER M3 ;
        RECT 2.784 9.708 2.816 12.216 ;
  LAYER M1 ;
        RECT 0.399 9.744 0.401 12.18 ;
  LAYER M1 ;
        RECT 0.479 9.744 0.481 12.18 ;
  LAYER M1 ;
        RECT 0.559 9.744 0.561 12.18 ;
  LAYER M1 ;
        RECT 0.639 9.744 0.641 12.18 ;
  LAYER M1 ;
        RECT 0.719 9.744 0.721 12.18 ;
  LAYER M1 ;
        RECT 0.799 9.744 0.801 12.18 ;
  LAYER M1 ;
        RECT 0.879 9.744 0.881 12.18 ;
  LAYER M1 ;
        RECT 0.959 9.744 0.961 12.18 ;
  LAYER M1 ;
        RECT 1.039 9.744 1.041 12.18 ;
  LAYER M1 ;
        RECT 1.119 9.744 1.121 12.18 ;
  LAYER M1 ;
        RECT 1.199 9.744 1.201 12.18 ;
  LAYER M1 ;
        RECT 1.279 9.744 1.281 12.18 ;
  LAYER M1 ;
        RECT 1.359 9.744 1.361 12.18 ;
  LAYER M1 ;
        RECT 1.439 9.744 1.441 12.18 ;
  LAYER M1 ;
        RECT 1.519 9.744 1.521 12.18 ;
  LAYER M1 ;
        RECT 1.599 9.744 1.601 12.18 ;
  LAYER M1 ;
        RECT 1.679 9.744 1.681 12.18 ;
  LAYER M1 ;
        RECT 1.759 9.744 1.761 12.18 ;
  LAYER M1 ;
        RECT 1.839 9.744 1.841 12.18 ;
  LAYER M1 ;
        RECT 1.919 9.744 1.921 12.18 ;
  LAYER M1 ;
        RECT 1.999 9.744 2.001 12.18 ;
  LAYER M1 ;
        RECT 2.079 9.744 2.081 12.18 ;
  LAYER M1 ;
        RECT 2.159 9.744 2.161 12.18 ;
  LAYER M1 ;
        RECT 2.239 9.744 2.241 12.18 ;
  LAYER M1 ;
        RECT 2.319 9.744 2.321 12.18 ;
  LAYER M1 ;
        RECT 2.399 9.744 2.401 12.18 ;
  LAYER M1 ;
        RECT 2.479 9.744 2.481 12.18 ;
  LAYER M1 ;
        RECT 2.559 9.744 2.561 12.18 ;
  LAYER M1 ;
        RECT 2.639 9.744 2.641 12.18 ;
  LAYER M1 ;
        RECT 2.719 9.744 2.721 12.18 ;
  LAYER M2 ;
        RECT 0.4 9.743 2.8 9.745 ;
  LAYER M2 ;
        RECT 0.4 9.827 2.8 9.829 ;
  LAYER M2 ;
        RECT 0.4 9.911 2.8 9.913 ;
  LAYER M2 ;
        RECT 0.4 9.995 2.8 9.997 ;
  LAYER M2 ;
        RECT 0.4 10.079 2.8 10.081 ;
  LAYER M2 ;
        RECT 0.4 10.163 2.8 10.165 ;
  LAYER M2 ;
        RECT 0.4 10.247 2.8 10.249 ;
  LAYER M2 ;
        RECT 0.4 10.331 2.8 10.333 ;
  LAYER M2 ;
        RECT 0.4 10.415 2.8 10.417 ;
  LAYER M2 ;
        RECT 0.4 10.499 2.8 10.501 ;
  LAYER M2 ;
        RECT 0.4 10.583 2.8 10.585 ;
  LAYER M2 ;
        RECT 0.4 10.667 2.8 10.669 ;
  LAYER M2 ;
        RECT 0.4 10.7505 2.8 10.7525 ;
  LAYER M2 ;
        RECT 0.4 10.835 2.8 10.837 ;
  LAYER M2 ;
        RECT 0.4 10.919 2.8 10.921 ;
  LAYER M2 ;
        RECT 0.4 11.003 2.8 11.005 ;
  LAYER M2 ;
        RECT 0.4 11.087 2.8 11.089 ;
  LAYER M2 ;
        RECT 0.4 11.171 2.8 11.173 ;
  LAYER M2 ;
        RECT 0.4 11.255 2.8 11.257 ;
  LAYER M2 ;
        RECT 0.4 11.339 2.8 11.341 ;
  LAYER M2 ;
        RECT 0.4 11.423 2.8 11.425 ;
  LAYER M2 ;
        RECT 0.4 11.507 2.8 11.509 ;
  LAYER M2 ;
        RECT 0.4 11.591 2.8 11.593 ;
  LAYER M2 ;
        RECT 0.4 11.675 2.8 11.677 ;
  LAYER M2 ;
        RECT 0.4 11.759 2.8 11.761 ;
  LAYER M2 ;
        RECT 0.4 11.843 2.8 11.845 ;
  LAYER M2 ;
        RECT 0.4 11.927 2.8 11.929 ;
  LAYER M2 ;
        RECT 0.4 12.011 2.8 12.013 ;
  LAYER M2 ;
        RECT 0.4 12.095 2.8 12.097 ;
  LAYER M1 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M1 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M1 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M1 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M1 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M1 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M1 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M1 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M1 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M1 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M1 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M1 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M1 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M1 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M1 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M1 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M1 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M1 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M1 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M1 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M1 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M1 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M1 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M1 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M1 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M1 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M1 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M1 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M1 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M1 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M1 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M1 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M1 ;
        RECT 2.432 12.648 2.464 15.156 ;
  LAYER M1 ;
        RECT 2.496 12.648 2.528 15.156 ;
  LAYER M1 ;
        RECT 2.56 12.648 2.592 15.156 ;
  LAYER M1 ;
        RECT 2.624 12.648 2.656 15.156 ;
  LAYER M1 ;
        RECT 2.688 12.648 2.72 15.156 ;
  LAYER M2 ;
        RECT 0.364 12.732 2.836 12.764 ;
  LAYER M2 ;
        RECT 0.364 12.796 2.836 12.828 ;
  LAYER M2 ;
        RECT 0.364 12.86 2.836 12.892 ;
  LAYER M2 ;
        RECT 0.364 12.924 2.836 12.956 ;
  LAYER M2 ;
        RECT 0.364 12.988 2.836 13.02 ;
  LAYER M2 ;
        RECT 0.364 13.052 2.836 13.084 ;
  LAYER M2 ;
        RECT 0.364 13.116 2.836 13.148 ;
  LAYER M2 ;
        RECT 0.364 13.18 2.836 13.212 ;
  LAYER M2 ;
        RECT 0.364 13.244 2.836 13.276 ;
  LAYER M2 ;
        RECT 0.364 13.308 2.836 13.34 ;
  LAYER M2 ;
        RECT 0.364 13.372 2.836 13.404 ;
  LAYER M2 ;
        RECT 0.364 13.436 2.836 13.468 ;
  LAYER M2 ;
        RECT 0.364 13.5 2.836 13.532 ;
  LAYER M2 ;
        RECT 0.364 13.564 2.836 13.596 ;
  LAYER M2 ;
        RECT 0.364 13.628 2.836 13.66 ;
  LAYER M2 ;
        RECT 0.364 13.692 2.836 13.724 ;
  LAYER M2 ;
        RECT 0.364 13.756 2.836 13.788 ;
  LAYER M2 ;
        RECT 0.364 13.82 2.836 13.852 ;
  LAYER M2 ;
        RECT 0.364 13.884 2.836 13.916 ;
  LAYER M2 ;
        RECT 0.364 13.948 2.836 13.98 ;
  LAYER M2 ;
        RECT 0.364 14.012 2.836 14.044 ;
  LAYER M2 ;
        RECT 0.364 14.076 2.836 14.108 ;
  LAYER M2 ;
        RECT 0.364 14.14 2.836 14.172 ;
  LAYER M2 ;
        RECT 0.364 14.204 2.836 14.236 ;
  LAYER M2 ;
        RECT 0.364 14.268 2.836 14.3 ;
  LAYER M2 ;
        RECT 0.364 14.332 2.836 14.364 ;
  LAYER M2 ;
        RECT 0.364 14.396 2.836 14.428 ;
  LAYER M2 ;
        RECT 0.364 14.46 2.836 14.492 ;
  LAYER M2 ;
        RECT 0.364 14.524 2.836 14.556 ;
  LAYER M2 ;
        RECT 0.364 14.588 2.836 14.62 ;
  LAYER M2 ;
        RECT 0.364 14.652 2.836 14.684 ;
  LAYER M2 ;
        RECT 0.364 14.716 2.836 14.748 ;
  LAYER M2 ;
        RECT 0.364 14.78 2.836 14.812 ;
  LAYER M2 ;
        RECT 0.364 14.844 2.836 14.876 ;
  LAYER M2 ;
        RECT 0.364 14.908 2.836 14.94 ;
  LAYER M2 ;
        RECT 0.364 14.972 2.836 15.004 ;
  LAYER M3 ;
        RECT 0.384 12.648 0.416 15.156 ;
  LAYER M3 ;
        RECT 0.448 12.648 0.48 15.156 ;
  LAYER M3 ;
        RECT 0.512 12.648 0.544 15.156 ;
  LAYER M3 ;
        RECT 0.576 12.648 0.608 15.156 ;
  LAYER M3 ;
        RECT 0.64 12.648 0.672 15.156 ;
  LAYER M3 ;
        RECT 0.704 12.648 0.736 15.156 ;
  LAYER M3 ;
        RECT 0.768 12.648 0.8 15.156 ;
  LAYER M3 ;
        RECT 0.832 12.648 0.864 15.156 ;
  LAYER M3 ;
        RECT 0.896 12.648 0.928 15.156 ;
  LAYER M3 ;
        RECT 0.96 12.648 0.992 15.156 ;
  LAYER M3 ;
        RECT 1.024 12.648 1.056 15.156 ;
  LAYER M3 ;
        RECT 1.088 12.648 1.12 15.156 ;
  LAYER M3 ;
        RECT 1.152 12.648 1.184 15.156 ;
  LAYER M3 ;
        RECT 1.216 12.648 1.248 15.156 ;
  LAYER M3 ;
        RECT 1.28 12.648 1.312 15.156 ;
  LAYER M3 ;
        RECT 1.344 12.648 1.376 15.156 ;
  LAYER M3 ;
        RECT 1.408 12.648 1.44 15.156 ;
  LAYER M3 ;
        RECT 1.472 12.648 1.504 15.156 ;
  LAYER M3 ;
        RECT 1.536 12.648 1.568 15.156 ;
  LAYER M3 ;
        RECT 1.6 12.648 1.632 15.156 ;
  LAYER M3 ;
        RECT 1.664 12.648 1.696 15.156 ;
  LAYER M3 ;
        RECT 1.728 12.648 1.76 15.156 ;
  LAYER M3 ;
        RECT 1.792 12.648 1.824 15.156 ;
  LAYER M3 ;
        RECT 1.856 12.648 1.888 15.156 ;
  LAYER M3 ;
        RECT 1.92 12.648 1.952 15.156 ;
  LAYER M3 ;
        RECT 1.984 12.648 2.016 15.156 ;
  LAYER M3 ;
        RECT 2.048 12.648 2.08 15.156 ;
  LAYER M3 ;
        RECT 2.112 12.648 2.144 15.156 ;
  LAYER M3 ;
        RECT 2.176 12.648 2.208 15.156 ;
  LAYER M3 ;
        RECT 2.24 12.648 2.272 15.156 ;
  LAYER M3 ;
        RECT 2.304 12.648 2.336 15.156 ;
  LAYER M3 ;
        RECT 2.368 12.648 2.4 15.156 ;
  LAYER M3 ;
        RECT 2.432 12.648 2.464 15.156 ;
  LAYER M3 ;
        RECT 2.496 12.648 2.528 15.156 ;
  LAYER M3 ;
        RECT 2.56 12.648 2.592 15.156 ;
  LAYER M3 ;
        RECT 2.624 12.648 2.656 15.156 ;
  LAYER M3 ;
        RECT 2.688 12.648 2.72 15.156 ;
  LAYER M3 ;
        RECT 2.784 12.648 2.816 15.156 ;
  LAYER M1 ;
        RECT 0.399 12.684 0.401 15.12 ;
  LAYER M1 ;
        RECT 0.479 12.684 0.481 15.12 ;
  LAYER M1 ;
        RECT 0.559 12.684 0.561 15.12 ;
  LAYER M1 ;
        RECT 0.639 12.684 0.641 15.12 ;
  LAYER M1 ;
        RECT 0.719 12.684 0.721 15.12 ;
  LAYER M1 ;
        RECT 0.799 12.684 0.801 15.12 ;
  LAYER M1 ;
        RECT 0.879 12.684 0.881 15.12 ;
  LAYER M1 ;
        RECT 0.959 12.684 0.961 15.12 ;
  LAYER M1 ;
        RECT 1.039 12.684 1.041 15.12 ;
  LAYER M1 ;
        RECT 1.119 12.684 1.121 15.12 ;
  LAYER M1 ;
        RECT 1.199 12.684 1.201 15.12 ;
  LAYER M1 ;
        RECT 1.279 12.684 1.281 15.12 ;
  LAYER M1 ;
        RECT 1.359 12.684 1.361 15.12 ;
  LAYER M1 ;
        RECT 1.439 12.684 1.441 15.12 ;
  LAYER M1 ;
        RECT 1.519 12.684 1.521 15.12 ;
  LAYER M1 ;
        RECT 1.599 12.684 1.601 15.12 ;
  LAYER M1 ;
        RECT 1.679 12.684 1.681 15.12 ;
  LAYER M1 ;
        RECT 1.759 12.684 1.761 15.12 ;
  LAYER M1 ;
        RECT 1.839 12.684 1.841 15.12 ;
  LAYER M1 ;
        RECT 1.919 12.684 1.921 15.12 ;
  LAYER M1 ;
        RECT 1.999 12.684 2.001 15.12 ;
  LAYER M1 ;
        RECT 2.079 12.684 2.081 15.12 ;
  LAYER M1 ;
        RECT 2.159 12.684 2.161 15.12 ;
  LAYER M1 ;
        RECT 2.239 12.684 2.241 15.12 ;
  LAYER M1 ;
        RECT 2.319 12.684 2.321 15.12 ;
  LAYER M1 ;
        RECT 2.399 12.684 2.401 15.12 ;
  LAYER M1 ;
        RECT 2.479 12.684 2.481 15.12 ;
  LAYER M1 ;
        RECT 2.559 12.684 2.561 15.12 ;
  LAYER M1 ;
        RECT 2.639 12.684 2.641 15.12 ;
  LAYER M1 ;
        RECT 2.719 12.684 2.721 15.12 ;
  LAYER M2 ;
        RECT 0.4 12.683 2.8 12.685 ;
  LAYER M2 ;
        RECT 0.4 12.767 2.8 12.769 ;
  LAYER M2 ;
        RECT 0.4 12.851 2.8 12.853 ;
  LAYER M2 ;
        RECT 0.4 12.935 2.8 12.937 ;
  LAYER M2 ;
        RECT 0.4 13.019 2.8 13.021 ;
  LAYER M2 ;
        RECT 0.4 13.103 2.8 13.105 ;
  LAYER M2 ;
        RECT 0.4 13.187 2.8 13.189 ;
  LAYER M2 ;
        RECT 0.4 13.271 2.8 13.273 ;
  LAYER M2 ;
        RECT 0.4 13.355 2.8 13.357 ;
  LAYER M2 ;
        RECT 0.4 13.439 2.8 13.441 ;
  LAYER M2 ;
        RECT 0.4 13.523 2.8 13.525 ;
  LAYER M2 ;
        RECT 0.4 13.607 2.8 13.609 ;
  LAYER M2 ;
        RECT 0.4 13.6905 2.8 13.6925 ;
  LAYER M2 ;
        RECT 0.4 13.775 2.8 13.777 ;
  LAYER M2 ;
        RECT 0.4 13.859 2.8 13.861 ;
  LAYER M2 ;
        RECT 0.4 13.943 2.8 13.945 ;
  LAYER M2 ;
        RECT 0.4 14.027 2.8 14.029 ;
  LAYER M2 ;
        RECT 0.4 14.111 2.8 14.113 ;
  LAYER M2 ;
        RECT 0.4 14.195 2.8 14.197 ;
  LAYER M2 ;
        RECT 0.4 14.279 2.8 14.281 ;
  LAYER M2 ;
        RECT 0.4 14.363 2.8 14.365 ;
  LAYER M2 ;
        RECT 0.4 14.447 2.8 14.449 ;
  LAYER M2 ;
        RECT 0.4 14.531 2.8 14.533 ;
  LAYER M2 ;
        RECT 0.4 14.615 2.8 14.617 ;
  LAYER M2 ;
        RECT 0.4 14.699 2.8 14.701 ;
  LAYER M2 ;
        RECT 0.4 14.783 2.8 14.785 ;
  LAYER M2 ;
        RECT 0.4 14.867 2.8 14.869 ;
  LAYER M2 ;
        RECT 0.4 14.951 2.8 14.953 ;
  LAYER M2 ;
        RECT 0.4 15.035 2.8 15.037 ;
  LAYER M1 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M1 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M1 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M1 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M1 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M1 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M1 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M1 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M1 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M1 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M1 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M1 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M1 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M1 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M1 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M1 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M1 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M1 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M1 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M1 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M1 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M1 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M1 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M1 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M1 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M1 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M1 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M1 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M1 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M1 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M1 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M1 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M1 ;
        RECT 2.432 15.588 2.464 18.096 ;
  LAYER M1 ;
        RECT 2.496 15.588 2.528 18.096 ;
  LAYER M1 ;
        RECT 2.56 15.588 2.592 18.096 ;
  LAYER M1 ;
        RECT 2.624 15.588 2.656 18.096 ;
  LAYER M1 ;
        RECT 2.688 15.588 2.72 18.096 ;
  LAYER M2 ;
        RECT 0.364 15.672 2.836 15.704 ;
  LAYER M2 ;
        RECT 0.364 15.736 2.836 15.768 ;
  LAYER M2 ;
        RECT 0.364 15.8 2.836 15.832 ;
  LAYER M2 ;
        RECT 0.364 15.864 2.836 15.896 ;
  LAYER M2 ;
        RECT 0.364 15.928 2.836 15.96 ;
  LAYER M2 ;
        RECT 0.364 15.992 2.836 16.024 ;
  LAYER M2 ;
        RECT 0.364 16.056 2.836 16.088 ;
  LAYER M2 ;
        RECT 0.364 16.12 2.836 16.152 ;
  LAYER M2 ;
        RECT 0.364 16.184 2.836 16.216 ;
  LAYER M2 ;
        RECT 0.364 16.248 2.836 16.28 ;
  LAYER M2 ;
        RECT 0.364 16.312 2.836 16.344 ;
  LAYER M2 ;
        RECT 0.364 16.376 2.836 16.408 ;
  LAYER M2 ;
        RECT 0.364 16.44 2.836 16.472 ;
  LAYER M2 ;
        RECT 0.364 16.504 2.836 16.536 ;
  LAYER M2 ;
        RECT 0.364 16.568 2.836 16.6 ;
  LAYER M2 ;
        RECT 0.364 16.632 2.836 16.664 ;
  LAYER M2 ;
        RECT 0.364 16.696 2.836 16.728 ;
  LAYER M2 ;
        RECT 0.364 16.76 2.836 16.792 ;
  LAYER M2 ;
        RECT 0.364 16.824 2.836 16.856 ;
  LAYER M2 ;
        RECT 0.364 16.888 2.836 16.92 ;
  LAYER M2 ;
        RECT 0.364 16.952 2.836 16.984 ;
  LAYER M2 ;
        RECT 0.364 17.016 2.836 17.048 ;
  LAYER M2 ;
        RECT 0.364 17.08 2.836 17.112 ;
  LAYER M2 ;
        RECT 0.364 17.144 2.836 17.176 ;
  LAYER M2 ;
        RECT 0.364 17.208 2.836 17.24 ;
  LAYER M2 ;
        RECT 0.364 17.272 2.836 17.304 ;
  LAYER M2 ;
        RECT 0.364 17.336 2.836 17.368 ;
  LAYER M2 ;
        RECT 0.364 17.4 2.836 17.432 ;
  LAYER M2 ;
        RECT 0.364 17.464 2.836 17.496 ;
  LAYER M2 ;
        RECT 0.364 17.528 2.836 17.56 ;
  LAYER M2 ;
        RECT 0.364 17.592 2.836 17.624 ;
  LAYER M2 ;
        RECT 0.364 17.656 2.836 17.688 ;
  LAYER M2 ;
        RECT 0.364 17.72 2.836 17.752 ;
  LAYER M2 ;
        RECT 0.364 17.784 2.836 17.816 ;
  LAYER M2 ;
        RECT 0.364 17.848 2.836 17.88 ;
  LAYER M2 ;
        RECT 0.364 17.912 2.836 17.944 ;
  LAYER M3 ;
        RECT 0.384 15.588 0.416 18.096 ;
  LAYER M3 ;
        RECT 0.448 15.588 0.48 18.096 ;
  LAYER M3 ;
        RECT 0.512 15.588 0.544 18.096 ;
  LAYER M3 ;
        RECT 0.576 15.588 0.608 18.096 ;
  LAYER M3 ;
        RECT 0.64 15.588 0.672 18.096 ;
  LAYER M3 ;
        RECT 0.704 15.588 0.736 18.096 ;
  LAYER M3 ;
        RECT 0.768 15.588 0.8 18.096 ;
  LAYER M3 ;
        RECT 0.832 15.588 0.864 18.096 ;
  LAYER M3 ;
        RECT 0.896 15.588 0.928 18.096 ;
  LAYER M3 ;
        RECT 0.96 15.588 0.992 18.096 ;
  LAYER M3 ;
        RECT 1.024 15.588 1.056 18.096 ;
  LAYER M3 ;
        RECT 1.088 15.588 1.12 18.096 ;
  LAYER M3 ;
        RECT 1.152 15.588 1.184 18.096 ;
  LAYER M3 ;
        RECT 1.216 15.588 1.248 18.096 ;
  LAYER M3 ;
        RECT 1.28 15.588 1.312 18.096 ;
  LAYER M3 ;
        RECT 1.344 15.588 1.376 18.096 ;
  LAYER M3 ;
        RECT 1.408 15.588 1.44 18.096 ;
  LAYER M3 ;
        RECT 1.472 15.588 1.504 18.096 ;
  LAYER M3 ;
        RECT 1.536 15.588 1.568 18.096 ;
  LAYER M3 ;
        RECT 1.6 15.588 1.632 18.096 ;
  LAYER M3 ;
        RECT 1.664 15.588 1.696 18.096 ;
  LAYER M3 ;
        RECT 1.728 15.588 1.76 18.096 ;
  LAYER M3 ;
        RECT 1.792 15.588 1.824 18.096 ;
  LAYER M3 ;
        RECT 1.856 15.588 1.888 18.096 ;
  LAYER M3 ;
        RECT 1.92 15.588 1.952 18.096 ;
  LAYER M3 ;
        RECT 1.984 15.588 2.016 18.096 ;
  LAYER M3 ;
        RECT 2.048 15.588 2.08 18.096 ;
  LAYER M3 ;
        RECT 2.112 15.588 2.144 18.096 ;
  LAYER M3 ;
        RECT 2.176 15.588 2.208 18.096 ;
  LAYER M3 ;
        RECT 2.24 15.588 2.272 18.096 ;
  LAYER M3 ;
        RECT 2.304 15.588 2.336 18.096 ;
  LAYER M3 ;
        RECT 2.368 15.588 2.4 18.096 ;
  LAYER M3 ;
        RECT 2.432 15.588 2.464 18.096 ;
  LAYER M3 ;
        RECT 2.496 15.588 2.528 18.096 ;
  LAYER M3 ;
        RECT 2.56 15.588 2.592 18.096 ;
  LAYER M3 ;
        RECT 2.624 15.588 2.656 18.096 ;
  LAYER M3 ;
        RECT 2.688 15.588 2.72 18.096 ;
  LAYER M3 ;
        RECT 2.784 15.588 2.816 18.096 ;
  LAYER M1 ;
        RECT 0.399 15.624 0.401 18.06 ;
  LAYER M1 ;
        RECT 0.479 15.624 0.481 18.06 ;
  LAYER M1 ;
        RECT 0.559 15.624 0.561 18.06 ;
  LAYER M1 ;
        RECT 0.639 15.624 0.641 18.06 ;
  LAYER M1 ;
        RECT 0.719 15.624 0.721 18.06 ;
  LAYER M1 ;
        RECT 0.799 15.624 0.801 18.06 ;
  LAYER M1 ;
        RECT 0.879 15.624 0.881 18.06 ;
  LAYER M1 ;
        RECT 0.959 15.624 0.961 18.06 ;
  LAYER M1 ;
        RECT 1.039 15.624 1.041 18.06 ;
  LAYER M1 ;
        RECT 1.119 15.624 1.121 18.06 ;
  LAYER M1 ;
        RECT 1.199 15.624 1.201 18.06 ;
  LAYER M1 ;
        RECT 1.279 15.624 1.281 18.06 ;
  LAYER M1 ;
        RECT 1.359 15.624 1.361 18.06 ;
  LAYER M1 ;
        RECT 1.439 15.624 1.441 18.06 ;
  LAYER M1 ;
        RECT 1.519 15.624 1.521 18.06 ;
  LAYER M1 ;
        RECT 1.599 15.624 1.601 18.06 ;
  LAYER M1 ;
        RECT 1.679 15.624 1.681 18.06 ;
  LAYER M1 ;
        RECT 1.759 15.624 1.761 18.06 ;
  LAYER M1 ;
        RECT 1.839 15.624 1.841 18.06 ;
  LAYER M1 ;
        RECT 1.919 15.624 1.921 18.06 ;
  LAYER M1 ;
        RECT 1.999 15.624 2.001 18.06 ;
  LAYER M1 ;
        RECT 2.079 15.624 2.081 18.06 ;
  LAYER M1 ;
        RECT 2.159 15.624 2.161 18.06 ;
  LAYER M1 ;
        RECT 2.239 15.624 2.241 18.06 ;
  LAYER M1 ;
        RECT 2.319 15.624 2.321 18.06 ;
  LAYER M1 ;
        RECT 2.399 15.624 2.401 18.06 ;
  LAYER M1 ;
        RECT 2.479 15.624 2.481 18.06 ;
  LAYER M1 ;
        RECT 2.559 15.624 2.561 18.06 ;
  LAYER M1 ;
        RECT 2.639 15.624 2.641 18.06 ;
  LAYER M1 ;
        RECT 2.719 15.624 2.721 18.06 ;
  LAYER M2 ;
        RECT 0.4 15.623 2.8 15.625 ;
  LAYER M2 ;
        RECT 0.4 15.707 2.8 15.709 ;
  LAYER M2 ;
        RECT 0.4 15.791 2.8 15.793 ;
  LAYER M2 ;
        RECT 0.4 15.875 2.8 15.877 ;
  LAYER M2 ;
        RECT 0.4 15.959 2.8 15.961 ;
  LAYER M2 ;
        RECT 0.4 16.043 2.8 16.045 ;
  LAYER M2 ;
        RECT 0.4 16.127 2.8 16.129 ;
  LAYER M2 ;
        RECT 0.4 16.211 2.8 16.213 ;
  LAYER M2 ;
        RECT 0.4 16.295 2.8 16.297 ;
  LAYER M2 ;
        RECT 0.4 16.379 2.8 16.381 ;
  LAYER M2 ;
        RECT 0.4 16.463 2.8 16.465 ;
  LAYER M2 ;
        RECT 0.4 16.547 2.8 16.549 ;
  LAYER M2 ;
        RECT 0.4 16.6305 2.8 16.6325 ;
  LAYER M2 ;
        RECT 0.4 16.715 2.8 16.717 ;
  LAYER M2 ;
        RECT 0.4 16.799 2.8 16.801 ;
  LAYER M2 ;
        RECT 0.4 16.883 2.8 16.885 ;
  LAYER M2 ;
        RECT 0.4 16.967 2.8 16.969 ;
  LAYER M2 ;
        RECT 0.4 17.051 2.8 17.053 ;
  LAYER M2 ;
        RECT 0.4 17.135 2.8 17.137 ;
  LAYER M2 ;
        RECT 0.4 17.219 2.8 17.221 ;
  LAYER M2 ;
        RECT 0.4 17.303 2.8 17.305 ;
  LAYER M2 ;
        RECT 0.4 17.387 2.8 17.389 ;
  LAYER M2 ;
        RECT 0.4 17.471 2.8 17.473 ;
  LAYER M2 ;
        RECT 0.4 17.555 2.8 17.557 ;
  LAYER M2 ;
        RECT 0.4 17.639 2.8 17.641 ;
  LAYER M2 ;
        RECT 0.4 17.723 2.8 17.725 ;
  LAYER M2 ;
        RECT 0.4 17.807 2.8 17.809 ;
  LAYER M2 ;
        RECT 0.4 17.891 2.8 17.893 ;
  LAYER M2 ;
        RECT 0.4 17.975 2.8 17.977 ;
  LAYER M1 ;
        RECT 3.264 0.888 3.296 3.396 ;
  LAYER M1 ;
        RECT 3.328 0.888 3.36 3.396 ;
  LAYER M1 ;
        RECT 3.392 0.888 3.424 3.396 ;
  LAYER M1 ;
        RECT 3.456 0.888 3.488 3.396 ;
  LAYER M1 ;
        RECT 3.52 0.888 3.552 3.396 ;
  LAYER M1 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M1 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M1 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M1 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M1 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M1 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M1 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M1 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M1 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M1 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M1 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M1 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M1 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M1 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M1 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M1 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M1 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M1 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M1 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M1 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M1 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M1 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M1 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M1 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M1 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M1 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M1 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M1 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M1 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M1 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M1 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M1 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M2 ;
        RECT 3.244 0.972 5.716 1.004 ;
  LAYER M2 ;
        RECT 3.244 1.036 5.716 1.068 ;
  LAYER M2 ;
        RECT 3.244 1.1 5.716 1.132 ;
  LAYER M2 ;
        RECT 3.244 1.164 5.716 1.196 ;
  LAYER M2 ;
        RECT 3.244 1.228 5.716 1.26 ;
  LAYER M2 ;
        RECT 3.244 1.292 5.716 1.324 ;
  LAYER M2 ;
        RECT 3.244 1.356 5.716 1.388 ;
  LAYER M2 ;
        RECT 3.244 1.42 5.716 1.452 ;
  LAYER M2 ;
        RECT 3.244 1.484 5.716 1.516 ;
  LAYER M2 ;
        RECT 3.244 1.548 5.716 1.58 ;
  LAYER M2 ;
        RECT 3.244 1.612 5.716 1.644 ;
  LAYER M2 ;
        RECT 3.244 1.676 5.716 1.708 ;
  LAYER M2 ;
        RECT 3.244 1.74 5.716 1.772 ;
  LAYER M2 ;
        RECT 3.244 1.804 5.716 1.836 ;
  LAYER M2 ;
        RECT 3.244 1.868 5.716 1.9 ;
  LAYER M2 ;
        RECT 3.244 1.932 5.716 1.964 ;
  LAYER M2 ;
        RECT 3.244 1.996 5.716 2.028 ;
  LAYER M2 ;
        RECT 3.244 2.06 5.716 2.092 ;
  LAYER M2 ;
        RECT 3.244 2.124 5.716 2.156 ;
  LAYER M2 ;
        RECT 3.244 2.188 5.716 2.22 ;
  LAYER M2 ;
        RECT 3.244 2.252 5.716 2.284 ;
  LAYER M2 ;
        RECT 3.244 2.316 5.716 2.348 ;
  LAYER M2 ;
        RECT 3.244 2.38 5.716 2.412 ;
  LAYER M2 ;
        RECT 3.244 2.444 5.716 2.476 ;
  LAYER M2 ;
        RECT 3.244 2.508 5.716 2.54 ;
  LAYER M2 ;
        RECT 3.244 2.572 5.716 2.604 ;
  LAYER M2 ;
        RECT 3.244 2.636 5.716 2.668 ;
  LAYER M2 ;
        RECT 3.244 2.7 5.716 2.732 ;
  LAYER M2 ;
        RECT 3.244 2.764 5.716 2.796 ;
  LAYER M2 ;
        RECT 3.244 2.828 5.716 2.86 ;
  LAYER M2 ;
        RECT 3.244 2.892 5.716 2.924 ;
  LAYER M2 ;
        RECT 3.244 2.956 5.716 2.988 ;
  LAYER M2 ;
        RECT 3.244 3.02 5.716 3.052 ;
  LAYER M2 ;
        RECT 3.244 3.084 5.716 3.116 ;
  LAYER M2 ;
        RECT 3.244 3.148 5.716 3.18 ;
  LAYER M2 ;
        RECT 3.244 3.212 5.716 3.244 ;
  LAYER M3 ;
        RECT 3.264 0.888 3.296 3.396 ;
  LAYER M3 ;
        RECT 3.328 0.888 3.36 3.396 ;
  LAYER M3 ;
        RECT 3.392 0.888 3.424 3.396 ;
  LAYER M3 ;
        RECT 3.456 0.888 3.488 3.396 ;
  LAYER M3 ;
        RECT 3.52 0.888 3.552 3.396 ;
  LAYER M3 ;
        RECT 3.584 0.888 3.616 3.396 ;
  LAYER M3 ;
        RECT 3.648 0.888 3.68 3.396 ;
  LAYER M3 ;
        RECT 3.712 0.888 3.744 3.396 ;
  LAYER M3 ;
        RECT 3.776 0.888 3.808 3.396 ;
  LAYER M3 ;
        RECT 3.84 0.888 3.872 3.396 ;
  LAYER M3 ;
        RECT 3.904 0.888 3.936 3.396 ;
  LAYER M3 ;
        RECT 3.968 0.888 4 3.396 ;
  LAYER M3 ;
        RECT 4.032 0.888 4.064 3.396 ;
  LAYER M3 ;
        RECT 4.096 0.888 4.128 3.396 ;
  LAYER M3 ;
        RECT 4.16 0.888 4.192 3.396 ;
  LAYER M3 ;
        RECT 4.224 0.888 4.256 3.396 ;
  LAYER M3 ;
        RECT 4.288 0.888 4.32 3.396 ;
  LAYER M3 ;
        RECT 4.352 0.888 4.384 3.396 ;
  LAYER M3 ;
        RECT 4.416 0.888 4.448 3.396 ;
  LAYER M3 ;
        RECT 4.48 0.888 4.512 3.396 ;
  LAYER M3 ;
        RECT 4.544 0.888 4.576 3.396 ;
  LAYER M3 ;
        RECT 4.608 0.888 4.64 3.396 ;
  LAYER M3 ;
        RECT 4.672 0.888 4.704 3.396 ;
  LAYER M3 ;
        RECT 4.736 0.888 4.768 3.396 ;
  LAYER M3 ;
        RECT 4.8 0.888 4.832 3.396 ;
  LAYER M3 ;
        RECT 4.864 0.888 4.896 3.396 ;
  LAYER M3 ;
        RECT 4.928 0.888 4.96 3.396 ;
  LAYER M3 ;
        RECT 4.992 0.888 5.024 3.396 ;
  LAYER M3 ;
        RECT 5.056 0.888 5.088 3.396 ;
  LAYER M3 ;
        RECT 5.12 0.888 5.152 3.396 ;
  LAYER M3 ;
        RECT 5.184 0.888 5.216 3.396 ;
  LAYER M3 ;
        RECT 5.248 0.888 5.28 3.396 ;
  LAYER M3 ;
        RECT 5.312 0.888 5.344 3.396 ;
  LAYER M3 ;
        RECT 5.376 0.888 5.408 3.396 ;
  LAYER M3 ;
        RECT 5.44 0.888 5.472 3.396 ;
  LAYER M3 ;
        RECT 5.504 0.888 5.536 3.396 ;
  LAYER M3 ;
        RECT 5.568 0.888 5.6 3.396 ;
  LAYER M3 ;
        RECT 5.664 0.888 5.696 3.396 ;
  LAYER M1 ;
        RECT 3.279 0.924 3.281 3.36 ;
  LAYER M1 ;
        RECT 3.359 0.924 3.361 3.36 ;
  LAYER M1 ;
        RECT 3.439 0.924 3.441 3.36 ;
  LAYER M1 ;
        RECT 3.519 0.924 3.521 3.36 ;
  LAYER M1 ;
        RECT 3.599 0.924 3.601 3.36 ;
  LAYER M1 ;
        RECT 3.679 0.924 3.681 3.36 ;
  LAYER M1 ;
        RECT 3.759 0.924 3.761 3.36 ;
  LAYER M1 ;
        RECT 3.839 0.924 3.841 3.36 ;
  LAYER M1 ;
        RECT 3.919 0.924 3.921 3.36 ;
  LAYER M1 ;
        RECT 3.999 0.924 4.001 3.36 ;
  LAYER M1 ;
        RECT 4.079 0.924 4.081 3.36 ;
  LAYER M1 ;
        RECT 4.159 0.924 4.161 3.36 ;
  LAYER M1 ;
        RECT 4.239 0.924 4.241 3.36 ;
  LAYER M1 ;
        RECT 4.319 0.924 4.321 3.36 ;
  LAYER M1 ;
        RECT 4.399 0.924 4.401 3.36 ;
  LAYER M1 ;
        RECT 4.479 0.924 4.481 3.36 ;
  LAYER M1 ;
        RECT 4.559 0.924 4.561 3.36 ;
  LAYER M1 ;
        RECT 4.639 0.924 4.641 3.36 ;
  LAYER M1 ;
        RECT 4.719 0.924 4.721 3.36 ;
  LAYER M1 ;
        RECT 4.799 0.924 4.801 3.36 ;
  LAYER M1 ;
        RECT 4.879 0.924 4.881 3.36 ;
  LAYER M1 ;
        RECT 4.959 0.924 4.961 3.36 ;
  LAYER M1 ;
        RECT 5.039 0.924 5.041 3.36 ;
  LAYER M1 ;
        RECT 5.119 0.924 5.121 3.36 ;
  LAYER M1 ;
        RECT 5.199 0.924 5.201 3.36 ;
  LAYER M1 ;
        RECT 5.279 0.924 5.281 3.36 ;
  LAYER M1 ;
        RECT 5.359 0.924 5.361 3.36 ;
  LAYER M1 ;
        RECT 5.439 0.924 5.441 3.36 ;
  LAYER M1 ;
        RECT 5.519 0.924 5.521 3.36 ;
  LAYER M1 ;
        RECT 5.599 0.924 5.601 3.36 ;
  LAYER M2 ;
        RECT 3.28 0.923 5.68 0.925 ;
  LAYER M2 ;
        RECT 3.28 1.007 5.68 1.009 ;
  LAYER M2 ;
        RECT 3.28 1.091 5.68 1.093 ;
  LAYER M2 ;
        RECT 3.28 1.175 5.68 1.177 ;
  LAYER M2 ;
        RECT 3.28 1.259 5.68 1.261 ;
  LAYER M2 ;
        RECT 3.28 1.343 5.68 1.345 ;
  LAYER M2 ;
        RECT 3.28 1.427 5.68 1.429 ;
  LAYER M2 ;
        RECT 3.28 1.511 5.68 1.513 ;
  LAYER M2 ;
        RECT 3.28 1.595 5.68 1.597 ;
  LAYER M2 ;
        RECT 3.28 1.679 5.68 1.681 ;
  LAYER M2 ;
        RECT 3.28 1.763 5.68 1.765 ;
  LAYER M2 ;
        RECT 3.28 1.847 5.68 1.849 ;
  LAYER M2 ;
        RECT 3.28 1.9305 5.68 1.9325 ;
  LAYER M2 ;
        RECT 3.28 2.015 5.68 2.017 ;
  LAYER M2 ;
        RECT 3.28 2.099 5.68 2.101 ;
  LAYER M2 ;
        RECT 3.28 2.183 5.68 2.185 ;
  LAYER M2 ;
        RECT 3.28 2.267 5.68 2.269 ;
  LAYER M2 ;
        RECT 3.28 2.351 5.68 2.353 ;
  LAYER M2 ;
        RECT 3.28 2.435 5.68 2.437 ;
  LAYER M2 ;
        RECT 3.28 2.519 5.68 2.521 ;
  LAYER M2 ;
        RECT 3.28 2.603 5.68 2.605 ;
  LAYER M2 ;
        RECT 3.28 2.687 5.68 2.689 ;
  LAYER M2 ;
        RECT 3.28 2.771 5.68 2.773 ;
  LAYER M2 ;
        RECT 3.28 2.855 5.68 2.857 ;
  LAYER M2 ;
        RECT 3.28 2.939 5.68 2.941 ;
  LAYER M2 ;
        RECT 3.28 3.023 5.68 3.025 ;
  LAYER M2 ;
        RECT 3.28 3.107 5.68 3.109 ;
  LAYER M2 ;
        RECT 3.28 3.191 5.68 3.193 ;
  LAYER M2 ;
        RECT 3.28 3.275 5.68 3.277 ;
  LAYER M1 ;
        RECT 3.264 3.828 3.296 6.336 ;
  LAYER M1 ;
        RECT 3.328 3.828 3.36 6.336 ;
  LAYER M1 ;
        RECT 3.392 3.828 3.424 6.336 ;
  LAYER M1 ;
        RECT 3.456 3.828 3.488 6.336 ;
  LAYER M1 ;
        RECT 3.52 3.828 3.552 6.336 ;
  LAYER M1 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M1 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M1 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M1 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M1 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M1 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M1 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M1 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M1 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M1 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M1 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M1 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M1 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M1 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M1 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M1 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M1 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M1 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M1 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M1 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M1 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M1 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M1 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M1 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M1 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M1 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M1 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M1 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M1 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M1 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M1 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M1 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M2 ;
        RECT 3.244 3.912 5.716 3.944 ;
  LAYER M2 ;
        RECT 3.244 3.976 5.716 4.008 ;
  LAYER M2 ;
        RECT 3.244 4.04 5.716 4.072 ;
  LAYER M2 ;
        RECT 3.244 4.104 5.716 4.136 ;
  LAYER M2 ;
        RECT 3.244 4.168 5.716 4.2 ;
  LAYER M2 ;
        RECT 3.244 4.232 5.716 4.264 ;
  LAYER M2 ;
        RECT 3.244 4.296 5.716 4.328 ;
  LAYER M2 ;
        RECT 3.244 4.36 5.716 4.392 ;
  LAYER M2 ;
        RECT 3.244 4.424 5.716 4.456 ;
  LAYER M2 ;
        RECT 3.244 4.488 5.716 4.52 ;
  LAYER M2 ;
        RECT 3.244 4.552 5.716 4.584 ;
  LAYER M2 ;
        RECT 3.244 4.616 5.716 4.648 ;
  LAYER M2 ;
        RECT 3.244 4.68 5.716 4.712 ;
  LAYER M2 ;
        RECT 3.244 4.744 5.716 4.776 ;
  LAYER M2 ;
        RECT 3.244 4.808 5.716 4.84 ;
  LAYER M2 ;
        RECT 3.244 4.872 5.716 4.904 ;
  LAYER M2 ;
        RECT 3.244 4.936 5.716 4.968 ;
  LAYER M2 ;
        RECT 3.244 5 5.716 5.032 ;
  LAYER M2 ;
        RECT 3.244 5.064 5.716 5.096 ;
  LAYER M2 ;
        RECT 3.244 5.128 5.716 5.16 ;
  LAYER M2 ;
        RECT 3.244 5.192 5.716 5.224 ;
  LAYER M2 ;
        RECT 3.244 5.256 5.716 5.288 ;
  LAYER M2 ;
        RECT 3.244 5.32 5.716 5.352 ;
  LAYER M2 ;
        RECT 3.244 5.384 5.716 5.416 ;
  LAYER M2 ;
        RECT 3.244 5.448 5.716 5.48 ;
  LAYER M2 ;
        RECT 3.244 5.512 5.716 5.544 ;
  LAYER M2 ;
        RECT 3.244 5.576 5.716 5.608 ;
  LAYER M2 ;
        RECT 3.244 5.64 5.716 5.672 ;
  LAYER M2 ;
        RECT 3.244 5.704 5.716 5.736 ;
  LAYER M2 ;
        RECT 3.244 5.768 5.716 5.8 ;
  LAYER M2 ;
        RECT 3.244 5.832 5.716 5.864 ;
  LAYER M2 ;
        RECT 3.244 5.896 5.716 5.928 ;
  LAYER M2 ;
        RECT 3.244 5.96 5.716 5.992 ;
  LAYER M2 ;
        RECT 3.244 6.024 5.716 6.056 ;
  LAYER M2 ;
        RECT 3.244 6.088 5.716 6.12 ;
  LAYER M2 ;
        RECT 3.244 6.152 5.716 6.184 ;
  LAYER M3 ;
        RECT 3.264 3.828 3.296 6.336 ;
  LAYER M3 ;
        RECT 3.328 3.828 3.36 6.336 ;
  LAYER M3 ;
        RECT 3.392 3.828 3.424 6.336 ;
  LAYER M3 ;
        RECT 3.456 3.828 3.488 6.336 ;
  LAYER M3 ;
        RECT 3.52 3.828 3.552 6.336 ;
  LAYER M3 ;
        RECT 3.584 3.828 3.616 6.336 ;
  LAYER M3 ;
        RECT 3.648 3.828 3.68 6.336 ;
  LAYER M3 ;
        RECT 3.712 3.828 3.744 6.336 ;
  LAYER M3 ;
        RECT 3.776 3.828 3.808 6.336 ;
  LAYER M3 ;
        RECT 3.84 3.828 3.872 6.336 ;
  LAYER M3 ;
        RECT 3.904 3.828 3.936 6.336 ;
  LAYER M3 ;
        RECT 3.968 3.828 4 6.336 ;
  LAYER M3 ;
        RECT 4.032 3.828 4.064 6.336 ;
  LAYER M3 ;
        RECT 4.096 3.828 4.128 6.336 ;
  LAYER M3 ;
        RECT 4.16 3.828 4.192 6.336 ;
  LAYER M3 ;
        RECT 4.224 3.828 4.256 6.336 ;
  LAYER M3 ;
        RECT 4.288 3.828 4.32 6.336 ;
  LAYER M3 ;
        RECT 4.352 3.828 4.384 6.336 ;
  LAYER M3 ;
        RECT 4.416 3.828 4.448 6.336 ;
  LAYER M3 ;
        RECT 4.48 3.828 4.512 6.336 ;
  LAYER M3 ;
        RECT 4.544 3.828 4.576 6.336 ;
  LAYER M3 ;
        RECT 4.608 3.828 4.64 6.336 ;
  LAYER M3 ;
        RECT 4.672 3.828 4.704 6.336 ;
  LAYER M3 ;
        RECT 4.736 3.828 4.768 6.336 ;
  LAYER M3 ;
        RECT 4.8 3.828 4.832 6.336 ;
  LAYER M3 ;
        RECT 4.864 3.828 4.896 6.336 ;
  LAYER M3 ;
        RECT 4.928 3.828 4.96 6.336 ;
  LAYER M3 ;
        RECT 4.992 3.828 5.024 6.336 ;
  LAYER M3 ;
        RECT 5.056 3.828 5.088 6.336 ;
  LAYER M3 ;
        RECT 5.12 3.828 5.152 6.336 ;
  LAYER M3 ;
        RECT 5.184 3.828 5.216 6.336 ;
  LAYER M3 ;
        RECT 5.248 3.828 5.28 6.336 ;
  LAYER M3 ;
        RECT 5.312 3.828 5.344 6.336 ;
  LAYER M3 ;
        RECT 5.376 3.828 5.408 6.336 ;
  LAYER M3 ;
        RECT 5.44 3.828 5.472 6.336 ;
  LAYER M3 ;
        RECT 5.504 3.828 5.536 6.336 ;
  LAYER M3 ;
        RECT 5.568 3.828 5.6 6.336 ;
  LAYER M3 ;
        RECT 5.664 3.828 5.696 6.336 ;
  LAYER M1 ;
        RECT 3.279 3.864 3.281 6.3 ;
  LAYER M1 ;
        RECT 3.359 3.864 3.361 6.3 ;
  LAYER M1 ;
        RECT 3.439 3.864 3.441 6.3 ;
  LAYER M1 ;
        RECT 3.519 3.864 3.521 6.3 ;
  LAYER M1 ;
        RECT 3.599 3.864 3.601 6.3 ;
  LAYER M1 ;
        RECT 3.679 3.864 3.681 6.3 ;
  LAYER M1 ;
        RECT 3.759 3.864 3.761 6.3 ;
  LAYER M1 ;
        RECT 3.839 3.864 3.841 6.3 ;
  LAYER M1 ;
        RECT 3.919 3.864 3.921 6.3 ;
  LAYER M1 ;
        RECT 3.999 3.864 4.001 6.3 ;
  LAYER M1 ;
        RECT 4.079 3.864 4.081 6.3 ;
  LAYER M1 ;
        RECT 4.159 3.864 4.161 6.3 ;
  LAYER M1 ;
        RECT 4.239 3.864 4.241 6.3 ;
  LAYER M1 ;
        RECT 4.319 3.864 4.321 6.3 ;
  LAYER M1 ;
        RECT 4.399 3.864 4.401 6.3 ;
  LAYER M1 ;
        RECT 4.479 3.864 4.481 6.3 ;
  LAYER M1 ;
        RECT 4.559 3.864 4.561 6.3 ;
  LAYER M1 ;
        RECT 4.639 3.864 4.641 6.3 ;
  LAYER M1 ;
        RECT 4.719 3.864 4.721 6.3 ;
  LAYER M1 ;
        RECT 4.799 3.864 4.801 6.3 ;
  LAYER M1 ;
        RECT 4.879 3.864 4.881 6.3 ;
  LAYER M1 ;
        RECT 4.959 3.864 4.961 6.3 ;
  LAYER M1 ;
        RECT 5.039 3.864 5.041 6.3 ;
  LAYER M1 ;
        RECT 5.119 3.864 5.121 6.3 ;
  LAYER M1 ;
        RECT 5.199 3.864 5.201 6.3 ;
  LAYER M1 ;
        RECT 5.279 3.864 5.281 6.3 ;
  LAYER M1 ;
        RECT 5.359 3.864 5.361 6.3 ;
  LAYER M1 ;
        RECT 5.439 3.864 5.441 6.3 ;
  LAYER M1 ;
        RECT 5.519 3.864 5.521 6.3 ;
  LAYER M1 ;
        RECT 5.599 3.864 5.601 6.3 ;
  LAYER M2 ;
        RECT 3.28 3.863 5.68 3.865 ;
  LAYER M2 ;
        RECT 3.28 3.947 5.68 3.949 ;
  LAYER M2 ;
        RECT 3.28 4.031 5.68 4.033 ;
  LAYER M2 ;
        RECT 3.28 4.115 5.68 4.117 ;
  LAYER M2 ;
        RECT 3.28 4.199 5.68 4.201 ;
  LAYER M2 ;
        RECT 3.28 4.283 5.68 4.285 ;
  LAYER M2 ;
        RECT 3.28 4.367 5.68 4.369 ;
  LAYER M2 ;
        RECT 3.28 4.451 5.68 4.453 ;
  LAYER M2 ;
        RECT 3.28 4.535 5.68 4.537 ;
  LAYER M2 ;
        RECT 3.28 4.619 5.68 4.621 ;
  LAYER M2 ;
        RECT 3.28 4.703 5.68 4.705 ;
  LAYER M2 ;
        RECT 3.28 4.787 5.68 4.789 ;
  LAYER M2 ;
        RECT 3.28 4.8705 5.68 4.8725 ;
  LAYER M2 ;
        RECT 3.28 4.955 5.68 4.957 ;
  LAYER M2 ;
        RECT 3.28 5.039 5.68 5.041 ;
  LAYER M2 ;
        RECT 3.28 5.123 5.68 5.125 ;
  LAYER M2 ;
        RECT 3.28 5.207 5.68 5.209 ;
  LAYER M2 ;
        RECT 3.28 5.291 5.68 5.293 ;
  LAYER M2 ;
        RECT 3.28 5.375 5.68 5.377 ;
  LAYER M2 ;
        RECT 3.28 5.459 5.68 5.461 ;
  LAYER M2 ;
        RECT 3.28 5.543 5.68 5.545 ;
  LAYER M2 ;
        RECT 3.28 5.627 5.68 5.629 ;
  LAYER M2 ;
        RECT 3.28 5.711 5.68 5.713 ;
  LAYER M2 ;
        RECT 3.28 5.795 5.68 5.797 ;
  LAYER M2 ;
        RECT 3.28 5.879 5.68 5.881 ;
  LAYER M2 ;
        RECT 3.28 5.963 5.68 5.965 ;
  LAYER M2 ;
        RECT 3.28 6.047 5.68 6.049 ;
  LAYER M2 ;
        RECT 3.28 6.131 5.68 6.133 ;
  LAYER M2 ;
        RECT 3.28 6.215 5.68 6.217 ;
  LAYER M1 ;
        RECT 3.264 6.768 3.296 9.276 ;
  LAYER M1 ;
        RECT 3.328 6.768 3.36 9.276 ;
  LAYER M1 ;
        RECT 3.392 6.768 3.424 9.276 ;
  LAYER M1 ;
        RECT 3.456 6.768 3.488 9.276 ;
  LAYER M1 ;
        RECT 3.52 6.768 3.552 9.276 ;
  LAYER M1 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M1 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M1 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M1 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M1 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M1 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M1 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M1 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M1 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M1 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M1 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M1 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M1 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M1 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M1 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M1 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M1 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M1 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M1 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M1 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M1 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M1 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M1 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M1 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M1 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M1 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M1 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M1 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M1 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M1 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M1 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M1 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M2 ;
        RECT 3.244 6.852 5.716 6.884 ;
  LAYER M2 ;
        RECT 3.244 6.916 5.716 6.948 ;
  LAYER M2 ;
        RECT 3.244 6.98 5.716 7.012 ;
  LAYER M2 ;
        RECT 3.244 7.044 5.716 7.076 ;
  LAYER M2 ;
        RECT 3.244 7.108 5.716 7.14 ;
  LAYER M2 ;
        RECT 3.244 7.172 5.716 7.204 ;
  LAYER M2 ;
        RECT 3.244 7.236 5.716 7.268 ;
  LAYER M2 ;
        RECT 3.244 7.3 5.716 7.332 ;
  LAYER M2 ;
        RECT 3.244 7.364 5.716 7.396 ;
  LAYER M2 ;
        RECT 3.244 7.428 5.716 7.46 ;
  LAYER M2 ;
        RECT 3.244 7.492 5.716 7.524 ;
  LAYER M2 ;
        RECT 3.244 7.556 5.716 7.588 ;
  LAYER M2 ;
        RECT 3.244 7.62 5.716 7.652 ;
  LAYER M2 ;
        RECT 3.244 7.684 5.716 7.716 ;
  LAYER M2 ;
        RECT 3.244 7.748 5.716 7.78 ;
  LAYER M2 ;
        RECT 3.244 7.812 5.716 7.844 ;
  LAYER M2 ;
        RECT 3.244 7.876 5.716 7.908 ;
  LAYER M2 ;
        RECT 3.244 7.94 5.716 7.972 ;
  LAYER M2 ;
        RECT 3.244 8.004 5.716 8.036 ;
  LAYER M2 ;
        RECT 3.244 8.068 5.716 8.1 ;
  LAYER M2 ;
        RECT 3.244 8.132 5.716 8.164 ;
  LAYER M2 ;
        RECT 3.244 8.196 5.716 8.228 ;
  LAYER M2 ;
        RECT 3.244 8.26 5.716 8.292 ;
  LAYER M2 ;
        RECT 3.244 8.324 5.716 8.356 ;
  LAYER M2 ;
        RECT 3.244 8.388 5.716 8.42 ;
  LAYER M2 ;
        RECT 3.244 8.452 5.716 8.484 ;
  LAYER M2 ;
        RECT 3.244 8.516 5.716 8.548 ;
  LAYER M2 ;
        RECT 3.244 8.58 5.716 8.612 ;
  LAYER M2 ;
        RECT 3.244 8.644 5.716 8.676 ;
  LAYER M2 ;
        RECT 3.244 8.708 5.716 8.74 ;
  LAYER M2 ;
        RECT 3.244 8.772 5.716 8.804 ;
  LAYER M2 ;
        RECT 3.244 8.836 5.716 8.868 ;
  LAYER M2 ;
        RECT 3.244 8.9 5.716 8.932 ;
  LAYER M2 ;
        RECT 3.244 8.964 5.716 8.996 ;
  LAYER M2 ;
        RECT 3.244 9.028 5.716 9.06 ;
  LAYER M2 ;
        RECT 3.244 9.092 5.716 9.124 ;
  LAYER M3 ;
        RECT 3.264 6.768 3.296 9.276 ;
  LAYER M3 ;
        RECT 3.328 6.768 3.36 9.276 ;
  LAYER M3 ;
        RECT 3.392 6.768 3.424 9.276 ;
  LAYER M3 ;
        RECT 3.456 6.768 3.488 9.276 ;
  LAYER M3 ;
        RECT 3.52 6.768 3.552 9.276 ;
  LAYER M3 ;
        RECT 3.584 6.768 3.616 9.276 ;
  LAYER M3 ;
        RECT 3.648 6.768 3.68 9.276 ;
  LAYER M3 ;
        RECT 3.712 6.768 3.744 9.276 ;
  LAYER M3 ;
        RECT 3.776 6.768 3.808 9.276 ;
  LAYER M3 ;
        RECT 3.84 6.768 3.872 9.276 ;
  LAYER M3 ;
        RECT 3.904 6.768 3.936 9.276 ;
  LAYER M3 ;
        RECT 3.968 6.768 4 9.276 ;
  LAYER M3 ;
        RECT 4.032 6.768 4.064 9.276 ;
  LAYER M3 ;
        RECT 4.096 6.768 4.128 9.276 ;
  LAYER M3 ;
        RECT 4.16 6.768 4.192 9.276 ;
  LAYER M3 ;
        RECT 4.224 6.768 4.256 9.276 ;
  LAYER M3 ;
        RECT 4.288 6.768 4.32 9.276 ;
  LAYER M3 ;
        RECT 4.352 6.768 4.384 9.276 ;
  LAYER M3 ;
        RECT 4.416 6.768 4.448 9.276 ;
  LAYER M3 ;
        RECT 4.48 6.768 4.512 9.276 ;
  LAYER M3 ;
        RECT 4.544 6.768 4.576 9.276 ;
  LAYER M3 ;
        RECT 4.608 6.768 4.64 9.276 ;
  LAYER M3 ;
        RECT 4.672 6.768 4.704 9.276 ;
  LAYER M3 ;
        RECT 4.736 6.768 4.768 9.276 ;
  LAYER M3 ;
        RECT 4.8 6.768 4.832 9.276 ;
  LAYER M3 ;
        RECT 4.864 6.768 4.896 9.276 ;
  LAYER M3 ;
        RECT 4.928 6.768 4.96 9.276 ;
  LAYER M3 ;
        RECT 4.992 6.768 5.024 9.276 ;
  LAYER M3 ;
        RECT 5.056 6.768 5.088 9.276 ;
  LAYER M3 ;
        RECT 5.12 6.768 5.152 9.276 ;
  LAYER M3 ;
        RECT 5.184 6.768 5.216 9.276 ;
  LAYER M3 ;
        RECT 5.248 6.768 5.28 9.276 ;
  LAYER M3 ;
        RECT 5.312 6.768 5.344 9.276 ;
  LAYER M3 ;
        RECT 5.376 6.768 5.408 9.276 ;
  LAYER M3 ;
        RECT 5.44 6.768 5.472 9.276 ;
  LAYER M3 ;
        RECT 5.504 6.768 5.536 9.276 ;
  LAYER M3 ;
        RECT 5.568 6.768 5.6 9.276 ;
  LAYER M3 ;
        RECT 5.664 6.768 5.696 9.276 ;
  LAYER M1 ;
        RECT 3.279 6.804 3.281 9.24 ;
  LAYER M1 ;
        RECT 3.359 6.804 3.361 9.24 ;
  LAYER M1 ;
        RECT 3.439 6.804 3.441 9.24 ;
  LAYER M1 ;
        RECT 3.519 6.804 3.521 9.24 ;
  LAYER M1 ;
        RECT 3.599 6.804 3.601 9.24 ;
  LAYER M1 ;
        RECT 3.679 6.804 3.681 9.24 ;
  LAYER M1 ;
        RECT 3.759 6.804 3.761 9.24 ;
  LAYER M1 ;
        RECT 3.839 6.804 3.841 9.24 ;
  LAYER M1 ;
        RECT 3.919 6.804 3.921 9.24 ;
  LAYER M1 ;
        RECT 3.999 6.804 4.001 9.24 ;
  LAYER M1 ;
        RECT 4.079 6.804 4.081 9.24 ;
  LAYER M1 ;
        RECT 4.159 6.804 4.161 9.24 ;
  LAYER M1 ;
        RECT 4.239 6.804 4.241 9.24 ;
  LAYER M1 ;
        RECT 4.319 6.804 4.321 9.24 ;
  LAYER M1 ;
        RECT 4.399 6.804 4.401 9.24 ;
  LAYER M1 ;
        RECT 4.479 6.804 4.481 9.24 ;
  LAYER M1 ;
        RECT 4.559 6.804 4.561 9.24 ;
  LAYER M1 ;
        RECT 4.639 6.804 4.641 9.24 ;
  LAYER M1 ;
        RECT 4.719 6.804 4.721 9.24 ;
  LAYER M1 ;
        RECT 4.799 6.804 4.801 9.24 ;
  LAYER M1 ;
        RECT 4.879 6.804 4.881 9.24 ;
  LAYER M1 ;
        RECT 4.959 6.804 4.961 9.24 ;
  LAYER M1 ;
        RECT 5.039 6.804 5.041 9.24 ;
  LAYER M1 ;
        RECT 5.119 6.804 5.121 9.24 ;
  LAYER M1 ;
        RECT 5.199 6.804 5.201 9.24 ;
  LAYER M1 ;
        RECT 5.279 6.804 5.281 9.24 ;
  LAYER M1 ;
        RECT 5.359 6.804 5.361 9.24 ;
  LAYER M1 ;
        RECT 5.439 6.804 5.441 9.24 ;
  LAYER M1 ;
        RECT 5.519 6.804 5.521 9.24 ;
  LAYER M1 ;
        RECT 5.599 6.804 5.601 9.24 ;
  LAYER M2 ;
        RECT 3.28 6.803 5.68 6.805 ;
  LAYER M2 ;
        RECT 3.28 6.887 5.68 6.889 ;
  LAYER M2 ;
        RECT 3.28 6.971 5.68 6.973 ;
  LAYER M2 ;
        RECT 3.28 7.055 5.68 7.057 ;
  LAYER M2 ;
        RECT 3.28 7.139 5.68 7.141 ;
  LAYER M2 ;
        RECT 3.28 7.223 5.68 7.225 ;
  LAYER M2 ;
        RECT 3.28 7.307 5.68 7.309 ;
  LAYER M2 ;
        RECT 3.28 7.391 5.68 7.393 ;
  LAYER M2 ;
        RECT 3.28 7.475 5.68 7.477 ;
  LAYER M2 ;
        RECT 3.28 7.559 5.68 7.561 ;
  LAYER M2 ;
        RECT 3.28 7.643 5.68 7.645 ;
  LAYER M2 ;
        RECT 3.28 7.727 5.68 7.729 ;
  LAYER M2 ;
        RECT 3.28 7.8105 5.68 7.8125 ;
  LAYER M2 ;
        RECT 3.28 7.895 5.68 7.897 ;
  LAYER M2 ;
        RECT 3.28 7.979 5.68 7.981 ;
  LAYER M2 ;
        RECT 3.28 8.063 5.68 8.065 ;
  LAYER M2 ;
        RECT 3.28 8.147 5.68 8.149 ;
  LAYER M2 ;
        RECT 3.28 8.231 5.68 8.233 ;
  LAYER M2 ;
        RECT 3.28 8.315 5.68 8.317 ;
  LAYER M2 ;
        RECT 3.28 8.399 5.68 8.401 ;
  LAYER M2 ;
        RECT 3.28 8.483 5.68 8.485 ;
  LAYER M2 ;
        RECT 3.28 8.567 5.68 8.569 ;
  LAYER M2 ;
        RECT 3.28 8.651 5.68 8.653 ;
  LAYER M2 ;
        RECT 3.28 8.735 5.68 8.737 ;
  LAYER M2 ;
        RECT 3.28 8.819 5.68 8.821 ;
  LAYER M2 ;
        RECT 3.28 8.903 5.68 8.905 ;
  LAYER M2 ;
        RECT 3.28 8.987 5.68 8.989 ;
  LAYER M2 ;
        RECT 3.28 9.071 5.68 9.073 ;
  LAYER M2 ;
        RECT 3.28 9.155 5.68 9.157 ;
  LAYER M1 ;
        RECT 3.264 9.708 3.296 12.216 ;
  LAYER M1 ;
        RECT 3.328 9.708 3.36 12.216 ;
  LAYER M1 ;
        RECT 3.392 9.708 3.424 12.216 ;
  LAYER M1 ;
        RECT 3.456 9.708 3.488 12.216 ;
  LAYER M1 ;
        RECT 3.52 9.708 3.552 12.216 ;
  LAYER M1 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M1 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M1 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M1 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M1 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M1 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M1 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M1 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M1 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M1 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M1 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M1 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M1 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M1 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M1 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M1 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M1 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M1 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M1 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M1 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M1 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M1 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M1 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M1 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M1 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M1 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M1 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M1 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M1 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M1 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M1 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M1 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M2 ;
        RECT 3.244 9.792 5.716 9.824 ;
  LAYER M2 ;
        RECT 3.244 9.856 5.716 9.888 ;
  LAYER M2 ;
        RECT 3.244 9.92 5.716 9.952 ;
  LAYER M2 ;
        RECT 3.244 9.984 5.716 10.016 ;
  LAYER M2 ;
        RECT 3.244 10.048 5.716 10.08 ;
  LAYER M2 ;
        RECT 3.244 10.112 5.716 10.144 ;
  LAYER M2 ;
        RECT 3.244 10.176 5.716 10.208 ;
  LAYER M2 ;
        RECT 3.244 10.24 5.716 10.272 ;
  LAYER M2 ;
        RECT 3.244 10.304 5.716 10.336 ;
  LAYER M2 ;
        RECT 3.244 10.368 5.716 10.4 ;
  LAYER M2 ;
        RECT 3.244 10.432 5.716 10.464 ;
  LAYER M2 ;
        RECT 3.244 10.496 5.716 10.528 ;
  LAYER M2 ;
        RECT 3.244 10.56 5.716 10.592 ;
  LAYER M2 ;
        RECT 3.244 10.624 5.716 10.656 ;
  LAYER M2 ;
        RECT 3.244 10.688 5.716 10.72 ;
  LAYER M2 ;
        RECT 3.244 10.752 5.716 10.784 ;
  LAYER M2 ;
        RECT 3.244 10.816 5.716 10.848 ;
  LAYER M2 ;
        RECT 3.244 10.88 5.716 10.912 ;
  LAYER M2 ;
        RECT 3.244 10.944 5.716 10.976 ;
  LAYER M2 ;
        RECT 3.244 11.008 5.716 11.04 ;
  LAYER M2 ;
        RECT 3.244 11.072 5.716 11.104 ;
  LAYER M2 ;
        RECT 3.244 11.136 5.716 11.168 ;
  LAYER M2 ;
        RECT 3.244 11.2 5.716 11.232 ;
  LAYER M2 ;
        RECT 3.244 11.264 5.716 11.296 ;
  LAYER M2 ;
        RECT 3.244 11.328 5.716 11.36 ;
  LAYER M2 ;
        RECT 3.244 11.392 5.716 11.424 ;
  LAYER M2 ;
        RECT 3.244 11.456 5.716 11.488 ;
  LAYER M2 ;
        RECT 3.244 11.52 5.716 11.552 ;
  LAYER M2 ;
        RECT 3.244 11.584 5.716 11.616 ;
  LAYER M2 ;
        RECT 3.244 11.648 5.716 11.68 ;
  LAYER M2 ;
        RECT 3.244 11.712 5.716 11.744 ;
  LAYER M2 ;
        RECT 3.244 11.776 5.716 11.808 ;
  LAYER M2 ;
        RECT 3.244 11.84 5.716 11.872 ;
  LAYER M2 ;
        RECT 3.244 11.904 5.716 11.936 ;
  LAYER M2 ;
        RECT 3.244 11.968 5.716 12 ;
  LAYER M2 ;
        RECT 3.244 12.032 5.716 12.064 ;
  LAYER M3 ;
        RECT 3.264 9.708 3.296 12.216 ;
  LAYER M3 ;
        RECT 3.328 9.708 3.36 12.216 ;
  LAYER M3 ;
        RECT 3.392 9.708 3.424 12.216 ;
  LAYER M3 ;
        RECT 3.456 9.708 3.488 12.216 ;
  LAYER M3 ;
        RECT 3.52 9.708 3.552 12.216 ;
  LAYER M3 ;
        RECT 3.584 9.708 3.616 12.216 ;
  LAYER M3 ;
        RECT 3.648 9.708 3.68 12.216 ;
  LAYER M3 ;
        RECT 3.712 9.708 3.744 12.216 ;
  LAYER M3 ;
        RECT 3.776 9.708 3.808 12.216 ;
  LAYER M3 ;
        RECT 3.84 9.708 3.872 12.216 ;
  LAYER M3 ;
        RECT 3.904 9.708 3.936 12.216 ;
  LAYER M3 ;
        RECT 3.968 9.708 4 12.216 ;
  LAYER M3 ;
        RECT 4.032 9.708 4.064 12.216 ;
  LAYER M3 ;
        RECT 4.096 9.708 4.128 12.216 ;
  LAYER M3 ;
        RECT 4.16 9.708 4.192 12.216 ;
  LAYER M3 ;
        RECT 4.224 9.708 4.256 12.216 ;
  LAYER M3 ;
        RECT 4.288 9.708 4.32 12.216 ;
  LAYER M3 ;
        RECT 4.352 9.708 4.384 12.216 ;
  LAYER M3 ;
        RECT 4.416 9.708 4.448 12.216 ;
  LAYER M3 ;
        RECT 4.48 9.708 4.512 12.216 ;
  LAYER M3 ;
        RECT 4.544 9.708 4.576 12.216 ;
  LAYER M3 ;
        RECT 4.608 9.708 4.64 12.216 ;
  LAYER M3 ;
        RECT 4.672 9.708 4.704 12.216 ;
  LAYER M3 ;
        RECT 4.736 9.708 4.768 12.216 ;
  LAYER M3 ;
        RECT 4.8 9.708 4.832 12.216 ;
  LAYER M3 ;
        RECT 4.864 9.708 4.896 12.216 ;
  LAYER M3 ;
        RECT 4.928 9.708 4.96 12.216 ;
  LAYER M3 ;
        RECT 4.992 9.708 5.024 12.216 ;
  LAYER M3 ;
        RECT 5.056 9.708 5.088 12.216 ;
  LAYER M3 ;
        RECT 5.12 9.708 5.152 12.216 ;
  LAYER M3 ;
        RECT 5.184 9.708 5.216 12.216 ;
  LAYER M3 ;
        RECT 5.248 9.708 5.28 12.216 ;
  LAYER M3 ;
        RECT 5.312 9.708 5.344 12.216 ;
  LAYER M3 ;
        RECT 5.376 9.708 5.408 12.216 ;
  LAYER M3 ;
        RECT 5.44 9.708 5.472 12.216 ;
  LAYER M3 ;
        RECT 5.504 9.708 5.536 12.216 ;
  LAYER M3 ;
        RECT 5.568 9.708 5.6 12.216 ;
  LAYER M3 ;
        RECT 5.664 9.708 5.696 12.216 ;
  LAYER M1 ;
        RECT 3.279 9.744 3.281 12.18 ;
  LAYER M1 ;
        RECT 3.359 9.744 3.361 12.18 ;
  LAYER M1 ;
        RECT 3.439 9.744 3.441 12.18 ;
  LAYER M1 ;
        RECT 3.519 9.744 3.521 12.18 ;
  LAYER M1 ;
        RECT 3.599 9.744 3.601 12.18 ;
  LAYER M1 ;
        RECT 3.679 9.744 3.681 12.18 ;
  LAYER M1 ;
        RECT 3.759 9.744 3.761 12.18 ;
  LAYER M1 ;
        RECT 3.839 9.744 3.841 12.18 ;
  LAYER M1 ;
        RECT 3.919 9.744 3.921 12.18 ;
  LAYER M1 ;
        RECT 3.999 9.744 4.001 12.18 ;
  LAYER M1 ;
        RECT 4.079 9.744 4.081 12.18 ;
  LAYER M1 ;
        RECT 4.159 9.744 4.161 12.18 ;
  LAYER M1 ;
        RECT 4.239 9.744 4.241 12.18 ;
  LAYER M1 ;
        RECT 4.319 9.744 4.321 12.18 ;
  LAYER M1 ;
        RECT 4.399 9.744 4.401 12.18 ;
  LAYER M1 ;
        RECT 4.479 9.744 4.481 12.18 ;
  LAYER M1 ;
        RECT 4.559 9.744 4.561 12.18 ;
  LAYER M1 ;
        RECT 4.639 9.744 4.641 12.18 ;
  LAYER M1 ;
        RECT 4.719 9.744 4.721 12.18 ;
  LAYER M1 ;
        RECT 4.799 9.744 4.801 12.18 ;
  LAYER M1 ;
        RECT 4.879 9.744 4.881 12.18 ;
  LAYER M1 ;
        RECT 4.959 9.744 4.961 12.18 ;
  LAYER M1 ;
        RECT 5.039 9.744 5.041 12.18 ;
  LAYER M1 ;
        RECT 5.119 9.744 5.121 12.18 ;
  LAYER M1 ;
        RECT 5.199 9.744 5.201 12.18 ;
  LAYER M1 ;
        RECT 5.279 9.744 5.281 12.18 ;
  LAYER M1 ;
        RECT 5.359 9.744 5.361 12.18 ;
  LAYER M1 ;
        RECT 5.439 9.744 5.441 12.18 ;
  LAYER M1 ;
        RECT 5.519 9.744 5.521 12.18 ;
  LAYER M1 ;
        RECT 5.599 9.744 5.601 12.18 ;
  LAYER M2 ;
        RECT 3.28 9.743 5.68 9.745 ;
  LAYER M2 ;
        RECT 3.28 9.827 5.68 9.829 ;
  LAYER M2 ;
        RECT 3.28 9.911 5.68 9.913 ;
  LAYER M2 ;
        RECT 3.28 9.995 5.68 9.997 ;
  LAYER M2 ;
        RECT 3.28 10.079 5.68 10.081 ;
  LAYER M2 ;
        RECT 3.28 10.163 5.68 10.165 ;
  LAYER M2 ;
        RECT 3.28 10.247 5.68 10.249 ;
  LAYER M2 ;
        RECT 3.28 10.331 5.68 10.333 ;
  LAYER M2 ;
        RECT 3.28 10.415 5.68 10.417 ;
  LAYER M2 ;
        RECT 3.28 10.499 5.68 10.501 ;
  LAYER M2 ;
        RECT 3.28 10.583 5.68 10.585 ;
  LAYER M2 ;
        RECT 3.28 10.667 5.68 10.669 ;
  LAYER M2 ;
        RECT 3.28 10.7505 5.68 10.7525 ;
  LAYER M2 ;
        RECT 3.28 10.835 5.68 10.837 ;
  LAYER M2 ;
        RECT 3.28 10.919 5.68 10.921 ;
  LAYER M2 ;
        RECT 3.28 11.003 5.68 11.005 ;
  LAYER M2 ;
        RECT 3.28 11.087 5.68 11.089 ;
  LAYER M2 ;
        RECT 3.28 11.171 5.68 11.173 ;
  LAYER M2 ;
        RECT 3.28 11.255 5.68 11.257 ;
  LAYER M2 ;
        RECT 3.28 11.339 5.68 11.341 ;
  LAYER M2 ;
        RECT 3.28 11.423 5.68 11.425 ;
  LAYER M2 ;
        RECT 3.28 11.507 5.68 11.509 ;
  LAYER M2 ;
        RECT 3.28 11.591 5.68 11.593 ;
  LAYER M2 ;
        RECT 3.28 11.675 5.68 11.677 ;
  LAYER M2 ;
        RECT 3.28 11.759 5.68 11.761 ;
  LAYER M2 ;
        RECT 3.28 11.843 5.68 11.845 ;
  LAYER M2 ;
        RECT 3.28 11.927 5.68 11.929 ;
  LAYER M2 ;
        RECT 3.28 12.011 5.68 12.013 ;
  LAYER M2 ;
        RECT 3.28 12.095 5.68 12.097 ;
  LAYER M1 ;
        RECT 3.264 12.648 3.296 15.156 ;
  LAYER M1 ;
        RECT 3.328 12.648 3.36 15.156 ;
  LAYER M1 ;
        RECT 3.392 12.648 3.424 15.156 ;
  LAYER M1 ;
        RECT 3.456 12.648 3.488 15.156 ;
  LAYER M1 ;
        RECT 3.52 12.648 3.552 15.156 ;
  LAYER M1 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M1 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M1 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M1 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M1 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M1 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M1 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M1 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M1 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M1 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M1 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M1 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M1 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M1 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M1 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M1 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M1 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M1 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M1 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M1 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M1 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M1 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M1 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M1 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M1 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M1 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M1 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M1 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M1 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M1 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M1 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M1 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M2 ;
        RECT 3.244 12.732 5.716 12.764 ;
  LAYER M2 ;
        RECT 3.244 12.796 5.716 12.828 ;
  LAYER M2 ;
        RECT 3.244 12.86 5.716 12.892 ;
  LAYER M2 ;
        RECT 3.244 12.924 5.716 12.956 ;
  LAYER M2 ;
        RECT 3.244 12.988 5.716 13.02 ;
  LAYER M2 ;
        RECT 3.244 13.052 5.716 13.084 ;
  LAYER M2 ;
        RECT 3.244 13.116 5.716 13.148 ;
  LAYER M2 ;
        RECT 3.244 13.18 5.716 13.212 ;
  LAYER M2 ;
        RECT 3.244 13.244 5.716 13.276 ;
  LAYER M2 ;
        RECT 3.244 13.308 5.716 13.34 ;
  LAYER M2 ;
        RECT 3.244 13.372 5.716 13.404 ;
  LAYER M2 ;
        RECT 3.244 13.436 5.716 13.468 ;
  LAYER M2 ;
        RECT 3.244 13.5 5.716 13.532 ;
  LAYER M2 ;
        RECT 3.244 13.564 5.716 13.596 ;
  LAYER M2 ;
        RECT 3.244 13.628 5.716 13.66 ;
  LAYER M2 ;
        RECT 3.244 13.692 5.716 13.724 ;
  LAYER M2 ;
        RECT 3.244 13.756 5.716 13.788 ;
  LAYER M2 ;
        RECT 3.244 13.82 5.716 13.852 ;
  LAYER M2 ;
        RECT 3.244 13.884 5.716 13.916 ;
  LAYER M2 ;
        RECT 3.244 13.948 5.716 13.98 ;
  LAYER M2 ;
        RECT 3.244 14.012 5.716 14.044 ;
  LAYER M2 ;
        RECT 3.244 14.076 5.716 14.108 ;
  LAYER M2 ;
        RECT 3.244 14.14 5.716 14.172 ;
  LAYER M2 ;
        RECT 3.244 14.204 5.716 14.236 ;
  LAYER M2 ;
        RECT 3.244 14.268 5.716 14.3 ;
  LAYER M2 ;
        RECT 3.244 14.332 5.716 14.364 ;
  LAYER M2 ;
        RECT 3.244 14.396 5.716 14.428 ;
  LAYER M2 ;
        RECT 3.244 14.46 5.716 14.492 ;
  LAYER M2 ;
        RECT 3.244 14.524 5.716 14.556 ;
  LAYER M2 ;
        RECT 3.244 14.588 5.716 14.62 ;
  LAYER M2 ;
        RECT 3.244 14.652 5.716 14.684 ;
  LAYER M2 ;
        RECT 3.244 14.716 5.716 14.748 ;
  LAYER M2 ;
        RECT 3.244 14.78 5.716 14.812 ;
  LAYER M2 ;
        RECT 3.244 14.844 5.716 14.876 ;
  LAYER M2 ;
        RECT 3.244 14.908 5.716 14.94 ;
  LAYER M2 ;
        RECT 3.244 14.972 5.716 15.004 ;
  LAYER M3 ;
        RECT 3.264 12.648 3.296 15.156 ;
  LAYER M3 ;
        RECT 3.328 12.648 3.36 15.156 ;
  LAYER M3 ;
        RECT 3.392 12.648 3.424 15.156 ;
  LAYER M3 ;
        RECT 3.456 12.648 3.488 15.156 ;
  LAYER M3 ;
        RECT 3.52 12.648 3.552 15.156 ;
  LAYER M3 ;
        RECT 3.584 12.648 3.616 15.156 ;
  LAYER M3 ;
        RECT 3.648 12.648 3.68 15.156 ;
  LAYER M3 ;
        RECT 3.712 12.648 3.744 15.156 ;
  LAYER M3 ;
        RECT 3.776 12.648 3.808 15.156 ;
  LAYER M3 ;
        RECT 3.84 12.648 3.872 15.156 ;
  LAYER M3 ;
        RECT 3.904 12.648 3.936 15.156 ;
  LAYER M3 ;
        RECT 3.968 12.648 4 15.156 ;
  LAYER M3 ;
        RECT 4.032 12.648 4.064 15.156 ;
  LAYER M3 ;
        RECT 4.096 12.648 4.128 15.156 ;
  LAYER M3 ;
        RECT 4.16 12.648 4.192 15.156 ;
  LAYER M3 ;
        RECT 4.224 12.648 4.256 15.156 ;
  LAYER M3 ;
        RECT 4.288 12.648 4.32 15.156 ;
  LAYER M3 ;
        RECT 4.352 12.648 4.384 15.156 ;
  LAYER M3 ;
        RECT 4.416 12.648 4.448 15.156 ;
  LAYER M3 ;
        RECT 4.48 12.648 4.512 15.156 ;
  LAYER M3 ;
        RECT 4.544 12.648 4.576 15.156 ;
  LAYER M3 ;
        RECT 4.608 12.648 4.64 15.156 ;
  LAYER M3 ;
        RECT 4.672 12.648 4.704 15.156 ;
  LAYER M3 ;
        RECT 4.736 12.648 4.768 15.156 ;
  LAYER M3 ;
        RECT 4.8 12.648 4.832 15.156 ;
  LAYER M3 ;
        RECT 4.864 12.648 4.896 15.156 ;
  LAYER M3 ;
        RECT 4.928 12.648 4.96 15.156 ;
  LAYER M3 ;
        RECT 4.992 12.648 5.024 15.156 ;
  LAYER M3 ;
        RECT 5.056 12.648 5.088 15.156 ;
  LAYER M3 ;
        RECT 5.12 12.648 5.152 15.156 ;
  LAYER M3 ;
        RECT 5.184 12.648 5.216 15.156 ;
  LAYER M3 ;
        RECT 5.248 12.648 5.28 15.156 ;
  LAYER M3 ;
        RECT 5.312 12.648 5.344 15.156 ;
  LAYER M3 ;
        RECT 5.376 12.648 5.408 15.156 ;
  LAYER M3 ;
        RECT 5.44 12.648 5.472 15.156 ;
  LAYER M3 ;
        RECT 5.504 12.648 5.536 15.156 ;
  LAYER M3 ;
        RECT 5.568 12.648 5.6 15.156 ;
  LAYER M3 ;
        RECT 5.664 12.648 5.696 15.156 ;
  LAYER M1 ;
        RECT 3.279 12.684 3.281 15.12 ;
  LAYER M1 ;
        RECT 3.359 12.684 3.361 15.12 ;
  LAYER M1 ;
        RECT 3.439 12.684 3.441 15.12 ;
  LAYER M1 ;
        RECT 3.519 12.684 3.521 15.12 ;
  LAYER M1 ;
        RECT 3.599 12.684 3.601 15.12 ;
  LAYER M1 ;
        RECT 3.679 12.684 3.681 15.12 ;
  LAYER M1 ;
        RECT 3.759 12.684 3.761 15.12 ;
  LAYER M1 ;
        RECT 3.839 12.684 3.841 15.12 ;
  LAYER M1 ;
        RECT 3.919 12.684 3.921 15.12 ;
  LAYER M1 ;
        RECT 3.999 12.684 4.001 15.12 ;
  LAYER M1 ;
        RECT 4.079 12.684 4.081 15.12 ;
  LAYER M1 ;
        RECT 4.159 12.684 4.161 15.12 ;
  LAYER M1 ;
        RECT 4.239 12.684 4.241 15.12 ;
  LAYER M1 ;
        RECT 4.319 12.684 4.321 15.12 ;
  LAYER M1 ;
        RECT 4.399 12.684 4.401 15.12 ;
  LAYER M1 ;
        RECT 4.479 12.684 4.481 15.12 ;
  LAYER M1 ;
        RECT 4.559 12.684 4.561 15.12 ;
  LAYER M1 ;
        RECT 4.639 12.684 4.641 15.12 ;
  LAYER M1 ;
        RECT 4.719 12.684 4.721 15.12 ;
  LAYER M1 ;
        RECT 4.799 12.684 4.801 15.12 ;
  LAYER M1 ;
        RECT 4.879 12.684 4.881 15.12 ;
  LAYER M1 ;
        RECT 4.959 12.684 4.961 15.12 ;
  LAYER M1 ;
        RECT 5.039 12.684 5.041 15.12 ;
  LAYER M1 ;
        RECT 5.119 12.684 5.121 15.12 ;
  LAYER M1 ;
        RECT 5.199 12.684 5.201 15.12 ;
  LAYER M1 ;
        RECT 5.279 12.684 5.281 15.12 ;
  LAYER M1 ;
        RECT 5.359 12.684 5.361 15.12 ;
  LAYER M1 ;
        RECT 5.439 12.684 5.441 15.12 ;
  LAYER M1 ;
        RECT 5.519 12.684 5.521 15.12 ;
  LAYER M1 ;
        RECT 5.599 12.684 5.601 15.12 ;
  LAYER M2 ;
        RECT 3.28 12.683 5.68 12.685 ;
  LAYER M2 ;
        RECT 3.28 12.767 5.68 12.769 ;
  LAYER M2 ;
        RECT 3.28 12.851 5.68 12.853 ;
  LAYER M2 ;
        RECT 3.28 12.935 5.68 12.937 ;
  LAYER M2 ;
        RECT 3.28 13.019 5.68 13.021 ;
  LAYER M2 ;
        RECT 3.28 13.103 5.68 13.105 ;
  LAYER M2 ;
        RECT 3.28 13.187 5.68 13.189 ;
  LAYER M2 ;
        RECT 3.28 13.271 5.68 13.273 ;
  LAYER M2 ;
        RECT 3.28 13.355 5.68 13.357 ;
  LAYER M2 ;
        RECT 3.28 13.439 5.68 13.441 ;
  LAYER M2 ;
        RECT 3.28 13.523 5.68 13.525 ;
  LAYER M2 ;
        RECT 3.28 13.607 5.68 13.609 ;
  LAYER M2 ;
        RECT 3.28 13.6905 5.68 13.6925 ;
  LAYER M2 ;
        RECT 3.28 13.775 5.68 13.777 ;
  LAYER M2 ;
        RECT 3.28 13.859 5.68 13.861 ;
  LAYER M2 ;
        RECT 3.28 13.943 5.68 13.945 ;
  LAYER M2 ;
        RECT 3.28 14.027 5.68 14.029 ;
  LAYER M2 ;
        RECT 3.28 14.111 5.68 14.113 ;
  LAYER M2 ;
        RECT 3.28 14.195 5.68 14.197 ;
  LAYER M2 ;
        RECT 3.28 14.279 5.68 14.281 ;
  LAYER M2 ;
        RECT 3.28 14.363 5.68 14.365 ;
  LAYER M2 ;
        RECT 3.28 14.447 5.68 14.449 ;
  LAYER M2 ;
        RECT 3.28 14.531 5.68 14.533 ;
  LAYER M2 ;
        RECT 3.28 14.615 5.68 14.617 ;
  LAYER M2 ;
        RECT 3.28 14.699 5.68 14.701 ;
  LAYER M2 ;
        RECT 3.28 14.783 5.68 14.785 ;
  LAYER M2 ;
        RECT 3.28 14.867 5.68 14.869 ;
  LAYER M2 ;
        RECT 3.28 14.951 5.68 14.953 ;
  LAYER M2 ;
        RECT 3.28 15.035 5.68 15.037 ;
  LAYER M1 ;
        RECT 3.264 15.588 3.296 18.096 ;
  LAYER M1 ;
        RECT 3.328 15.588 3.36 18.096 ;
  LAYER M1 ;
        RECT 3.392 15.588 3.424 18.096 ;
  LAYER M1 ;
        RECT 3.456 15.588 3.488 18.096 ;
  LAYER M1 ;
        RECT 3.52 15.588 3.552 18.096 ;
  LAYER M1 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M1 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M1 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M1 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M1 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M1 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M1 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M1 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M1 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M1 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M1 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M1 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M1 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M1 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M1 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M1 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M1 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M1 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M1 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M1 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M1 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M1 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M1 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M1 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M1 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M1 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M1 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M1 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M1 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M1 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M1 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M1 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M2 ;
        RECT 3.244 15.672 5.716 15.704 ;
  LAYER M2 ;
        RECT 3.244 15.736 5.716 15.768 ;
  LAYER M2 ;
        RECT 3.244 15.8 5.716 15.832 ;
  LAYER M2 ;
        RECT 3.244 15.864 5.716 15.896 ;
  LAYER M2 ;
        RECT 3.244 15.928 5.716 15.96 ;
  LAYER M2 ;
        RECT 3.244 15.992 5.716 16.024 ;
  LAYER M2 ;
        RECT 3.244 16.056 5.716 16.088 ;
  LAYER M2 ;
        RECT 3.244 16.12 5.716 16.152 ;
  LAYER M2 ;
        RECT 3.244 16.184 5.716 16.216 ;
  LAYER M2 ;
        RECT 3.244 16.248 5.716 16.28 ;
  LAYER M2 ;
        RECT 3.244 16.312 5.716 16.344 ;
  LAYER M2 ;
        RECT 3.244 16.376 5.716 16.408 ;
  LAYER M2 ;
        RECT 3.244 16.44 5.716 16.472 ;
  LAYER M2 ;
        RECT 3.244 16.504 5.716 16.536 ;
  LAYER M2 ;
        RECT 3.244 16.568 5.716 16.6 ;
  LAYER M2 ;
        RECT 3.244 16.632 5.716 16.664 ;
  LAYER M2 ;
        RECT 3.244 16.696 5.716 16.728 ;
  LAYER M2 ;
        RECT 3.244 16.76 5.716 16.792 ;
  LAYER M2 ;
        RECT 3.244 16.824 5.716 16.856 ;
  LAYER M2 ;
        RECT 3.244 16.888 5.716 16.92 ;
  LAYER M2 ;
        RECT 3.244 16.952 5.716 16.984 ;
  LAYER M2 ;
        RECT 3.244 17.016 5.716 17.048 ;
  LAYER M2 ;
        RECT 3.244 17.08 5.716 17.112 ;
  LAYER M2 ;
        RECT 3.244 17.144 5.716 17.176 ;
  LAYER M2 ;
        RECT 3.244 17.208 5.716 17.24 ;
  LAYER M2 ;
        RECT 3.244 17.272 5.716 17.304 ;
  LAYER M2 ;
        RECT 3.244 17.336 5.716 17.368 ;
  LAYER M2 ;
        RECT 3.244 17.4 5.716 17.432 ;
  LAYER M2 ;
        RECT 3.244 17.464 5.716 17.496 ;
  LAYER M2 ;
        RECT 3.244 17.528 5.716 17.56 ;
  LAYER M2 ;
        RECT 3.244 17.592 5.716 17.624 ;
  LAYER M2 ;
        RECT 3.244 17.656 5.716 17.688 ;
  LAYER M2 ;
        RECT 3.244 17.72 5.716 17.752 ;
  LAYER M2 ;
        RECT 3.244 17.784 5.716 17.816 ;
  LAYER M2 ;
        RECT 3.244 17.848 5.716 17.88 ;
  LAYER M2 ;
        RECT 3.244 17.912 5.716 17.944 ;
  LAYER M3 ;
        RECT 3.264 15.588 3.296 18.096 ;
  LAYER M3 ;
        RECT 3.328 15.588 3.36 18.096 ;
  LAYER M3 ;
        RECT 3.392 15.588 3.424 18.096 ;
  LAYER M3 ;
        RECT 3.456 15.588 3.488 18.096 ;
  LAYER M3 ;
        RECT 3.52 15.588 3.552 18.096 ;
  LAYER M3 ;
        RECT 3.584 15.588 3.616 18.096 ;
  LAYER M3 ;
        RECT 3.648 15.588 3.68 18.096 ;
  LAYER M3 ;
        RECT 3.712 15.588 3.744 18.096 ;
  LAYER M3 ;
        RECT 3.776 15.588 3.808 18.096 ;
  LAYER M3 ;
        RECT 3.84 15.588 3.872 18.096 ;
  LAYER M3 ;
        RECT 3.904 15.588 3.936 18.096 ;
  LAYER M3 ;
        RECT 3.968 15.588 4 18.096 ;
  LAYER M3 ;
        RECT 4.032 15.588 4.064 18.096 ;
  LAYER M3 ;
        RECT 4.096 15.588 4.128 18.096 ;
  LAYER M3 ;
        RECT 4.16 15.588 4.192 18.096 ;
  LAYER M3 ;
        RECT 4.224 15.588 4.256 18.096 ;
  LAYER M3 ;
        RECT 4.288 15.588 4.32 18.096 ;
  LAYER M3 ;
        RECT 4.352 15.588 4.384 18.096 ;
  LAYER M3 ;
        RECT 4.416 15.588 4.448 18.096 ;
  LAYER M3 ;
        RECT 4.48 15.588 4.512 18.096 ;
  LAYER M3 ;
        RECT 4.544 15.588 4.576 18.096 ;
  LAYER M3 ;
        RECT 4.608 15.588 4.64 18.096 ;
  LAYER M3 ;
        RECT 4.672 15.588 4.704 18.096 ;
  LAYER M3 ;
        RECT 4.736 15.588 4.768 18.096 ;
  LAYER M3 ;
        RECT 4.8 15.588 4.832 18.096 ;
  LAYER M3 ;
        RECT 4.864 15.588 4.896 18.096 ;
  LAYER M3 ;
        RECT 4.928 15.588 4.96 18.096 ;
  LAYER M3 ;
        RECT 4.992 15.588 5.024 18.096 ;
  LAYER M3 ;
        RECT 5.056 15.588 5.088 18.096 ;
  LAYER M3 ;
        RECT 5.12 15.588 5.152 18.096 ;
  LAYER M3 ;
        RECT 5.184 15.588 5.216 18.096 ;
  LAYER M3 ;
        RECT 5.248 15.588 5.28 18.096 ;
  LAYER M3 ;
        RECT 5.312 15.588 5.344 18.096 ;
  LAYER M3 ;
        RECT 5.376 15.588 5.408 18.096 ;
  LAYER M3 ;
        RECT 5.44 15.588 5.472 18.096 ;
  LAYER M3 ;
        RECT 5.504 15.588 5.536 18.096 ;
  LAYER M3 ;
        RECT 5.568 15.588 5.6 18.096 ;
  LAYER M3 ;
        RECT 5.664 15.588 5.696 18.096 ;
  LAYER M1 ;
        RECT 3.279 15.624 3.281 18.06 ;
  LAYER M1 ;
        RECT 3.359 15.624 3.361 18.06 ;
  LAYER M1 ;
        RECT 3.439 15.624 3.441 18.06 ;
  LAYER M1 ;
        RECT 3.519 15.624 3.521 18.06 ;
  LAYER M1 ;
        RECT 3.599 15.624 3.601 18.06 ;
  LAYER M1 ;
        RECT 3.679 15.624 3.681 18.06 ;
  LAYER M1 ;
        RECT 3.759 15.624 3.761 18.06 ;
  LAYER M1 ;
        RECT 3.839 15.624 3.841 18.06 ;
  LAYER M1 ;
        RECT 3.919 15.624 3.921 18.06 ;
  LAYER M1 ;
        RECT 3.999 15.624 4.001 18.06 ;
  LAYER M1 ;
        RECT 4.079 15.624 4.081 18.06 ;
  LAYER M1 ;
        RECT 4.159 15.624 4.161 18.06 ;
  LAYER M1 ;
        RECT 4.239 15.624 4.241 18.06 ;
  LAYER M1 ;
        RECT 4.319 15.624 4.321 18.06 ;
  LAYER M1 ;
        RECT 4.399 15.624 4.401 18.06 ;
  LAYER M1 ;
        RECT 4.479 15.624 4.481 18.06 ;
  LAYER M1 ;
        RECT 4.559 15.624 4.561 18.06 ;
  LAYER M1 ;
        RECT 4.639 15.624 4.641 18.06 ;
  LAYER M1 ;
        RECT 4.719 15.624 4.721 18.06 ;
  LAYER M1 ;
        RECT 4.799 15.624 4.801 18.06 ;
  LAYER M1 ;
        RECT 4.879 15.624 4.881 18.06 ;
  LAYER M1 ;
        RECT 4.959 15.624 4.961 18.06 ;
  LAYER M1 ;
        RECT 5.039 15.624 5.041 18.06 ;
  LAYER M1 ;
        RECT 5.119 15.624 5.121 18.06 ;
  LAYER M1 ;
        RECT 5.199 15.624 5.201 18.06 ;
  LAYER M1 ;
        RECT 5.279 15.624 5.281 18.06 ;
  LAYER M1 ;
        RECT 5.359 15.624 5.361 18.06 ;
  LAYER M1 ;
        RECT 5.439 15.624 5.441 18.06 ;
  LAYER M1 ;
        RECT 5.519 15.624 5.521 18.06 ;
  LAYER M1 ;
        RECT 5.599 15.624 5.601 18.06 ;
  LAYER M2 ;
        RECT 3.28 15.623 5.68 15.625 ;
  LAYER M2 ;
        RECT 3.28 15.707 5.68 15.709 ;
  LAYER M2 ;
        RECT 3.28 15.791 5.68 15.793 ;
  LAYER M2 ;
        RECT 3.28 15.875 5.68 15.877 ;
  LAYER M2 ;
        RECT 3.28 15.959 5.68 15.961 ;
  LAYER M2 ;
        RECT 3.28 16.043 5.68 16.045 ;
  LAYER M2 ;
        RECT 3.28 16.127 5.68 16.129 ;
  LAYER M2 ;
        RECT 3.28 16.211 5.68 16.213 ;
  LAYER M2 ;
        RECT 3.28 16.295 5.68 16.297 ;
  LAYER M2 ;
        RECT 3.28 16.379 5.68 16.381 ;
  LAYER M2 ;
        RECT 3.28 16.463 5.68 16.465 ;
  LAYER M2 ;
        RECT 3.28 16.547 5.68 16.549 ;
  LAYER M2 ;
        RECT 3.28 16.6305 5.68 16.6325 ;
  LAYER M2 ;
        RECT 3.28 16.715 5.68 16.717 ;
  LAYER M2 ;
        RECT 3.28 16.799 5.68 16.801 ;
  LAYER M2 ;
        RECT 3.28 16.883 5.68 16.885 ;
  LAYER M2 ;
        RECT 3.28 16.967 5.68 16.969 ;
  LAYER M2 ;
        RECT 3.28 17.051 5.68 17.053 ;
  LAYER M2 ;
        RECT 3.28 17.135 5.68 17.137 ;
  LAYER M2 ;
        RECT 3.28 17.219 5.68 17.221 ;
  LAYER M2 ;
        RECT 3.28 17.303 5.68 17.305 ;
  LAYER M2 ;
        RECT 3.28 17.387 5.68 17.389 ;
  LAYER M2 ;
        RECT 3.28 17.471 5.68 17.473 ;
  LAYER M2 ;
        RECT 3.28 17.555 5.68 17.557 ;
  LAYER M2 ;
        RECT 3.28 17.639 5.68 17.641 ;
  LAYER M2 ;
        RECT 3.28 17.723 5.68 17.725 ;
  LAYER M2 ;
        RECT 3.28 17.807 5.68 17.809 ;
  LAYER M2 ;
        RECT 3.28 17.891 5.68 17.893 ;
  LAYER M2 ;
        RECT 3.28 17.975 5.68 17.977 ;
  LAYER M1 ;
        RECT 6.144 0.888 6.176 3.396 ;
  LAYER M1 ;
        RECT 6.208 0.888 6.24 3.396 ;
  LAYER M1 ;
        RECT 6.272 0.888 6.304 3.396 ;
  LAYER M1 ;
        RECT 6.336 0.888 6.368 3.396 ;
  LAYER M1 ;
        RECT 6.4 0.888 6.432 3.396 ;
  LAYER M1 ;
        RECT 6.464 0.888 6.496 3.396 ;
  LAYER M1 ;
        RECT 6.528 0.888 6.56 3.396 ;
  LAYER M1 ;
        RECT 6.592 0.888 6.624 3.396 ;
  LAYER M1 ;
        RECT 6.656 0.888 6.688 3.396 ;
  LAYER M1 ;
        RECT 6.72 0.888 6.752 3.396 ;
  LAYER M1 ;
        RECT 6.784 0.888 6.816 3.396 ;
  LAYER M1 ;
        RECT 6.848 0.888 6.88 3.396 ;
  LAYER M1 ;
        RECT 6.912 0.888 6.944 3.396 ;
  LAYER M1 ;
        RECT 6.976 0.888 7.008 3.396 ;
  LAYER M1 ;
        RECT 7.04 0.888 7.072 3.396 ;
  LAYER M1 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M1 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M1 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M1 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M1 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M1 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M1 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M1 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M1 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M1 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M1 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M1 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M1 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M1 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M1 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M1 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M1 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M1 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M1 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M1 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M1 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M1 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M2 ;
        RECT 6.124 0.972 8.596 1.004 ;
  LAYER M2 ;
        RECT 6.124 1.036 8.596 1.068 ;
  LAYER M2 ;
        RECT 6.124 1.1 8.596 1.132 ;
  LAYER M2 ;
        RECT 6.124 1.164 8.596 1.196 ;
  LAYER M2 ;
        RECT 6.124 1.228 8.596 1.26 ;
  LAYER M2 ;
        RECT 6.124 1.292 8.596 1.324 ;
  LAYER M2 ;
        RECT 6.124 1.356 8.596 1.388 ;
  LAYER M2 ;
        RECT 6.124 1.42 8.596 1.452 ;
  LAYER M2 ;
        RECT 6.124 1.484 8.596 1.516 ;
  LAYER M2 ;
        RECT 6.124 1.548 8.596 1.58 ;
  LAYER M2 ;
        RECT 6.124 1.612 8.596 1.644 ;
  LAYER M2 ;
        RECT 6.124 1.676 8.596 1.708 ;
  LAYER M2 ;
        RECT 6.124 1.74 8.596 1.772 ;
  LAYER M2 ;
        RECT 6.124 1.804 8.596 1.836 ;
  LAYER M2 ;
        RECT 6.124 1.868 8.596 1.9 ;
  LAYER M2 ;
        RECT 6.124 1.932 8.596 1.964 ;
  LAYER M2 ;
        RECT 6.124 1.996 8.596 2.028 ;
  LAYER M2 ;
        RECT 6.124 2.06 8.596 2.092 ;
  LAYER M2 ;
        RECT 6.124 2.124 8.596 2.156 ;
  LAYER M2 ;
        RECT 6.124 2.188 8.596 2.22 ;
  LAYER M2 ;
        RECT 6.124 2.252 8.596 2.284 ;
  LAYER M2 ;
        RECT 6.124 2.316 8.596 2.348 ;
  LAYER M2 ;
        RECT 6.124 2.38 8.596 2.412 ;
  LAYER M2 ;
        RECT 6.124 2.444 8.596 2.476 ;
  LAYER M2 ;
        RECT 6.124 2.508 8.596 2.54 ;
  LAYER M2 ;
        RECT 6.124 2.572 8.596 2.604 ;
  LAYER M2 ;
        RECT 6.124 2.636 8.596 2.668 ;
  LAYER M2 ;
        RECT 6.124 2.7 8.596 2.732 ;
  LAYER M2 ;
        RECT 6.124 2.764 8.596 2.796 ;
  LAYER M2 ;
        RECT 6.124 2.828 8.596 2.86 ;
  LAYER M2 ;
        RECT 6.124 2.892 8.596 2.924 ;
  LAYER M2 ;
        RECT 6.124 2.956 8.596 2.988 ;
  LAYER M2 ;
        RECT 6.124 3.02 8.596 3.052 ;
  LAYER M2 ;
        RECT 6.124 3.084 8.596 3.116 ;
  LAYER M2 ;
        RECT 6.124 3.148 8.596 3.18 ;
  LAYER M2 ;
        RECT 6.124 3.212 8.596 3.244 ;
  LAYER M3 ;
        RECT 6.144 0.888 6.176 3.396 ;
  LAYER M3 ;
        RECT 6.208 0.888 6.24 3.396 ;
  LAYER M3 ;
        RECT 6.272 0.888 6.304 3.396 ;
  LAYER M3 ;
        RECT 6.336 0.888 6.368 3.396 ;
  LAYER M3 ;
        RECT 6.4 0.888 6.432 3.396 ;
  LAYER M3 ;
        RECT 6.464 0.888 6.496 3.396 ;
  LAYER M3 ;
        RECT 6.528 0.888 6.56 3.396 ;
  LAYER M3 ;
        RECT 6.592 0.888 6.624 3.396 ;
  LAYER M3 ;
        RECT 6.656 0.888 6.688 3.396 ;
  LAYER M3 ;
        RECT 6.72 0.888 6.752 3.396 ;
  LAYER M3 ;
        RECT 6.784 0.888 6.816 3.396 ;
  LAYER M3 ;
        RECT 6.848 0.888 6.88 3.396 ;
  LAYER M3 ;
        RECT 6.912 0.888 6.944 3.396 ;
  LAYER M3 ;
        RECT 6.976 0.888 7.008 3.396 ;
  LAYER M3 ;
        RECT 7.04 0.888 7.072 3.396 ;
  LAYER M3 ;
        RECT 7.104 0.888 7.136 3.396 ;
  LAYER M3 ;
        RECT 7.168 0.888 7.2 3.396 ;
  LAYER M3 ;
        RECT 7.232 0.888 7.264 3.396 ;
  LAYER M3 ;
        RECT 7.296 0.888 7.328 3.396 ;
  LAYER M3 ;
        RECT 7.36 0.888 7.392 3.396 ;
  LAYER M3 ;
        RECT 7.424 0.888 7.456 3.396 ;
  LAYER M3 ;
        RECT 7.488 0.888 7.52 3.396 ;
  LAYER M3 ;
        RECT 7.552 0.888 7.584 3.396 ;
  LAYER M3 ;
        RECT 7.616 0.888 7.648 3.396 ;
  LAYER M3 ;
        RECT 7.68 0.888 7.712 3.396 ;
  LAYER M3 ;
        RECT 7.744 0.888 7.776 3.396 ;
  LAYER M3 ;
        RECT 7.808 0.888 7.84 3.396 ;
  LAYER M3 ;
        RECT 7.872 0.888 7.904 3.396 ;
  LAYER M3 ;
        RECT 7.936 0.888 7.968 3.396 ;
  LAYER M3 ;
        RECT 8 0.888 8.032 3.396 ;
  LAYER M3 ;
        RECT 8.064 0.888 8.096 3.396 ;
  LAYER M3 ;
        RECT 8.128 0.888 8.16 3.396 ;
  LAYER M3 ;
        RECT 8.192 0.888 8.224 3.396 ;
  LAYER M3 ;
        RECT 8.256 0.888 8.288 3.396 ;
  LAYER M3 ;
        RECT 8.32 0.888 8.352 3.396 ;
  LAYER M3 ;
        RECT 8.384 0.888 8.416 3.396 ;
  LAYER M3 ;
        RECT 8.448 0.888 8.48 3.396 ;
  LAYER M3 ;
        RECT 8.544 0.888 8.576 3.396 ;
  LAYER M1 ;
        RECT 6.159 0.924 6.161 3.36 ;
  LAYER M1 ;
        RECT 6.239 0.924 6.241 3.36 ;
  LAYER M1 ;
        RECT 6.319 0.924 6.321 3.36 ;
  LAYER M1 ;
        RECT 6.399 0.924 6.401 3.36 ;
  LAYER M1 ;
        RECT 6.479 0.924 6.481 3.36 ;
  LAYER M1 ;
        RECT 6.559 0.924 6.561 3.36 ;
  LAYER M1 ;
        RECT 6.639 0.924 6.641 3.36 ;
  LAYER M1 ;
        RECT 6.719 0.924 6.721 3.36 ;
  LAYER M1 ;
        RECT 6.799 0.924 6.801 3.36 ;
  LAYER M1 ;
        RECT 6.879 0.924 6.881 3.36 ;
  LAYER M1 ;
        RECT 6.959 0.924 6.961 3.36 ;
  LAYER M1 ;
        RECT 7.039 0.924 7.041 3.36 ;
  LAYER M1 ;
        RECT 7.119 0.924 7.121 3.36 ;
  LAYER M1 ;
        RECT 7.199 0.924 7.201 3.36 ;
  LAYER M1 ;
        RECT 7.279 0.924 7.281 3.36 ;
  LAYER M1 ;
        RECT 7.359 0.924 7.361 3.36 ;
  LAYER M1 ;
        RECT 7.439 0.924 7.441 3.36 ;
  LAYER M1 ;
        RECT 7.519 0.924 7.521 3.36 ;
  LAYER M1 ;
        RECT 7.599 0.924 7.601 3.36 ;
  LAYER M1 ;
        RECT 7.679 0.924 7.681 3.36 ;
  LAYER M1 ;
        RECT 7.759 0.924 7.761 3.36 ;
  LAYER M1 ;
        RECT 7.839 0.924 7.841 3.36 ;
  LAYER M1 ;
        RECT 7.919 0.924 7.921 3.36 ;
  LAYER M1 ;
        RECT 7.999 0.924 8.001 3.36 ;
  LAYER M1 ;
        RECT 8.079 0.924 8.081 3.36 ;
  LAYER M1 ;
        RECT 8.159 0.924 8.161 3.36 ;
  LAYER M1 ;
        RECT 8.239 0.924 8.241 3.36 ;
  LAYER M1 ;
        RECT 8.319 0.924 8.321 3.36 ;
  LAYER M1 ;
        RECT 8.399 0.924 8.401 3.36 ;
  LAYER M1 ;
        RECT 8.479 0.924 8.481 3.36 ;
  LAYER M2 ;
        RECT 6.16 0.923 8.56 0.925 ;
  LAYER M2 ;
        RECT 6.16 1.007 8.56 1.009 ;
  LAYER M2 ;
        RECT 6.16 1.091 8.56 1.093 ;
  LAYER M2 ;
        RECT 6.16 1.175 8.56 1.177 ;
  LAYER M2 ;
        RECT 6.16 1.259 8.56 1.261 ;
  LAYER M2 ;
        RECT 6.16 1.343 8.56 1.345 ;
  LAYER M2 ;
        RECT 6.16 1.427 8.56 1.429 ;
  LAYER M2 ;
        RECT 6.16 1.511 8.56 1.513 ;
  LAYER M2 ;
        RECT 6.16 1.595 8.56 1.597 ;
  LAYER M2 ;
        RECT 6.16 1.679 8.56 1.681 ;
  LAYER M2 ;
        RECT 6.16 1.763 8.56 1.765 ;
  LAYER M2 ;
        RECT 6.16 1.847 8.56 1.849 ;
  LAYER M2 ;
        RECT 6.16 1.9305 8.56 1.9325 ;
  LAYER M2 ;
        RECT 6.16 2.015 8.56 2.017 ;
  LAYER M2 ;
        RECT 6.16 2.099 8.56 2.101 ;
  LAYER M2 ;
        RECT 6.16 2.183 8.56 2.185 ;
  LAYER M2 ;
        RECT 6.16 2.267 8.56 2.269 ;
  LAYER M2 ;
        RECT 6.16 2.351 8.56 2.353 ;
  LAYER M2 ;
        RECT 6.16 2.435 8.56 2.437 ;
  LAYER M2 ;
        RECT 6.16 2.519 8.56 2.521 ;
  LAYER M2 ;
        RECT 6.16 2.603 8.56 2.605 ;
  LAYER M2 ;
        RECT 6.16 2.687 8.56 2.689 ;
  LAYER M2 ;
        RECT 6.16 2.771 8.56 2.773 ;
  LAYER M2 ;
        RECT 6.16 2.855 8.56 2.857 ;
  LAYER M2 ;
        RECT 6.16 2.939 8.56 2.941 ;
  LAYER M2 ;
        RECT 6.16 3.023 8.56 3.025 ;
  LAYER M2 ;
        RECT 6.16 3.107 8.56 3.109 ;
  LAYER M2 ;
        RECT 6.16 3.191 8.56 3.193 ;
  LAYER M2 ;
        RECT 6.16 3.275 8.56 3.277 ;
  LAYER M1 ;
        RECT 6.144 3.828 6.176 6.336 ;
  LAYER M1 ;
        RECT 6.208 3.828 6.24 6.336 ;
  LAYER M1 ;
        RECT 6.272 3.828 6.304 6.336 ;
  LAYER M1 ;
        RECT 6.336 3.828 6.368 6.336 ;
  LAYER M1 ;
        RECT 6.4 3.828 6.432 6.336 ;
  LAYER M1 ;
        RECT 6.464 3.828 6.496 6.336 ;
  LAYER M1 ;
        RECT 6.528 3.828 6.56 6.336 ;
  LAYER M1 ;
        RECT 6.592 3.828 6.624 6.336 ;
  LAYER M1 ;
        RECT 6.656 3.828 6.688 6.336 ;
  LAYER M1 ;
        RECT 6.72 3.828 6.752 6.336 ;
  LAYER M1 ;
        RECT 6.784 3.828 6.816 6.336 ;
  LAYER M1 ;
        RECT 6.848 3.828 6.88 6.336 ;
  LAYER M1 ;
        RECT 6.912 3.828 6.944 6.336 ;
  LAYER M1 ;
        RECT 6.976 3.828 7.008 6.336 ;
  LAYER M1 ;
        RECT 7.04 3.828 7.072 6.336 ;
  LAYER M1 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M1 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M1 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M1 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M1 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M1 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M1 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M1 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M1 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M1 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M1 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M1 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M1 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M1 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M1 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M1 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M1 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M1 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M1 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M1 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M1 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M1 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M2 ;
        RECT 6.124 3.912 8.596 3.944 ;
  LAYER M2 ;
        RECT 6.124 3.976 8.596 4.008 ;
  LAYER M2 ;
        RECT 6.124 4.04 8.596 4.072 ;
  LAYER M2 ;
        RECT 6.124 4.104 8.596 4.136 ;
  LAYER M2 ;
        RECT 6.124 4.168 8.596 4.2 ;
  LAYER M2 ;
        RECT 6.124 4.232 8.596 4.264 ;
  LAYER M2 ;
        RECT 6.124 4.296 8.596 4.328 ;
  LAYER M2 ;
        RECT 6.124 4.36 8.596 4.392 ;
  LAYER M2 ;
        RECT 6.124 4.424 8.596 4.456 ;
  LAYER M2 ;
        RECT 6.124 4.488 8.596 4.52 ;
  LAYER M2 ;
        RECT 6.124 4.552 8.596 4.584 ;
  LAYER M2 ;
        RECT 6.124 4.616 8.596 4.648 ;
  LAYER M2 ;
        RECT 6.124 4.68 8.596 4.712 ;
  LAYER M2 ;
        RECT 6.124 4.744 8.596 4.776 ;
  LAYER M2 ;
        RECT 6.124 4.808 8.596 4.84 ;
  LAYER M2 ;
        RECT 6.124 4.872 8.596 4.904 ;
  LAYER M2 ;
        RECT 6.124 4.936 8.596 4.968 ;
  LAYER M2 ;
        RECT 6.124 5 8.596 5.032 ;
  LAYER M2 ;
        RECT 6.124 5.064 8.596 5.096 ;
  LAYER M2 ;
        RECT 6.124 5.128 8.596 5.16 ;
  LAYER M2 ;
        RECT 6.124 5.192 8.596 5.224 ;
  LAYER M2 ;
        RECT 6.124 5.256 8.596 5.288 ;
  LAYER M2 ;
        RECT 6.124 5.32 8.596 5.352 ;
  LAYER M2 ;
        RECT 6.124 5.384 8.596 5.416 ;
  LAYER M2 ;
        RECT 6.124 5.448 8.596 5.48 ;
  LAYER M2 ;
        RECT 6.124 5.512 8.596 5.544 ;
  LAYER M2 ;
        RECT 6.124 5.576 8.596 5.608 ;
  LAYER M2 ;
        RECT 6.124 5.64 8.596 5.672 ;
  LAYER M2 ;
        RECT 6.124 5.704 8.596 5.736 ;
  LAYER M2 ;
        RECT 6.124 5.768 8.596 5.8 ;
  LAYER M2 ;
        RECT 6.124 5.832 8.596 5.864 ;
  LAYER M2 ;
        RECT 6.124 5.896 8.596 5.928 ;
  LAYER M2 ;
        RECT 6.124 5.96 8.596 5.992 ;
  LAYER M2 ;
        RECT 6.124 6.024 8.596 6.056 ;
  LAYER M2 ;
        RECT 6.124 6.088 8.596 6.12 ;
  LAYER M2 ;
        RECT 6.124 6.152 8.596 6.184 ;
  LAYER M3 ;
        RECT 6.144 3.828 6.176 6.336 ;
  LAYER M3 ;
        RECT 6.208 3.828 6.24 6.336 ;
  LAYER M3 ;
        RECT 6.272 3.828 6.304 6.336 ;
  LAYER M3 ;
        RECT 6.336 3.828 6.368 6.336 ;
  LAYER M3 ;
        RECT 6.4 3.828 6.432 6.336 ;
  LAYER M3 ;
        RECT 6.464 3.828 6.496 6.336 ;
  LAYER M3 ;
        RECT 6.528 3.828 6.56 6.336 ;
  LAYER M3 ;
        RECT 6.592 3.828 6.624 6.336 ;
  LAYER M3 ;
        RECT 6.656 3.828 6.688 6.336 ;
  LAYER M3 ;
        RECT 6.72 3.828 6.752 6.336 ;
  LAYER M3 ;
        RECT 6.784 3.828 6.816 6.336 ;
  LAYER M3 ;
        RECT 6.848 3.828 6.88 6.336 ;
  LAYER M3 ;
        RECT 6.912 3.828 6.944 6.336 ;
  LAYER M3 ;
        RECT 6.976 3.828 7.008 6.336 ;
  LAYER M3 ;
        RECT 7.04 3.828 7.072 6.336 ;
  LAYER M3 ;
        RECT 7.104 3.828 7.136 6.336 ;
  LAYER M3 ;
        RECT 7.168 3.828 7.2 6.336 ;
  LAYER M3 ;
        RECT 7.232 3.828 7.264 6.336 ;
  LAYER M3 ;
        RECT 7.296 3.828 7.328 6.336 ;
  LAYER M3 ;
        RECT 7.36 3.828 7.392 6.336 ;
  LAYER M3 ;
        RECT 7.424 3.828 7.456 6.336 ;
  LAYER M3 ;
        RECT 7.488 3.828 7.52 6.336 ;
  LAYER M3 ;
        RECT 7.552 3.828 7.584 6.336 ;
  LAYER M3 ;
        RECT 7.616 3.828 7.648 6.336 ;
  LAYER M3 ;
        RECT 7.68 3.828 7.712 6.336 ;
  LAYER M3 ;
        RECT 7.744 3.828 7.776 6.336 ;
  LAYER M3 ;
        RECT 7.808 3.828 7.84 6.336 ;
  LAYER M3 ;
        RECT 7.872 3.828 7.904 6.336 ;
  LAYER M3 ;
        RECT 7.936 3.828 7.968 6.336 ;
  LAYER M3 ;
        RECT 8 3.828 8.032 6.336 ;
  LAYER M3 ;
        RECT 8.064 3.828 8.096 6.336 ;
  LAYER M3 ;
        RECT 8.128 3.828 8.16 6.336 ;
  LAYER M3 ;
        RECT 8.192 3.828 8.224 6.336 ;
  LAYER M3 ;
        RECT 8.256 3.828 8.288 6.336 ;
  LAYER M3 ;
        RECT 8.32 3.828 8.352 6.336 ;
  LAYER M3 ;
        RECT 8.384 3.828 8.416 6.336 ;
  LAYER M3 ;
        RECT 8.448 3.828 8.48 6.336 ;
  LAYER M3 ;
        RECT 8.544 3.828 8.576 6.336 ;
  LAYER M1 ;
        RECT 6.159 3.864 6.161 6.3 ;
  LAYER M1 ;
        RECT 6.239 3.864 6.241 6.3 ;
  LAYER M1 ;
        RECT 6.319 3.864 6.321 6.3 ;
  LAYER M1 ;
        RECT 6.399 3.864 6.401 6.3 ;
  LAYER M1 ;
        RECT 6.479 3.864 6.481 6.3 ;
  LAYER M1 ;
        RECT 6.559 3.864 6.561 6.3 ;
  LAYER M1 ;
        RECT 6.639 3.864 6.641 6.3 ;
  LAYER M1 ;
        RECT 6.719 3.864 6.721 6.3 ;
  LAYER M1 ;
        RECT 6.799 3.864 6.801 6.3 ;
  LAYER M1 ;
        RECT 6.879 3.864 6.881 6.3 ;
  LAYER M1 ;
        RECT 6.959 3.864 6.961 6.3 ;
  LAYER M1 ;
        RECT 7.039 3.864 7.041 6.3 ;
  LAYER M1 ;
        RECT 7.119 3.864 7.121 6.3 ;
  LAYER M1 ;
        RECT 7.199 3.864 7.201 6.3 ;
  LAYER M1 ;
        RECT 7.279 3.864 7.281 6.3 ;
  LAYER M1 ;
        RECT 7.359 3.864 7.361 6.3 ;
  LAYER M1 ;
        RECT 7.439 3.864 7.441 6.3 ;
  LAYER M1 ;
        RECT 7.519 3.864 7.521 6.3 ;
  LAYER M1 ;
        RECT 7.599 3.864 7.601 6.3 ;
  LAYER M1 ;
        RECT 7.679 3.864 7.681 6.3 ;
  LAYER M1 ;
        RECT 7.759 3.864 7.761 6.3 ;
  LAYER M1 ;
        RECT 7.839 3.864 7.841 6.3 ;
  LAYER M1 ;
        RECT 7.919 3.864 7.921 6.3 ;
  LAYER M1 ;
        RECT 7.999 3.864 8.001 6.3 ;
  LAYER M1 ;
        RECT 8.079 3.864 8.081 6.3 ;
  LAYER M1 ;
        RECT 8.159 3.864 8.161 6.3 ;
  LAYER M1 ;
        RECT 8.239 3.864 8.241 6.3 ;
  LAYER M1 ;
        RECT 8.319 3.864 8.321 6.3 ;
  LAYER M1 ;
        RECT 8.399 3.864 8.401 6.3 ;
  LAYER M1 ;
        RECT 8.479 3.864 8.481 6.3 ;
  LAYER M2 ;
        RECT 6.16 3.863 8.56 3.865 ;
  LAYER M2 ;
        RECT 6.16 3.947 8.56 3.949 ;
  LAYER M2 ;
        RECT 6.16 4.031 8.56 4.033 ;
  LAYER M2 ;
        RECT 6.16 4.115 8.56 4.117 ;
  LAYER M2 ;
        RECT 6.16 4.199 8.56 4.201 ;
  LAYER M2 ;
        RECT 6.16 4.283 8.56 4.285 ;
  LAYER M2 ;
        RECT 6.16 4.367 8.56 4.369 ;
  LAYER M2 ;
        RECT 6.16 4.451 8.56 4.453 ;
  LAYER M2 ;
        RECT 6.16 4.535 8.56 4.537 ;
  LAYER M2 ;
        RECT 6.16 4.619 8.56 4.621 ;
  LAYER M2 ;
        RECT 6.16 4.703 8.56 4.705 ;
  LAYER M2 ;
        RECT 6.16 4.787 8.56 4.789 ;
  LAYER M2 ;
        RECT 6.16 4.8705 8.56 4.8725 ;
  LAYER M2 ;
        RECT 6.16 4.955 8.56 4.957 ;
  LAYER M2 ;
        RECT 6.16 5.039 8.56 5.041 ;
  LAYER M2 ;
        RECT 6.16 5.123 8.56 5.125 ;
  LAYER M2 ;
        RECT 6.16 5.207 8.56 5.209 ;
  LAYER M2 ;
        RECT 6.16 5.291 8.56 5.293 ;
  LAYER M2 ;
        RECT 6.16 5.375 8.56 5.377 ;
  LAYER M2 ;
        RECT 6.16 5.459 8.56 5.461 ;
  LAYER M2 ;
        RECT 6.16 5.543 8.56 5.545 ;
  LAYER M2 ;
        RECT 6.16 5.627 8.56 5.629 ;
  LAYER M2 ;
        RECT 6.16 5.711 8.56 5.713 ;
  LAYER M2 ;
        RECT 6.16 5.795 8.56 5.797 ;
  LAYER M2 ;
        RECT 6.16 5.879 8.56 5.881 ;
  LAYER M2 ;
        RECT 6.16 5.963 8.56 5.965 ;
  LAYER M2 ;
        RECT 6.16 6.047 8.56 6.049 ;
  LAYER M2 ;
        RECT 6.16 6.131 8.56 6.133 ;
  LAYER M2 ;
        RECT 6.16 6.215 8.56 6.217 ;
  LAYER M1 ;
        RECT 6.144 6.768 6.176 9.276 ;
  LAYER M1 ;
        RECT 6.208 6.768 6.24 9.276 ;
  LAYER M1 ;
        RECT 6.272 6.768 6.304 9.276 ;
  LAYER M1 ;
        RECT 6.336 6.768 6.368 9.276 ;
  LAYER M1 ;
        RECT 6.4 6.768 6.432 9.276 ;
  LAYER M1 ;
        RECT 6.464 6.768 6.496 9.276 ;
  LAYER M1 ;
        RECT 6.528 6.768 6.56 9.276 ;
  LAYER M1 ;
        RECT 6.592 6.768 6.624 9.276 ;
  LAYER M1 ;
        RECT 6.656 6.768 6.688 9.276 ;
  LAYER M1 ;
        RECT 6.72 6.768 6.752 9.276 ;
  LAYER M1 ;
        RECT 6.784 6.768 6.816 9.276 ;
  LAYER M1 ;
        RECT 6.848 6.768 6.88 9.276 ;
  LAYER M1 ;
        RECT 6.912 6.768 6.944 9.276 ;
  LAYER M1 ;
        RECT 6.976 6.768 7.008 9.276 ;
  LAYER M1 ;
        RECT 7.04 6.768 7.072 9.276 ;
  LAYER M1 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M1 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M1 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M1 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M1 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M1 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M1 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M1 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M1 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M1 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M1 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M1 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M1 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M1 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M1 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M1 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M1 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M1 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M1 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M1 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M1 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M1 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M2 ;
        RECT 6.124 6.852 8.596 6.884 ;
  LAYER M2 ;
        RECT 6.124 6.916 8.596 6.948 ;
  LAYER M2 ;
        RECT 6.124 6.98 8.596 7.012 ;
  LAYER M2 ;
        RECT 6.124 7.044 8.596 7.076 ;
  LAYER M2 ;
        RECT 6.124 7.108 8.596 7.14 ;
  LAYER M2 ;
        RECT 6.124 7.172 8.596 7.204 ;
  LAYER M2 ;
        RECT 6.124 7.236 8.596 7.268 ;
  LAYER M2 ;
        RECT 6.124 7.3 8.596 7.332 ;
  LAYER M2 ;
        RECT 6.124 7.364 8.596 7.396 ;
  LAYER M2 ;
        RECT 6.124 7.428 8.596 7.46 ;
  LAYER M2 ;
        RECT 6.124 7.492 8.596 7.524 ;
  LAYER M2 ;
        RECT 6.124 7.556 8.596 7.588 ;
  LAYER M2 ;
        RECT 6.124 7.62 8.596 7.652 ;
  LAYER M2 ;
        RECT 6.124 7.684 8.596 7.716 ;
  LAYER M2 ;
        RECT 6.124 7.748 8.596 7.78 ;
  LAYER M2 ;
        RECT 6.124 7.812 8.596 7.844 ;
  LAYER M2 ;
        RECT 6.124 7.876 8.596 7.908 ;
  LAYER M2 ;
        RECT 6.124 7.94 8.596 7.972 ;
  LAYER M2 ;
        RECT 6.124 8.004 8.596 8.036 ;
  LAYER M2 ;
        RECT 6.124 8.068 8.596 8.1 ;
  LAYER M2 ;
        RECT 6.124 8.132 8.596 8.164 ;
  LAYER M2 ;
        RECT 6.124 8.196 8.596 8.228 ;
  LAYER M2 ;
        RECT 6.124 8.26 8.596 8.292 ;
  LAYER M2 ;
        RECT 6.124 8.324 8.596 8.356 ;
  LAYER M2 ;
        RECT 6.124 8.388 8.596 8.42 ;
  LAYER M2 ;
        RECT 6.124 8.452 8.596 8.484 ;
  LAYER M2 ;
        RECT 6.124 8.516 8.596 8.548 ;
  LAYER M2 ;
        RECT 6.124 8.58 8.596 8.612 ;
  LAYER M2 ;
        RECT 6.124 8.644 8.596 8.676 ;
  LAYER M2 ;
        RECT 6.124 8.708 8.596 8.74 ;
  LAYER M2 ;
        RECT 6.124 8.772 8.596 8.804 ;
  LAYER M2 ;
        RECT 6.124 8.836 8.596 8.868 ;
  LAYER M2 ;
        RECT 6.124 8.9 8.596 8.932 ;
  LAYER M2 ;
        RECT 6.124 8.964 8.596 8.996 ;
  LAYER M2 ;
        RECT 6.124 9.028 8.596 9.06 ;
  LAYER M2 ;
        RECT 6.124 9.092 8.596 9.124 ;
  LAYER M3 ;
        RECT 6.144 6.768 6.176 9.276 ;
  LAYER M3 ;
        RECT 6.208 6.768 6.24 9.276 ;
  LAYER M3 ;
        RECT 6.272 6.768 6.304 9.276 ;
  LAYER M3 ;
        RECT 6.336 6.768 6.368 9.276 ;
  LAYER M3 ;
        RECT 6.4 6.768 6.432 9.276 ;
  LAYER M3 ;
        RECT 6.464 6.768 6.496 9.276 ;
  LAYER M3 ;
        RECT 6.528 6.768 6.56 9.276 ;
  LAYER M3 ;
        RECT 6.592 6.768 6.624 9.276 ;
  LAYER M3 ;
        RECT 6.656 6.768 6.688 9.276 ;
  LAYER M3 ;
        RECT 6.72 6.768 6.752 9.276 ;
  LAYER M3 ;
        RECT 6.784 6.768 6.816 9.276 ;
  LAYER M3 ;
        RECT 6.848 6.768 6.88 9.276 ;
  LAYER M3 ;
        RECT 6.912 6.768 6.944 9.276 ;
  LAYER M3 ;
        RECT 6.976 6.768 7.008 9.276 ;
  LAYER M3 ;
        RECT 7.04 6.768 7.072 9.276 ;
  LAYER M3 ;
        RECT 7.104 6.768 7.136 9.276 ;
  LAYER M3 ;
        RECT 7.168 6.768 7.2 9.276 ;
  LAYER M3 ;
        RECT 7.232 6.768 7.264 9.276 ;
  LAYER M3 ;
        RECT 7.296 6.768 7.328 9.276 ;
  LAYER M3 ;
        RECT 7.36 6.768 7.392 9.276 ;
  LAYER M3 ;
        RECT 7.424 6.768 7.456 9.276 ;
  LAYER M3 ;
        RECT 7.488 6.768 7.52 9.276 ;
  LAYER M3 ;
        RECT 7.552 6.768 7.584 9.276 ;
  LAYER M3 ;
        RECT 7.616 6.768 7.648 9.276 ;
  LAYER M3 ;
        RECT 7.68 6.768 7.712 9.276 ;
  LAYER M3 ;
        RECT 7.744 6.768 7.776 9.276 ;
  LAYER M3 ;
        RECT 7.808 6.768 7.84 9.276 ;
  LAYER M3 ;
        RECT 7.872 6.768 7.904 9.276 ;
  LAYER M3 ;
        RECT 7.936 6.768 7.968 9.276 ;
  LAYER M3 ;
        RECT 8 6.768 8.032 9.276 ;
  LAYER M3 ;
        RECT 8.064 6.768 8.096 9.276 ;
  LAYER M3 ;
        RECT 8.128 6.768 8.16 9.276 ;
  LAYER M3 ;
        RECT 8.192 6.768 8.224 9.276 ;
  LAYER M3 ;
        RECT 8.256 6.768 8.288 9.276 ;
  LAYER M3 ;
        RECT 8.32 6.768 8.352 9.276 ;
  LAYER M3 ;
        RECT 8.384 6.768 8.416 9.276 ;
  LAYER M3 ;
        RECT 8.448 6.768 8.48 9.276 ;
  LAYER M3 ;
        RECT 8.544 6.768 8.576 9.276 ;
  LAYER M1 ;
        RECT 6.159 6.804 6.161 9.24 ;
  LAYER M1 ;
        RECT 6.239 6.804 6.241 9.24 ;
  LAYER M1 ;
        RECT 6.319 6.804 6.321 9.24 ;
  LAYER M1 ;
        RECT 6.399 6.804 6.401 9.24 ;
  LAYER M1 ;
        RECT 6.479 6.804 6.481 9.24 ;
  LAYER M1 ;
        RECT 6.559 6.804 6.561 9.24 ;
  LAYER M1 ;
        RECT 6.639 6.804 6.641 9.24 ;
  LAYER M1 ;
        RECT 6.719 6.804 6.721 9.24 ;
  LAYER M1 ;
        RECT 6.799 6.804 6.801 9.24 ;
  LAYER M1 ;
        RECT 6.879 6.804 6.881 9.24 ;
  LAYER M1 ;
        RECT 6.959 6.804 6.961 9.24 ;
  LAYER M1 ;
        RECT 7.039 6.804 7.041 9.24 ;
  LAYER M1 ;
        RECT 7.119 6.804 7.121 9.24 ;
  LAYER M1 ;
        RECT 7.199 6.804 7.201 9.24 ;
  LAYER M1 ;
        RECT 7.279 6.804 7.281 9.24 ;
  LAYER M1 ;
        RECT 7.359 6.804 7.361 9.24 ;
  LAYER M1 ;
        RECT 7.439 6.804 7.441 9.24 ;
  LAYER M1 ;
        RECT 7.519 6.804 7.521 9.24 ;
  LAYER M1 ;
        RECT 7.599 6.804 7.601 9.24 ;
  LAYER M1 ;
        RECT 7.679 6.804 7.681 9.24 ;
  LAYER M1 ;
        RECT 7.759 6.804 7.761 9.24 ;
  LAYER M1 ;
        RECT 7.839 6.804 7.841 9.24 ;
  LAYER M1 ;
        RECT 7.919 6.804 7.921 9.24 ;
  LAYER M1 ;
        RECT 7.999 6.804 8.001 9.24 ;
  LAYER M1 ;
        RECT 8.079 6.804 8.081 9.24 ;
  LAYER M1 ;
        RECT 8.159 6.804 8.161 9.24 ;
  LAYER M1 ;
        RECT 8.239 6.804 8.241 9.24 ;
  LAYER M1 ;
        RECT 8.319 6.804 8.321 9.24 ;
  LAYER M1 ;
        RECT 8.399 6.804 8.401 9.24 ;
  LAYER M1 ;
        RECT 8.479 6.804 8.481 9.24 ;
  LAYER M2 ;
        RECT 6.16 6.803 8.56 6.805 ;
  LAYER M2 ;
        RECT 6.16 6.887 8.56 6.889 ;
  LAYER M2 ;
        RECT 6.16 6.971 8.56 6.973 ;
  LAYER M2 ;
        RECT 6.16 7.055 8.56 7.057 ;
  LAYER M2 ;
        RECT 6.16 7.139 8.56 7.141 ;
  LAYER M2 ;
        RECT 6.16 7.223 8.56 7.225 ;
  LAYER M2 ;
        RECT 6.16 7.307 8.56 7.309 ;
  LAYER M2 ;
        RECT 6.16 7.391 8.56 7.393 ;
  LAYER M2 ;
        RECT 6.16 7.475 8.56 7.477 ;
  LAYER M2 ;
        RECT 6.16 7.559 8.56 7.561 ;
  LAYER M2 ;
        RECT 6.16 7.643 8.56 7.645 ;
  LAYER M2 ;
        RECT 6.16 7.727 8.56 7.729 ;
  LAYER M2 ;
        RECT 6.16 7.8105 8.56 7.8125 ;
  LAYER M2 ;
        RECT 6.16 7.895 8.56 7.897 ;
  LAYER M2 ;
        RECT 6.16 7.979 8.56 7.981 ;
  LAYER M2 ;
        RECT 6.16 8.063 8.56 8.065 ;
  LAYER M2 ;
        RECT 6.16 8.147 8.56 8.149 ;
  LAYER M2 ;
        RECT 6.16 8.231 8.56 8.233 ;
  LAYER M2 ;
        RECT 6.16 8.315 8.56 8.317 ;
  LAYER M2 ;
        RECT 6.16 8.399 8.56 8.401 ;
  LAYER M2 ;
        RECT 6.16 8.483 8.56 8.485 ;
  LAYER M2 ;
        RECT 6.16 8.567 8.56 8.569 ;
  LAYER M2 ;
        RECT 6.16 8.651 8.56 8.653 ;
  LAYER M2 ;
        RECT 6.16 8.735 8.56 8.737 ;
  LAYER M2 ;
        RECT 6.16 8.819 8.56 8.821 ;
  LAYER M2 ;
        RECT 6.16 8.903 8.56 8.905 ;
  LAYER M2 ;
        RECT 6.16 8.987 8.56 8.989 ;
  LAYER M2 ;
        RECT 6.16 9.071 8.56 9.073 ;
  LAYER M2 ;
        RECT 6.16 9.155 8.56 9.157 ;
  LAYER M1 ;
        RECT 6.144 9.708 6.176 12.216 ;
  LAYER M1 ;
        RECT 6.208 9.708 6.24 12.216 ;
  LAYER M1 ;
        RECT 6.272 9.708 6.304 12.216 ;
  LAYER M1 ;
        RECT 6.336 9.708 6.368 12.216 ;
  LAYER M1 ;
        RECT 6.4 9.708 6.432 12.216 ;
  LAYER M1 ;
        RECT 6.464 9.708 6.496 12.216 ;
  LAYER M1 ;
        RECT 6.528 9.708 6.56 12.216 ;
  LAYER M1 ;
        RECT 6.592 9.708 6.624 12.216 ;
  LAYER M1 ;
        RECT 6.656 9.708 6.688 12.216 ;
  LAYER M1 ;
        RECT 6.72 9.708 6.752 12.216 ;
  LAYER M1 ;
        RECT 6.784 9.708 6.816 12.216 ;
  LAYER M1 ;
        RECT 6.848 9.708 6.88 12.216 ;
  LAYER M1 ;
        RECT 6.912 9.708 6.944 12.216 ;
  LAYER M1 ;
        RECT 6.976 9.708 7.008 12.216 ;
  LAYER M1 ;
        RECT 7.04 9.708 7.072 12.216 ;
  LAYER M1 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M1 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M1 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M1 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M1 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M1 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M1 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M1 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M1 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M1 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M1 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M1 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M1 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M1 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M1 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M1 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M1 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M1 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M1 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M1 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M1 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M1 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M2 ;
        RECT 6.124 9.792 8.596 9.824 ;
  LAYER M2 ;
        RECT 6.124 9.856 8.596 9.888 ;
  LAYER M2 ;
        RECT 6.124 9.92 8.596 9.952 ;
  LAYER M2 ;
        RECT 6.124 9.984 8.596 10.016 ;
  LAYER M2 ;
        RECT 6.124 10.048 8.596 10.08 ;
  LAYER M2 ;
        RECT 6.124 10.112 8.596 10.144 ;
  LAYER M2 ;
        RECT 6.124 10.176 8.596 10.208 ;
  LAYER M2 ;
        RECT 6.124 10.24 8.596 10.272 ;
  LAYER M2 ;
        RECT 6.124 10.304 8.596 10.336 ;
  LAYER M2 ;
        RECT 6.124 10.368 8.596 10.4 ;
  LAYER M2 ;
        RECT 6.124 10.432 8.596 10.464 ;
  LAYER M2 ;
        RECT 6.124 10.496 8.596 10.528 ;
  LAYER M2 ;
        RECT 6.124 10.56 8.596 10.592 ;
  LAYER M2 ;
        RECT 6.124 10.624 8.596 10.656 ;
  LAYER M2 ;
        RECT 6.124 10.688 8.596 10.72 ;
  LAYER M2 ;
        RECT 6.124 10.752 8.596 10.784 ;
  LAYER M2 ;
        RECT 6.124 10.816 8.596 10.848 ;
  LAYER M2 ;
        RECT 6.124 10.88 8.596 10.912 ;
  LAYER M2 ;
        RECT 6.124 10.944 8.596 10.976 ;
  LAYER M2 ;
        RECT 6.124 11.008 8.596 11.04 ;
  LAYER M2 ;
        RECT 6.124 11.072 8.596 11.104 ;
  LAYER M2 ;
        RECT 6.124 11.136 8.596 11.168 ;
  LAYER M2 ;
        RECT 6.124 11.2 8.596 11.232 ;
  LAYER M2 ;
        RECT 6.124 11.264 8.596 11.296 ;
  LAYER M2 ;
        RECT 6.124 11.328 8.596 11.36 ;
  LAYER M2 ;
        RECT 6.124 11.392 8.596 11.424 ;
  LAYER M2 ;
        RECT 6.124 11.456 8.596 11.488 ;
  LAYER M2 ;
        RECT 6.124 11.52 8.596 11.552 ;
  LAYER M2 ;
        RECT 6.124 11.584 8.596 11.616 ;
  LAYER M2 ;
        RECT 6.124 11.648 8.596 11.68 ;
  LAYER M2 ;
        RECT 6.124 11.712 8.596 11.744 ;
  LAYER M2 ;
        RECT 6.124 11.776 8.596 11.808 ;
  LAYER M2 ;
        RECT 6.124 11.84 8.596 11.872 ;
  LAYER M2 ;
        RECT 6.124 11.904 8.596 11.936 ;
  LAYER M2 ;
        RECT 6.124 11.968 8.596 12 ;
  LAYER M2 ;
        RECT 6.124 12.032 8.596 12.064 ;
  LAYER M3 ;
        RECT 6.144 9.708 6.176 12.216 ;
  LAYER M3 ;
        RECT 6.208 9.708 6.24 12.216 ;
  LAYER M3 ;
        RECT 6.272 9.708 6.304 12.216 ;
  LAYER M3 ;
        RECT 6.336 9.708 6.368 12.216 ;
  LAYER M3 ;
        RECT 6.4 9.708 6.432 12.216 ;
  LAYER M3 ;
        RECT 6.464 9.708 6.496 12.216 ;
  LAYER M3 ;
        RECT 6.528 9.708 6.56 12.216 ;
  LAYER M3 ;
        RECT 6.592 9.708 6.624 12.216 ;
  LAYER M3 ;
        RECT 6.656 9.708 6.688 12.216 ;
  LAYER M3 ;
        RECT 6.72 9.708 6.752 12.216 ;
  LAYER M3 ;
        RECT 6.784 9.708 6.816 12.216 ;
  LAYER M3 ;
        RECT 6.848 9.708 6.88 12.216 ;
  LAYER M3 ;
        RECT 6.912 9.708 6.944 12.216 ;
  LAYER M3 ;
        RECT 6.976 9.708 7.008 12.216 ;
  LAYER M3 ;
        RECT 7.04 9.708 7.072 12.216 ;
  LAYER M3 ;
        RECT 7.104 9.708 7.136 12.216 ;
  LAYER M3 ;
        RECT 7.168 9.708 7.2 12.216 ;
  LAYER M3 ;
        RECT 7.232 9.708 7.264 12.216 ;
  LAYER M3 ;
        RECT 7.296 9.708 7.328 12.216 ;
  LAYER M3 ;
        RECT 7.36 9.708 7.392 12.216 ;
  LAYER M3 ;
        RECT 7.424 9.708 7.456 12.216 ;
  LAYER M3 ;
        RECT 7.488 9.708 7.52 12.216 ;
  LAYER M3 ;
        RECT 7.552 9.708 7.584 12.216 ;
  LAYER M3 ;
        RECT 7.616 9.708 7.648 12.216 ;
  LAYER M3 ;
        RECT 7.68 9.708 7.712 12.216 ;
  LAYER M3 ;
        RECT 7.744 9.708 7.776 12.216 ;
  LAYER M3 ;
        RECT 7.808 9.708 7.84 12.216 ;
  LAYER M3 ;
        RECT 7.872 9.708 7.904 12.216 ;
  LAYER M3 ;
        RECT 7.936 9.708 7.968 12.216 ;
  LAYER M3 ;
        RECT 8 9.708 8.032 12.216 ;
  LAYER M3 ;
        RECT 8.064 9.708 8.096 12.216 ;
  LAYER M3 ;
        RECT 8.128 9.708 8.16 12.216 ;
  LAYER M3 ;
        RECT 8.192 9.708 8.224 12.216 ;
  LAYER M3 ;
        RECT 8.256 9.708 8.288 12.216 ;
  LAYER M3 ;
        RECT 8.32 9.708 8.352 12.216 ;
  LAYER M3 ;
        RECT 8.384 9.708 8.416 12.216 ;
  LAYER M3 ;
        RECT 8.448 9.708 8.48 12.216 ;
  LAYER M3 ;
        RECT 8.544 9.708 8.576 12.216 ;
  LAYER M1 ;
        RECT 6.159 9.744 6.161 12.18 ;
  LAYER M1 ;
        RECT 6.239 9.744 6.241 12.18 ;
  LAYER M1 ;
        RECT 6.319 9.744 6.321 12.18 ;
  LAYER M1 ;
        RECT 6.399 9.744 6.401 12.18 ;
  LAYER M1 ;
        RECT 6.479 9.744 6.481 12.18 ;
  LAYER M1 ;
        RECT 6.559 9.744 6.561 12.18 ;
  LAYER M1 ;
        RECT 6.639 9.744 6.641 12.18 ;
  LAYER M1 ;
        RECT 6.719 9.744 6.721 12.18 ;
  LAYER M1 ;
        RECT 6.799 9.744 6.801 12.18 ;
  LAYER M1 ;
        RECT 6.879 9.744 6.881 12.18 ;
  LAYER M1 ;
        RECT 6.959 9.744 6.961 12.18 ;
  LAYER M1 ;
        RECT 7.039 9.744 7.041 12.18 ;
  LAYER M1 ;
        RECT 7.119 9.744 7.121 12.18 ;
  LAYER M1 ;
        RECT 7.199 9.744 7.201 12.18 ;
  LAYER M1 ;
        RECT 7.279 9.744 7.281 12.18 ;
  LAYER M1 ;
        RECT 7.359 9.744 7.361 12.18 ;
  LAYER M1 ;
        RECT 7.439 9.744 7.441 12.18 ;
  LAYER M1 ;
        RECT 7.519 9.744 7.521 12.18 ;
  LAYER M1 ;
        RECT 7.599 9.744 7.601 12.18 ;
  LAYER M1 ;
        RECT 7.679 9.744 7.681 12.18 ;
  LAYER M1 ;
        RECT 7.759 9.744 7.761 12.18 ;
  LAYER M1 ;
        RECT 7.839 9.744 7.841 12.18 ;
  LAYER M1 ;
        RECT 7.919 9.744 7.921 12.18 ;
  LAYER M1 ;
        RECT 7.999 9.744 8.001 12.18 ;
  LAYER M1 ;
        RECT 8.079 9.744 8.081 12.18 ;
  LAYER M1 ;
        RECT 8.159 9.744 8.161 12.18 ;
  LAYER M1 ;
        RECT 8.239 9.744 8.241 12.18 ;
  LAYER M1 ;
        RECT 8.319 9.744 8.321 12.18 ;
  LAYER M1 ;
        RECT 8.399 9.744 8.401 12.18 ;
  LAYER M1 ;
        RECT 8.479 9.744 8.481 12.18 ;
  LAYER M2 ;
        RECT 6.16 9.743 8.56 9.745 ;
  LAYER M2 ;
        RECT 6.16 9.827 8.56 9.829 ;
  LAYER M2 ;
        RECT 6.16 9.911 8.56 9.913 ;
  LAYER M2 ;
        RECT 6.16 9.995 8.56 9.997 ;
  LAYER M2 ;
        RECT 6.16 10.079 8.56 10.081 ;
  LAYER M2 ;
        RECT 6.16 10.163 8.56 10.165 ;
  LAYER M2 ;
        RECT 6.16 10.247 8.56 10.249 ;
  LAYER M2 ;
        RECT 6.16 10.331 8.56 10.333 ;
  LAYER M2 ;
        RECT 6.16 10.415 8.56 10.417 ;
  LAYER M2 ;
        RECT 6.16 10.499 8.56 10.501 ;
  LAYER M2 ;
        RECT 6.16 10.583 8.56 10.585 ;
  LAYER M2 ;
        RECT 6.16 10.667 8.56 10.669 ;
  LAYER M2 ;
        RECT 6.16 10.7505 8.56 10.7525 ;
  LAYER M2 ;
        RECT 6.16 10.835 8.56 10.837 ;
  LAYER M2 ;
        RECT 6.16 10.919 8.56 10.921 ;
  LAYER M2 ;
        RECT 6.16 11.003 8.56 11.005 ;
  LAYER M2 ;
        RECT 6.16 11.087 8.56 11.089 ;
  LAYER M2 ;
        RECT 6.16 11.171 8.56 11.173 ;
  LAYER M2 ;
        RECT 6.16 11.255 8.56 11.257 ;
  LAYER M2 ;
        RECT 6.16 11.339 8.56 11.341 ;
  LAYER M2 ;
        RECT 6.16 11.423 8.56 11.425 ;
  LAYER M2 ;
        RECT 6.16 11.507 8.56 11.509 ;
  LAYER M2 ;
        RECT 6.16 11.591 8.56 11.593 ;
  LAYER M2 ;
        RECT 6.16 11.675 8.56 11.677 ;
  LAYER M2 ;
        RECT 6.16 11.759 8.56 11.761 ;
  LAYER M2 ;
        RECT 6.16 11.843 8.56 11.845 ;
  LAYER M2 ;
        RECT 6.16 11.927 8.56 11.929 ;
  LAYER M2 ;
        RECT 6.16 12.011 8.56 12.013 ;
  LAYER M2 ;
        RECT 6.16 12.095 8.56 12.097 ;
  LAYER M1 ;
        RECT 6.144 12.648 6.176 15.156 ;
  LAYER M1 ;
        RECT 6.208 12.648 6.24 15.156 ;
  LAYER M1 ;
        RECT 6.272 12.648 6.304 15.156 ;
  LAYER M1 ;
        RECT 6.336 12.648 6.368 15.156 ;
  LAYER M1 ;
        RECT 6.4 12.648 6.432 15.156 ;
  LAYER M1 ;
        RECT 6.464 12.648 6.496 15.156 ;
  LAYER M1 ;
        RECT 6.528 12.648 6.56 15.156 ;
  LAYER M1 ;
        RECT 6.592 12.648 6.624 15.156 ;
  LAYER M1 ;
        RECT 6.656 12.648 6.688 15.156 ;
  LAYER M1 ;
        RECT 6.72 12.648 6.752 15.156 ;
  LAYER M1 ;
        RECT 6.784 12.648 6.816 15.156 ;
  LAYER M1 ;
        RECT 6.848 12.648 6.88 15.156 ;
  LAYER M1 ;
        RECT 6.912 12.648 6.944 15.156 ;
  LAYER M1 ;
        RECT 6.976 12.648 7.008 15.156 ;
  LAYER M1 ;
        RECT 7.04 12.648 7.072 15.156 ;
  LAYER M1 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M1 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M1 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M1 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M1 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M1 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M1 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M1 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M1 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M1 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M1 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M1 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M1 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M1 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M1 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M1 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M1 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M1 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M1 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M1 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M1 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M1 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M2 ;
        RECT 6.124 12.732 8.596 12.764 ;
  LAYER M2 ;
        RECT 6.124 12.796 8.596 12.828 ;
  LAYER M2 ;
        RECT 6.124 12.86 8.596 12.892 ;
  LAYER M2 ;
        RECT 6.124 12.924 8.596 12.956 ;
  LAYER M2 ;
        RECT 6.124 12.988 8.596 13.02 ;
  LAYER M2 ;
        RECT 6.124 13.052 8.596 13.084 ;
  LAYER M2 ;
        RECT 6.124 13.116 8.596 13.148 ;
  LAYER M2 ;
        RECT 6.124 13.18 8.596 13.212 ;
  LAYER M2 ;
        RECT 6.124 13.244 8.596 13.276 ;
  LAYER M2 ;
        RECT 6.124 13.308 8.596 13.34 ;
  LAYER M2 ;
        RECT 6.124 13.372 8.596 13.404 ;
  LAYER M2 ;
        RECT 6.124 13.436 8.596 13.468 ;
  LAYER M2 ;
        RECT 6.124 13.5 8.596 13.532 ;
  LAYER M2 ;
        RECT 6.124 13.564 8.596 13.596 ;
  LAYER M2 ;
        RECT 6.124 13.628 8.596 13.66 ;
  LAYER M2 ;
        RECT 6.124 13.692 8.596 13.724 ;
  LAYER M2 ;
        RECT 6.124 13.756 8.596 13.788 ;
  LAYER M2 ;
        RECT 6.124 13.82 8.596 13.852 ;
  LAYER M2 ;
        RECT 6.124 13.884 8.596 13.916 ;
  LAYER M2 ;
        RECT 6.124 13.948 8.596 13.98 ;
  LAYER M2 ;
        RECT 6.124 14.012 8.596 14.044 ;
  LAYER M2 ;
        RECT 6.124 14.076 8.596 14.108 ;
  LAYER M2 ;
        RECT 6.124 14.14 8.596 14.172 ;
  LAYER M2 ;
        RECT 6.124 14.204 8.596 14.236 ;
  LAYER M2 ;
        RECT 6.124 14.268 8.596 14.3 ;
  LAYER M2 ;
        RECT 6.124 14.332 8.596 14.364 ;
  LAYER M2 ;
        RECT 6.124 14.396 8.596 14.428 ;
  LAYER M2 ;
        RECT 6.124 14.46 8.596 14.492 ;
  LAYER M2 ;
        RECT 6.124 14.524 8.596 14.556 ;
  LAYER M2 ;
        RECT 6.124 14.588 8.596 14.62 ;
  LAYER M2 ;
        RECT 6.124 14.652 8.596 14.684 ;
  LAYER M2 ;
        RECT 6.124 14.716 8.596 14.748 ;
  LAYER M2 ;
        RECT 6.124 14.78 8.596 14.812 ;
  LAYER M2 ;
        RECT 6.124 14.844 8.596 14.876 ;
  LAYER M2 ;
        RECT 6.124 14.908 8.596 14.94 ;
  LAYER M2 ;
        RECT 6.124 14.972 8.596 15.004 ;
  LAYER M3 ;
        RECT 6.144 12.648 6.176 15.156 ;
  LAYER M3 ;
        RECT 6.208 12.648 6.24 15.156 ;
  LAYER M3 ;
        RECT 6.272 12.648 6.304 15.156 ;
  LAYER M3 ;
        RECT 6.336 12.648 6.368 15.156 ;
  LAYER M3 ;
        RECT 6.4 12.648 6.432 15.156 ;
  LAYER M3 ;
        RECT 6.464 12.648 6.496 15.156 ;
  LAYER M3 ;
        RECT 6.528 12.648 6.56 15.156 ;
  LAYER M3 ;
        RECT 6.592 12.648 6.624 15.156 ;
  LAYER M3 ;
        RECT 6.656 12.648 6.688 15.156 ;
  LAYER M3 ;
        RECT 6.72 12.648 6.752 15.156 ;
  LAYER M3 ;
        RECT 6.784 12.648 6.816 15.156 ;
  LAYER M3 ;
        RECT 6.848 12.648 6.88 15.156 ;
  LAYER M3 ;
        RECT 6.912 12.648 6.944 15.156 ;
  LAYER M3 ;
        RECT 6.976 12.648 7.008 15.156 ;
  LAYER M3 ;
        RECT 7.04 12.648 7.072 15.156 ;
  LAYER M3 ;
        RECT 7.104 12.648 7.136 15.156 ;
  LAYER M3 ;
        RECT 7.168 12.648 7.2 15.156 ;
  LAYER M3 ;
        RECT 7.232 12.648 7.264 15.156 ;
  LAYER M3 ;
        RECT 7.296 12.648 7.328 15.156 ;
  LAYER M3 ;
        RECT 7.36 12.648 7.392 15.156 ;
  LAYER M3 ;
        RECT 7.424 12.648 7.456 15.156 ;
  LAYER M3 ;
        RECT 7.488 12.648 7.52 15.156 ;
  LAYER M3 ;
        RECT 7.552 12.648 7.584 15.156 ;
  LAYER M3 ;
        RECT 7.616 12.648 7.648 15.156 ;
  LAYER M3 ;
        RECT 7.68 12.648 7.712 15.156 ;
  LAYER M3 ;
        RECT 7.744 12.648 7.776 15.156 ;
  LAYER M3 ;
        RECT 7.808 12.648 7.84 15.156 ;
  LAYER M3 ;
        RECT 7.872 12.648 7.904 15.156 ;
  LAYER M3 ;
        RECT 7.936 12.648 7.968 15.156 ;
  LAYER M3 ;
        RECT 8 12.648 8.032 15.156 ;
  LAYER M3 ;
        RECT 8.064 12.648 8.096 15.156 ;
  LAYER M3 ;
        RECT 8.128 12.648 8.16 15.156 ;
  LAYER M3 ;
        RECT 8.192 12.648 8.224 15.156 ;
  LAYER M3 ;
        RECT 8.256 12.648 8.288 15.156 ;
  LAYER M3 ;
        RECT 8.32 12.648 8.352 15.156 ;
  LAYER M3 ;
        RECT 8.384 12.648 8.416 15.156 ;
  LAYER M3 ;
        RECT 8.448 12.648 8.48 15.156 ;
  LAYER M3 ;
        RECT 8.544 12.648 8.576 15.156 ;
  LAYER M1 ;
        RECT 6.159 12.684 6.161 15.12 ;
  LAYER M1 ;
        RECT 6.239 12.684 6.241 15.12 ;
  LAYER M1 ;
        RECT 6.319 12.684 6.321 15.12 ;
  LAYER M1 ;
        RECT 6.399 12.684 6.401 15.12 ;
  LAYER M1 ;
        RECT 6.479 12.684 6.481 15.12 ;
  LAYER M1 ;
        RECT 6.559 12.684 6.561 15.12 ;
  LAYER M1 ;
        RECT 6.639 12.684 6.641 15.12 ;
  LAYER M1 ;
        RECT 6.719 12.684 6.721 15.12 ;
  LAYER M1 ;
        RECT 6.799 12.684 6.801 15.12 ;
  LAYER M1 ;
        RECT 6.879 12.684 6.881 15.12 ;
  LAYER M1 ;
        RECT 6.959 12.684 6.961 15.12 ;
  LAYER M1 ;
        RECT 7.039 12.684 7.041 15.12 ;
  LAYER M1 ;
        RECT 7.119 12.684 7.121 15.12 ;
  LAYER M1 ;
        RECT 7.199 12.684 7.201 15.12 ;
  LAYER M1 ;
        RECT 7.279 12.684 7.281 15.12 ;
  LAYER M1 ;
        RECT 7.359 12.684 7.361 15.12 ;
  LAYER M1 ;
        RECT 7.439 12.684 7.441 15.12 ;
  LAYER M1 ;
        RECT 7.519 12.684 7.521 15.12 ;
  LAYER M1 ;
        RECT 7.599 12.684 7.601 15.12 ;
  LAYER M1 ;
        RECT 7.679 12.684 7.681 15.12 ;
  LAYER M1 ;
        RECT 7.759 12.684 7.761 15.12 ;
  LAYER M1 ;
        RECT 7.839 12.684 7.841 15.12 ;
  LAYER M1 ;
        RECT 7.919 12.684 7.921 15.12 ;
  LAYER M1 ;
        RECT 7.999 12.684 8.001 15.12 ;
  LAYER M1 ;
        RECT 8.079 12.684 8.081 15.12 ;
  LAYER M1 ;
        RECT 8.159 12.684 8.161 15.12 ;
  LAYER M1 ;
        RECT 8.239 12.684 8.241 15.12 ;
  LAYER M1 ;
        RECT 8.319 12.684 8.321 15.12 ;
  LAYER M1 ;
        RECT 8.399 12.684 8.401 15.12 ;
  LAYER M1 ;
        RECT 8.479 12.684 8.481 15.12 ;
  LAYER M2 ;
        RECT 6.16 12.683 8.56 12.685 ;
  LAYER M2 ;
        RECT 6.16 12.767 8.56 12.769 ;
  LAYER M2 ;
        RECT 6.16 12.851 8.56 12.853 ;
  LAYER M2 ;
        RECT 6.16 12.935 8.56 12.937 ;
  LAYER M2 ;
        RECT 6.16 13.019 8.56 13.021 ;
  LAYER M2 ;
        RECT 6.16 13.103 8.56 13.105 ;
  LAYER M2 ;
        RECT 6.16 13.187 8.56 13.189 ;
  LAYER M2 ;
        RECT 6.16 13.271 8.56 13.273 ;
  LAYER M2 ;
        RECT 6.16 13.355 8.56 13.357 ;
  LAYER M2 ;
        RECT 6.16 13.439 8.56 13.441 ;
  LAYER M2 ;
        RECT 6.16 13.523 8.56 13.525 ;
  LAYER M2 ;
        RECT 6.16 13.607 8.56 13.609 ;
  LAYER M2 ;
        RECT 6.16 13.6905 8.56 13.6925 ;
  LAYER M2 ;
        RECT 6.16 13.775 8.56 13.777 ;
  LAYER M2 ;
        RECT 6.16 13.859 8.56 13.861 ;
  LAYER M2 ;
        RECT 6.16 13.943 8.56 13.945 ;
  LAYER M2 ;
        RECT 6.16 14.027 8.56 14.029 ;
  LAYER M2 ;
        RECT 6.16 14.111 8.56 14.113 ;
  LAYER M2 ;
        RECT 6.16 14.195 8.56 14.197 ;
  LAYER M2 ;
        RECT 6.16 14.279 8.56 14.281 ;
  LAYER M2 ;
        RECT 6.16 14.363 8.56 14.365 ;
  LAYER M2 ;
        RECT 6.16 14.447 8.56 14.449 ;
  LAYER M2 ;
        RECT 6.16 14.531 8.56 14.533 ;
  LAYER M2 ;
        RECT 6.16 14.615 8.56 14.617 ;
  LAYER M2 ;
        RECT 6.16 14.699 8.56 14.701 ;
  LAYER M2 ;
        RECT 6.16 14.783 8.56 14.785 ;
  LAYER M2 ;
        RECT 6.16 14.867 8.56 14.869 ;
  LAYER M2 ;
        RECT 6.16 14.951 8.56 14.953 ;
  LAYER M2 ;
        RECT 6.16 15.035 8.56 15.037 ;
  LAYER M1 ;
        RECT 6.144 15.588 6.176 18.096 ;
  LAYER M1 ;
        RECT 6.208 15.588 6.24 18.096 ;
  LAYER M1 ;
        RECT 6.272 15.588 6.304 18.096 ;
  LAYER M1 ;
        RECT 6.336 15.588 6.368 18.096 ;
  LAYER M1 ;
        RECT 6.4 15.588 6.432 18.096 ;
  LAYER M1 ;
        RECT 6.464 15.588 6.496 18.096 ;
  LAYER M1 ;
        RECT 6.528 15.588 6.56 18.096 ;
  LAYER M1 ;
        RECT 6.592 15.588 6.624 18.096 ;
  LAYER M1 ;
        RECT 6.656 15.588 6.688 18.096 ;
  LAYER M1 ;
        RECT 6.72 15.588 6.752 18.096 ;
  LAYER M1 ;
        RECT 6.784 15.588 6.816 18.096 ;
  LAYER M1 ;
        RECT 6.848 15.588 6.88 18.096 ;
  LAYER M1 ;
        RECT 6.912 15.588 6.944 18.096 ;
  LAYER M1 ;
        RECT 6.976 15.588 7.008 18.096 ;
  LAYER M1 ;
        RECT 7.04 15.588 7.072 18.096 ;
  LAYER M1 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M1 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M1 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M1 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M1 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M1 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M1 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M1 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M1 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M1 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M1 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M1 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M1 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M1 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M1 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M1 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M1 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M1 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M1 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M1 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M1 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M1 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M2 ;
        RECT 6.124 15.672 8.596 15.704 ;
  LAYER M2 ;
        RECT 6.124 15.736 8.596 15.768 ;
  LAYER M2 ;
        RECT 6.124 15.8 8.596 15.832 ;
  LAYER M2 ;
        RECT 6.124 15.864 8.596 15.896 ;
  LAYER M2 ;
        RECT 6.124 15.928 8.596 15.96 ;
  LAYER M2 ;
        RECT 6.124 15.992 8.596 16.024 ;
  LAYER M2 ;
        RECT 6.124 16.056 8.596 16.088 ;
  LAYER M2 ;
        RECT 6.124 16.12 8.596 16.152 ;
  LAYER M2 ;
        RECT 6.124 16.184 8.596 16.216 ;
  LAYER M2 ;
        RECT 6.124 16.248 8.596 16.28 ;
  LAYER M2 ;
        RECT 6.124 16.312 8.596 16.344 ;
  LAYER M2 ;
        RECT 6.124 16.376 8.596 16.408 ;
  LAYER M2 ;
        RECT 6.124 16.44 8.596 16.472 ;
  LAYER M2 ;
        RECT 6.124 16.504 8.596 16.536 ;
  LAYER M2 ;
        RECT 6.124 16.568 8.596 16.6 ;
  LAYER M2 ;
        RECT 6.124 16.632 8.596 16.664 ;
  LAYER M2 ;
        RECT 6.124 16.696 8.596 16.728 ;
  LAYER M2 ;
        RECT 6.124 16.76 8.596 16.792 ;
  LAYER M2 ;
        RECT 6.124 16.824 8.596 16.856 ;
  LAYER M2 ;
        RECT 6.124 16.888 8.596 16.92 ;
  LAYER M2 ;
        RECT 6.124 16.952 8.596 16.984 ;
  LAYER M2 ;
        RECT 6.124 17.016 8.596 17.048 ;
  LAYER M2 ;
        RECT 6.124 17.08 8.596 17.112 ;
  LAYER M2 ;
        RECT 6.124 17.144 8.596 17.176 ;
  LAYER M2 ;
        RECT 6.124 17.208 8.596 17.24 ;
  LAYER M2 ;
        RECT 6.124 17.272 8.596 17.304 ;
  LAYER M2 ;
        RECT 6.124 17.336 8.596 17.368 ;
  LAYER M2 ;
        RECT 6.124 17.4 8.596 17.432 ;
  LAYER M2 ;
        RECT 6.124 17.464 8.596 17.496 ;
  LAYER M2 ;
        RECT 6.124 17.528 8.596 17.56 ;
  LAYER M2 ;
        RECT 6.124 17.592 8.596 17.624 ;
  LAYER M2 ;
        RECT 6.124 17.656 8.596 17.688 ;
  LAYER M2 ;
        RECT 6.124 17.72 8.596 17.752 ;
  LAYER M2 ;
        RECT 6.124 17.784 8.596 17.816 ;
  LAYER M2 ;
        RECT 6.124 17.848 8.596 17.88 ;
  LAYER M2 ;
        RECT 6.124 17.912 8.596 17.944 ;
  LAYER M3 ;
        RECT 6.144 15.588 6.176 18.096 ;
  LAYER M3 ;
        RECT 6.208 15.588 6.24 18.096 ;
  LAYER M3 ;
        RECT 6.272 15.588 6.304 18.096 ;
  LAYER M3 ;
        RECT 6.336 15.588 6.368 18.096 ;
  LAYER M3 ;
        RECT 6.4 15.588 6.432 18.096 ;
  LAYER M3 ;
        RECT 6.464 15.588 6.496 18.096 ;
  LAYER M3 ;
        RECT 6.528 15.588 6.56 18.096 ;
  LAYER M3 ;
        RECT 6.592 15.588 6.624 18.096 ;
  LAYER M3 ;
        RECT 6.656 15.588 6.688 18.096 ;
  LAYER M3 ;
        RECT 6.72 15.588 6.752 18.096 ;
  LAYER M3 ;
        RECT 6.784 15.588 6.816 18.096 ;
  LAYER M3 ;
        RECT 6.848 15.588 6.88 18.096 ;
  LAYER M3 ;
        RECT 6.912 15.588 6.944 18.096 ;
  LAYER M3 ;
        RECT 6.976 15.588 7.008 18.096 ;
  LAYER M3 ;
        RECT 7.04 15.588 7.072 18.096 ;
  LAYER M3 ;
        RECT 7.104 15.588 7.136 18.096 ;
  LAYER M3 ;
        RECT 7.168 15.588 7.2 18.096 ;
  LAYER M3 ;
        RECT 7.232 15.588 7.264 18.096 ;
  LAYER M3 ;
        RECT 7.296 15.588 7.328 18.096 ;
  LAYER M3 ;
        RECT 7.36 15.588 7.392 18.096 ;
  LAYER M3 ;
        RECT 7.424 15.588 7.456 18.096 ;
  LAYER M3 ;
        RECT 7.488 15.588 7.52 18.096 ;
  LAYER M3 ;
        RECT 7.552 15.588 7.584 18.096 ;
  LAYER M3 ;
        RECT 7.616 15.588 7.648 18.096 ;
  LAYER M3 ;
        RECT 7.68 15.588 7.712 18.096 ;
  LAYER M3 ;
        RECT 7.744 15.588 7.776 18.096 ;
  LAYER M3 ;
        RECT 7.808 15.588 7.84 18.096 ;
  LAYER M3 ;
        RECT 7.872 15.588 7.904 18.096 ;
  LAYER M3 ;
        RECT 7.936 15.588 7.968 18.096 ;
  LAYER M3 ;
        RECT 8 15.588 8.032 18.096 ;
  LAYER M3 ;
        RECT 8.064 15.588 8.096 18.096 ;
  LAYER M3 ;
        RECT 8.128 15.588 8.16 18.096 ;
  LAYER M3 ;
        RECT 8.192 15.588 8.224 18.096 ;
  LAYER M3 ;
        RECT 8.256 15.588 8.288 18.096 ;
  LAYER M3 ;
        RECT 8.32 15.588 8.352 18.096 ;
  LAYER M3 ;
        RECT 8.384 15.588 8.416 18.096 ;
  LAYER M3 ;
        RECT 8.448 15.588 8.48 18.096 ;
  LAYER M3 ;
        RECT 8.544 15.588 8.576 18.096 ;
  LAYER M1 ;
        RECT 6.159 15.624 6.161 18.06 ;
  LAYER M1 ;
        RECT 6.239 15.624 6.241 18.06 ;
  LAYER M1 ;
        RECT 6.319 15.624 6.321 18.06 ;
  LAYER M1 ;
        RECT 6.399 15.624 6.401 18.06 ;
  LAYER M1 ;
        RECT 6.479 15.624 6.481 18.06 ;
  LAYER M1 ;
        RECT 6.559 15.624 6.561 18.06 ;
  LAYER M1 ;
        RECT 6.639 15.624 6.641 18.06 ;
  LAYER M1 ;
        RECT 6.719 15.624 6.721 18.06 ;
  LAYER M1 ;
        RECT 6.799 15.624 6.801 18.06 ;
  LAYER M1 ;
        RECT 6.879 15.624 6.881 18.06 ;
  LAYER M1 ;
        RECT 6.959 15.624 6.961 18.06 ;
  LAYER M1 ;
        RECT 7.039 15.624 7.041 18.06 ;
  LAYER M1 ;
        RECT 7.119 15.624 7.121 18.06 ;
  LAYER M1 ;
        RECT 7.199 15.624 7.201 18.06 ;
  LAYER M1 ;
        RECT 7.279 15.624 7.281 18.06 ;
  LAYER M1 ;
        RECT 7.359 15.624 7.361 18.06 ;
  LAYER M1 ;
        RECT 7.439 15.624 7.441 18.06 ;
  LAYER M1 ;
        RECT 7.519 15.624 7.521 18.06 ;
  LAYER M1 ;
        RECT 7.599 15.624 7.601 18.06 ;
  LAYER M1 ;
        RECT 7.679 15.624 7.681 18.06 ;
  LAYER M1 ;
        RECT 7.759 15.624 7.761 18.06 ;
  LAYER M1 ;
        RECT 7.839 15.624 7.841 18.06 ;
  LAYER M1 ;
        RECT 7.919 15.624 7.921 18.06 ;
  LAYER M1 ;
        RECT 7.999 15.624 8.001 18.06 ;
  LAYER M1 ;
        RECT 8.079 15.624 8.081 18.06 ;
  LAYER M1 ;
        RECT 8.159 15.624 8.161 18.06 ;
  LAYER M1 ;
        RECT 8.239 15.624 8.241 18.06 ;
  LAYER M1 ;
        RECT 8.319 15.624 8.321 18.06 ;
  LAYER M1 ;
        RECT 8.399 15.624 8.401 18.06 ;
  LAYER M1 ;
        RECT 8.479 15.624 8.481 18.06 ;
  LAYER M2 ;
        RECT 6.16 15.623 8.56 15.625 ;
  LAYER M2 ;
        RECT 6.16 15.707 8.56 15.709 ;
  LAYER M2 ;
        RECT 6.16 15.791 8.56 15.793 ;
  LAYER M2 ;
        RECT 6.16 15.875 8.56 15.877 ;
  LAYER M2 ;
        RECT 6.16 15.959 8.56 15.961 ;
  LAYER M2 ;
        RECT 6.16 16.043 8.56 16.045 ;
  LAYER M2 ;
        RECT 6.16 16.127 8.56 16.129 ;
  LAYER M2 ;
        RECT 6.16 16.211 8.56 16.213 ;
  LAYER M2 ;
        RECT 6.16 16.295 8.56 16.297 ;
  LAYER M2 ;
        RECT 6.16 16.379 8.56 16.381 ;
  LAYER M2 ;
        RECT 6.16 16.463 8.56 16.465 ;
  LAYER M2 ;
        RECT 6.16 16.547 8.56 16.549 ;
  LAYER M2 ;
        RECT 6.16 16.6305 8.56 16.6325 ;
  LAYER M2 ;
        RECT 6.16 16.715 8.56 16.717 ;
  LAYER M2 ;
        RECT 6.16 16.799 8.56 16.801 ;
  LAYER M2 ;
        RECT 6.16 16.883 8.56 16.885 ;
  LAYER M2 ;
        RECT 6.16 16.967 8.56 16.969 ;
  LAYER M2 ;
        RECT 6.16 17.051 8.56 17.053 ;
  LAYER M2 ;
        RECT 6.16 17.135 8.56 17.137 ;
  LAYER M2 ;
        RECT 6.16 17.219 8.56 17.221 ;
  LAYER M2 ;
        RECT 6.16 17.303 8.56 17.305 ;
  LAYER M2 ;
        RECT 6.16 17.387 8.56 17.389 ;
  LAYER M2 ;
        RECT 6.16 17.471 8.56 17.473 ;
  LAYER M2 ;
        RECT 6.16 17.555 8.56 17.557 ;
  LAYER M2 ;
        RECT 6.16 17.639 8.56 17.641 ;
  LAYER M2 ;
        RECT 6.16 17.723 8.56 17.725 ;
  LAYER M2 ;
        RECT 6.16 17.807 8.56 17.809 ;
  LAYER M2 ;
        RECT 6.16 17.891 8.56 17.893 ;
  LAYER M2 ;
        RECT 6.16 17.975 8.56 17.977 ;
  LAYER M1 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M1 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M1 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M1 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M1 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M1 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M1 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M1 ;
        RECT 9.472 0.888 9.504 3.396 ;
  LAYER M1 ;
        RECT 9.536 0.888 9.568 3.396 ;
  LAYER M1 ;
        RECT 9.6 0.888 9.632 3.396 ;
  LAYER M1 ;
        RECT 9.664 0.888 9.696 3.396 ;
  LAYER M1 ;
        RECT 9.728 0.888 9.76 3.396 ;
  LAYER M1 ;
        RECT 9.792 0.888 9.824 3.396 ;
  LAYER M1 ;
        RECT 9.856 0.888 9.888 3.396 ;
  LAYER M1 ;
        RECT 9.92 0.888 9.952 3.396 ;
  LAYER M1 ;
        RECT 9.984 0.888 10.016 3.396 ;
  LAYER M1 ;
        RECT 10.048 0.888 10.08 3.396 ;
  LAYER M1 ;
        RECT 10.112 0.888 10.144 3.396 ;
  LAYER M1 ;
        RECT 10.176 0.888 10.208 3.396 ;
  LAYER M1 ;
        RECT 10.24 0.888 10.272 3.396 ;
  LAYER M1 ;
        RECT 10.304 0.888 10.336 3.396 ;
  LAYER M1 ;
        RECT 10.368 0.888 10.4 3.396 ;
  LAYER M1 ;
        RECT 10.432 0.888 10.464 3.396 ;
  LAYER M1 ;
        RECT 10.496 0.888 10.528 3.396 ;
  LAYER M1 ;
        RECT 10.56 0.888 10.592 3.396 ;
  LAYER M1 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M1 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M1 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M1 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M1 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M1 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M1 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M1 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M1 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M1 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M1 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M1 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M2 ;
        RECT 9.004 0.972 11.476 1.004 ;
  LAYER M2 ;
        RECT 9.004 1.036 11.476 1.068 ;
  LAYER M2 ;
        RECT 9.004 1.1 11.476 1.132 ;
  LAYER M2 ;
        RECT 9.004 1.164 11.476 1.196 ;
  LAYER M2 ;
        RECT 9.004 1.228 11.476 1.26 ;
  LAYER M2 ;
        RECT 9.004 1.292 11.476 1.324 ;
  LAYER M2 ;
        RECT 9.004 1.356 11.476 1.388 ;
  LAYER M2 ;
        RECT 9.004 1.42 11.476 1.452 ;
  LAYER M2 ;
        RECT 9.004 1.484 11.476 1.516 ;
  LAYER M2 ;
        RECT 9.004 1.548 11.476 1.58 ;
  LAYER M2 ;
        RECT 9.004 1.612 11.476 1.644 ;
  LAYER M2 ;
        RECT 9.004 1.676 11.476 1.708 ;
  LAYER M2 ;
        RECT 9.004 1.74 11.476 1.772 ;
  LAYER M2 ;
        RECT 9.004 1.804 11.476 1.836 ;
  LAYER M2 ;
        RECT 9.004 1.868 11.476 1.9 ;
  LAYER M2 ;
        RECT 9.004 1.932 11.476 1.964 ;
  LAYER M2 ;
        RECT 9.004 1.996 11.476 2.028 ;
  LAYER M2 ;
        RECT 9.004 2.06 11.476 2.092 ;
  LAYER M2 ;
        RECT 9.004 2.124 11.476 2.156 ;
  LAYER M2 ;
        RECT 9.004 2.188 11.476 2.22 ;
  LAYER M2 ;
        RECT 9.004 2.252 11.476 2.284 ;
  LAYER M2 ;
        RECT 9.004 2.316 11.476 2.348 ;
  LAYER M2 ;
        RECT 9.004 2.38 11.476 2.412 ;
  LAYER M2 ;
        RECT 9.004 2.444 11.476 2.476 ;
  LAYER M2 ;
        RECT 9.004 2.508 11.476 2.54 ;
  LAYER M2 ;
        RECT 9.004 2.572 11.476 2.604 ;
  LAYER M2 ;
        RECT 9.004 2.636 11.476 2.668 ;
  LAYER M2 ;
        RECT 9.004 2.7 11.476 2.732 ;
  LAYER M2 ;
        RECT 9.004 2.764 11.476 2.796 ;
  LAYER M2 ;
        RECT 9.004 2.828 11.476 2.86 ;
  LAYER M2 ;
        RECT 9.004 2.892 11.476 2.924 ;
  LAYER M2 ;
        RECT 9.004 2.956 11.476 2.988 ;
  LAYER M2 ;
        RECT 9.004 3.02 11.476 3.052 ;
  LAYER M2 ;
        RECT 9.004 3.084 11.476 3.116 ;
  LAYER M2 ;
        RECT 9.004 3.148 11.476 3.18 ;
  LAYER M2 ;
        RECT 9.004 3.212 11.476 3.244 ;
  LAYER M3 ;
        RECT 9.024 0.888 9.056 3.396 ;
  LAYER M3 ;
        RECT 9.088 0.888 9.12 3.396 ;
  LAYER M3 ;
        RECT 9.152 0.888 9.184 3.396 ;
  LAYER M3 ;
        RECT 9.216 0.888 9.248 3.396 ;
  LAYER M3 ;
        RECT 9.28 0.888 9.312 3.396 ;
  LAYER M3 ;
        RECT 9.344 0.888 9.376 3.396 ;
  LAYER M3 ;
        RECT 9.408 0.888 9.44 3.396 ;
  LAYER M3 ;
        RECT 9.472 0.888 9.504 3.396 ;
  LAYER M3 ;
        RECT 9.536 0.888 9.568 3.396 ;
  LAYER M3 ;
        RECT 9.6 0.888 9.632 3.396 ;
  LAYER M3 ;
        RECT 9.664 0.888 9.696 3.396 ;
  LAYER M3 ;
        RECT 9.728 0.888 9.76 3.396 ;
  LAYER M3 ;
        RECT 9.792 0.888 9.824 3.396 ;
  LAYER M3 ;
        RECT 9.856 0.888 9.888 3.396 ;
  LAYER M3 ;
        RECT 9.92 0.888 9.952 3.396 ;
  LAYER M3 ;
        RECT 9.984 0.888 10.016 3.396 ;
  LAYER M3 ;
        RECT 10.048 0.888 10.08 3.396 ;
  LAYER M3 ;
        RECT 10.112 0.888 10.144 3.396 ;
  LAYER M3 ;
        RECT 10.176 0.888 10.208 3.396 ;
  LAYER M3 ;
        RECT 10.24 0.888 10.272 3.396 ;
  LAYER M3 ;
        RECT 10.304 0.888 10.336 3.396 ;
  LAYER M3 ;
        RECT 10.368 0.888 10.4 3.396 ;
  LAYER M3 ;
        RECT 10.432 0.888 10.464 3.396 ;
  LAYER M3 ;
        RECT 10.496 0.888 10.528 3.396 ;
  LAYER M3 ;
        RECT 10.56 0.888 10.592 3.396 ;
  LAYER M3 ;
        RECT 10.624 0.888 10.656 3.396 ;
  LAYER M3 ;
        RECT 10.688 0.888 10.72 3.396 ;
  LAYER M3 ;
        RECT 10.752 0.888 10.784 3.396 ;
  LAYER M3 ;
        RECT 10.816 0.888 10.848 3.396 ;
  LAYER M3 ;
        RECT 10.88 0.888 10.912 3.396 ;
  LAYER M3 ;
        RECT 10.944 0.888 10.976 3.396 ;
  LAYER M3 ;
        RECT 11.008 0.888 11.04 3.396 ;
  LAYER M3 ;
        RECT 11.072 0.888 11.104 3.396 ;
  LAYER M3 ;
        RECT 11.136 0.888 11.168 3.396 ;
  LAYER M3 ;
        RECT 11.2 0.888 11.232 3.396 ;
  LAYER M3 ;
        RECT 11.264 0.888 11.296 3.396 ;
  LAYER M3 ;
        RECT 11.328 0.888 11.36 3.396 ;
  LAYER M3 ;
        RECT 11.424 0.888 11.456 3.396 ;
  LAYER M1 ;
        RECT 9.039 0.924 9.041 3.36 ;
  LAYER M1 ;
        RECT 9.119 0.924 9.121 3.36 ;
  LAYER M1 ;
        RECT 9.199 0.924 9.201 3.36 ;
  LAYER M1 ;
        RECT 9.279 0.924 9.281 3.36 ;
  LAYER M1 ;
        RECT 9.359 0.924 9.361 3.36 ;
  LAYER M1 ;
        RECT 9.439 0.924 9.441 3.36 ;
  LAYER M1 ;
        RECT 9.519 0.924 9.521 3.36 ;
  LAYER M1 ;
        RECT 9.599 0.924 9.601 3.36 ;
  LAYER M1 ;
        RECT 9.679 0.924 9.681 3.36 ;
  LAYER M1 ;
        RECT 9.759 0.924 9.761 3.36 ;
  LAYER M1 ;
        RECT 9.839 0.924 9.841 3.36 ;
  LAYER M1 ;
        RECT 9.919 0.924 9.921 3.36 ;
  LAYER M1 ;
        RECT 9.999 0.924 10.001 3.36 ;
  LAYER M1 ;
        RECT 10.079 0.924 10.081 3.36 ;
  LAYER M1 ;
        RECT 10.159 0.924 10.161 3.36 ;
  LAYER M1 ;
        RECT 10.239 0.924 10.241 3.36 ;
  LAYER M1 ;
        RECT 10.319 0.924 10.321 3.36 ;
  LAYER M1 ;
        RECT 10.399 0.924 10.401 3.36 ;
  LAYER M1 ;
        RECT 10.479 0.924 10.481 3.36 ;
  LAYER M1 ;
        RECT 10.559 0.924 10.561 3.36 ;
  LAYER M1 ;
        RECT 10.639 0.924 10.641 3.36 ;
  LAYER M1 ;
        RECT 10.719 0.924 10.721 3.36 ;
  LAYER M1 ;
        RECT 10.799 0.924 10.801 3.36 ;
  LAYER M1 ;
        RECT 10.879 0.924 10.881 3.36 ;
  LAYER M1 ;
        RECT 10.959 0.924 10.961 3.36 ;
  LAYER M1 ;
        RECT 11.039 0.924 11.041 3.36 ;
  LAYER M1 ;
        RECT 11.119 0.924 11.121 3.36 ;
  LAYER M1 ;
        RECT 11.199 0.924 11.201 3.36 ;
  LAYER M1 ;
        RECT 11.279 0.924 11.281 3.36 ;
  LAYER M1 ;
        RECT 11.359 0.924 11.361 3.36 ;
  LAYER M2 ;
        RECT 9.04 0.923 11.44 0.925 ;
  LAYER M2 ;
        RECT 9.04 1.007 11.44 1.009 ;
  LAYER M2 ;
        RECT 9.04 1.091 11.44 1.093 ;
  LAYER M2 ;
        RECT 9.04 1.175 11.44 1.177 ;
  LAYER M2 ;
        RECT 9.04 1.259 11.44 1.261 ;
  LAYER M2 ;
        RECT 9.04 1.343 11.44 1.345 ;
  LAYER M2 ;
        RECT 9.04 1.427 11.44 1.429 ;
  LAYER M2 ;
        RECT 9.04 1.511 11.44 1.513 ;
  LAYER M2 ;
        RECT 9.04 1.595 11.44 1.597 ;
  LAYER M2 ;
        RECT 9.04 1.679 11.44 1.681 ;
  LAYER M2 ;
        RECT 9.04 1.763 11.44 1.765 ;
  LAYER M2 ;
        RECT 9.04 1.847 11.44 1.849 ;
  LAYER M2 ;
        RECT 9.04 1.9305 11.44 1.9325 ;
  LAYER M2 ;
        RECT 9.04 2.015 11.44 2.017 ;
  LAYER M2 ;
        RECT 9.04 2.099 11.44 2.101 ;
  LAYER M2 ;
        RECT 9.04 2.183 11.44 2.185 ;
  LAYER M2 ;
        RECT 9.04 2.267 11.44 2.269 ;
  LAYER M2 ;
        RECT 9.04 2.351 11.44 2.353 ;
  LAYER M2 ;
        RECT 9.04 2.435 11.44 2.437 ;
  LAYER M2 ;
        RECT 9.04 2.519 11.44 2.521 ;
  LAYER M2 ;
        RECT 9.04 2.603 11.44 2.605 ;
  LAYER M2 ;
        RECT 9.04 2.687 11.44 2.689 ;
  LAYER M2 ;
        RECT 9.04 2.771 11.44 2.773 ;
  LAYER M2 ;
        RECT 9.04 2.855 11.44 2.857 ;
  LAYER M2 ;
        RECT 9.04 2.939 11.44 2.941 ;
  LAYER M2 ;
        RECT 9.04 3.023 11.44 3.025 ;
  LAYER M2 ;
        RECT 9.04 3.107 11.44 3.109 ;
  LAYER M2 ;
        RECT 9.04 3.191 11.44 3.193 ;
  LAYER M2 ;
        RECT 9.04 3.275 11.44 3.277 ;
  LAYER M1 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M1 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M1 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M1 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M1 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M1 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M1 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M1 ;
        RECT 9.472 3.828 9.504 6.336 ;
  LAYER M1 ;
        RECT 9.536 3.828 9.568 6.336 ;
  LAYER M1 ;
        RECT 9.6 3.828 9.632 6.336 ;
  LAYER M1 ;
        RECT 9.664 3.828 9.696 6.336 ;
  LAYER M1 ;
        RECT 9.728 3.828 9.76 6.336 ;
  LAYER M1 ;
        RECT 9.792 3.828 9.824 6.336 ;
  LAYER M1 ;
        RECT 9.856 3.828 9.888 6.336 ;
  LAYER M1 ;
        RECT 9.92 3.828 9.952 6.336 ;
  LAYER M1 ;
        RECT 9.984 3.828 10.016 6.336 ;
  LAYER M1 ;
        RECT 10.048 3.828 10.08 6.336 ;
  LAYER M1 ;
        RECT 10.112 3.828 10.144 6.336 ;
  LAYER M1 ;
        RECT 10.176 3.828 10.208 6.336 ;
  LAYER M1 ;
        RECT 10.24 3.828 10.272 6.336 ;
  LAYER M1 ;
        RECT 10.304 3.828 10.336 6.336 ;
  LAYER M1 ;
        RECT 10.368 3.828 10.4 6.336 ;
  LAYER M1 ;
        RECT 10.432 3.828 10.464 6.336 ;
  LAYER M1 ;
        RECT 10.496 3.828 10.528 6.336 ;
  LAYER M1 ;
        RECT 10.56 3.828 10.592 6.336 ;
  LAYER M1 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M1 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M1 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M1 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M1 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M1 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M1 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M1 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M1 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M1 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M1 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M1 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M2 ;
        RECT 9.004 3.912 11.476 3.944 ;
  LAYER M2 ;
        RECT 9.004 3.976 11.476 4.008 ;
  LAYER M2 ;
        RECT 9.004 4.04 11.476 4.072 ;
  LAYER M2 ;
        RECT 9.004 4.104 11.476 4.136 ;
  LAYER M2 ;
        RECT 9.004 4.168 11.476 4.2 ;
  LAYER M2 ;
        RECT 9.004 4.232 11.476 4.264 ;
  LAYER M2 ;
        RECT 9.004 4.296 11.476 4.328 ;
  LAYER M2 ;
        RECT 9.004 4.36 11.476 4.392 ;
  LAYER M2 ;
        RECT 9.004 4.424 11.476 4.456 ;
  LAYER M2 ;
        RECT 9.004 4.488 11.476 4.52 ;
  LAYER M2 ;
        RECT 9.004 4.552 11.476 4.584 ;
  LAYER M2 ;
        RECT 9.004 4.616 11.476 4.648 ;
  LAYER M2 ;
        RECT 9.004 4.68 11.476 4.712 ;
  LAYER M2 ;
        RECT 9.004 4.744 11.476 4.776 ;
  LAYER M2 ;
        RECT 9.004 4.808 11.476 4.84 ;
  LAYER M2 ;
        RECT 9.004 4.872 11.476 4.904 ;
  LAYER M2 ;
        RECT 9.004 4.936 11.476 4.968 ;
  LAYER M2 ;
        RECT 9.004 5 11.476 5.032 ;
  LAYER M2 ;
        RECT 9.004 5.064 11.476 5.096 ;
  LAYER M2 ;
        RECT 9.004 5.128 11.476 5.16 ;
  LAYER M2 ;
        RECT 9.004 5.192 11.476 5.224 ;
  LAYER M2 ;
        RECT 9.004 5.256 11.476 5.288 ;
  LAYER M2 ;
        RECT 9.004 5.32 11.476 5.352 ;
  LAYER M2 ;
        RECT 9.004 5.384 11.476 5.416 ;
  LAYER M2 ;
        RECT 9.004 5.448 11.476 5.48 ;
  LAYER M2 ;
        RECT 9.004 5.512 11.476 5.544 ;
  LAYER M2 ;
        RECT 9.004 5.576 11.476 5.608 ;
  LAYER M2 ;
        RECT 9.004 5.64 11.476 5.672 ;
  LAYER M2 ;
        RECT 9.004 5.704 11.476 5.736 ;
  LAYER M2 ;
        RECT 9.004 5.768 11.476 5.8 ;
  LAYER M2 ;
        RECT 9.004 5.832 11.476 5.864 ;
  LAYER M2 ;
        RECT 9.004 5.896 11.476 5.928 ;
  LAYER M2 ;
        RECT 9.004 5.96 11.476 5.992 ;
  LAYER M2 ;
        RECT 9.004 6.024 11.476 6.056 ;
  LAYER M2 ;
        RECT 9.004 6.088 11.476 6.12 ;
  LAYER M2 ;
        RECT 9.004 6.152 11.476 6.184 ;
  LAYER M3 ;
        RECT 9.024 3.828 9.056 6.336 ;
  LAYER M3 ;
        RECT 9.088 3.828 9.12 6.336 ;
  LAYER M3 ;
        RECT 9.152 3.828 9.184 6.336 ;
  LAYER M3 ;
        RECT 9.216 3.828 9.248 6.336 ;
  LAYER M3 ;
        RECT 9.28 3.828 9.312 6.336 ;
  LAYER M3 ;
        RECT 9.344 3.828 9.376 6.336 ;
  LAYER M3 ;
        RECT 9.408 3.828 9.44 6.336 ;
  LAYER M3 ;
        RECT 9.472 3.828 9.504 6.336 ;
  LAYER M3 ;
        RECT 9.536 3.828 9.568 6.336 ;
  LAYER M3 ;
        RECT 9.6 3.828 9.632 6.336 ;
  LAYER M3 ;
        RECT 9.664 3.828 9.696 6.336 ;
  LAYER M3 ;
        RECT 9.728 3.828 9.76 6.336 ;
  LAYER M3 ;
        RECT 9.792 3.828 9.824 6.336 ;
  LAYER M3 ;
        RECT 9.856 3.828 9.888 6.336 ;
  LAYER M3 ;
        RECT 9.92 3.828 9.952 6.336 ;
  LAYER M3 ;
        RECT 9.984 3.828 10.016 6.336 ;
  LAYER M3 ;
        RECT 10.048 3.828 10.08 6.336 ;
  LAYER M3 ;
        RECT 10.112 3.828 10.144 6.336 ;
  LAYER M3 ;
        RECT 10.176 3.828 10.208 6.336 ;
  LAYER M3 ;
        RECT 10.24 3.828 10.272 6.336 ;
  LAYER M3 ;
        RECT 10.304 3.828 10.336 6.336 ;
  LAYER M3 ;
        RECT 10.368 3.828 10.4 6.336 ;
  LAYER M3 ;
        RECT 10.432 3.828 10.464 6.336 ;
  LAYER M3 ;
        RECT 10.496 3.828 10.528 6.336 ;
  LAYER M3 ;
        RECT 10.56 3.828 10.592 6.336 ;
  LAYER M3 ;
        RECT 10.624 3.828 10.656 6.336 ;
  LAYER M3 ;
        RECT 10.688 3.828 10.72 6.336 ;
  LAYER M3 ;
        RECT 10.752 3.828 10.784 6.336 ;
  LAYER M3 ;
        RECT 10.816 3.828 10.848 6.336 ;
  LAYER M3 ;
        RECT 10.88 3.828 10.912 6.336 ;
  LAYER M3 ;
        RECT 10.944 3.828 10.976 6.336 ;
  LAYER M3 ;
        RECT 11.008 3.828 11.04 6.336 ;
  LAYER M3 ;
        RECT 11.072 3.828 11.104 6.336 ;
  LAYER M3 ;
        RECT 11.136 3.828 11.168 6.336 ;
  LAYER M3 ;
        RECT 11.2 3.828 11.232 6.336 ;
  LAYER M3 ;
        RECT 11.264 3.828 11.296 6.336 ;
  LAYER M3 ;
        RECT 11.328 3.828 11.36 6.336 ;
  LAYER M3 ;
        RECT 11.424 3.828 11.456 6.336 ;
  LAYER M1 ;
        RECT 9.039 3.864 9.041 6.3 ;
  LAYER M1 ;
        RECT 9.119 3.864 9.121 6.3 ;
  LAYER M1 ;
        RECT 9.199 3.864 9.201 6.3 ;
  LAYER M1 ;
        RECT 9.279 3.864 9.281 6.3 ;
  LAYER M1 ;
        RECT 9.359 3.864 9.361 6.3 ;
  LAYER M1 ;
        RECT 9.439 3.864 9.441 6.3 ;
  LAYER M1 ;
        RECT 9.519 3.864 9.521 6.3 ;
  LAYER M1 ;
        RECT 9.599 3.864 9.601 6.3 ;
  LAYER M1 ;
        RECT 9.679 3.864 9.681 6.3 ;
  LAYER M1 ;
        RECT 9.759 3.864 9.761 6.3 ;
  LAYER M1 ;
        RECT 9.839 3.864 9.841 6.3 ;
  LAYER M1 ;
        RECT 9.919 3.864 9.921 6.3 ;
  LAYER M1 ;
        RECT 9.999 3.864 10.001 6.3 ;
  LAYER M1 ;
        RECT 10.079 3.864 10.081 6.3 ;
  LAYER M1 ;
        RECT 10.159 3.864 10.161 6.3 ;
  LAYER M1 ;
        RECT 10.239 3.864 10.241 6.3 ;
  LAYER M1 ;
        RECT 10.319 3.864 10.321 6.3 ;
  LAYER M1 ;
        RECT 10.399 3.864 10.401 6.3 ;
  LAYER M1 ;
        RECT 10.479 3.864 10.481 6.3 ;
  LAYER M1 ;
        RECT 10.559 3.864 10.561 6.3 ;
  LAYER M1 ;
        RECT 10.639 3.864 10.641 6.3 ;
  LAYER M1 ;
        RECT 10.719 3.864 10.721 6.3 ;
  LAYER M1 ;
        RECT 10.799 3.864 10.801 6.3 ;
  LAYER M1 ;
        RECT 10.879 3.864 10.881 6.3 ;
  LAYER M1 ;
        RECT 10.959 3.864 10.961 6.3 ;
  LAYER M1 ;
        RECT 11.039 3.864 11.041 6.3 ;
  LAYER M1 ;
        RECT 11.119 3.864 11.121 6.3 ;
  LAYER M1 ;
        RECT 11.199 3.864 11.201 6.3 ;
  LAYER M1 ;
        RECT 11.279 3.864 11.281 6.3 ;
  LAYER M1 ;
        RECT 11.359 3.864 11.361 6.3 ;
  LAYER M2 ;
        RECT 9.04 3.863 11.44 3.865 ;
  LAYER M2 ;
        RECT 9.04 3.947 11.44 3.949 ;
  LAYER M2 ;
        RECT 9.04 4.031 11.44 4.033 ;
  LAYER M2 ;
        RECT 9.04 4.115 11.44 4.117 ;
  LAYER M2 ;
        RECT 9.04 4.199 11.44 4.201 ;
  LAYER M2 ;
        RECT 9.04 4.283 11.44 4.285 ;
  LAYER M2 ;
        RECT 9.04 4.367 11.44 4.369 ;
  LAYER M2 ;
        RECT 9.04 4.451 11.44 4.453 ;
  LAYER M2 ;
        RECT 9.04 4.535 11.44 4.537 ;
  LAYER M2 ;
        RECT 9.04 4.619 11.44 4.621 ;
  LAYER M2 ;
        RECT 9.04 4.703 11.44 4.705 ;
  LAYER M2 ;
        RECT 9.04 4.787 11.44 4.789 ;
  LAYER M2 ;
        RECT 9.04 4.8705 11.44 4.8725 ;
  LAYER M2 ;
        RECT 9.04 4.955 11.44 4.957 ;
  LAYER M2 ;
        RECT 9.04 5.039 11.44 5.041 ;
  LAYER M2 ;
        RECT 9.04 5.123 11.44 5.125 ;
  LAYER M2 ;
        RECT 9.04 5.207 11.44 5.209 ;
  LAYER M2 ;
        RECT 9.04 5.291 11.44 5.293 ;
  LAYER M2 ;
        RECT 9.04 5.375 11.44 5.377 ;
  LAYER M2 ;
        RECT 9.04 5.459 11.44 5.461 ;
  LAYER M2 ;
        RECT 9.04 5.543 11.44 5.545 ;
  LAYER M2 ;
        RECT 9.04 5.627 11.44 5.629 ;
  LAYER M2 ;
        RECT 9.04 5.711 11.44 5.713 ;
  LAYER M2 ;
        RECT 9.04 5.795 11.44 5.797 ;
  LAYER M2 ;
        RECT 9.04 5.879 11.44 5.881 ;
  LAYER M2 ;
        RECT 9.04 5.963 11.44 5.965 ;
  LAYER M2 ;
        RECT 9.04 6.047 11.44 6.049 ;
  LAYER M2 ;
        RECT 9.04 6.131 11.44 6.133 ;
  LAYER M2 ;
        RECT 9.04 6.215 11.44 6.217 ;
  LAYER M1 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M1 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M1 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M1 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M1 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M1 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M1 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M1 ;
        RECT 9.472 6.768 9.504 9.276 ;
  LAYER M1 ;
        RECT 9.536 6.768 9.568 9.276 ;
  LAYER M1 ;
        RECT 9.6 6.768 9.632 9.276 ;
  LAYER M1 ;
        RECT 9.664 6.768 9.696 9.276 ;
  LAYER M1 ;
        RECT 9.728 6.768 9.76 9.276 ;
  LAYER M1 ;
        RECT 9.792 6.768 9.824 9.276 ;
  LAYER M1 ;
        RECT 9.856 6.768 9.888 9.276 ;
  LAYER M1 ;
        RECT 9.92 6.768 9.952 9.276 ;
  LAYER M1 ;
        RECT 9.984 6.768 10.016 9.276 ;
  LAYER M1 ;
        RECT 10.048 6.768 10.08 9.276 ;
  LAYER M1 ;
        RECT 10.112 6.768 10.144 9.276 ;
  LAYER M1 ;
        RECT 10.176 6.768 10.208 9.276 ;
  LAYER M1 ;
        RECT 10.24 6.768 10.272 9.276 ;
  LAYER M1 ;
        RECT 10.304 6.768 10.336 9.276 ;
  LAYER M1 ;
        RECT 10.368 6.768 10.4 9.276 ;
  LAYER M1 ;
        RECT 10.432 6.768 10.464 9.276 ;
  LAYER M1 ;
        RECT 10.496 6.768 10.528 9.276 ;
  LAYER M1 ;
        RECT 10.56 6.768 10.592 9.276 ;
  LAYER M1 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M1 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M1 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M1 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M1 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M1 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M1 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M1 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M1 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M1 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M1 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M1 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M2 ;
        RECT 9.004 6.852 11.476 6.884 ;
  LAYER M2 ;
        RECT 9.004 6.916 11.476 6.948 ;
  LAYER M2 ;
        RECT 9.004 6.98 11.476 7.012 ;
  LAYER M2 ;
        RECT 9.004 7.044 11.476 7.076 ;
  LAYER M2 ;
        RECT 9.004 7.108 11.476 7.14 ;
  LAYER M2 ;
        RECT 9.004 7.172 11.476 7.204 ;
  LAYER M2 ;
        RECT 9.004 7.236 11.476 7.268 ;
  LAYER M2 ;
        RECT 9.004 7.3 11.476 7.332 ;
  LAYER M2 ;
        RECT 9.004 7.364 11.476 7.396 ;
  LAYER M2 ;
        RECT 9.004 7.428 11.476 7.46 ;
  LAYER M2 ;
        RECT 9.004 7.492 11.476 7.524 ;
  LAYER M2 ;
        RECT 9.004 7.556 11.476 7.588 ;
  LAYER M2 ;
        RECT 9.004 7.62 11.476 7.652 ;
  LAYER M2 ;
        RECT 9.004 7.684 11.476 7.716 ;
  LAYER M2 ;
        RECT 9.004 7.748 11.476 7.78 ;
  LAYER M2 ;
        RECT 9.004 7.812 11.476 7.844 ;
  LAYER M2 ;
        RECT 9.004 7.876 11.476 7.908 ;
  LAYER M2 ;
        RECT 9.004 7.94 11.476 7.972 ;
  LAYER M2 ;
        RECT 9.004 8.004 11.476 8.036 ;
  LAYER M2 ;
        RECT 9.004 8.068 11.476 8.1 ;
  LAYER M2 ;
        RECT 9.004 8.132 11.476 8.164 ;
  LAYER M2 ;
        RECT 9.004 8.196 11.476 8.228 ;
  LAYER M2 ;
        RECT 9.004 8.26 11.476 8.292 ;
  LAYER M2 ;
        RECT 9.004 8.324 11.476 8.356 ;
  LAYER M2 ;
        RECT 9.004 8.388 11.476 8.42 ;
  LAYER M2 ;
        RECT 9.004 8.452 11.476 8.484 ;
  LAYER M2 ;
        RECT 9.004 8.516 11.476 8.548 ;
  LAYER M2 ;
        RECT 9.004 8.58 11.476 8.612 ;
  LAYER M2 ;
        RECT 9.004 8.644 11.476 8.676 ;
  LAYER M2 ;
        RECT 9.004 8.708 11.476 8.74 ;
  LAYER M2 ;
        RECT 9.004 8.772 11.476 8.804 ;
  LAYER M2 ;
        RECT 9.004 8.836 11.476 8.868 ;
  LAYER M2 ;
        RECT 9.004 8.9 11.476 8.932 ;
  LAYER M2 ;
        RECT 9.004 8.964 11.476 8.996 ;
  LAYER M2 ;
        RECT 9.004 9.028 11.476 9.06 ;
  LAYER M2 ;
        RECT 9.004 9.092 11.476 9.124 ;
  LAYER M3 ;
        RECT 9.024 6.768 9.056 9.276 ;
  LAYER M3 ;
        RECT 9.088 6.768 9.12 9.276 ;
  LAYER M3 ;
        RECT 9.152 6.768 9.184 9.276 ;
  LAYER M3 ;
        RECT 9.216 6.768 9.248 9.276 ;
  LAYER M3 ;
        RECT 9.28 6.768 9.312 9.276 ;
  LAYER M3 ;
        RECT 9.344 6.768 9.376 9.276 ;
  LAYER M3 ;
        RECT 9.408 6.768 9.44 9.276 ;
  LAYER M3 ;
        RECT 9.472 6.768 9.504 9.276 ;
  LAYER M3 ;
        RECT 9.536 6.768 9.568 9.276 ;
  LAYER M3 ;
        RECT 9.6 6.768 9.632 9.276 ;
  LAYER M3 ;
        RECT 9.664 6.768 9.696 9.276 ;
  LAYER M3 ;
        RECT 9.728 6.768 9.76 9.276 ;
  LAYER M3 ;
        RECT 9.792 6.768 9.824 9.276 ;
  LAYER M3 ;
        RECT 9.856 6.768 9.888 9.276 ;
  LAYER M3 ;
        RECT 9.92 6.768 9.952 9.276 ;
  LAYER M3 ;
        RECT 9.984 6.768 10.016 9.276 ;
  LAYER M3 ;
        RECT 10.048 6.768 10.08 9.276 ;
  LAYER M3 ;
        RECT 10.112 6.768 10.144 9.276 ;
  LAYER M3 ;
        RECT 10.176 6.768 10.208 9.276 ;
  LAYER M3 ;
        RECT 10.24 6.768 10.272 9.276 ;
  LAYER M3 ;
        RECT 10.304 6.768 10.336 9.276 ;
  LAYER M3 ;
        RECT 10.368 6.768 10.4 9.276 ;
  LAYER M3 ;
        RECT 10.432 6.768 10.464 9.276 ;
  LAYER M3 ;
        RECT 10.496 6.768 10.528 9.276 ;
  LAYER M3 ;
        RECT 10.56 6.768 10.592 9.276 ;
  LAYER M3 ;
        RECT 10.624 6.768 10.656 9.276 ;
  LAYER M3 ;
        RECT 10.688 6.768 10.72 9.276 ;
  LAYER M3 ;
        RECT 10.752 6.768 10.784 9.276 ;
  LAYER M3 ;
        RECT 10.816 6.768 10.848 9.276 ;
  LAYER M3 ;
        RECT 10.88 6.768 10.912 9.276 ;
  LAYER M3 ;
        RECT 10.944 6.768 10.976 9.276 ;
  LAYER M3 ;
        RECT 11.008 6.768 11.04 9.276 ;
  LAYER M3 ;
        RECT 11.072 6.768 11.104 9.276 ;
  LAYER M3 ;
        RECT 11.136 6.768 11.168 9.276 ;
  LAYER M3 ;
        RECT 11.2 6.768 11.232 9.276 ;
  LAYER M3 ;
        RECT 11.264 6.768 11.296 9.276 ;
  LAYER M3 ;
        RECT 11.328 6.768 11.36 9.276 ;
  LAYER M3 ;
        RECT 11.424 6.768 11.456 9.276 ;
  LAYER M1 ;
        RECT 9.039 6.804 9.041 9.24 ;
  LAYER M1 ;
        RECT 9.119 6.804 9.121 9.24 ;
  LAYER M1 ;
        RECT 9.199 6.804 9.201 9.24 ;
  LAYER M1 ;
        RECT 9.279 6.804 9.281 9.24 ;
  LAYER M1 ;
        RECT 9.359 6.804 9.361 9.24 ;
  LAYER M1 ;
        RECT 9.439 6.804 9.441 9.24 ;
  LAYER M1 ;
        RECT 9.519 6.804 9.521 9.24 ;
  LAYER M1 ;
        RECT 9.599 6.804 9.601 9.24 ;
  LAYER M1 ;
        RECT 9.679 6.804 9.681 9.24 ;
  LAYER M1 ;
        RECT 9.759 6.804 9.761 9.24 ;
  LAYER M1 ;
        RECT 9.839 6.804 9.841 9.24 ;
  LAYER M1 ;
        RECT 9.919 6.804 9.921 9.24 ;
  LAYER M1 ;
        RECT 9.999 6.804 10.001 9.24 ;
  LAYER M1 ;
        RECT 10.079 6.804 10.081 9.24 ;
  LAYER M1 ;
        RECT 10.159 6.804 10.161 9.24 ;
  LAYER M1 ;
        RECT 10.239 6.804 10.241 9.24 ;
  LAYER M1 ;
        RECT 10.319 6.804 10.321 9.24 ;
  LAYER M1 ;
        RECT 10.399 6.804 10.401 9.24 ;
  LAYER M1 ;
        RECT 10.479 6.804 10.481 9.24 ;
  LAYER M1 ;
        RECT 10.559 6.804 10.561 9.24 ;
  LAYER M1 ;
        RECT 10.639 6.804 10.641 9.24 ;
  LAYER M1 ;
        RECT 10.719 6.804 10.721 9.24 ;
  LAYER M1 ;
        RECT 10.799 6.804 10.801 9.24 ;
  LAYER M1 ;
        RECT 10.879 6.804 10.881 9.24 ;
  LAYER M1 ;
        RECT 10.959 6.804 10.961 9.24 ;
  LAYER M1 ;
        RECT 11.039 6.804 11.041 9.24 ;
  LAYER M1 ;
        RECT 11.119 6.804 11.121 9.24 ;
  LAYER M1 ;
        RECT 11.199 6.804 11.201 9.24 ;
  LAYER M1 ;
        RECT 11.279 6.804 11.281 9.24 ;
  LAYER M1 ;
        RECT 11.359 6.804 11.361 9.24 ;
  LAYER M2 ;
        RECT 9.04 6.803 11.44 6.805 ;
  LAYER M2 ;
        RECT 9.04 6.887 11.44 6.889 ;
  LAYER M2 ;
        RECT 9.04 6.971 11.44 6.973 ;
  LAYER M2 ;
        RECT 9.04 7.055 11.44 7.057 ;
  LAYER M2 ;
        RECT 9.04 7.139 11.44 7.141 ;
  LAYER M2 ;
        RECT 9.04 7.223 11.44 7.225 ;
  LAYER M2 ;
        RECT 9.04 7.307 11.44 7.309 ;
  LAYER M2 ;
        RECT 9.04 7.391 11.44 7.393 ;
  LAYER M2 ;
        RECT 9.04 7.475 11.44 7.477 ;
  LAYER M2 ;
        RECT 9.04 7.559 11.44 7.561 ;
  LAYER M2 ;
        RECT 9.04 7.643 11.44 7.645 ;
  LAYER M2 ;
        RECT 9.04 7.727 11.44 7.729 ;
  LAYER M2 ;
        RECT 9.04 7.8105 11.44 7.8125 ;
  LAYER M2 ;
        RECT 9.04 7.895 11.44 7.897 ;
  LAYER M2 ;
        RECT 9.04 7.979 11.44 7.981 ;
  LAYER M2 ;
        RECT 9.04 8.063 11.44 8.065 ;
  LAYER M2 ;
        RECT 9.04 8.147 11.44 8.149 ;
  LAYER M2 ;
        RECT 9.04 8.231 11.44 8.233 ;
  LAYER M2 ;
        RECT 9.04 8.315 11.44 8.317 ;
  LAYER M2 ;
        RECT 9.04 8.399 11.44 8.401 ;
  LAYER M2 ;
        RECT 9.04 8.483 11.44 8.485 ;
  LAYER M2 ;
        RECT 9.04 8.567 11.44 8.569 ;
  LAYER M2 ;
        RECT 9.04 8.651 11.44 8.653 ;
  LAYER M2 ;
        RECT 9.04 8.735 11.44 8.737 ;
  LAYER M2 ;
        RECT 9.04 8.819 11.44 8.821 ;
  LAYER M2 ;
        RECT 9.04 8.903 11.44 8.905 ;
  LAYER M2 ;
        RECT 9.04 8.987 11.44 8.989 ;
  LAYER M2 ;
        RECT 9.04 9.071 11.44 9.073 ;
  LAYER M2 ;
        RECT 9.04 9.155 11.44 9.157 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M1 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M1 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M1 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M1 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M1 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M1 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M1 ;
        RECT 9.472 9.708 9.504 12.216 ;
  LAYER M1 ;
        RECT 9.536 9.708 9.568 12.216 ;
  LAYER M1 ;
        RECT 9.6 9.708 9.632 12.216 ;
  LAYER M1 ;
        RECT 9.664 9.708 9.696 12.216 ;
  LAYER M1 ;
        RECT 9.728 9.708 9.76 12.216 ;
  LAYER M1 ;
        RECT 9.792 9.708 9.824 12.216 ;
  LAYER M1 ;
        RECT 9.856 9.708 9.888 12.216 ;
  LAYER M1 ;
        RECT 9.92 9.708 9.952 12.216 ;
  LAYER M1 ;
        RECT 9.984 9.708 10.016 12.216 ;
  LAYER M1 ;
        RECT 10.048 9.708 10.08 12.216 ;
  LAYER M1 ;
        RECT 10.112 9.708 10.144 12.216 ;
  LAYER M1 ;
        RECT 10.176 9.708 10.208 12.216 ;
  LAYER M1 ;
        RECT 10.24 9.708 10.272 12.216 ;
  LAYER M1 ;
        RECT 10.304 9.708 10.336 12.216 ;
  LAYER M1 ;
        RECT 10.368 9.708 10.4 12.216 ;
  LAYER M1 ;
        RECT 10.432 9.708 10.464 12.216 ;
  LAYER M1 ;
        RECT 10.496 9.708 10.528 12.216 ;
  LAYER M1 ;
        RECT 10.56 9.708 10.592 12.216 ;
  LAYER M1 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M1 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M1 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M1 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M1 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M1 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M1 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M1 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M1 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M1 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M1 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M1 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M2 ;
        RECT 9.004 9.792 11.476 9.824 ;
  LAYER M2 ;
        RECT 9.004 9.856 11.476 9.888 ;
  LAYER M2 ;
        RECT 9.004 9.92 11.476 9.952 ;
  LAYER M2 ;
        RECT 9.004 9.984 11.476 10.016 ;
  LAYER M2 ;
        RECT 9.004 10.048 11.476 10.08 ;
  LAYER M2 ;
        RECT 9.004 10.112 11.476 10.144 ;
  LAYER M2 ;
        RECT 9.004 10.176 11.476 10.208 ;
  LAYER M2 ;
        RECT 9.004 10.24 11.476 10.272 ;
  LAYER M2 ;
        RECT 9.004 10.304 11.476 10.336 ;
  LAYER M2 ;
        RECT 9.004 10.368 11.476 10.4 ;
  LAYER M2 ;
        RECT 9.004 10.432 11.476 10.464 ;
  LAYER M2 ;
        RECT 9.004 10.496 11.476 10.528 ;
  LAYER M2 ;
        RECT 9.004 10.56 11.476 10.592 ;
  LAYER M2 ;
        RECT 9.004 10.624 11.476 10.656 ;
  LAYER M2 ;
        RECT 9.004 10.688 11.476 10.72 ;
  LAYER M2 ;
        RECT 9.004 10.752 11.476 10.784 ;
  LAYER M2 ;
        RECT 9.004 10.816 11.476 10.848 ;
  LAYER M2 ;
        RECT 9.004 10.88 11.476 10.912 ;
  LAYER M2 ;
        RECT 9.004 10.944 11.476 10.976 ;
  LAYER M2 ;
        RECT 9.004 11.008 11.476 11.04 ;
  LAYER M2 ;
        RECT 9.004 11.072 11.476 11.104 ;
  LAYER M2 ;
        RECT 9.004 11.136 11.476 11.168 ;
  LAYER M2 ;
        RECT 9.004 11.2 11.476 11.232 ;
  LAYER M2 ;
        RECT 9.004 11.264 11.476 11.296 ;
  LAYER M2 ;
        RECT 9.004 11.328 11.476 11.36 ;
  LAYER M2 ;
        RECT 9.004 11.392 11.476 11.424 ;
  LAYER M2 ;
        RECT 9.004 11.456 11.476 11.488 ;
  LAYER M2 ;
        RECT 9.004 11.52 11.476 11.552 ;
  LAYER M2 ;
        RECT 9.004 11.584 11.476 11.616 ;
  LAYER M2 ;
        RECT 9.004 11.648 11.476 11.68 ;
  LAYER M2 ;
        RECT 9.004 11.712 11.476 11.744 ;
  LAYER M2 ;
        RECT 9.004 11.776 11.476 11.808 ;
  LAYER M2 ;
        RECT 9.004 11.84 11.476 11.872 ;
  LAYER M2 ;
        RECT 9.004 11.904 11.476 11.936 ;
  LAYER M2 ;
        RECT 9.004 11.968 11.476 12 ;
  LAYER M2 ;
        RECT 9.004 12.032 11.476 12.064 ;
  LAYER M3 ;
        RECT 9.024 9.708 9.056 12.216 ;
  LAYER M3 ;
        RECT 9.088 9.708 9.12 12.216 ;
  LAYER M3 ;
        RECT 9.152 9.708 9.184 12.216 ;
  LAYER M3 ;
        RECT 9.216 9.708 9.248 12.216 ;
  LAYER M3 ;
        RECT 9.28 9.708 9.312 12.216 ;
  LAYER M3 ;
        RECT 9.344 9.708 9.376 12.216 ;
  LAYER M3 ;
        RECT 9.408 9.708 9.44 12.216 ;
  LAYER M3 ;
        RECT 9.472 9.708 9.504 12.216 ;
  LAYER M3 ;
        RECT 9.536 9.708 9.568 12.216 ;
  LAYER M3 ;
        RECT 9.6 9.708 9.632 12.216 ;
  LAYER M3 ;
        RECT 9.664 9.708 9.696 12.216 ;
  LAYER M3 ;
        RECT 9.728 9.708 9.76 12.216 ;
  LAYER M3 ;
        RECT 9.792 9.708 9.824 12.216 ;
  LAYER M3 ;
        RECT 9.856 9.708 9.888 12.216 ;
  LAYER M3 ;
        RECT 9.92 9.708 9.952 12.216 ;
  LAYER M3 ;
        RECT 9.984 9.708 10.016 12.216 ;
  LAYER M3 ;
        RECT 10.048 9.708 10.08 12.216 ;
  LAYER M3 ;
        RECT 10.112 9.708 10.144 12.216 ;
  LAYER M3 ;
        RECT 10.176 9.708 10.208 12.216 ;
  LAYER M3 ;
        RECT 10.24 9.708 10.272 12.216 ;
  LAYER M3 ;
        RECT 10.304 9.708 10.336 12.216 ;
  LAYER M3 ;
        RECT 10.368 9.708 10.4 12.216 ;
  LAYER M3 ;
        RECT 10.432 9.708 10.464 12.216 ;
  LAYER M3 ;
        RECT 10.496 9.708 10.528 12.216 ;
  LAYER M3 ;
        RECT 10.56 9.708 10.592 12.216 ;
  LAYER M3 ;
        RECT 10.624 9.708 10.656 12.216 ;
  LAYER M3 ;
        RECT 10.688 9.708 10.72 12.216 ;
  LAYER M3 ;
        RECT 10.752 9.708 10.784 12.216 ;
  LAYER M3 ;
        RECT 10.816 9.708 10.848 12.216 ;
  LAYER M3 ;
        RECT 10.88 9.708 10.912 12.216 ;
  LAYER M3 ;
        RECT 10.944 9.708 10.976 12.216 ;
  LAYER M3 ;
        RECT 11.008 9.708 11.04 12.216 ;
  LAYER M3 ;
        RECT 11.072 9.708 11.104 12.216 ;
  LAYER M3 ;
        RECT 11.136 9.708 11.168 12.216 ;
  LAYER M3 ;
        RECT 11.2 9.708 11.232 12.216 ;
  LAYER M3 ;
        RECT 11.264 9.708 11.296 12.216 ;
  LAYER M3 ;
        RECT 11.328 9.708 11.36 12.216 ;
  LAYER M3 ;
        RECT 11.424 9.708 11.456 12.216 ;
  LAYER M1 ;
        RECT 9.039 9.744 9.041 12.18 ;
  LAYER M1 ;
        RECT 9.119 9.744 9.121 12.18 ;
  LAYER M1 ;
        RECT 9.199 9.744 9.201 12.18 ;
  LAYER M1 ;
        RECT 9.279 9.744 9.281 12.18 ;
  LAYER M1 ;
        RECT 9.359 9.744 9.361 12.18 ;
  LAYER M1 ;
        RECT 9.439 9.744 9.441 12.18 ;
  LAYER M1 ;
        RECT 9.519 9.744 9.521 12.18 ;
  LAYER M1 ;
        RECT 9.599 9.744 9.601 12.18 ;
  LAYER M1 ;
        RECT 9.679 9.744 9.681 12.18 ;
  LAYER M1 ;
        RECT 9.759 9.744 9.761 12.18 ;
  LAYER M1 ;
        RECT 9.839 9.744 9.841 12.18 ;
  LAYER M1 ;
        RECT 9.919 9.744 9.921 12.18 ;
  LAYER M1 ;
        RECT 9.999 9.744 10.001 12.18 ;
  LAYER M1 ;
        RECT 10.079 9.744 10.081 12.18 ;
  LAYER M1 ;
        RECT 10.159 9.744 10.161 12.18 ;
  LAYER M1 ;
        RECT 10.239 9.744 10.241 12.18 ;
  LAYER M1 ;
        RECT 10.319 9.744 10.321 12.18 ;
  LAYER M1 ;
        RECT 10.399 9.744 10.401 12.18 ;
  LAYER M1 ;
        RECT 10.479 9.744 10.481 12.18 ;
  LAYER M1 ;
        RECT 10.559 9.744 10.561 12.18 ;
  LAYER M1 ;
        RECT 10.639 9.744 10.641 12.18 ;
  LAYER M1 ;
        RECT 10.719 9.744 10.721 12.18 ;
  LAYER M1 ;
        RECT 10.799 9.744 10.801 12.18 ;
  LAYER M1 ;
        RECT 10.879 9.744 10.881 12.18 ;
  LAYER M1 ;
        RECT 10.959 9.744 10.961 12.18 ;
  LAYER M1 ;
        RECT 11.039 9.744 11.041 12.18 ;
  LAYER M1 ;
        RECT 11.119 9.744 11.121 12.18 ;
  LAYER M1 ;
        RECT 11.199 9.744 11.201 12.18 ;
  LAYER M1 ;
        RECT 11.279 9.744 11.281 12.18 ;
  LAYER M1 ;
        RECT 11.359 9.744 11.361 12.18 ;
  LAYER M2 ;
        RECT 9.04 9.743 11.44 9.745 ;
  LAYER M2 ;
        RECT 9.04 9.827 11.44 9.829 ;
  LAYER M2 ;
        RECT 9.04 9.911 11.44 9.913 ;
  LAYER M2 ;
        RECT 9.04 9.995 11.44 9.997 ;
  LAYER M2 ;
        RECT 9.04 10.079 11.44 10.081 ;
  LAYER M2 ;
        RECT 9.04 10.163 11.44 10.165 ;
  LAYER M2 ;
        RECT 9.04 10.247 11.44 10.249 ;
  LAYER M2 ;
        RECT 9.04 10.331 11.44 10.333 ;
  LAYER M2 ;
        RECT 9.04 10.415 11.44 10.417 ;
  LAYER M2 ;
        RECT 9.04 10.499 11.44 10.501 ;
  LAYER M2 ;
        RECT 9.04 10.583 11.44 10.585 ;
  LAYER M2 ;
        RECT 9.04 10.667 11.44 10.669 ;
  LAYER M2 ;
        RECT 9.04 10.7505 11.44 10.7525 ;
  LAYER M2 ;
        RECT 9.04 10.835 11.44 10.837 ;
  LAYER M2 ;
        RECT 9.04 10.919 11.44 10.921 ;
  LAYER M2 ;
        RECT 9.04 11.003 11.44 11.005 ;
  LAYER M2 ;
        RECT 9.04 11.087 11.44 11.089 ;
  LAYER M2 ;
        RECT 9.04 11.171 11.44 11.173 ;
  LAYER M2 ;
        RECT 9.04 11.255 11.44 11.257 ;
  LAYER M2 ;
        RECT 9.04 11.339 11.44 11.341 ;
  LAYER M2 ;
        RECT 9.04 11.423 11.44 11.425 ;
  LAYER M2 ;
        RECT 9.04 11.507 11.44 11.509 ;
  LAYER M2 ;
        RECT 9.04 11.591 11.44 11.593 ;
  LAYER M2 ;
        RECT 9.04 11.675 11.44 11.677 ;
  LAYER M2 ;
        RECT 9.04 11.759 11.44 11.761 ;
  LAYER M2 ;
        RECT 9.04 11.843 11.44 11.845 ;
  LAYER M2 ;
        RECT 9.04 11.927 11.44 11.929 ;
  LAYER M2 ;
        RECT 9.04 12.011 11.44 12.013 ;
  LAYER M2 ;
        RECT 9.04 12.095 11.44 12.097 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M1 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M1 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M1 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M1 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M1 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M1 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M1 ;
        RECT 9.472 12.648 9.504 15.156 ;
  LAYER M1 ;
        RECT 9.536 12.648 9.568 15.156 ;
  LAYER M1 ;
        RECT 9.6 12.648 9.632 15.156 ;
  LAYER M1 ;
        RECT 9.664 12.648 9.696 15.156 ;
  LAYER M1 ;
        RECT 9.728 12.648 9.76 15.156 ;
  LAYER M1 ;
        RECT 9.792 12.648 9.824 15.156 ;
  LAYER M1 ;
        RECT 9.856 12.648 9.888 15.156 ;
  LAYER M1 ;
        RECT 9.92 12.648 9.952 15.156 ;
  LAYER M1 ;
        RECT 9.984 12.648 10.016 15.156 ;
  LAYER M1 ;
        RECT 10.048 12.648 10.08 15.156 ;
  LAYER M1 ;
        RECT 10.112 12.648 10.144 15.156 ;
  LAYER M1 ;
        RECT 10.176 12.648 10.208 15.156 ;
  LAYER M1 ;
        RECT 10.24 12.648 10.272 15.156 ;
  LAYER M1 ;
        RECT 10.304 12.648 10.336 15.156 ;
  LAYER M1 ;
        RECT 10.368 12.648 10.4 15.156 ;
  LAYER M1 ;
        RECT 10.432 12.648 10.464 15.156 ;
  LAYER M1 ;
        RECT 10.496 12.648 10.528 15.156 ;
  LAYER M1 ;
        RECT 10.56 12.648 10.592 15.156 ;
  LAYER M1 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M1 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M1 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M1 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M1 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M1 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M1 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M1 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M1 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M1 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M1 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M1 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M2 ;
        RECT 9.004 12.732 11.476 12.764 ;
  LAYER M2 ;
        RECT 9.004 12.796 11.476 12.828 ;
  LAYER M2 ;
        RECT 9.004 12.86 11.476 12.892 ;
  LAYER M2 ;
        RECT 9.004 12.924 11.476 12.956 ;
  LAYER M2 ;
        RECT 9.004 12.988 11.476 13.02 ;
  LAYER M2 ;
        RECT 9.004 13.052 11.476 13.084 ;
  LAYER M2 ;
        RECT 9.004 13.116 11.476 13.148 ;
  LAYER M2 ;
        RECT 9.004 13.18 11.476 13.212 ;
  LAYER M2 ;
        RECT 9.004 13.244 11.476 13.276 ;
  LAYER M2 ;
        RECT 9.004 13.308 11.476 13.34 ;
  LAYER M2 ;
        RECT 9.004 13.372 11.476 13.404 ;
  LAYER M2 ;
        RECT 9.004 13.436 11.476 13.468 ;
  LAYER M2 ;
        RECT 9.004 13.5 11.476 13.532 ;
  LAYER M2 ;
        RECT 9.004 13.564 11.476 13.596 ;
  LAYER M2 ;
        RECT 9.004 13.628 11.476 13.66 ;
  LAYER M2 ;
        RECT 9.004 13.692 11.476 13.724 ;
  LAYER M2 ;
        RECT 9.004 13.756 11.476 13.788 ;
  LAYER M2 ;
        RECT 9.004 13.82 11.476 13.852 ;
  LAYER M2 ;
        RECT 9.004 13.884 11.476 13.916 ;
  LAYER M2 ;
        RECT 9.004 13.948 11.476 13.98 ;
  LAYER M2 ;
        RECT 9.004 14.012 11.476 14.044 ;
  LAYER M2 ;
        RECT 9.004 14.076 11.476 14.108 ;
  LAYER M2 ;
        RECT 9.004 14.14 11.476 14.172 ;
  LAYER M2 ;
        RECT 9.004 14.204 11.476 14.236 ;
  LAYER M2 ;
        RECT 9.004 14.268 11.476 14.3 ;
  LAYER M2 ;
        RECT 9.004 14.332 11.476 14.364 ;
  LAYER M2 ;
        RECT 9.004 14.396 11.476 14.428 ;
  LAYER M2 ;
        RECT 9.004 14.46 11.476 14.492 ;
  LAYER M2 ;
        RECT 9.004 14.524 11.476 14.556 ;
  LAYER M2 ;
        RECT 9.004 14.588 11.476 14.62 ;
  LAYER M2 ;
        RECT 9.004 14.652 11.476 14.684 ;
  LAYER M2 ;
        RECT 9.004 14.716 11.476 14.748 ;
  LAYER M2 ;
        RECT 9.004 14.78 11.476 14.812 ;
  LAYER M2 ;
        RECT 9.004 14.844 11.476 14.876 ;
  LAYER M2 ;
        RECT 9.004 14.908 11.476 14.94 ;
  LAYER M2 ;
        RECT 9.004 14.972 11.476 15.004 ;
  LAYER M3 ;
        RECT 9.024 12.648 9.056 15.156 ;
  LAYER M3 ;
        RECT 9.088 12.648 9.12 15.156 ;
  LAYER M3 ;
        RECT 9.152 12.648 9.184 15.156 ;
  LAYER M3 ;
        RECT 9.216 12.648 9.248 15.156 ;
  LAYER M3 ;
        RECT 9.28 12.648 9.312 15.156 ;
  LAYER M3 ;
        RECT 9.344 12.648 9.376 15.156 ;
  LAYER M3 ;
        RECT 9.408 12.648 9.44 15.156 ;
  LAYER M3 ;
        RECT 9.472 12.648 9.504 15.156 ;
  LAYER M3 ;
        RECT 9.536 12.648 9.568 15.156 ;
  LAYER M3 ;
        RECT 9.6 12.648 9.632 15.156 ;
  LAYER M3 ;
        RECT 9.664 12.648 9.696 15.156 ;
  LAYER M3 ;
        RECT 9.728 12.648 9.76 15.156 ;
  LAYER M3 ;
        RECT 9.792 12.648 9.824 15.156 ;
  LAYER M3 ;
        RECT 9.856 12.648 9.888 15.156 ;
  LAYER M3 ;
        RECT 9.92 12.648 9.952 15.156 ;
  LAYER M3 ;
        RECT 9.984 12.648 10.016 15.156 ;
  LAYER M3 ;
        RECT 10.048 12.648 10.08 15.156 ;
  LAYER M3 ;
        RECT 10.112 12.648 10.144 15.156 ;
  LAYER M3 ;
        RECT 10.176 12.648 10.208 15.156 ;
  LAYER M3 ;
        RECT 10.24 12.648 10.272 15.156 ;
  LAYER M3 ;
        RECT 10.304 12.648 10.336 15.156 ;
  LAYER M3 ;
        RECT 10.368 12.648 10.4 15.156 ;
  LAYER M3 ;
        RECT 10.432 12.648 10.464 15.156 ;
  LAYER M3 ;
        RECT 10.496 12.648 10.528 15.156 ;
  LAYER M3 ;
        RECT 10.56 12.648 10.592 15.156 ;
  LAYER M3 ;
        RECT 10.624 12.648 10.656 15.156 ;
  LAYER M3 ;
        RECT 10.688 12.648 10.72 15.156 ;
  LAYER M3 ;
        RECT 10.752 12.648 10.784 15.156 ;
  LAYER M3 ;
        RECT 10.816 12.648 10.848 15.156 ;
  LAYER M3 ;
        RECT 10.88 12.648 10.912 15.156 ;
  LAYER M3 ;
        RECT 10.944 12.648 10.976 15.156 ;
  LAYER M3 ;
        RECT 11.008 12.648 11.04 15.156 ;
  LAYER M3 ;
        RECT 11.072 12.648 11.104 15.156 ;
  LAYER M3 ;
        RECT 11.136 12.648 11.168 15.156 ;
  LAYER M3 ;
        RECT 11.2 12.648 11.232 15.156 ;
  LAYER M3 ;
        RECT 11.264 12.648 11.296 15.156 ;
  LAYER M3 ;
        RECT 11.328 12.648 11.36 15.156 ;
  LAYER M3 ;
        RECT 11.424 12.648 11.456 15.156 ;
  LAYER M1 ;
        RECT 9.039 12.684 9.041 15.12 ;
  LAYER M1 ;
        RECT 9.119 12.684 9.121 15.12 ;
  LAYER M1 ;
        RECT 9.199 12.684 9.201 15.12 ;
  LAYER M1 ;
        RECT 9.279 12.684 9.281 15.12 ;
  LAYER M1 ;
        RECT 9.359 12.684 9.361 15.12 ;
  LAYER M1 ;
        RECT 9.439 12.684 9.441 15.12 ;
  LAYER M1 ;
        RECT 9.519 12.684 9.521 15.12 ;
  LAYER M1 ;
        RECT 9.599 12.684 9.601 15.12 ;
  LAYER M1 ;
        RECT 9.679 12.684 9.681 15.12 ;
  LAYER M1 ;
        RECT 9.759 12.684 9.761 15.12 ;
  LAYER M1 ;
        RECT 9.839 12.684 9.841 15.12 ;
  LAYER M1 ;
        RECT 9.919 12.684 9.921 15.12 ;
  LAYER M1 ;
        RECT 9.999 12.684 10.001 15.12 ;
  LAYER M1 ;
        RECT 10.079 12.684 10.081 15.12 ;
  LAYER M1 ;
        RECT 10.159 12.684 10.161 15.12 ;
  LAYER M1 ;
        RECT 10.239 12.684 10.241 15.12 ;
  LAYER M1 ;
        RECT 10.319 12.684 10.321 15.12 ;
  LAYER M1 ;
        RECT 10.399 12.684 10.401 15.12 ;
  LAYER M1 ;
        RECT 10.479 12.684 10.481 15.12 ;
  LAYER M1 ;
        RECT 10.559 12.684 10.561 15.12 ;
  LAYER M1 ;
        RECT 10.639 12.684 10.641 15.12 ;
  LAYER M1 ;
        RECT 10.719 12.684 10.721 15.12 ;
  LAYER M1 ;
        RECT 10.799 12.684 10.801 15.12 ;
  LAYER M1 ;
        RECT 10.879 12.684 10.881 15.12 ;
  LAYER M1 ;
        RECT 10.959 12.684 10.961 15.12 ;
  LAYER M1 ;
        RECT 11.039 12.684 11.041 15.12 ;
  LAYER M1 ;
        RECT 11.119 12.684 11.121 15.12 ;
  LAYER M1 ;
        RECT 11.199 12.684 11.201 15.12 ;
  LAYER M1 ;
        RECT 11.279 12.684 11.281 15.12 ;
  LAYER M1 ;
        RECT 11.359 12.684 11.361 15.12 ;
  LAYER M2 ;
        RECT 9.04 12.683 11.44 12.685 ;
  LAYER M2 ;
        RECT 9.04 12.767 11.44 12.769 ;
  LAYER M2 ;
        RECT 9.04 12.851 11.44 12.853 ;
  LAYER M2 ;
        RECT 9.04 12.935 11.44 12.937 ;
  LAYER M2 ;
        RECT 9.04 13.019 11.44 13.021 ;
  LAYER M2 ;
        RECT 9.04 13.103 11.44 13.105 ;
  LAYER M2 ;
        RECT 9.04 13.187 11.44 13.189 ;
  LAYER M2 ;
        RECT 9.04 13.271 11.44 13.273 ;
  LAYER M2 ;
        RECT 9.04 13.355 11.44 13.357 ;
  LAYER M2 ;
        RECT 9.04 13.439 11.44 13.441 ;
  LAYER M2 ;
        RECT 9.04 13.523 11.44 13.525 ;
  LAYER M2 ;
        RECT 9.04 13.607 11.44 13.609 ;
  LAYER M2 ;
        RECT 9.04 13.6905 11.44 13.6925 ;
  LAYER M2 ;
        RECT 9.04 13.775 11.44 13.777 ;
  LAYER M2 ;
        RECT 9.04 13.859 11.44 13.861 ;
  LAYER M2 ;
        RECT 9.04 13.943 11.44 13.945 ;
  LAYER M2 ;
        RECT 9.04 14.027 11.44 14.029 ;
  LAYER M2 ;
        RECT 9.04 14.111 11.44 14.113 ;
  LAYER M2 ;
        RECT 9.04 14.195 11.44 14.197 ;
  LAYER M2 ;
        RECT 9.04 14.279 11.44 14.281 ;
  LAYER M2 ;
        RECT 9.04 14.363 11.44 14.365 ;
  LAYER M2 ;
        RECT 9.04 14.447 11.44 14.449 ;
  LAYER M2 ;
        RECT 9.04 14.531 11.44 14.533 ;
  LAYER M2 ;
        RECT 9.04 14.615 11.44 14.617 ;
  LAYER M2 ;
        RECT 9.04 14.699 11.44 14.701 ;
  LAYER M2 ;
        RECT 9.04 14.783 11.44 14.785 ;
  LAYER M2 ;
        RECT 9.04 14.867 11.44 14.869 ;
  LAYER M2 ;
        RECT 9.04 14.951 11.44 14.953 ;
  LAYER M2 ;
        RECT 9.04 15.035 11.44 15.037 ;
  LAYER M1 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M1 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M1 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M1 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M1 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M1 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M1 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M1 ;
        RECT 9.472 15.588 9.504 18.096 ;
  LAYER M1 ;
        RECT 9.536 15.588 9.568 18.096 ;
  LAYER M1 ;
        RECT 9.6 15.588 9.632 18.096 ;
  LAYER M1 ;
        RECT 9.664 15.588 9.696 18.096 ;
  LAYER M1 ;
        RECT 9.728 15.588 9.76 18.096 ;
  LAYER M1 ;
        RECT 9.792 15.588 9.824 18.096 ;
  LAYER M1 ;
        RECT 9.856 15.588 9.888 18.096 ;
  LAYER M1 ;
        RECT 9.92 15.588 9.952 18.096 ;
  LAYER M1 ;
        RECT 9.984 15.588 10.016 18.096 ;
  LAYER M1 ;
        RECT 10.048 15.588 10.08 18.096 ;
  LAYER M1 ;
        RECT 10.112 15.588 10.144 18.096 ;
  LAYER M1 ;
        RECT 10.176 15.588 10.208 18.096 ;
  LAYER M1 ;
        RECT 10.24 15.588 10.272 18.096 ;
  LAYER M1 ;
        RECT 10.304 15.588 10.336 18.096 ;
  LAYER M1 ;
        RECT 10.368 15.588 10.4 18.096 ;
  LAYER M1 ;
        RECT 10.432 15.588 10.464 18.096 ;
  LAYER M1 ;
        RECT 10.496 15.588 10.528 18.096 ;
  LAYER M1 ;
        RECT 10.56 15.588 10.592 18.096 ;
  LAYER M1 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M1 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M1 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M1 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M1 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M1 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M1 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M1 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M1 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M1 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M1 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M1 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M2 ;
        RECT 9.004 15.672 11.476 15.704 ;
  LAYER M2 ;
        RECT 9.004 15.736 11.476 15.768 ;
  LAYER M2 ;
        RECT 9.004 15.8 11.476 15.832 ;
  LAYER M2 ;
        RECT 9.004 15.864 11.476 15.896 ;
  LAYER M2 ;
        RECT 9.004 15.928 11.476 15.96 ;
  LAYER M2 ;
        RECT 9.004 15.992 11.476 16.024 ;
  LAYER M2 ;
        RECT 9.004 16.056 11.476 16.088 ;
  LAYER M2 ;
        RECT 9.004 16.12 11.476 16.152 ;
  LAYER M2 ;
        RECT 9.004 16.184 11.476 16.216 ;
  LAYER M2 ;
        RECT 9.004 16.248 11.476 16.28 ;
  LAYER M2 ;
        RECT 9.004 16.312 11.476 16.344 ;
  LAYER M2 ;
        RECT 9.004 16.376 11.476 16.408 ;
  LAYER M2 ;
        RECT 9.004 16.44 11.476 16.472 ;
  LAYER M2 ;
        RECT 9.004 16.504 11.476 16.536 ;
  LAYER M2 ;
        RECT 9.004 16.568 11.476 16.6 ;
  LAYER M2 ;
        RECT 9.004 16.632 11.476 16.664 ;
  LAYER M2 ;
        RECT 9.004 16.696 11.476 16.728 ;
  LAYER M2 ;
        RECT 9.004 16.76 11.476 16.792 ;
  LAYER M2 ;
        RECT 9.004 16.824 11.476 16.856 ;
  LAYER M2 ;
        RECT 9.004 16.888 11.476 16.92 ;
  LAYER M2 ;
        RECT 9.004 16.952 11.476 16.984 ;
  LAYER M2 ;
        RECT 9.004 17.016 11.476 17.048 ;
  LAYER M2 ;
        RECT 9.004 17.08 11.476 17.112 ;
  LAYER M2 ;
        RECT 9.004 17.144 11.476 17.176 ;
  LAYER M2 ;
        RECT 9.004 17.208 11.476 17.24 ;
  LAYER M2 ;
        RECT 9.004 17.272 11.476 17.304 ;
  LAYER M2 ;
        RECT 9.004 17.336 11.476 17.368 ;
  LAYER M2 ;
        RECT 9.004 17.4 11.476 17.432 ;
  LAYER M2 ;
        RECT 9.004 17.464 11.476 17.496 ;
  LAYER M2 ;
        RECT 9.004 17.528 11.476 17.56 ;
  LAYER M2 ;
        RECT 9.004 17.592 11.476 17.624 ;
  LAYER M2 ;
        RECT 9.004 17.656 11.476 17.688 ;
  LAYER M2 ;
        RECT 9.004 17.72 11.476 17.752 ;
  LAYER M2 ;
        RECT 9.004 17.784 11.476 17.816 ;
  LAYER M2 ;
        RECT 9.004 17.848 11.476 17.88 ;
  LAYER M2 ;
        RECT 9.004 17.912 11.476 17.944 ;
  LAYER M3 ;
        RECT 9.024 15.588 9.056 18.096 ;
  LAYER M3 ;
        RECT 9.088 15.588 9.12 18.096 ;
  LAYER M3 ;
        RECT 9.152 15.588 9.184 18.096 ;
  LAYER M3 ;
        RECT 9.216 15.588 9.248 18.096 ;
  LAYER M3 ;
        RECT 9.28 15.588 9.312 18.096 ;
  LAYER M3 ;
        RECT 9.344 15.588 9.376 18.096 ;
  LAYER M3 ;
        RECT 9.408 15.588 9.44 18.096 ;
  LAYER M3 ;
        RECT 9.472 15.588 9.504 18.096 ;
  LAYER M3 ;
        RECT 9.536 15.588 9.568 18.096 ;
  LAYER M3 ;
        RECT 9.6 15.588 9.632 18.096 ;
  LAYER M3 ;
        RECT 9.664 15.588 9.696 18.096 ;
  LAYER M3 ;
        RECT 9.728 15.588 9.76 18.096 ;
  LAYER M3 ;
        RECT 9.792 15.588 9.824 18.096 ;
  LAYER M3 ;
        RECT 9.856 15.588 9.888 18.096 ;
  LAYER M3 ;
        RECT 9.92 15.588 9.952 18.096 ;
  LAYER M3 ;
        RECT 9.984 15.588 10.016 18.096 ;
  LAYER M3 ;
        RECT 10.048 15.588 10.08 18.096 ;
  LAYER M3 ;
        RECT 10.112 15.588 10.144 18.096 ;
  LAYER M3 ;
        RECT 10.176 15.588 10.208 18.096 ;
  LAYER M3 ;
        RECT 10.24 15.588 10.272 18.096 ;
  LAYER M3 ;
        RECT 10.304 15.588 10.336 18.096 ;
  LAYER M3 ;
        RECT 10.368 15.588 10.4 18.096 ;
  LAYER M3 ;
        RECT 10.432 15.588 10.464 18.096 ;
  LAYER M3 ;
        RECT 10.496 15.588 10.528 18.096 ;
  LAYER M3 ;
        RECT 10.56 15.588 10.592 18.096 ;
  LAYER M3 ;
        RECT 10.624 15.588 10.656 18.096 ;
  LAYER M3 ;
        RECT 10.688 15.588 10.72 18.096 ;
  LAYER M3 ;
        RECT 10.752 15.588 10.784 18.096 ;
  LAYER M3 ;
        RECT 10.816 15.588 10.848 18.096 ;
  LAYER M3 ;
        RECT 10.88 15.588 10.912 18.096 ;
  LAYER M3 ;
        RECT 10.944 15.588 10.976 18.096 ;
  LAYER M3 ;
        RECT 11.008 15.588 11.04 18.096 ;
  LAYER M3 ;
        RECT 11.072 15.588 11.104 18.096 ;
  LAYER M3 ;
        RECT 11.136 15.588 11.168 18.096 ;
  LAYER M3 ;
        RECT 11.2 15.588 11.232 18.096 ;
  LAYER M3 ;
        RECT 11.264 15.588 11.296 18.096 ;
  LAYER M3 ;
        RECT 11.328 15.588 11.36 18.096 ;
  LAYER M3 ;
        RECT 11.424 15.588 11.456 18.096 ;
  LAYER M1 ;
        RECT 9.039 15.624 9.041 18.06 ;
  LAYER M1 ;
        RECT 9.119 15.624 9.121 18.06 ;
  LAYER M1 ;
        RECT 9.199 15.624 9.201 18.06 ;
  LAYER M1 ;
        RECT 9.279 15.624 9.281 18.06 ;
  LAYER M1 ;
        RECT 9.359 15.624 9.361 18.06 ;
  LAYER M1 ;
        RECT 9.439 15.624 9.441 18.06 ;
  LAYER M1 ;
        RECT 9.519 15.624 9.521 18.06 ;
  LAYER M1 ;
        RECT 9.599 15.624 9.601 18.06 ;
  LAYER M1 ;
        RECT 9.679 15.624 9.681 18.06 ;
  LAYER M1 ;
        RECT 9.759 15.624 9.761 18.06 ;
  LAYER M1 ;
        RECT 9.839 15.624 9.841 18.06 ;
  LAYER M1 ;
        RECT 9.919 15.624 9.921 18.06 ;
  LAYER M1 ;
        RECT 9.999 15.624 10.001 18.06 ;
  LAYER M1 ;
        RECT 10.079 15.624 10.081 18.06 ;
  LAYER M1 ;
        RECT 10.159 15.624 10.161 18.06 ;
  LAYER M1 ;
        RECT 10.239 15.624 10.241 18.06 ;
  LAYER M1 ;
        RECT 10.319 15.624 10.321 18.06 ;
  LAYER M1 ;
        RECT 10.399 15.624 10.401 18.06 ;
  LAYER M1 ;
        RECT 10.479 15.624 10.481 18.06 ;
  LAYER M1 ;
        RECT 10.559 15.624 10.561 18.06 ;
  LAYER M1 ;
        RECT 10.639 15.624 10.641 18.06 ;
  LAYER M1 ;
        RECT 10.719 15.624 10.721 18.06 ;
  LAYER M1 ;
        RECT 10.799 15.624 10.801 18.06 ;
  LAYER M1 ;
        RECT 10.879 15.624 10.881 18.06 ;
  LAYER M1 ;
        RECT 10.959 15.624 10.961 18.06 ;
  LAYER M1 ;
        RECT 11.039 15.624 11.041 18.06 ;
  LAYER M1 ;
        RECT 11.119 15.624 11.121 18.06 ;
  LAYER M1 ;
        RECT 11.199 15.624 11.201 18.06 ;
  LAYER M1 ;
        RECT 11.279 15.624 11.281 18.06 ;
  LAYER M1 ;
        RECT 11.359 15.624 11.361 18.06 ;
  LAYER M2 ;
        RECT 9.04 15.623 11.44 15.625 ;
  LAYER M2 ;
        RECT 9.04 15.707 11.44 15.709 ;
  LAYER M2 ;
        RECT 9.04 15.791 11.44 15.793 ;
  LAYER M2 ;
        RECT 9.04 15.875 11.44 15.877 ;
  LAYER M2 ;
        RECT 9.04 15.959 11.44 15.961 ;
  LAYER M2 ;
        RECT 9.04 16.043 11.44 16.045 ;
  LAYER M2 ;
        RECT 9.04 16.127 11.44 16.129 ;
  LAYER M2 ;
        RECT 9.04 16.211 11.44 16.213 ;
  LAYER M2 ;
        RECT 9.04 16.295 11.44 16.297 ;
  LAYER M2 ;
        RECT 9.04 16.379 11.44 16.381 ;
  LAYER M2 ;
        RECT 9.04 16.463 11.44 16.465 ;
  LAYER M2 ;
        RECT 9.04 16.547 11.44 16.549 ;
  LAYER M2 ;
        RECT 9.04 16.6305 11.44 16.6325 ;
  LAYER M2 ;
        RECT 9.04 16.715 11.44 16.717 ;
  LAYER M2 ;
        RECT 9.04 16.799 11.44 16.801 ;
  LAYER M2 ;
        RECT 9.04 16.883 11.44 16.885 ;
  LAYER M2 ;
        RECT 9.04 16.967 11.44 16.969 ;
  LAYER M2 ;
        RECT 9.04 17.051 11.44 17.053 ;
  LAYER M2 ;
        RECT 9.04 17.135 11.44 17.137 ;
  LAYER M2 ;
        RECT 9.04 17.219 11.44 17.221 ;
  LAYER M2 ;
        RECT 9.04 17.303 11.44 17.305 ;
  LAYER M2 ;
        RECT 9.04 17.387 11.44 17.389 ;
  LAYER M2 ;
        RECT 9.04 17.471 11.44 17.473 ;
  LAYER M2 ;
        RECT 9.04 17.555 11.44 17.557 ;
  LAYER M2 ;
        RECT 9.04 17.639 11.44 17.641 ;
  LAYER M2 ;
        RECT 9.04 17.723 11.44 17.725 ;
  LAYER M2 ;
        RECT 9.04 17.807 11.44 17.809 ;
  LAYER M2 ;
        RECT 9.04 17.891 11.44 17.893 ;
  LAYER M2 ;
        RECT 9.04 17.975 11.44 17.977 ;
  LAYER M1 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M1 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M1 ;
        RECT 12.032 0.888 12.064 3.396 ;
  LAYER M1 ;
        RECT 12.096 0.888 12.128 3.396 ;
  LAYER M1 ;
        RECT 12.16 0.888 12.192 3.396 ;
  LAYER M1 ;
        RECT 12.224 0.888 12.256 3.396 ;
  LAYER M1 ;
        RECT 12.288 0.888 12.32 3.396 ;
  LAYER M1 ;
        RECT 12.352 0.888 12.384 3.396 ;
  LAYER M1 ;
        RECT 12.416 0.888 12.448 3.396 ;
  LAYER M1 ;
        RECT 12.48 0.888 12.512 3.396 ;
  LAYER M1 ;
        RECT 12.544 0.888 12.576 3.396 ;
  LAYER M1 ;
        RECT 12.608 0.888 12.64 3.396 ;
  LAYER M1 ;
        RECT 12.672 0.888 12.704 3.396 ;
  LAYER M1 ;
        RECT 12.736 0.888 12.768 3.396 ;
  LAYER M1 ;
        RECT 12.8 0.888 12.832 3.396 ;
  LAYER M1 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M1 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M1 ;
        RECT 12.992 0.888 13.024 3.396 ;
  LAYER M1 ;
        RECT 13.056 0.888 13.088 3.396 ;
  LAYER M1 ;
        RECT 13.12 0.888 13.152 3.396 ;
  LAYER M1 ;
        RECT 13.184 0.888 13.216 3.396 ;
  LAYER M1 ;
        RECT 13.248 0.888 13.28 3.396 ;
  LAYER M1 ;
        RECT 13.312 0.888 13.344 3.396 ;
  LAYER M1 ;
        RECT 13.376 0.888 13.408 3.396 ;
  LAYER M1 ;
        RECT 13.44 0.888 13.472 3.396 ;
  LAYER M1 ;
        RECT 13.504 0.888 13.536 3.396 ;
  LAYER M1 ;
        RECT 13.568 0.888 13.6 3.396 ;
  LAYER M1 ;
        RECT 13.632 0.888 13.664 3.396 ;
  LAYER M1 ;
        RECT 13.696 0.888 13.728 3.396 ;
  LAYER M1 ;
        RECT 13.76 0.888 13.792 3.396 ;
  LAYER M1 ;
        RECT 13.824 0.888 13.856 3.396 ;
  LAYER M1 ;
        RECT 13.888 0.888 13.92 3.396 ;
  LAYER M1 ;
        RECT 13.952 0.888 13.984 3.396 ;
  LAYER M1 ;
        RECT 14.016 0.888 14.048 3.396 ;
  LAYER M1 ;
        RECT 14.08 0.888 14.112 3.396 ;
  LAYER M1 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M1 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M2 ;
        RECT 11.884 0.972 14.356 1.004 ;
  LAYER M2 ;
        RECT 11.884 1.036 14.356 1.068 ;
  LAYER M2 ;
        RECT 11.884 1.1 14.356 1.132 ;
  LAYER M2 ;
        RECT 11.884 1.164 14.356 1.196 ;
  LAYER M2 ;
        RECT 11.884 1.228 14.356 1.26 ;
  LAYER M2 ;
        RECT 11.884 1.292 14.356 1.324 ;
  LAYER M2 ;
        RECT 11.884 1.356 14.356 1.388 ;
  LAYER M2 ;
        RECT 11.884 1.42 14.356 1.452 ;
  LAYER M2 ;
        RECT 11.884 1.484 14.356 1.516 ;
  LAYER M2 ;
        RECT 11.884 1.548 14.356 1.58 ;
  LAYER M2 ;
        RECT 11.884 1.612 14.356 1.644 ;
  LAYER M2 ;
        RECT 11.884 1.676 14.356 1.708 ;
  LAYER M2 ;
        RECT 11.884 1.74 14.356 1.772 ;
  LAYER M2 ;
        RECT 11.884 1.804 14.356 1.836 ;
  LAYER M2 ;
        RECT 11.884 1.868 14.356 1.9 ;
  LAYER M2 ;
        RECT 11.884 1.932 14.356 1.964 ;
  LAYER M2 ;
        RECT 11.884 1.996 14.356 2.028 ;
  LAYER M2 ;
        RECT 11.884 2.06 14.356 2.092 ;
  LAYER M2 ;
        RECT 11.884 2.124 14.356 2.156 ;
  LAYER M2 ;
        RECT 11.884 2.188 14.356 2.22 ;
  LAYER M2 ;
        RECT 11.884 2.252 14.356 2.284 ;
  LAYER M2 ;
        RECT 11.884 2.316 14.356 2.348 ;
  LAYER M2 ;
        RECT 11.884 2.38 14.356 2.412 ;
  LAYER M2 ;
        RECT 11.884 2.444 14.356 2.476 ;
  LAYER M2 ;
        RECT 11.884 2.508 14.356 2.54 ;
  LAYER M2 ;
        RECT 11.884 2.572 14.356 2.604 ;
  LAYER M2 ;
        RECT 11.884 2.636 14.356 2.668 ;
  LAYER M2 ;
        RECT 11.884 2.7 14.356 2.732 ;
  LAYER M2 ;
        RECT 11.884 2.764 14.356 2.796 ;
  LAYER M2 ;
        RECT 11.884 2.828 14.356 2.86 ;
  LAYER M2 ;
        RECT 11.884 2.892 14.356 2.924 ;
  LAYER M2 ;
        RECT 11.884 2.956 14.356 2.988 ;
  LAYER M2 ;
        RECT 11.884 3.02 14.356 3.052 ;
  LAYER M2 ;
        RECT 11.884 3.084 14.356 3.116 ;
  LAYER M2 ;
        RECT 11.884 3.148 14.356 3.18 ;
  LAYER M2 ;
        RECT 11.884 3.212 14.356 3.244 ;
  LAYER M3 ;
        RECT 11.904 0.888 11.936 3.396 ;
  LAYER M3 ;
        RECT 11.968 0.888 12 3.396 ;
  LAYER M3 ;
        RECT 12.032 0.888 12.064 3.396 ;
  LAYER M3 ;
        RECT 12.096 0.888 12.128 3.396 ;
  LAYER M3 ;
        RECT 12.16 0.888 12.192 3.396 ;
  LAYER M3 ;
        RECT 12.224 0.888 12.256 3.396 ;
  LAYER M3 ;
        RECT 12.288 0.888 12.32 3.396 ;
  LAYER M3 ;
        RECT 12.352 0.888 12.384 3.396 ;
  LAYER M3 ;
        RECT 12.416 0.888 12.448 3.396 ;
  LAYER M3 ;
        RECT 12.48 0.888 12.512 3.396 ;
  LAYER M3 ;
        RECT 12.544 0.888 12.576 3.396 ;
  LAYER M3 ;
        RECT 12.608 0.888 12.64 3.396 ;
  LAYER M3 ;
        RECT 12.672 0.888 12.704 3.396 ;
  LAYER M3 ;
        RECT 12.736 0.888 12.768 3.396 ;
  LAYER M3 ;
        RECT 12.8 0.888 12.832 3.396 ;
  LAYER M3 ;
        RECT 12.864 0.888 12.896 3.396 ;
  LAYER M3 ;
        RECT 12.928 0.888 12.96 3.396 ;
  LAYER M3 ;
        RECT 12.992 0.888 13.024 3.396 ;
  LAYER M3 ;
        RECT 13.056 0.888 13.088 3.396 ;
  LAYER M3 ;
        RECT 13.12 0.888 13.152 3.396 ;
  LAYER M3 ;
        RECT 13.184 0.888 13.216 3.396 ;
  LAYER M3 ;
        RECT 13.248 0.888 13.28 3.396 ;
  LAYER M3 ;
        RECT 13.312 0.888 13.344 3.396 ;
  LAYER M3 ;
        RECT 13.376 0.888 13.408 3.396 ;
  LAYER M3 ;
        RECT 13.44 0.888 13.472 3.396 ;
  LAYER M3 ;
        RECT 13.504 0.888 13.536 3.396 ;
  LAYER M3 ;
        RECT 13.568 0.888 13.6 3.396 ;
  LAYER M3 ;
        RECT 13.632 0.888 13.664 3.396 ;
  LAYER M3 ;
        RECT 13.696 0.888 13.728 3.396 ;
  LAYER M3 ;
        RECT 13.76 0.888 13.792 3.396 ;
  LAYER M3 ;
        RECT 13.824 0.888 13.856 3.396 ;
  LAYER M3 ;
        RECT 13.888 0.888 13.92 3.396 ;
  LAYER M3 ;
        RECT 13.952 0.888 13.984 3.396 ;
  LAYER M3 ;
        RECT 14.016 0.888 14.048 3.396 ;
  LAYER M3 ;
        RECT 14.08 0.888 14.112 3.396 ;
  LAYER M3 ;
        RECT 14.144 0.888 14.176 3.396 ;
  LAYER M3 ;
        RECT 14.208 0.888 14.24 3.396 ;
  LAYER M3 ;
        RECT 14.304 0.888 14.336 3.396 ;
  LAYER M1 ;
        RECT 11.919 0.924 11.921 3.36 ;
  LAYER M1 ;
        RECT 11.999 0.924 12.001 3.36 ;
  LAYER M1 ;
        RECT 12.079 0.924 12.081 3.36 ;
  LAYER M1 ;
        RECT 12.159 0.924 12.161 3.36 ;
  LAYER M1 ;
        RECT 12.239 0.924 12.241 3.36 ;
  LAYER M1 ;
        RECT 12.319 0.924 12.321 3.36 ;
  LAYER M1 ;
        RECT 12.399 0.924 12.401 3.36 ;
  LAYER M1 ;
        RECT 12.479 0.924 12.481 3.36 ;
  LAYER M1 ;
        RECT 12.559 0.924 12.561 3.36 ;
  LAYER M1 ;
        RECT 12.639 0.924 12.641 3.36 ;
  LAYER M1 ;
        RECT 12.719 0.924 12.721 3.36 ;
  LAYER M1 ;
        RECT 12.799 0.924 12.801 3.36 ;
  LAYER M1 ;
        RECT 12.879 0.924 12.881 3.36 ;
  LAYER M1 ;
        RECT 12.959 0.924 12.961 3.36 ;
  LAYER M1 ;
        RECT 13.039 0.924 13.041 3.36 ;
  LAYER M1 ;
        RECT 13.119 0.924 13.121 3.36 ;
  LAYER M1 ;
        RECT 13.199 0.924 13.201 3.36 ;
  LAYER M1 ;
        RECT 13.279 0.924 13.281 3.36 ;
  LAYER M1 ;
        RECT 13.359 0.924 13.361 3.36 ;
  LAYER M1 ;
        RECT 13.439 0.924 13.441 3.36 ;
  LAYER M1 ;
        RECT 13.519 0.924 13.521 3.36 ;
  LAYER M1 ;
        RECT 13.599 0.924 13.601 3.36 ;
  LAYER M1 ;
        RECT 13.679 0.924 13.681 3.36 ;
  LAYER M1 ;
        RECT 13.759 0.924 13.761 3.36 ;
  LAYER M1 ;
        RECT 13.839 0.924 13.841 3.36 ;
  LAYER M1 ;
        RECT 13.919 0.924 13.921 3.36 ;
  LAYER M1 ;
        RECT 13.999 0.924 14.001 3.36 ;
  LAYER M1 ;
        RECT 14.079 0.924 14.081 3.36 ;
  LAYER M1 ;
        RECT 14.159 0.924 14.161 3.36 ;
  LAYER M1 ;
        RECT 14.239 0.924 14.241 3.36 ;
  LAYER M2 ;
        RECT 11.92 0.923 14.32 0.925 ;
  LAYER M2 ;
        RECT 11.92 1.007 14.32 1.009 ;
  LAYER M2 ;
        RECT 11.92 1.091 14.32 1.093 ;
  LAYER M2 ;
        RECT 11.92 1.175 14.32 1.177 ;
  LAYER M2 ;
        RECT 11.92 1.259 14.32 1.261 ;
  LAYER M2 ;
        RECT 11.92 1.343 14.32 1.345 ;
  LAYER M2 ;
        RECT 11.92 1.427 14.32 1.429 ;
  LAYER M2 ;
        RECT 11.92 1.511 14.32 1.513 ;
  LAYER M2 ;
        RECT 11.92 1.595 14.32 1.597 ;
  LAYER M2 ;
        RECT 11.92 1.679 14.32 1.681 ;
  LAYER M2 ;
        RECT 11.92 1.763 14.32 1.765 ;
  LAYER M2 ;
        RECT 11.92 1.847 14.32 1.849 ;
  LAYER M2 ;
        RECT 11.92 1.9305 14.32 1.9325 ;
  LAYER M2 ;
        RECT 11.92 2.015 14.32 2.017 ;
  LAYER M2 ;
        RECT 11.92 2.099 14.32 2.101 ;
  LAYER M2 ;
        RECT 11.92 2.183 14.32 2.185 ;
  LAYER M2 ;
        RECT 11.92 2.267 14.32 2.269 ;
  LAYER M2 ;
        RECT 11.92 2.351 14.32 2.353 ;
  LAYER M2 ;
        RECT 11.92 2.435 14.32 2.437 ;
  LAYER M2 ;
        RECT 11.92 2.519 14.32 2.521 ;
  LAYER M2 ;
        RECT 11.92 2.603 14.32 2.605 ;
  LAYER M2 ;
        RECT 11.92 2.687 14.32 2.689 ;
  LAYER M2 ;
        RECT 11.92 2.771 14.32 2.773 ;
  LAYER M2 ;
        RECT 11.92 2.855 14.32 2.857 ;
  LAYER M2 ;
        RECT 11.92 2.939 14.32 2.941 ;
  LAYER M2 ;
        RECT 11.92 3.023 14.32 3.025 ;
  LAYER M2 ;
        RECT 11.92 3.107 14.32 3.109 ;
  LAYER M2 ;
        RECT 11.92 3.191 14.32 3.193 ;
  LAYER M2 ;
        RECT 11.92 3.275 14.32 3.277 ;
  LAYER M1 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M1 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M1 ;
        RECT 12.032 3.828 12.064 6.336 ;
  LAYER M1 ;
        RECT 12.096 3.828 12.128 6.336 ;
  LAYER M1 ;
        RECT 12.16 3.828 12.192 6.336 ;
  LAYER M1 ;
        RECT 12.224 3.828 12.256 6.336 ;
  LAYER M1 ;
        RECT 12.288 3.828 12.32 6.336 ;
  LAYER M1 ;
        RECT 12.352 3.828 12.384 6.336 ;
  LAYER M1 ;
        RECT 12.416 3.828 12.448 6.336 ;
  LAYER M1 ;
        RECT 12.48 3.828 12.512 6.336 ;
  LAYER M1 ;
        RECT 12.544 3.828 12.576 6.336 ;
  LAYER M1 ;
        RECT 12.608 3.828 12.64 6.336 ;
  LAYER M1 ;
        RECT 12.672 3.828 12.704 6.336 ;
  LAYER M1 ;
        RECT 12.736 3.828 12.768 6.336 ;
  LAYER M1 ;
        RECT 12.8 3.828 12.832 6.336 ;
  LAYER M1 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M1 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M1 ;
        RECT 12.992 3.828 13.024 6.336 ;
  LAYER M1 ;
        RECT 13.056 3.828 13.088 6.336 ;
  LAYER M1 ;
        RECT 13.12 3.828 13.152 6.336 ;
  LAYER M1 ;
        RECT 13.184 3.828 13.216 6.336 ;
  LAYER M1 ;
        RECT 13.248 3.828 13.28 6.336 ;
  LAYER M1 ;
        RECT 13.312 3.828 13.344 6.336 ;
  LAYER M1 ;
        RECT 13.376 3.828 13.408 6.336 ;
  LAYER M1 ;
        RECT 13.44 3.828 13.472 6.336 ;
  LAYER M1 ;
        RECT 13.504 3.828 13.536 6.336 ;
  LAYER M1 ;
        RECT 13.568 3.828 13.6 6.336 ;
  LAYER M1 ;
        RECT 13.632 3.828 13.664 6.336 ;
  LAYER M1 ;
        RECT 13.696 3.828 13.728 6.336 ;
  LAYER M1 ;
        RECT 13.76 3.828 13.792 6.336 ;
  LAYER M1 ;
        RECT 13.824 3.828 13.856 6.336 ;
  LAYER M1 ;
        RECT 13.888 3.828 13.92 6.336 ;
  LAYER M1 ;
        RECT 13.952 3.828 13.984 6.336 ;
  LAYER M1 ;
        RECT 14.016 3.828 14.048 6.336 ;
  LAYER M1 ;
        RECT 14.08 3.828 14.112 6.336 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M1 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M2 ;
        RECT 11.884 3.912 14.356 3.944 ;
  LAYER M2 ;
        RECT 11.884 3.976 14.356 4.008 ;
  LAYER M2 ;
        RECT 11.884 4.04 14.356 4.072 ;
  LAYER M2 ;
        RECT 11.884 4.104 14.356 4.136 ;
  LAYER M2 ;
        RECT 11.884 4.168 14.356 4.2 ;
  LAYER M2 ;
        RECT 11.884 4.232 14.356 4.264 ;
  LAYER M2 ;
        RECT 11.884 4.296 14.356 4.328 ;
  LAYER M2 ;
        RECT 11.884 4.36 14.356 4.392 ;
  LAYER M2 ;
        RECT 11.884 4.424 14.356 4.456 ;
  LAYER M2 ;
        RECT 11.884 4.488 14.356 4.52 ;
  LAYER M2 ;
        RECT 11.884 4.552 14.356 4.584 ;
  LAYER M2 ;
        RECT 11.884 4.616 14.356 4.648 ;
  LAYER M2 ;
        RECT 11.884 4.68 14.356 4.712 ;
  LAYER M2 ;
        RECT 11.884 4.744 14.356 4.776 ;
  LAYER M2 ;
        RECT 11.884 4.808 14.356 4.84 ;
  LAYER M2 ;
        RECT 11.884 4.872 14.356 4.904 ;
  LAYER M2 ;
        RECT 11.884 4.936 14.356 4.968 ;
  LAYER M2 ;
        RECT 11.884 5 14.356 5.032 ;
  LAYER M2 ;
        RECT 11.884 5.064 14.356 5.096 ;
  LAYER M2 ;
        RECT 11.884 5.128 14.356 5.16 ;
  LAYER M2 ;
        RECT 11.884 5.192 14.356 5.224 ;
  LAYER M2 ;
        RECT 11.884 5.256 14.356 5.288 ;
  LAYER M2 ;
        RECT 11.884 5.32 14.356 5.352 ;
  LAYER M2 ;
        RECT 11.884 5.384 14.356 5.416 ;
  LAYER M2 ;
        RECT 11.884 5.448 14.356 5.48 ;
  LAYER M2 ;
        RECT 11.884 5.512 14.356 5.544 ;
  LAYER M2 ;
        RECT 11.884 5.576 14.356 5.608 ;
  LAYER M2 ;
        RECT 11.884 5.64 14.356 5.672 ;
  LAYER M2 ;
        RECT 11.884 5.704 14.356 5.736 ;
  LAYER M2 ;
        RECT 11.884 5.768 14.356 5.8 ;
  LAYER M2 ;
        RECT 11.884 5.832 14.356 5.864 ;
  LAYER M2 ;
        RECT 11.884 5.896 14.356 5.928 ;
  LAYER M2 ;
        RECT 11.884 5.96 14.356 5.992 ;
  LAYER M2 ;
        RECT 11.884 6.024 14.356 6.056 ;
  LAYER M2 ;
        RECT 11.884 6.088 14.356 6.12 ;
  LAYER M2 ;
        RECT 11.884 6.152 14.356 6.184 ;
  LAYER M3 ;
        RECT 11.904 3.828 11.936 6.336 ;
  LAYER M3 ;
        RECT 11.968 3.828 12 6.336 ;
  LAYER M3 ;
        RECT 12.032 3.828 12.064 6.336 ;
  LAYER M3 ;
        RECT 12.096 3.828 12.128 6.336 ;
  LAYER M3 ;
        RECT 12.16 3.828 12.192 6.336 ;
  LAYER M3 ;
        RECT 12.224 3.828 12.256 6.336 ;
  LAYER M3 ;
        RECT 12.288 3.828 12.32 6.336 ;
  LAYER M3 ;
        RECT 12.352 3.828 12.384 6.336 ;
  LAYER M3 ;
        RECT 12.416 3.828 12.448 6.336 ;
  LAYER M3 ;
        RECT 12.48 3.828 12.512 6.336 ;
  LAYER M3 ;
        RECT 12.544 3.828 12.576 6.336 ;
  LAYER M3 ;
        RECT 12.608 3.828 12.64 6.336 ;
  LAYER M3 ;
        RECT 12.672 3.828 12.704 6.336 ;
  LAYER M3 ;
        RECT 12.736 3.828 12.768 6.336 ;
  LAYER M3 ;
        RECT 12.8 3.828 12.832 6.336 ;
  LAYER M3 ;
        RECT 12.864 3.828 12.896 6.336 ;
  LAYER M3 ;
        RECT 12.928 3.828 12.96 6.336 ;
  LAYER M3 ;
        RECT 12.992 3.828 13.024 6.336 ;
  LAYER M3 ;
        RECT 13.056 3.828 13.088 6.336 ;
  LAYER M3 ;
        RECT 13.12 3.828 13.152 6.336 ;
  LAYER M3 ;
        RECT 13.184 3.828 13.216 6.336 ;
  LAYER M3 ;
        RECT 13.248 3.828 13.28 6.336 ;
  LAYER M3 ;
        RECT 13.312 3.828 13.344 6.336 ;
  LAYER M3 ;
        RECT 13.376 3.828 13.408 6.336 ;
  LAYER M3 ;
        RECT 13.44 3.828 13.472 6.336 ;
  LAYER M3 ;
        RECT 13.504 3.828 13.536 6.336 ;
  LAYER M3 ;
        RECT 13.568 3.828 13.6 6.336 ;
  LAYER M3 ;
        RECT 13.632 3.828 13.664 6.336 ;
  LAYER M3 ;
        RECT 13.696 3.828 13.728 6.336 ;
  LAYER M3 ;
        RECT 13.76 3.828 13.792 6.336 ;
  LAYER M3 ;
        RECT 13.824 3.828 13.856 6.336 ;
  LAYER M3 ;
        RECT 13.888 3.828 13.92 6.336 ;
  LAYER M3 ;
        RECT 13.952 3.828 13.984 6.336 ;
  LAYER M3 ;
        RECT 14.016 3.828 14.048 6.336 ;
  LAYER M3 ;
        RECT 14.08 3.828 14.112 6.336 ;
  LAYER M3 ;
        RECT 14.144 3.828 14.176 6.336 ;
  LAYER M3 ;
        RECT 14.208 3.828 14.24 6.336 ;
  LAYER M3 ;
        RECT 14.304 3.828 14.336 6.336 ;
  LAYER M1 ;
        RECT 11.919 3.864 11.921 6.3 ;
  LAYER M1 ;
        RECT 11.999 3.864 12.001 6.3 ;
  LAYER M1 ;
        RECT 12.079 3.864 12.081 6.3 ;
  LAYER M1 ;
        RECT 12.159 3.864 12.161 6.3 ;
  LAYER M1 ;
        RECT 12.239 3.864 12.241 6.3 ;
  LAYER M1 ;
        RECT 12.319 3.864 12.321 6.3 ;
  LAYER M1 ;
        RECT 12.399 3.864 12.401 6.3 ;
  LAYER M1 ;
        RECT 12.479 3.864 12.481 6.3 ;
  LAYER M1 ;
        RECT 12.559 3.864 12.561 6.3 ;
  LAYER M1 ;
        RECT 12.639 3.864 12.641 6.3 ;
  LAYER M1 ;
        RECT 12.719 3.864 12.721 6.3 ;
  LAYER M1 ;
        RECT 12.799 3.864 12.801 6.3 ;
  LAYER M1 ;
        RECT 12.879 3.864 12.881 6.3 ;
  LAYER M1 ;
        RECT 12.959 3.864 12.961 6.3 ;
  LAYER M1 ;
        RECT 13.039 3.864 13.041 6.3 ;
  LAYER M1 ;
        RECT 13.119 3.864 13.121 6.3 ;
  LAYER M1 ;
        RECT 13.199 3.864 13.201 6.3 ;
  LAYER M1 ;
        RECT 13.279 3.864 13.281 6.3 ;
  LAYER M1 ;
        RECT 13.359 3.864 13.361 6.3 ;
  LAYER M1 ;
        RECT 13.439 3.864 13.441 6.3 ;
  LAYER M1 ;
        RECT 13.519 3.864 13.521 6.3 ;
  LAYER M1 ;
        RECT 13.599 3.864 13.601 6.3 ;
  LAYER M1 ;
        RECT 13.679 3.864 13.681 6.3 ;
  LAYER M1 ;
        RECT 13.759 3.864 13.761 6.3 ;
  LAYER M1 ;
        RECT 13.839 3.864 13.841 6.3 ;
  LAYER M1 ;
        RECT 13.919 3.864 13.921 6.3 ;
  LAYER M1 ;
        RECT 13.999 3.864 14.001 6.3 ;
  LAYER M1 ;
        RECT 14.079 3.864 14.081 6.3 ;
  LAYER M1 ;
        RECT 14.159 3.864 14.161 6.3 ;
  LAYER M1 ;
        RECT 14.239 3.864 14.241 6.3 ;
  LAYER M2 ;
        RECT 11.92 3.863 14.32 3.865 ;
  LAYER M2 ;
        RECT 11.92 3.947 14.32 3.949 ;
  LAYER M2 ;
        RECT 11.92 4.031 14.32 4.033 ;
  LAYER M2 ;
        RECT 11.92 4.115 14.32 4.117 ;
  LAYER M2 ;
        RECT 11.92 4.199 14.32 4.201 ;
  LAYER M2 ;
        RECT 11.92 4.283 14.32 4.285 ;
  LAYER M2 ;
        RECT 11.92 4.367 14.32 4.369 ;
  LAYER M2 ;
        RECT 11.92 4.451 14.32 4.453 ;
  LAYER M2 ;
        RECT 11.92 4.535 14.32 4.537 ;
  LAYER M2 ;
        RECT 11.92 4.619 14.32 4.621 ;
  LAYER M2 ;
        RECT 11.92 4.703 14.32 4.705 ;
  LAYER M2 ;
        RECT 11.92 4.787 14.32 4.789 ;
  LAYER M2 ;
        RECT 11.92 4.8705 14.32 4.8725 ;
  LAYER M2 ;
        RECT 11.92 4.955 14.32 4.957 ;
  LAYER M2 ;
        RECT 11.92 5.039 14.32 5.041 ;
  LAYER M2 ;
        RECT 11.92 5.123 14.32 5.125 ;
  LAYER M2 ;
        RECT 11.92 5.207 14.32 5.209 ;
  LAYER M2 ;
        RECT 11.92 5.291 14.32 5.293 ;
  LAYER M2 ;
        RECT 11.92 5.375 14.32 5.377 ;
  LAYER M2 ;
        RECT 11.92 5.459 14.32 5.461 ;
  LAYER M2 ;
        RECT 11.92 5.543 14.32 5.545 ;
  LAYER M2 ;
        RECT 11.92 5.627 14.32 5.629 ;
  LAYER M2 ;
        RECT 11.92 5.711 14.32 5.713 ;
  LAYER M2 ;
        RECT 11.92 5.795 14.32 5.797 ;
  LAYER M2 ;
        RECT 11.92 5.879 14.32 5.881 ;
  LAYER M2 ;
        RECT 11.92 5.963 14.32 5.965 ;
  LAYER M2 ;
        RECT 11.92 6.047 14.32 6.049 ;
  LAYER M2 ;
        RECT 11.92 6.131 14.32 6.133 ;
  LAYER M2 ;
        RECT 11.92 6.215 14.32 6.217 ;
  LAYER M1 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M1 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M1 ;
        RECT 12.032 6.768 12.064 9.276 ;
  LAYER M1 ;
        RECT 12.096 6.768 12.128 9.276 ;
  LAYER M1 ;
        RECT 12.16 6.768 12.192 9.276 ;
  LAYER M1 ;
        RECT 12.224 6.768 12.256 9.276 ;
  LAYER M1 ;
        RECT 12.288 6.768 12.32 9.276 ;
  LAYER M1 ;
        RECT 12.352 6.768 12.384 9.276 ;
  LAYER M1 ;
        RECT 12.416 6.768 12.448 9.276 ;
  LAYER M1 ;
        RECT 12.48 6.768 12.512 9.276 ;
  LAYER M1 ;
        RECT 12.544 6.768 12.576 9.276 ;
  LAYER M1 ;
        RECT 12.608 6.768 12.64 9.276 ;
  LAYER M1 ;
        RECT 12.672 6.768 12.704 9.276 ;
  LAYER M1 ;
        RECT 12.736 6.768 12.768 9.276 ;
  LAYER M1 ;
        RECT 12.8 6.768 12.832 9.276 ;
  LAYER M1 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M1 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M1 ;
        RECT 12.992 6.768 13.024 9.276 ;
  LAYER M1 ;
        RECT 13.056 6.768 13.088 9.276 ;
  LAYER M1 ;
        RECT 13.12 6.768 13.152 9.276 ;
  LAYER M1 ;
        RECT 13.184 6.768 13.216 9.276 ;
  LAYER M1 ;
        RECT 13.248 6.768 13.28 9.276 ;
  LAYER M1 ;
        RECT 13.312 6.768 13.344 9.276 ;
  LAYER M1 ;
        RECT 13.376 6.768 13.408 9.276 ;
  LAYER M1 ;
        RECT 13.44 6.768 13.472 9.276 ;
  LAYER M1 ;
        RECT 13.504 6.768 13.536 9.276 ;
  LAYER M1 ;
        RECT 13.568 6.768 13.6 9.276 ;
  LAYER M1 ;
        RECT 13.632 6.768 13.664 9.276 ;
  LAYER M1 ;
        RECT 13.696 6.768 13.728 9.276 ;
  LAYER M1 ;
        RECT 13.76 6.768 13.792 9.276 ;
  LAYER M1 ;
        RECT 13.824 6.768 13.856 9.276 ;
  LAYER M1 ;
        RECT 13.888 6.768 13.92 9.276 ;
  LAYER M1 ;
        RECT 13.952 6.768 13.984 9.276 ;
  LAYER M1 ;
        RECT 14.016 6.768 14.048 9.276 ;
  LAYER M1 ;
        RECT 14.08 6.768 14.112 9.276 ;
  LAYER M1 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M1 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M2 ;
        RECT 11.884 6.852 14.356 6.884 ;
  LAYER M2 ;
        RECT 11.884 6.916 14.356 6.948 ;
  LAYER M2 ;
        RECT 11.884 6.98 14.356 7.012 ;
  LAYER M2 ;
        RECT 11.884 7.044 14.356 7.076 ;
  LAYER M2 ;
        RECT 11.884 7.108 14.356 7.14 ;
  LAYER M2 ;
        RECT 11.884 7.172 14.356 7.204 ;
  LAYER M2 ;
        RECT 11.884 7.236 14.356 7.268 ;
  LAYER M2 ;
        RECT 11.884 7.3 14.356 7.332 ;
  LAYER M2 ;
        RECT 11.884 7.364 14.356 7.396 ;
  LAYER M2 ;
        RECT 11.884 7.428 14.356 7.46 ;
  LAYER M2 ;
        RECT 11.884 7.492 14.356 7.524 ;
  LAYER M2 ;
        RECT 11.884 7.556 14.356 7.588 ;
  LAYER M2 ;
        RECT 11.884 7.62 14.356 7.652 ;
  LAYER M2 ;
        RECT 11.884 7.684 14.356 7.716 ;
  LAYER M2 ;
        RECT 11.884 7.748 14.356 7.78 ;
  LAYER M2 ;
        RECT 11.884 7.812 14.356 7.844 ;
  LAYER M2 ;
        RECT 11.884 7.876 14.356 7.908 ;
  LAYER M2 ;
        RECT 11.884 7.94 14.356 7.972 ;
  LAYER M2 ;
        RECT 11.884 8.004 14.356 8.036 ;
  LAYER M2 ;
        RECT 11.884 8.068 14.356 8.1 ;
  LAYER M2 ;
        RECT 11.884 8.132 14.356 8.164 ;
  LAYER M2 ;
        RECT 11.884 8.196 14.356 8.228 ;
  LAYER M2 ;
        RECT 11.884 8.26 14.356 8.292 ;
  LAYER M2 ;
        RECT 11.884 8.324 14.356 8.356 ;
  LAYER M2 ;
        RECT 11.884 8.388 14.356 8.42 ;
  LAYER M2 ;
        RECT 11.884 8.452 14.356 8.484 ;
  LAYER M2 ;
        RECT 11.884 8.516 14.356 8.548 ;
  LAYER M2 ;
        RECT 11.884 8.58 14.356 8.612 ;
  LAYER M2 ;
        RECT 11.884 8.644 14.356 8.676 ;
  LAYER M2 ;
        RECT 11.884 8.708 14.356 8.74 ;
  LAYER M2 ;
        RECT 11.884 8.772 14.356 8.804 ;
  LAYER M2 ;
        RECT 11.884 8.836 14.356 8.868 ;
  LAYER M2 ;
        RECT 11.884 8.9 14.356 8.932 ;
  LAYER M2 ;
        RECT 11.884 8.964 14.356 8.996 ;
  LAYER M2 ;
        RECT 11.884 9.028 14.356 9.06 ;
  LAYER M2 ;
        RECT 11.884 9.092 14.356 9.124 ;
  LAYER M3 ;
        RECT 11.904 6.768 11.936 9.276 ;
  LAYER M3 ;
        RECT 11.968 6.768 12 9.276 ;
  LAYER M3 ;
        RECT 12.032 6.768 12.064 9.276 ;
  LAYER M3 ;
        RECT 12.096 6.768 12.128 9.276 ;
  LAYER M3 ;
        RECT 12.16 6.768 12.192 9.276 ;
  LAYER M3 ;
        RECT 12.224 6.768 12.256 9.276 ;
  LAYER M3 ;
        RECT 12.288 6.768 12.32 9.276 ;
  LAYER M3 ;
        RECT 12.352 6.768 12.384 9.276 ;
  LAYER M3 ;
        RECT 12.416 6.768 12.448 9.276 ;
  LAYER M3 ;
        RECT 12.48 6.768 12.512 9.276 ;
  LAYER M3 ;
        RECT 12.544 6.768 12.576 9.276 ;
  LAYER M3 ;
        RECT 12.608 6.768 12.64 9.276 ;
  LAYER M3 ;
        RECT 12.672 6.768 12.704 9.276 ;
  LAYER M3 ;
        RECT 12.736 6.768 12.768 9.276 ;
  LAYER M3 ;
        RECT 12.8 6.768 12.832 9.276 ;
  LAYER M3 ;
        RECT 12.864 6.768 12.896 9.276 ;
  LAYER M3 ;
        RECT 12.928 6.768 12.96 9.276 ;
  LAYER M3 ;
        RECT 12.992 6.768 13.024 9.276 ;
  LAYER M3 ;
        RECT 13.056 6.768 13.088 9.276 ;
  LAYER M3 ;
        RECT 13.12 6.768 13.152 9.276 ;
  LAYER M3 ;
        RECT 13.184 6.768 13.216 9.276 ;
  LAYER M3 ;
        RECT 13.248 6.768 13.28 9.276 ;
  LAYER M3 ;
        RECT 13.312 6.768 13.344 9.276 ;
  LAYER M3 ;
        RECT 13.376 6.768 13.408 9.276 ;
  LAYER M3 ;
        RECT 13.44 6.768 13.472 9.276 ;
  LAYER M3 ;
        RECT 13.504 6.768 13.536 9.276 ;
  LAYER M3 ;
        RECT 13.568 6.768 13.6 9.276 ;
  LAYER M3 ;
        RECT 13.632 6.768 13.664 9.276 ;
  LAYER M3 ;
        RECT 13.696 6.768 13.728 9.276 ;
  LAYER M3 ;
        RECT 13.76 6.768 13.792 9.276 ;
  LAYER M3 ;
        RECT 13.824 6.768 13.856 9.276 ;
  LAYER M3 ;
        RECT 13.888 6.768 13.92 9.276 ;
  LAYER M3 ;
        RECT 13.952 6.768 13.984 9.276 ;
  LAYER M3 ;
        RECT 14.016 6.768 14.048 9.276 ;
  LAYER M3 ;
        RECT 14.08 6.768 14.112 9.276 ;
  LAYER M3 ;
        RECT 14.144 6.768 14.176 9.276 ;
  LAYER M3 ;
        RECT 14.208 6.768 14.24 9.276 ;
  LAYER M3 ;
        RECT 14.304 6.768 14.336 9.276 ;
  LAYER M1 ;
        RECT 11.919 6.804 11.921 9.24 ;
  LAYER M1 ;
        RECT 11.999 6.804 12.001 9.24 ;
  LAYER M1 ;
        RECT 12.079 6.804 12.081 9.24 ;
  LAYER M1 ;
        RECT 12.159 6.804 12.161 9.24 ;
  LAYER M1 ;
        RECT 12.239 6.804 12.241 9.24 ;
  LAYER M1 ;
        RECT 12.319 6.804 12.321 9.24 ;
  LAYER M1 ;
        RECT 12.399 6.804 12.401 9.24 ;
  LAYER M1 ;
        RECT 12.479 6.804 12.481 9.24 ;
  LAYER M1 ;
        RECT 12.559 6.804 12.561 9.24 ;
  LAYER M1 ;
        RECT 12.639 6.804 12.641 9.24 ;
  LAYER M1 ;
        RECT 12.719 6.804 12.721 9.24 ;
  LAYER M1 ;
        RECT 12.799 6.804 12.801 9.24 ;
  LAYER M1 ;
        RECT 12.879 6.804 12.881 9.24 ;
  LAYER M1 ;
        RECT 12.959 6.804 12.961 9.24 ;
  LAYER M1 ;
        RECT 13.039 6.804 13.041 9.24 ;
  LAYER M1 ;
        RECT 13.119 6.804 13.121 9.24 ;
  LAYER M1 ;
        RECT 13.199 6.804 13.201 9.24 ;
  LAYER M1 ;
        RECT 13.279 6.804 13.281 9.24 ;
  LAYER M1 ;
        RECT 13.359 6.804 13.361 9.24 ;
  LAYER M1 ;
        RECT 13.439 6.804 13.441 9.24 ;
  LAYER M1 ;
        RECT 13.519 6.804 13.521 9.24 ;
  LAYER M1 ;
        RECT 13.599 6.804 13.601 9.24 ;
  LAYER M1 ;
        RECT 13.679 6.804 13.681 9.24 ;
  LAYER M1 ;
        RECT 13.759 6.804 13.761 9.24 ;
  LAYER M1 ;
        RECT 13.839 6.804 13.841 9.24 ;
  LAYER M1 ;
        RECT 13.919 6.804 13.921 9.24 ;
  LAYER M1 ;
        RECT 13.999 6.804 14.001 9.24 ;
  LAYER M1 ;
        RECT 14.079 6.804 14.081 9.24 ;
  LAYER M1 ;
        RECT 14.159 6.804 14.161 9.24 ;
  LAYER M1 ;
        RECT 14.239 6.804 14.241 9.24 ;
  LAYER M2 ;
        RECT 11.92 6.803 14.32 6.805 ;
  LAYER M2 ;
        RECT 11.92 6.887 14.32 6.889 ;
  LAYER M2 ;
        RECT 11.92 6.971 14.32 6.973 ;
  LAYER M2 ;
        RECT 11.92 7.055 14.32 7.057 ;
  LAYER M2 ;
        RECT 11.92 7.139 14.32 7.141 ;
  LAYER M2 ;
        RECT 11.92 7.223 14.32 7.225 ;
  LAYER M2 ;
        RECT 11.92 7.307 14.32 7.309 ;
  LAYER M2 ;
        RECT 11.92 7.391 14.32 7.393 ;
  LAYER M2 ;
        RECT 11.92 7.475 14.32 7.477 ;
  LAYER M2 ;
        RECT 11.92 7.559 14.32 7.561 ;
  LAYER M2 ;
        RECT 11.92 7.643 14.32 7.645 ;
  LAYER M2 ;
        RECT 11.92 7.727 14.32 7.729 ;
  LAYER M2 ;
        RECT 11.92 7.8105 14.32 7.8125 ;
  LAYER M2 ;
        RECT 11.92 7.895 14.32 7.897 ;
  LAYER M2 ;
        RECT 11.92 7.979 14.32 7.981 ;
  LAYER M2 ;
        RECT 11.92 8.063 14.32 8.065 ;
  LAYER M2 ;
        RECT 11.92 8.147 14.32 8.149 ;
  LAYER M2 ;
        RECT 11.92 8.231 14.32 8.233 ;
  LAYER M2 ;
        RECT 11.92 8.315 14.32 8.317 ;
  LAYER M2 ;
        RECT 11.92 8.399 14.32 8.401 ;
  LAYER M2 ;
        RECT 11.92 8.483 14.32 8.485 ;
  LAYER M2 ;
        RECT 11.92 8.567 14.32 8.569 ;
  LAYER M2 ;
        RECT 11.92 8.651 14.32 8.653 ;
  LAYER M2 ;
        RECT 11.92 8.735 14.32 8.737 ;
  LAYER M2 ;
        RECT 11.92 8.819 14.32 8.821 ;
  LAYER M2 ;
        RECT 11.92 8.903 14.32 8.905 ;
  LAYER M2 ;
        RECT 11.92 8.987 14.32 8.989 ;
  LAYER M2 ;
        RECT 11.92 9.071 14.32 9.073 ;
  LAYER M2 ;
        RECT 11.92 9.155 14.32 9.157 ;
  LAYER M1 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M1 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M1 ;
        RECT 12.032 9.708 12.064 12.216 ;
  LAYER M1 ;
        RECT 12.096 9.708 12.128 12.216 ;
  LAYER M1 ;
        RECT 12.16 9.708 12.192 12.216 ;
  LAYER M1 ;
        RECT 12.224 9.708 12.256 12.216 ;
  LAYER M1 ;
        RECT 12.288 9.708 12.32 12.216 ;
  LAYER M1 ;
        RECT 12.352 9.708 12.384 12.216 ;
  LAYER M1 ;
        RECT 12.416 9.708 12.448 12.216 ;
  LAYER M1 ;
        RECT 12.48 9.708 12.512 12.216 ;
  LAYER M1 ;
        RECT 12.544 9.708 12.576 12.216 ;
  LAYER M1 ;
        RECT 12.608 9.708 12.64 12.216 ;
  LAYER M1 ;
        RECT 12.672 9.708 12.704 12.216 ;
  LAYER M1 ;
        RECT 12.736 9.708 12.768 12.216 ;
  LAYER M1 ;
        RECT 12.8 9.708 12.832 12.216 ;
  LAYER M1 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M1 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M1 ;
        RECT 12.992 9.708 13.024 12.216 ;
  LAYER M1 ;
        RECT 13.056 9.708 13.088 12.216 ;
  LAYER M1 ;
        RECT 13.12 9.708 13.152 12.216 ;
  LAYER M1 ;
        RECT 13.184 9.708 13.216 12.216 ;
  LAYER M1 ;
        RECT 13.248 9.708 13.28 12.216 ;
  LAYER M1 ;
        RECT 13.312 9.708 13.344 12.216 ;
  LAYER M1 ;
        RECT 13.376 9.708 13.408 12.216 ;
  LAYER M1 ;
        RECT 13.44 9.708 13.472 12.216 ;
  LAYER M1 ;
        RECT 13.504 9.708 13.536 12.216 ;
  LAYER M1 ;
        RECT 13.568 9.708 13.6 12.216 ;
  LAYER M1 ;
        RECT 13.632 9.708 13.664 12.216 ;
  LAYER M1 ;
        RECT 13.696 9.708 13.728 12.216 ;
  LAYER M1 ;
        RECT 13.76 9.708 13.792 12.216 ;
  LAYER M1 ;
        RECT 13.824 9.708 13.856 12.216 ;
  LAYER M1 ;
        RECT 13.888 9.708 13.92 12.216 ;
  LAYER M1 ;
        RECT 13.952 9.708 13.984 12.216 ;
  LAYER M1 ;
        RECT 14.016 9.708 14.048 12.216 ;
  LAYER M1 ;
        RECT 14.08 9.708 14.112 12.216 ;
  LAYER M1 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M1 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M2 ;
        RECT 11.884 9.792 14.356 9.824 ;
  LAYER M2 ;
        RECT 11.884 9.856 14.356 9.888 ;
  LAYER M2 ;
        RECT 11.884 9.92 14.356 9.952 ;
  LAYER M2 ;
        RECT 11.884 9.984 14.356 10.016 ;
  LAYER M2 ;
        RECT 11.884 10.048 14.356 10.08 ;
  LAYER M2 ;
        RECT 11.884 10.112 14.356 10.144 ;
  LAYER M2 ;
        RECT 11.884 10.176 14.356 10.208 ;
  LAYER M2 ;
        RECT 11.884 10.24 14.356 10.272 ;
  LAYER M2 ;
        RECT 11.884 10.304 14.356 10.336 ;
  LAYER M2 ;
        RECT 11.884 10.368 14.356 10.4 ;
  LAYER M2 ;
        RECT 11.884 10.432 14.356 10.464 ;
  LAYER M2 ;
        RECT 11.884 10.496 14.356 10.528 ;
  LAYER M2 ;
        RECT 11.884 10.56 14.356 10.592 ;
  LAYER M2 ;
        RECT 11.884 10.624 14.356 10.656 ;
  LAYER M2 ;
        RECT 11.884 10.688 14.356 10.72 ;
  LAYER M2 ;
        RECT 11.884 10.752 14.356 10.784 ;
  LAYER M2 ;
        RECT 11.884 10.816 14.356 10.848 ;
  LAYER M2 ;
        RECT 11.884 10.88 14.356 10.912 ;
  LAYER M2 ;
        RECT 11.884 10.944 14.356 10.976 ;
  LAYER M2 ;
        RECT 11.884 11.008 14.356 11.04 ;
  LAYER M2 ;
        RECT 11.884 11.072 14.356 11.104 ;
  LAYER M2 ;
        RECT 11.884 11.136 14.356 11.168 ;
  LAYER M2 ;
        RECT 11.884 11.2 14.356 11.232 ;
  LAYER M2 ;
        RECT 11.884 11.264 14.356 11.296 ;
  LAYER M2 ;
        RECT 11.884 11.328 14.356 11.36 ;
  LAYER M2 ;
        RECT 11.884 11.392 14.356 11.424 ;
  LAYER M2 ;
        RECT 11.884 11.456 14.356 11.488 ;
  LAYER M2 ;
        RECT 11.884 11.52 14.356 11.552 ;
  LAYER M2 ;
        RECT 11.884 11.584 14.356 11.616 ;
  LAYER M2 ;
        RECT 11.884 11.648 14.356 11.68 ;
  LAYER M2 ;
        RECT 11.884 11.712 14.356 11.744 ;
  LAYER M2 ;
        RECT 11.884 11.776 14.356 11.808 ;
  LAYER M2 ;
        RECT 11.884 11.84 14.356 11.872 ;
  LAYER M2 ;
        RECT 11.884 11.904 14.356 11.936 ;
  LAYER M2 ;
        RECT 11.884 11.968 14.356 12 ;
  LAYER M2 ;
        RECT 11.884 12.032 14.356 12.064 ;
  LAYER M3 ;
        RECT 11.904 9.708 11.936 12.216 ;
  LAYER M3 ;
        RECT 11.968 9.708 12 12.216 ;
  LAYER M3 ;
        RECT 12.032 9.708 12.064 12.216 ;
  LAYER M3 ;
        RECT 12.096 9.708 12.128 12.216 ;
  LAYER M3 ;
        RECT 12.16 9.708 12.192 12.216 ;
  LAYER M3 ;
        RECT 12.224 9.708 12.256 12.216 ;
  LAYER M3 ;
        RECT 12.288 9.708 12.32 12.216 ;
  LAYER M3 ;
        RECT 12.352 9.708 12.384 12.216 ;
  LAYER M3 ;
        RECT 12.416 9.708 12.448 12.216 ;
  LAYER M3 ;
        RECT 12.48 9.708 12.512 12.216 ;
  LAYER M3 ;
        RECT 12.544 9.708 12.576 12.216 ;
  LAYER M3 ;
        RECT 12.608 9.708 12.64 12.216 ;
  LAYER M3 ;
        RECT 12.672 9.708 12.704 12.216 ;
  LAYER M3 ;
        RECT 12.736 9.708 12.768 12.216 ;
  LAYER M3 ;
        RECT 12.8 9.708 12.832 12.216 ;
  LAYER M3 ;
        RECT 12.864 9.708 12.896 12.216 ;
  LAYER M3 ;
        RECT 12.928 9.708 12.96 12.216 ;
  LAYER M3 ;
        RECT 12.992 9.708 13.024 12.216 ;
  LAYER M3 ;
        RECT 13.056 9.708 13.088 12.216 ;
  LAYER M3 ;
        RECT 13.12 9.708 13.152 12.216 ;
  LAYER M3 ;
        RECT 13.184 9.708 13.216 12.216 ;
  LAYER M3 ;
        RECT 13.248 9.708 13.28 12.216 ;
  LAYER M3 ;
        RECT 13.312 9.708 13.344 12.216 ;
  LAYER M3 ;
        RECT 13.376 9.708 13.408 12.216 ;
  LAYER M3 ;
        RECT 13.44 9.708 13.472 12.216 ;
  LAYER M3 ;
        RECT 13.504 9.708 13.536 12.216 ;
  LAYER M3 ;
        RECT 13.568 9.708 13.6 12.216 ;
  LAYER M3 ;
        RECT 13.632 9.708 13.664 12.216 ;
  LAYER M3 ;
        RECT 13.696 9.708 13.728 12.216 ;
  LAYER M3 ;
        RECT 13.76 9.708 13.792 12.216 ;
  LAYER M3 ;
        RECT 13.824 9.708 13.856 12.216 ;
  LAYER M3 ;
        RECT 13.888 9.708 13.92 12.216 ;
  LAYER M3 ;
        RECT 13.952 9.708 13.984 12.216 ;
  LAYER M3 ;
        RECT 14.016 9.708 14.048 12.216 ;
  LAYER M3 ;
        RECT 14.08 9.708 14.112 12.216 ;
  LAYER M3 ;
        RECT 14.144 9.708 14.176 12.216 ;
  LAYER M3 ;
        RECT 14.208 9.708 14.24 12.216 ;
  LAYER M3 ;
        RECT 14.304 9.708 14.336 12.216 ;
  LAYER M1 ;
        RECT 11.919 9.744 11.921 12.18 ;
  LAYER M1 ;
        RECT 11.999 9.744 12.001 12.18 ;
  LAYER M1 ;
        RECT 12.079 9.744 12.081 12.18 ;
  LAYER M1 ;
        RECT 12.159 9.744 12.161 12.18 ;
  LAYER M1 ;
        RECT 12.239 9.744 12.241 12.18 ;
  LAYER M1 ;
        RECT 12.319 9.744 12.321 12.18 ;
  LAYER M1 ;
        RECT 12.399 9.744 12.401 12.18 ;
  LAYER M1 ;
        RECT 12.479 9.744 12.481 12.18 ;
  LAYER M1 ;
        RECT 12.559 9.744 12.561 12.18 ;
  LAYER M1 ;
        RECT 12.639 9.744 12.641 12.18 ;
  LAYER M1 ;
        RECT 12.719 9.744 12.721 12.18 ;
  LAYER M1 ;
        RECT 12.799 9.744 12.801 12.18 ;
  LAYER M1 ;
        RECT 12.879 9.744 12.881 12.18 ;
  LAYER M1 ;
        RECT 12.959 9.744 12.961 12.18 ;
  LAYER M1 ;
        RECT 13.039 9.744 13.041 12.18 ;
  LAYER M1 ;
        RECT 13.119 9.744 13.121 12.18 ;
  LAYER M1 ;
        RECT 13.199 9.744 13.201 12.18 ;
  LAYER M1 ;
        RECT 13.279 9.744 13.281 12.18 ;
  LAYER M1 ;
        RECT 13.359 9.744 13.361 12.18 ;
  LAYER M1 ;
        RECT 13.439 9.744 13.441 12.18 ;
  LAYER M1 ;
        RECT 13.519 9.744 13.521 12.18 ;
  LAYER M1 ;
        RECT 13.599 9.744 13.601 12.18 ;
  LAYER M1 ;
        RECT 13.679 9.744 13.681 12.18 ;
  LAYER M1 ;
        RECT 13.759 9.744 13.761 12.18 ;
  LAYER M1 ;
        RECT 13.839 9.744 13.841 12.18 ;
  LAYER M1 ;
        RECT 13.919 9.744 13.921 12.18 ;
  LAYER M1 ;
        RECT 13.999 9.744 14.001 12.18 ;
  LAYER M1 ;
        RECT 14.079 9.744 14.081 12.18 ;
  LAYER M1 ;
        RECT 14.159 9.744 14.161 12.18 ;
  LAYER M1 ;
        RECT 14.239 9.744 14.241 12.18 ;
  LAYER M2 ;
        RECT 11.92 9.743 14.32 9.745 ;
  LAYER M2 ;
        RECT 11.92 9.827 14.32 9.829 ;
  LAYER M2 ;
        RECT 11.92 9.911 14.32 9.913 ;
  LAYER M2 ;
        RECT 11.92 9.995 14.32 9.997 ;
  LAYER M2 ;
        RECT 11.92 10.079 14.32 10.081 ;
  LAYER M2 ;
        RECT 11.92 10.163 14.32 10.165 ;
  LAYER M2 ;
        RECT 11.92 10.247 14.32 10.249 ;
  LAYER M2 ;
        RECT 11.92 10.331 14.32 10.333 ;
  LAYER M2 ;
        RECT 11.92 10.415 14.32 10.417 ;
  LAYER M2 ;
        RECT 11.92 10.499 14.32 10.501 ;
  LAYER M2 ;
        RECT 11.92 10.583 14.32 10.585 ;
  LAYER M2 ;
        RECT 11.92 10.667 14.32 10.669 ;
  LAYER M2 ;
        RECT 11.92 10.7505 14.32 10.7525 ;
  LAYER M2 ;
        RECT 11.92 10.835 14.32 10.837 ;
  LAYER M2 ;
        RECT 11.92 10.919 14.32 10.921 ;
  LAYER M2 ;
        RECT 11.92 11.003 14.32 11.005 ;
  LAYER M2 ;
        RECT 11.92 11.087 14.32 11.089 ;
  LAYER M2 ;
        RECT 11.92 11.171 14.32 11.173 ;
  LAYER M2 ;
        RECT 11.92 11.255 14.32 11.257 ;
  LAYER M2 ;
        RECT 11.92 11.339 14.32 11.341 ;
  LAYER M2 ;
        RECT 11.92 11.423 14.32 11.425 ;
  LAYER M2 ;
        RECT 11.92 11.507 14.32 11.509 ;
  LAYER M2 ;
        RECT 11.92 11.591 14.32 11.593 ;
  LAYER M2 ;
        RECT 11.92 11.675 14.32 11.677 ;
  LAYER M2 ;
        RECT 11.92 11.759 14.32 11.761 ;
  LAYER M2 ;
        RECT 11.92 11.843 14.32 11.845 ;
  LAYER M2 ;
        RECT 11.92 11.927 14.32 11.929 ;
  LAYER M2 ;
        RECT 11.92 12.011 14.32 12.013 ;
  LAYER M2 ;
        RECT 11.92 12.095 14.32 12.097 ;
  LAYER M1 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M1 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M1 ;
        RECT 12.032 12.648 12.064 15.156 ;
  LAYER M1 ;
        RECT 12.096 12.648 12.128 15.156 ;
  LAYER M1 ;
        RECT 12.16 12.648 12.192 15.156 ;
  LAYER M1 ;
        RECT 12.224 12.648 12.256 15.156 ;
  LAYER M1 ;
        RECT 12.288 12.648 12.32 15.156 ;
  LAYER M1 ;
        RECT 12.352 12.648 12.384 15.156 ;
  LAYER M1 ;
        RECT 12.416 12.648 12.448 15.156 ;
  LAYER M1 ;
        RECT 12.48 12.648 12.512 15.156 ;
  LAYER M1 ;
        RECT 12.544 12.648 12.576 15.156 ;
  LAYER M1 ;
        RECT 12.608 12.648 12.64 15.156 ;
  LAYER M1 ;
        RECT 12.672 12.648 12.704 15.156 ;
  LAYER M1 ;
        RECT 12.736 12.648 12.768 15.156 ;
  LAYER M1 ;
        RECT 12.8 12.648 12.832 15.156 ;
  LAYER M1 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M1 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M1 ;
        RECT 12.992 12.648 13.024 15.156 ;
  LAYER M1 ;
        RECT 13.056 12.648 13.088 15.156 ;
  LAYER M1 ;
        RECT 13.12 12.648 13.152 15.156 ;
  LAYER M1 ;
        RECT 13.184 12.648 13.216 15.156 ;
  LAYER M1 ;
        RECT 13.248 12.648 13.28 15.156 ;
  LAYER M1 ;
        RECT 13.312 12.648 13.344 15.156 ;
  LAYER M1 ;
        RECT 13.376 12.648 13.408 15.156 ;
  LAYER M1 ;
        RECT 13.44 12.648 13.472 15.156 ;
  LAYER M1 ;
        RECT 13.504 12.648 13.536 15.156 ;
  LAYER M1 ;
        RECT 13.568 12.648 13.6 15.156 ;
  LAYER M1 ;
        RECT 13.632 12.648 13.664 15.156 ;
  LAYER M1 ;
        RECT 13.696 12.648 13.728 15.156 ;
  LAYER M1 ;
        RECT 13.76 12.648 13.792 15.156 ;
  LAYER M1 ;
        RECT 13.824 12.648 13.856 15.156 ;
  LAYER M1 ;
        RECT 13.888 12.648 13.92 15.156 ;
  LAYER M1 ;
        RECT 13.952 12.648 13.984 15.156 ;
  LAYER M1 ;
        RECT 14.016 12.648 14.048 15.156 ;
  LAYER M1 ;
        RECT 14.08 12.648 14.112 15.156 ;
  LAYER M1 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M1 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M2 ;
        RECT 11.884 12.732 14.356 12.764 ;
  LAYER M2 ;
        RECT 11.884 12.796 14.356 12.828 ;
  LAYER M2 ;
        RECT 11.884 12.86 14.356 12.892 ;
  LAYER M2 ;
        RECT 11.884 12.924 14.356 12.956 ;
  LAYER M2 ;
        RECT 11.884 12.988 14.356 13.02 ;
  LAYER M2 ;
        RECT 11.884 13.052 14.356 13.084 ;
  LAYER M2 ;
        RECT 11.884 13.116 14.356 13.148 ;
  LAYER M2 ;
        RECT 11.884 13.18 14.356 13.212 ;
  LAYER M2 ;
        RECT 11.884 13.244 14.356 13.276 ;
  LAYER M2 ;
        RECT 11.884 13.308 14.356 13.34 ;
  LAYER M2 ;
        RECT 11.884 13.372 14.356 13.404 ;
  LAYER M2 ;
        RECT 11.884 13.436 14.356 13.468 ;
  LAYER M2 ;
        RECT 11.884 13.5 14.356 13.532 ;
  LAYER M2 ;
        RECT 11.884 13.564 14.356 13.596 ;
  LAYER M2 ;
        RECT 11.884 13.628 14.356 13.66 ;
  LAYER M2 ;
        RECT 11.884 13.692 14.356 13.724 ;
  LAYER M2 ;
        RECT 11.884 13.756 14.356 13.788 ;
  LAYER M2 ;
        RECT 11.884 13.82 14.356 13.852 ;
  LAYER M2 ;
        RECT 11.884 13.884 14.356 13.916 ;
  LAYER M2 ;
        RECT 11.884 13.948 14.356 13.98 ;
  LAYER M2 ;
        RECT 11.884 14.012 14.356 14.044 ;
  LAYER M2 ;
        RECT 11.884 14.076 14.356 14.108 ;
  LAYER M2 ;
        RECT 11.884 14.14 14.356 14.172 ;
  LAYER M2 ;
        RECT 11.884 14.204 14.356 14.236 ;
  LAYER M2 ;
        RECT 11.884 14.268 14.356 14.3 ;
  LAYER M2 ;
        RECT 11.884 14.332 14.356 14.364 ;
  LAYER M2 ;
        RECT 11.884 14.396 14.356 14.428 ;
  LAYER M2 ;
        RECT 11.884 14.46 14.356 14.492 ;
  LAYER M2 ;
        RECT 11.884 14.524 14.356 14.556 ;
  LAYER M2 ;
        RECT 11.884 14.588 14.356 14.62 ;
  LAYER M2 ;
        RECT 11.884 14.652 14.356 14.684 ;
  LAYER M2 ;
        RECT 11.884 14.716 14.356 14.748 ;
  LAYER M2 ;
        RECT 11.884 14.78 14.356 14.812 ;
  LAYER M2 ;
        RECT 11.884 14.844 14.356 14.876 ;
  LAYER M2 ;
        RECT 11.884 14.908 14.356 14.94 ;
  LAYER M2 ;
        RECT 11.884 14.972 14.356 15.004 ;
  LAYER M3 ;
        RECT 11.904 12.648 11.936 15.156 ;
  LAYER M3 ;
        RECT 11.968 12.648 12 15.156 ;
  LAYER M3 ;
        RECT 12.032 12.648 12.064 15.156 ;
  LAYER M3 ;
        RECT 12.096 12.648 12.128 15.156 ;
  LAYER M3 ;
        RECT 12.16 12.648 12.192 15.156 ;
  LAYER M3 ;
        RECT 12.224 12.648 12.256 15.156 ;
  LAYER M3 ;
        RECT 12.288 12.648 12.32 15.156 ;
  LAYER M3 ;
        RECT 12.352 12.648 12.384 15.156 ;
  LAYER M3 ;
        RECT 12.416 12.648 12.448 15.156 ;
  LAYER M3 ;
        RECT 12.48 12.648 12.512 15.156 ;
  LAYER M3 ;
        RECT 12.544 12.648 12.576 15.156 ;
  LAYER M3 ;
        RECT 12.608 12.648 12.64 15.156 ;
  LAYER M3 ;
        RECT 12.672 12.648 12.704 15.156 ;
  LAYER M3 ;
        RECT 12.736 12.648 12.768 15.156 ;
  LAYER M3 ;
        RECT 12.8 12.648 12.832 15.156 ;
  LAYER M3 ;
        RECT 12.864 12.648 12.896 15.156 ;
  LAYER M3 ;
        RECT 12.928 12.648 12.96 15.156 ;
  LAYER M3 ;
        RECT 12.992 12.648 13.024 15.156 ;
  LAYER M3 ;
        RECT 13.056 12.648 13.088 15.156 ;
  LAYER M3 ;
        RECT 13.12 12.648 13.152 15.156 ;
  LAYER M3 ;
        RECT 13.184 12.648 13.216 15.156 ;
  LAYER M3 ;
        RECT 13.248 12.648 13.28 15.156 ;
  LAYER M3 ;
        RECT 13.312 12.648 13.344 15.156 ;
  LAYER M3 ;
        RECT 13.376 12.648 13.408 15.156 ;
  LAYER M3 ;
        RECT 13.44 12.648 13.472 15.156 ;
  LAYER M3 ;
        RECT 13.504 12.648 13.536 15.156 ;
  LAYER M3 ;
        RECT 13.568 12.648 13.6 15.156 ;
  LAYER M3 ;
        RECT 13.632 12.648 13.664 15.156 ;
  LAYER M3 ;
        RECT 13.696 12.648 13.728 15.156 ;
  LAYER M3 ;
        RECT 13.76 12.648 13.792 15.156 ;
  LAYER M3 ;
        RECT 13.824 12.648 13.856 15.156 ;
  LAYER M3 ;
        RECT 13.888 12.648 13.92 15.156 ;
  LAYER M3 ;
        RECT 13.952 12.648 13.984 15.156 ;
  LAYER M3 ;
        RECT 14.016 12.648 14.048 15.156 ;
  LAYER M3 ;
        RECT 14.08 12.648 14.112 15.156 ;
  LAYER M3 ;
        RECT 14.144 12.648 14.176 15.156 ;
  LAYER M3 ;
        RECT 14.208 12.648 14.24 15.156 ;
  LAYER M3 ;
        RECT 14.304 12.648 14.336 15.156 ;
  LAYER M1 ;
        RECT 11.919 12.684 11.921 15.12 ;
  LAYER M1 ;
        RECT 11.999 12.684 12.001 15.12 ;
  LAYER M1 ;
        RECT 12.079 12.684 12.081 15.12 ;
  LAYER M1 ;
        RECT 12.159 12.684 12.161 15.12 ;
  LAYER M1 ;
        RECT 12.239 12.684 12.241 15.12 ;
  LAYER M1 ;
        RECT 12.319 12.684 12.321 15.12 ;
  LAYER M1 ;
        RECT 12.399 12.684 12.401 15.12 ;
  LAYER M1 ;
        RECT 12.479 12.684 12.481 15.12 ;
  LAYER M1 ;
        RECT 12.559 12.684 12.561 15.12 ;
  LAYER M1 ;
        RECT 12.639 12.684 12.641 15.12 ;
  LAYER M1 ;
        RECT 12.719 12.684 12.721 15.12 ;
  LAYER M1 ;
        RECT 12.799 12.684 12.801 15.12 ;
  LAYER M1 ;
        RECT 12.879 12.684 12.881 15.12 ;
  LAYER M1 ;
        RECT 12.959 12.684 12.961 15.12 ;
  LAYER M1 ;
        RECT 13.039 12.684 13.041 15.12 ;
  LAYER M1 ;
        RECT 13.119 12.684 13.121 15.12 ;
  LAYER M1 ;
        RECT 13.199 12.684 13.201 15.12 ;
  LAYER M1 ;
        RECT 13.279 12.684 13.281 15.12 ;
  LAYER M1 ;
        RECT 13.359 12.684 13.361 15.12 ;
  LAYER M1 ;
        RECT 13.439 12.684 13.441 15.12 ;
  LAYER M1 ;
        RECT 13.519 12.684 13.521 15.12 ;
  LAYER M1 ;
        RECT 13.599 12.684 13.601 15.12 ;
  LAYER M1 ;
        RECT 13.679 12.684 13.681 15.12 ;
  LAYER M1 ;
        RECT 13.759 12.684 13.761 15.12 ;
  LAYER M1 ;
        RECT 13.839 12.684 13.841 15.12 ;
  LAYER M1 ;
        RECT 13.919 12.684 13.921 15.12 ;
  LAYER M1 ;
        RECT 13.999 12.684 14.001 15.12 ;
  LAYER M1 ;
        RECT 14.079 12.684 14.081 15.12 ;
  LAYER M1 ;
        RECT 14.159 12.684 14.161 15.12 ;
  LAYER M1 ;
        RECT 14.239 12.684 14.241 15.12 ;
  LAYER M2 ;
        RECT 11.92 12.683 14.32 12.685 ;
  LAYER M2 ;
        RECT 11.92 12.767 14.32 12.769 ;
  LAYER M2 ;
        RECT 11.92 12.851 14.32 12.853 ;
  LAYER M2 ;
        RECT 11.92 12.935 14.32 12.937 ;
  LAYER M2 ;
        RECT 11.92 13.019 14.32 13.021 ;
  LAYER M2 ;
        RECT 11.92 13.103 14.32 13.105 ;
  LAYER M2 ;
        RECT 11.92 13.187 14.32 13.189 ;
  LAYER M2 ;
        RECT 11.92 13.271 14.32 13.273 ;
  LAYER M2 ;
        RECT 11.92 13.355 14.32 13.357 ;
  LAYER M2 ;
        RECT 11.92 13.439 14.32 13.441 ;
  LAYER M2 ;
        RECT 11.92 13.523 14.32 13.525 ;
  LAYER M2 ;
        RECT 11.92 13.607 14.32 13.609 ;
  LAYER M2 ;
        RECT 11.92 13.6905 14.32 13.6925 ;
  LAYER M2 ;
        RECT 11.92 13.775 14.32 13.777 ;
  LAYER M2 ;
        RECT 11.92 13.859 14.32 13.861 ;
  LAYER M2 ;
        RECT 11.92 13.943 14.32 13.945 ;
  LAYER M2 ;
        RECT 11.92 14.027 14.32 14.029 ;
  LAYER M2 ;
        RECT 11.92 14.111 14.32 14.113 ;
  LAYER M2 ;
        RECT 11.92 14.195 14.32 14.197 ;
  LAYER M2 ;
        RECT 11.92 14.279 14.32 14.281 ;
  LAYER M2 ;
        RECT 11.92 14.363 14.32 14.365 ;
  LAYER M2 ;
        RECT 11.92 14.447 14.32 14.449 ;
  LAYER M2 ;
        RECT 11.92 14.531 14.32 14.533 ;
  LAYER M2 ;
        RECT 11.92 14.615 14.32 14.617 ;
  LAYER M2 ;
        RECT 11.92 14.699 14.32 14.701 ;
  LAYER M2 ;
        RECT 11.92 14.783 14.32 14.785 ;
  LAYER M2 ;
        RECT 11.92 14.867 14.32 14.869 ;
  LAYER M2 ;
        RECT 11.92 14.951 14.32 14.953 ;
  LAYER M2 ;
        RECT 11.92 15.035 14.32 15.037 ;
  LAYER M1 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M1 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M1 ;
        RECT 12.032 15.588 12.064 18.096 ;
  LAYER M1 ;
        RECT 12.096 15.588 12.128 18.096 ;
  LAYER M1 ;
        RECT 12.16 15.588 12.192 18.096 ;
  LAYER M1 ;
        RECT 12.224 15.588 12.256 18.096 ;
  LAYER M1 ;
        RECT 12.288 15.588 12.32 18.096 ;
  LAYER M1 ;
        RECT 12.352 15.588 12.384 18.096 ;
  LAYER M1 ;
        RECT 12.416 15.588 12.448 18.096 ;
  LAYER M1 ;
        RECT 12.48 15.588 12.512 18.096 ;
  LAYER M1 ;
        RECT 12.544 15.588 12.576 18.096 ;
  LAYER M1 ;
        RECT 12.608 15.588 12.64 18.096 ;
  LAYER M1 ;
        RECT 12.672 15.588 12.704 18.096 ;
  LAYER M1 ;
        RECT 12.736 15.588 12.768 18.096 ;
  LAYER M1 ;
        RECT 12.8 15.588 12.832 18.096 ;
  LAYER M1 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M1 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M1 ;
        RECT 12.992 15.588 13.024 18.096 ;
  LAYER M1 ;
        RECT 13.056 15.588 13.088 18.096 ;
  LAYER M1 ;
        RECT 13.12 15.588 13.152 18.096 ;
  LAYER M1 ;
        RECT 13.184 15.588 13.216 18.096 ;
  LAYER M1 ;
        RECT 13.248 15.588 13.28 18.096 ;
  LAYER M1 ;
        RECT 13.312 15.588 13.344 18.096 ;
  LAYER M1 ;
        RECT 13.376 15.588 13.408 18.096 ;
  LAYER M1 ;
        RECT 13.44 15.588 13.472 18.096 ;
  LAYER M1 ;
        RECT 13.504 15.588 13.536 18.096 ;
  LAYER M1 ;
        RECT 13.568 15.588 13.6 18.096 ;
  LAYER M1 ;
        RECT 13.632 15.588 13.664 18.096 ;
  LAYER M1 ;
        RECT 13.696 15.588 13.728 18.096 ;
  LAYER M1 ;
        RECT 13.76 15.588 13.792 18.096 ;
  LAYER M1 ;
        RECT 13.824 15.588 13.856 18.096 ;
  LAYER M1 ;
        RECT 13.888 15.588 13.92 18.096 ;
  LAYER M1 ;
        RECT 13.952 15.588 13.984 18.096 ;
  LAYER M1 ;
        RECT 14.016 15.588 14.048 18.096 ;
  LAYER M1 ;
        RECT 14.08 15.588 14.112 18.096 ;
  LAYER M1 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M1 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M2 ;
        RECT 11.884 15.672 14.356 15.704 ;
  LAYER M2 ;
        RECT 11.884 15.736 14.356 15.768 ;
  LAYER M2 ;
        RECT 11.884 15.8 14.356 15.832 ;
  LAYER M2 ;
        RECT 11.884 15.864 14.356 15.896 ;
  LAYER M2 ;
        RECT 11.884 15.928 14.356 15.96 ;
  LAYER M2 ;
        RECT 11.884 15.992 14.356 16.024 ;
  LAYER M2 ;
        RECT 11.884 16.056 14.356 16.088 ;
  LAYER M2 ;
        RECT 11.884 16.12 14.356 16.152 ;
  LAYER M2 ;
        RECT 11.884 16.184 14.356 16.216 ;
  LAYER M2 ;
        RECT 11.884 16.248 14.356 16.28 ;
  LAYER M2 ;
        RECT 11.884 16.312 14.356 16.344 ;
  LAYER M2 ;
        RECT 11.884 16.376 14.356 16.408 ;
  LAYER M2 ;
        RECT 11.884 16.44 14.356 16.472 ;
  LAYER M2 ;
        RECT 11.884 16.504 14.356 16.536 ;
  LAYER M2 ;
        RECT 11.884 16.568 14.356 16.6 ;
  LAYER M2 ;
        RECT 11.884 16.632 14.356 16.664 ;
  LAYER M2 ;
        RECT 11.884 16.696 14.356 16.728 ;
  LAYER M2 ;
        RECT 11.884 16.76 14.356 16.792 ;
  LAYER M2 ;
        RECT 11.884 16.824 14.356 16.856 ;
  LAYER M2 ;
        RECT 11.884 16.888 14.356 16.92 ;
  LAYER M2 ;
        RECT 11.884 16.952 14.356 16.984 ;
  LAYER M2 ;
        RECT 11.884 17.016 14.356 17.048 ;
  LAYER M2 ;
        RECT 11.884 17.08 14.356 17.112 ;
  LAYER M2 ;
        RECT 11.884 17.144 14.356 17.176 ;
  LAYER M2 ;
        RECT 11.884 17.208 14.356 17.24 ;
  LAYER M2 ;
        RECT 11.884 17.272 14.356 17.304 ;
  LAYER M2 ;
        RECT 11.884 17.336 14.356 17.368 ;
  LAYER M2 ;
        RECT 11.884 17.4 14.356 17.432 ;
  LAYER M2 ;
        RECT 11.884 17.464 14.356 17.496 ;
  LAYER M2 ;
        RECT 11.884 17.528 14.356 17.56 ;
  LAYER M2 ;
        RECT 11.884 17.592 14.356 17.624 ;
  LAYER M2 ;
        RECT 11.884 17.656 14.356 17.688 ;
  LAYER M2 ;
        RECT 11.884 17.72 14.356 17.752 ;
  LAYER M2 ;
        RECT 11.884 17.784 14.356 17.816 ;
  LAYER M2 ;
        RECT 11.884 17.848 14.356 17.88 ;
  LAYER M2 ;
        RECT 11.884 17.912 14.356 17.944 ;
  LAYER M3 ;
        RECT 11.904 15.588 11.936 18.096 ;
  LAYER M3 ;
        RECT 11.968 15.588 12 18.096 ;
  LAYER M3 ;
        RECT 12.032 15.588 12.064 18.096 ;
  LAYER M3 ;
        RECT 12.096 15.588 12.128 18.096 ;
  LAYER M3 ;
        RECT 12.16 15.588 12.192 18.096 ;
  LAYER M3 ;
        RECT 12.224 15.588 12.256 18.096 ;
  LAYER M3 ;
        RECT 12.288 15.588 12.32 18.096 ;
  LAYER M3 ;
        RECT 12.352 15.588 12.384 18.096 ;
  LAYER M3 ;
        RECT 12.416 15.588 12.448 18.096 ;
  LAYER M3 ;
        RECT 12.48 15.588 12.512 18.096 ;
  LAYER M3 ;
        RECT 12.544 15.588 12.576 18.096 ;
  LAYER M3 ;
        RECT 12.608 15.588 12.64 18.096 ;
  LAYER M3 ;
        RECT 12.672 15.588 12.704 18.096 ;
  LAYER M3 ;
        RECT 12.736 15.588 12.768 18.096 ;
  LAYER M3 ;
        RECT 12.8 15.588 12.832 18.096 ;
  LAYER M3 ;
        RECT 12.864 15.588 12.896 18.096 ;
  LAYER M3 ;
        RECT 12.928 15.588 12.96 18.096 ;
  LAYER M3 ;
        RECT 12.992 15.588 13.024 18.096 ;
  LAYER M3 ;
        RECT 13.056 15.588 13.088 18.096 ;
  LAYER M3 ;
        RECT 13.12 15.588 13.152 18.096 ;
  LAYER M3 ;
        RECT 13.184 15.588 13.216 18.096 ;
  LAYER M3 ;
        RECT 13.248 15.588 13.28 18.096 ;
  LAYER M3 ;
        RECT 13.312 15.588 13.344 18.096 ;
  LAYER M3 ;
        RECT 13.376 15.588 13.408 18.096 ;
  LAYER M3 ;
        RECT 13.44 15.588 13.472 18.096 ;
  LAYER M3 ;
        RECT 13.504 15.588 13.536 18.096 ;
  LAYER M3 ;
        RECT 13.568 15.588 13.6 18.096 ;
  LAYER M3 ;
        RECT 13.632 15.588 13.664 18.096 ;
  LAYER M3 ;
        RECT 13.696 15.588 13.728 18.096 ;
  LAYER M3 ;
        RECT 13.76 15.588 13.792 18.096 ;
  LAYER M3 ;
        RECT 13.824 15.588 13.856 18.096 ;
  LAYER M3 ;
        RECT 13.888 15.588 13.92 18.096 ;
  LAYER M3 ;
        RECT 13.952 15.588 13.984 18.096 ;
  LAYER M3 ;
        RECT 14.016 15.588 14.048 18.096 ;
  LAYER M3 ;
        RECT 14.08 15.588 14.112 18.096 ;
  LAYER M3 ;
        RECT 14.144 15.588 14.176 18.096 ;
  LAYER M3 ;
        RECT 14.208 15.588 14.24 18.096 ;
  LAYER M3 ;
        RECT 14.304 15.588 14.336 18.096 ;
  LAYER M1 ;
        RECT 11.919 15.624 11.921 18.06 ;
  LAYER M1 ;
        RECT 11.999 15.624 12.001 18.06 ;
  LAYER M1 ;
        RECT 12.079 15.624 12.081 18.06 ;
  LAYER M1 ;
        RECT 12.159 15.624 12.161 18.06 ;
  LAYER M1 ;
        RECT 12.239 15.624 12.241 18.06 ;
  LAYER M1 ;
        RECT 12.319 15.624 12.321 18.06 ;
  LAYER M1 ;
        RECT 12.399 15.624 12.401 18.06 ;
  LAYER M1 ;
        RECT 12.479 15.624 12.481 18.06 ;
  LAYER M1 ;
        RECT 12.559 15.624 12.561 18.06 ;
  LAYER M1 ;
        RECT 12.639 15.624 12.641 18.06 ;
  LAYER M1 ;
        RECT 12.719 15.624 12.721 18.06 ;
  LAYER M1 ;
        RECT 12.799 15.624 12.801 18.06 ;
  LAYER M1 ;
        RECT 12.879 15.624 12.881 18.06 ;
  LAYER M1 ;
        RECT 12.959 15.624 12.961 18.06 ;
  LAYER M1 ;
        RECT 13.039 15.624 13.041 18.06 ;
  LAYER M1 ;
        RECT 13.119 15.624 13.121 18.06 ;
  LAYER M1 ;
        RECT 13.199 15.624 13.201 18.06 ;
  LAYER M1 ;
        RECT 13.279 15.624 13.281 18.06 ;
  LAYER M1 ;
        RECT 13.359 15.624 13.361 18.06 ;
  LAYER M1 ;
        RECT 13.439 15.624 13.441 18.06 ;
  LAYER M1 ;
        RECT 13.519 15.624 13.521 18.06 ;
  LAYER M1 ;
        RECT 13.599 15.624 13.601 18.06 ;
  LAYER M1 ;
        RECT 13.679 15.624 13.681 18.06 ;
  LAYER M1 ;
        RECT 13.759 15.624 13.761 18.06 ;
  LAYER M1 ;
        RECT 13.839 15.624 13.841 18.06 ;
  LAYER M1 ;
        RECT 13.919 15.624 13.921 18.06 ;
  LAYER M1 ;
        RECT 13.999 15.624 14.001 18.06 ;
  LAYER M1 ;
        RECT 14.079 15.624 14.081 18.06 ;
  LAYER M1 ;
        RECT 14.159 15.624 14.161 18.06 ;
  LAYER M1 ;
        RECT 14.239 15.624 14.241 18.06 ;
  LAYER M2 ;
        RECT 11.92 15.623 14.32 15.625 ;
  LAYER M2 ;
        RECT 11.92 15.707 14.32 15.709 ;
  LAYER M2 ;
        RECT 11.92 15.791 14.32 15.793 ;
  LAYER M2 ;
        RECT 11.92 15.875 14.32 15.877 ;
  LAYER M2 ;
        RECT 11.92 15.959 14.32 15.961 ;
  LAYER M2 ;
        RECT 11.92 16.043 14.32 16.045 ;
  LAYER M2 ;
        RECT 11.92 16.127 14.32 16.129 ;
  LAYER M2 ;
        RECT 11.92 16.211 14.32 16.213 ;
  LAYER M2 ;
        RECT 11.92 16.295 14.32 16.297 ;
  LAYER M2 ;
        RECT 11.92 16.379 14.32 16.381 ;
  LAYER M2 ;
        RECT 11.92 16.463 14.32 16.465 ;
  LAYER M2 ;
        RECT 11.92 16.547 14.32 16.549 ;
  LAYER M2 ;
        RECT 11.92 16.6305 14.32 16.6325 ;
  LAYER M2 ;
        RECT 11.92 16.715 14.32 16.717 ;
  LAYER M2 ;
        RECT 11.92 16.799 14.32 16.801 ;
  LAYER M2 ;
        RECT 11.92 16.883 14.32 16.885 ;
  LAYER M2 ;
        RECT 11.92 16.967 14.32 16.969 ;
  LAYER M2 ;
        RECT 11.92 17.051 14.32 17.053 ;
  LAYER M2 ;
        RECT 11.92 17.135 14.32 17.137 ;
  LAYER M2 ;
        RECT 11.92 17.219 14.32 17.221 ;
  LAYER M2 ;
        RECT 11.92 17.303 14.32 17.305 ;
  LAYER M2 ;
        RECT 11.92 17.387 14.32 17.389 ;
  LAYER M2 ;
        RECT 11.92 17.471 14.32 17.473 ;
  LAYER M2 ;
        RECT 11.92 17.555 14.32 17.557 ;
  LAYER M2 ;
        RECT 11.92 17.639 14.32 17.641 ;
  LAYER M2 ;
        RECT 11.92 17.723 14.32 17.725 ;
  LAYER M2 ;
        RECT 11.92 17.807 14.32 17.809 ;
  LAYER M2 ;
        RECT 11.92 17.891 14.32 17.893 ;
  LAYER M2 ;
        RECT 11.92 17.975 14.32 17.977 ;
  END 
END Cap_60fF_Cap_60fF
