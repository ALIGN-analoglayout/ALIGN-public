MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 15.36 BY 21.924 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
      LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
      LAYER M1 ;
        RECT 12.384 21.468 12.416 21.54 ;
      LAYER M2 ;
        RECT 12.364 21.488 12.436 21.52 ;
      LAYER M2 ;
        RECT 2.8 21.488 12.4 21.52 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
      LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
      LAYER M1 ;
        RECT 9.024 0.384 9.056 0.456 ;
      LAYER M2 ;
        RECT 9.004 0.404 9.076 0.436 ;
      LAYER M2 ;
        RECT 5.84 0.404 9.04 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.144 21.636 6.176 21.708 ;
      LAYER M2 ;
        RECT 6.124 21.656 6.196 21.688 ;
      LAYER M1 ;
        RECT 9.344 21.636 9.376 21.708 ;
      LAYER M2 ;
        RECT 9.324 21.656 9.396 21.688 ;
      LAYER M2 ;
        RECT 6.16 21.656 9.36 21.688 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.624 0.216 2.656 0.288 ;
      LAYER M2 ;
        RECT 2.604 0.236 2.676 0.268 ;
      LAYER M1 ;
        RECT 12.224 0.216 12.256 0.288 ;
      LAYER M2 ;
        RECT 12.204 0.236 12.276 0.268 ;
      LAYER M2 ;
        RECT 2.64 0.236 12.24 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.864 6.768 8.896 6.84 ;
  LAYER M2 ;
        RECT 8.844 6.788 8.916 6.82 ;
  LAYER M2 ;
        RECT 5.84 6.788 8.88 6.82 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 6.84 ;
  LAYER M2 ;
        RECT 5.804 6.788 5.876 6.82 ;
  LAYER M1 ;
        RECT 8.864 12.648 8.896 12.72 ;
  LAYER M2 ;
        RECT 8.844 12.668 8.916 12.7 ;
  LAYER M2 ;
        RECT 5.84 12.668 8.88 12.7 ;
  LAYER M1 ;
        RECT 5.824 12.648 5.856 12.72 ;
  LAYER M2 ;
        RECT 5.804 12.668 5.876 12.7 ;
  LAYER M1 ;
        RECT 5.664 9.708 5.696 9.78 ;
  LAYER M2 ;
        RECT 5.644 9.728 5.716 9.76 ;
  LAYER M1 ;
        RECT 5.664 9.576 5.696 9.744 ;
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M2 ;
        RECT 5.68 9.56 5.84 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 5.664 6.768 5.696 6.84 ;
  LAYER M2 ;
        RECT 5.644 6.788 5.716 6.82 ;
  LAYER M1 ;
        RECT 5.664 6.636 5.696 6.804 ;
  LAYER M1 ;
        RECT 5.664 6.6 5.696 6.672 ;
  LAYER M2 ;
        RECT 5.644 6.62 5.716 6.652 ;
  LAYER M2 ;
        RECT 5.68 6.62 5.84 6.652 ;
  LAYER M1 ;
        RECT 5.824 6.6 5.856 6.672 ;
  LAYER M2 ;
        RECT 5.804 6.62 5.876 6.652 ;
  LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
  LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 0.588 ;
  LAYER M1 ;
        RECT 5.824 0.588 5.856 12.684 ;
  LAYER M1 ;
        RECT 12.064 9.708 12.096 9.78 ;
  LAYER M2 ;
        RECT 12.044 9.728 12.116 9.76 ;
  LAYER M2 ;
        RECT 9.04 9.728 12.08 9.76 ;
  LAYER M1 ;
        RECT 9.024 9.708 9.056 9.78 ;
  LAYER M2 ;
        RECT 9.004 9.728 9.076 9.76 ;
  LAYER M1 ;
        RECT 12.064 12.648 12.096 12.72 ;
  LAYER M2 ;
        RECT 12.044 12.668 12.116 12.7 ;
  LAYER M2 ;
        RECT 9.04 12.668 12.08 12.7 ;
  LAYER M1 ;
        RECT 9.024 12.648 9.056 12.72 ;
  LAYER M2 ;
        RECT 9.004 12.668 9.076 12.7 ;
  LAYER M1 ;
        RECT 9.024 0.384 9.056 0.456 ;
  LAYER M2 ;
        RECT 9.004 0.404 9.076 0.436 ;
  LAYER M1 ;
        RECT 9.024 0.42 9.056 0.588 ;
  LAYER M1 ;
        RECT 9.024 0.588 9.056 12.684 ;
  LAYER M2 ;
        RECT 5.84 0.404 9.04 0.436 ;
  LAYER M1 ;
        RECT 5.664 12.648 5.696 12.72 ;
  LAYER M2 ;
        RECT 5.644 12.668 5.716 12.7 ;
  LAYER M2 ;
        RECT 2.64 12.668 5.68 12.7 ;
  LAYER M1 ;
        RECT 2.624 12.648 2.656 12.72 ;
  LAYER M2 ;
        RECT 2.604 12.668 2.676 12.7 ;
  LAYER M1 ;
        RECT 5.664 15.588 5.696 15.66 ;
  LAYER M2 ;
        RECT 5.644 15.608 5.716 15.64 ;
  LAYER M2 ;
        RECT 2.64 15.608 5.68 15.64 ;
  LAYER M1 ;
        RECT 2.624 15.588 2.656 15.66 ;
  LAYER M2 ;
        RECT 2.604 15.608 2.676 15.64 ;
  LAYER M1 ;
        RECT 2.624 0.216 2.656 0.288 ;
  LAYER M2 ;
        RECT 2.604 0.236 2.676 0.268 ;
  LAYER M1 ;
        RECT 2.624 0.252 2.656 0.588 ;
  LAYER M1 ;
        RECT 2.624 0.588 2.656 15.624 ;
  LAYER M1 ;
        RECT 12.064 6.768 12.096 6.84 ;
  LAYER M2 ;
        RECT 12.044 6.788 12.116 6.82 ;
  LAYER M1 ;
        RECT 12.064 6.636 12.096 6.804 ;
  LAYER M1 ;
        RECT 12.064 6.6 12.096 6.672 ;
  LAYER M2 ;
        RECT 12.044 6.62 12.116 6.652 ;
  LAYER M2 ;
        RECT 12.08 6.62 12.24 6.652 ;
  LAYER M1 ;
        RECT 12.224 6.6 12.256 6.672 ;
  LAYER M2 ;
        RECT 12.204 6.62 12.276 6.652 ;
  LAYER M1 ;
        RECT 12.064 3.828 12.096 3.9 ;
  LAYER M2 ;
        RECT 12.044 3.848 12.116 3.88 ;
  LAYER M1 ;
        RECT 12.064 3.696 12.096 3.864 ;
  LAYER M1 ;
        RECT 12.064 3.66 12.096 3.732 ;
  LAYER M2 ;
        RECT 12.044 3.68 12.116 3.712 ;
  LAYER M2 ;
        RECT 12.08 3.68 12.24 3.712 ;
  LAYER M1 ;
        RECT 12.224 3.66 12.256 3.732 ;
  LAYER M2 ;
        RECT 12.204 3.68 12.276 3.712 ;
  LAYER M1 ;
        RECT 12.224 0.216 12.256 0.288 ;
  LAYER M2 ;
        RECT 12.204 0.236 12.276 0.268 ;
  LAYER M1 ;
        RECT 12.224 0.252 12.256 0.588 ;
  LAYER M1 ;
        RECT 12.224 0.588 12.256 6.636 ;
  LAYER M2 ;
        RECT 2.64 0.236 12.24 0.268 ;
  LAYER M1 ;
        RECT 8.864 15.588 8.896 15.66 ;
  LAYER M2 ;
        RECT 8.844 15.608 8.916 15.64 ;
  LAYER M2 ;
        RECT 5.68 15.608 8.88 15.64 ;
  LAYER M1 ;
        RECT 5.664 15.588 5.696 15.66 ;
  LAYER M2 ;
        RECT 5.644 15.608 5.716 15.64 ;
  LAYER M1 ;
        RECT 8.864 3.828 8.896 3.9 ;
  LAYER M2 ;
        RECT 8.844 3.848 8.916 3.88 ;
  LAYER M2 ;
        RECT 8.88 3.848 12.08 3.88 ;
  LAYER M1 ;
        RECT 12.064 3.828 12.096 3.9 ;
  LAYER M2 ;
        RECT 12.044 3.848 12.116 3.88 ;
  LAYER M1 ;
        RECT 5.664 0.888 5.696 0.96 ;
  LAYER M2 ;
        RECT 5.644 0.908 5.716 0.94 ;
  LAYER M1 ;
        RECT 5.664 0.756 5.696 0.924 ;
  LAYER M1 ;
        RECT 5.664 0.72 5.696 0.792 ;
  LAYER M2 ;
        RECT 5.644 0.74 5.716 0.772 ;
  LAYER M2 ;
        RECT 5.68 0.74 6 0.772 ;
  LAYER M1 ;
        RECT 5.984 0.72 6.016 0.792 ;
  LAYER M2 ;
        RECT 5.964 0.74 6.036 0.772 ;
  LAYER M1 ;
        RECT 5.664 3.828 5.696 3.9 ;
  LAYER M2 ;
        RECT 5.644 3.848 5.716 3.88 ;
  LAYER M1 ;
        RECT 5.664 3.696 5.696 3.864 ;
  LAYER M1 ;
        RECT 5.664 3.66 5.696 3.732 ;
  LAYER M2 ;
        RECT 5.644 3.68 5.716 3.712 ;
  LAYER M2 ;
        RECT 5.68 3.68 6 3.712 ;
  LAYER M1 ;
        RECT 5.984 3.66 6.016 3.732 ;
  LAYER M2 ;
        RECT 5.964 3.68 6.036 3.712 ;
  LAYER M1 ;
        RECT 5.664 18.528 5.696 18.6 ;
  LAYER M2 ;
        RECT 5.644 18.548 5.716 18.58 ;
  LAYER M1 ;
        RECT 5.664 18.396 5.696 18.564 ;
  LAYER M1 ;
        RECT 5.664 18.36 5.696 18.432 ;
  LAYER M2 ;
        RECT 5.644 18.38 5.716 18.412 ;
  LAYER M2 ;
        RECT 5.68 18.38 6 18.412 ;
  LAYER M1 ;
        RECT 5.984 18.36 6.016 18.432 ;
  LAYER M2 ;
        RECT 5.964 18.38 6.036 18.412 ;
  LAYER M1 ;
        RECT 8.864 0.888 8.896 0.96 ;
  LAYER M2 ;
        RECT 8.844 0.908 8.916 0.94 ;
  LAYER M2 ;
        RECT 6 0.908 8.88 0.94 ;
  LAYER M1 ;
        RECT 5.984 0.888 6.016 0.96 ;
  LAYER M2 ;
        RECT 5.964 0.908 6.036 0.94 ;
  LAYER M1 ;
        RECT 8.864 9.708 8.896 9.78 ;
  LAYER M2 ;
        RECT 8.844 9.728 8.916 9.76 ;
  LAYER M2 ;
        RECT 6 9.728 8.88 9.76 ;
  LAYER M1 ;
        RECT 5.984 9.708 6.016 9.78 ;
  LAYER M2 ;
        RECT 5.964 9.728 6.036 9.76 ;
  LAYER M1 ;
        RECT 8.864 18.528 8.896 18.6 ;
  LAYER M2 ;
        RECT 8.844 18.548 8.916 18.58 ;
  LAYER M2 ;
        RECT 6 18.548 8.88 18.58 ;
  LAYER M1 ;
        RECT 5.984 18.528 6.016 18.6 ;
  LAYER M2 ;
        RECT 5.964 18.548 6.036 18.58 ;
  LAYER M1 ;
        RECT 5.984 0.048 6.016 0.12 ;
  LAYER M2 ;
        RECT 5.964 0.068 6.036 0.1 ;
  LAYER M1 ;
        RECT 5.984 0.084 6.016 0.588 ;
  LAYER M1 ;
        RECT 5.984 0.588 6.016 18.564 ;
  LAYER M1 ;
        RECT 12.064 0.888 12.096 0.96 ;
  LAYER M2 ;
        RECT 12.044 0.908 12.116 0.94 ;
  LAYER M2 ;
        RECT 9.2 0.908 12.08 0.94 ;
  LAYER M1 ;
        RECT 9.184 0.888 9.216 0.96 ;
  LAYER M2 ;
        RECT 9.164 0.908 9.236 0.94 ;
  LAYER M1 ;
        RECT 12.064 15.588 12.096 15.66 ;
  LAYER M2 ;
        RECT 12.044 15.608 12.116 15.64 ;
  LAYER M2 ;
        RECT 9.2 15.608 12.08 15.64 ;
  LAYER M1 ;
        RECT 9.184 15.588 9.216 15.66 ;
  LAYER M2 ;
        RECT 9.164 15.608 9.236 15.64 ;
  LAYER M1 ;
        RECT 12.064 18.528 12.096 18.6 ;
  LAYER M2 ;
        RECT 12.044 18.548 12.116 18.58 ;
  LAYER M2 ;
        RECT 9.2 18.548 12.08 18.58 ;
  LAYER M1 ;
        RECT 9.184 18.528 9.216 18.6 ;
  LAYER M2 ;
        RECT 9.164 18.548 9.236 18.58 ;
  LAYER M1 ;
        RECT 9.184 0.048 9.216 0.12 ;
  LAYER M2 ;
        RECT 9.164 0.068 9.236 0.1 ;
  LAYER M1 ;
        RECT 9.184 0.084 9.216 0.588 ;
  LAYER M1 ;
        RECT 9.184 0.588 9.216 18.564 ;
  LAYER M2 ;
        RECT 6 0.068 9.2 0.1 ;
  LAYER M1 ;
        RECT 2.464 18.528 2.496 18.6 ;
  LAYER M2 ;
        RECT 2.444 18.548 2.516 18.58 ;
  LAYER M2 ;
        RECT 2.48 18.548 5.68 18.58 ;
  LAYER M1 ;
        RECT 5.664 18.528 5.696 18.6 ;
  LAYER M2 ;
        RECT 5.644 18.548 5.716 18.58 ;
  LAYER M1 ;
        RECT 2.464 15.588 2.496 15.66 ;
  LAYER M2 ;
        RECT 2.444 15.608 2.516 15.64 ;
  LAYER M1 ;
        RECT 2.464 15.624 2.496 18.564 ;
  LAYER M1 ;
        RECT 2.464 18.528 2.496 18.6 ;
  LAYER M2 ;
        RECT 2.444 18.548 2.516 18.58 ;
  LAYER M1 ;
        RECT 2.464 12.648 2.496 12.72 ;
  LAYER M2 ;
        RECT 2.444 12.668 2.516 12.7 ;
  LAYER M1 ;
        RECT 2.464 12.684 2.496 15.624 ;
  LAYER M1 ;
        RECT 2.464 15.588 2.496 15.66 ;
  LAYER M2 ;
        RECT 2.444 15.608 2.516 15.64 ;
  LAYER M1 ;
        RECT 2.464 9.708 2.496 9.78 ;
  LAYER M2 ;
        RECT 2.444 9.728 2.516 9.76 ;
  LAYER M1 ;
        RECT 2.464 9.744 2.496 12.684 ;
  LAYER M1 ;
        RECT 2.464 12.648 2.496 12.72 ;
  LAYER M2 ;
        RECT 2.444 12.668 2.516 12.7 ;
  LAYER M1 ;
        RECT 2.464 6.768 2.496 6.84 ;
  LAYER M2 ;
        RECT 2.444 6.788 2.516 6.82 ;
  LAYER M1 ;
        RECT 2.464 6.804 2.496 9.744 ;
  LAYER M1 ;
        RECT 2.464 9.708 2.496 9.78 ;
  LAYER M2 ;
        RECT 2.444 9.728 2.516 9.76 ;
  LAYER M1 ;
        RECT 2.464 3.828 2.496 3.9 ;
  LAYER M2 ;
        RECT 2.444 3.848 2.516 3.88 ;
  LAYER M1 ;
        RECT 2.464 3.864 2.496 6.804 ;
  LAYER M1 ;
        RECT 2.464 6.768 2.496 6.84 ;
  LAYER M2 ;
        RECT 2.444 6.788 2.516 6.82 ;
  LAYER M1 ;
        RECT 2.464 0.888 2.496 0.96 ;
  LAYER M2 ;
        RECT 2.444 0.908 2.516 0.94 ;
  LAYER M1 ;
        RECT 2.464 0.924 2.496 3.864 ;
  LAYER M1 ;
        RECT 2.464 3.828 2.496 3.9 ;
  LAYER M2 ;
        RECT 2.444 3.848 2.516 3.88 ;
  LAYER M1 ;
        RECT 15.264 18.528 15.296 18.6 ;
  LAYER M2 ;
        RECT 15.244 18.548 15.316 18.58 ;
  LAYER M2 ;
        RECT 12.08 18.548 15.28 18.58 ;
  LAYER M1 ;
        RECT 12.064 18.528 12.096 18.6 ;
  LAYER M2 ;
        RECT 12.044 18.548 12.116 18.58 ;
  LAYER M1 ;
        RECT 15.264 15.588 15.296 15.66 ;
  LAYER M2 ;
        RECT 15.244 15.608 15.316 15.64 ;
  LAYER M2 ;
        RECT 12.08 15.608 15.28 15.64 ;
  LAYER M1 ;
        RECT 12.064 15.588 12.096 15.66 ;
  LAYER M2 ;
        RECT 12.044 15.608 12.116 15.64 ;
  LAYER M1 ;
        RECT 15.264 12.648 15.296 12.72 ;
  LAYER M2 ;
        RECT 15.244 12.668 15.316 12.7 ;
  LAYER M1 ;
        RECT 15.264 12.684 15.296 15.624 ;
  LAYER M1 ;
        RECT 15.264 15.588 15.296 15.66 ;
  LAYER M2 ;
        RECT 15.244 15.608 15.316 15.64 ;
  LAYER M1 ;
        RECT 15.264 9.708 15.296 9.78 ;
  LAYER M2 ;
        RECT 15.244 9.728 15.316 9.76 ;
  LAYER M1 ;
        RECT 15.264 9.744 15.296 12.684 ;
  LAYER M1 ;
        RECT 15.264 12.648 15.296 12.72 ;
  LAYER M2 ;
        RECT 15.244 12.668 15.316 12.7 ;
  LAYER M1 ;
        RECT 15.264 6.768 15.296 6.84 ;
  LAYER M2 ;
        RECT 15.244 6.788 15.316 6.82 ;
  LAYER M1 ;
        RECT 15.264 6.804 15.296 9.744 ;
  LAYER M1 ;
        RECT 15.264 9.708 15.296 9.78 ;
  LAYER M2 ;
        RECT 15.244 9.728 15.316 9.76 ;
  LAYER M1 ;
        RECT 15.264 3.828 15.296 3.9 ;
  LAYER M2 ;
        RECT 15.244 3.848 15.316 3.88 ;
  LAYER M1 ;
        RECT 15.264 3.864 15.296 6.804 ;
  LAYER M1 ;
        RECT 15.264 6.768 15.296 6.84 ;
  LAYER M2 ;
        RECT 15.244 6.788 15.316 6.82 ;
  LAYER M1 ;
        RECT 15.264 0.888 15.296 0.96 ;
  LAYER M2 ;
        RECT 15.244 0.908 15.316 0.94 ;
  LAYER M1 ;
        RECT 15.264 0.924 15.296 3.864 ;
  LAYER M1 ;
        RECT 15.264 3.828 15.296 3.9 ;
  LAYER M2 ;
        RECT 15.244 3.848 15.316 3.88 ;
  LAYER M1 ;
        RECT 3.264 12.144 3.296 12.216 ;
  LAYER M2 ;
        RECT 3.244 12.164 3.316 12.196 ;
  LAYER M2 ;
        RECT 2.8 12.164 3.28 12.196 ;
  LAYER M1 ;
        RECT 2.784 12.144 2.816 12.216 ;
  LAYER M2 ;
        RECT 2.764 12.164 2.836 12.196 ;
  LAYER M1 ;
        RECT 3.264 9.204 3.296 9.276 ;
  LAYER M2 ;
        RECT 3.244 9.224 3.316 9.256 ;
  LAYER M2 ;
        RECT 2.8 9.224 3.28 9.256 ;
  LAYER M1 ;
        RECT 2.784 9.204 2.816 9.276 ;
  LAYER M2 ;
        RECT 2.764 9.224 2.836 9.256 ;
  LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
  LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
  LAYER M1 ;
        RECT 2.784 21.336 2.816 21.504 ;
  LAYER M1 ;
        RECT 2.784 9.24 2.816 21.336 ;
  LAYER M1 ;
        RECT 9.664 12.144 9.696 12.216 ;
  LAYER M2 ;
        RECT 9.644 12.164 9.716 12.196 ;
  LAYER M1 ;
        RECT 9.664 12.18 9.696 12.348 ;
  LAYER M1 ;
        RECT 9.664 12.312 9.696 12.384 ;
  LAYER M2 ;
        RECT 9.644 12.332 9.716 12.364 ;
  LAYER M2 ;
        RECT 9.68 12.332 12.4 12.364 ;
  LAYER M1 ;
        RECT 12.384 12.312 12.416 12.384 ;
  LAYER M2 ;
        RECT 12.364 12.332 12.436 12.364 ;
  LAYER M1 ;
        RECT 9.664 15.084 9.696 15.156 ;
  LAYER M2 ;
        RECT 9.644 15.104 9.716 15.136 ;
  LAYER M1 ;
        RECT 9.664 15.12 9.696 15.288 ;
  LAYER M1 ;
        RECT 9.664 15.252 9.696 15.324 ;
  LAYER M2 ;
        RECT 9.644 15.272 9.716 15.304 ;
  LAYER M2 ;
        RECT 9.68 15.272 12.4 15.304 ;
  LAYER M1 ;
        RECT 12.384 15.252 12.416 15.324 ;
  LAYER M2 ;
        RECT 12.364 15.272 12.436 15.304 ;
  LAYER M1 ;
        RECT 12.384 21.468 12.416 21.54 ;
  LAYER M2 ;
        RECT 12.364 21.488 12.436 21.52 ;
  LAYER M1 ;
        RECT 12.384 21.336 12.416 21.504 ;
  LAYER M1 ;
        RECT 12.384 12.348 12.416 21.336 ;
  LAYER M2 ;
        RECT 2.8 21.488 12.4 21.52 ;
  LAYER M1 ;
        RECT 6.464 9.204 6.496 9.276 ;
  LAYER M2 ;
        RECT 6.444 9.224 6.516 9.256 ;
  LAYER M2 ;
        RECT 3.28 9.224 6.48 9.256 ;
  LAYER M1 ;
        RECT 3.264 9.204 3.296 9.276 ;
  LAYER M2 ;
        RECT 3.244 9.224 3.316 9.256 ;
  LAYER M1 ;
        RECT 6.464 15.084 6.496 15.156 ;
  LAYER M2 ;
        RECT 6.444 15.104 6.516 15.136 ;
  LAYER M2 ;
        RECT 6.48 15.104 9.68 15.136 ;
  LAYER M1 ;
        RECT 9.664 15.084 9.696 15.156 ;
  LAYER M2 ;
        RECT 9.644 15.104 9.716 15.136 ;
  LAYER M1 ;
        RECT 3.264 15.084 3.296 15.156 ;
  LAYER M2 ;
        RECT 3.244 15.104 3.316 15.136 ;
  LAYER M1 ;
        RECT 3.264 15.12 3.296 15.288 ;
  LAYER M1 ;
        RECT 3.264 15.252 3.296 15.324 ;
  LAYER M2 ;
        RECT 3.244 15.272 3.316 15.304 ;
  LAYER M2 ;
        RECT 3.28 15.272 6.16 15.304 ;
  LAYER M1 ;
        RECT 6.144 15.252 6.176 15.324 ;
  LAYER M2 ;
        RECT 6.124 15.272 6.196 15.304 ;
  LAYER M1 ;
        RECT 6.464 6.264 6.496 6.336 ;
  LAYER M2 ;
        RECT 6.444 6.284 6.516 6.316 ;
  LAYER M2 ;
        RECT 6.16 6.284 6.48 6.316 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M1 ;
        RECT 6.464 18.024 6.496 18.096 ;
  LAYER M2 ;
        RECT 6.444 18.044 6.516 18.076 ;
  LAYER M2 ;
        RECT 6.16 18.044 6.48 18.076 ;
  LAYER M1 ;
        RECT 6.144 18.024 6.176 18.096 ;
  LAYER M2 ;
        RECT 6.124 18.044 6.196 18.076 ;
  LAYER M1 ;
        RECT 3.264 18.024 3.296 18.096 ;
  LAYER M2 ;
        RECT 3.244 18.044 3.316 18.076 ;
  LAYER M1 ;
        RECT 3.264 18.06 3.296 18.228 ;
  LAYER M1 ;
        RECT 3.264 18.192 3.296 18.264 ;
  LAYER M2 ;
        RECT 3.244 18.212 3.316 18.244 ;
  LAYER M2 ;
        RECT 3.28 18.212 6.16 18.244 ;
  LAYER M1 ;
        RECT 6.144 18.192 6.176 18.264 ;
  LAYER M2 ;
        RECT 6.124 18.212 6.196 18.244 ;
  LAYER M1 ;
        RECT 6.144 21.636 6.176 21.708 ;
  LAYER M2 ;
        RECT 6.124 21.656 6.196 21.688 ;
  LAYER M1 ;
        RECT 6.144 21.336 6.176 21.672 ;
  LAYER M1 ;
        RECT 6.144 6.3 6.176 21.336 ;
  LAYER M1 ;
        RECT 9.664 9.204 9.696 9.276 ;
  LAYER M2 ;
        RECT 9.644 9.224 9.716 9.256 ;
  LAYER M2 ;
        RECT 9.36 9.224 9.68 9.256 ;
  LAYER M1 ;
        RECT 9.344 9.204 9.376 9.276 ;
  LAYER M2 ;
        RECT 9.324 9.224 9.396 9.256 ;
  LAYER M1 ;
        RECT 9.664 6.264 9.696 6.336 ;
  LAYER M2 ;
        RECT 9.644 6.284 9.716 6.316 ;
  LAYER M2 ;
        RECT 9.36 6.284 9.68 6.316 ;
  LAYER M1 ;
        RECT 9.344 6.264 9.376 6.336 ;
  LAYER M2 ;
        RECT 9.324 6.284 9.396 6.316 ;
  LAYER M1 ;
        RECT 9.344 21.636 9.376 21.708 ;
  LAYER M2 ;
        RECT 9.324 21.656 9.396 21.688 ;
  LAYER M1 ;
        RECT 9.344 21.336 9.376 21.672 ;
  LAYER M1 ;
        RECT 9.344 6.3 9.376 21.336 ;
  LAYER M2 ;
        RECT 6.16 21.656 9.36 21.688 ;
  LAYER M1 ;
        RECT 3.264 3.324 3.296 3.396 ;
  LAYER M2 ;
        RECT 3.244 3.344 3.316 3.376 ;
  LAYER M1 ;
        RECT 3.264 3.36 3.296 3.528 ;
  LAYER M1 ;
        RECT 3.264 3.492 3.296 3.564 ;
  LAYER M2 ;
        RECT 3.244 3.512 3.316 3.544 ;
  LAYER M2 ;
        RECT 3.28 3.512 6.32 3.544 ;
  LAYER M1 ;
        RECT 6.304 3.492 6.336 3.564 ;
  LAYER M2 ;
        RECT 6.284 3.512 6.356 3.544 ;
  LAYER M1 ;
        RECT 3.264 6.264 3.296 6.336 ;
  LAYER M2 ;
        RECT 3.244 6.284 3.316 6.316 ;
  LAYER M1 ;
        RECT 3.264 6.3 3.296 6.468 ;
  LAYER M1 ;
        RECT 3.264 6.432 3.296 6.504 ;
  LAYER M2 ;
        RECT 3.244 6.452 3.316 6.484 ;
  LAYER M2 ;
        RECT 3.28 6.452 6.32 6.484 ;
  LAYER M1 ;
        RECT 6.304 6.432 6.336 6.504 ;
  LAYER M2 ;
        RECT 6.284 6.452 6.356 6.484 ;
  LAYER M1 ;
        RECT 3.264 20.964 3.296 21.036 ;
  LAYER M2 ;
        RECT 3.244 20.984 3.316 21.016 ;
  LAYER M1 ;
        RECT 3.264 21 3.296 21.168 ;
  LAYER M1 ;
        RECT 3.264 21.132 3.296 21.204 ;
  LAYER M2 ;
        RECT 3.244 21.152 3.316 21.184 ;
  LAYER M2 ;
        RECT 3.28 21.152 6.32 21.184 ;
  LAYER M1 ;
        RECT 6.304 21.132 6.336 21.204 ;
  LAYER M2 ;
        RECT 6.284 21.152 6.356 21.184 ;
  LAYER M1 ;
        RECT 6.464 3.324 6.496 3.396 ;
  LAYER M2 ;
        RECT 6.444 3.344 6.516 3.376 ;
  LAYER M2 ;
        RECT 6.32 3.344 6.48 3.376 ;
  LAYER M1 ;
        RECT 6.304 3.324 6.336 3.396 ;
  LAYER M2 ;
        RECT 6.284 3.344 6.356 3.376 ;
  LAYER M1 ;
        RECT 6.464 12.144 6.496 12.216 ;
  LAYER M2 ;
        RECT 6.444 12.164 6.516 12.196 ;
  LAYER M2 ;
        RECT 6.32 12.164 6.48 12.196 ;
  LAYER M1 ;
        RECT 6.304 12.144 6.336 12.216 ;
  LAYER M2 ;
        RECT 6.284 12.164 6.356 12.196 ;
  LAYER M1 ;
        RECT 6.464 20.964 6.496 21.036 ;
  LAYER M2 ;
        RECT 6.444 20.984 6.516 21.016 ;
  LAYER M2 ;
        RECT 6.32 20.984 6.48 21.016 ;
  LAYER M1 ;
        RECT 6.304 20.964 6.336 21.036 ;
  LAYER M2 ;
        RECT 6.284 20.984 6.356 21.016 ;
  LAYER M1 ;
        RECT 6.304 21.804 6.336 21.876 ;
  LAYER M2 ;
        RECT 6.284 21.824 6.356 21.856 ;
  LAYER M1 ;
        RECT 6.304 21.336 6.336 21.84 ;
  LAYER M1 ;
        RECT 6.304 3.36 6.336 21.336 ;
  LAYER M1 ;
        RECT 9.664 3.324 9.696 3.396 ;
  LAYER M2 ;
        RECT 9.644 3.344 9.716 3.376 ;
  LAYER M2 ;
        RECT 9.52 3.344 9.68 3.376 ;
  LAYER M1 ;
        RECT 9.504 3.324 9.536 3.396 ;
  LAYER M2 ;
        RECT 9.484 3.344 9.556 3.376 ;
  LAYER M1 ;
        RECT 9.664 18.024 9.696 18.096 ;
  LAYER M2 ;
        RECT 9.644 18.044 9.716 18.076 ;
  LAYER M2 ;
        RECT 9.52 18.044 9.68 18.076 ;
  LAYER M1 ;
        RECT 9.504 18.024 9.536 18.096 ;
  LAYER M2 ;
        RECT 9.484 18.044 9.556 18.076 ;
  LAYER M1 ;
        RECT 9.664 20.964 9.696 21.036 ;
  LAYER M2 ;
        RECT 9.644 20.984 9.716 21.016 ;
  LAYER M2 ;
        RECT 9.52 20.984 9.68 21.016 ;
  LAYER M1 ;
        RECT 9.504 20.964 9.536 21.036 ;
  LAYER M2 ;
        RECT 9.484 20.984 9.556 21.016 ;
  LAYER M1 ;
        RECT 9.504 21.804 9.536 21.876 ;
  LAYER M2 ;
        RECT 9.484 21.824 9.556 21.856 ;
  LAYER M1 ;
        RECT 9.504 21.336 9.536 21.84 ;
  LAYER M1 ;
        RECT 9.504 3.36 9.536 21.336 ;
  LAYER M2 ;
        RECT 6.32 21.824 9.52 21.856 ;
  LAYER M1 ;
        RECT 0.064 20.964 0.096 21.036 ;
  LAYER M2 ;
        RECT 0.044 20.984 0.116 21.016 ;
  LAYER M2 ;
        RECT 0.08 20.984 3.28 21.016 ;
  LAYER M1 ;
        RECT 3.264 20.964 3.296 21.036 ;
  LAYER M2 ;
        RECT 3.244 20.984 3.316 21.016 ;
  LAYER M1 ;
        RECT 0.064 18.024 0.096 18.096 ;
  LAYER M2 ;
        RECT 0.044 18.044 0.116 18.076 ;
  LAYER M1 ;
        RECT 0.064 18.06 0.096 21 ;
  LAYER M1 ;
        RECT 0.064 20.964 0.096 21.036 ;
  LAYER M2 ;
        RECT 0.044 20.984 0.116 21.016 ;
  LAYER M1 ;
        RECT 0.064 15.084 0.096 15.156 ;
  LAYER M2 ;
        RECT 0.044 15.104 0.116 15.136 ;
  LAYER M1 ;
        RECT 0.064 15.12 0.096 18.06 ;
  LAYER M1 ;
        RECT 0.064 18.024 0.096 18.096 ;
  LAYER M2 ;
        RECT 0.044 18.044 0.116 18.076 ;
  LAYER M1 ;
        RECT 0.064 12.144 0.096 12.216 ;
  LAYER M2 ;
        RECT 0.044 12.164 0.116 12.196 ;
  LAYER M1 ;
        RECT 0.064 12.18 0.096 15.12 ;
  LAYER M1 ;
        RECT 0.064 15.084 0.096 15.156 ;
  LAYER M2 ;
        RECT 0.044 15.104 0.116 15.136 ;
  LAYER M1 ;
        RECT 0.064 9.204 0.096 9.276 ;
  LAYER M2 ;
        RECT 0.044 9.224 0.116 9.256 ;
  LAYER M1 ;
        RECT 0.064 9.24 0.096 12.18 ;
  LAYER M1 ;
        RECT 0.064 12.144 0.096 12.216 ;
  LAYER M2 ;
        RECT 0.044 12.164 0.116 12.196 ;
  LAYER M1 ;
        RECT 0.064 6.264 0.096 6.336 ;
  LAYER M2 ;
        RECT 0.044 6.284 0.116 6.316 ;
  LAYER M1 ;
        RECT 0.064 6.3 0.096 9.24 ;
  LAYER M1 ;
        RECT 0.064 9.204 0.096 9.276 ;
  LAYER M2 ;
        RECT 0.044 9.224 0.116 9.256 ;
  LAYER M1 ;
        RECT 0.064 3.324 0.096 3.396 ;
  LAYER M2 ;
        RECT 0.044 3.344 0.116 3.376 ;
  LAYER M1 ;
        RECT 0.064 3.36 0.096 6.3 ;
  LAYER M1 ;
        RECT 0.064 6.264 0.096 6.336 ;
  LAYER M2 ;
        RECT 0.044 6.284 0.116 6.316 ;
  LAYER M1 ;
        RECT 12.864 20.964 12.896 21.036 ;
  LAYER M2 ;
        RECT 12.844 20.984 12.916 21.016 ;
  LAYER M2 ;
        RECT 9.68 20.984 12.88 21.016 ;
  LAYER M1 ;
        RECT 9.664 20.964 9.696 21.036 ;
  LAYER M2 ;
        RECT 9.644 20.984 9.716 21.016 ;
  LAYER M1 ;
        RECT 12.864 18.024 12.896 18.096 ;
  LAYER M2 ;
        RECT 12.844 18.044 12.916 18.076 ;
  LAYER M2 ;
        RECT 9.68 18.044 12.88 18.076 ;
  LAYER M1 ;
        RECT 9.664 18.024 9.696 18.096 ;
  LAYER M2 ;
        RECT 9.644 18.044 9.716 18.076 ;
  LAYER M1 ;
        RECT 12.864 15.084 12.896 15.156 ;
  LAYER M2 ;
        RECT 12.844 15.104 12.916 15.136 ;
  LAYER M1 ;
        RECT 12.864 15.12 12.896 18.06 ;
  LAYER M1 ;
        RECT 12.864 18.024 12.896 18.096 ;
  LAYER M2 ;
        RECT 12.844 18.044 12.916 18.076 ;
  LAYER M1 ;
        RECT 12.864 12.144 12.896 12.216 ;
  LAYER M2 ;
        RECT 12.844 12.164 12.916 12.196 ;
  LAYER M1 ;
        RECT 12.864 12.18 12.896 15.12 ;
  LAYER M1 ;
        RECT 12.864 15.084 12.896 15.156 ;
  LAYER M2 ;
        RECT 12.844 15.104 12.916 15.136 ;
  LAYER M1 ;
        RECT 12.864 9.204 12.896 9.276 ;
  LAYER M2 ;
        RECT 12.844 9.224 12.916 9.256 ;
  LAYER M1 ;
        RECT 12.864 9.24 12.896 12.18 ;
  LAYER M1 ;
        RECT 12.864 12.144 12.896 12.216 ;
  LAYER M2 ;
        RECT 12.844 12.164 12.916 12.196 ;
  LAYER M1 ;
        RECT 12.864 6.264 12.896 6.336 ;
  LAYER M2 ;
        RECT 12.844 6.284 12.916 6.316 ;
  LAYER M1 ;
        RECT 12.864 6.3 12.896 9.24 ;
  LAYER M1 ;
        RECT 12.864 9.204 12.896 9.276 ;
  LAYER M2 ;
        RECT 12.844 9.224 12.916 9.256 ;
  LAYER M1 ;
        RECT 12.864 3.324 12.896 3.396 ;
  LAYER M2 ;
        RECT 12.844 3.344 12.916 3.376 ;
  LAYER M1 ;
        RECT 12.864 3.36 12.896 6.3 ;
  LAYER M1 ;
        RECT 12.864 6.264 12.896 6.336 ;
  LAYER M2 ;
        RECT 12.844 6.284 12.916 6.316 ;
  LAYER M1 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M2 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M3 ;
        RECT 0.08 0.924 2.48 3.36 ;
  LAYER M1 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M2 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M3 ;
        RECT 0.08 3.864 2.48 6.3 ;
  LAYER M1 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M2 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M3 ;
        RECT 0.08 6.804 2.48 9.24 ;
  LAYER M1 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M2 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M3 ;
        RECT 0.08 9.744 2.48 12.18 ;
  LAYER M1 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M2 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M3 ;
        RECT 0.08 12.684 2.48 15.12 ;
  LAYER M1 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M2 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M3 ;
        RECT 0.08 15.624 2.48 18.06 ;
  LAYER M1 ;
        RECT 0.08 18.564 2.48 21 ;
  LAYER M2 ;
        RECT 0.08 18.564 2.48 21 ;
  LAYER M3 ;
        RECT 0.08 18.564 2.48 21 ;
  LAYER M1 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M2 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M3 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M1 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M2 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M3 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M1 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M2 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M3 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M1 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M2 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M3 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M1 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M2 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M3 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M1 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M2 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M3 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M1 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M2 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M3 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M1 ;
        RECT 6.48 0.924 8.88 3.36 ;
  LAYER M2 ;
        RECT 6.48 0.924 8.88 3.36 ;
  LAYER M3 ;
        RECT 6.48 0.924 8.88 3.36 ;
  LAYER M1 ;
        RECT 6.48 3.864 8.88 6.3 ;
  LAYER M2 ;
        RECT 6.48 3.864 8.88 6.3 ;
  LAYER M3 ;
        RECT 6.48 3.864 8.88 6.3 ;
  LAYER M1 ;
        RECT 6.48 6.804 8.88 9.24 ;
  LAYER M2 ;
        RECT 6.48 6.804 8.88 9.24 ;
  LAYER M3 ;
        RECT 6.48 6.804 8.88 9.24 ;
  LAYER M1 ;
        RECT 6.48 9.744 8.88 12.18 ;
  LAYER M2 ;
        RECT 6.48 9.744 8.88 12.18 ;
  LAYER M3 ;
        RECT 6.48 9.744 8.88 12.18 ;
  LAYER M1 ;
        RECT 6.48 12.684 8.88 15.12 ;
  LAYER M2 ;
        RECT 6.48 12.684 8.88 15.12 ;
  LAYER M3 ;
        RECT 6.48 12.684 8.88 15.12 ;
  LAYER M1 ;
        RECT 6.48 15.624 8.88 18.06 ;
  LAYER M2 ;
        RECT 6.48 15.624 8.88 18.06 ;
  LAYER M3 ;
        RECT 6.48 15.624 8.88 18.06 ;
  LAYER M1 ;
        RECT 6.48 18.564 8.88 21 ;
  LAYER M2 ;
        RECT 6.48 18.564 8.88 21 ;
  LAYER M3 ;
        RECT 6.48 18.564 8.88 21 ;
  LAYER M1 ;
        RECT 9.68 0.924 12.08 3.36 ;
  LAYER M2 ;
        RECT 9.68 0.924 12.08 3.36 ;
  LAYER M3 ;
        RECT 9.68 0.924 12.08 3.36 ;
  LAYER M1 ;
        RECT 9.68 3.864 12.08 6.3 ;
  LAYER M2 ;
        RECT 9.68 3.864 12.08 6.3 ;
  LAYER M3 ;
        RECT 9.68 3.864 12.08 6.3 ;
  LAYER M1 ;
        RECT 9.68 6.804 12.08 9.24 ;
  LAYER M2 ;
        RECT 9.68 6.804 12.08 9.24 ;
  LAYER M3 ;
        RECT 9.68 6.804 12.08 9.24 ;
  LAYER M1 ;
        RECT 9.68 9.744 12.08 12.18 ;
  LAYER M2 ;
        RECT 9.68 9.744 12.08 12.18 ;
  LAYER M3 ;
        RECT 9.68 9.744 12.08 12.18 ;
  LAYER M1 ;
        RECT 9.68 12.684 12.08 15.12 ;
  LAYER M2 ;
        RECT 9.68 12.684 12.08 15.12 ;
  LAYER M3 ;
        RECT 9.68 12.684 12.08 15.12 ;
  LAYER M1 ;
        RECT 9.68 15.624 12.08 18.06 ;
  LAYER M2 ;
        RECT 9.68 15.624 12.08 18.06 ;
  LAYER M3 ;
        RECT 9.68 15.624 12.08 18.06 ;
  LAYER M1 ;
        RECT 9.68 18.564 12.08 21 ;
  LAYER M2 ;
        RECT 9.68 18.564 12.08 21 ;
  LAYER M3 ;
        RECT 9.68 18.564 12.08 21 ;
  LAYER M1 ;
        RECT 12.88 0.924 15.28 3.36 ;
  LAYER M2 ;
        RECT 12.88 0.924 15.28 3.36 ;
  LAYER M3 ;
        RECT 12.88 0.924 15.28 3.36 ;
  LAYER M1 ;
        RECT 12.88 3.864 15.28 6.3 ;
  LAYER M2 ;
        RECT 12.88 3.864 15.28 6.3 ;
  LAYER M3 ;
        RECT 12.88 3.864 15.28 6.3 ;
  LAYER M1 ;
        RECT 12.88 6.804 15.28 9.24 ;
  LAYER M2 ;
        RECT 12.88 6.804 15.28 9.24 ;
  LAYER M3 ;
        RECT 12.88 6.804 15.28 9.24 ;
  LAYER M1 ;
        RECT 12.88 9.744 15.28 12.18 ;
  LAYER M2 ;
        RECT 12.88 9.744 15.28 12.18 ;
  LAYER M3 ;
        RECT 12.88 9.744 15.28 12.18 ;
  LAYER M1 ;
        RECT 12.88 12.684 15.28 15.12 ;
  LAYER M2 ;
        RECT 12.88 12.684 15.28 15.12 ;
  LAYER M3 ;
        RECT 12.88 12.684 15.28 15.12 ;
  LAYER M1 ;
        RECT 12.88 15.624 15.28 18.06 ;
  LAYER M2 ;
        RECT 12.88 15.624 15.28 18.06 ;
  LAYER M3 ;
        RECT 12.88 15.624 15.28 18.06 ;
  LAYER M1 ;
        RECT 12.88 18.564 15.28 21 ;
  LAYER M2 ;
        RECT 12.88 18.564 15.28 21 ;
  LAYER M3 ;
        RECT 12.88 18.564 15.28 21 ;
  END 
END Cap_60fF_Cap_60fF
