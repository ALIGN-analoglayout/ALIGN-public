MACRO Cap_30fF_Cap_30fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_30fF 0 0 ;
  SIZE 12.24 BY 16.884 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 16.428 3.232 16.5 ;
      LAYER M2 ;
        RECT 3.18 16.448 3.252 16.48 ;
      LAYER M1 ;
        RECT 9.216 16.428 9.248 16.5 ;
      LAYER M2 ;
        RECT 9.196 16.448 9.268 16.48 ;
      LAYER M2 ;
        RECT 3.216 16.448 9.232 16.48 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
      LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 16.596 6.208 16.668 ;
      LAYER M2 ;
        RECT 6.156 16.616 6.228 16.648 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
      LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M2 ;
        RECT 6.032 7.208 8.784 7.24 ;
  LAYER M1 ;
        RECT 6.016 7.188 6.048 7.26 ;
  LAYER M2 ;
        RECT 5.996 7.208 6.068 7.24 ;
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.164 5.824 10.332 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M2 ;
        RECT 6.032 4.1 8.784 4.132 ;
  LAYER M1 ;
        RECT 6.016 4.08 6.048 4.152 ;
  LAYER M2 ;
        RECT 5.996 4.1 6.068 4.132 ;
  LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
  LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
  LAYER M1 ;
        RECT 6.016 0.42 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 10.164 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M2 ;
        RECT 3.056 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 3.04 7.188 3.072 7.26 ;
  LAYER M2 ;
        RECT 3.02 7.208 3.092 7.24 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M2 ;
        RECT 3.056 4.1 5.808 4.132 ;
  LAYER M1 ;
        RECT 3.04 4.08 3.072 4.152 ;
  LAYER M2 ;
        RECT 3.02 4.1 3.092 4.132 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 7.224 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M1 ;
        RECT 8.768 10.164 8.8 10.332 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M2 ;
        RECT 8.784 10.148 9.008 10.18 ;
  LAYER M1 ;
        RECT 8.992 10.128 9.024 10.2 ;
  LAYER M2 ;
        RECT 8.972 10.148 9.044 10.18 ;
  LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
  LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
  LAYER M1 ;
        RECT 8.992 0.252 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 10.164 ;
  LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 2.832 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 2.832 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 2.832 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 2.832 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 2.832 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 13.44 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.84 11.776 1.008 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M2 ;
        RECT 11.76 0.824 11.984 0.856 ;
  LAYER M1 ;
        RECT 11.968 0.804 12 0.876 ;
  LAYER M2 ;
        RECT 11.948 0.824 12.02 0.856 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M1 ;
        RECT 11.744 3.948 11.776 4.116 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 11.76 3.932 11.984 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M1 ;
        RECT 11.744 7.056 11.776 7.224 ;
  LAYER M1 ;
        RECT 11.744 7.02 11.776 7.092 ;
  LAYER M2 ;
        RECT 11.724 7.04 11.796 7.072 ;
  LAYER M2 ;
        RECT 11.76 7.04 11.984 7.072 ;
  LAYER M1 ;
        RECT 11.968 7.02 12 7.092 ;
  LAYER M2 ;
        RECT 11.948 7.04 12.02 7.072 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M1 ;
        RECT 11.744 10.164 11.776 10.332 ;
  LAYER M1 ;
        RECT 11.744 10.128 11.776 10.2 ;
  LAYER M2 ;
        RECT 11.724 10.148 11.796 10.18 ;
  LAYER M2 ;
        RECT 11.76 10.148 11.984 10.18 ;
  LAYER M1 ;
        RECT 11.968 10.128 12 10.2 ;
  LAYER M2 ;
        RECT 11.948 10.148 12.02 10.18 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 13.476 ;
  LAYER M2 ;
        RECT 11.724 13.424 11.796 13.456 ;
  LAYER M1 ;
        RECT 11.744 13.272 11.776 13.44 ;
  LAYER M1 ;
        RECT 11.744 13.236 11.776 13.308 ;
  LAYER M2 ;
        RECT 11.724 13.256 11.796 13.288 ;
  LAYER M2 ;
        RECT 11.76 13.256 11.984 13.288 ;
  LAYER M1 ;
        RECT 11.968 13.236 12 13.308 ;
  LAYER M2 ;
        RECT 11.948 13.256 12.02 13.288 ;
  LAYER M1 ;
        RECT 11.968 0.048 12 0.12 ;
  LAYER M2 ;
        RECT 11.948 0.068 12.02 0.1 ;
  LAYER M1 ;
        RECT 11.968 0.084 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 13.272 ;
  LAYER M2 ;
        RECT 0.08 0.068 11.984 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 2.832 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M2 ;
        RECT 2.832 13.424 5.808 13.456 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M2 ;
        RECT 5.808 13.424 8.784 13.456 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.2 16.428 3.232 16.5 ;
  LAYER M2 ;
        RECT 3.18 16.448 3.252 16.48 ;
  LAYER M1 ;
        RECT 3.2 16.212 3.232 16.464 ;
  LAYER M1 ;
        RECT 3.2 12.768 3.232 16.212 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M1 ;
        RECT 6.416 9.644 9.168 9.676 ;
  LAYER M1 ;
        RECT 9.152 9.624 9.184 9.696 ;
  LAYER M2 ;
        RECT 9.132 9.644 9.204 9.676 ;
  LAYER M2 ;
        RECT 9.168 9.644 9.232 9.676 ;
  LAYER M1 ;
        RECT 9.216 9.624 9.248 9.696 ;
  LAYER M2 ;
        RECT 9.196 9.644 9.268 9.676 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M1 ;
        RECT 6.416 6.536 9.168 6.568 ;
  LAYER M1 ;
        RECT 9.152 6.516 9.184 6.588 ;
  LAYER M2 ;
        RECT 9.132 6.536 9.204 6.568 ;
  LAYER M2 ;
        RECT 9.168 6.536 9.232 6.568 ;
  LAYER M1 ;
        RECT 9.216 6.516 9.248 6.588 ;
  LAYER M2 ;
        RECT 9.196 6.536 9.268 6.568 ;
  LAYER M1 ;
        RECT 9.216 16.428 9.248 16.5 ;
  LAYER M2 ;
        RECT 9.196 16.448 9.268 16.48 ;
  LAYER M1 ;
        RECT 9.216 16.212 9.248 16.464 ;
  LAYER M1 ;
        RECT 9.216 6.72 9.248 16.212 ;
  LAYER M2 ;
        RECT 3.216 16.448 9.232 16.48 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M1 ;
        RECT 3.44 9.644 6.192 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M2 ;
        RECT 6.192 9.644 6.256 9.676 ;
  LAYER M1 ;
        RECT 6.24 9.624 6.272 9.696 ;
  LAYER M2 ;
        RECT 6.22 9.644 6.292 9.676 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M1 ;
        RECT 3.44 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.256 6.568 ;
  LAYER M1 ;
        RECT 6.24 6.516 6.272 6.588 ;
  LAYER M2 ;
        RECT 6.22 6.536 6.292 6.568 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 6.192 12.752 6.416 12.784 ;
  LAYER M1 ;
        RECT 6.176 12.732 6.208 12.804 ;
  LAYER M2 ;
        RECT 6.156 12.752 6.228 12.784 ;
  LAYER M1 ;
        RECT 6.176 16.596 6.208 16.668 ;
  LAYER M2 ;
        RECT 6.156 16.616 6.228 16.648 ;
  LAYER M1 ;
        RECT 6.176 16.212 6.208 16.632 ;
  LAYER M1 ;
        RECT 6.176 6.72 6.208 16.212 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.464 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.224 16.764 0.256 16.836 ;
  LAYER M2 ;
        RECT 0.204 16.784 0.276 16.816 ;
  LAYER M1 ;
        RECT 0.224 16.212 0.256 16.8 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 16.212 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 9.392 3.428 12.144 3.46 ;
  LAYER M1 ;
        RECT 12.128 3.408 12.16 3.48 ;
  LAYER M2 ;
        RECT 12.108 3.428 12.18 3.46 ;
  LAYER M2 ;
        RECT 12.144 3.428 12.208 3.46 ;
  LAYER M1 ;
        RECT 12.192 3.408 12.224 3.48 ;
  LAYER M2 ;
        RECT 12.172 3.428 12.244 3.46 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.392 6.536 12.144 6.568 ;
  LAYER M1 ;
        RECT 12.128 6.516 12.16 6.588 ;
  LAYER M2 ;
        RECT 12.108 6.536 12.18 6.568 ;
  LAYER M2 ;
        RECT 12.144 6.536 12.208 6.568 ;
  LAYER M1 ;
        RECT 12.192 6.516 12.224 6.588 ;
  LAYER M2 ;
        RECT 12.172 6.536 12.244 6.568 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M1 ;
        RECT 9.392 9.644 12.144 9.676 ;
  LAYER M1 ;
        RECT 12.128 9.624 12.16 9.696 ;
  LAYER M2 ;
        RECT 12.108 9.644 12.18 9.676 ;
  LAYER M2 ;
        RECT 12.144 9.644 12.208 9.676 ;
  LAYER M1 ;
        RECT 12.192 9.624 12.224 9.696 ;
  LAYER M2 ;
        RECT 12.172 9.644 12.244 9.676 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M1 ;
        RECT 9.392 12.752 12.144 12.784 ;
  LAYER M1 ;
        RECT 12.128 12.732 12.16 12.804 ;
  LAYER M2 ;
        RECT 12.108 12.752 12.18 12.784 ;
  LAYER M2 ;
        RECT 12.144 12.752 12.208 12.784 ;
  LAYER M1 ;
        RECT 12.192 12.732 12.224 12.804 ;
  LAYER M2 ;
        RECT 12.172 12.752 12.244 12.784 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M1 ;
        RECT 9.392 15.86 12.144 15.892 ;
  LAYER M1 ;
        RECT 12.128 15.84 12.16 15.912 ;
  LAYER M2 ;
        RECT 12.108 15.86 12.18 15.892 ;
  LAYER M2 ;
        RECT 12.144 15.86 12.208 15.892 ;
  LAYER M1 ;
        RECT 12.192 15.84 12.224 15.912 ;
  LAYER M2 ;
        RECT 12.172 15.86 12.244 15.892 ;
  LAYER M1 ;
        RECT 12.192 16.764 12.224 16.836 ;
  LAYER M2 ;
        RECT 12.172 16.784 12.244 16.816 ;
  LAYER M1 ;
        RECT 12.192 16.212 12.224 16.8 ;
  LAYER M1 ;
        RECT 12.192 3.612 12.224 16.212 ;
  LAYER M2 ;
        RECT 0.24 16.784 12.208 16.816 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 0.464 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M2 ;
        RECT 3.44 15.86 6.416 15.892 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M3 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M3 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M3 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M3 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M2 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M1 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M3 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M3 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M3 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M3 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M3 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M2 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M1 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M3 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M3 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M3 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M3 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M3 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M2 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M1 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M3 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M3 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M3 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M3 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M3 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M2 ;
        RECT 9.328 13.356 11.824 15.96 ;
  END 
END Cap_30fF_Cap_30fF
