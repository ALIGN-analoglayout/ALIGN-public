MACRO test
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 2.5600 BY 1.6800 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
      LAYER M2 ;
        RECT 0.2040 0.9080 2.3560 0.9400 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
      LAYER M2 ;
        RECT 1.0040 0.9920 1.5560 1.0240 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 1.5560 0.2680 ;
      LAYER M2 ;
        RECT 0.3640 1.0760 2.1960 1.1080 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 2.2760 0.3520 ;
      LAYER M2 ;
        RECT 0.9240 1.1600 1.6360 1.1920 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4040 1.6360 0.4360 ;
      LAYER M2 ;
        RECT 0.2840 1.2440 2.2760 1.2760 ;
    END
  END GB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER V0 ;
      RECT 0.2240 0.2360 0.2560 0.2680 ;
    LAYER V0 ;
      RECT 0.2240 0.3620 0.2560 0.3940 ;
    LAYER V0 ;
      RECT 0.2240 0.4880 0.2560 0.5200 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER V0 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V0 ;
      RECT 2.3040 0.3620 2.3360 0.3940 ;
    LAYER V0 ;
      RECT 2.3040 0.4880 2.3360 0.5200 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER V0 ;
      RECT 0.8640 0.2360 0.8960 0.2680 ;
    LAYER V0 ;
      RECT 0.8640 0.3620 0.8960 0.3940 ;
    LAYER V0 ;
      RECT 0.8640 0.4880 0.8960 0.5200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER V0 ;
      RECT 1.6640 0.2360 1.6960 0.2680 ;
    LAYER V0 ;
      RECT 1.6640 0.3620 1.6960 0.3940 ;
    LAYER V0 ;
      RECT 1.6640 0.4880 1.6960 0.5200 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER V0 ;
      RECT 0.3840 0.2360 0.4160 0.2680 ;
    LAYER V0 ;
      RECT 0.3840 0.3620 0.4160 0.3940 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 0.4160 0.5200 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER V0 ;
      RECT 2.1440 0.2360 2.1760 0.2680 ;
    LAYER V0 ;
      RECT 2.1440 0.3620 2.1760 0.3940 ;
    LAYER V0 ;
      RECT 2.1440 0.4880 2.1760 0.5200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER V0 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V0 ;
      RECT 1.0240 0.3620 1.0560 0.3940 ;
    LAYER V0 ;
      RECT 1.0240 0.4880 1.0560 0.5200 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER V0 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER V0 ;
      RECT 1.5040 0.3620 1.5360 0.3940 ;
    LAYER V0 ;
      RECT 1.5040 0.4880 1.5360 0.5200 ;
    LAYER M3 ;
      RECT 1.2600 0.0480 1.3000 0.1200 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 2.3040 0.0680 2.3360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.6640 0.0680 1.6960 0.1000 ;
    LAYER M3 ;
      RECT 1.1800 0.1320 1.2200 0.2040 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 2.1440 0.1520 2.1760 0.1840 ;
    LAYER M3 ;
      RECT 1.3400 0.2160 1.3800 0.2880 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.5040 0.2360 1.5360 0.2680 ;
    LAYER M3 ;
      RECT 1.1000 0.3000 1.1400 0.3720 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V1 ;
      RECT 0.3040 0.3200 0.3360 0.3520 ;
    LAYER V1 ;
      RECT 2.2240 0.3200 2.2560 0.3520 ;
    LAYER M3 ;
      RECT 1.4200 0.3840 1.4600 0.4560 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V1 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V1 ;
      RECT 1.5840 0.4040 1.6160 0.4360 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER V0 ;
      RECT 0.2240 1.0760 0.2560 1.1080 ;
    LAYER V0 ;
      RECT 0.2240 1.2020 0.2560 1.2340 ;
    LAYER V0 ;
      RECT 0.2240 1.3280 0.2560 1.3600 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER V0 ;
      RECT 2.3040 1.0760 2.3360 1.1080 ;
    LAYER V0 ;
      RECT 2.3040 1.2020 2.3360 1.2340 ;
    LAYER V0 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER V0 ;
      RECT 0.8640 1.0760 0.8960 1.1080 ;
    LAYER V0 ;
      RECT 0.8640 1.2020 0.8960 1.2340 ;
    LAYER V0 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER V0 ;
      RECT 1.6640 1.0760 1.6960 1.1080 ;
    LAYER V0 ;
      RECT 1.6640 1.2020 1.6960 1.2340 ;
    LAYER V0 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER V0 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V0 ;
      RECT 0.3840 1.2020 0.4160 1.2340 ;
    LAYER V0 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER V0 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER V0 ;
      RECT 2.1440 1.2020 2.1760 1.2340 ;
    LAYER V0 ;
      RECT 2.1440 1.3280 2.1760 1.3600 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER V0 ;
      RECT 1.0240 1.0760 1.0560 1.1080 ;
    LAYER V0 ;
      RECT 1.0240 1.2020 1.0560 1.2340 ;
    LAYER V0 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER V0 ;
      RECT 1.5040 1.0760 1.5360 1.1080 ;
    LAYER V0 ;
      RECT 1.5040 1.2020 1.5360 1.2340 ;
    LAYER V0 ;
      RECT 1.5040 1.3280 1.5360 1.3600 ;
    LAYER M3 ;
      RECT 1.2600 0.0480 1.3000 0.9600 ;
    LAYER V2 ;
      RECT 1.2600 0.0680 1.3000 0.1000 ;
    LAYER V2 ;
      RECT 1.2600 0.9080 1.3000 0.9400 ;
    LAYER V1 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V1 ;
      RECT 2.3040 0.9080 2.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.8640 0.9080 0.8960 0.9400 ;
    LAYER V1 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER M3 ;
      RECT 1.1800 0.1320 1.2200 1.0440 ;
    LAYER V2 ;
      RECT 1.1800 0.1520 1.2200 0.1840 ;
    LAYER V2 ;
      RECT 1.1800 0.9920 1.2200 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.5040 0.9920 1.5360 1.0240 ;
    LAYER M3 ;
      RECT 1.3400 0.2160 1.3800 1.1280 ;
    LAYER V2 ;
      RECT 1.3400 0.2360 1.3800 0.2680 ;
    LAYER V2 ;
      RECT 1.3400 1.0760 1.3800 1.1080 ;
    LAYER V1 ;
      RECT 0.3840 1.0760 0.4160 1.1080 ;
    LAYER V1 ;
      RECT 2.1440 1.0760 2.1760 1.1080 ;
    LAYER M3 ;
      RECT 1.1000 0.3000 1.1400 1.2120 ;
    LAYER V2 ;
      RECT 1.1000 0.3200 1.1400 0.3520 ;
    LAYER V2 ;
      RECT 1.1000 1.1600 1.1400 1.1920 ;
    LAYER V1 ;
      RECT 0.9440 1.1600 0.9760 1.1920 ;
    LAYER V1 ;
      RECT 1.5840 1.1600 1.6160 1.1920 ;
    LAYER M3 ;
      RECT 1.4200 0.3840 1.4600 1.2960 ;
    LAYER V2 ;
      RECT 1.4200 0.4040 1.4600 0.4360 ;
    LAYER V2 ;
      RECT 1.4200 1.2440 1.4600 1.2760 ;
    LAYER V1 ;
      RECT 0.3040 1.2440 0.3360 1.2760 ;
    LAYER V1 ;
      RECT 2.2240 1.2440 2.2560 1.2760 ;
  END
END test
