MACRO DCL_PMOS_nfin60_n12_X5_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_nfin60_n12_X5_Y1_RVT 0 0 ;
  SIZE 1.2800 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 0.9600 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.0760 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 1.4960 0.9960 1.5280 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.9960 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.9960 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V2 ;
      RECT 0.4640 0.0680 0.4960 0.1000 ;
    LAYER V2 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.5440 0.1520 0.5760 0.1840 ;
    LAYER V2 ;
      RECT 0.5440 0.9080 0.5760 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
  END
END DCL_PMOS_nfin60_n12_X5_Y1_RVT
MACRO SCM_NMOS_nfin10_n12_X1_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin10_n12_X1_Y1_RVT 0 0 ;
  SIZE 0.8000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.2360 0.5160 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.5960 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.5160 1.5280 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 0.5160 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 0.1520 0.3560 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V2 ;
      RECT 0.2240 0.1520 0.2560 0.1840 ;
    LAYER V2 ;
      RECT 0.2240 0.9080 0.2560 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
  END
END SCM_NMOS_nfin10_n12_X1_Y1_RVT
MACRO SCM_NMOS_nfin24_n12_X2_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin24_n12_X2_Y1_RVT 0 0 ;
  SIZE 1.1200 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.0480 0.3400 1.5480 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.1320 0.4200 0.9600 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 0.6760 0.2680 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2840 1.4960 0.8360 1.5280 ;
    LAYER M2 ;
      RECT 0.2840 0.9080 0.8360 0.9400 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 0.8360 0.1840 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.2360 0.6560 0.2680 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.1520 0.8160 0.1840 ;
    LAYER V1 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V2 ;
      RECT 0.3040 0.0680 0.3360 0.1000 ;
    LAYER V2 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V2 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V2 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
  END
END SCM_NMOS_nfin24_n12_X2_Y1_RVT
MACRO Switch_PMOS_nfin240_n12_X5_Y4_ST2_RVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin240_n12_X5_Y4_ST2_RVT 0 0 ;
  SIZE 2.0800 BY 5.3760 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.0480 0.8200 5.0760 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8600 0.1320 0.9000 3.7320 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9400 0.8880 0.9800 4.4880 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.4000 0.4160 3.1440 ;
    LAYER M1 ;
      RECT 0.3840 3.2400 0.4160 3.4800 ;
    LAYER M1 ;
      RECT 0.3840 3.5760 0.4160 4.3200 ;
    LAYER M1 ;
      RECT 0.3840 4.4160 0.4160 4.6560 ;
    LAYER M1 ;
      RECT 0.3840 4.9200 0.4160 5.1600 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.2240 2.4000 0.2560 3.1440 ;
    LAYER M1 ;
      RECT 0.2240 3.5760 0.2560 4.3200 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 2.4000 0.5760 3.1440 ;
    LAYER M1 ;
      RECT 0.5440 3.5760 0.5760 4.3200 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.4000 0.7360 3.1440 ;
    LAYER M1 ;
      RECT 0.7040 3.2400 0.7360 3.4800 ;
    LAYER M1 ;
      RECT 0.7040 3.5760 0.7360 4.3200 ;
    LAYER M1 ;
      RECT 0.7040 4.4160 0.7360 4.6560 ;
    LAYER M1 ;
      RECT 0.7040 4.9200 0.7360 5.1600 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 0.8640 2.4000 0.8960 3.1440 ;
    LAYER M1 ;
      RECT 0.8640 3.5760 0.8960 4.3200 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.1280 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.0640 1.0560 2.3040 ;
    LAYER M1 ;
      RECT 1.0240 2.4000 1.0560 3.1440 ;
    LAYER M1 ;
      RECT 1.0240 3.2400 1.0560 3.4800 ;
    LAYER M1 ;
      RECT 1.0240 3.5760 1.0560 4.3200 ;
    LAYER M1 ;
      RECT 1.0240 4.4160 1.0560 4.6560 ;
    LAYER M1 ;
      RECT 1.0240 4.9200 1.0560 5.1600 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.1840 2.4000 1.2160 3.1440 ;
    LAYER M1 ;
      RECT 1.1840 3.5760 1.2160 4.3200 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.8880 1.3760 1.1280 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 2.0640 1.3760 2.3040 ;
    LAYER M1 ;
      RECT 1.3440 2.4000 1.3760 3.1440 ;
    LAYER M1 ;
      RECT 1.3440 3.2400 1.3760 3.4800 ;
    LAYER M1 ;
      RECT 1.3440 3.5760 1.3760 4.3200 ;
    LAYER M1 ;
      RECT 1.3440 4.4160 1.3760 4.6560 ;
    LAYER M1 ;
      RECT 1.3440 4.9200 1.3760 5.1600 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M1 ;
      RECT 1.5040 2.4000 1.5360 3.1440 ;
    LAYER M1 ;
      RECT 1.5040 3.5760 1.5360 4.3200 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.1280 ;
    LAYER M1 ;
      RECT 1.6640 1.2240 1.6960 1.9680 ;
    LAYER M1 ;
      RECT 1.6640 2.0640 1.6960 2.3040 ;
    LAYER M1 ;
      RECT 1.6640 2.4000 1.6960 3.1440 ;
    LAYER M1 ;
      RECT 1.6640 3.2400 1.6960 3.4800 ;
    LAYER M1 ;
      RECT 1.6640 3.5760 1.6960 4.3200 ;
    LAYER M1 ;
      RECT 1.6640 4.4160 1.6960 4.6560 ;
    LAYER M1 ;
      RECT 1.6640 4.9200 1.6960 5.1600 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.8240 1.2240 1.8560 1.9680 ;
    LAYER M1 ;
      RECT 1.8240 2.4000 1.8560 3.1440 ;
    LAYER M1 ;
      RECT 1.8240 3.5760 1.8560 4.3200 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.8760 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 1.7160 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.8760 1.2760 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 1.7160 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 1.7160 2.1160 ;
    LAYER M2 ;
      RECT 0.2040 2.4200 1.8760 2.4520 ;
    LAYER M2 ;
      RECT 0.3640 2.5040 1.7160 2.5360 ;
    LAYER M2 ;
      RECT 0.3640 3.2600 1.7160 3.2920 ;
    LAYER M2 ;
      RECT 0.2040 3.5960 1.8760 3.6280 ;
    LAYER M2 ;
      RECT 0.3640 5.0240 1.7160 5.0560 ;
    LAYER M2 ;
      RECT 0.3640 3.6800 1.7160 3.7120 ;
    LAYER M2 ;
      RECT 0.3640 4.4360 1.7160 4.4680 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 2.4200 0.2560 2.4520 ;
    LAYER V1 ;
      RECT 0.2240 3.5960 0.2560 3.6280 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 2.4200 0.5760 2.4520 ;
    LAYER V1 ;
      RECT 0.5440 3.5960 0.5760 3.6280 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 2.4200 0.8960 2.4520 ;
    LAYER V1 ;
      RECT 0.8640 3.5960 0.8960 3.6280 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 2.4200 1.2160 2.4520 ;
    LAYER V1 ;
      RECT 1.1840 3.5960 1.2160 3.6280 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 2.4200 1.5360 2.4520 ;
    LAYER V1 ;
      RECT 1.5040 3.5960 1.5360 3.6280 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 1.2440 1.8560 1.2760 ;
    LAYER V1 ;
      RECT 1.8240 2.4200 1.8560 2.4520 ;
    LAYER V1 ;
      RECT 1.8240 3.5960 1.8560 3.6280 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.5040 0.4160 2.5360 ;
    LAYER V1 ;
      RECT 0.3840 3.2600 0.4160 3.2920 ;
    LAYER V1 ;
      RECT 0.3840 3.6800 0.4160 3.7120 ;
    LAYER V1 ;
      RECT 0.3840 4.4360 0.4160 4.4680 ;
    LAYER V1 ;
      RECT 0.3840 5.0240 0.4160 5.0560 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.5040 0.7360 2.5360 ;
    LAYER V1 ;
      RECT 0.7040 3.2600 0.7360 3.2920 ;
    LAYER V1 ;
      RECT 0.7040 3.6800 0.7360 3.7120 ;
    LAYER V1 ;
      RECT 0.7040 4.4360 0.7360 4.4680 ;
    LAYER V1 ;
      RECT 0.7040 5.0240 0.7360 5.0560 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V1 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER V1 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V1 ;
      RECT 1.0240 2.5040 1.0560 2.5360 ;
    LAYER V1 ;
      RECT 1.0240 3.2600 1.0560 3.2920 ;
    LAYER V1 ;
      RECT 1.0240 3.6800 1.0560 3.7120 ;
    LAYER V1 ;
      RECT 1.0240 4.4360 1.0560 4.4680 ;
    LAYER V1 ;
      RECT 1.0240 5.0240 1.0560 5.0560 ;
    LAYER V1 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V1 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V1 ;
      RECT 1.3440 1.3280 1.3760 1.3600 ;
    LAYER V1 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V1 ;
      RECT 1.3440 2.5040 1.3760 2.5360 ;
    LAYER V1 ;
      RECT 1.3440 3.2600 1.3760 3.2920 ;
    LAYER V1 ;
      RECT 1.3440 3.6800 1.3760 3.7120 ;
    LAYER V1 ;
      RECT 1.3440 4.4360 1.3760 4.4680 ;
    LAYER V1 ;
      RECT 1.3440 5.0240 1.3760 5.0560 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V1 ;
      RECT 1.6640 1.3280 1.6960 1.3600 ;
    LAYER V1 ;
      RECT 1.6640 2.0840 1.6960 2.1160 ;
    LAYER V1 ;
      RECT 1.6640 2.5040 1.6960 2.5360 ;
    LAYER V1 ;
      RECT 1.6640 3.2600 1.6960 3.2920 ;
    LAYER V1 ;
      RECT 1.6640 3.6800 1.6960 3.7120 ;
    LAYER V1 ;
      RECT 1.6640 4.4360 1.6960 4.4680 ;
    LAYER V1 ;
      RECT 1.6640 5.0240 1.6960 5.0560 ;
    LAYER V2 ;
      RECT 0.7840 0.0680 0.8160 0.1000 ;
    LAYER V2 ;
      RECT 0.7840 1.2440 0.8160 1.2760 ;
    LAYER V2 ;
      RECT 0.7840 2.4200 0.8160 2.4520 ;
    LAYER V2 ;
      RECT 0.7840 3.5960 0.8160 3.6280 ;
    LAYER V2 ;
      RECT 0.7840 5.0240 0.8160 5.0560 ;
    LAYER V2 ;
      RECT 0.8640 0.1520 0.8960 0.1840 ;
    LAYER V2 ;
      RECT 0.8640 1.3280 0.8960 1.3600 ;
    LAYER V2 ;
      RECT 0.8640 2.5040 0.8960 2.5360 ;
    LAYER V2 ;
      RECT 0.8640 3.6800 0.8960 3.7120 ;
    LAYER V2 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V2 ;
      RECT 0.9440 2.0840 0.9760 2.1160 ;
    LAYER V2 ;
      RECT 0.9440 3.2600 0.9760 3.2920 ;
    LAYER V2 ;
      RECT 0.9440 4.4360 0.9760 4.4680 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.7560 0.4160 2.7880 ;
    LAYER V0 ;
      RECT 0.3840 2.8820 0.4160 2.9140 ;
    LAYER V0 ;
      RECT 0.3840 3.0080 0.4160 3.0400 ;
    LAYER V0 ;
      RECT 0.3840 3.2600 0.4160 3.2920 ;
    LAYER V0 ;
      RECT 0.3840 3.9320 0.4160 3.9640 ;
    LAYER V0 ;
      RECT 0.3840 4.0580 0.4160 4.0900 ;
    LAYER V0 ;
      RECT 0.3840 4.1840 0.4160 4.2160 ;
    LAYER V0 ;
      RECT 0.3840 4.4360 0.4160 4.4680 ;
    LAYER V0 ;
      RECT 0.3840 5.0240 0.4160 5.0560 ;
    LAYER V0 ;
      RECT 0.3840 5.0240 0.4160 5.0560 ;
    LAYER V0 ;
      RECT 0.3840 5.0240 0.4160 5.0560 ;
    LAYER V0 ;
      RECT 0.3840 5.0240 0.4160 5.0560 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.2240 2.7560 0.2560 2.7880 ;
    LAYER V0 ;
      RECT 0.2240 2.8820 0.2560 2.9140 ;
    LAYER V0 ;
      RECT 0.2240 3.0080 0.2560 3.0400 ;
    LAYER V0 ;
      RECT 0.2240 3.9320 0.2560 3.9640 ;
    LAYER V0 ;
      RECT 0.2240 4.0580 0.2560 4.0900 ;
    LAYER V0 ;
      RECT 0.2240 4.1840 0.2560 4.2160 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.7560 0.5760 2.7880 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 2.8820 0.5760 2.9140 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.0080 0.5760 3.0400 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 3.9320 0.5760 3.9640 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.0580 0.5760 4.0900 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.5440 4.1840 0.5760 4.2160 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.7560 0.7360 2.7880 ;
    LAYER V0 ;
      RECT 0.7040 2.8820 0.7360 2.9140 ;
    LAYER V0 ;
      RECT 0.7040 3.0080 0.7360 3.0400 ;
    LAYER V0 ;
      RECT 0.7040 3.2600 0.7360 3.2920 ;
    LAYER V0 ;
      RECT 0.7040 3.9320 0.7360 3.9640 ;
    LAYER V0 ;
      RECT 0.7040 4.0580 0.7360 4.0900 ;
    LAYER V0 ;
      RECT 0.7040 4.1840 0.7360 4.2160 ;
    LAYER V0 ;
      RECT 0.7040 4.4360 0.7360 4.4680 ;
    LAYER V0 ;
      RECT 0.7040 5.0240 0.7360 5.0560 ;
    LAYER V0 ;
      RECT 0.7040 5.0240 0.7360 5.0560 ;
    LAYER V0 ;
      RECT 0.7040 5.0240 0.7360 5.0560 ;
    LAYER V0 ;
      RECT 0.7040 5.0240 0.7360 5.0560 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.7560 0.8960 2.7880 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 2.8820 0.8960 2.9140 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.0080 0.8960 3.0400 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 3.9320 0.8960 3.9640 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.0580 0.8960 4.0900 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 0.8640 4.1840 0.8960 4.2160 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V0 ;
      RECT 1.0240 2.7560 1.0560 2.7880 ;
    LAYER V0 ;
      RECT 1.0240 2.8820 1.0560 2.9140 ;
    LAYER V0 ;
      RECT 1.0240 3.0080 1.0560 3.0400 ;
    LAYER V0 ;
      RECT 1.0240 3.2600 1.0560 3.2920 ;
    LAYER V0 ;
      RECT 1.0240 3.9320 1.0560 3.9640 ;
    LAYER V0 ;
      RECT 1.0240 4.0580 1.0560 4.0900 ;
    LAYER V0 ;
      RECT 1.0240 4.1840 1.0560 4.2160 ;
    LAYER V0 ;
      RECT 1.0240 4.4360 1.0560 4.4680 ;
    LAYER V0 ;
      RECT 1.0240 5.0240 1.0560 5.0560 ;
    LAYER V0 ;
      RECT 1.0240 5.0240 1.0560 5.0560 ;
    LAYER V0 ;
      RECT 1.0240 5.0240 1.0560 5.0560 ;
    LAYER V0 ;
      RECT 1.0240 5.0240 1.0560 5.0560 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 2.7560 1.2160 2.7880 ;
    LAYER V0 ;
      RECT 1.1840 2.7560 1.2160 2.7880 ;
    LAYER V0 ;
      RECT 1.1840 2.8820 1.2160 2.9140 ;
    LAYER V0 ;
      RECT 1.1840 2.8820 1.2160 2.9140 ;
    LAYER V0 ;
      RECT 1.1840 3.0080 1.2160 3.0400 ;
    LAYER V0 ;
      RECT 1.1840 3.0080 1.2160 3.0400 ;
    LAYER V0 ;
      RECT 1.1840 3.9320 1.2160 3.9640 ;
    LAYER V0 ;
      RECT 1.1840 3.9320 1.2160 3.9640 ;
    LAYER V0 ;
      RECT 1.1840 4.0580 1.2160 4.0900 ;
    LAYER V0 ;
      RECT 1.1840 4.0580 1.2160 4.0900 ;
    LAYER V0 ;
      RECT 1.1840 4.1840 1.2160 4.2160 ;
    LAYER V0 ;
      RECT 1.1840 4.1840 1.2160 4.2160 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V0 ;
      RECT 1.3440 2.7560 1.3760 2.7880 ;
    LAYER V0 ;
      RECT 1.3440 2.8820 1.3760 2.9140 ;
    LAYER V0 ;
      RECT 1.3440 3.0080 1.3760 3.0400 ;
    LAYER V0 ;
      RECT 1.3440 3.2600 1.3760 3.2920 ;
    LAYER V0 ;
      RECT 1.3440 3.9320 1.3760 3.9640 ;
    LAYER V0 ;
      RECT 1.3440 4.0580 1.3760 4.0900 ;
    LAYER V0 ;
      RECT 1.3440 4.1840 1.3760 4.2160 ;
    LAYER V0 ;
      RECT 1.3440 4.4360 1.3760 4.4680 ;
    LAYER V0 ;
      RECT 1.3440 5.0240 1.3760 5.0560 ;
    LAYER V0 ;
      RECT 1.3440 5.0240 1.3760 5.0560 ;
    LAYER V0 ;
      RECT 1.3440 5.0240 1.3760 5.0560 ;
    LAYER V0 ;
      RECT 1.3440 5.0240 1.3760 5.0560 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5040 2.7560 1.5360 2.7880 ;
    LAYER V0 ;
      RECT 1.5040 2.7560 1.5360 2.7880 ;
    LAYER V0 ;
      RECT 1.5040 2.8820 1.5360 2.9140 ;
    LAYER V0 ;
      RECT 1.5040 2.8820 1.5360 2.9140 ;
    LAYER V0 ;
      RECT 1.5040 3.0080 1.5360 3.0400 ;
    LAYER V0 ;
      RECT 1.5040 3.0080 1.5360 3.0400 ;
    LAYER V0 ;
      RECT 1.5040 3.9320 1.5360 3.9640 ;
    LAYER V0 ;
      RECT 1.5040 3.9320 1.5360 3.9640 ;
    LAYER V0 ;
      RECT 1.5040 4.0580 1.5360 4.0900 ;
    LAYER V0 ;
      RECT 1.5040 4.0580 1.5360 4.0900 ;
    LAYER V0 ;
      RECT 1.5040 4.1840 1.5360 4.2160 ;
    LAYER V0 ;
      RECT 1.5040 4.1840 1.5360 4.2160 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.6640 2.0840 1.6960 2.1160 ;
    LAYER V0 ;
      RECT 1.6640 2.7560 1.6960 2.7880 ;
    LAYER V0 ;
      RECT 1.6640 2.8820 1.6960 2.9140 ;
    LAYER V0 ;
      RECT 1.6640 3.0080 1.6960 3.0400 ;
    LAYER V0 ;
      RECT 1.6640 3.2600 1.6960 3.2920 ;
    LAYER V0 ;
      RECT 1.6640 3.9320 1.6960 3.9640 ;
    LAYER V0 ;
      RECT 1.6640 4.0580 1.6960 4.0900 ;
    LAYER V0 ;
      RECT 1.6640 4.1840 1.6960 4.2160 ;
    LAYER V0 ;
      RECT 1.6640 4.4360 1.6960 4.4680 ;
    LAYER V0 ;
      RECT 1.6640 5.0240 1.6960 5.0560 ;
    LAYER V0 ;
      RECT 1.6640 5.0240 1.6960 5.0560 ;
    LAYER V0 ;
      RECT 1.6640 5.0240 1.6960 5.0560 ;
    LAYER V0 ;
      RECT 1.6640 5.0240 1.6960 5.0560 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.8240 2.7560 1.8560 2.7880 ;
    LAYER V0 ;
      RECT 1.8240 2.8820 1.8560 2.9140 ;
    LAYER V0 ;
      RECT 1.8240 3.0080 1.8560 3.0400 ;
    LAYER V0 ;
      RECT 1.8240 3.9320 1.8560 3.9640 ;
    LAYER V0 ;
      RECT 1.8240 4.0580 1.8560 4.0900 ;
    LAYER V0 ;
      RECT 1.8240 4.1840 1.8560 4.2160 ;
  END
END Switch_PMOS_nfin240_n12_X5_Y4_ST2_RVT
MACRO DP_NMOS_B_nfin28_n12_X3_Y1_RVT
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin28_n12_X3_Y1_RVT 0 0 ;
  SIZE 1.4400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 1.2360 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.1520 0.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.2360 1.1560 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.9080 0.9960 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.4440 0.9920 1.1560 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 1.4960 1.1560 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.0480 0.4960 0.7920 ;
    LAYER M1 ;
      RECT 0.4640 0.8880 0.4960 1.1280 ;
    LAYER M1 ;
      RECT 0.4640 1.3920 0.4960 1.6320 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.0480 0.6560 0.7920 ;
    LAYER M1 ;
      RECT 0.6240 0.8880 0.6560 1.1280 ;
    LAYER M1 ;
      RECT 0.6240 1.3920 0.6560 1.6320 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.0480 0.8160 0.7920 ;
    LAYER M1 ;
      RECT 0.7840 0.8880 0.8160 1.1280 ;
    LAYER M1 ;
      RECT 0.7840 1.3920 0.8160 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7920 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.1280 ;
    LAYER M1 ;
      RECT 0.9440 1.3920 0.9760 1.6320 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.0480 1.1360 0.7920 ;
    LAYER M1 ;
      RECT 1.1040 0.8880 1.1360 1.1280 ;
    LAYER M1 ;
      RECT 1.1040 1.3920 1.1360 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.7040 0.0680 0.7360 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.0240 0.0680 1.0560 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 0.6240 0.1520 0.6560 0.1840 ;
    LAYER V1 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V1 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V1 ;
      RECT 0.9440 0.1520 0.9760 0.1840 ;
    LAYER V1 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V1 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.7840 0.2360 0.8160 0.2680 ;
    LAYER V1 ;
      RECT 0.7840 0.9920 0.8160 1.0240 ;
    LAYER V1 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V1 ;
      RECT 0.4640 0.2360 0.4960 0.2680 ;
    LAYER V1 ;
      RECT 0.4640 0.9920 0.4960 1.0240 ;
    LAYER V1 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V1 ;
      RECT 1.1040 0.2360 1.1360 0.2680 ;
    LAYER V1 ;
      RECT 1.1040 0.9920 1.1360 1.0240 ;
    LAYER V1 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.4040 0.4960 0.4360 ;
    LAYER V0 ;
      RECT 0.4640 0.5300 0.4960 0.5620 ;
    LAYER V0 ;
      RECT 0.4640 0.6560 0.4960 0.6880 ;
    LAYER V0 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V0 ;
      RECT 0.4640 1.4960 0.4960 1.5280 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.4040 0.6560 0.4360 ;
    LAYER V0 ;
      RECT 0.6240 0.5300 0.6560 0.5620 ;
    LAYER V0 ;
      RECT 0.6240 0.6560 0.6560 0.6880 ;
    LAYER V0 ;
      RECT 0.6240 0.9080 0.6560 0.9400 ;
    LAYER V0 ;
      RECT 0.6240 1.4960 0.6560 1.5280 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.4040 0.8160 0.4360 ;
    LAYER V0 ;
      RECT 0.7840 0.5300 0.8160 0.5620 ;
    LAYER V0 ;
      RECT 0.7840 0.6560 0.8160 0.6880 ;
    LAYER V0 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V0 ;
      RECT 0.7840 1.4960 0.8160 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.4040 0.9760 0.4360 ;
    LAYER V0 ;
      RECT 0.9440 0.5300 0.9760 0.5620 ;
    LAYER V0 ;
      RECT 0.9440 0.6560 0.9760 0.6880 ;
    LAYER V0 ;
      RECT 0.9440 0.9080 0.9760 0.9400 ;
    LAYER V0 ;
      RECT 0.9440 1.4960 0.9760 1.5280 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.4040 1.1360 0.4360 ;
    LAYER V0 ;
      RECT 1.1040 0.5300 1.1360 0.5620 ;
    LAYER V0 ;
      RECT 1.1040 0.6560 1.1360 0.6880 ;
    LAYER V0 ;
      RECT 1.1040 0.9080 1.1360 0.9400 ;
    LAYER V0 ;
      RECT 1.1040 1.4960 1.1360 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
  END
END DP_NMOS_B_nfin28_n12_X3_Y1_RVT
