MACRO SCM_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT 0 0 ;
  SIZE 3.0400 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2600 0.0480 1.3000 2.7240 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3400 0.1320 1.3800 2.1360 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4200 0.2160 1.4600 1.4640 ;
    END
  END DB
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.1280 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.0640 1.0560 2.3040 ;
    LAYER M1 ;
      RECT 1.0240 2.5680 1.0560 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.8880 1.3760 1.1280 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 2.0640 1.3760 2.3040 ;
    LAYER M1 ;
      RECT 1.3440 2.5680 1.3760 2.8080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.1280 ;
    LAYER M1 ;
      RECT 1.6640 1.2240 1.6960 1.9680 ;
    LAYER M1 ;
      RECT 1.6640 2.0640 1.6960 2.3040 ;
    LAYER M1 ;
      RECT 1.6640 2.5680 1.6960 2.8080 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.8240 1.2240 1.8560 1.9680 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 1.9840 0.8880 2.0160 1.1280 ;
    LAYER M1 ;
      RECT 1.9840 1.2240 2.0160 1.9680 ;
    LAYER M1 ;
      RECT 1.9840 2.0640 2.0160 2.3040 ;
    LAYER M1 ;
      RECT 1.9840 2.5680 2.0160 2.8080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.1440 1.2240 2.1760 1.9680 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.1280 ;
    LAYER M1 ;
      RECT 2.3040 1.2240 2.3360 1.9680 ;
    LAYER M1 ;
      RECT 2.3040 2.0640 2.3360 2.3040 ;
    LAYER M1 ;
      RECT 2.3040 2.5680 2.3360 2.8080 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER M1 ;
      RECT 2.4640 1.2240 2.4960 1.9680 ;
    LAYER M1 ;
      RECT 2.6240 0.0480 2.6560 0.7920 ;
    LAYER M1 ;
      RECT 2.6240 0.8880 2.6560 1.1280 ;
    LAYER M1 ;
      RECT 2.6240 1.2240 2.6560 1.9680 ;
    LAYER M1 ;
      RECT 2.6240 2.0640 2.6560 2.3040 ;
    LAYER M1 ;
      RECT 2.6240 2.5680 2.6560 2.8080 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER M1 ;
      RECT 2.7840 1.2240 2.8160 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 2.6760 0.9400 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.6760 0.1840 ;
    LAYER M2 ;
      RECT 0.6840 0.2360 2.3560 0.2680 ;
    LAYER M2 ;
      RECT 0.3640 2.6720 2.6760 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 2.8360 1.2760 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 2.6760 2.1160 ;
    LAYER M2 ;
      RECT 0.6840 1.3280 2.3560 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 1.4120 2.6760 1.4440 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 1.2440 2.8160 1.2760 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 1.2440 1.8560 1.2760 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 1.2440 2.1760 1.2760 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 1.2440 2.4960 1.2760 ;
    LAYER V1 ;
      RECT 2.6240 0.1520 2.6560 0.1840 ;
    LAYER V1 ;
      RECT 2.6240 0.9080 2.6560 0.9400 ;
    LAYER V1 ;
      RECT 2.6240 1.4120 2.6560 1.4440 ;
    LAYER V1 ;
      RECT 2.6240 2.0840 2.6560 2.1160 ;
    LAYER V1 ;
      RECT 2.6240 2.6720 2.6560 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.4120 0.4160 1.4440 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V1 ;
      RECT 0.7040 0.2360 0.7360 0.2680 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V1 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER V1 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V1 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V1 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V1 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V1 ;
      RECT 1.3440 1.4120 1.3760 1.4440 ;
    LAYER V1 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V1 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V1 ;
      RECT 1.6640 1.4120 1.6960 1.4440 ;
    LAYER V1 ;
      RECT 1.6640 2.0840 1.6960 2.1160 ;
    LAYER V1 ;
      RECT 1.6640 2.6720 1.6960 2.7040 ;
    LAYER V1 ;
      RECT 1.9840 0.2360 2.0160 0.2680 ;
    LAYER V1 ;
      RECT 1.9840 0.9080 2.0160 0.9400 ;
    LAYER V1 ;
      RECT 1.9840 1.3280 2.0160 1.3600 ;
    LAYER V1 ;
      RECT 1.9840 2.0840 2.0160 2.1160 ;
    LAYER V1 ;
      RECT 1.9840 2.6720 2.0160 2.7040 ;
    LAYER V1 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V1 ;
      RECT 2.3040 0.9080 2.3360 0.9400 ;
    LAYER V1 ;
      RECT 2.3040 1.3280 2.3360 1.3600 ;
    LAYER V1 ;
      RECT 2.3040 2.0840 2.3360 2.1160 ;
    LAYER V1 ;
      RECT 2.3040 2.6720 2.3360 2.7040 ;
    LAYER V2 ;
      RECT 1.2640 0.0680 1.2960 0.1000 ;
    LAYER V2 ;
      RECT 1.2640 1.2440 1.2960 1.2760 ;
    LAYER V2 ;
      RECT 1.2640 2.6720 1.2960 2.7040 ;
    LAYER V2 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V2 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V2 ;
      RECT 1.3440 1.3280 1.3760 1.3600 ;
    LAYER V2 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V2 ;
      RECT 1.4240 0.2360 1.4560 0.2680 ;
    LAYER V2 ;
      RECT 1.4240 1.4120 1.4560 1.4440 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V0 ;
      RECT 1.6640 1.5800 1.6960 1.6120 ;
    LAYER V0 ;
      RECT 1.6640 1.7060 1.6960 1.7380 ;
    LAYER V0 ;
      RECT 1.6640 1.8320 1.6960 1.8640 ;
    LAYER V0 ;
      RECT 1.6640 2.0840 1.6960 2.1160 ;
    LAYER V0 ;
      RECT 1.6640 2.6720 1.6960 2.7040 ;
    LAYER V0 ;
      RECT 1.6640 2.6720 1.6960 2.7040 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.5800 1.8560 1.6120 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.7060 1.8560 1.7380 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.8240 1.8320 1.8560 1.8640 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.9080 2.0160 0.9400 ;
    LAYER V0 ;
      RECT 1.9840 1.5800 2.0160 1.6120 ;
    LAYER V0 ;
      RECT 1.9840 1.7060 2.0160 1.7380 ;
    LAYER V0 ;
      RECT 1.9840 1.8320 2.0160 1.8640 ;
    LAYER V0 ;
      RECT 1.9840 2.0840 2.0160 2.1160 ;
    LAYER V0 ;
      RECT 1.9840 2.6720 2.0160 2.7040 ;
    LAYER V0 ;
      RECT 1.9840 2.6720 2.0160 2.7040 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.5800 2.1760 1.6120 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.7060 2.1760 1.7380 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.1440 1.8320 2.1760 1.8640 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.9080 2.3360 0.9400 ;
    LAYER V0 ;
      RECT 2.3040 1.5800 2.3360 1.6120 ;
    LAYER V0 ;
      RECT 2.3040 1.7060 2.3360 1.7380 ;
    LAYER V0 ;
      RECT 2.3040 1.8320 2.3360 1.8640 ;
    LAYER V0 ;
      RECT 2.3040 2.0840 2.3360 2.1160 ;
    LAYER V0 ;
      RECT 2.3040 2.6720 2.3360 2.7040 ;
    LAYER V0 ;
      RECT 2.3040 2.6720 2.3360 2.7040 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.5800 2.4960 1.6120 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.7060 2.4960 1.7380 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.4640 1.8320 2.4960 1.8640 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.9080 2.6560 0.9400 ;
    LAYER V0 ;
      RECT 2.6240 1.5800 2.6560 1.6120 ;
    LAYER V0 ;
      RECT 2.6240 1.7060 2.6560 1.7380 ;
    LAYER V0 ;
      RECT 2.6240 1.8320 2.6560 1.8640 ;
    LAYER V0 ;
      RECT 2.6240 2.0840 2.6560 2.1160 ;
    LAYER V0 ;
      RECT 2.6240 2.6720 2.6560 2.7040 ;
    LAYER V0 ;
      RECT 2.6240 2.6720 2.6560 2.7040 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.7840 1.5800 2.8160 1.6120 ;
    LAYER V0 ;
      RECT 2.7840 1.7060 2.8160 1.7380 ;
    LAYER V0 ;
      RECT 2.7840 1.8320 2.8160 1.8640 ;
  END
END SCM_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
MACRO DCL_PMOS_nfin6_m8_n12_X2_Y2_ST2_LVT
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_nfin6_m8_n12_X2_Y2_ST2_LVT 0 0 ;
  SIZE 1.1200 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 2.1360 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 0.7560 0.9400 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 0.7560 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 2.6720 0.7560 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 0.9160 1.2760 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 0.7560 2.1160 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 0.7560 1.3600 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V2 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V2 ;
      RECT 0.3840 1.2440 0.4160 1.2760 ;
    LAYER V2 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V2 ;
      RECT 0.4640 0.1520 0.4960 0.1840 ;
    LAYER V2 ;
      RECT 0.4640 0.9080 0.4960 0.9400 ;
    LAYER V2 ;
      RECT 0.4640 1.3280 0.4960 1.3600 ;
    LAYER V2 ;
      RECT 0.4640 2.0840 0.4960 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
  END
END DCL_PMOS_nfin6_m8_n12_X2_Y2_ST2_LVT
MACRO DP_NMOS_B_nfin6_m16_n12_X8_Y1_ST2_LVT
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_nfin6_m16_n12_X8_Y1_ST2_LVT 0 0 ;
  SIZE 5.6000 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 5.3960 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 5.2360 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6840 0.2360 4.9160 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.9080 5.2360 0.9400 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.6840 0.9920 4.9160 1.0240 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 1.4960 5.2360 1.5280 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.3920 0.4160 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.3920 0.7360 1.6320 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.1280 ;
    LAYER M1 ;
      RECT 1.0240 1.3920 1.0560 1.6320 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.8880 1.3760 1.1280 ;
    LAYER M1 ;
      RECT 1.3440 1.3920 1.3760 1.6320 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7920 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.1280 ;
    LAYER M1 ;
      RECT 1.6640 1.3920 1.6960 1.6320 ;
    LAYER M1 ;
      RECT 1.8240 0.0480 1.8560 0.7920 ;
    LAYER M1 ;
      RECT 1.9840 0.0480 2.0160 0.7920 ;
    LAYER M1 ;
      RECT 1.9840 0.8880 2.0160 1.1280 ;
    LAYER M1 ;
      RECT 1.9840 1.3920 2.0160 1.6320 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7920 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.1280 ;
    LAYER M1 ;
      RECT 2.3040 1.3920 2.3360 1.6320 ;
    LAYER M1 ;
      RECT 2.4640 0.0480 2.4960 0.7920 ;
    LAYER M1 ;
      RECT 2.6240 0.0480 2.6560 0.7920 ;
    LAYER M1 ;
      RECT 2.6240 0.8880 2.6560 1.1280 ;
    LAYER M1 ;
      RECT 2.6240 1.3920 2.6560 1.6320 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7920 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7920 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.1280 ;
    LAYER M1 ;
      RECT 2.9440 1.3920 2.9760 1.6320 ;
    LAYER M1 ;
      RECT 3.1040 0.0480 3.1360 0.7920 ;
    LAYER M1 ;
      RECT 3.2640 0.0480 3.2960 0.7920 ;
    LAYER M1 ;
      RECT 3.2640 0.8880 3.2960 1.1280 ;
    LAYER M1 ;
      RECT 3.2640 1.3920 3.2960 1.6320 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7920 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7920 ;
    LAYER M1 ;
      RECT 3.5840 0.8880 3.6160 1.1280 ;
    LAYER M1 ;
      RECT 3.5840 1.3920 3.6160 1.6320 ;
    LAYER M1 ;
      RECT 3.7440 0.0480 3.7760 0.7920 ;
    LAYER M1 ;
      RECT 3.9040 0.0480 3.9360 0.7920 ;
    LAYER M1 ;
      RECT 3.9040 0.8880 3.9360 1.1280 ;
    LAYER M1 ;
      RECT 3.9040 1.3920 3.9360 1.6320 ;
    LAYER M1 ;
      RECT 4.0640 0.0480 4.0960 0.7920 ;
    LAYER M1 ;
      RECT 4.2240 0.0480 4.2560 0.7920 ;
    LAYER M1 ;
      RECT 4.2240 0.8880 4.2560 1.1280 ;
    LAYER M1 ;
      RECT 4.2240 1.3920 4.2560 1.6320 ;
    LAYER M1 ;
      RECT 4.3840 0.0480 4.4160 0.7920 ;
    LAYER M1 ;
      RECT 4.5440 0.0480 4.5760 0.7920 ;
    LAYER M1 ;
      RECT 4.5440 0.8880 4.5760 1.1280 ;
    LAYER M1 ;
      RECT 4.5440 1.3920 4.5760 1.6320 ;
    LAYER M1 ;
      RECT 4.7040 0.0480 4.7360 0.7920 ;
    LAYER M1 ;
      RECT 4.8640 0.0480 4.8960 0.7920 ;
    LAYER M1 ;
      RECT 4.8640 0.8880 4.8960 1.1280 ;
    LAYER M1 ;
      RECT 4.8640 1.3920 4.8960 1.6320 ;
    LAYER M1 ;
      RECT 5.0240 0.0480 5.0560 0.7920 ;
    LAYER M1 ;
      RECT 5.1840 0.0480 5.2160 0.7920 ;
    LAYER M1 ;
      RECT 5.1840 0.8880 5.2160 1.1280 ;
    LAYER M1 ;
      RECT 5.1840 1.3920 5.2160 1.6320 ;
    LAYER M1 ;
      RECT 5.3440 0.0480 5.3760 0.7920 ;
    LAYER V1 ;
      RECT 5.3440 0.0680 5.3760 0.1000 ;
    LAYER V1 ;
      RECT 2.7840 0.0680 2.8160 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 3.1040 0.0680 3.1360 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 4.7040 0.0680 4.7360 0.1000 ;
    LAYER V1 ;
      RECT 3.4240 0.0680 3.4560 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 3.7440 0.0680 3.7760 0.1000 ;
    LAYER V1 ;
      RECT 4.0640 0.0680 4.0960 0.1000 ;
    LAYER V1 ;
      RECT 1.8240 0.0680 1.8560 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 4.3840 0.0680 4.4160 0.1000 ;
    LAYER V1 ;
      RECT 2.1440 0.0680 2.1760 0.1000 ;
    LAYER V1 ;
      RECT 5.0240 0.0680 5.0560 0.1000 ;
    LAYER V1 ;
      RECT 2.4640 0.0680 2.4960 0.1000 ;
    LAYER V1 ;
      RECT 2.6240 0.1520 2.6560 0.1840 ;
    LAYER V1 ;
      RECT 2.6240 0.9080 2.6560 0.9400 ;
    LAYER V1 ;
      RECT 2.6240 1.4960 2.6560 1.5280 ;
    LAYER V1 ;
      RECT 5.1840 0.1520 5.2160 0.1840 ;
    LAYER V1 ;
      RECT 5.1840 0.9080 5.2160 0.9400 ;
    LAYER V1 ;
      RECT 5.1840 1.4960 5.2160 1.5280 ;
    LAYER V1 ;
      RECT 2.9440 0.1520 2.9760 0.1840 ;
    LAYER V1 ;
      RECT 2.9440 0.9080 2.9760 0.9400 ;
    LAYER V1 ;
      RECT 2.9440 1.4960 2.9760 1.5280 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.4960 0.4160 1.5280 ;
    LAYER V1 ;
      RECT 3.9040 0.1520 3.9360 0.1840 ;
    LAYER V1 ;
      RECT 3.9040 0.9080 3.9360 0.9400 ;
    LAYER V1 ;
      RECT 3.9040 1.4960 3.9360 1.5280 ;
    LAYER V1 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V1 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V1 ;
      RECT 1.3440 1.4960 1.3760 1.5280 ;
    LAYER V1 ;
      RECT 1.6640 0.1520 1.6960 0.1840 ;
    LAYER V1 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V1 ;
      RECT 1.6640 1.4960 1.6960 1.5280 ;
    LAYER V1 ;
      RECT 4.2240 0.1520 4.2560 0.1840 ;
    LAYER V1 ;
      RECT 4.2240 0.9080 4.2560 0.9400 ;
    LAYER V1 ;
      RECT 4.2240 1.4960 4.2560 1.5280 ;
    LAYER V1 ;
      RECT 0.7040 0.2360 0.7360 0.2680 ;
    LAYER V1 ;
      RECT 0.7040 0.9920 0.7360 1.0240 ;
    LAYER V1 ;
      RECT 0.7040 1.4960 0.7360 1.5280 ;
    LAYER V1 ;
      RECT 3.2640 0.2360 3.2960 0.2680 ;
    LAYER V1 ;
      RECT 3.2640 0.9920 3.2960 1.0240 ;
    LAYER V1 ;
      RECT 3.2640 1.4960 3.2960 1.5280 ;
    LAYER V1 ;
      RECT 3.5840 0.2360 3.6160 0.2680 ;
    LAYER V1 ;
      RECT 3.5840 0.9920 3.6160 1.0240 ;
    LAYER V1 ;
      RECT 3.5840 1.4960 3.6160 1.5280 ;
    LAYER V1 ;
      RECT 1.0240 0.2360 1.0560 0.2680 ;
    LAYER V1 ;
      RECT 1.0240 0.9920 1.0560 1.0240 ;
    LAYER V1 ;
      RECT 1.0240 1.4960 1.0560 1.5280 ;
    LAYER V1 ;
      RECT 2.3040 0.2360 2.3360 0.2680 ;
    LAYER V1 ;
      RECT 2.3040 0.9920 2.3360 1.0240 ;
    LAYER V1 ;
      RECT 2.3040 1.4960 2.3360 1.5280 ;
    LAYER V1 ;
      RECT 1.9840 0.2360 2.0160 0.2680 ;
    LAYER V1 ;
      RECT 1.9840 0.9920 2.0160 1.0240 ;
    LAYER V1 ;
      RECT 1.9840 1.4960 2.0160 1.5280 ;
    LAYER V1 ;
      RECT 4.8640 0.2360 4.8960 0.2680 ;
    LAYER V1 ;
      RECT 4.8640 0.9920 4.8960 1.0240 ;
    LAYER V1 ;
      RECT 4.8640 1.4960 4.8960 1.5280 ;
    LAYER V1 ;
      RECT 4.5440 0.2360 4.5760 0.2680 ;
    LAYER V1 ;
      RECT 4.5440 0.9920 4.5760 1.0240 ;
    LAYER V1 ;
      RECT 4.5440 1.4960 4.5760 1.5280 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.4960 0.4160 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.4960 0.7360 1.5280 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 1.0240 1.4960 1.0560 1.5280 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V0 ;
      RECT 1.3440 1.4960 1.3760 1.5280 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.4040 1.6960 0.4360 ;
    LAYER V0 ;
      RECT 1.6640 0.5300 1.6960 0.5620 ;
    LAYER V0 ;
      RECT 1.6640 0.6560 1.6960 0.6880 ;
    LAYER V0 ;
      RECT 1.6640 0.9080 1.6960 0.9400 ;
    LAYER V0 ;
      RECT 1.6640 1.4960 1.6960 1.5280 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.4040 1.8560 0.4360 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.5300 1.8560 0.5620 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.8240 0.6560 1.8560 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.4040 2.0160 0.4360 ;
    LAYER V0 ;
      RECT 1.9840 0.5300 2.0160 0.5620 ;
    LAYER V0 ;
      RECT 1.9840 0.6560 2.0160 0.6880 ;
    LAYER V0 ;
      RECT 1.9840 0.9080 2.0160 0.9400 ;
    LAYER V0 ;
      RECT 1.9840 1.4960 2.0160 1.5280 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.4040 2.1760 0.4360 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.5300 2.1760 0.5620 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.1440 0.6560 2.1760 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.4040 2.3360 0.4360 ;
    LAYER V0 ;
      RECT 2.3040 0.5300 2.3360 0.5620 ;
    LAYER V0 ;
      RECT 2.3040 0.6560 2.3360 0.6880 ;
    LAYER V0 ;
      RECT 2.3040 0.9080 2.3360 0.9400 ;
    LAYER V0 ;
      RECT 2.3040 1.4960 2.3360 1.5280 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.4040 2.4960 0.4360 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.5300 2.4960 0.5620 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.4640 0.6560 2.4960 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.4040 2.6560 0.4360 ;
    LAYER V0 ;
      RECT 2.6240 0.5300 2.6560 0.5620 ;
    LAYER V0 ;
      RECT 2.6240 0.6560 2.6560 0.6880 ;
    LAYER V0 ;
      RECT 2.6240 0.9080 2.6560 0.9400 ;
    LAYER V0 ;
      RECT 2.6240 1.4960 2.6560 1.5280 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.4040 2.8160 0.4360 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.5300 2.8160 0.5620 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.7840 0.6560 2.8160 0.6880 ;
    LAYER V0 ;
      RECT 2.9440 0.4040 2.9760 0.4360 ;
    LAYER V0 ;
      RECT 2.9440 0.5300 2.9760 0.5620 ;
    LAYER V0 ;
      RECT 2.9440 0.6560 2.9760 0.6880 ;
    LAYER V0 ;
      RECT 2.9440 0.9080 2.9760 0.9400 ;
    LAYER V0 ;
      RECT 2.9440 1.4960 2.9760 1.5280 ;
    LAYER V0 ;
      RECT 3.1040 0.4040 3.1360 0.4360 ;
    LAYER V0 ;
      RECT 3.1040 0.4040 3.1360 0.4360 ;
    LAYER V0 ;
      RECT 3.1040 0.5300 3.1360 0.5620 ;
    LAYER V0 ;
      RECT 3.1040 0.5300 3.1360 0.5620 ;
    LAYER V0 ;
      RECT 3.1040 0.6560 3.1360 0.6880 ;
    LAYER V0 ;
      RECT 3.1040 0.6560 3.1360 0.6880 ;
    LAYER V0 ;
      RECT 3.2640 0.4040 3.2960 0.4360 ;
    LAYER V0 ;
      RECT 3.2640 0.5300 3.2960 0.5620 ;
    LAYER V0 ;
      RECT 3.2640 0.6560 3.2960 0.6880 ;
    LAYER V0 ;
      RECT 3.2640 0.9080 3.2960 0.9400 ;
    LAYER V0 ;
      RECT 3.2640 1.4960 3.2960 1.5280 ;
    LAYER V0 ;
      RECT 3.4240 0.4040 3.4560 0.4360 ;
    LAYER V0 ;
      RECT 3.4240 0.4040 3.4560 0.4360 ;
    LAYER V0 ;
      RECT 3.4240 0.5300 3.4560 0.5620 ;
    LAYER V0 ;
      RECT 3.4240 0.5300 3.4560 0.5620 ;
    LAYER V0 ;
      RECT 3.4240 0.6560 3.4560 0.6880 ;
    LAYER V0 ;
      RECT 3.4240 0.6560 3.4560 0.6880 ;
    LAYER V0 ;
      RECT 3.5840 0.4040 3.6160 0.4360 ;
    LAYER V0 ;
      RECT 3.5840 0.5300 3.6160 0.5620 ;
    LAYER V0 ;
      RECT 3.5840 0.6560 3.6160 0.6880 ;
    LAYER V0 ;
      RECT 3.5840 0.9080 3.6160 0.9400 ;
    LAYER V0 ;
      RECT 3.5840 1.4960 3.6160 1.5280 ;
    LAYER V0 ;
      RECT 3.7440 0.4040 3.7760 0.4360 ;
    LAYER V0 ;
      RECT 3.7440 0.4040 3.7760 0.4360 ;
    LAYER V0 ;
      RECT 3.7440 0.5300 3.7760 0.5620 ;
    LAYER V0 ;
      RECT 3.7440 0.5300 3.7760 0.5620 ;
    LAYER V0 ;
      RECT 3.7440 0.6560 3.7760 0.6880 ;
    LAYER V0 ;
      RECT 3.7440 0.6560 3.7760 0.6880 ;
    LAYER V0 ;
      RECT 3.9040 0.4040 3.9360 0.4360 ;
    LAYER V0 ;
      RECT 3.9040 0.5300 3.9360 0.5620 ;
    LAYER V0 ;
      RECT 3.9040 0.6560 3.9360 0.6880 ;
    LAYER V0 ;
      RECT 3.9040 0.9080 3.9360 0.9400 ;
    LAYER V0 ;
      RECT 3.9040 1.4960 3.9360 1.5280 ;
    LAYER V0 ;
      RECT 4.0640 0.4040 4.0960 0.4360 ;
    LAYER V0 ;
      RECT 4.0640 0.4040 4.0960 0.4360 ;
    LAYER V0 ;
      RECT 4.0640 0.5300 4.0960 0.5620 ;
    LAYER V0 ;
      RECT 4.0640 0.5300 4.0960 0.5620 ;
    LAYER V0 ;
      RECT 4.0640 0.6560 4.0960 0.6880 ;
    LAYER V0 ;
      RECT 4.0640 0.6560 4.0960 0.6880 ;
    LAYER V0 ;
      RECT 4.2240 0.4040 4.2560 0.4360 ;
    LAYER V0 ;
      RECT 4.2240 0.5300 4.2560 0.5620 ;
    LAYER V0 ;
      RECT 4.2240 0.6560 4.2560 0.6880 ;
    LAYER V0 ;
      RECT 4.2240 0.9080 4.2560 0.9400 ;
    LAYER V0 ;
      RECT 4.2240 1.4960 4.2560 1.5280 ;
    LAYER V0 ;
      RECT 4.3840 0.4040 4.4160 0.4360 ;
    LAYER V0 ;
      RECT 4.3840 0.4040 4.4160 0.4360 ;
    LAYER V0 ;
      RECT 4.3840 0.5300 4.4160 0.5620 ;
    LAYER V0 ;
      RECT 4.3840 0.5300 4.4160 0.5620 ;
    LAYER V0 ;
      RECT 4.3840 0.6560 4.4160 0.6880 ;
    LAYER V0 ;
      RECT 4.3840 0.6560 4.4160 0.6880 ;
    LAYER V0 ;
      RECT 4.5440 0.4040 4.5760 0.4360 ;
    LAYER V0 ;
      RECT 4.5440 0.5300 4.5760 0.5620 ;
    LAYER V0 ;
      RECT 4.5440 0.6560 4.5760 0.6880 ;
    LAYER V0 ;
      RECT 4.5440 0.9080 4.5760 0.9400 ;
    LAYER V0 ;
      RECT 4.5440 1.4960 4.5760 1.5280 ;
    LAYER V0 ;
      RECT 4.7040 0.4040 4.7360 0.4360 ;
    LAYER V0 ;
      RECT 4.7040 0.4040 4.7360 0.4360 ;
    LAYER V0 ;
      RECT 4.7040 0.5300 4.7360 0.5620 ;
    LAYER V0 ;
      RECT 4.7040 0.5300 4.7360 0.5620 ;
    LAYER V0 ;
      RECT 4.7040 0.6560 4.7360 0.6880 ;
    LAYER V0 ;
      RECT 4.7040 0.6560 4.7360 0.6880 ;
    LAYER V0 ;
      RECT 4.8640 0.4040 4.8960 0.4360 ;
    LAYER V0 ;
      RECT 4.8640 0.5300 4.8960 0.5620 ;
    LAYER V0 ;
      RECT 4.8640 0.6560 4.8960 0.6880 ;
    LAYER V0 ;
      RECT 4.8640 0.9080 4.8960 0.9400 ;
    LAYER V0 ;
      RECT 4.8640 1.4960 4.8960 1.5280 ;
    LAYER V0 ;
      RECT 5.0240 0.4040 5.0560 0.4360 ;
    LAYER V0 ;
      RECT 5.0240 0.4040 5.0560 0.4360 ;
    LAYER V0 ;
      RECT 5.0240 0.5300 5.0560 0.5620 ;
    LAYER V0 ;
      RECT 5.0240 0.5300 5.0560 0.5620 ;
    LAYER V0 ;
      RECT 5.0240 0.6560 5.0560 0.6880 ;
    LAYER V0 ;
      RECT 5.0240 0.6560 5.0560 0.6880 ;
    LAYER V0 ;
      RECT 5.1840 0.4040 5.2160 0.4360 ;
    LAYER V0 ;
      RECT 5.1840 0.5300 5.2160 0.5620 ;
    LAYER V0 ;
      RECT 5.1840 0.6560 5.2160 0.6880 ;
    LAYER V0 ;
      RECT 5.1840 0.9080 5.2160 0.9400 ;
    LAYER V0 ;
      RECT 5.1840 1.4960 5.2160 1.5280 ;
    LAYER V0 ;
      RECT 5.3440 0.4040 5.3760 0.4360 ;
    LAYER V0 ;
      RECT 5.3440 0.5300 5.3760 0.5620 ;
    LAYER V0 ;
      RECT 5.3440 0.6560 5.3760 0.6880 ;
  END
END DP_NMOS_B_nfin6_m16_n12_X8_Y1_ST2_LVT
MACRO Switch_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT 0 0 ;
  SIZE 1.7600 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.0480 0.6600 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7000 0.1320 0.7400 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.8880 0.8200 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.1280 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.0640 1.0560 2.3040 ;
    LAYER M1 ;
      RECT 1.0240 2.5680 1.0560 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.8880 1.3760 1.1280 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 2.0640 1.3760 2.3040 ;
    LAYER M1 ;
      RECT 1.3440 2.5680 1.3760 2.8080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.3960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 1.3960 0.9400 ;
    LAYER M2 ;
      RECT 0.3640 2.6720 1.3960 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.5560 1.2760 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 1.3960 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 1.3960 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V1 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER V1 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V1 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V1 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V1 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V1 ;
      RECT 1.3440 1.3280 1.3760 1.3600 ;
    LAYER V1 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V1 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V2 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER V2 ;
      RECT 0.6240 1.2440 0.6560 1.2760 ;
    LAYER V2 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V2 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V2 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V2 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V2 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
  END
END Switch_NMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
MACRO Switch_PMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_nfin6_m16_n12_X4_Y2_ST2_LVT 0 0 ;
  SIZE 1.7600 BY 3.0240 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.0480 0.6600 2.7240 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7000 0.1320 0.7400 1.3800 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.8880 0.8200 2.1360 ;
    END
  END G
  OBS
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.1280 ;
    LAYER M1 ;
      RECT 0.3840 1.2240 0.4160 1.9680 ;
    LAYER M1 ;
      RECT 0.3840 2.0640 0.4160 2.3040 ;
    LAYER M1 ;
      RECT 0.3840 2.5680 0.4160 2.8080 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.2240 1.2240 0.2560 1.9680 ;
    LAYER M1 ;
      RECT 0.5440 0.0480 0.5760 0.7920 ;
    LAYER M1 ;
      RECT 0.5440 1.2240 0.5760 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 0.0480 0.7360 0.7920 ;
    LAYER M1 ;
      RECT 0.7040 0.8880 0.7360 1.1280 ;
    LAYER M1 ;
      RECT 0.7040 1.2240 0.7360 1.9680 ;
    LAYER M1 ;
      RECT 0.7040 2.0640 0.7360 2.3040 ;
    LAYER M1 ;
      RECT 0.7040 2.5680 0.7360 2.8080 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7920 ;
    LAYER M1 ;
      RECT 0.8640 1.2240 0.8960 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7920 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.1280 ;
    LAYER M1 ;
      RECT 1.0240 1.2240 1.0560 1.9680 ;
    LAYER M1 ;
      RECT 1.0240 2.0640 1.0560 2.3040 ;
    LAYER M1 ;
      RECT 1.0240 2.5680 1.0560 2.8080 ;
    LAYER M1 ;
      RECT 1.1840 0.0480 1.2160 0.7920 ;
    LAYER M1 ;
      RECT 1.1840 1.2240 1.2160 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 0.0480 1.3760 0.7920 ;
    LAYER M1 ;
      RECT 1.3440 0.8880 1.3760 1.1280 ;
    LAYER M1 ;
      RECT 1.3440 1.2240 1.3760 1.9680 ;
    LAYER M1 ;
      RECT 1.3440 2.0640 1.3760 2.3040 ;
    LAYER M1 ;
      RECT 1.3440 2.5680 1.3760 2.8080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7920 ;
    LAYER M1 ;
      RECT 1.5040 1.2240 1.5360 1.9680 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.3960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.9080 1.3960 0.9400 ;
    LAYER M2 ;
      RECT 0.3640 2.6720 1.3960 2.7040 ;
    LAYER M2 ;
      RECT 0.2040 1.2440 1.5560 1.2760 ;
    LAYER M2 ;
      RECT 0.3640 1.3280 1.3960 1.3600 ;
    LAYER M2 ;
      RECT 0.3640 2.0840 1.3960 2.1160 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.2240 1.2440 0.2560 1.2760 ;
    LAYER V1 ;
      RECT 0.5440 0.0680 0.5760 0.1000 ;
    LAYER V1 ;
      RECT 0.5440 1.2440 0.5760 1.2760 ;
    LAYER V1 ;
      RECT 0.8640 0.0680 0.8960 0.1000 ;
    LAYER V1 ;
      RECT 0.8640 1.2440 0.8960 1.2760 ;
    LAYER V1 ;
      RECT 1.1840 0.0680 1.2160 0.1000 ;
    LAYER V1 ;
      RECT 1.1840 1.2440 1.2160 1.2760 ;
    LAYER V1 ;
      RECT 1.5040 0.0680 1.5360 0.1000 ;
    LAYER V1 ;
      RECT 1.5040 1.2440 1.5360 1.2760 ;
    LAYER V1 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V1 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V1 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V1 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V1 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V1 ;
      RECT 0.3840 0.1520 0.4160 0.1840 ;
    LAYER V1 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V1 ;
      RECT 0.3840 1.3280 0.4160 1.3600 ;
    LAYER V1 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V1 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V1 ;
      RECT 1.0240 0.1520 1.0560 0.1840 ;
    LAYER V1 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V1 ;
      RECT 1.0240 1.3280 1.0560 1.3600 ;
    LAYER V1 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V1 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V1 ;
      RECT 1.3440 0.1520 1.3760 0.1840 ;
    LAYER V1 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V1 ;
      RECT 1.3440 1.3280 1.3760 1.3600 ;
    LAYER V1 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V1 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V2 ;
      RECT 0.6240 0.0680 0.6560 0.1000 ;
    LAYER V2 ;
      RECT 0.6240 1.2440 0.6560 1.2760 ;
    LAYER V2 ;
      RECT 0.6240 2.6720 0.6560 2.7040 ;
    LAYER V2 ;
      RECT 0.7040 0.1520 0.7360 0.1840 ;
    LAYER V2 ;
      RECT 0.7040 1.3280 0.7360 1.3600 ;
    LAYER V2 ;
      RECT 0.7840 0.9080 0.8160 0.9400 ;
    LAYER V2 ;
      RECT 0.7840 2.0840 0.8160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 0.4160 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 1.5800 0.4160 1.6120 ;
    LAYER V0 ;
      RECT 0.3840 1.7060 0.4160 1.7380 ;
    LAYER V0 ;
      RECT 0.3840 1.8320 0.4160 1.8640 ;
    LAYER V0 ;
      RECT 0.3840 2.0840 0.4160 2.1160 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.3840 2.6720 0.4160 2.7040 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.2240 1.5800 0.2560 1.6120 ;
    LAYER V0 ;
      RECT 0.2240 1.7060 0.2560 1.7380 ;
    LAYER V0 ;
      RECT 0.2240 1.8320 0.2560 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.4040 0.5760 0.4360 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.5300 0.5760 0.5620 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 0.6560 0.5760 0.6880 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.5800 0.5760 1.6120 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.7060 0.5760 1.7380 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.5440 1.8320 0.5760 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 0.4040 0.7360 0.4360 ;
    LAYER V0 ;
      RECT 0.7040 0.5300 0.7360 0.5620 ;
    LAYER V0 ;
      RECT 0.7040 0.6560 0.7360 0.6880 ;
    LAYER V0 ;
      RECT 0.7040 0.9080 0.7360 0.9400 ;
    LAYER V0 ;
      RECT 0.7040 1.5800 0.7360 1.6120 ;
    LAYER V0 ;
      RECT 0.7040 1.7060 0.7360 1.7380 ;
    LAYER V0 ;
      RECT 0.7040 1.8320 0.7360 1.8640 ;
    LAYER V0 ;
      RECT 0.7040 2.0840 0.7360 2.1160 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.7040 2.6720 0.7360 2.7040 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.4040 0.8960 0.4360 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.5300 0.8960 0.5620 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 0.6560 0.8960 0.6880 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.5800 0.8960 1.6120 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.7060 0.8960 1.7380 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 0.8640 1.8320 0.8960 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 1.0240 0.5300 1.0560 0.5620 ;
    LAYER V0 ;
      RECT 1.0240 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 1.0240 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 1.0240 1.5800 1.0560 1.6120 ;
    LAYER V0 ;
      RECT 1.0240 1.7060 1.0560 1.7380 ;
    LAYER V0 ;
      RECT 1.0240 1.8320 1.0560 1.8640 ;
    LAYER V0 ;
      RECT 1.0240 2.0840 1.0560 2.1160 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.0240 2.6720 1.0560 2.7040 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.4040 1.2160 0.4360 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.5300 1.2160 0.5620 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 0.6560 1.2160 0.6880 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.5800 1.2160 1.6120 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.7060 1.2160 1.7380 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.1840 1.8320 1.2160 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 0.4040 1.3760 0.4360 ;
    LAYER V0 ;
      RECT 1.3440 0.5300 1.3760 0.5620 ;
    LAYER V0 ;
      RECT 1.3440 0.6560 1.3760 0.6880 ;
    LAYER V0 ;
      RECT 1.3440 0.9080 1.3760 0.9400 ;
    LAYER V0 ;
      RECT 1.3440 1.5800 1.3760 1.6120 ;
    LAYER V0 ;
      RECT 1.3440 1.7060 1.3760 1.7380 ;
    LAYER V0 ;
      RECT 1.3440 1.8320 1.3760 1.8640 ;
    LAYER V0 ;
      RECT 1.3440 2.0840 1.3760 2.1160 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.3440 2.6720 1.3760 2.7040 ;
    LAYER V0 ;
      RECT 1.5040 0.4040 1.5360 0.4360 ;
    LAYER V0 ;
      RECT 1.5040 0.5300 1.5360 0.5620 ;
    LAYER V0 ;
      RECT 1.5040 0.6560 1.5360 0.6880 ;
    LAYER V0 ;
      RECT 1.5040 1.5800 1.5360 1.6120 ;
    LAYER V0 ;
      RECT 1.5040 1.7060 1.5360 1.7380 ;
    LAYER V0 ;
      RECT 1.5040 1.8320 1.5360 1.8640 ;
  END
END Switch_PMOS_nfin6_m16_n12_X4_Y2_ST2_LVT
MACRO Dummy_NMOS_nfin6_m1_n12_X1_Y1_LVT
  ORIGIN 0 0 ;
  FOREIGN Dummy_NMOS_nfin6_m1_n12_X1_Y1_LVT 0 0 ;
  SIZE 0.6400 BY 1.8480 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 1.5480 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1240 0.1520 0.3560 0.1840 ;
    END
  END D
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7920 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.1280 ;
    LAYER M1 ;
      RECT 0.3040 1.3920 0.3360 1.6320 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7920 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7920 ;
    LAYER M2 ;
      RECT 0.1240 0.9080 0.3560 0.9400 ;
    LAYER M2 ;
      RECT 0.1240 1.4960 0.3560 1.5280 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.4360 0.1000 ;
    LAYER V1 ;
      RECT 0.3040 0.1520 0.3360 0.1840 ;
    LAYER V1 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V1 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V1 ;
      RECT 0.2240 0.0680 0.2560 0.1000 ;
    LAYER V1 ;
      RECT 0.3840 0.0680 0.4160 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 0.0680 0.1760 0.1000 ;
    LAYER V2 ;
      RECT 0.1440 0.9080 0.1760 0.9400 ;
    LAYER V2 ;
      RECT 0.1440 1.4960 0.1760 1.5280 ;
    LAYER V0 ;
      RECT 0.3040 0.4040 0.3360 0.4360 ;
    LAYER V0 ;
      RECT 0.3040 0.5300 0.3360 0.5620 ;
    LAYER V0 ;
      RECT 0.3040 0.6560 0.3360 0.6880 ;
    LAYER V0 ;
      RECT 0.3040 0.9080 0.3360 0.9400 ;
    LAYER V0 ;
      RECT 0.3040 1.4960 0.3360 1.5280 ;
    LAYER V0 ;
      RECT 0.2240 0.4040 0.2560 0.4360 ;
    LAYER V0 ;
      RECT 0.2240 0.5300 0.2560 0.5620 ;
    LAYER V0 ;
      RECT 0.2240 0.6560 0.2560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.4040 0.4160 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.5300 0.4160 0.5620 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 0.4160 0.6880 ;
  END
END Dummy_NMOS_nfin6_m1_n12_X1_Y1_LVT
