MACRO guard_ring
  ORIGIN 0 0 ;
  FOREIGN guard_ring 0 0 ;
  SIZE 1.4400 BY 1.4280 ;
  PIN Body
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3440 0.3360 1.0960 1.0920 ;
    END
  END Body
  OBS
    LAYER V0 ;
      RECT 0.3840 0.4040 1.0560 0.4360 ;
    LAYER V0 ;
      RECT 0.3840 0.4880 1.0560 0.5200 ;
    LAYER V0 ;
      RECT 0.3840 0.5720 1.0560 0.6040 ;
    LAYER V0 ;
      RECT 0.3840 0.6560 1.0560 0.6880 ;
    LAYER V0 ;
      RECT 0.3840 0.7400 1.0560 0.7720 ;
    LAYER V0 ;
      RECT 0.3840 0.8240 1.0560 0.8560 ;
    LAYER V0 ;
      RECT 0.3840 0.9080 1.0560 0.9400 ;
    LAYER V0 ;
      RECT 0.3840 0.9920 1.0560 1.0240 ;
  END
END guard_ring