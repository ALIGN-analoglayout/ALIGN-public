.subckt powertrain_cell ond vcc vout
mmp0 vout ond vcc vcc p w=180n l=40n nfin=4 nf=8 m=4
.ends

.subckt powertrain_thermo on_d[63] on_d[62] on_d[61] on_d[60] on_d[59]
+ on_d[58] on_d[57] on_d[56] on_d[55] on_d[54] on_d[53] on_d[52] on_d[51] on_d[50]
+ on_d[49] on_d[48] on_d[47] on_d[46] on_d[45] on_d[44] on_d[43] on_d[42] on_d[41]
+ on_d[40] on_d[39] on_d[38] on_d[37] on_d[36] on_d[35] on_d[34] on_d[33] on_d[32]
+ on_d[31] on_d[30] on_d[29] on_d[28] on_d[27] on_d[26] on_d[25] on_d[24] on_d[23]
+ on_d[22] on_d[21] on_d[20] on_d[19] on_d[18] on_d[17] on_d[16] on_d[15] on_d[14]
+ on_d[13] on_d[12] on_d[11] on_d[10] on_d[9] on_d[8] on_d[7] on_d[6] on_d[5] on_d[4]
+ on_d[3] on_d[2] on_d[1] on_d[0] vcc vout
xu_pmos_title[63] on_d[63] vcc vout powertrain_cell
xu_pmos_title[62] on_d[62] vcc vout powertrain_cell
xu_pmos_title[61] on_d[61] vcc vout powertrain_cell
xu_pmos_title[60] on_d[60] vcc vout powertrain_cell
xu_pmos_title[59] on_d[59] vcc vout powertrain_cell
xu_pmos_title[58] on_d[58] vcc vout powertrain_cell
xu_pmos_title[57] on_d[57] vcc vout powertrain_cell
xu_pmos_title[56] on_d[56] vcc vout powertrain_cell
xu_pmos_title[55] on_d[55] vcc vout powertrain_cell
xu_pmos_title[54] on_d[54] vcc vout powertrain_cell
xu_pmos_title[53] on_d[53] vcc vout powertrain_cell
xu_pmos_title[52] on_d[52] vcc vout powertrain_cell
xu_pmos_title[51] on_d[51] vcc vout powertrain_cell
xu_pmos_title[50] on_d[50] vcc vout powertrain_cell
xu_pmos_title[49] on_d[49] vcc vout powertrain_cell
xu_pmos_title[48] on_d[48] vcc vout powertrain_cell
xu_pmos_title[47] on_d[47] vcc vout powertrain_cell
xu_pmos_title[46] on_d[46] vcc vout powertrain_cell
xu_pmos_title[45] on_d[45] vcc vout powertrain_cell
xu_pmos_title[44] on_d[44] vcc vout powertrain_cell
xu_pmos_title[43] on_d[43] vcc vout powertrain_cell
xu_pmos_title[42] on_d[42] vcc vout powertrain_cell
xu_pmos_title[41] on_d[41] vcc vout powertrain_cell
xu_pmos_title[40] on_d[40] vcc vout powertrain_cell
xu_pmos_title[39] on_d[39] vcc vout powertrain_cell
xu_pmos_title[38] on_d[38] vcc vout powertrain_cell
xu_pmos_title[37] on_d[37] vcc vout powertrain_cell
xu_pmos_title[36] on_d[36] vcc vout powertrain_cell
xu_pmos_title[35] on_d[35] vcc vout powertrain_cell
xu_pmos_title[34] on_d[34] vcc vout powertrain_cell
xu_pmos_title[33] on_d[33] vcc vout powertrain_cell
xu_pmos_title[32] on_d[32] vcc vout powertrain_cell
xu_pmos_title[31] on_d[31] vcc vout powertrain_cell
xu_pmos_title[30] on_d[30] vcc vout powertrain_cell
xu_pmos_title[29] on_d[29] vcc vout powertrain_cell
xu_pmos_title[28] on_d[28] vcc vout powertrain_cell
xu_pmos_title[27] on_d[27] vcc vout powertrain_cell
xu_pmos_title[26] on_d[26] vcc vout powertrain_cell
xu_pmos_title[25] on_d[25] vcc vout powertrain_cell
xu_pmos_title[24] on_d[24] vcc vout powertrain_cell
xu_pmos_title[23] on_d[23] vcc vout powertrain_cell
xu_pmos_title[22] on_d[22] vcc vout powertrain_cell
xu_pmos_title[21] on_d[21] vcc vout powertrain_cell
xu_pmos_title[20] on_d[20] vcc vout powertrain_cell
xu_pmos_title[19] on_d[19] vcc vout powertrain_cell
xu_pmos_title[18] on_d[18] vcc vout powertrain_cell
xu_pmos_title[17] on_d[17] vcc vout powertrain_cell
xu_pmos_title[16] on_d[16] vcc vout powertrain_cell
xu_pmos_title[15] on_d[15] vcc vout powertrain_cell
xu_pmos_title[14] on_d[14] vcc vout powertrain_cell
xu_pmos_title[13] on_d[13] vcc vout powertrain_cell
xu_pmos_title[12] on_d[12] vcc vout powertrain_cell
xu_pmos_title[11] on_d[11] vcc vout powertrain_cell
xu_pmos_title[10] on_d[10] vcc vout powertrain_cell
xu_pmos_title[9] on_d[9] vcc vout powertrain_cell
xu_pmos_title[8] on_d[8] vcc vout powertrain_cell
xu_pmos_title[7] on_d[7] vcc vout powertrain_cell
xu_pmos_title[6] on_d[6] vcc vout powertrain_cell
xu_pmos_title[5] on_d[5] vcc vout powertrain_cell
xu_pmos_title[4] on_d[4] vcc vout powertrain_cell
xu_pmos_title[3] on_d[3] vcc vout powertrain_cell
xu_pmos_title[2] on_d[2] vcc vout powertrain_cell
xu_pmos_title[1] on_d[1] vcc vout powertrain_cell
xu_pmos_title[0] on_d[0] vcc vout powertrain_cell
.ends


