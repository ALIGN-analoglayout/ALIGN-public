MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 11.84 BY 24.864 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 24.408 3.136 24.48 ;
      LAYER M2 ;
        RECT 3.084 24.428 3.156 24.46 ;
      LAYER M1 ;
        RECT 8.864 24.408 8.896 24.48 ;
      LAYER M2 ;
        RECT 8.844 24.428 8.916 24.46 ;
      LAYER M2 ;
        RECT 3.12 24.428 8.88 24.46 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
      LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.984 24.576 6.016 24.648 ;
      LAYER M2 ;
        RECT 5.964 24.596 6.036 24.628 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
      LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
      LAYER M1 ;
        RECT 8.704 0.216 8.736 0.288 ;
      LAYER M2 ;
        RECT 8.684 0.236 8.756 0.268 ;
      LAYER M2 ;
        RECT 2.96 0.236 8.72 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 5.664 9.708 5.696 9.78 ;
  LAYER M2 ;
        RECT 5.644 9.728 5.716 9.76 ;
  LAYER M1 ;
        RECT 5.664 9.576 5.696 9.744 ;
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M2 ;
        RECT 5.68 9.56 5.84 9.592 ;
  LAYER M1 ;
        RECT 5.824 9.54 5.856 9.612 ;
  LAYER M2 ;
        RECT 5.804 9.56 5.876 9.592 ;
  LAYER M1 ;
        RECT 8.544 12.648 8.576 12.72 ;
  LAYER M2 ;
        RECT 8.524 12.668 8.596 12.7 ;
  LAYER M2 ;
        RECT 5.84 12.668 8.56 12.7 ;
  LAYER M1 ;
        RECT 5.824 12.648 5.856 12.72 ;
  LAYER M2 ;
        RECT 5.804 12.668 5.876 12.7 ;
  LAYER M1 ;
        RECT 5.664 12.648 5.696 12.72 ;
  LAYER M2 ;
        RECT 5.644 12.668 5.716 12.7 ;
  LAYER M1 ;
        RECT 5.664 12.516 5.696 12.684 ;
  LAYER M1 ;
        RECT 5.664 12.48 5.696 12.552 ;
  LAYER M2 ;
        RECT 5.644 12.5 5.716 12.532 ;
  LAYER M2 ;
        RECT 5.68 12.5 5.84 12.532 ;
  LAYER M1 ;
        RECT 5.824 12.48 5.856 12.552 ;
  LAYER M2 ;
        RECT 5.804 12.5 5.876 12.532 ;
  LAYER M1 ;
        RECT 8.544 9.708 8.576 9.78 ;
  LAYER M2 ;
        RECT 8.524 9.728 8.596 9.76 ;
  LAYER M2 ;
        RECT 5.84 9.728 8.56 9.76 ;
  LAYER M1 ;
        RECT 5.824 9.708 5.856 9.78 ;
  LAYER M2 ;
        RECT 5.804 9.728 5.876 9.76 ;
  LAYER M1 ;
        RECT 5.664 15.588 5.696 15.66 ;
  LAYER M2 ;
        RECT 5.644 15.608 5.716 15.64 ;
  LAYER M1 ;
        RECT 5.664 15.456 5.696 15.624 ;
  LAYER M1 ;
        RECT 5.664 15.42 5.696 15.492 ;
  LAYER M2 ;
        RECT 5.644 15.44 5.716 15.472 ;
  LAYER M2 ;
        RECT 5.68 15.44 5.84 15.472 ;
  LAYER M1 ;
        RECT 5.824 15.42 5.856 15.492 ;
  LAYER M2 ;
        RECT 5.804 15.44 5.876 15.472 ;
  LAYER M1 ;
        RECT 8.544 6.768 8.576 6.84 ;
  LAYER M2 ;
        RECT 8.524 6.788 8.596 6.82 ;
  LAYER M2 ;
        RECT 5.84 6.788 8.56 6.82 ;
  LAYER M1 ;
        RECT 5.824 6.768 5.856 6.84 ;
  LAYER M2 ;
        RECT 5.804 6.788 5.876 6.82 ;
  LAYER M1 ;
        RECT 5.824 0.384 5.856 0.456 ;
  LAYER M2 ;
        RECT 5.804 0.404 5.876 0.436 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 0.588 ;
  LAYER M1 ;
        RECT 5.824 0.588 5.856 15.456 ;
  LAYER M1 ;
        RECT 5.664 6.768 5.696 6.84 ;
  LAYER M2 ;
        RECT 5.644 6.788 5.716 6.82 ;
  LAYER M2 ;
        RECT 2.96 6.788 5.68 6.82 ;
  LAYER M1 ;
        RECT 2.944 6.768 2.976 6.84 ;
  LAYER M2 ;
        RECT 2.924 6.788 2.996 6.82 ;
  LAYER M1 ;
        RECT 5.664 18.528 5.696 18.6 ;
  LAYER M2 ;
        RECT 5.644 18.548 5.716 18.58 ;
  LAYER M2 ;
        RECT 2.96 18.548 5.68 18.58 ;
  LAYER M1 ;
        RECT 2.944 18.528 2.976 18.6 ;
  LAYER M2 ;
        RECT 2.924 18.548 2.996 18.58 ;
  LAYER M1 ;
        RECT 5.664 3.828 5.696 3.9 ;
  LAYER M2 ;
        RECT 5.644 3.848 5.716 3.88 ;
  LAYER M2 ;
        RECT 2.96 3.848 5.68 3.88 ;
  LAYER M1 ;
        RECT 2.944 3.828 2.976 3.9 ;
  LAYER M2 ;
        RECT 2.924 3.848 2.996 3.88 ;
  LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
  LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
  LAYER M1 ;
        RECT 2.944 0.252 2.976 0.588 ;
  LAYER M1 ;
        RECT 2.944 0.588 2.976 18.564 ;
  LAYER M1 ;
        RECT 8.544 15.588 8.576 15.66 ;
  LAYER M2 ;
        RECT 8.524 15.608 8.596 15.64 ;
  LAYER M1 ;
        RECT 8.544 15.456 8.576 15.624 ;
  LAYER M1 ;
        RECT 8.544 15.42 8.576 15.492 ;
  LAYER M2 ;
        RECT 8.524 15.44 8.596 15.472 ;
  LAYER M2 ;
        RECT 8.56 15.44 8.72 15.472 ;
  LAYER M1 ;
        RECT 8.704 15.42 8.736 15.492 ;
  LAYER M2 ;
        RECT 8.684 15.44 8.756 15.472 ;
  LAYER M1 ;
        RECT 8.544 3.828 8.576 3.9 ;
  LAYER M2 ;
        RECT 8.524 3.848 8.596 3.88 ;
  LAYER M1 ;
        RECT 8.544 3.696 8.576 3.864 ;
  LAYER M1 ;
        RECT 8.544 3.66 8.576 3.732 ;
  LAYER M2 ;
        RECT 8.524 3.68 8.596 3.712 ;
  LAYER M2 ;
        RECT 8.56 3.68 8.72 3.712 ;
  LAYER M1 ;
        RECT 8.704 3.66 8.736 3.732 ;
  LAYER M2 ;
        RECT 8.684 3.68 8.756 3.712 ;
  LAYER M1 ;
        RECT 8.544 18.528 8.576 18.6 ;
  LAYER M2 ;
        RECT 8.524 18.548 8.596 18.58 ;
  LAYER M1 ;
        RECT 8.544 18.396 8.576 18.564 ;
  LAYER M1 ;
        RECT 8.544 18.36 8.576 18.432 ;
  LAYER M2 ;
        RECT 8.524 18.38 8.596 18.412 ;
  LAYER M2 ;
        RECT 8.56 18.38 8.72 18.412 ;
  LAYER M1 ;
        RECT 8.704 18.36 8.736 18.432 ;
  LAYER M2 ;
        RECT 8.684 18.38 8.756 18.412 ;
  LAYER M1 ;
        RECT 8.704 0.216 8.736 0.288 ;
  LAYER M2 ;
        RECT 8.684 0.236 8.756 0.268 ;
  LAYER M1 ;
        RECT 8.704 0.252 8.736 0.588 ;
  LAYER M1 ;
        RECT 8.704 0.588 8.736 18.396 ;
  LAYER M2 ;
        RECT 2.96 0.236 8.72 0.268 ;
  LAYER M1 ;
        RECT 2.784 0.888 2.816 0.96 ;
  LAYER M2 ;
        RECT 2.764 0.908 2.836 0.94 ;
  LAYER M2 ;
        RECT 0.08 0.908 2.8 0.94 ;
  LAYER M1 ;
        RECT 0.064 0.888 0.096 0.96 ;
  LAYER M2 ;
        RECT 0.044 0.908 0.116 0.94 ;
  LAYER M1 ;
        RECT 2.784 3.828 2.816 3.9 ;
  LAYER M2 ;
        RECT 2.764 3.848 2.836 3.88 ;
  LAYER M2 ;
        RECT 0.08 3.848 2.8 3.88 ;
  LAYER M1 ;
        RECT 0.064 3.828 0.096 3.9 ;
  LAYER M2 ;
        RECT 0.044 3.848 0.116 3.88 ;
  LAYER M1 ;
        RECT 2.784 6.768 2.816 6.84 ;
  LAYER M2 ;
        RECT 2.764 6.788 2.836 6.82 ;
  LAYER M2 ;
        RECT 0.08 6.788 2.8 6.82 ;
  LAYER M1 ;
        RECT 0.064 6.768 0.096 6.84 ;
  LAYER M2 ;
        RECT 0.044 6.788 0.116 6.82 ;
  LAYER M1 ;
        RECT 2.784 9.708 2.816 9.78 ;
  LAYER M2 ;
        RECT 2.764 9.728 2.836 9.76 ;
  LAYER M2 ;
        RECT 0.08 9.728 2.8 9.76 ;
  LAYER M1 ;
        RECT 0.064 9.708 0.096 9.78 ;
  LAYER M2 ;
        RECT 0.044 9.728 0.116 9.76 ;
  LAYER M1 ;
        RECT 2.784 12.648 2.816 12.72 ;
  LAYER M2 ;
        RECT 2.764 12.668 2.836 12.7 ;
  LAYER M2 ;
        RECT 0.08 12.668 2.8 12.7 ;
  LAYER M1 ;
        RECT 0.064 12.648 0.096 12.72 ;
  LAYER M2 ;
        RECT 0.044 12.668 0.116 12.7 ;
  LAYER M1 ;
        RECT 2.784 15.588 2.816 15.66 ;
  LAYER M2 ;
        RECT 2.764 15.608 2.836 15.64 ;
  LAYER M2 ;
        RECT 0.08 15.608 2.8 15.64 ;
  LAYER M1 ;
        RECT 0.064 15.588 0.096 15.66 ;
  LAYER M2 ;
        RECT 0.044 15.608 0.116 15.64 ;
  LAYER M1 ;
        RECT 2.784 18.528 2.816 18.6 ;
  LAYER M2 ;
        RECT 2.764 18.548 2.836 18.58 ;
  LAYER M2 ;
        RECT 0.08 18.548 2.8 18.58 ;
  LAYER M1 ;
        RECT 0.064 18.528 0.096 18.6 ;
  LAYER M2 ;
        RECT 0.044 18.548 0.116 18.58 ;
  LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
  LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
  LAYER M2 ;
        RECT 0.08 21.488 2.8 21.52 ;
  LAYER M1 ;
        RECT 0.064 21.468 0.096 21.54 ;
  LAYER M2 ;
        RECT 0.044 21.488 0.116 21.52 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.588 ;
  LAYER M1 ;
        RECT 0.064 0.588 0.096 21.504 ;
  LAYER M1 ;
        RECT 11.424 0.888 11.456 0.96 ;
  LAYER M2 ;
        RECT 11.404 0.908 11.476 0.94 ;
  LAYER M1 ;
        RECT 11.424 0.756 11.456 0.924 ;
  LAYER M1 ;
        RECT 11.424 0.72 11.456 0.792 ;
  LAYER M2 ;
        RECT 11.404 0.74 11.476 0.772 ;
  LAYER M2 ;
        RECT 11.44 0.74 11.6 0.772 ;
  LAYER M1 ;
        RECT 11.584 0.72 11.616 0.792 ;
  LAYER M2 ;
        RECT 11.564 0.74 11.636 0.772 ;
  LAYER M1 ;
        RECT 11.424 3.828 11.456 3.9 ;
  LAYER M2 ;
        RECT 11.404 3.848 11.476 3.88 ;
  LAYER M1 ;
        RECT 11.424 3.696 11.456 3.864 ;
  LAYER M1 ;
        RECT 11.424 3.66 11.456 3.732 ;
  LAYER M2 ;
        RECT 11.404 3.68 11.476 3.712 ;
  LAYER M2 ;
        RECT 11.44 3.68 11.6 3.712 ;
  LAYER M1 ;
        RECT 11.584 3.66 11.616 3.732 ;
  LAYER M2 ;
        RECT 11.564 3.68 11.636 3.712 ;
  LAYER M1 ;
        RECT 11.424 6.768 11.456 6.84 ;
  LAYER M2 ;
        RECT 11.404 6.788 11.476 6.82 ;
  LAYER M1 ;
        RECT 11.424 6.636 11.456 6.804 ;
  LAYER M1 ;
        RECT 11.424 6.6 11.456 6.672 ;
  LAYER M2 ;
        RECT 11.404 6.62 11.476 6.652 ;
  LAYER M2 ;
        RECT 11.44 6.62 11.6 6.652 ;
  LAYER M1 ;
        RECT 11.584 6.6 11.616 6.672 ;
  LAYER M2 ;
        RECT 11.564 6.62 11.636 6.652 ;
  LAYER M1 ;
        RECT 11.424 9.708 11.456 9.78 ;
  LAYER M2 ;
        RECT 11.404 9.728 11.476 9.76 ;
  LAYER M1 ;
        RECT 11.424 9.576 11.456 9.744 ;
  LAYER M1 ;
        RECT 11.424 9.54 11.456 9.612 ;
  LAYER M2 ;
        RECT 11.404 9.56 11.476 9.592 ;
  LAYER M2 ;
        RECT 11.44 9.56 11.6 9.592 ;
  LAYER M1 ;
        RECT 11.584 9.54 11.616 9.612 ;
  LAYER M2 ;
        RECT 11.564 9.56 11.636 9.592 ;
  LAYER M1 ;
        RECT 11.424 12.648 11.456 12.72 ;
  LAYER M2 ;
        RECT 11.404 12.668 11.476 12.7 ;
  LAYER M1 ;
        RECT 11.424 12.516 11.456 12.684 ;
  LAYER M1 ;
        RECT 11.424 12.48 11.456 12.552 ;
  LAYER M2 ;
        RECT 11.404 12.5 11.476 12.532 ;
  LAYER M2 ;
        RECT 11.44 12.5 11.6 12.532 ;
  LAYER M1 ;
        RECT 11.584 12.48 11.616 12.552 ;
  LAYER M2 ;
        RECT 11.564 12.5 11.636 12.532 ;
  LAYER M1 ;
        RECT 11.424 15.588 11.456 15.66 ;
  LAYER M2 ;
        RECT 11.404 15.608 11.476 15.64 ;
  LAYER M1 ;
        RECT 11.424 15.456 11.456 15.624 ;
  LAYER M1 ;
        RECT 11.424 15.42 11.456 15.492 ;
  LAYER M2 ;
        RECT 11.404 15.44 11.476 15.472 ;
  LAYER M2 ;
        RECT 11.44 15.44 11.6 15.472 ;
  LAYER M1 ;
        RECT 11.584 15.42 11.616 15.492 ;
  LAYER M2 ;
        RECT 11.564 15.44 11.636 15.472 ;
  LAYER M1 ;
        RECT 11.424 18.528 11.456 18.6 ;
  LAYER M2 ;
        RECT 11.404 18.548 11.476 18.58 ;
  LAYER M1 ;
        RECT 11.424 18.396 11.456 18.564 ;
  LAYER M1 ;
        RECT 11.424 18.36 11.456 18.432 ;
  LAYER M2 ;
        RECT 11.404 18.38 11.476 18.412 ;
  LAYER M2 ;
        RECT 11.44 18.38 11.6 18.412 ;
  LAYER M1 ;
        RECT 11.584 18.36 11.616 18.432 ;
  LAYER M2 ;
        RECT 11.564 18.38 11.636 18.412 ;
  LAYER M1 ;
        RECT 11.424 21.468 11.456 21.54 ;
  LAYER M2 ;
        RECT 11.404 21.488 11.476 21.52 ;
  LAYER M1 ;
        RECT 11.424 21.336 11.456 21.504 ;
  LAYER M1 ;
        RECT 11.424 21.3 11.456 21.372 ;
  LAYER M2 ;
        RECT 11.404 21.32 11.476 21.352 ;
  LAYER M2 ;
        RECT 11.44 21.32 11.6 21.352 ;
  LAYER M1 ;
        RECT 11.584 21.3 11.616 21.372 ;
  LAYER M2 ;
        RECT 11.564 21.32 11.636 21.352 ;
  LAYER M1 ;
        RECT 11.584 0.048 11.616 0.12 ;
  LAYER M2 ;
        RECT 11.564 0.068 11.636 0.1 ;
  LAYER M1 ;
        RECT 11.584 0.084 11.616 0.588 ;
  LAYER M1 ;
        RECT 11.584 0.588 11.616 21.336 ;
  LAYER M2 ;
        RECT 0.08 0.068 11.6 0.1 ;
  LAYER M1 ;
        RECT 5.664 0.888 5.696 0.96 ;
  LAYER M2 ;
        RECT 5.644 0.908 5.716 0.94 ;
  LAYER M2 ;
        RECT 2.8 0.908 5.68 0.94 ;
  LAYER M1 ;
        RECT 2.784 0.888 2.816 0.96 ;
  LAYER M2 ;
        RECT 2.764 0.908 2.836 0.94 ;
  LAYER M1 ;
        RECT 5.664 21.468 5.696 21.54 ;
  LAYER M2 ;
        RECT 5.644 21.488 5.716 21.52 ;
  LAYER M2 ;
        RECT 2.8 21.488 5.68 21.52 ;
  LAYER M1 ;
        RECT 2.784 21.468 2.816 21.54 ;
  LAYER M2 ;
        RECT 2.764 21.488 2.836 21.52 ;
  LAYER M1 ;
        RECT 8.544 21.468 8.576 21.54 ;
  LAYER M2 ;
        RECT 8.524 21.488 8.596 21.52 ;
  LAYER M2 ;
        RECT 5.68 21.488 8.56 21.52 ;
  LAYER M1 ;
        RECT 5.664 21.468 5.696 21.54 ;
  LAYER M2 ;
        RECT 5.644 21.488 5.716 21.52 ;
  LAYER M1 ;
        RECT 8.544 0.888 8.576 0.96 ;
  LAYER M2 ;
        RECT 8.524 0.908 8.596 0.94 ;
  LAYER M2 ;
        RECT 8.56 0.908 11.44 0.94 ;
  LAYER M1 ;
        RECT 11.424 0.888 11.456 0.96 ;
  LAYER M2 ;
        RECT 11.404 0.908 11.476 0.94 ;
  LAYER M1 ;
        RECT 3.264 12.144 3.296 12.216 ;
  LAYER M2 ;
        RECT 3.244 12.164 3.316 12.196 ;
  LAYER M2 ;
        RECT 3.12 12.164 3.28 12.196 ;
  LAYER M1 ;
        RECT 3.104 12.144 3.136 12.216 ;
  LAYER M2 ;
        RECT 3.084 12.164 3.156 12.196 ;
  LAYER M1 ;
        RECT 3.264 15.084 3.296 15.156 ;
  LAYER M2 ;
        RECT 3.244 15.104 3.316 15.136 ;
  LAYER M2 ;
        RECT 3.12 15.104 3.28 15.136 ;
  LAYER M1 ;
        RECT 3.104 15.084 3.136 15.156 ;
  LAYER M2 ;
        RECT 3.084 15.104 3.156 15.136 ;
  LAYER M1 ;
        RECT 3.264 18.024 3.296 18.096 ;
  LAYER M2 ;
        RECT 3.244 18.044 3.316 18.076 ;
  LAYER M2 ;
        RECT 3.12 18.044 3.28 18.076 ;
  LAYER M1 ;
        RECT 3.104 18.024 3.136 18.096 ;
  LAYER M2 ;
        RECT 3.084 18.044 3.156 18.076 ;
  LAYER M1 ;
        RECT 3.104 24.408 3.136 24.48 ;
  LAYER M2 ;
        RECT 3.084 24.428 3.156 24.46 ;
  LAYER M1 ;
        RECT 3.104 24.276 3.136 24.444 ;
  LAYER M1 ;
        RECT 3.104 12.18 3.136 24.276 ;
  LAYER M1 ;
        RECT 6.144 15.084 6.176 15.156 ;
  LAYER M2 ;
        RECT 6.124 15.104 6.196 15.136 ;
  LAYER M1 ;
        RECT 6.144 15.12 6.176 15.288 ;
  LAYER M1 ;
        RECT 6.144 15.252 6.176 15.324 ;
  LAYER M2 ;
        RECT 6.124 15.272 6.196 15.304 ;
  LAYER M2 ;
        RECT 6.16 15.272 8.88 15.304 ;
  LAYER M1 ;
        RECT 8.864 15.252 8.896 15.324 ;
  LAYER M2 ;
        RECT 8.844 15.272 8.916 15.304 ;
  LAYER M1 ;
        RECT 6.144 12.144 6.176 12.216 ;
  LAYER M2 ;
        RECT 6.124 12.164 6.196 12.196 ;
  LAYER M1 ;
        RECT 6.144 12.18 6.176 12.348 ;
  LAYER M1 ;
        RECT 6.144 12.312 6.176 12.384 ;
  LAYER M2 ;
        RECT 6.124 12.332 6.196 12.364 ;
  LAYER M2 ;
        RECT 6.16 12.332 8.88 12.364 ;
  LAYER M1 ;
        RECT 8.864 12.312 8.896 12.384 ;
  LAYER M2 ;
        RECT 8.844 12.332 8.916 12.364 ;
  LAYER M1 ;
        RECT 6.144 9.204 6.176 9.276 ;
  LAYER M2 ;
        RECT 6.124 9.224 6.196 9.256 ;
  LAYER M1 ;
        RECT 6.144 9.24 6.176 9.408 ;
  LAYER M1 ;
        RECT 6.144 9.372 6.176 9.444 ;
  LAYER M2 ;
        RECT 6.124 9.392 6.196 9.424 ;
  LAYER M2 ;
        RECT 6.16 9.392 8.88 9.424 ;
  LAYER M1 ;
        RECT 8.864 9.372 8.896 9.444 ;
  LAYER M2 ;
        RECT 8.844 9.392 8.916 9.424 ;
  LAYER M1 ;
        RECT 8.864 24.408 8.896 24.48 ;
  LAYER M2 ;
        RECT 8.844 24.428 8.916 24.46 ;
  LAYER M1 ;
        RECT 8.864 24.276 8.896 24.444 ;
  LAYER M1 ;
        RECT 8.864 9.408 8.896 24.276 ;
  LAYER M2 ;
        RECT 3.12 24.428 8.88 24.46 ;
  LAYER M1 ;
        RECT 3.264 9.204 3.296 9.276 ;
  LAYER M2 ;
        RECT 3.244 9.224 3.316 9.256 ;
  LAYER M1 ;
        RECT 3.264 9.24 3.296 9.408 ;
  LAYER M1 ;
        RECT 3.264 9.372 3.296 9.444 ;
  LAYER M2 ;
        RECT 3.244 9.392 3.316 9.424 ;
  LAYER M2 ;
        RECT 3.28 9.392 6 9.424 ;
  LAYER M1 ;
        RECT 5.984 9.372 6.016 9.444 ;
  LAYER M2 ;
        RECT 5.964 9.392 6.036 9.424 ;
  LAYER M1 ;
        RECT 6.144 18.024 6.176 18.096 ;
  LAYER M2 ;
        RECT 6.124 18.044 6.196 18.076 ;
  LAYER M2 ;
        RECT 6 18.044 6.16 18.076 ;
  LAYER M1 ;
        RECT 5.984 18.024 6.016 18.096 ;
  LAYER M2 ;
        RECT 5.964 18.044 6.036 18.076 ;
  LAYER M1 ;
        RECT 3.264 20.964 3.296 21.036 ;
  LAYER M2 ;
        RECT 3.244 20.984 3.316 21.016 ;
  LAYER M1 ;
        RECT 3.264 21 3.296 21.168 ;
  LAYER M1 ;
        RECT 3.264 21.132 3.296 21.204 ;
  LAYER M2 ;
        RECT 3.244 21.152 3.316 21.184 ;
  LAYER M2 ;
        RECT 3.28 21.152 6 21.184 ;
  LAYER M1 ;
        RECT 5.984 21.132 6.016 21.204 ;
  LAYER M2 ;
        RECT 5.964 21.152 6.036 21.184 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M2 ;
        RECT 6 6.284 6.16 6.316 ;
  LAYER M1 ;
        RECT 5.984 6.264 6.016 6.336 ;
  LAYER M2 ;
        RECT 5.964 6.284 6.036 6.316 ;
  LAYER M1 ;
        RECT 3.264 6.264 3.296 6.336 ;
  LAYER M2 ;
        RECT 3.244 6.284 3.316 6.316 ;
  LAYER M1 ;
        RECT 3.264 6.3 3.296 6.468 ;
  LAYER M1 ;
        RECT 3.264 6.432 3.296 6.504 ;
  LAYER M2 ;
        RECT 3.244 6.452 3.316 6.484 ;
  LAYER M2 ;
        RECT 3.28 6.452 6 6.484 ;
  LAYER M1 ;
        RECT 5.984 6.432 6.016 6.504 ;
  LAYER M2 ;
        RECT 5.964 6.452 6.036 6.484 ;
  LAYER M1 ;
        RECT 6.144 20.964 6.176 21.036 ;
  LAYER M2 ;
        RECT 6.124 20.984 6.196 21.016 ;
  LAYER M2 ;
        RECT 6 20.984 6.16 21.016 ;
  LAYER M1 ;
        RECT 5.984 20.964 6.016 21.036 ;
  LAYER M2 ;
        RECT 5.964 20.984 6.036 21.016 ;
  LAYER M1 ;
        RECT 5.984 24.576 6.016 24.648 ;
  LAYER M2 ;
        RECT 5.964 24.596 6.036 24.628 ;
  LAYER M1 ;
        RECT 5.984 24.276 6.016 24.612 ;
  LAYER M1 ;
        RECT 5.984 6.3 6.016 24.276 ;
  LAYER M1 ;
        RECT 0.384 3.324 0.416 3.396 ;
  LAYER M2 ;
        RECT 0.364 3.344 0.436 3.376 ;
  LAYER M2 ;
        RECT 0.24 3.344 0.4 3.376 ;
  LAYER M1 ;
        RECT 0.224 3.324 0.256 3.396 ;
  LAYER M2 ;
        RECT 0.204 3.344 0.276 3.376 ;
  LAYER M1 ;
        RECT 0.384 6.264 0.416 6.336 ;
  LAYER M2 ;
        RECT 0.364 6.284 0.436 6.316 ;
  LAYER M2 ;
        RECT 0.24 6.284 0.4 6.316 ;
  LAYER M1 ;
        RECT 0.224 6.264 0.256 6.336 ;
  LAYER M2 ;
        RECT 0.204 6.284 0.276 6.316 ;
  LAYER M1 ;
        RECT 0.384 9.204 0.416 9.276 ;
  LAYER M2 ;
        RECT 0.364 9.224 0.436 9.256 ;
  LAYER M2 ;
        RECT 0.24 9.224 0.4 9.256 ;
  LAYER M1 ;
        RECT 0.224 9.204 0.256 9.276 ;
  LAYER M2 ;
        RECT 0.204 9.224 0.276 9.256 ;
  LAYER M1 ;
        RECT 0.384 12.144 0.416 12.216 ;
  LAYER M2 ;
        RECT 0.364 12.164 0.436 12.196 ;
  LAYER M2 ;
        RECT 0.24 12.164 0.4 12.196 ;
  LAYER M1 ;
        RECT 0.224 12.144 0.256 12.216 ;
  LAYER M2 ;
        RECT 0.204 12.164 0.276 12.196 ;
  LAYER M1 ;
        RECT 0.384 15.084 0.416 15.156 ;
  LAYER M2 ;
        RECT 0.364 15.104 0.436 15.136 ;
  LAYER M2 ;
        RECT 0.24 15.104 0.4 15.136 ;
  LAYER M1 ;
        RECT 0.224 15.084 0.256 15.156 ;
  LAYER M2 ;
        RECT 0.204 15.104 0.276 15.136 ;
  LAYER M1 ;
        RECT 0.384 18.024 0.416 18.096 ;
  LAYER M2 ;
        RECT 0.364 18.044 0.436 18.076 ;
  LAYER M2 ;
        RECT 0.24 18.044 0.4 18.076 ;
  LAYER M1 ;
        RECT 0.224 18.024 0.256 18.096 ;
  LAYER M2 ;
        RECT 0.204 18.044 0.276 18.076 ;
  LAYER M1 ;
        RECT 0.384 20.964 0.416 21.036 ;
  LAYER M2 ;
        RECT 0.364 20.984 0.436 21.016 ;
  LAYER M2 ;
        RECT 0.24 20.984 0.4 21.016 ;
  LAYER M1 ;
        RECT 0.224 20.964 0.256 21.036 ;
  LAYER M2 ;
        RECT 0.204 20.984 0.276 21.016 ;
  LAYER M1 ;
        RECT 0.384 23.904 0.416 23.976 ;
  LAYER M2 ;
        RECT 0.364 23.924 0.436 23.956 ;
  LAYER M2 ;
        RECT 0.24 23.924 0.4 23.956 ;
  LAYER M1 ;
        RECT 0.224 23.904 0.256 23.976 ;
  LAYER M2 ;
        RECT 0.204 23.924 0.276 23.956 ;
  LAYER M1 ;
        RECT 0.224 24.744 0.256 24.816 ;
  LAYER M2 ;
        RECT 0.204 24.764 0.276 24.796 ;
  LAYER M1 ;
        RECT 0.224 24.276 0.256 24.78 ;
  LAYER M1 ;
        RECT 0.224 3.36 0.256 24.276 ;
  LAYER M1 ;
        RECT 9.024 3.324 9.056 3.396 ;
  LAYER M2 ;
        RECT 9.004 3.344 9.076 3.376 ;
  LAYER M1 ;
        RECT 9.024 3.36 9.056 3.528 ;
  LAYER M1 ;
        RECT 9.024 3.492 9.056 3.564 ;
  LAYER M2 ;
        RECT 9.004 3.512 9.076 3.544 ;
  LAYER M2 ;
        RECT 9.04 3.512 11.76 3.544 ;
  LAYER M1 ;
        RECT 11.744 3.492 11.776 3.564 ;
  LAYER M2 ;
        RECT 11.724 3.512 11.796 3.544 ;
  LAYER M1 ;
        RECT 9.024 6.264 9.056 6.336 ;
  LAYER M2 ;
        RECT 9.004 6.284 9.076 6.316 ;
  LAYER M1 ;
        RECT 9.024 6.3 9.056 6.468 ;
  LAYER M1 ;
        RECT 9.024 6.432 9.056 6.504 ;
  LAYER M2 ;
        RECT 9.004 6.452 9.076 6.484 ;
  LAYER M2 ;
        RECT 9.04 6.452 11.76 6.484 ;
  LAYER M1 ;
        RECT 11.744 6.432 11.776 6.504 ;
  LAYER M2 ;
        RECT 11.724 6.452 11.796 6.484 ;
  LAYER M1 ;
        RECT 9.024 9.204 9.056 9.276 ;
  LAYER M2 ;
        RECT 9.004 9.224 9.076 9.256 ;
  LAYER M1 ;
        RECT 9.024 9.24 9.056 9.408 ;
  LAYER M1 ;
        RECT 9.024 9.372 9.056 9.444 ;
  LAYER M2 ;
        RECT 9.004 9.392 9.076 9.424 ;
  LAYER M2 ;
        RECT 9.04 9.392 11.76 9.424 ;
  LAYER M1 ;
        RECT 11.744 9.372 11.776 9.444 ;
  LAYER M2 ;
        RECT 11.724 9.392 11.796 9.424 ;
  LAYER M1 ;
        RECT 9.024 12.144 9.056 12.216 ;
  LAYER M2 ;
        RECT 9.004 12.164 9.076 12.196 ;
  LAYER M1 ;
        RECT 9.024 12.18 9.056 12.348 ;
  LAYER M1 ;
        RECT 9.024 12.312 9.056 12.384 ;
  LAYER M2 ;
        RECT 9.004 12.332 9.076 12.364 ;
  LAYER M2 ;
        RECT 9.04 12.332 11.76 12.364 ;
  LAYER M1 ;
        RECT 11.744 12.312 11.776 12.384 ;
  LAYER M2 ;
        RECT 11.724 12.332 11.796 12.364 ;
  LAYER M1 ;
        RECT 9.024 15.084 9.056 15.156 ;
  LAYER M2 ;
        RECT 9.004 15.104 9.076 15.136 ;
  LAYER M1 ;
        RECT 9.024 15.12 9.056 15.288 ;
  LAYER M1 ;
        RECT 9.024 15.252 9.056 15.324 ;
  LAYER M2 ;
        RECT 9.004 15.272 9.076 15.304 ;
  LAYER M2 ;
        RECT 9.04 15.272 11.76 15.304 ;
  LAYER M1 ;
        RECT 11.744 15.252 11.776 15.324 ;
  LAYER M2 ;
        RECT 11.724 15.272 11.796 15.304 ;
  LAYER M1 ;
        RECT 9.024 18.024 9.056 18.096 ;
  LAYER M2 ;
        RECT 9.004 18.044 9.076 18.076 ;
  LAYER M1 ;
        RECT 9.024 18.06 9.056 18.228 ;
  LAYER M1 ;
        RECT 9.024 18.192 9.056 18.264 ;
  LAYER M2 ;
        RECT 9.004 18.212 9.076 18.244 ;
  LAYER M2 ;
        RECT 9.04 18.212 11.76 18.244 ;
  LAYER M1 ;
        RECT 11.744 18.192 11.776 18.264 ;
  LAYER M2 ;
        RECT 11.724 18.212 11.796 18.244 ;
  LAYER M1 ;
        RECT 9.024 20.964 9.056 21.036 ;
  LAYER M2 ;
        RECT 9.004 20.984 9.076 21.016 ;
  LAYER M1 ;
        RECT 9.024 21 9.056 21.168 ;
  LAYER M1 ;
        RECT 9.024 21.132 9.056 21.204 ;
  LAYER M2 ;
        RECT 9.004 21.152 9.076 21.184 ;
  LAYER M2 ;
        RECT 9.04 21.152 11.76 21.184 ;
  LAYER M1 ;
        RECT 11.744 21.132 11.776 21.204 ;
  LAYER M2 ;
        RECT 11.724 21.152 11.796 21.184 ;
  LAYER M1 ;
        RECT 9.024 23.904 9.056 23.976 ;
  LAYER M2 ;
        RECT 9.004 23.924 9.076 23.956 ;
  LAYER M1 ;
        RECT 9.024 23.94 9.056 24.108 ;
  LAYER M1 ;
        RECT 9.024 24.072 9.056 24.144 ;
  LAYER M2 ;
        RECT 9.004 24.092 9.076 24.124 ;
  LAYER M2 ;
        RECT 9.04 24.092 11.76 24.124 ;
  LAYER M1 ;
        RECT 11.744 24.072 11.776 24.144 ;
  LAYER M2 ;
        RECT 11.724 24.092 11.796 24.124 ;
  LAYER M1 ;
        RECT 11.744 24.744 11.776 24.816 ;
  LAYER M2 ;
        RECT 11.724 24.764 11.796 24.796 ;
  LAYER M1 ;
        RECT 11.744 24.276 11.776 24.78 ;
  LAYER M1 ;
        RECT 11.744 3.528 11.776 24.276 ;
  LAYER M2 ;
        RECT 0.24 24.764 11.76 24.796 ;
  LAYER M1 ;
        RECT 3.264 3.324 3.296 3.396 ;
  LAYER M2 ;
        RECT 3.244 3.344 3.316 3.376 ;
  LAYER M2 ;
        RECT 0.4 3.344 3.28 3.376 ;
  LAYER M1 ;
        RECT 0.384 3.324 0.416 3.396 ;
  LAYER M2 ;
        RECT 0.364 3.344 0.436 3.376 ;
  LAYER M1 ;
        RECT 3.264 23.904 3.296 23.976 ;
  LAYER M2 ;
        RECT 3.244 23.924 3.316 23.956 ;
  LAYER M2 ;
        RECT 0.4 23.924 3.28 23.956 ;
  LAYER M1 ;
        RECT 0.384 23.904 0.416 23.976 ;
  LAYER M2 ;
        RECT 0.364 23.924 0.436 23.956 ;
  LAYER M1 ;
        RECT 6.144 23.904 6.176 23.976 ;
  LAYER M2 ;
        RECT 6.124 23.924 6.196 23.956 ;
  LAYER M2 ;
        RECT 3.28 23.924 6.16 23.956 ;
  LAYER M1 ;
        RECT 3.264 23.904 3.296 23.976 ;
  LAYER M2 ;
        RECT 3.244 23.924 3.316 23.956 ;
  LAYER M1 ;
        RECT 6.144 3.324 6.176 3.396 ;
  LAYER M2 ;
        RECT 6.124 3.344 6.196 3.376 ;
  LAYER M2 ;
        RECT 6.16 3.344 9.04 3.376 ;
  LAYER M1 ;
        RECT 9.024 3.324 9.056 3.396 ;
  LAYER M2 ;
        RECT 9.004 3.344 9.076 3.376 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.8 3.36 ;
  LAYER M1 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M3 ;
        RECT 0.4 3.864 2.8 6.3 ;
  LAYER M1 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M2 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M3 ;
        RECT 0.4 6.804 2.8 9.24 ;
  LAYER M1 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M2 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M3 ;
        RECT 0.4 9.744 2.8 12.18 ;
  LAYER M1 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M2 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M3 ;
        RECT 0.4 12.684 2.8 15.12 ;
  LAYER M1 ;
        RECT 0.4 15.624 2.8 18.06 ;
  LAYER M2 ;
        RECT 0.4 15.624 2.8 18.06 ;
  LAYER M3 ;
        RECT 0.4 15.624 2.8 18.06 ;
  LAYER M1 ;
        RECT 0.4 18.564 2.8 21 ;
  LAYER M2 ;
        RECT 0.4 18.564 2.8 21 ;
  LAYER M3 ;
        RECT 0.4 18.564 2.8 21 ;
  LAYER M1 ;
        RECT 0.4 21.504 2.8 23.94 ;
  LAYER M2 ;
        RECT 0.4 21.504 2.8 23.94 ;
  LAYER M3 ;
        RECT 0.4 21.504 2.8 23.94 ;
  LAYER M1 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M2 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M3 ;
        RECT 3.28 0.924 5.68 3.36 ;
  LAYER M1 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M2 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M3 ;
        RECT 3.28 3.864 5.68 6.3 ;
  LAYER M1 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M2 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M3 ;
        RECT 3.28 6.804 5.68 9.24 ;
  LAYER M1 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M2 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M3 ;
        RECT 3.28 9.744 5.68 12.18 ;
  LAYER M1 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M2 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M3 ;
        RECT 3.28 12.684 5.68 15.12 ;
  LAYER M1 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M2 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M3 ;
        RECT 3.28 15.624 5.68 18.06 ;
  LAYER M1 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M2 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M3 ;
        RECT 3.28 18.564 5.68 21 ;
  LAYER M1 ;
        RECT 3.28 21.504 5.68 23.94 ;
  LAYER M2 ;
        RECT 3.28 21.504 5.68 23.94 ;
  LAYER M3 ;
        RECT 3.28 21.504 5.68 23.94 ;
  LAYER M1 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M2 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M3 ;
        RECT 6.16 0.924 8.56 3.36 ;
  LAYER M1 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M2 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M3 ;
        RECT 6.16 3.864 8.56 6.3 ;
  LAYER M1 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M2 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M3 ;
        RECT 6.16 6.804 8.56 9.24 ;
  LAYER M1 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M2 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M3 ;
        RECT 6.16 9.744 8.56 12.18 ;
  LAYER M1 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M2 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M3 ;
        RECT 6.16 12.684 8.56 15.12 ;
  LAYER M1 ;
        RECT 6.16 15.624 8.56 18.06 ;
  LAYER M2 ;
        RECT 6.16 15.624 8.56 18.06 ;
  LAYER M3 ;
        RECT 6.16 15.624 8.56 18.06 ;
  LAYER M1 ;
        RECT 6.16 18.564 8.56 21 ;
  LAYER M2 ;
        RECT 6.16 18.564 8.56 21 ;
  LAYER M3 ;
        RECT 6.16 18.564 8.56 21 ;
  LAYER M1 ;
        RECT 6.16 21.504 8.56 23.94 ;
  LAYER M2 ;
        RECT 6.16 21.504 8.56 23.94 ;
  LAYER M3 ;
        RECT 6.16 21.504 8.56 23.94 ;
  LAYER M1 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M2 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M3 ;
        RECT 9.04 0.924 11.44 3.36 ;
  LAYER M1 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M2 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M3 ;
        RECT 9.04 3.864 11.44 6.3 ;
  LAYER M1 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M2 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M3 ;
        RECT 9.04 6.804 11.44 9.24 ;
  LAYER M1 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M2 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M3 ;
        RECT 9.04 9.744 11.44 12.18 ;
  LAYER M1 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M2 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M3 ;
        RECT 9.04 12.684 11.44 15.12 ;
  LAYER M1 ;
        RECT 9.04 15.624 11.44 18.06 ;
  LAYER M2 ;
        RECT 9.04 15.624 11.44 18.06 ;
  LAYER M3 ;
        RECT 9.04 15.624 11.44 18.06 ;
  LAYER M1 ;
        RECT 9.04 18.564 11.44 21 ;
  LAYER M2 ;
        RECT 9.04 18.564 11.44 21 ;
  LAYER M3 ;
        RECT 9.04 18.564 11.44 21 ;
  LAYER M1 ;
        RECT 9.04 21.504 11.44 23.94 ;
  LAYER M2 ;
        RECT 9.04 21.504 11.44 23.94 ;
  LAYER M3 ;
        RECT 9.04 21.504 11.44 23.94 ;
  END 
END Cap_60fF_Cap_60fF
