MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 12 BY 16.548 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 16.26 3.232 16.332 ;
      LAYER M2 ;
        RECT 3.18 16.28 3.252 16.312 ;
      LAYER M1 ;
        RECT 9.152 16.26 9.184 16.332 ;
      LAYER M2 ;
        RECT 9.132 16.28 9.204 16.312 ;
      LAYER M2 ;
        RECT 3.216 16.28 9.168 16.312 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
      LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.792 7.02 5.824 7.092 ;
  LAYER M2 ;
        RECT 5.772 7.04 5.844 7.072 ;
  LAYER M1 ;
        RECT 5.792 6.888 5.824 7.056 ;
  LAYER M1 ;
        RECT 5.792 6.852 5.824 6.924 ;
  LAYER M2 ;
        RECT 5.772 6.872 5.844 6.904 ;
  LAYER M2 ;
        RECT 5.808 6.872 6.032 6.904 ;
  LAYER M1 ;
        RECT 6.016 6.852 6.048 6.924 ;
  LAYER M2 ;
        RECT 5.996 6.872 6.068 6.904 ;
  LAYER M1 ;
        RECT 8.768 7.02 8.8 7.092 ;
  LAYER M2 ;
        RECT 8.748 7.04 8.82 7.072 ;
  LAYER M2 ;
        RECT 6.032 7.04 8.784 7.072 ;
  LAYER M1 ;
        RECT 6.016 7.02 6.048 7.092 ;
  LAYER M2 ;
        RECT 5.996 7.04 6.068 7.072 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M1 ;
        RECT 5.792 9.996 5.824 10.164 ;
  LAYER M1 ;
        RECT 5.792 9.96 5.824 10.032 ;
  LAYER M2 ;
        RECT 5.772 9.98 5.844 10.012 ;
  LAYER M2 ;
        RECT 5.808 9.98 6.032 10.012 ;
  LAYER M1 ;
        RECT 6.016 9.96 6.048 10.032 ;
  LAYER M2 ;
        RECT 5.996 9.98 6.068 10.012 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 6.032 3.932 8.784 3.964 ;
  LAYER M1 ;
        RECT 6.016 3.912 6.048 3.984 ;
  LAYER M2 ;
        RECT 5.996 3.932 6.068 3.964 ;
  LAYER M1 ;
        RECT 5.792 3.912 5.824 3.984 ;
  LAYER M2 ;
        RECT 5.772 3.932 5.844 3.964 ;
  LAYER M1 ;
        RECT 5.792 3.78 5.824 3.948 ;
  LAYER M1 ;
        RECT 5.792 3.744 5.824 3.816 ;
  LAYER M2 ;
        RECT 5.772 3.764 5.844 3.796 ;
  LAYER M2 ;
        RECT 5.808 3.764 6.032 3.796 ;
  LAYER M1 ;
        RECT 6.016 3.744 6.048 3.816 ;
  LAYER M2 ;
        RECT 5.996 3.764 6.068 3.796 ;
  LAYER M1 ;
        RECT 8.768 10.128 8.8 10.2 ;
  LAYER M2 ;
        RECT 8.748 10.148 8.82 10.18 ;
  LAYER M2 ;
        RECT 6.032 10.148 8.784 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 6.016 0.216 6.048 0.288 ;
  LAYER M2 ;
        RECT 5.996 0.236 6.068 0.268 ;
  LAYER M1 ;
        RECT 6.016 0.252 6.048 0.504 ;
  LAYER M1 ;
        RECT 6.016 0.504 6.048 10.164 ;
  LAYER M1 ;
        RECT 2.816 0.804 2.848 0.876 ;
  LAYER M2 ;
        RECT 2.796 0.824 2.868 0.856 ;
  LAYER M1 ;
        RECT 2.816 0.672 2.848 0.84 ;
  LAYER M1 ;
        RECT 2.816 0.636 2.848 0.708 ;
  LAYER M2 ;
        RECT 2.796 0.656 2.868 0.688 ;
  LAYER M2 ;
        RECT 2.832 0.656 3.056 0.688 ;
  LAYER M1 ;
        RECT 3.04 0.636 3.072 0.708 ;
  LAYER M2 ;
        RECT 3.02 0.656 3.092 0.688 ;
  LAYER M1 ;
        RECT 2.816 3.912 2.848 3.984 ;
  LAYER M2 ;
        RECT 2.796 3.932 2.868 3.964 ;
  LAYER M1 ;
        RECT 2.816 3.78 2.848 3.948 ;
  LAYER M1 ;
        RECT 2.816 3.744 2.848 3.816 ;
  LAYER M2 ;
        RECT 2.796 3.764 2.868 3.796 ;
  LAYER M2 ;
        RECT 2.832 3.764 3.056 3.796 ;
  LAYER M1 ;
        RECT 3.04 3.744 3.072 3.816 ;
  LAYER M2 ;
        RECT 3.02 3.764 3.092 3.796 ;
  LAYER M1 ;
        RECT 2.816 7.02 2.848 7.092 ;
  LAYER M2 ;
        RECT 2.796 7.04 2.868 7.072 ;
  LAYER M1 ;
        RECT 2.816 6.888 2.848 7.056 ;
  LAYER M1 ;
        RECT 2.816 6.852 2.848 6.924 ;
  LAYER M2 ;
        RECT 2.796 6.872 2.868 6.904 ;
  LAYER M2 ;
        RECT 2.832 6.872 3.056 6.904 ;
  LAYER M1 ;
        RECT 3.04 6.852 3.072 6.924 ;
  LAYER M2 ;
        RECT 3.02 6.872 3.092 6.904 ;
  LAYER M1 ;
        RECT 2.816 10.128 2.848 10.2 ;
  LAYER M2 ;
        RECT 2.796 10.148 2.868 10.18 ;
  LAYER M1 ;
        RECT 2.816 9.996 2.848 10.164 ;
  LAYER M1 ;
        RECT 2.816 9.96 2.848 10.032 ;
  LAYER M2 ;
        RECT 2.796 9.98 2.868 10.012 ;
  LAYER M2 ;
        RECT 2.832 9.98 3.056 10.012 ;
  LAYER M1 ;
        RECT 3.04 9.96 3.072 10.032 ;
  LAYER M2 ;
        RECT 3.02 9.98 3.092 10.012 ;
  LAYER M1 ;
        RECT 2.816 13.236 2.848 13.308 ;
  LAYER M2 ;
        RECT 2.796 13.256 2.868 13.288 ;
  LAYER M1 ;
        RECT 2.816 13.104 2.848 13.272 ;
  LAYER M1 ;
        RECT 2.816 13.068 2.848 13.14 ;
  LAYER M2 ;
        RECT 2.796 13.088 2.868 13.12 ;
  LAYER M2 ;
        RECT 2.832 13.088 3.056 13.12 ;
  LAYER M1 ;
        RECT 3.04 13.068 3.072 13.14 ;
  LAYER M2 ;
        RECT 3.02 13.088 3.092 13.12 ;
  LAYER M1 ;
        RECT 5.792 0.804 5.824 0.876 ;
  LAYER M2 ;
        RECT 5.772 0.824 5.844 0.856 ;
  LAYER M2 ;
        RECT 3.056 0.824 5.808 0.856 ;
  LAYER M1 ;
        RECT 3.04 0.804 3.072 0.876 ;
  LAYER M2 ;
        RECT 3.02 0.824 3.092 0.856 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M2 ;
        RECT 3.056 13.256 5.808 13.288 ;
  LAYER M1 ;
        RECT 3.04 13.236 3.072 13.308 ;
  LAYER M2 ;
        RECT 3.02 13.256 3.092 13.288 ;
  LAYER M1 ;
        RECT 3.04 0.048 3.072 0.12 ;
  LAYER M2 ;
        RECT 3.02 0.068 3.092 0.1 ;
  LAYER M1 ;
        RECT 3.04 0.084 3.072 0.504 ;
  LAYER M1 ;
        RECT 3.04 0.504 3.072 13.272 ;
  LAYER M1 ;
        RECT 8.768 0.804 8.8 0.876 ;
  LAYER M2 ;
        RECT 8.748 0.824 8.82 0.856 ;
  LAYER M1 ;
        RECT 8.768 0.672 8.8 0.84 ;
  LAYER M1 ;
        RECT 8.768 0.636 8.8 0.708 ;
  LAYER M2 ;
        RECT 8.748 0.656 8.82 0.688 ;
  LAYER M2 ;
        RECT 8.784 0.656 9.008 0.688 ;
  LAYER M1 ;
        RECT 8.992 0.636 9.024 0.708 ;
  LAYER M2 ;
        RECT 8.972 0.656 9.044 0.688 ;
  LAYER M1 ;
        RECT 8.768 13.236 8.8 13.308 ;
  LAYER M2 ;
        RECT 8.748 13.256 8.82 13.288 ;
  LAYER M1 ;
        RECT 8.768 13.104 8.8 13.272 ;
  LAYER M1 ;
        RECT 8.768 13.068 8.8 13.14 ;
  LAYER M2 ;
        RECT 8.748 13.088 8.82 13.12 ;
  LAYER M2 ;
        RECT 8.784 13.088 9.008 13.12 ;
  LAYER M1 ;
        RECT 8.992 13.068 9.024 13.14 ;
  LAYER M2 ;
        RECT 8.972 13.088 9.044 13.12 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M2 ;
        RECT 9.008 0.824 11.76 0.856 ;
  LAYER M1 ;
        RECT 8.992 0.804 9.024 0.876 ;
  LAYER M2 ;
        RECT 8.972 0.824 9.044 0.856 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 9.008 3.932 11.76 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 11.744 7.02 11.776 7.092 ;
  LAYER M2 ;
        RECT 11.724 7.04 11.796 7.072 ;
  LAYER M2 ;
        RECT 9.008 7.04 11.76 7.072 ;
  LAYER M1 ;
        RECT 8.992 7.02 9.024 7.092 ;
  LAYER M2 ;
        RECT 8.972 7.04 9.044 7.072 ;
  LAYER M1 ;
        RECT 11.744 10.128 11.776 10.2 ;
  LAYER M2 ;
        RECT 11.724 10.148 11.796 10.18 ;
  LAYER M2 ;
        RECT 9.008 10.148 11.76 10.18 ;
  LAYER M1 ;
        RECT 8.992 10.128 9.024 10.2 ;
  LAYER M2 ;
        RECT 8.972 10.148 9.044 10.18 ;
  LAYER M1 ;
        RECT 11.744 13.236 11.776 13.308 ;
  LAYER M2 ;
        RECT 11.724 13.256 11.796 13.288 ;
  LAYER M2 ;
        RECT 9.008 13.256 11.76 13.288 ;
  LAYER M1 ;
        RECT 8.992 13.236 9.024 13.308 ;
  LAYER M2 ;
        RECT 8.972 13.256 9.044 13.288 ;
  LAYER M1 ;
        RECT 8.992 0.048 9.024 0.12 ;
  LAYER M2 ;
        RECT 8.972 0.068 9.044 0.1 ;
  LAYER M1 ;
        RECT 8.992 0.084 9.024 0.504 ;
  LAYER M1 ;
        RECT 8.992 0.504 9.024 13.272 ;
  LAYER M2 ;
        RECT 3.056 0.068 9.008 0.1 ;
  LAYER M1 ;
        RECT 3.424 9.456 3.456 9.528 ;
  LAYER M2 ;
        RECT 3.404 9.476 3.476 9.508 ;
  LAYER M2 ;
        RECT 3.216 9.476 3.44 9.508 ;
  LAYER M1 ;
        RECT 3.2 9.456 3.232 9.528 ;
  LAYER M2 ;
        RECT 3.18 9.476 3.252 9.508 ;
  LAYER M1 ;
        RECT 3.424 12.564 3.456 12.636 ;
  LAYER M2 ;
        RECT 3.404 12.584 3.476 12.616 ;
  LAYER M2 ;
        RECT 3.216 12.584 3.44 12.616 ;
  LAYER M1 ;
        RECT 3.2 12.564 3.232 12.636 ;
  LAYER M2 ;
        RECT 3.18 12.584 3.252 12.616 ;
  LAYER M1 ;
        RECT 3.424 6.348 3.456 6.42 ;
  LAYER M2 ;
        RECT 3.404 6.368 3.476 6.4 ;
  LAYER M2 ;
        RECT 3.216 6.368 3.44 6.4 ;
  LAYER M1 ;
        RECT 3.2 6.348 3.232 6.42 ;
  LAYER M2 ;
        RECT 3.18 6.368 3.252 6.4 ;
  LAYER M1 ;
        RECT 3.2 16.26 3.232 16.332 ;
  LAYER M2 ;
        RECT 3.18 16.28 3.252 16.312 ;
  LAYER M1 ;
        RECT 3.2 16.044 3.232 16.296 ;
  LAYER M1 ;
        RECT 3.2 6.384 3.232 16.044 ;
  LAYER M1 ;
        RECT 6.4 9.456 6.432 9.528 ;
  LAYER M2 ;
        RECT 6.38 9.476 6.452 9.508 ;
  LAYER M1 ;
        RECT 6.4 9.492 6.432 9.66 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M2 ;
        RECT 6.416 9.644 9.168 9.676 ;
  LAYER M1 ;
        RECT 9.152 9.624 9.184 9.696 ;
  LAYER M2 ;
        RECT 9.132 9.644 9.204 9.676 ;
  LAYER M1 ;
        RECT 6.4 6.348 6.432 6.42 ;
  LAYER M2 ;
        RECT 6.38 6.368 6.452 6.4 ;
  LAYER M1 ;
        RECT 6.4 6.384 6.432 6.552 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.416 6.536 9.168 6.568 ;
  LAYER M1 ;
        RECT 9.152 6.516 9.184 6.588 ;
  LAYER M2 ;
        RECT 9.132 6.536 9.204 6.568 ;
  LAYER M1 ;
        RECT 6.4 12.564 6.432 12.636 ;
  LAYER M2 ;
        RECT 6.38 12.584 6.452 12.616 ;
  LAYER M1 ;
        RECT 6.4 12.6 6.432 12.768 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M2 ;
        RECT 6.416 12.752 9.168 12.784 ;
  LAYER M1 ;
        RECT 9.152 12.732 9.184 12.804 ;
  LAYER M2 ;
        RECT 9.132 12.752 9.204 12.784 ;
  LAYER M1 ;
        RECT 9.152 16.26 9.184 16.332 ;
  LAYER M2 ;
        RECT 9.132 16.28 9.204 16.312 ;
  LAYER M1 ;
        RECT 9.152 16.044 9.184 16.296 ;
  LAYER M1 ;
        RECT 9.152 6.552 9.184 16.044 ;
  LAYER M2 ;
        RECT 3.216 16.28 9.168 16.312 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M2 ;
        RECT 0.08 3.26 0.464 3.292 ;
  LAYER M1 ;
        RECT 0.064 3.24 0.096 3.312 ;
  LAYER M2 ;
        RECT 0.044 3.26 0.116 3.292 ;
  LAYER M1 ;
        RECT 0.448 6.348 0.48 6.42 ;
  LAYER M2 ;
        RECT 0.428 6.368 0.5 6.4 ;
  LAYER M2 ;
        RECT 0.08 6.368 0.464 6.4 ;
  LAYER M1 ;
        RECT 0.064 6.348 0.096 6.42 ;
  LAYER M2 ;
        RECT 0.044 6.368 0.116 6.4 ;
  LAYER M1 ;
        RECT 0.448 9.456 0.48 9.528 ;
  LAYER M2 ;
        RECT 0.428 9.476 0.5 9.508 ;
  LAYER M2 ;
        RECT 0.08 9.476 0.464 9.508 ;
  LAYER M1 ;
        RECT 0.064 9.456 0.096 9.528 ;
  LAYER M2 ;
        RECT 0.044 9.476 0.116 9.508 ;
  LAYER M1 ;
        RECT 0.448 12.564 0.48 12.636 ;
  LAYER M2 ;
        RECT 0.428 12.584 0.5 12.616 ;
  LAYER M2 ;
        RECT 0.08 12.584 0.464 12.616 ;
  LAYER M1 ;
        RECT 0.064 12.564 0.096 12.636 ;
  LAYER M2 ;
        RECT 0.044 12.584 0.116 12.616 ;
  LAYER M1 ;
        RECT 0.448 15.672 0.48 15.744 ;
  LAYER M2 ;
        RECT 0.428 15.692 0.5 15.724 ;
  LAYER M2 ;
        RECT 0.08 15.692 0.464 15.724 ;
  LAYER M1 ;
        RECT 0.064 15.672 0.096 15.744 ;
  LAYER M2 ;
        RECT 0.044 15.692 0.116 15.724 ;
  LAYER M1 ;
        RECT 0.064 16.428 0.096 16.5 ;
  LAYER M2 ;
        RECT 0.044 16.448 0.116 16.48 ;
  LAYER M1 ;
        RECT 0.064 16.044 0.096 16.464 ;
  LAYER M1 ;
        RECT 0.064 3.276 0.096 16.044 ;
  LAYER M1 ;
        RECT 9.376 3.24 9.408 3.312 ;
  LAYER M2 ;
        RECT 9.356 3.26 9.428 3.292 ;
  LAYER M1 ;
        RECT 9.376 3.276 9.408 3.444 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M2 ;
        RECT 9.392 3.428 11.984 3.46 ;
  LAYER M1 ;
        RECT 11.968 3.408 12 3.48 ;
  LAYER M2 ;
        RECT 11.948 3.428 12.02 3.46 ;
  LAYER M1 ;
        RECT 9.376 6.348 9.408 6.42 ;
  LAYER M2 ;
        RECT 9.356 6.368 9.428 6.4 ;
  LAYER M1 ;
        RECT 9.376 6.384 9.408 6.552 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M2 ;
        RECT 9.392 6.536 11.984 6.568 ;
  LAYER M1 ;
        RECT 11.968 6.516 12 6.588 ;
  LAYER M2 ;
        RECT 11.948 6.536 12.02 6.568 ;
  LAYER M1 ;
        RECT 9.376 9.456 9.408 9.528 ;
  LAYER M2 ;
        RECT 9.356 9.476 9.428 9.508 ;
  LAYER M1 ;
        RECT 9.376 9.492 9.408 9.66 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M2 ;
        RECT 9.392 9.644 11.984 9.676 ;
  LAYER M1 ;
        RECT 11.968 9.624 12 9.696 ;
  LAYER M2 ;
        RECT 11.948 9.644 12.02 9.676 ;
  LAYER M1 ;
        RECT 9.376 12.564 9.408 12.636 ;
  LAYER M2 ;
        RECT 9.356 12.584 9.428 12.616 ;
  LAYER M1 ;
        RECT 9.376 12.6 9.408 12.768 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M2 ;
        RECT 9.392 12.752 11.984 12.784 ;
  LAYER M1 ;
        RECT 11.968 12.732 12 12.804 ;
  LAYER M2 ;
        RECT 11.948 12.752 12.02 12.784 ;
  LAYER M1 ;
        RECT 9.376 15.672 9.408 15.744 ;
  LAYER M2 ;
        RECT 9.356 15.692 9.428 15.724 ;
  LAYER M1 ;
        RECT 9.376 15.708 9.408 15.876 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M2 ;
        RECT 9.392 15.86 11.984 15.892 ;
  LAYER M1 ;
        RECT 11.968 15.84 12 15.912 ;
  LAYER M2 ;
        RECT 11.948 15.86 12.02 15.892 ;
  LAYER M1 ;
        RECT 11.968 16.428 12 16.5 ;
  LAYER M2 ;
        RECT 11.948 16.448 12.02 16.48 ;
  LAYER M1 ;
        RECT 11.968 16.044 12 16.464 ;
  LAYER M1 ;
        RECT 11.968 3.444 12 16.044 ;
  LAYER M2 ;
        RECT 0.08 16.448 11.984 16.48 ;
  LAYER M1 ;
        RECT 3.424 3.24 3.456 3.312 ;
  LAYER M2 ;
        RECT 3.404 3.26 3.476 3.292 ;
  LAYER M2 ;
        RECT 0.464 3.26 3.44 3.292 ;
  LAYER M1 ;
        RECT 0.448 3.24 0.48 3.312 ;
  LAYER M2 ;
        RECT 0.428 3.26 0.5 3.292 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M2 ;
        RECT 0.464 15.692 3.44 15.724 ;
  LAYER M1 ;
        RECT 0.448 15.672 0.48 15.744 ;
  LAYER M2 ;
        RECT 0.428 15.692 0.5 15.724 ;
  LAYER M1 ;
        RECT 6.4 15.672 6.432 15.744 ;
  LAYER M2 ;
        RECT 6.38 15.692 6.452 15.724 ;
  LAYER M2 ;
        RECT 3.44 15.692 6.416 15.724 ;
  LAYER M1 ;
        RECT 3.424 15.672 3.456 15.744 ;
  LAYER M2 ;
        RECT 3.404 15.692 3.476 15.724 ;
  LAYER M1 ;
        RECT 6.4 3.24 6.432 3.312 ;
  LAYER M2 ;
        RECT 6.38 3.26 6.452 3.292 ;
  LAYER M2 ;
        RECT 6.416 3.26 9.392 3.292 ;
  LAYER M1 ;
        RECT 9.376 3.24 9.408 3.312 ;
  LAYER M2 ;
        RECT 9.356 3.26 9.428 3.292 ;
  LAYER M1 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M3 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.896 3.36 ;
  LAYER M1 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M3 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M2 ;
        RECT 0.4 3.864 2.896 6.468 ;
  LAYER M1 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M3 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M2 ;
        RECT 0.4 6.972 2.896 9.576 ;
  LAYER M1 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M3 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M2 ;
        RECT 0.4 10.08 2.896 12.684 ;
  LAYER M1 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M3 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M2 ;
        RECT 0.4 13.188 2.896 15.792 ;
  LAYER M1 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M3 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M2 ;
        RECT 3.376 0.756 5.872 3.36 ;
  LAYER M1 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M3 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M2 ;
        RECT 3.376 3.864 5.872 6.468 ;
  LAYER M1 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M3 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M2 ;
        RECT 3.376 6.972 5.872 9.576 ;
  LAYER M1 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M3 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M2 ;
        RECT 3.376 10.08 5.872 12.684 ;
  LAYER M1 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M3 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M2 ;
        RECT 3.376 13.188 5.872 15.792 ;
  LAYER M1 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M3 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M2 ;
        RECT 6.352 0.756 8.848 3.36 ;
  LAYER M1 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M3 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M2 ;
        RECT 6.352 3.864 8.848 6.468 ;
  LAYER M1 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M3 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M2 ;
        RECT 6.352 6.972 8.848 9.576 ;
  LAYER M1 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M3 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M2 ;
        RECT 6.352 10.08 8.848 12.684 ;
  LAYER M1 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M3 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M2 ;
        RECT 6.352 13.188 8.848 15.792 ;
  LAYER M1 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M3 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M2 ;
        RECT 9.328 0.756 11.824 3.36 ;
  LAYER M1 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M3 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M2 ;
        RECT 9.328 3.864 11.824 6.468 ;
  LAYER M1 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M3 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M2 ;
        RECT 9.328 6.972 11.824 9.576 ;
  LAYER M1 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M3 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M2 ;
        RECT 9.328 10.08 11.824 12.684 ;
  LAYER M1 ;
        RECT 9.328 13.188 11.824 15.792 ;
  LAYER M3 ;
        RECT 9.328 13.188 11.824 15.792 ;
  LAYER M2 ;
        RECT 9.328 13.188 11.824 15.792 ;
  END 
END Cap_60fF
