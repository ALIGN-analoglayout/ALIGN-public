
.subckt Sanitized_Coarse_Comp_CK VCTIN DVDD DVSS OUTNC OUTPC VALIDC ST_FINE CKSBT CKC
XI67 net07 VCTIN DVDD DVSS net09 PINVD0YVT
XI46 net30 VCTIN DVDD DVSS net29 PINVD0YVT
XI21 net33 VCTIN DVDD DVSS net32 PINVD0YVT
XI12 net34 VCTIN DVDD DVSS net33 PINVD0YVT
XI47 net31 VCTIN DVDD DVSS net30 PINVD0YVT
XI0 net29 net07 DVDD DVSS INVD0HVT
XI22 net32 net31 DVDD DVSS INVD0HVT
XI3 OUTNC OUTPC VALIDC DVDD DVSS ND2D3LVT
XI218 VALIDC ST_FINE CKSBT net34 DVDD DVSS NR3D1LVT
XI65 net09 CKC DVDD DVSS INVD2LVT
.ends Sanitized_Coarse_Comp_CK

.subckt PINVD0YVT I P VDD VSS ZN
xMM4 ZN I net11 VSS Switch_NMOS_n12_X1_Y1
xMM1 net11 P VSS VSS Switch_NMOS_n12_X1_Y1
xMM3 net09 VSS VDD VDD Switch_PMOS_n12_X1_Y1
xMM0 ZN I net09 VDD Switch_PMOS_n12_X1_Y1
.ends PINVD0YVT

.subckt Switch_NMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_NMOS_n12_X1_Y1

.subckt Switch_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends Switch_PMOS_n12_X1_Y1

.subckt INVD0HVT I ZN VDD VSS
xMMU1_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD0HVT

.subckt CMC_NMOS_S_n12_X1_Y1 B DA G S DB
xM0 DA G S B Switch_NMOS_n12_X1_Y1
xM1 DB G S B Switch_NMOS_n12_X1_Y1
.ends CMC_NMOS_S_n12_X1_Y1

.subckt ND2D3LVT A1 A2 ZN VDD VSS
xMMU3_1_M_u3 ZN A1 net20 VSS Switch_NMOS_n12_X1_Y1
xMMU3_2_M_u4 net13 A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMMU3_0_M_u3 ZN A1 net21 VSS Switch_NMOS_n12_X1_Y1
xMMU3_2_M_u3 ZN A1 net13 VSS Switch_NMOS_n12_X1_Y1
xMMU3_2_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU3_1_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU3_0_M_u2 ZN A2 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU3_0_M_u1 ZN A1 VDD VDD Switch_PMOS_n12_X1_Y1
xMMU3_1_M_u4_MMU3_0_M_u4 net20 A2 VSS net21 VSS CMC_NMOS_S_n12_X1_Y1
.ends ND2D3LVT

.subckt CMC_NMOS_S_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends CMC_NMOS_S_n12_X1_Y1

.subckt CMC_PMOS_S_n12_X1_Y1 B DA G S DB
xM0 DA G S B Switch_PMOS_n12_X1_Y1
xM1 DB G S B Switch_PMOS_n12_X1_Y1
.ends CMC_PMOS_S_n12_X1_Y1

.subckt CMC_PMOS_n12_X1_Y1 B DA G SA DB SB
xM0 DA G SA B Switch_PMOS_n12_X1_Y1
xM1 DB G SB B Switch_PMOS_n12_X1_Y1
.ends CMC_PMOS_n12_X1_Y1

.subckt NR3D1LVT A1 A2 A3 ZN VDD VSS
xMMI1_1 ZN A1 net5 VDD Switch_PMOS_n12_X1_Y1
xMMI1_0 ZN A1 net9 VDD Switch_PMOS_n12_X1_Y1
xMMI3 ZN A1 VSS VSS Switch_NMOS_n12_X1_Y1
xMMI2 ZN A2 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u4 ZN A3 VSS VSS Switch_NMOS_n12_X1_Y1
xMM_u1_1_MM_u1_0 net1 A3 VDD net17 VDD CMC_PMOS_S_n12_X1_Y1
xMMI0_1_MMI0_0 net5 A2 net1 net9 net17 VDD CMC_PMOS_n12_X1_Y1
.ends NR3D1LVT

.subckt CMC_PMOS_S_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends CMC_PMOS_S_n12_X1_Y1

.subckt CMC_PMOS_n12_X1_Y1 D G S B
m0 D G S1 B nmos_rvt  l=1e-08 w=1e-08 m=1
m1 S1 G S B nmos_rvt  l=1e-08 w=1e-08 m=1
.ends CMC_PMOS_n12_X1_Y1

.subckt INVD2LVT I ZN VDD VSS
xMMU1_0_M_u2 ZN I VSS VSS Switch_NMOS_n12_X1_Y1
xMMU1_0_M_u3 ZN I VDD VDD Switch_PMOS_n12_X1_Y1
.ends INVD2LVT
