MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 8.96 BY 24.528 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.104 24.24 3.136 24.312 ;
      LAYER M2 ;
        RECT 3.084 24.26 3.156 24.292 ;
      LAYER M1 ;
        RECT 5.984 24.24 6.016 24.312 ;
      LAYER M2 ;
        RECT 5.964 24.26 6.036 24.292 ;
      LAYER M2 ;
        RECT 3.12 24.26 6 24.292 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
      LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
      LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
      LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
      LAYER M2 ;
        RECT 2.96 0.236 5.84 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M2 ;
        RECT 2.96 9.56 5.68 9.592 ;
  LAYER M1 ;
        RECT 2.944 9.54 2.976 9.612 ;
  LAYER M2 ;
        RECT 2.924 9.56 2.996 9.592 ;
  LAYER M1 ;
        RECT 5.664 12.48 5.696 12.552 ;
  LAYER M2 ;
        RECT 5.644 12.5 5.716 12.532 ;
  LAYER M2 ;
        RECT 2.96 12.5 5.68 12.532 ;
  LAYER M1 ;
        RECT 2.944 12.48 2.976 12.552 ;
  LAYER M2 ;
        RECT 2.924 12.5 2.996 12.532 ;
  LAYER M1 ;
        RECT 5.664 6.6 5.696 6.672 ;
  LAYER M2 ;
        RECT 5.644 6.62 5.716 6.652 ;
  LAYER M2 ;
        RECT 2.96 6.62 5.68 6.652 ;
  LAYER M1 ;
        RECT 2.944 6.6 2.976 6.672 ;
  LAYER M2 ;
        RECT 2.924 6.62 2.996 6.652 ;
  LAYER M1 ;
        RECT 5.664 15.42 5.696 15.492 ;
  LAYER M2 ;
        RECT 5.644 15.44 5.716 15.472 ;
  LAYER M2 ;
        RECT 2.96 15.44 5.68 15.472 ;
  LAYER M1 ;
        RECT 2.944 15.42 2.976 15.492 ;
  LAYER M2 ;
        RECT 2.924 15.44 2.996 15.472 ;
  LAYER M1 ;
        RECT 5.664 3.66 5.696 3.732 ;
  LAYER M2 ;
        RECT 5.644 3.68 5.716 3.712 ;
  LAYER M2 ;
        RECT 2.96 3.68 5.68 3.712 ;
  LAYER M1 ;
        RECT 2.944 3.66 2.976 3.732 ;
  LAYER M2 ;
        RECT 2.924 3.68 2.996 3.712 ;
  LAYER M1 ;
        RECT 5.664 18.36 5.696 18.432 ;
  LAYER M2 ;
        RECT 5.644 18.38 5.716 18.412 ;
  LAYER M2 ;
        RECT 2.96 18.38 5.68 18.412 ;
  LAYER M1 ;
        RECT 2.944 18.36 2.976 18.432 ;
  LAYER M2 ;
        RECT 2.924 18.38 2.996 18.412 ;
  LAYER M1 ;
        RECT 2.944 0.216 2.976 0.288 ;
  LAYER M2 ;
        RECT 2.924 0.236 2.996 0.268 ;
  LAYER M1 ;
        RECT 2.944 0.252 2.976 0.42 ;
  LAYER M1 ;
        RECT 2.944 0.42 2.976 18.396 ;
  LAYER M1 ;
        RECT 5.664 9.54 5.696 9.612 ;
  LAYER M2 ;
        RECT 5.644 9.56 5.716 9.592 ;
  LAYER M1 ;
        RECT 5.664 9.408 5.696 9.576 ;
  LAYER M1 ;
        RECT 5.664 9.372 5.696 9.444 ;
  LAYER M2 ;
        RECT 5.644 9.392 5.716 9.424 ;
  LAYER M2 ;
        RECT 5.68 9.392 5.84 9.424 ;
  LAYER M1 ;
        RECT 5.824 9.372 5.856 9.444 ;
  LAYER M2 ;
        RECT 5.804 9.392 5.876 9.424 ;
  LAYER M1 ;
        RECT 5.664 12.48 5.696 12.552 ;
  LAYER M2 ;
        RECT 5.644 12.5 5.716 12.532 ;
  LAYER M1 ;
        RECT 5.664 12.348 5.696 12.516 ;
  LAYER M1 ;
        RECT 5.664 12.312 5.696 12.384 ;
  LAYER M2 ;
        RECT 5.644 12.332 5.716 12.364 ;
  LAYER M2 ;
        RECT 5.68 12.332 5.84 12.364 ;
  LAYER M1 ;
        RECT 5.824 12.312 5.856 12.384 ;
  LAYER M2 ;
        RECT 5.804 12.332 5.876 12.364 ;
  LAYER M1 ;
        RECT 5.664 6.6 5.696 6.672 ;
  LAYER M2 ;
        RECT 5.644 6.62 5.716 6.652 ;
  LAYER M1 ;
        RECT 5.664 6.468 5.696 6.636 ;
  LAYER M1 ;
        RECT 5.664 6.432 5.696 6.504 ;
  LAYER M2 ;
        RECT 5.644 6.452 5.716 6.484 ;
  LAYER M2 ;
        RECT 5.68 6.452 5.84 6.484 ;
  LAYER M1 ;
        RECT 5.824 6.432 5.856 6.504 ;
  LAYER M2 ;
        RECT 5.804 6.452 5.876 6.484 ;
  LAYER M1 ;
        RECT 5.664 15.42 5.696 15.492 ;
  LAYER M2 ;
        RECT 5.644 15.44 5.716 15.472 ;
  LAYER M1 ;
        RECT 5.664 15.288 5.696 15.456 ;
  LAYER M1 ;
        RECT 5.664 15.252 5.696 15.324 ;
  LAYER M2 ;
        RECT 5.644 15.272 5.716 15.304 ;
  LAYER M2 ;
        RECT 5.68 15.272 5.84 15.304 ;
  LAYER M1 ;
        RECT 5.824 15.252 5.856 15.324 ;
  LAYER M2 ;
        RECT 5.804 15.272 5.876 15.304 ;
  LAYER M1 ;
        RECT 5.664 3.66 5.696 3.732 ;
  LAYER M2 ;
        RECT 5.644 3.68 5.716 3.712 ;
  LAYER M1 ;
        RECT 5.664 3.528 5.696 3.696 ;
  LAYER M1 ;
        RECT 5.664 3.492 5.696 3.564 ;
  LAYER M2 ;
        RECT 5.644 3.512 5.716 3.544 ;
  LAYER M2 ;
        RECT 5.68 3.512 5.84 3.544 ;
  LAYER M1 ;
        RECT 5.824 3.492 5.856 3.564 ;
  LAYER M2 ;
        RECT 5.804 3.512 5.876 3.544 ;
  LAYER M1 ;
        RECT 5.664 18.36 5.696 18.432 ;
  LAYER M2 ;
        RECT 5.644 18.38 5.716 18.412 ;
  LAYER M1 ;
        RECT 5.664 18.228 5.696 18.396 ;
  LAYER M1 ;
        RECT 5.664 18.192 5.696 18.264 ;
  LAYER M2 ;
        RECT 5.644 18.212 5.716 18.244 ;
  LAYER M2 ;
        RECT 5.68 18.212 5.84 18.244 ;
  LAYER M1 ;
        RECT 5.824 18.192 5.856 18.264 ;
  LAYER M2 ;
        RECT 5.804 18.212 5.876 18.244 ;
  LAYER M1 ;
        RECT 5.824 0.216 5.856 0.288 ;
  LAYER M2 ;
        RECT 5.804 0.236 5.876 0.268 ;
  LAYER M1 ;
        RECT 5.824 0.252 5.856 0.42 ;
  LAYER M1 ;
        RECT 5.824 0.42 5.856 18.228 ;
  LAYER M2 ;
        RECT 2.96 0.236 5.84 0.268 ;
  LAYER M1 ;
        RECT 2.784 0.72 2.816 0.792 ;
  LAYER M2 ;
        RECT 2.764 0.74 2.836 0.772 ;
  LAYER M2 ;
        RECT 0.08 0.74 2.8 0.772 ;
  LAYER M1 ;
        RECT 0.064 0.72 0.096 0.792 ;
  LAYER M2 ;
        RECT 0.044 0.74 0.116 0.772 ;
  LAYER M1 ;
        RECT 2.784 3.66 2.816 3.732 ;
  LAYER M2 ;
        RECT 2.764 3.68 2.836 3.712 ;
  LAYER M2 ;
        RECT 0.08 3.68 2.8 3.712 ;
  LAYER M1 ;
        RECT 0.064 3.66 0.096 3.732 ;
  LAYER M2 ;
        RECT 0.044 3.68 0.116 3.712 ;
  LAYER M1 ;
        RECT 2.784 6.6 2.816 6.672 ;
  LAYER M2 ;
        RECT 2.764 6.62 2.836 6.652 ;
  LAYER M2 ;
        RECT 0.08 6.62 2.8 6.652 ;
  LAYER M1 ;
        RECT 0.064 6.6 0.096 6.672 ;
  LAYER M2 ;
        RECT 0.044 6.62 0.116 6.652 ;
  LAYER M1 ;
        RECT 2.784 9.54 2.816 9.612 ;
  LAYER M2 ;
        RECT 2.764 9.56 2.836 9.592 ;
  LAYER M2 ;
        RECT 0.08 9.56 2.8 9.592 ;
  LAYER M1 ;
        RECT 0.064 9.54 0.096 9.612 ;
  LAYER M2 ;
        RECT 0.044 9.56 0.116 9.592 ;
  LAYER M1 ;
        RECT 2.784 12.48 2.816 12.552 ;
  LAYER M2 ;
        RECT 2.764 12.5 2.836 12.532 ;
  LAYER M2 ;
        RECT 0.08 12.5 2.8 12.532 ;
  LAYER M1 ;
        RECT 0.064 12.48 0.096 12.552 ;
  LAYER M2 ;
        RECT 0.044 12.5 0.116 12.532 ;
  LAYER M1 ;
        RECT 2.784 15.42 2.816 15.492 ;
  LAYER M2 ;
        RECT 2.764 15.44 2.836 15.472 ;
  LAYER M2 ;
        RECT 0.08 15.44 2.8 15.472 ;
  LAYER M1 ;
        RECT 0.064 15.42 0.096 15.492 ;
  LAYER M2 ;
        RECT 0.044 15.44 0.116 15.472 ;
  LAYER M1 ;
        RECT 2.784 18.36 2.816 18.432 ;
  LAYER M2 ;
        RECT 2.764 18.38 2.836 18.412 ;
  LAYER M2 ;
        RECT 0.08 18.38 2.8 18.412 ;
  LAYER M1 ;
        RECT 0.064 18.36 0.096 18.432 ;
  LAYER M2 ;
        RECT 0.044 18.38 0.116 18.412 ;
  LAYER M1 ;
        RECT 2.784 21.3 2.816 21.372 ;
  LAYER M2 ;
        RECT 2.764 21.32 2.836 21.352 ;
  LAYER M2 ;
        RECT 0.08 21.32 2.8 21.352 ;
  LAYER M1 ;
        RECT 0.064 21.3 0.096 21.372 ;
  LAYER M2 ;
        RECT 0.044 21.32 0.116 21.352 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.42 ;
  LAYER M1 ;
        RECT 0.064 0.42 0.096 21.336 ;
  LAYER M1 ;
        RECT 8.544 0.72 8.576 0.792 ;
  LAYER M2 ;
        RECT 8.524 0.74 8.596 0.772 ;
  LAYER M1 ;
        RECT 8.544 0.588 8.576 0.756 ;
  LAYER M1 ;
        RECT 8.544 0.552 8.576 0.624 ;
  LAYER M2 ;
        RECT 8.524 0.572 8.596 0.604 ;
  LAYER M2 ;
        RECT 8.56 0.572 8.72 0.604 ;
  LAYER M1 ;
        RECT 8.704 0.552 8.736 0.624 ;
  LAYER M2 ;
        RECT 8.684 0.572 8.756 0.604 ;
  LAYER M1 ;
        RECT 8.544 3.66 8.576 3.732 ;
  LAYER M2 ;
        RECT 8.524 3.68 8.596 3.712 ;
  LAYER M1 ;
        RECT 8.544 3.528 8.576 3.696 ;
  LAYER M1 ;
        RECT 8.544 3.492 8.576 3.564 ;
  LAYER M2 ;
        RECT 8.524 3.512 8.596 3.544 ;
  LAYER M2 ;
        RECT 8.56 3.512 8.72 3.544 ;
  LAYER M1 ;
        RECT 8.704 3.492 8.736 3.564 ;
  LAYER M2 ;
        RECT 8.684 3.512 8.756 3.544 ;
  LAYER M1 ;
        RECT 8.544 6.6 8.576 6.672 ;
  LAYER M2 ;
        RECT 8.524 6.62 8.596 6.652 ;
  LAYER M1 ;
        RECT 8.544 6.468 8.576 6.636 ;
  LAYER M1 ;
        RECT 8.544 6.432 8.576 6.504 ;
  LAYER M2 ;
        RECT 8.524 6.452 8.596 6.484 ;
  LAYER M2 ;
        RECT 8.56 6.452 8.72 6.484 ;
  LAYER M1 ;
        RECT 8.704 6.432 8.736 6.504 ;
  LAYER M2 ;
        RECT 8.684 6.452 8.756 6.484 ;
  LAYER M1 ;
        RECT 8.544 9.54 8.576 9.612 ;
  LAYER M2 ;
        RECT 8.524 9.56 8.596 9.592 ;
  LAYER M1 ;
        RECT 8.544 9.408 8.576 9.576 ;
  LAYER M1 ;
        RECT 8.544 9.372 8.576 9.444 ;
  LAYER M2 ;
        RECT 8.524 9.392 8.596 9.424 ;
  LAYER M2 ;
        RECT 8.56 9.392 8.72 9.424 ;
  LAYER M1 ;
        RECT 8.704 9.372 8.736 9.444 ;
  LAYER M2 ;
        RECT 8.684 9.392 8.756 9.424 ;
  LAYER M1 ;
        RECT 8.544 12.48 8.576 12.552 ;
  LAYER M2 ;
        RECT 8.524 12.5 8.596 12.532 ;
  LAYER M1 ;
        RECT 8.544 12.348 8.576 12.516 ;
  LAYER M1 ;
        RECT 8.544 12.312 8.576 12.384 ;
  LAYER M2 ;
        RECT 8.524 12.332 8.596 12.364 ;
  LAYER M2 ;
        RECT 8.56 12.332 8.72 12.364 ;
  LAYER M1 ;
        RECT 8.704 12.312 8.736 12.384 ;
  LAYER M2 ;
        RECT 8.684 12.332 8.756 12.364 ;
  LAYER M1 ;
        RECT 8.544 15.42 8.576 15.492 ;
  LAYER M2 ;
        RECT 8.524 15.44 8.596 15.472 ;
  LAYER M1 ;
        RECT 8.544 15.288 8.576 15.456 ;
  LAYER M1 ;
        RECT 8.544 15.252 8.576 15.324 ;
  LAYER M2 ;
        RECT 8.524 15.272 8.596 15.304 ;
  LAYER M2 ;
        RECT 8.56 15.272 8.72 15.304 ;
  LAYER M1 ;
        RECT 8.704 15.252 8.736 15.324 ;
  LAYER M2 ;
        RECT 8.684 15.272 8.756 15.304 ;
  LAYER M1 ;
        RECT 8.544 18.36 8.576 18.432 ;
  LAYER M2 ;
        RECT 8.524 18.38 8.596 18.412 ;
  LAYER M1 ;
        RECT 8.544 18.228 8.576 18.396 ;
  LAYER M1 ;
        RECT 8.544 18.192 8.576 18.264 ;
  LAYER M2 ;
        RECT 8.524 18.212 8.596 18.244 ;
  LAYER M2 ;
        RECT 8.56 18.212 8.72 18.244 ;
  LAYER M1 ;
        RECT 8.704 18.192 8.736 18.264 ;
  LAYER M2 ;
        RECT 8.684 18.212 8.756 18.244 ;
  LAYER M1 ;
        RECT 8.544 21.3 8.576 21.372 ;
  LAYER M2 ;
        RECT 8.524 21.32 8.596 21.352 ;
  LAYER M1 ;
        RECT 8.544 21.168 8.576 21.336 ;
  LAYER M1 ;
        RECT 8.544 21.132 8.576 21.204 ;
  LAYER M2 ;
        RECT 8.524 21.152 8.596 21.184 ;
  LAYER M2 ;
        RECT 8.56 21.152 8.72 21.184 ;
  LAYER M1 ;
        RECT 8.704 21.132 8.736 21.204 ;
  LAYER M2 ;
        RECT 8.684 21.152 8.756 21.184 ;
  LAYER M1 ;
        RECT 8.704 0.048 8.736 0.12 ;
  LAYER M2 ;
        RECT 8.684 0.068 8.756 0.1 ;
  LAYER M1 ;
        RECT 8.704 0.084 8.736 0.42 ;
  LAYER M1 ;
        RECT 8.704 0.42 8.736 21.168 ;
  LAYER M2 ;
        RECT 0.08 0.068 8.72 0.1 ;
  LAYER M1 ;
        RECT 5.664 0.72 5.696 0.792 ;
  LAYER M2 ;
        RECT 5.644 0.74 5.716 0.772 ;
  LAYER M2 ;
        RECT 2.8 0.74 5.68 0.772 ;
  LAYER M1 ;
        RECT 2.784 0.72 2.816 0.792 ;
  LAYER M2 ;
        RECT 2.764 0.74 2.836 0.772 ;
  LAYER M1 ;
        RECT 5.664 21.3 5.696 21.372 ;
  LAYER M2 ;
        RECT 5.644 21.32 5.716 21.352 ;
  LAYER M2 ;
        RECT 2.8 21.32 5.68 21.352 ;
  LAYER M1 ;
        RECT 2.784 21.3 2.816 21.372 ;
  LAYER M2 ;
        RECT 2.764 21.32 2.836 21.352 ;
  LAYER M1 ;
        RECT 3.264 11.976 3.296 12.048 ;
  LAYER M2 ;
        RECT 3.244 11.996 3.316 12.028 ;
  LAYER M2 ;
        RECT 3.12 11.996 3.28 12.028 ;
  LAYER M1 ;
        RECT 3.104 11.976 3.136 12.048 ;
  LAYER M2 ;
        RECT 3.084 11.996 3.156 12.028 ;
  LAYER M1 ;
        RECT 3.264 14.916 3.296 14.988 ;
  LAYER M2 ;
        RECT 3.244 14.936 3.316 14.968 ;
  LAYER M2 ;
        RECT 3.12 14.936 3.28 14.968 ;
  LAYER M1 ;
        RECT 3.104 14.916 3.136 14.988 ;
  LAYER M2 ;
        RECT 3.084 14.936 3.156 14.968 ;
  LAYER M1 ;
        RECT 3.264 9.036 3.296 9.108 ;
  LAYER M2 ;
        RECT 3.244 9.056 3.316 9.088 ;
  LAYER M2 ;
        RECT 3.12 9.056 3.28 9.088 ;
  LAYER M1 ;
        RECT 3.104 9.036 3.136 9.108 ;
  LAYER M2 ;
        RECT 3.084 9.056 3.156 9.088 ;
  LAYER M1 ;
        RECT 3.264 17.856 3.296 17.928 ;
  LAYER M2 ;
        RECT 3.244 17.876 3.316 17.908 ;
  LAYER M2 ;
        RECT 3.12 17.876 3.28 17.908 ;
  LAYER M1 ;
        RECT 3.104 17.856 3.136 17.928 ;
  LAYER M2 ;
        RECT 3.084 17.876 3.156 17.908 ;
  LAYER M1 ;
        RECT 3.264 6.096 3.296 6.168 ;
  LAYER M2 ;
        RECT 3.244 6.116 3.316 6.148 ;
  LAYER M2 ;
        RECT 3.12 6.116 3.28 6.148 ;
  LAYER M1 ;
        RECT 3.104 6.096 3.136 6.168 ;
  LAYER M2 ;
        RECT 3.084 6.116 3.156 6.148 ;
  LAYER M1 ;
        RECT 3.264 20.796 3.296 20.868 ;
  LAYER M2 ;
        RECT 3.244 20.816 3.316 20.848 ;
  LAYER M2 ;
        RECT 3.12 20.816 3.28 20.848 ;
  LAYER M1 ;
        RECT 3.104 20.796 3.136 20.868 ;
  LAYER M2 ;
        RECT 3.084 20.816 3.156 20.848 ;
  LAYER M1 ;
        RECT 3.104 24.24 3.136 24.312 ;
  LAYER M2 ;
        RECT 3.084 24.26 3.156 24.292 ;
  LAYER M1 ;
        RECT 3.104 24.108 3.136 24.276 ;
  LAYER M1 ;
        RECT 3.104 6.132 3.136 24.108 ;
  LAYER M1 ;
        RECT 3.264 11.976 3.296 12.048 ;
  LAYER M2 ;
        RECT 3.244 11.996 3.316 12.028 ;
  LAYER M1 ;
        RECT 3.264 12.012 3.296 12.18 ;
  LAYER M1 ;
        RECT 3.264 12.144 3.296 12.216 ;
  LAYER M2 ;
        RECT 3.244 12.164 3.316 12.196 ;
  LAYER M2 ;
        RECT 3.28 12.164 6 12.196 ;
  LAYER M1 ;
        RECT 5.984 12.144 6.016 12.216 ;
  LAYER M2 ;
        RECT 5.964 12.164 6.036 12.196 ;
  LAYER M1 ;
        RECT 3.264 14.916 3.296 14.988 ;
  LAYER M2 ;
        RECT 3.244 14.936 3.316 14.968 ;
  LAYER M1 ;
        RECT 3.264 14.952 3.296 15.12 ;
  LAYER M1 ;
        RECT 3.264 15.084 3.296 15.156 ;
  LAYER M2 ;
        RECT 3.244 15.104 3.316 15.136 ;
  LAYER M2 ;
        RECT 3.28 15.104 6 15.136 ;
  LAYER M1 ;
        RECT 5.984 15.084 6.016 15.156 ;
  LAYER M2 ;
        RECT 5.964 15.104 6.036 15.136 ;
  LAYER M1 ;
        RECT 3.264 9.036 3.296 9.108 ;
  LAYER M2 ;
        RECT 3.244 9.056 3.316 9.088 ;
  LAYER M1 ;
        RECT 3.264 9.072 3.296 9.24 ;
  LAYER M1 ;
        RECT 3.264 9.204 3.296 9.276 ;
  LAYER M2 ;
        RECT 3.244 9.224 3.316 9.256 ;
  LAYER M2 ;
        RECT 3.28 9.224 6 9.256 ;
  LAYER M1 ;
        RECT 5.984 9.204 6.016 9.276 ;
  LAYER M2 ;
        RECT 5.964 9.224 6.036 9.256 ;
  LAYER M1 ;
        RECT 3.264 17.856 3.296 17.928 ;
  LAYER M2 ;
        RECT 3.244 17.876 3.316 17.908 ;
  LAYER M1 ;
        RECT 3.264 17.892 3.296 18.06 ;
  LAYER M1 ;
        RECT 3.264 18.024 3.296 18.096 ;
  LAYER M2 ;
        RECT 3.244 18.044 3.316 18.076 ;
  LAYER M2 ;
        RECT 3.28 18.044 6 18.076 ;
  LAYER M1 ;
        RECT 5.984 18.024 6.016 18.096 ;
  LAYER M2 ;
        RECT 5.964 18.044 6.036 18.076 ;
  LAYER M1 ;
        RECT 3.264 6.096 3.296 6.168 ;
  LAYER M2 ;
        RECT 3.244 6.116 3.316 6.148 ;
  LAYER M1 ;
        RECT 3.264 6.132 3.296 6.3 ;
  LAYER M1 ;
        RECT 3.264 6.264 3.296 6.336 ;
  LAYER M2 ;
        RECT 3.244 6.284 3.316 6.316 ;
  LAYER M2 ;
        RECT 3.28 6.284 6 6.316 ;
  LAYER M1 ;
        RECT 5.984 6.264 6.016 6.336 ;
  LAYER M2 ;
        RECT 5.964 6.284 6.036 6.316 ;
  LAYER M1 ;
        RECT 3.264 20.796 3.296 20.868 ;
  LAYER M2 ;
        RECT 3.244 20.816 3.316 20.848 ;
  LAYER M1 ;
        RECT 3.264 20.832 3.296 21 ;
  LAYER M1 ;
        RECT 3.264 20.964 3.296 21.036 ;
  LAYER M2 ;
        RECT 3.244 20.984 3.316 21.016 ;
  LAYER M2 ;
        RECT 3.28 20.984 6 21.016 ;
  LAYER M1 ;
        RECT 5.984 20.964 6.016 21.036 ;
  LAYER M2 ;
        RECT 5.964 20.984 6.036 21.016 ;
  LAYER M1 ;
        RECT 5.984 24.24 6.016 24.312 ;
  LAYER M2 ;
        RECT 5.964 24.26 6.036 24.292 ;
  LAYER M1 ;
        RECT 5.984 24.108 6.016 24.276 ;
  LAYER M1 ;
        RECT 5.984 6.3 6.016 24.108 ;
  LAYER M2 ;
        RECT 3.12 24.26 6 24.292 ;
  LAYER M1 ;
        RECT 0.384 3.156 0.416 3.228 ;
  LAYER M2 ;
        RECT 0.364 3.176 0.436 3.208 ;
  LAYER M2 ;
        RECT 0.24 3.176 0.4 3.208 ;
  LAYER M1 ;
        RECT 0.224 3.156 0.256 3.228 ;
  LAYER M2 ;
        RECT 0.204 3.176 0.276 3.208 ;
  LAYER M1 ;
        RECT 0.384 6.096 0.416 6.168 ;
  LAYER M2 ;
        RECT 0.364 6.116 0.436 6.148 ;
  LAYER M2 ;
        RECT 0.24 6.116 0.4 6.148 ;
  LAYER M1 ;
        RECT 0.224 6.096 0.256 6.168 ;
  LAYER M2 ;
        RECT 0.204 6.116 0.276 6.148 ;
  LAYER M1 ;
        RECT 0.384 9.036 0.416 9.108 ;
  LAYER M2 ;
        RECT 0.364 9.056 0.436 9.088 ;
  LAYER M2 ;
        RECT 0.24 9.056 0.4 9.088 ;
  LAYER M1 ;
        RECT 0.224 9.036 0.256 9.108 ;
  LAYER M2 ;
        RECT 0.204 9.056 0.276 9.088 ;
  LAYER M1 ;
        RECT 0.384 11.976 0.416 12.048 ;
  LAYER M2 ;
        RECT 0.364 11.996 0.436 12.028 ;
  LAYER M2 ;
        RECT 0.24 11.996 0.4 12.028 ;
  LAYER M1 ;
        RECT 0.224 11.976 0.256 12.048 ;
  LAYER M2 ;
        RECT 0.204 11.996 0.276 12.028 ;
  LAYER M1 ;
        RECT 0.384 14.916 0.416 14.988 ;
  LAYER M2 ;
        RECT 0.364 14.936 0.436 14.968 ;
  LAYER M2 ;
        RECT 0.24 14.936 0.4 14.968 ;
  LAYER M1 ;
        RECT 0.224 14.916 0.256 14.988 ;
  LAYER M2 ;
        RECT 0.204 14.936 0.276 14.968 ;
  LAYER M1 ;
        RECT 0.384 17.856 0.416 17.928 ;
  LAYER M2 ;
        RECT 0.364 17.876 0.436 17.908 ;
  LAYER M2 ;
        RECT 0.24 17.876 0.4 17.908 ;
  LAYER M1 ;
        RECT 0.224 17.856 0.256 17.928 ;
  LAYER M2 ;
        RECT 0.204 17.876 0.276 17.908 ;
  LAYER M1 ;
        RECT 0.384 20.796 0.416 20.868 ;
  LAYER M2 ;
        RECT 0.364 20.816 0.436 20.848 ;
  LAYER M2 ;
        RECT 0.24 20.816 0.4 20.848 ;
  LAYER M1 ;
        RECT 0.224 20.796 0.256 20.868 ;
  LAYER M2 ;
        RECT 0.204 20.816 0.276 20.848 ;
  LAYER M1 ;
        RECT 0.384 23.736 0.416 23.808 ;
  LAYER M2 ;
        RECT 0.364 23.756 0.436 23.788 ;
  LAYER M2 ;
        RECT 0.24 23.756 0.4 23.788 ;
  LAYER M1 ;
        RECT 0.224 23.736 0.256 23.808 ;
  LAYER M2 ;
        RECT 0.204 23.756 0.276 23.788 ;
  LAYER M1 ;
        RECT 0.224 24.408 0.256 24.48 ;
  LAYER M2 ;
        RECT 0.204 24.428 0.276 24.46 ;
  LAYER M1 ;
        RECT 0.224 24.108 0.256 24.444 ;
  LAYER M1 ;
        RECT 0.224 3.192 0.256 24.108 ;
  LAYER M1 ;
        RECT 6.144 3.156 6.176 3.228 ;
  LAYER M2 ;
        RECT 6.124 3.176 6.196 3.208 ;
  LAYER M1 ;
        RECT 6.144 3.192 6.176 3.36 ;
  LAYER M1 ;
        RECT 6.144 3.324 6.176 3.396 ;
  LAYER M2 ;
        RECT 6.124 3.344 6.196 3.376 ;
  LAYER M2 ;
        RECT 6.16 3.344 8.88 3.376 ;
  LAYER M1 ;
        RECT 8.864 3.324 8.896 3.396 ;
  LAYER M2 ;
        RECT 8.844 3.344 8.916 3.376 ;
  LAYER M1 ;
        RECT 6.144 6.096 6.176 6.168 ;
  LAYER M2 ;
        RECT 6.124 6.116 6.196 6.148 ;
  LAYER M1 ;
        RECT 6.144 6.132 6.176 6.3 ;
  LAYER M1 ;
        RECT 6.144 6.264 6.176 6.336 ;
  LAYER M2 ;
        RECT 6.124 6.284 6.196 6.316 ;
  LAYER M2 ;
        RECT 6.16 6.284 8.88 6.316 ;
  LAYER M1 ;
        RECT 8.864 6.264 8.896 6.336 ;
  LAYER M2 ;
        RECT 8.844 6.284 8.916 6.316 ;
  LAYER M1 ;
        RECT 6.144 9.036 6.176 9.108 ;
  LAYER M2 ;
        RECT 6.124 9.056 6.196 9.088 ;
  LAYER M1 ;
        RECT 6.144 9.072 6.176 9.24 ;
  LAYER M1 ;
        RECT 6.144 9.204 6.176 9.276 ;
  LAYER M2 ;
        RECT 6.124 9.224 6.196 9.256 ;
  LAYER M2 ;
        RECT 6.16 9.224 8.88 9.256 ;
  LAYER M1 ;
        RECT 8.864 9.204 8.896 9.276 ;
  LAYER M2 ;
        RECT 8.844 9.224 8.916 9.256 ;
  LAYER M1 ;
        RECT 6.144 11.976 6.176 12.048 ;
  LAYER M2 ;
        RECT 6.124 11.996 6.196 12.028 ;
  LAYER M1 ;
        RECT 6.144 12.012 6.176 12.18 ;
  LAYER M1 ;
        RECT 6.144 12.144 6.176 12.216 ;
  LAYER M2 ;
        RECT 6.124 12.164 6.196 12.196 ;
  LAYER M2 ;
        RECT 6.16 12.164 8.88 12.196 ;
  LAYER M1 ;
        RECT 8.864 12.144 8.896 12.216 ;
  LAYER M2 ;
        RECT 8.844 12.164 8.916 12.196 ;
  LAYER M1 ;
        RECT 6.144 14.916 6.176 14.988 ;
  LAYER M2 ;
        RECT 6.124 14.936 6.196 14.968 ;
  LAYER M1 ;
        RECT 6.144 14.952 6.176 15.12 ;
  LAYER M1 ;
        RECT 6.144 15.084 6.176 15.156 ;
  LAYER M2 ;
        RECT 6.124 15.104 6.196 15.136 ;
  LAYER M2 ;
        RECT 6.16 15.104 8.88 15.136 ;
  LAYER M1 ;
        RECT 8.864 15.084 8.896 15.156 ;
  LAYER M2 ;
        RECT 8.844 15.104 8.916 15.136 ;
  LAYER M1 ;
        RECT 6.144 17.856 6.176 17.928 ;
  LAYER M2 ;
        RECT 6.124 17.876 6.196 17.908 ;
  LAYER M1 ;
        RECT 6.144 17.892 6.176 18.06 ;
  LAYER M1 ;
        RECT 6.144 18.024 6.176 18.096 ;
  LAYER M2 ;
        RECT 6.124 18.044 6.196 18.076 ;
  LAYER M2 ;
        RECT 6.16 18.044 8.88 18.076 ;
  LAYER M1 ;
        RECT 8.864 18.024 8.896 18.096 ;
  LAYER M2 ;
        RECT 8.844 18.044 8.916 18.076 ;
  LAYER M1 ;
        RECT 6.144 20.796 6.176 20.868 ;
  LAYER M2 ;
        RECT 6.124 20.816 6.196 20.848 ;
  LAYER M1 ;
        RECT 6.144 20.832 6.176 21 ;
  LAYER M1 ;
        RECT 6.144 20.964 6.176 21.036 ;
  LAYER M2 ;
        RECT 6.124 20.984 6.196 21.016 ;
  LAYER M2 ;
        RECT 6.16 20.984 8.88 21.016 ;
  LAYER M1 ;
        RECT 8.864 20.964 8.896 21.036 ;
  LAYER M2 ;
        RECT 8.844 20.984 8.916 21.016 ;
  LAYER M1 ;
        RECT 6.144 23.736 6.176 23.808 ;
  LAYER M2 ;
        RECT 6.124 23.756 6.196 23.788 ;
  LAYER M1 ;
        RECT 6.144 23.772 6.176 23.94 ;
  LAYER M1 ;
        RECT 6.144 23.904 6.176 23.976 ;
  LAYER M2 ;
        RECT 6.124 23.924 6.196 23.956 ;
  LAYER M2 ;
        RECT 6.16 23.924 8.88 23.956 ;
  LAYER M1 ;
        RECT 8.864 23.904 8.896 23.976 ;
  LAYER M2 ;
        RECT 8.844 23.924 8.916 23.956 ;
  LAYER M1 ;
        RECT 8.864 24.408 8.896 24.48 ;
  LAYER M2 ;
        RECT 8.844 24.428 8.916 24.46 ;
  LAYER M1 ;
        RECT 8.864 24.108 8.896 24.444 ;
  LAYER M1 ;
        RECT 8.864 3.36 8.896 24.108 ;
  LAYER M2 ;
        RECT 0.24 24.428 8.88 24.46 ;
  LAYER M1 ;
        RECT 3.264 3.156 3.296 3.228 ;
  LAYER M2 ;
        RECT 3.244 3.176 3.316 3.208 ;
  LAYER M2 ;
        RECT 0.4 3.176 3.28 3.208 ;
  LAYER M1 ;
        RECT 0.384 3.156 0.416 3.228 ;
  LAYER M2 ;
        RECT 0.364 3.176 0.436 3.208 ;
  LAYER M1 ;
        RECT 3.264 23.736 3.296 23.808 ;
  LAYER M2 ;
        RECT 3.244 23.756 3.316 23.788 ;
  LAYER M2 ;
        RECT 0.4 23.756 3.28 23.788 ;
  LAYER M1 ;
        RECT 0.384 23.736 0.416 23.808 ;
  LAYER M2 ;
        RECT 0.364 23.756 0.436 23.788 ;
  LAYER M1 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M2 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M3 ;
        RECT 0.4 0.756 2.8 3.192 ;
  LAYER M1 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M2 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M3 ;
        RECT 0.4 3.696 2.8 6.132 ;
  LAYER M1 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M2 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M3 ;
        RECT 0.4 6.636 2.8 9.072 ;
  LAYER M1 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M2 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M3 ;
        RECT 0.4 9.576 2.8 12.012 ;
  LAYER M1 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M2 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M3 ;
        RECT 0.4 12.516 2.8 14.952 ;
  LAYER M1 ;
        RECT 0.4 15.456 2.8 17.892 ;
  LAYER M2 ;
        RECT 0.4 15.456 2.8 17.892 ;
  LAYER M3 ;
        RECT 0.4 15.456 2.8 17.892 ;
  LAYER M1 ;
        RECT 0.4 18.396 2.8 20.832 ;
  LAYER M2 ;
        RECT 0.4 18.396 2.8 20.832 ;
  LAYER M3 ;
        RECT 0.4 18.396 2.8 20.832 ;
  LAYER M1 ;
        RECT 0.4 21.336 2.8 23.772 ;
  LAYER M2 ;
        RECT 0.4 21.336 2.8 23.772 ;
  LAYER M3 ;
        RECT 0.4 21.336 2.8 23.772 ;
  LAYER M1 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M2 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M3 ;
        RECT 3.28 0.756 5.68 3.192 ;
  LAYER M1 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M2 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M3 ;
        RECT 3.28 3.696 5.68 6.132 ;
  LAYER M1 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M2 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M3 ;
        RECT 3.28 6.636 5.68 9.072 ;
  LAYER M1 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M2 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M3 ;
        RECT 3.28 9.576 5.68 12.012 ;
  LAYER M1 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M2 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M3 ;
        RECT 3.28 12.516 5.68 14.952 ;
  LAYER M1 ;
        RECT 3.28 15.456 5.68 17.892 ;
  LAYER M2 ;
        RECT 3.28 15.456 5.68 17.892 ;
  LAYER M3 ;
        RECT 3.28 15.456 5.68 17.892 ;
  LAYER M1 ;
        RECT 3.28 18.396 5.68 20.832 ;
  LAYER M2 ;
        RECT 3.28 18.396 5.68 20.832 ;
  LAYER M3 ;
        RECT 3.28 18.396 5.68 20.832 ;
  LAYER M1 ;
        RECT 3.28 21.336 5.68 23.772 ;
  LAYER M2 ;
        RECT 3.28 21.336 5.68 23.772 ;
  LAYER M3 ;
        RECT 3.28 21.336 5.68 23.772 ;
  LAYER M1 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M2 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M3 ;
        RECT 6.16 0.756 8.56 3.192 ;
  LAYER M1 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M2 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M3 ;
        RECT 6.16 3.696 8.56 6.132 ;
  LAYER M1 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M2 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M3 ;
        RECT 6.16 6.636 8.56 9.072 ;
  LAYER M1 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M2 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M3 ;
        RECT 6.16 9.576 8.56 12.012 ;
  LAYER M1 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M2 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M3 ;
        RECT 6.16 12.516 8.56 14.952 ;
  LAYER M1 ;
        RECT 6.16 15.456 8.56 17.892 ;
  LAYER M2 ;
        RECT 6.16 15.456 8.56 17.892 ;
  LAYER M3 ;
        RECT 6.16 15.456 8.56 17.892 ;
  LAYER M1 ;
        RECT 6.16 18.396 8.56 20.832 ;
  LAYER M2 ;
        RECT 6.16 18.396 8.56 20.832 ;
  LAYER M3 ;
        RECT 6.16 18.396 8.56 20.832 ;
  LAYER M1 ;
        RECT 6.16 21.336 8.56 23.772 ;
  LAYER M2 ;
        RECT 6.16 21.336 8.56 23.772 ;
  LAYER M3 ;
        RECT 6.16 21.336 8.56 23.772 ;
  END 
END Cap_60fF
