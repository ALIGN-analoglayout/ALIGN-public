MACRO Cap_60fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF_Cap_60fF 0 0 ;
  SIZE 12.16 BY 26.208 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 25.752 3.232 25.824 ;
      LAYER M2 ;
        RECT 3.18 25.772 3.252 25.804 ;
      LAYER M1 ;
        RECT 9.152 25.752 9.184 25.824 ;
      LAYER M2 ;
        RECT 9.132 25.772 9.204 25.804 ;
      LAYER M2 ;
        RECT 3.216 25.772 9.168 25.804 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
      LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 25.92 6.208 25.992 ;
      LAYER M2 ;
        RECT 6.156 25.94 6.228 25.972 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
      LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
      LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
      LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
      LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 5.792 10.296 5.824 10.368 ;
  LAYER M2 ;
        RECT 5.772 10.316 5.844 10.348 ;
  LAYER M1 ;
        RECT 5.792 10.164 5.824 10.332 ;
  LAYER M1 ;
        RECT 5.792 10.128 5.824 10.2 ;
  LAYER M2 ;
        RECT 5.772 10.148 5.844 10.18 ;
  LAYER M2 ;
        RECT 5.808 10.148 6.032 10.18 ;
  LAYER M1 ;
        RECT 6.016 10.128 6.048 10.2 ;
  LAYER M2 ;
        RECT 5.996 10.148 6.068 10.18 ;
  LAYER M1 ;
        RECT 8.768 13.404 8.8 13.476 ;
  LAYER M2 ;
        RECT 8.748 13.424 8.82 13.456 ;
  LAYER M2 ;
        RECT 6.032 13.424 8.784 13.456 ;
  LAYER M1 ;
        RECT 6.016 13.404 6.048 13.476 ;
  LAYER M2 ;
        RECT 5.996 13.424 6.068 13.456 ;
  LAYER M1 ;
        RECT 5.792 13.404 5.824 13.476 ;
  LAYER M2 ;
        RECT 5.772 13.424 5.844 13.456 ;
  LAYER M1 ;
        RECT 5.792 13.272 5.824 13.44 ;
  LAYER M1 ;
        RECT 5.792 13.236 5.824 13.308 ;
  LAYER M2 ;
        RECT 5.772 13.256 5.844 13.288 ;
  LAYER M2 ;
        RECT 5.808 13.256 6.032 13.288 ;
  LAYER M1 ;
        RECT 6.016 13.236 6.048 13.308 ;
  LAYER M2 ;
        RECT 5.996 13.256 6.068 13.288 ;
  LAYER M1 ;
        RECT 8.768 10.296 8.8 10.368 ;
  LAYER M2 ;
        RECT 8.748 10.316 8.82 10.348 ;
  LAYER M2 ;
        RECT 6.032 10.316 8.784 10.348 ;
  LAYER M1 ;
        RECT 6.016 10.296 6.048 10.368 ;
  LAYER M2 ;
        RECT 5.996 10.316 6.068 10.348 ;
  LAYER M1 ;
        RECT 5.792 16.512 5.824 16.584 ;
  LAYER M2 ;
        RECT 5.772 16.532 5.844 16.564 ;
  LAYER M1 ;
        RECT 5.792 16.38 5.824 16.548 ;
  LAYER M1 ;
        RECT 5.792 16.344 5.824 16.416 ;
  LAYER M2 ;
        RECT 5.772 16.364 5.844 16.396 ;
  LAYER M2 ;
        RECT 5.808 16.364 6.032 16.396 ;
  LAYER M1 ;
        RECT 6.016 16.344 6.048 16.416 ;
  LAYER M2 ;
        RECT 5.996 16.364 6.068 16.396 ;
  LAYER M1 ;
        RECT 8.768 7.188 8.8 7.26 ;
  LAYER M2 ;
        RECT 8.748 7.208 8.82 7.24 ;
  LAYER M2 ;
        RECT 6.032 7.208 8.784 7.24 ;
  LAYER M1 ;
        RECT 6.016 7.188 6.048 7.26 ;
  LAYER M2 ;
        RECT 5.996 7.208 6.068 7.24 ;
  LAYER M1 ;
        RECT 6.016 0.384 6.048 0.456 ;
  LAYER M2 ;
        RECT 5.996 0.404 6.068 0.436 ;
  LAYER M1 ;
        RECT 6.016 0.42 6.048 0.672 ;
  LAYER M1 ;
        RECT 6.016 0.672 6.048 16.38 ;
  LAYER M1 ;
        RECT 5.792 7.188 5.824 7.26 ;
  LAYER M2 ;
        RECT 5.772 7.208 5.844 7.24 ;
  LAYER M2 ;
        RECT 3.056 7.208 5.808 7.24 ;
  LAYER M1 ;
        RECT 3.04 7.188 3.072 7.26 ;
  LAYER M2 ;
        RECT 3.02 7.208 3.092 7.24 ;
  LAYER M1 ;
        RECT 5.792 19.62 5.824 19.692 ;
  LAYER M2 ;
        RECT 5.772 19.64 5.844 19.672 ;
  LAYER M2 ;
        RECT 3.056 19.64 5.808 19.672 ;
  LAYER M1 ;
        RECT 3.04 19.62 3.072 19.692 ;
  LAYER M2 ;
        RECT 3.02 19.64 3.092 19.672 ;
  LAYER M1 ;
        RECT 5.792 4.08 5.824 4.152 ;
  LAYER M2 ;
        RECT 5.772 4.1 5.844 4.132 ;
  LAYER M2 ;
        RECT 3.056 4.1 5.808 4.132 ;
  LAYER M1 ;
        RECT 3.04 4.08 3.072 4.152 ;
  LAYER M2 ;
        RECT 3.02 4.1 3.092 4.132 ;
  LAYER M1 ;
        RECT 3.04 0.216 3.072 0.288 ;
  LAYER M2 ;
        RECT 3.02 0.236 3.092 0.268 ;
  LAYER M1 ;
        RECT 3.04 0.252 3.072 0.672 ;
  LAYER M1 ;
        RECT 3.04 0.672 3.072 19.656 ;
  LAYER M1 ;
        RECT 8.768 16.512 8.8 16.584 ;
  LAYER M2 ;
        RECT 8.748 16.532 8.82 16.564 ;
  LAYER M1 ;
        RECT 8.768 16.38 8.8 16.548 ;
  LAYER M1 ;
        RECT 8.768 16.344 8.8 16.416 ;
  LAYER M2 ;
        RECT 8.748 16.364 8.82 16.396 ;
  LAYER M2 ;
        RECT 8.784 16.364 9.008 16.396 ;
  LAYER M1 ;
        RECT 8.992 16.344 9.024 16.416 ;
  LAYER M2 ;
        RECT 8.972 16.364 9.044 16.396 ;
  LAYER M1 ;
        RECT 8.768 4.08 8.8 4.152 ;
  LAYER M2 ;
        RECT 8.748 4.1 8.82 4.132 ;
  LAYER M1 ;
        RECT 8.768 3.948 8.8 4.116 ;
  LAYER M1 ;
        RECT 8.768 3.912 8.8 3.984 ;
  LAYER M2 ;
        RECT 8.748 3.932 8.82 3.964 ;
  LAYER M2 ;
        RECT 8.784 3.932 9.008 3.964 ;
  LAYER M1 ;
        RECT 8.992 3.912 9.024 3.984 ;
  LAYER M2 ;
        RECT 8.972 3.932 9.044 3.964 ;
  LAYER M1 ;
        RECT 8.768 19.62 8.8 19.692 ;
  LAYER M2 ;
        RECT 8.748 19.64 8.82 19.672 ;
  LAYER M1 ;
        RECT 8.768 19.488 8.8 19.656 ;
  LAYER M1 ;
        RECT 8.768 19.452 8.8 19.524 ;
  LAYER M2 ;
        RECT 8.748 19.472 8.82 19.504 ;
  LAYER M2 ;
        RECT 8.784 19.472 9.008 19.504 ;
  LAYER M1 ;
        RECT 8.992 19.452 9.024 19.524 ;
  LAYER M2 ;
        RECT 8.972 19.472 9.044 19.504 ;
  LAYER M1 ;
        RECT 8.992 0.216 9.024 0.288 ;
  LAYER M2 ;
        RECT 8.972 0.236 9.044 0.268 ;
  LAYER M1 ;
        RECT 8.992 0.252 9.024 0.672 ;
  LAYER M1 ;
        RECT 8.992 0.672 9.024 19.488 ;
  LAYER M2 ;
        RECT 3.056 0.236 9.008 0.268 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 2.832 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 2.816 4.08 2.848 4.152 ;
  LAYER M2 ;
        RECT 2.796 4.1 2.868 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 2.832 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 2.816 7.188 2.848 7.26 ;
  LAYER M2 ;
        RECT 2.796 7.208 2.868 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 2.832 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 2.816 10.296 2.848 10.368 ;
  LAYER M2 ;
        RECT 2.796 10.316 2.868 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 2.832 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 2.816 13.404 2.848 13.476 ;
  LAYER M2 ;
        RECT 2.796 13.424 2.868 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 2.832 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 2.816 16.512 2.848 16.584 ;
  LAYER M2 ;
        RECT 2.796 16.532 2.868 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 2.832 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 2.816 19.62 2.848 19.692 ;
  LAYER M2 ;
        RECT 2.796 19.64 2.868 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 2.832 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 2.816 22.728 2.848 22.8 ;
  LAYER M2 ;
        RECT 2.796 22.748 2.868 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 2.832 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 22.764 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.84 11.776 1.008 ;
  LAYER M1 ;
        RECT 11.744 0.804 11.776 0.876 ;
  LAYER M2 ;
        RECT 11.724 0.824 11.796 0.856 ;
  LAYER M2 ;
        RECT 11.76 0.824 11.984 0.856 ;
  LAYER M1 ;
        RECT 11.968 0.804 12 0.876 ;
  LAYER M2 ;
        RECT 11.948 0.824 12.02 0.856 ;
  LAYER M1 ;
        RECT 11.744 4.08 11.776 4.152 ;
  LAYER M2 ;
        RECT 11.724 4.1 11.796 4.132 ;
  LAYER M1 ;
        RECT 11.744 3.948 11.776 4.116 ;
  LAYER M1 ;
        RECT 11.744 3.912 11.776 3.984 ;
  LAYER M2 ;
        RECT 11.724 3.932 11.796 3.964 ;
  LAYER M2 ;
        RECT 11.76 3.932 11.984 3.964 ;
  LAYER M1 ;
        RECT 11.968 3.912 12 3.984 ;
  LAYER M2 ;
        RECT 11.948 3.932 12.02 3.964 ;
  LAYER M1 ;
        RECT 11.744 7.188 11.776 7.26 ;
  LAYER M2 ;
        RECT 11.724 7.208 11.796 7.24 ;
  LAYER M1 ;
        RECT 11.744 7.056 11.776 7.224 ;
  LAYER M1 ;
        RECT 11.744 7.02 11.776 7.092 ;
  LAYER M2 ;
        RECT 11.724 7.04 11.796 7.072 ;
  LAYER M2 ;
        RECT 11.76 7.04 11.984 7.072 ;
  LAYER M1 ;
        RECT 11.968 7.02 12 7.092 ;
  LAYER M2 ;
        RECT 11.948 7.04 12.02 7.072 ;
  LAYER M1 ;
        RECT 11.744 10.296 11.776 10.368 ;
  LAYER M2 ;
        RECT 11.724 10.316 11.796 10.348 ;
  LAYER M1 ;
        RECT 11.744 10.164 11.776 10.332 ;
  LAYER M1 ;
        RECT 11.744 10.128 11.776 10.2 ;
  LAYER M2 ;
        RECT 11.724 10.148 11.796 10.18 ;
  LAYER M2 ;
        RECT 11.76 10.148 11.984 10.18 ;
  LAYER M1 ;
        RECT 11.968 10.128 12 10.2 ;
  LAYER M2 ;
        RECT 11.948 10.148 12.02 10.18 ;
  LAYER M1 ;
        RECT 11.744 13.404 11.776 13.476 ;
  LAYER M2 ;
        RECT 11.724 13.424 11.796 13.456 ;
  LAYER M1 ;
        RECT 11.744 13.272 11.776 13.44 ;
  LAYER M1 ;
        RECT 11.744 13.236 11.776 13.308 ;
  LAYER M2 ;
        RECT 11.724 13.256 11.796 13.288 ;
  LAYER M2 ;
        RECT 11.76 13.256 11.984 13.288 ;
  LAYER M1 ;
        RECT 11.968 13.236 12 13.308 ;
  LAYER M2 ;
        RECT 11.948 13.256 12.02 13.288 ;
  LAYER M1 ;
        RECT 11.744 16.512 11.776 16.584 ;
  LAYER M2 ;
        RECT 11.724 16.532 11.796 16.564 ;
  LAYER M1 ;
        RECT 11.744 16.38 11.776 16.548 ;
  LAYER M1 ;
        RECT 11.744 16.344 11.776 16.416 ;
  LAYER M2 ;
        RECT 11.724 16.364 11.796 16.396 ;
  LAYER M2 ;
        RECT 11.76 16.364 11.984 16.396 ;
  LAYER M1 ;
        RECT 11.968 16.344 12 16.416 ;
  LAYER M2 ;
        RECT 11.948 16.364 12.02 16.396 ;
  LAYER M1 ;
        RECT 11.744 19.62 11.776 19.692 ;
  LAYER M2 ;
        RECT 11.724 19.64 11.796 19.672 ;
  LAYER M1 ;
        RECT 11.744 19.488 11.776 19.656 ;
  LAYER M1 ;
        RECT 11.744 19.452 11.776 19.524 ;
  LAYER M2 ;
        RECT 11.724 19.472 11.796 19.504 ;
  LAYER M2 ;
        RECT 11.76 19.472 11.984 19.504 ;
  LAYER M1 ;
        RECT 11.968 19.452 12 19.524 ;
  LAYER M2 ;
        RECT 11.948 19.472 12.02 19.504 ;
  LAYER M1 ;
        RECT 11.744 22.728 11.776 22.8 ;
  LAYER M2 ;
        RECT 11.724 22.748 11.796 22.78 ;
  LAYER M1 ;
        RECT 11.744 22.596 11.776 22.764 ;
  LAYER M1 ;
        RECT 11.744 22.56 11.776 22.632 ;
  LAYER M2 ;
        RECT 11.724 22.58 11.796 22.612 ;
  LAYER M2 ;
        RECT 11.76 22.58 11.984 22.612 ;
  LAYER M1 ;
        RECT 11.968 22.56 12 22.632 ;
  LAYER M2 ;
        RECT 11.948 22.58 12.02 22.612 ;
  LAYER M1 ;
        RECT 11.968 0.048 12 0.12 ;
  LAYER M2 ;
        RECT 11.948 0.068 12.02 0.1 ;
  LAYER M1 ;
        RECT 11.968 0.084 12 0.672 ;
  LAYER M1 ;
        RECT 11.968 0.672 12 22.596 ;
  LAYER M2 ;
        RECT 0.08 0.068 11.984 0.1 ;
  LAYER M1 ;
        RECT 5.792 0.972 5.824 1.044 ;
  LAYER M2 ;
        RECT 5.772 0.992 5.844 1.024 ;
  LAYER M2 ;
        RECT 2.832 0.992 5.808 1.024 ;
  LAYER M1 ;
        RECT 2.816 0.972 2.848 1.044 ;
  LAYER M2 ;
        RECT 2.796 0.992 2.868 1.024 ;
  LAYER M1 ;
        RECT 5.792 22.728 5.824 22.8 ;
  LAYER M2 ;
        RECT 5.772 22.748 5.844 22.78 ;
  LAYER M2 ;
        RECT 2.832 22.748 5.808 22.78 ;
  LAYER M1 ;
        RECT 2.816 22.728 2.848 22.8 ;
  LAYER M2 ;
        RECT 2.796 22.748 2.868 22.78 ;
  LAYER M1 ;
        RECT 8.768 22.728 8.8 22.8 ;
  LAYER M2 ;
        RECT 8.748 22.748 8.82 22.78 ;
  LAYER M2 ;
        RECT 5.808 22.748 8.784 22.78 ;
  LAYER M1 ;
        RECT 5.792 22.728 5.824 22.8 ;
  LAYER M2 ;
        RECT 5.772 22.748 5.844 22.78 ;
  LAYER M1 ;
        RECT 8.768 0.972 8.8 1.044 ;
  LAYER M2 ;
        RECT 8.748 0.992 8.82 1.024 ;
  LAYER M2 ;
        RECT 8.784 0.992 11.76 1.024 ;
  LAYER M1 ;
        RECT 11.744 0.972 11.776 1.044 ;
  LAYER M2 ;
        RECT 11.724 0.992 11.796 1.024 ;
  LAYER M1 ;
        RECT 3.424 12.732 3.456 12.804 ;
  LAYER M2 ;
        RECT 3.404 12.752 3.476 12.784 ;
  LAYER M2 ;
        RECT 3.216 12.752 3.44 12.784 ;
  LAYER M1 ;
        RECT 3.2 12.732 3.232 12.804 ;
  LAYER M2 ;
        RECT 3.18 12.752 3.252 12.784 ;
  LAYER M1 ;
        RECT 3.424 15.84 3.456 15.912 ;
  LAYER M2 ;
        RECT 3.404 15.86 3.476 15.892 ;
  LAYER M2 ;
        RECT 3.216 15.86 3.44 15.892 ;
  LAYER M1 ;
        RECT 3.2 15.84 3.232 15.912 ;
  LAYER M2 ;
        RECT 3.18 15.86 3.252 15.892 ;
  LAYER M1 ;
        RECT 3.424 18.948 3.456 19.02 ;
  LAYER M2 ;
        RECT 3.404 18.968 3.476 19 ;
  LAYER M2 ;
        RECT 3.216 18.968 3.44 19 ;
  LAYER M1 ;
        RECT 3.2 18.948 3.232 19.02 ;
  LAYER M2 ;
        RECT 3.18 18.968 3.252 19 ;
  LAYER M1 ;
        RECT 3.2 25.752 3.232 25.824 ;
  LAYER M2 ;
        RECT 3.18 25.772 3.252 25.804 ;
  LAYER M1 ;
        RECT 3.2 25.536 3.232 25.788 ;
  LAYER M1 ;
        RECT 3.2 12.768 3.232 25.536 ;
  LAYER M1 ;
        RECT 6.4 15.84 6.432 15.912 ;
  LAYER M2 ;
        RECT 6.38 15.86 6.452 15.892 ;
  LAYER M1 ;
        RECT 6.4 15.876 6.432 16.044 ;
  LAYER M1 ;
        RECT 6.4 16.008 6.432 16.08 ;
  LAYER M2 ;
        RECT 6.38 16.028 6.452 16.06 ;
  LAYER M2 ;
        RECT 6.416 16.028 9.168 16.06 ;
  LAYER M1 ;
        RECT 9.152 16.008 9.184 16.08 ;
  LAYER M2 ;
        RECT 9.132 16.028 9.204 16.06 ;
  LAYER M1 ;
        RECT 6.4 12.732 6.432 12.804 ;
  LAYER M2 ;
        RECT 6.38 12.752 6.452 12.784 ;
  LAYER M1 ;
        RECT 6.4 12.768 6.432 12.936 ;
  LAYER M1 ;
        RECT 6.4 12.9 6.432 12.972 ;
  LAYER M2 ;
        RECT 6.38 12.92 6.452 12.952 ;
  LAYER M2 ;
        RECT 6.416 12.92 9.168 12.952 ;
  LAYER M1 ;
        RECT 9.152 12.9 9.184 12.972 ;
  LAYER M2 ;
        RECT 9.132 12.92 9.204 12.952 ;
  LAYER M1 ;
        RECT 6.4 9.624 6.432 9.696 ;
  LAYER M2 ;
        RECT 6.38 9.644 6.452 9.676 ;
  LAYER M1 ;
        RECT 6.4 9.66 6.432 9.828 ;
  LAYER M1 ;
        RECT 6.4 9.792 6.432 9.864 ;
  LAYER M2 ;
        RECT 6.38 9.812 6.452 9.844 ;
  LAYER M2 ;
        RECT 6.416 9.812 9.168 9.844 ;
  LAYER M1 ;
        RECT 9.152 9.792 9.184 9.864 ;
  LAYER M2 ;
        RECT 9.132 9.812 9.204 9.844 ;
  LAYER M1 ;
        RECT 9.152 25.752 9.184 25.824 ;
  LAYER M2 ;
        RECT 9.132 25.772 9.204 25.804 ;
  LAYER M1 ;
        RECT 9.152 25.536 9.184 25.788 ;
  LAYER M1 ;
        RECT 9.152 9.828 9.184 25.536 ;
  LAYER M2 ;
        RECT 3.216 25.772 9.168 25.804 ;
  LAYER M1 ;
        RECT 3.424 9.624 3.456 9.696 ;
  LAYER M2 ;
        RECT 3.404 9.644 3.476 9.676 ;
  LAYER M1 ;
        RECT 3.424 9.66 3.456 9.828 ;
  LAYER M1 ;
        RECT 3.424 9.792 3.456 9.864 ;
  LAYER M2 ;
        RECT 3.404 9.812 3.476 9.844 ;
  LAYER M2 ;
        RECT 3.44 9.812 6.192 9.844 ;
  LAYER M1 ;
        RECT 6.176 9.792 6.208 9.864 ;
  LAYER M2 ;
        RECT 6.156 9.812 6.228 9.844 ;
  LAYER M1 ;
        RECT 6.4 18.948 6.432 19.02 ;
  LAYER M2 ;
        RECT 6.38 18.968 6.452 19 ;
  LAYER M2 ;
        RECT 6.192 18.968 6.416 19 ;
  LAYER M1 ;
        RECT 6.176 18.948 6.208 19.02 ;
  LAYER M2 ;
        RECT 6.156 18.968 6.228 19 ;
  LAYER M1 ;
        RECT 3.424 22.056 3.456 22.128 ;
  LAYER M2 ;
        RECT 3.404 22.076 3.476 22.108 ;
  LAYER M1 ;
        RECT 3.424 22.092 3.456 22.26 ;
  LAYER M1 ;
        RECT 3.424 22.224 3.456 22.296 ;
  LAYER M2 ;
        RECT 3.404 22.244 3.476 22.276 ;
  LAYER M2 ;
        RECT 3.44 22.244 6.192 22.276 ;
  LAYER M1 ;
        RECT 6.176 22.224 6.208 22.296 ;
  LAYER M2 ;
        RECT 6.156 22.244 6.228 22.276 ;
  LAYER M1 ;
        RECT 6.4 6.516 6.432 6.588 ;
  LAYER M2 ;
        RECT 6.38 6.536 6.452 6.568 ;
  LAYER M2 ;
        RECT 6.192 6.536 6.416 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 3.424 6.516 3.456 6.588 ;
  LAYER M2 ;
        RECT 3.404 6.536 3.476 6.568 ;
  LAYER M1 ;
        RECT 3.424 6.552 3.456 6.72 ;
  LAYER M1 ;
        RECT 3.424 6.684 3.456 6.756 ;
  LAYER M2 ;
        RECT 3.404 6.704 3.476 6.736 ;
  LAYER M2 ;
        RECT 3.44 6.704 6.192 6.736 ;
  LAYER M1 ;
        RECT 6.176 6.684 6.208 6.756 ;
  LAYER M2 ;
        RECT 6.156 6.704 6.228 6.736 ;
  LAYER M1 ;
        RECT 6.4 22.056 6.432 22.128 ;
  LAYER M2 ;
        RECT 6.38 22.076 6.452 22.108 ;
  LAYER M2 ;
        RECT 6.192 22.076 6.416 22.108 ;
  LAYER M1 ;
        RECT 6.176 22.056 6.208 22.128 ;
  LAYER M2 ;
        RECT 6.156 22.076 6.228 22.108 ;
  LAYER M1 ;
        RECT 6.176 25.92 6.208 25.992 ;
  LAYER M2 ;
        RECT 6.156 25.94 6.228 25.972 ;
  LAYER M1 ;
        RECT 6.176 25.536 6.208 25.956 ;
  LAYER M1 ;
        RECT 6.176 6.552 6.208 25.536 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.464 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.448 6.516 0.48 6.588 ;
  LAYER M2 ;
        RECT 0.428 6.536 0.5 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.464 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.448 9.624 0.48 9.696 ;
  LAYER M2 ;
        RECT 0.428 9.644 0.5 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.464 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.448 12.732 0.48 12.804 ;
  LAYER M2 ;
        RECT 0.428 12.752 0.5 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.464 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.448 15.84 0.48 15.912 ;
  LAYER M2 ;
        RECT 0.428 15.86 0.5 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.464 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.448 18.948 0.48 19.02 ;
  LAYER M2 ;
        RECT 0.428 18.968 0.5 19 ;
  LAYER M2 ;
        RECT 0.24 18.968 0.464 19 ;
  LAYER M1 ;
        RECT 0.224 18.948 0.256 19.02 ;
  LAYER M2 ;
        RECT 0.204 18.968 0.276 19 ;
  LAYER M1 ;
        RECT 0.448 22.056 0.48 22.128 ;
  LAYER M2 ;
        RECT 0.428 22.076 0.5 22.108 ;
  LAYER M2 ;
        RECT 0.24 22.076 0.464 22.108 ;
  LAYER M1 ;
        RECT 0.224 22.056 0.256 22.128 ;
  LAYER M2 ;
        RECT 0.204 22.076 0.276 22.108 ;
  LAYER M1 ;
        RECT 0.448 25.164 0.48 25.236 ;
  LAYER M2 ;
        RECT 0.428 25.184 0.5 25.216 ;
  LAYER M2 ;
        RECT 0.24 25.184 0.464 25.216 ;
  LAYER M1 ;
        RECT 0.224 25.164 0.256 25.236 ;
  LAYER M2 ;
        RECT 0.204 25.184 0.276 25.216 ;
  LAYER M1 ;
        RECT 0.224 26.088 0.256 26.16 ;
  LAYER M2 ;
        RECT 0.204 26.108 0.276 26.14 ;
  LAYER M1 ;
        RECT 0.224 25.536 0.256 26.124 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 25.536 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.444 9.408 3.612 ;
  LAYER M1 ;
        RECT 9.376 3.576 9.408 3.648 ;
  LAYER M2 ;
        RECT 9.356 3.596 9.428 3.628 ;
  LAYER M2 ;
        RECT 9.392 3.596 12.144 3.628 ;
  LAYER M1 ;
        RECT 12.128 3.576 12.16 3.648 ;
  LAYER M2 ;
        RECT 12.108 3.596 12.18 3.628 ;
  LAYER M1 ;
        RECT 9.376 6.516 9.408 6.588 ;
  LAYER M2 ;
        RECT 9.356 6.536 9.428 6.568 ;
  LAYER M1 ;
        RECT 9.376 6.552 9.408 6.72 ;
  LAYER M1 ;
        RECT 9.376 6.684 9.408 6.756 ;
  LAYER M2 ;
        RECT 9.356 6.704 9.428 6.736 ;
  LAYER M2 ;
        RECT 9.392 6.704 12.144 6.736 ;
  LAYER M1 ;
        RECT 12.128 6.684 12.16 6.756 ;
  LAYER M2 ;
        RECT 12.108 6.704 12.18 6.736 ;
  LAYER M1 ;
        RECT 9.376 9.624 9.408 9.696 ;
  LAYER M2 ;
        RECT 9.356 9.644 9.428 9.676 ;
  LAYER M1 ;
        RECT 9.376 9.66 9.408 9.828 ;
  LAYER M1 ;
        RECT 9.376 9.792 9.408 9.864 ;
  LAYER M2 ;
        RECT 9.356 9.812 9.428 9.844 ;
  LAYER M2 ;
        RECT 9.392 9.812 12.144 9.844 ;
  LAYER M1 ;
        RECT 12.128 9.792 12.16 9.864 ;
  LAYER M2 ;
        RECT 12.108 9.812 12.18 9.844 ;
  LAYER M1 ;
        RECT 9.376 12.732 9.408 12.804 ;
  LAYER M2 ;
        RECT 9.356 12.752 9.428 12.784 ;
  LAYER M1 ;
        RECT 9.376 12.768 9.408 12.936 ;
  LAYER M1 ;
        RECT 9.376 12.9 9.408 12.972 ;
  LAYER M2 ;
        RECT 9.356 12.92 9.428 12.952 ;
  LAYER M2 ;
        RECT 9.392 12.92 12.144 12.952 ;
  LAYER M1 ;
        RECT 12.128 12.9 12.16 12.972 ;
  LAYER M2 ;
        RECT 12.108 12.92 12.18 12.952 ;
  LAYER M1 ;
        RECT 9.376 15.84 9.408 15.912 ;
  LAYER M2 ;
        RECT 9.356 15.86 9.428 15.892 ;
  LAYER M1 ;
        RECT 9.376 15.876 9.408 16.044 ;
  LAYER M1 ;
        RECT 9.376 16.008 9.408 16.08 ;
  LAYER M2 ;
        RECT 9.356 16.028 9.428 16.06 ;
  LAYER M2 ;
        RECT 9.392 16.028 12.144 16.06 ;
  LAYER M1 ;
        RECT 12.128 16.008 12.16 16.08 ;
  LAYER M2 ;
        RECT 12.108 16.028 12.18 16.06 ;
  LAYER M1 ;
        RECT 9.376 18.948 9.408 19.02 ;
  LAYER M2 ;
        RECT 9.356 18.968 9.428 19 ;
  LAYER M1 ;
        RECT 9.376 18.984 9.408 19.152 ;
  LAYER M1 ;
        RECT 9.376 19.116 9.408 19.188 ;
  LAYER M2 ;
        RECT 9.356 19.136 9.428 19.168 ;
  LAYER M2 ;
        RECT 9.392 19.136 12.144 19.168 ;
  LAYER M1 ;
        RECT 12.128 19.116 12.16 19.188 ;
  LAYER M2 ;
        RECT 12.108 19.136 12.18 19.168 ;
  LAYER M1 ;
        RECT 9.376 22.056 9.408 22.128 ;
  LAYER M2 ;
        RECT 9.356 22.076 9.428 22.108 ;
  LAYER M1 ;
        RECT 9.376 22.092 9.408 22.26 ;
  LAYER M1 ;
        RECT 9.376 22.224 9.408 22.296 ;
  LAYER M2 ;
        RECT 9.356 22.244 9.428 22.276 ;
  LAYER M2 ;
        RECT 9.392 22.244 12.144 22.276 ;
  LAYER M1 ;
        RECT 12.128 22.224 12.16 22.296 ;
  LAYER M2 ;
        RECT 12.108 22.244 12.18 22.276 ;
  LAYER M1 ;
        RECT 9.376 25.164 9.408 25.236 ;
  LAYER M2 ;
        RECT 9.356 25.184 9.428 25.216 ;
  LAYER M1 ;
        RECT 9.376 25.2 9.408 25.368 ;
  LAYER M1 ;
        RECT 9.376 25.332 9.408 25.404 ;
  LAYER M2 ;
        RECT 9.356 25.352 9.428 25.384 ;
  LAYER M2 ;
        RECT 9.392 25.352 12.144 25.384 ;
  LAYER M1 ;
        RECT 12.128 25.332 12.16 25.404 ;
  LAYER M2 ;
        RECT 12.108 25.352 12.18 25.384 ;
  LAYER M1 ;
        RECT 12.128 26.088 12.16 26.16 ;
  LAYER M2 ;
        RECT 12.108 26.108 12.18 26.14 ;
  LAYER M1 ;
        RECT 12.128 25.536 12.16 26.124 ;
  LAYER M1 ;
        RECT 12.128 3.612 12.16 25.536 ;
  LAYER M2 ;
        RECT 0.24 26.108 12.144 26.14 ;
  LAYER M1 ;
        RECT 3.424 3.408 3.456 3.48 ;
  LAYER M2 ;
        RECT 3.404 3.428 3.476 3.46 ;
  LAYER M2 ;
        RECT 0.464 3.428 3.44 3.46 ;
  LAYER M1 ;
        RECT 0.448 3.408 0.48 3.48 ;
  LAYER M2 ;
        RECT 0.428 3.428 0.5 3.46 ;
  LAYER M1 ;
        RECT 3.424 25.164 3.456 25.236 ;
  LAYER M2 ;
        RECT 3.404 25.184 3.476 25.216 ;
  LAYER M2 ;
        RECT 0.464 25.184 3.44 25.216 ;
  LAYER M1 ;
        RECT 0.448 25.164 0.48 25.236 ;
  LAYER M2 ;
        RECT 0.428 25.184 0.5 25.216 ;
  LAYER M1 ;
        RECT 6.4 25.164 6.432 25.236 ;
  LAYER M2 ;
        RECT 6.38 25.184 6.452 25.216 ;
  LAYER M2 ;
        RECT 3.44 25.184 6.416 25.216 ;
  LAYER M1 ;
        RECT 3.424 25.164 3.456 25.236 ;
  LAYER M2 ;
        RECT 3.404 25.184 3.476 25.216 ;
  LAYER M1 ;
        RECT 6.4 3.408 6.432 3.48 ;
  LAYER M2 ;
        RECT 6.38 3.428 6.452 3.46 ;
  LAYER M2 ;
        RECT 6.416 3.428 9.392 3.46 ;
  LAYER M1 ;
        RECT 9.376 3.408 9.408 3.48 ;
  LAYER M2 ;
        RECT 9.356 3.428 9.428 3.46 ;
  LAYER M1 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M3 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M2 ;
        RECT 0.4 0.924 2.896 3.528 ;
  LAYER M1 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M3 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M2 ;
        RECT 0.4 4.032 2.896 6.636 ;
  LAYER M1 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M3 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M2 ;
        RECT 0.4 7.14 2.896 9.744 ;
  LAYER M1 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M3 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M2 ;
        RECT 0.4 10.248 2.896 12.852 ;
  LAYER M1 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M3 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M2 ;
        RECT 0.4 13.356 2.896 15.96 ;
  LAYER M1 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M3 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M2 ;
        RECT 0.4 16.464 2.896 19.068 ;
  LAYER M1 ;
        RECT 0.4 19.572 2.896 22.176 ;
  LAYER M3 ;
        RECT 0.4 19.572 2.896 22.176 ;
  LAYER M2 ;
        RECT 0.4 19.572 2.896 22.176 ;
  LAYER M1 ;
        RECT 0.4 22.68 2.896 25.284 ;
  LAYER M3 ;
        RECT 0.4 22.68 2.896 25.284 ;
  LAYER M2 ;
        RECT 0.4 22.68 2.896 25.284 ;
  LAYER M1 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M3 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M2 ;
        RECT 3.376 0.924 5.872 3.528 ;
  LAYER M1 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M3 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M2 ;
        RECT 3.376 4.032 5.872 6.636 ;
  LAYER M1 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M3 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M2 ;
        RECT 3.376 7.14 5.872 9.744 ;
  LAYER M1 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M3 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M2 ;
        RECT 3.376 10.248 5.872 12.852 ;
  LAYER M1 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M3 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M2 ;
        RECT 3.376 13.356 5.872 15.96 ;
  LAYER M1 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M3 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M2 ;
        RECT 3.376 16.464 5.872 19.068 ;
  LAYER M1 ;
        RECT 3.376 19.572 5.872 22.176 ;
  LAYER M3 ;
        RECT 3.376 19.572 5.872 22.176 ;
  LAYER M2 ;
        RECT 3.376 19.572 5.872 22.176 ;
  LAYER M1 ;
        RECT 3.376 22.68 5.872 25.284 ;
  LAYER M3 ;
        RECT 3.376 22.68 5.872 25.284 ;
  LAYER M2 ;
        RECT 3.376 22.68 5.872 25.284 ;
  LAYER M1 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M3 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M2 ;
        RECT 6.352 0.924 8.848 3.528 ;
  LAYER M1 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M3 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M2 ;
        RECT 6.352 4.032 8.848 6.636 ;
  LAYER M1 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M3 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M2 ;
        RECT 6.352 7.14 8.848 9.744 ;
  LAYER M1 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M3 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M2 ;
        RECT 6.352 10.248 8.848 12.852 ;
  LAYER M1 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M3 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M2 ;
        RECT 6.352 13.356 8.848 15.96 ;
  LAYER M1 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M3 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M2 ;
        RECT 6.352 16.464 8.848 19.068 ;
  LAYER M1 ;
        RECT 6.352 19.572 8.848 22.176 ;
  LAYER M3 ;
        RECT 6.352 19.572 8.848 22.176 ;
  LAYER M2 ;
        RECT 6.352 19.572 8.848 22.176 ;
  LAYER M1 ;
        RECT 6.352 22.68 8.848 25.284 ;
  LAYER M3 ;
        RECT 6.352 22.68 8.848 25.284 ;
  LAYER M2 ;
        RECT 6.352 22.68 8.848 25.284 ;
  LAYER M1 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M3 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M2 ;
        RECT 9.328 0.924 11.824 3.528 ;
  LAYER M1 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M3 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M2 ;
        RECT 9.328 4.032 11.824 6.636 ;
  LAYER M1 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M3 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M2 ;
        RECT 9.328 7.14 11.824 9.744 ;
  LAYER M1 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M3 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M2 ;
        RECT 9.328 10.248 11.824 12.852 ;
  LAYER M1 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M3 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M2 ;
        RECT 9.328 13.356 11.824 15.96 ;
  LAYER M1 ;
        RECT 9.328 16.464 11.824 19.068 ;
  LAYER M3 ;
        RECT 9.328 16.464 11.824 19.068 ;
  LAYER M2 ;
        RECT 9.328 16.464 11.824 19.068 ;
  LAYER M1 ;
        RECT 9.328 19.572 11.824 22.176 ;
  LAYER M3 ;
        RECT 9.328 19.572 11.824 22.176 ;
  LAYER M2 ;
        RECT 9.328 19.572 11.824 22.176 ;
  LAYER M1 ;
        RECT 9.328 22.68 11.824 25.284 ;
  LAYER M3 ;
        RECT 9.328 22.68 11.824 25.284 ;
  LAYER M2 ;
        RECT 9.328 22.68 11.824 25.284 ;
  END 
END Cap_60fF_Cap_60fF
