MACRO Cap_30fF_Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_30fF_Cap_60fF 0 0 ;
  SIZE 10.16 BY 35.532 ;
  PIN MINUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.68 35.076 3.712 35.148 ;
      LAYER M2 ;
        RECT 3.66 35.096 3.732 35.128 ;
      LAYER M1 ;
        RECT 6.976 35.076 7.008 35.148 ;
      LAYER M2 ;
        RECT 6.956 35.096 7.028 35.128 ;
      LAYER M2 ;
        RECT 3.696 35.096 6.992 35.128 ;
    END
  END MINUS1
  PIN PLUS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
      LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
      LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
      LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
      LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
    END
  END PLUS1
  PIN MINUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.84 35.244 3.872 35.316 ;
      LAYER M2 ;
        RECT 3.82 35.264 3.892 35.296 ;
      LAYER M1 ;
        RECT 7.136 35.244 7.168 35.316 ;
      LAYER M2 ;
        RECT 7.116 35.264 7.188 35.296 ;
      LAYER M2 ;
        RECT 3.856 35.264 7.152 35.296 ;
    END
  END MINUS2
  PIN PLUS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
      LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
      LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
      LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
      LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
    END
  END PLUS2
  OBS 
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M2 ;
        RECT 3.376 16.532 6.448 16.564 ;
  LAYER M1 ;
        RECT 3.36 16.512 3.392 16.584 ;
  LAYER M2 ;
        RECT 3.34 16.532 3.412 16.564 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M2 ;
        RECT 3.376 4.1 6.448 4.132 ;
  LAYER M1 ;
        RECT 3.36 4.08 3.392 4.152 ;
  LAYER M2 ;
        RECT 3.34 4.1 3.412 4.132 ;
  LAYER M1 ;
        RECT 6.432 28.944 6.464 29.016 ;
  LAYER M2 ;
        RECT 6.412 28.964 6.484 28.996 ;
  LAYER M2 ;
        RECT 3.376 28.964 6.448 28.996 ;
  LAYER M1 ;
        RECT 3.36 28.944 3.392 29.016 ;
  LAYER M2 ;
        RECT 3.34 28.964 3.412 28.996 ;
  LAYER M1 ;
        RECT 3.36 0.384 3.392 0.456 ;
  LAYER M2 ;
        RECT 3.34 0.404 3.412 0.436 ;
  LAYER M1 ;
        RECT 3.36 0.42 3.392 0.672 ;
  LAYER M1 ;
        RECT 3.36 0.672 3.392 28.98 ;
  LAYER M1 ;
        RECT 6.432 16.512 6.464 16.584 ;
  LAYER M2 ;
        RECT 6.412 16.532 6.484 16.564 ;
  LAYER M1 ;
        RECT 6.432 16.38 6.464 16.548 ;
  LAYER M1 ;
        RECT 6.432 16.344 6.464 16.416 ;
  LAYER M2 ;
        RECT 6.412 16.364 6.484 16.396 ;
  LAYER M2 ;
        RECT 6.448 16.364 6.672 16.396 ;
  LAYER M1 ;
        RECT 6.656 16.344 6.688 16.416 ;
  LAYER M2 ;
        RECT 6.636 16.364 6.708 16.396 ;
  LAYER M1 ;
        RECT 6.432 4.08 6.464 4.152 ;
  LAYER M2 ;
        RECT 6.412 4.1 6.484 4.132 ;
  LAYER M1 ;
        RECT 6.432 3.948 6.464 4.116 ;
  LAYER M1 ;
        RECT 6.432 3.912 6.464 3.984 ;
  LAYER M2 ;
        RECT 6.412 3.932 6.484 3.964 ;
  LAYER M2 ;
        RECT 6.448 3.932 6.672 3.964 ;
  LAYER M1 ;
        RECT 6.656 3.912 6.688 3.984 ;
  LAYER M2 ;
        RECT 6.636 3.932 6.708 3.964 ;
  LAYER M1 ;
        RECT 6.432 28.944 6.464 29.016 ;
  LAYER M2 ;
        RECT 6.412 28.964 6.484 28.996 ;
  LAYER M1 ;
        RECT 6.432 28.812 6.464 28.98 ;
  LAYER M1 ;
        RECT 6.432 28.776 6.464 28.848 ;
  LAYER M2 ;
        RECT 6.412 28.796 6.484 28.828 ;
  LAYER M2 ;
        RECT 6.448 28.796 6.672 28.828 ;
  LAYER M1 ;
        RECT 6.656 28.776 6.688 28.848 ;
  LAYER M2 ;
        RECT 6.636 28.796 6.708 28.828 ;
  LAYER M1 ;
        RECT 6.656 0.384 6.688 0.456 ;
  LAYER M2 ;
        RECT 6.636 0.404 6.708 0.436 ;
  LAYER M1 ;
        RECT 6.656 0.42 6.688 0.672 ;
  LAYER M1 ;
        RECT 6.656 0.672 6.688 28.812 ;
  LAYER M2 ;
        RECT 3.376 0.404 6.672 0.436 ;
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M2 ;
        RECT 3.536 13.424 6.448 13.456 ;
  LAYER M1 ;
        RECT 3.52 13.404 3.552 13.476 ;
  LAYER M2 ;
        RECT 3.5 13.424 3.572 13.456 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M2 ;
        RECT 3.536 19.64 6.448 19.672 ;
  LAYER M1 ;
        RECT 3.52 19.62 3.552 19.692 ;
  LAYER M2 ;
        RECT 3.5 19.64 3.572 19.672 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M2 ;
        RECT 3.536 10.316 6.448 10.348 ;
  LAYER M1 ;
        RECT 3.52 10.296 3.552 10.368 ;
  LAYER M2 ;
        RECT 3.5 10.316 3.572 10.348 ;
  LAYER M1 ;
        RECT 6.432 22.728 6.464 22.8 ;
  LAYER M2 ;
        RECT 6.412 22.748 6.484 22.78 ;
  LAYER M2 ;
        RECT 3.536 22.748 6.448 22.78 ;
  LAYER M1 ;
        RECT 3.52 22.728 3.552 22.8 ;
  LAYER M2 ;
        RECT 3.5 22.748 3.572 22.78 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M2 ;
        RECT 3.536 7.208 6.448 7.24 ;
  LAYER M1 ;
        RECT 3.52 7.188 3.552 7.26 ;
  LAYER M2 ;
        RECT 3.5 7.208 3.572 7.24 ;
  LAYER M1 ;
        RECT 6.432 25.836 6.464 25.908 ;
  LAYER M2 ;
        RECT 6.412 25.856 6.484 25.888 ;
  LAYER M2 ;
        RECT 3.536 25.856 6.448 25.888 ;
  LAYER M1 ;
        RECT 3.52 25.836 3.552 25.908 ;
  LAYER M2 ;
        RECT 3.5 25.856 3.572 25.888 ;
  LAYER M1 ;
        RECT 3.52 0.216 3.552 0.288 ;
  LAYER M2 ;
        RECT 3.5 0.236 3.572 0.268 ;
  LAYER M1 ;
        RECT 3.52 0.252 3.552 0.672 ;
  LAYER M1 ;
        RECT 3.52 0.672 3.552 25.872 ;
  LAYER M1 ;
        RECT 6.432 13.404 6.464 13.476 ;
  LAYER M2 ;
        RECT 6.412 13.424 6.484 13.456 ;
  LAYER M1 ;
        RECT 6.432 13.272 6.464 13.44 ;
  LAYER M1 ;
        RECT 6.432 13.236 6.464 13.308 ;
  LAYER M2 ;
        RECT 6.412 13.256 6.484 13.288 ;
  LAYER M2 ;
        RECT 6.448 13.256 6.832 13.288 ;
  LAYER M1 ;
        RECT 6.816 13.236 6.848 13.308 ;
  LAYER M2 ;
        RECT 6.796 13.256 6.868 13.288 ;
  LAYER M1 ;
        RECT 6.432 19.62 6.464 19.692 ;
  LAYER M2 ;
        RECT 6.412 19.64 6.484 19.672 ;
  LAYER M1 ;
        RECT 6.432 19.488 6.464 19.656 ;
  LAYER M1 ;
        RECT 6.432 19.452 6.464 19.524 ;
  LAYER M2 ;
        RECT 6.412 19.472 6.484 19.504 ;
  LAYER M2 ;
        RECT 6.448 19.472 6.832 19.504 ;
  LAYER M1 ;
        RECT 6.816 19.452 6.848 19.524 ;
  LAYER M2 ;
        RECT 6.796 19.472 6.868 19.504 ;
  LAYER M1 ;
        RECT 6.432 10.296 6.464 10.368 ;
  LAYER M2 ;
        RECT 6.412 10.316 6.484 10.348 ;
  LAYER M1 ;
        RECT 6.432 10.164 6.464 10.332 ;
  LAYER M1 ;
        RECT 6.432 10.128 6.464 10.2 ;
  LAYER M2 ;
        RECT 6.412 10.148 6.484 10.18 ;
  LAYER M2 ;
        RECT 6.448 10.148 6.832 10.18 ;
  LAYER M1 ;
        RECT 6.816 10.128 6.848 10.2 ;
  LAYER M2 ;
        RECT 6.796 10.148 6.868 10.18 ;
  LAYER M1 ;
        RECT 6.432 22.728 6.464 22.8 ;
  LAYER M2 ;
        RECT 6.412 22.748 6.484 22.78 ;
  LAYER M1 ;
        RECT 6.432 22.596 6.464 22.764 ;
  LAYER M1 ;
        RECT 6.432 22.56 6.464 22.632 ;
  LAYER M2 ;
        RECT 6.412 22.58 6.484 22.612 ;
  LAYER M2 ;
        RECT 6.448 22.58 6.832 22.612 ;
  LAYER M1 ;
        RECT 6.816 22.56 6.848 22.632 ;
  LAYER M2 ;
        RECT 6.796 22.58 6.868 22.612 ;
  LAYER M1 ;
        RECT 6.432 7.188 6.464 7.26 ;
  LAYER M2 ;
        RECT 6.412 7.208 6.484 7.24 ;
  LAYER M1 ;
        RECT 6.432 7.056 6.464 7.224 ;
  LAYER M1 ;
        RECT 6.432 7.02 6.464 7.092 ;
  LAYER M2 ;
        RECT 6.412 7.04 6.484 7.072 ;
  LAYER M2 ;
        RECT 6.448 7.04 6.832 7.072 ;
  LAYER M1 ;
        RECT 6.816 7.02 6.848 7.092 ;
  LAYER M2 ;
        RECT 6.796 7.04 6.868 7.072 ;
  LAYER M1 ;
        RECT 6.432 25.836 6.464 25.908 ;
  LAYER M2 ;
        RECT 6.412 25.856 6.484 25.888 ;
  LAYER M1 ;
        RECT 6.432 25.704 6.464 25.872 ;
  LAYER M1 ;
        RECT 6.432 25.668 6.464 25.74 ;
  LAYER M2 ;
        RECT 6.412 25.688 6.484 25.72 ;
  LAYER M2 ;
        RECT 6.448 25.688 6.832 25.72 ;
  LAYER M1 ;
        RECT 6.816 25.668 6.848 25.74 ;
  LAYER M2 ;
        RECT 6.796 25.688 6.868 25.72 ;
  LAYER M1 ;
        RECT 6.816 0.216 6.848 0.288 ;
  LAYER M2 ;
        RECT 6.796 0.236 6.868 0.268 ;
  LAYER M1 ;
        RECT 6.816 0.252 6.848 0.672 ;
  LAYER M1 ;
        RECT 6.816 0.672 6.848 25.704 ;
  LAYER M2 ;
        RECT 3.536 0.236 6.832 0.268 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M2 ;
        RECT 0.08 0.992 3.152 1.024 ;
  LAYER M1 ;
        RECT 0.064 0.972 0.096 1.044 ;
  LAYER M2 ;
        RECT 0.044 0.992 0.116 1.024 ;
  LAYER M1 ;
        RECT 3.136 4.08 3.168 4.152 ;
  LAYER M2 ;
        RECT 3.116 4.1 3.188 4.132 ;
  LAYER M2 ;
        RECT 0.08 4.1 3.152 4.132 ;
  LAYER M1 ;
        RECT 0.064 4.08 0.096 4.152 ;
  LAYER M2 ;
        RECT 0.044 4.1 0.116 4.132 ;
  LAYER M1 ;
        RECT 3.136 7.188 3.168 7.26 ;
  LAYER M2 ;
        RECT 3.116 7.208 3.188 7.24 ;
  LAYER M2 ;
        RECT 0.08 7.208 3.152 7.24 ;
  LAYER M1 ;
        RECT 0.064 7.188 0.096 7.26 ;
  LAYER M2 ;
        RECT 0.044 7.208 0.116 7.24 ;
  LAYER M1 ;
        RECT 3.136 10.296 3.168 10.368 ;
  LAYER M2 ;
        RECT 3.116 10.316 3.188 10.348 ;
  LAYER M2 ;
        RECT 0.08 10.316 3.152 10.348 ;
  LAYER M1 ;
        RECT 0.064 10.296 0.096 10.368 ;
  LAYER M2 ;
        RECT 0.044 10.316 0.116 10.348 ;
  LAYER M1 ;
        RECT 3.136 13.404 3.168 13.476 ;
  LAYER M2 ;
        RECT 3.116 13.424 3.188 13.456 ;
  LAYER M2 ;
        RECT 0.08 13.424 3.152 13.456 ;
  LAYER M1 ;
        RECT 0.064 13.404 0.096 13.476 ;
  LAYER M2 ;
        RECT 0.044 13.424 0.116 13.456 ;
  LAYER M1 ;
        RECT 3.136 16.512 3.168 16.584 ;
  LAYER M2 ;
        RECT 3.116 16.532 3.188 16.564 ;
  LAYER M2 ;
        RECT 0.08 16.532 3.152 16.564 ;
  LAYER M1 ;
        RECT 0.064 16.512 0.096 16.584 ;
  LAYER M2 ;
        RECT 0.044 16.532 0.116 16.564 ;
  LAYER M1 ;
        RECT 3.136 19.62 3.168 19.692 ;
  LAYER M2 ;
        RECT 3.116 19.64 3.188 19.672 ;
  LAYER M2 ;
        RECT 0.08 19.64 3.152 19.672 ;
  LAYER M1 ;
        RECT 0.064 19.62 0.096 19.692 ;
  LAYER M2 ;
        RECT 0.044 19.64 0.116 19.672 ;
  LAYER M1 ;
        RECT 3.136 22.728 3.168 22.8 ;
  LAYER M2 ;
        RECT 3.116 22.748 3.188 22.78 ;
  LAYER M2 ;
        RECT 0.08 22.748 3.152 22.78 ;
  LAYER M1 ;
        RECT 0.064 22.728 0.096 22.8 ;
  LAYER M2 ;
        RECT 0.044 22.748 0.116 22.78 ;
  LAYER M1 ;
        RECT 3.136 25.836 3.168 25.908 ;
  LAYER M2 ;
        RECT 3.116 25.856 3.188 25.888 ;
  LAYER M2 ;
        RECT 0.08 25.856 3.152 25.888 ;
  LAYER M1 ;
        RECT 0.064 25.836 0.096 25.908 ;
  LAYER M2 ;
        RECT 0.044 25.856 0.116 25.888 ;
  LAYER M1 ;
        RECT 3.136 28.944 3.168 29.016 ;
  LAYER M2 ;
        RECT 3.116 28.964 3.188 28.996 ;
  LAYER M2 ;
        RECT 0.08 28.964 3.152 28.996 ;
  LAYER M1 ;
        RECT 0.064 28.944 0.096 29.016 ;
  LAYER M2 ;
        RECT 0.044 28.964 0.116 28.996 ;
  LAYER M1 ;
        RECT 3.136 32.052 3.168 32.124 ;
  LAYER M2 ;
        RECT 3.116 32.072 3.188 32.104 ;
  LAYER M2 ;
        RECT 0.08 32.072 3.152 32.104 ;
  LAYER M1 ;
        RECT 0.064 32.052 0.096 32.124 ;
  LAYER M2 ;
        RECT 0.044 32.072 0.116 32.104 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 0.12 ;
  LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
  LAYER M1 ;
        RECT 0.064 0.084 0.096 0.672 ;
  LAYER M1 ;
        RECT 0.064 0.672 0.096 32.088 ;
  LAYER M1 ;
        RECT 9.728 0.972 9.76 1.044 ;
  LAYER M2 ;
        RECT 9.708 0.992 9.78 1.024 ;
  LAYER M1 ;
        RECT 9.728 0.84 9.76 1.008 ;
  LAYER M1 ;
        RECT 9.728 0.804 9.76 0.876 ;
  LAYER M2 ;
        RECT 9.708 0.824 9.78 0.856 ;
  LAYER M2 ;
        RECT 9.744 0.824 9.968 0.856 ;
  LAYER M1 ;
        RECT 9.952 0.804 9.984 0.876 ;
  LAYER M2 ;
        RECT 9.932 0.824 10.004 0.856 ;
  LAYER M1 ;
        RECT 9.728 4.08 9.76 4.152 ;
  LAYER M2 ;
        RECT 9.708 4.1 9.78 4.132 ;
  LAYER M1 ;
        RECT 9.728 3.948 9.76 4.116 ;
  LAYER M1 ;
        RECT 9.728 3.912 9.76 3.984 ;
  LAYER M2 ;
        RECT 9.708 3.932 9.78 3.964 ;
  LAYER M2 ;
        RECT 9.744 3.932 9.968 3.964 ;
  LAYER M1 ;
        RECT 9.952 3.912 9.984 3.984 ;
  LAYER M2 ;
        RECT 9.932 3.932 10.004 3.964 ;
  LAYER M1 ;
        RECT 9.728 7.188 9.76 7.26 ;
  LAYER M2 ;
        RECT 9.708 7.208 9.78 7.24 ;
  LAYER M1 ;
        RECT 9.728 7.056 9.76 7.224 ;
  LAYER M1 ;
        RECT 9.728 7.02 9.76 7.092 ;
  LAYER M2 ;
        RECT 9.708 7.04 9.78 7.072 ;
  LAYER M2 ;
        RECT 9.744 7.04 9.968 7.072 ;
  LAYER M1 ;
        RECT 9.952 7.02 9.984 7.092 ;
  LAYER M2 ;
        RECT 9.932 7.04 10.004 7.072 ;
  LAYER M1 ;
        RECT 9.728 10.296 9.76 10.368 ;
  LAYER M2 ;
        RECT 9.708 10.316 9.78 10.348 ;
  LAYER M1 ;
        RECT 9.728 10.164 9.76 10.332 ;
  LAYER M1 ;
        RECT 9.728 10.128 9.76 10.2 ;
  LAYER M2 ;
        RECT 9.708 10.148 9.78 10.18 ;
  LAYER M2 ;
        RECT 9.744 10.148 9.968 10.18 ;
  LAYER M1 ;
        RECT 9.952 10.128 9.984 10.2 ;
  LAYER M2 ;
        RECT 9.932 10.148 10.004 10.18 ;
  LAYER M1 ;
        RECT 9.728 13.404 9.76 13.476 ;
  LAYER M2 ;
        RECT 9.708 13.424 9.78 13.456 ;
  LAYER M1 ;
        RECT 9.728 13.272 9.76 13.44 ;
  LAYER M1 ;
        RECT 9.728 13.236 9.76 13.308 ;
  LAYER M2 ;
        RECT 9.708 13.256 9.78 13.288 ;
  LAYER M2 ;
        RECT 9.744 13.256 9.968 13.288 ;
  LAYER M1 ;
        RECT 9.952 13.236 9.984 13.308 ;
  LAYER M2 ;
        RECT 9.932 13.256 10.004 13.288 ;
  LAYER M1 ;
        RECT 9.728 16.512 9.76 16.584 ;
  LAYER M2 ;
        RECT 9.708 16.532 9.78 16.564 ;
  LAYER M1 ;
        RECT 9.728 16.38 9.76 16.548 ;
  LAYER M1 ;
        RECT 9.728 16.344 9.76 16.416 ;
  LAYER M2 ;
        RECT 9.708 16.364 9.78 16.396 ;
  LAYER M2 ;
        RECT 9.744 16.364 9.968 16.396 ;
  LAYER M1 ;
        RECT 9.952 16.344 9.984 16.416 ;
  LAYER M2 ;
        RECT 9.932 16.364 10.004 16.396 ;
  LAYER M1 ;
        RECT 9.728 19.62 9.76 19.692 ;
  LAYER M2 ;
        RECT 9.708 19.64 9.78 19.672 ;
  LAYER M1 ;
        RECT 9.728 19.488 9.76 19.656 ;
  LAYER M1 ;
        RECT 9.728 19.452 9.76 19.524 ;
  LAYER M2 ;
        RECT 9.708 19.472 9.78 19.504 ;
  LAYER M2 ;
        RECT 9.744 19.472 9.968 19.504 ;
  LAYER M1 ;
        RECT 9.952 19.452 9.984 19.524 ;
  LAYER M2 ;
        RECT 9.932 19.472 10.004 19.504 ;
  LAYER M1 ;
        RECT 9.728 22.728 9.76 22.8 ;
  LAYER M2 ;
        RECT 9.708 22.748 9.78 22.78 ;
  LAYER M1 ;
        RECT 9.728 22.596 9.76 22.764 ;
  LAYER M1 ;
        RECT 9.728 22.56 9.76 22.632 ;
  LAYER M2 ;
        RECT 9.708 22.58 9.78 22.612 ;
  LAYER M2 ;
        RECT 9.744 22.58 9.968 22.612 ;
  LAYER M1 ;
        RECT 9.952 22.56 9.984 22.632 ;
  LAYER M2 ;
        RECT 9.932 22.58 10.004 22.612 ;
  LAYER M1 ;
        RECT 9.728 25.836 9.76 25.908 ;
  LAYER M2 ;
        RECT 9.708 25.856 9.78 25.888 ;
  LAYER M1 ;
        RECT 9.728 25.704 9.76 25.872 ;
  LAYER M1 ;
        RECT 9.728 25.668 9.76 25.74 ;
  LAYER M2 ;
        RECT 9.708 25.688 9.78 25.72 ;
  LAYER M2 ;
        RECT 9.744 25.688 9.968 25.72 ;
  LAYER M1 ;
        RECT 9.952 25.668 9.984 25.74 ;
  LAYER M2 ;
        RECT 9.932 25.688 10.004 25.72 ;
  LAYER M1 ;
        RECT 9.728 28.944 9.76 29.016 ;
  LAYER M2 ;
        RECT 9.708 28.964 9.78 28.996 ;
  LAYER M1 ;
        RECT 9.728 28.812 9.76 28.98 ;
  LAYER M1 ;
        RECT 9.728 28.776 9.76 28.848 ;
  LAYER M2 ;
        RECT 9.708 28.796 9.78 28.828 ;
  LAYER M2 ;
        RECT 9.744 28.796 9.968 28.828 ;
  LAYER M1 ;
        RECT 9.952 28.776 9.984 28.848 ;
  LAYER M2 ;
        RECT 9.932 28.796 10.004 28.828 ;
  LAYER M1 ;
        RECT 9.728 32.052 9.76 32.124 ;
  LAYER M2 ;
        RECT 9.708 32.072 9.78 32.104 ;
  LAYER M1 ;
        RECT 9.728 31.92 9.76 32.088 ;
  LAYER M1 ;
        RECT 9.728 31.884 9.76 31.956 ;
  LAYER M2 ;
        RECT 9.708 31.904 9.78 31.936 ;
  LAYER M2 ;
        RECT 9.744 31.904 9.968 31.936 ;
  LAYER M1 ;
        RECT 9.952 31.884 9.984 31.956 ;
  LAYER M2 ;
        RECT 9.932 31.904 10.004 31.936 ;
  LAYER M1 ;
        RECT 9.952 0.048 9.984 0.12 ;
  LAYER M2 ;
        RECT 9.932 0.068 10.004 0.1 ;
  LAYER M1 ;
        RECT 9.952 0.084 9.984 0.672 ;
  LAYER M1 ;
        RECT 9.952 0.672 9.984 31.92 ;
  LAYER M2 ;
        RECT 0.08 0.068 9.968 0.1 ;
  LAYER M1 ;
        RECT 6.432 0.972 6.464 1.044 ;
  LAYER M2 ;
        RECT 6.412 0.992 6.484 1.024 ;
  LAYER M2 ;
        RECT 3.152 0.992 6.448 1.024 ;
  LAYER M1 ;
        RECT 3.136 0.972 3.168 1.044 ;
  LAYER M2 ;
        RECT 3.116 0.992 3.188 1.024 ;
  LAYER M1 ;
        RECT 6.432 32.052 6.464 32.124 ;
  LAYER M2 ;
        RECT 6.412 32.072 6.484 32.104 ;
  LAYER M2 ;
        RECT 3.152 32.072 6.448 32.104 ;
  LAYER M1 ;
        RECT 3.136 32.052 3.168 32.124 ;
  LAYER M2 ;
        RECT 3.116 32.072 3.188 32.104 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M2 ;
        RECT 3.696 18.968 4.08 19 ;
  LAYER M1 ;
        RECT 3.68 18.948 3.712 19.02 ;
  LAYER M2 ;
        RECT 3.66 18.968 3.732 19 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M2 ;
        RECT 3.696 6.536 4.08 6.568 ;
  LAYER M1 ;
        RECT 3.68 6.516 3.712 6.588 ;
  LAYER M2 ;
        RECT 3.66 6.536 3.732 6.568 ;
  LAYER M1 ;
        RECT 4.064 31.38 4.096 31.452 ;
  LAYER M2 ;
        RECT 4.044 31.4 4.116 31.432 ;
  LAYER M2 ;
        RECT 3.696 31.4 4.08 31.432 ;
  LAYER M1 ;
        RECT 3.68 31.38 3.712 31.452 ;
  LAYER M2 ;
        RECT 3.66 31.4 3.732 31.432 ;
  LAYER M1 ;
        RECT 3.68 35.076 3.712 35.148 ;
  LAYER M2 ;
        RECT 3.66 35.096 3.732 35.128 ;
  LAYER M1 ;
        RECT 3.68 34.86 3.712 35.112 ;
  LAYER M1 ;
        RECT 3.68 6.552 3.712 34.86 ;
  LAYER M1 ;
        RECT 4.064 18.948 4.096 19.02 ;
  LAYER M2 ;
        RECT 4.044 18.968 4.116 19 ;
  LAYER M1 ;
        RECT 4.064 18.984 4.096 19.152 ;
  LAYER M1 ;
        RECT 4.064 19.116 4.096 19.188 ;
  LAYER M2 ;
        RECT 4.044 19.136 4.116 19.168 ;
  LAYER M2 ;
        RECT 4.08 19.136 6.992 19.168 ;
  LAYER M1 ;
        RECT 6.976 19.116 7.008 19.188 ;
  LAYER M2 ;
        RECT 6.956 19.136 7.028 19.168 ;
  LAYER M1 ;
        RECT 4.064 6.516 4.096 6.588 ;
  LAYER M2 ;
        RECT 4.044 6.536 4.116 6.568 ;
  LAYER M1 ;
        RECT 4.064 6.552 4.096 6.72 ;
  LAYER M1 ;
        RECT 4.064 6.684 4.096 6.756 ;
  LAYER M2 ;
        RECT 4.044 6.704 4.116 6.736 ;
  LAYER M2 ;
        RECT 4.08 6.704 6.992 6.736 ;
  LAYER M1 ;
        RECT 6.976 6.684 7.008 6.756 ;
  LAYER M2 ;
        RECT 6.956 6.704 7.028 6.736 ;
  LAYER M1 ;
        RECT 4.064 31.38 4.096 31.452 ;
  LAYER M2 ;
        RECT 4.044 31.4 4.116 31.432 ;
  LAYER M1 ;
        RECT 4.064 31.416 4.096 31.584 ;
  LAYER M1 ;
        RECT 4.064 31.548 4.096 31.62 ;
  LAYER M2 ;
        RECT 4.044 31.568 4.116 31.6 ;
  LAYER M2 ;
        RECT 4.08 31.568 6.992 31.6 ;
  LAYER M1 ;
        RECT 6.976 31.548 7.008 31.62 ;
  LAYER M2 ;
        RECT 6.956 31.568 7.028 31.6 ;
  LAYER M1 ;
        RECT 6.976 35.076 7.008 35.148 ;
  LAYER M2 ;
        RECT 6.956 35.096 7.028 35.128 ;
  LAYER M1 ;
        RECT 6.976 34.86 7.008 35.112 ;
  LAYER M1 ;
        RECT 6.976 6.72 7.008 34.86 ;
  LAYER M2 ;
        RECT 3.696 35.096 6.992 35.128 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M2 ;
        RECT 3.856 15.86 4.08 15.892 ;
  LAYER M1 ;
        RECT 3.84 15.84 3.872 15.912 ;
  LAYER M2 ;
        RECT 3.82 15.86 3.892 15.892 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M2 ;
        RECT 3.856 22.076 4.08 22.108 ;
  LAYER M1 ;
        RECT 3.84 22.056 3.872 22.128 ;
  LAYER M2 ;
        RECT 3.82 22.076 3.892 22.108 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M2 ;
        RECT 3.856 12.752 4.08 12.784 ;
  LAYER M1 ;
        RECT 3.84 12.732 3.872 12.804 ;
  LAYER M2 ;
        RECT 3.82 12.752 3.892 12.784 ;
  LAYER M1 ;
        RECT 4.064 25.164 4.096 25.236 ;
  LAYER M2 ;
        RECT 4.044 25.184 4.116 25.216 ;
  LAYER M2 ;
        RECT 3.856 25.184 4.08 25.216 ;
  LAYER M1 ;
        RECT 3.84 25.164 3.872 25.236 ;
  LAYER M2 ;
        RECT 3.82 25.184 3.892 25.216 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M2 ;
        RECT 3.856 9.644 4.08 9.676 ;
  LAYER M1 ;
        RECT 3.84 9.624 3.872 9.696 ;
  LAYER M2 ;
        RECT 3.82 9.644 3.892 9.676 ;
  LAYER M1 ;
        RECT 4.064 28.272 4.096 28.344 ;
  LAYER M2 ;
        RECT 4.044 28.292 4.116 28.324 ;
  LAYER M2 ;
        RECT 3.856 28.292 4.08 28.324 ;
  LAYER M1 ;
        RECT 3.84 28.272 3.872 28.344 ;
  LAYER M2 ;
        RECT 3.82 28.292 3.892 28.324 ;
  LAYER M1 ;
        RECT 3.84 35.244 3.872 35.316 ;
  LAYER M2 ;
        RECT 3.82 35.264 3.892 35.296 ;
  LAYER M1 ;
        RECT 3.84 34.86 3.872 35.28 ;
  LAYER M1 ;
        RECT 3.84 9.66 3.872 34.86 ;
  LAYER M1 ;
        RECT 4.064 15.84 4.096 15.912 ;
  LAYER M2 ;
        RECT 4.044 15.86 4.116 15.892 ;
  LAYER M1 ;
        RECT 4.064 15.876 4.096 16.044 ;
  LAYER M1 ;
        RECT 4.064 16.008 4.096 16.08 ;
  LAYER M2 ;
        RECT 4.044 16.028 4.116 16.06 ;
  LAYER M2 ;
        RECT 4.08 16.028 7.152 16.06 ;
  LAYER M1 ;
        RECT 7.136 16.008 7.168 16.08 ;
  LAYER M2 ;
        RECT 7.116 16.028 7.188 16.06 ;
  LAYER M1 ;
        RECT 4.064 22.056 4.096 22.128 ;
  LAYER M2 ;
        RECT 4.044 22.076 4.116 22.108 ;
  LAYER M1 ;
        RECT 4.064 22.092 4.096 22.26 ;
  LAYER M1 ;
        RECT 4.064 22.224 4.096 22.296 ;
  LAYER M2 ;
        RECT 4.044 22.244 4.116 22.276 ;
  LAYER M2 ;
        RECT 4.08 22.244 7.152 22.276 ;
  LAYER M1 ;
        RECT 7.136 22.224 7.168 22.296 ;
  LAYER M2 ;
        RECT 7.116 22.244 7.188 22.276 ;
  LAYER M1 ;
        RECT 4.064 12.732 4.096 12.804 ;
  LAYER M2 ;
        RECT 4.044 12.752 4.116 12.784 ;
  LAYER M1 ;
        RECT 4.064 12.768 4.096 12.936 ;
  LAYER M1 ;
        RECT 4.064 12.9 4.096 12.972 ;
  LAYER M2 ;
        RECT 4.044 12.92 4.116 12.952 ;
  LAYER M2 ;
        RECT 4.08 12.92 7.152 12.952 ;
  LAYER M1 ;
        RECT 7.136 12.9 7.168 12.972 ;
  LAYER M2 ;
        RECT 7.116 12.92 7.188 12.952 ;
  LAYER M1 ;
        RECT 4.064 25.164 4.096 25.236 ;
  LAYER M2 ;
        RECT 4.044 25.184 4.116 25.216 ;
  LAYER M1 ;
        RECT 4.064 25.2 4.096 25.368 ;
  LAYER M1 ;
        RECT 4.064 25.332 4.096 25.404 ;
  LAYER M2 ;
        RECT 4.044 25.352 4.116 25.384 ;
  LAYER M2 ;
        RECT 4.08 25.352 7.152 25.384 ;
  LAYER M1 ;
        RECT 7.136 25.332 7.168 25.404 ;
  LAYER M2 ;
        RECT 7.116 25.352 7.188 25.384 ;
  LAYER M1 ;
        RECT 4.064 9.624 4.096 9.696 ;
  LAYER M2 ;
        RECT 4.044 9.644 4.116 9.676 ;
  LAYER M1 ;
        RECT 4.064 9.66 4.096 9.828 ;
  LAYER M1 ;
        RECT 4.064 9.792 4.096 9.864 ;
  LAYER M2 ;
        RECT 4.044 9.812 4.116 9.844 ;
  LAYER M2 ;
        RECT 4.08 9.812 7.152 9.844 ;
  LAYER M1 ;
        RECT 7.136 9.792 7.168 9.864 ;
  LAYER M2 ;
        RECT 7.116 9.812 7.188 9.844 ;
  LAYER M1 ;
        RECT 4.064 28.272 4.096 28.344 ;
  LAYER M2 ;
        RECT 4.044 28.292 4.116 28.324 ;
  LAYER M1 ;
        RECT 4.064 28.308 4.096 28.476 ;
  LAYER M1 ;
        RECT 4.064 28.44 4.096 28.512 ;
  LAYER M2 ;
        RECT 4.044 28.46 4.116 28.492 ;
  LAYER M2 ;
        RECT 4.08 28.46 7.152 28.492 ;
  LAYER M1 ;
        RECT 7.136 28.44 7.168 28.512 ;
  LAYER M2 ;
        RECT 7.116 28.46 7.188 28.492 ;
  LAYER M1 ;
        RECT 7.136 35.244 7.168 35.316 ;
  LAYER M2 ;
        RECT 7.116 35.264 7.188 35.296 ;
  LAYER M1 ;
        RECT 7.136 34.86 7.168 35.28 ;
  LAYER M1 ;
        RECT 7.136 9.828 7.168 34.86 ;
  LAYER M2 ;
        RECT 3.856 35.264 7.152 35.296 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M2 ;
        RECT 0.24 3.428 0.784 3.46 ;
  LAYER M1 ;
        RECT 0.224 3.408 0.256 3.48 ;
  LAYER M2 ;
        RECT 0.204 3.428 0.276 3.46 ;
  LAYER M1 ;
        RECT 0.768 6.516 0.8 6.588 ;
  LAYER M2 ;
        RECT 0.748 6.536 0.82 6.568 ;
  LAYER M2 ;
        RECT 0.24 6.536 0.784 6.568 ;
  LAYER M1 ;
        RECT 0.224 6.516 0.256 6.588 ;
  LAYER M2 ;
        RECT 0.204 6.536 0.276 6.568 ;
  LAYER M1 ;
        RECT 0.768 9.624 0.8 9.696 ;
  LAYER M2 ;
        RECT 0.748 9.644 0.82 9.676 ;
  LAYER M2 ;
        RECT 0.24 9.644 0.784 9.676 ;
  LAYER M1 ;
        RECT 0.224 9.624 0.256 9.696 ;
  LAYER M2 ;
        RECT 0.204 9.644 0.276 9.676 ;
  LAYER M1 ;
        RECT 0.768 12.732 0.8 12.804 ;
  LAYER M2 ;
        RECT 0.748 12.752 0.82 12.784 ;
  LAYER M2 ;
        RECT 0.24 12.752 0.784 12.784 ;
  LAYER M1 ;
        RECT 0.224 12.732 0.256 12.804 ;
  LAYER M2 ;
        RECT 0.204 12.752 0.276 12.784 ;
  LAYER M1 ;
        RECT 0.768 15.84 0.8 15.912 ;
  LAYER M2 ;
        RECT 0.748 15.86 0.82 15.892 ;
  LAYER M2 ;
        RECT 0.24 15.86 0.784 15.892 ;
  LAYER M1 ;
        RECT 0.224 15.84 0.256 15.912 ;
  LAYER M2 ;
        RECT 0.204 15.86 0.276 15.892 ;
  LAYER M1 ;
        RECT 0.768 18.948 0.8 19.02 ;
  LAYER M2 ;
        RECT 0.748 18.968 0.82 19 ;
  LAYER M2 ;
        RECT 0.24 18.968 0.784 19 ;
  LAYER M1 ;
        RECT 0.224 18.948 0.256 19.02 ;
  LAYER M2 ;
        RECT 0.204 18.968 0.276 19 ;
  LAYER M1 ;
        RECT 0.768 22.056 0.8 22.128 ;
  LAYER M2 ;
        RECT 0.748 22.076 0.82 22.108 ;
  LAYER M2 ;
        RECT 0.24 22.076 0.784 22.108 ;
  LAYER M1 ;
        RECT 0.224 22.056 0.256 22.128 ;
  LAYER M2 ;
        RECT 0.204 22.076 0.276 22.108 ;
  LAYER M1 ;
        RECT 0.768 25.164 0.8 25.236 ;
  LAYER M2 ;
        RECT 0.748 25.184 0.82 25.216 ;
  LAYER M2 ;
        RECT 0.24 25.184 0.784 25.216 ;
  LAYER M1 ;
        RECT 0.224 25.164 0.256 25.236 ;
  LAYER M2 ;
        RECT 0.204 25.184 0.276 25.216 ;
  LAYER M1 ;
        RECT 0.768 28.272 0.8 28.344 ;
  LAYER M2 ;
        RECT 0.748 28.292 0.82 28.324 ;
  LAYER M2 ;
        RECT 0.24 28.292 0.784 28.324 ;
  LAYER M1 ;
        RECT 0.224 28.272 0.256 28.344 ;
  LAYER M2 ;
        RECT 0.204 28.292 0.276 28.324 ;
  LAYER M1 ;
        RECT 0.768 31.38 0.8 31.452 ;
  LAYER M2 ;
        RECT 0.748 31.4 0.82 31.432 ;
  LAYER M2 ;
        RECT 0.24 31.4 0.784 31.432 ;
  LAYER M1 ;
        RECT 0.224 31.38 0.256 31.452 ;
  LAYER M2 ;
        RECT 0.204 31.4 0.276 31.432 ;
  LAYER M1 ;
        RECT 0.768 34.488 0.8 34.56 ;
  LAYER M2 ;
        RECT 0.748 34.508 0.82 34.54 ;
  LAYER M2 ;
        RECT 0.24 34.508 0.784 34.54 ;
  LAYER M1 ;
        RECT 0.224 34.488 0.256 34.56 ;
  LAYER M2 ;
        RECT 0.204 34.508 0.276 34.54 ;
  LAYER M1 ;
        RECT 0.224 35.412 0.256 35.484 ;
  LAYER M2 ;
        RECT 0.204 35.432 0.276 35.464 ;
  LAYER M1 ;
        RECT 0.224 34.86 0.256 35.448 ;
  LAYER M1 ;
        RECT 0.224 3.444 0.256 34.86 ;
  LAYER M1 ;
        RECT 7.36 3.408 7.392 3.48 ;
  LAYER M2 ;
        RECT 7.34 3.428 7.412 3.46 ;
  LAYER M1 ;
        RECT 7.36 3.444 7.392 3.612 ;
  LAYER M1 ;
        RECT 7.36 3.576 7.392 3.648 ;
  LAYER M2 ;
        RECT 7.34 3.596 7.412 3.628 ;
  LAYER M2 ;
        RECT 7.376 3.596 10.128 3.628 ;
  LAYER M1 ;
        RECT 10.112 3.576 10.144 3.648 ;
  LAYER M2 ;
        RECT 10.092 3.596 10.164 3.628 ;
  LAYER M1 ;
        RECT 7.36 6.516 7.392 6.588 ;
  LAYER M2 ;
        RECT 7.34 6.536 7.412 6.568 ;
  LAYER M1 ;
        RECT 7.36 6.552 7.392 6.72 ;
  LAYER M1 ;
        RECT 7.36 6.684 7.392 6.756 ;
  LAYER M2 ;
        RECT 7.34 6.704 7.412 6.736 ;
  LAYER M2 ;
        RECT 7.376 6.704 10.128 6.736 ;
  LAYER M1 ;
        RECT 10.112 6.684 10.144 6.756 ;
  LAYER M2 ;
        RECT 10.092 6.704 10.164 6.736 ;
  LAYER M1 ;
        RECT 7.36 9.624 7.392 9.696 ;
  LAYER M2 ;
        RECT 7.34 9.644 7.412 9.676 ;
  LAYER M1 ;
        RECT 7.36 9.66 7.392 9.828 ;
  LAYER M1 ;
        RECT 7.36 9.792 7.392 9.864 ;
  LAYER M2 ;
        RECT 7.34 9.812 7.412 9.844 ;
  LAYER M2 ;
        RECT 7.376 9.812 10.128 9.844 ;
  LAYER M1 ;
        RECT 10.112 9.792 10.144 9.864 ;
  LAYER M2 ;
        RECT 10.092 9.812 10.164 9.844 ;
  LAYER M1 ;
        RECT 7.36 12.732 7.392 12.804 ;
  LAYER M2 ;
        RECT 7.34 12.752 7.412 12.784 ;
  LAYER M1 ;
        RECT 7.36 12.768 7.392 12.936 ;
  LAYER M1 ;
        RECT 7.36 12.9 7.392 12.972 ;
  LAYER M2 ;
        RECT 7.34 12.92 7.412 12.952 ;
  LAYER M2 ;
        RECT 7.376 12.92 10.128 12.952 ;
  LAYER M1 ;
        RECT 10.112 12.9 10.144 12.972 ;
  LAYER M2 ;
        RECT 10.092 12.92 10.164 12.952 ;
  LAYER M1 ;
        RECT 7.36 15.84 7.392 15.912 ;
  LAYER M2 ;
        RECT 7.34 15.86 7.412 15.892 ;
  LAYER M1 ;
        RECT 7.36 15.876 7.392 16.044 ;
  LAYER M1 ;
        RECT 7.36 16.008 7.392 16.08 ;
  LAYER M2 ;
        RECT 7.34 16.028 7.412 16.06 ;
  LAYER M2 ;
        RECT 7.376 16.028 10.128 16.06 ;
  LAYER M1 ;
        RECT 10.112 16.008 10.144 16.08 ;
  LAYER M2 ;
        RECT 10.092 16.028 10.164 16.06 ;
  LAYER M1 ;
        RECT 7.36 18.948 7.392 19.02 ;
  LAYER M2 ;
        RECT 7.34 18.968 7.412 19 ;
  LAYER M1 ;
        RECT 7.36 18.984 7.392 19.152 ;
  LAYER M1 ;
        RECT 7.36 19.116 7.392 19.188 ;
  LAYER M2 ;
        RECT 7.34 19.136 7.412 19.168 ;
  LAYER M2 ;
        RECT 7.376 19.136 10.128 19.168 ;
  LAYER M1 ;
        RECT 10.112 19.116 10.144 19.188 ;
  LAYER M2 ;
        RECT 10.092 19.136 10.164 19.168 ;
  LAYER M1 ;
        RECT 7.36 22.056 7.392 22.128 ;
  LAYER M2 ;
        RECT 7.34 22.076 7.412 22.108 ;
  LAYER M1 ;
        RECT 7.36 22.092 7.392 22.26 ;
  LAYER M1 ;
        RECT 7.36 22.224 7.392 22.296 ;
  LAYER M2 ;
        RECT 7.34 22.244 7.412 22.276 ;
  LAYER M2 ;
        RECT 7.376 22.244 10.128 22.276 ;
  LAYER M1 ;
        RECT 10.112 22.224 10.144 22.296 ;
  LAYER M2 ;
        RECT 10.092 22.244 10.164 22.276 ;
  LAYER M1 ;
        RECT 7.36 25.164 7.392 25.236 ;
  LAYER M2 ;
        RECT 7.34 25.184 7.412 25.216 ;
  LAYER M1 ;
        RECT 7.36 25.2 7.392 25.368 ;
  LAYER M1 ;
        RECT 7.36 25.332 7.392 25.404 ;
  LAYER M2 ;
        RECT 7.34 25.352 7.412 25.384 ;
  LAYER M2 ;
        RECT 7.376 25.352 10.128 25.384 ;
  LAYER M1 ;
        RECT 10.112 25.332 10.144 25.404 ;
  LAYER M2 ;
        RECT 10.092 25.352 10.164 25.384 ;
  LAYER M1 ;
        RECT 7.36 28.272 7.392 28.344 ;
  LAYER M2 ;
        RECT 7.34 28.292 7.412 28.324 ;
  LAYER M1 ;
        RECT 7.36 28.308 7.392 28.476 ;
  LAYER M1 ;
        RECT 7.36 28.44 7.392 28.512 ;
  LAYER M2 ;
        RECT 7.34 28.46 7.412 28.492 ;
  LAYER M2 ;
        RECT 7.376 28.46 10.128 28.492 ;
  LAYER M1 ;
        RECT 10.112 28.44 10.144 28.512 ;
  LAYER M2 ;
        RECT 10.092 28.46 10.164 28.492 ;
  LAYER M1 ;
        RECT 7.36 31.38 7.392 31.452 ;
  LAYER M2 ;
        RECT 7.34 31.4 7.412 31.432 ;
  LAYER M1 ;
        RECT 7.36 31.416 7.392 31.584 ;
  LAYER M1 ;
        RECT 7.36 31.548 7.392 31.62 ;
  LAYER M2 ;
        RECT 7.34 31.568 7.412 31.6 ;
  LAYER M2 ;
        RECT 7.376 31.568 10.128 31.6 ;
  LAYER M1 ;
        RECT 10.112 31.548 10.144 31.62 ;
  LAYER M2 ;
        RECT 10.092 31.568 10.164 31.6 ;
  LAYER M1 ;
        RECT 7.36 34.488 7.392 34.56 ;
  LAYER M2 ;
        RECT 7.34 34.508 7.412 34.54 ;
  LAYER M1 ;
        RECT 7.36 34.524 7.392 34.692 ;
  LAYER M1 ;
        RECT 7.36 34.656 7.392 34.728 ;
  LAYER M2 ;
        RECT 7.34 34.676 7.412 34.708 ;
  LAYER M2 ;
        RECT 7.376 34.676 10.128 34.708 ;
  LAYER M1 ;
        RECT 10.112 34.656 10.144 34.728 ;
  LAYER M2 ;
        RECT 10.092 34.676 10.164 34.708 ;
  LAYER M1 ;
        RECT 10.112 35.412 10.144 35.484 ;
  LAYER M2 ;
        RECT 10.092 35.432 10.164 35.464 ;
  LAYER M1 ;
        RECT 10.112 34.86 10.144 35.448 ;
  LAYER M1 ;
        RECT 10.112 3.612 10.144 34.86 ;
  LAYER M2 ;
        RECT 0.24 35.432 10.128 35.464 ;
  LAYER M1 ;
        RECT 4.064 3.408 4.096 3.48 ;
  LAYER M2 ;
        RECT 4.044 3.428 4.116 3.46 ;
  LAYER M2 ;
        RECT 0.784 3.428 4.08 3.46 ;
  LAYER M1 ;
        RECT 0.768 3.408 0.8 3.48 ;
  LAYER M2 ;
        RECT 0.748 3.428 0.82 3.46 ;
  LAYER M1 ;
        RECT 4.064 34.488 4.096 34.56 ;
  LAYER M2 ;
        RECT 4.044 34.508 4.116 34.54 ;
  LAYER M2 ;
        RECT 0.784 34.508 4.08 34.54 ;
  LAYER M1 ;
        RECT 0.768 34.488 0.8 34.56 ;
  LAYER M2 ;
        RECT 0.748 34.508 0.82 34.54 ;
  LAYER M1 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M3 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M2 ;
        RECT 0.72 0.924 3.216 3.528 ;
  LAYER M1 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M3 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M2 ;
        RECT 0.72 4.032 3.216 6.636 ;
  LAYER M1 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M3 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M2 ;
        RECT 0.72 7.14 3.216 9.744 ;
  LAYER M1 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M3 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M2 ;
        RECT 0.72 10.248 3.216 12.852 ;
  LAYER M1 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M3 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M2 ;
        RECT 0.72 13.356 3.216 15.96 ;
  LAYER M1 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M3 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M2 ;
        RECT 0.72 16.464 3.216 19.068 ;
  LAYER M1 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M3 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M2 ;
        RECT 0.72 19.572 3.216 22.176 ;
  LAYER M1 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M3 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M2 ;
        RECT 0.72 22.68 3.216 25.284 ;
  LAYER M1 ;
        RECT 0.72 25.788 3.216 28.392 ;
  LAYER M3 ;
        RECT 0.72 25.788 3.216 28.392 ;
  LAYER M2 ;
        RECT 0.72 25.788 3.216 28.392 ;
  LAYER M1 ;
        RECT 0.72 28.896 3.216 31.5 ;
  LAYER M3 ;
        RECT 0.72 28.896 3.216 31.5 ;
  LAYER M2 ;
        RECT 0.72 28.896 3.216 31.5 ;
  LAYER M1 ;
        RECT 0.72 32.004 3.216 34.608 ;
  LAYER M3 ;
        RECT 0.72 32.004 3.216 34.608 ;
  LAYER M2 ;
        RECT 0.72 32.004 3.216 34.608 ;
  LAYER M1 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M3 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M2 ;
        RECT 4.016 0.924 6.512 3.528 ;
  LAYER M1 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M3 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M2 ;
        RECT 4.016 4.032 6.512 6.636 ;
  LAYER M1 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M3 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M2 ;
        RECT 4.016 7.14 6.512 9.744 ;
  LAYER M1 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M3 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M2 ;
        RECT 4.016 10.248 6.512 12.852 ;
  LAYER M1 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M3 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M2 ;
        RECT 4.016 13.356 6.512 15.96 ;
  LAYER M1 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M3 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M2 ;
        RECT 4.016 16.464 6.512 19.068 ;
  LAYER M1 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M3 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M2 ;
        RECT 4.016 19.572 6.512 22.176 ;
  LAYER M1 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M3 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M2 ;
        RECT 4.016 22.68 6.512 25.284 ;
  LAYER M1 ;
        RECT 4.016 25.788 6.512 28.392 ;
  LAYER M3 ;
        RECT 4.016 25.788 6.512 28.392 ;
  LAYER M2 ;
        RECT 4.016 25.788 6.512 28.392 ;
  LAYER M1 ;
        RECT 4.016 28.896 6.512 31.5 ;
  LAYER M3 ;
        RECT 4.016 28.896 6.512 31.5 ;
  LAYER M2 ;
        RECT 4.016 28.896 6.512 31.5 ;
  LAYER M1 ;
        RECT 4.016 32.004 6.512 34.608 ;
  LAYER M3 ;
        RECT 4.016 32.004 6.512 34.608 ;
  LAYER M2 ;
        RECT 4.016 32.004 6.512 34.608 ;
  LAYER M1 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M3 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M2 ;
        RECT 7.312 0.924 9.808 3.528 ;
  LAYER M1 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M3 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M2 ;
        RECT 7.312 4.032 9.808 6.636 ;
  LAYER M1 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M3 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M2 ;
        RECT 7.312 7.14 9.808 9.744 ;
  LAYER M1 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M3 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M2 ;
        RECT 7.312 10.248 9.808 12.852 ;
  LAYER M1 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M3 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M2 ;
        RECT 7.312 13.356 9.808 15.96 ;
  LAYER M1 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M3 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M2 ;
        RECT 7.312 16.464 9.808 19.068 ;
  LAYER M1 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M3 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M2 ;
        RECT 7.312 19.572 9.808 22.176 ;
  LAYER M1 ;
        RECT 7.312 22.68 9.808 25.284 ;
  LAYER M3 ;
        RECT 7.312 22.68 9.808 25.284 ;
  LAYER M2 ;
        RECT 7.312 22.68 9.808 25.284 ;
  LAYER M1 ;
        RECT 7.312 25.788 9.808 28.392 ;
  LAYER M3 ;
        RECT 7.312 25.788 9.808 28.392 ;
  LAYER M2 ;
        RECT 7.312 25.788 9.808 28.392 ;
  LAYER M1 ;
        RECT 7.312 28.896 9.808 31.5 ;
  LAYER M3 ;
        RECT 7.312 28.896 9.808 31.5 ;
  LAYER M2 ;
        RECT 7.312 28.896 9.808 31.5 ;
  LAYER M1 ;
        RECT 7.312 32.004 9.808 34.608 ;
  LAYER M3 ;
        RECT 7.312 32.004 9.808 34.608 ;
  LAYER M2 ;
        RECT 7.312 32.004 9.808 34.608 ;
  END 
END Cap_30fF_Cap_60fF
