MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 12 BY 19.656 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 3.2 19.368 3.232 19.44 ;
      LAYER M2 ;
        RECT 3.18 19.388 3.252 19.42 ;
      LAYER M1 ;
        RECT 9.152 19.368 9.184 19.44 ;
      LAYER M2 ;
        RECT 9.132 19.388 9.204 19.42 ;
      LAYER M2 ;
        RECT 3.216 19.388 9.168 19.42 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
      LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 5.728 7.02 5.76 7.092 ;
  LAYER M2 ;
        RECT 5.708 7.04 5.78 7.072 ;
  LAYER M1 ;
        RECT 5.728 6.888 5.76 7.056 ;
  LAYER M1 ;
        RECT 5.728 6.852 5.76 6.924 ;
  LAYER M2 ;
        RECT 5.708 6.872 5.78 6.904 ;
  LAYER M2 ;
        RECT 5.744 6.872 5.904 6.904 ;
  LAYER M1 ;
        RECT 5.888 6.852 5.92 6.924 ;
  LAYER M2 ;
        RECT 5.868 6.872 5.94 6.904 ;
  LAYER M1 ;
        RECT 8.704 10.128 8.736 10.2 ;
  LAYER M2 ;
        RECT 8.684 10.148 8.756 10.18 ;
  LAYER M2 ;
        RECT 5.904 10.148 8.72 10.18 ;
  LAYER M1 ;
        RECT 5.888 10.128 5.92 10.2 ;
  LAYER M2 ;
        RECT 5.868 10.148 5.94 10.18 ;
  LAYER M1 ;
        RECT 5.728 10.128 5.76 10.2 ;
  LAYER M2 ;
        RECT 5.708 10.148 5.78 10.18 ;
  LAYER M1 ;
        RECT 5.728 9.996 5.76 10.164 ;
  LAYER M1 ;
        RECT 5.728 9.96 5.76 10.032 ;
  LAYER M2 ;
        RECT 5.708 9.98 5.78 10.012 ;
  LAYER M2 ;
        RECT 5.744 9.98 5.904 10.012 ;
  LAYER M1 ;
        RECT 5.888 9.96 5.92 10.032 ;
  LAYER M2 ;
        RECT 5.868 9.98 5.94 10.012 ;
  LAYER M1 ;
        RECT 8.704 7.02 8.736 7.092 ;
  LAYER M2 ;
        RECT 8.684 7.04 8.756 7.072 ;
  LAYER M2 ;
        RECT 5.904 7.04 8.72 7.072 ;
  LAYER M1 ;
        RECT 5.888 7.02 5.92 7.092 ;
  LAYER M2 ;
        RECT 5.868 7.04 5.94 7.072 ;
  LAYER M1 ;
        RECT 5.728 13.236 5.76 13.308 ;
  LAYER M2 ;
        RECT 5.708 13.256 5.78 13.288 ;
  LAYER M1 ;
        RECT 5.728 13.104 5.76 13.272 ;
  LAYER M1 ;
        RECT 5.728 13.068 5.76 13.14 ;
  LAYER M2 ;
        RECT 5.708 13.088 5.78 13.12 ;
  LAYER M2 ;
        RECT 5.744 13.088 5.904 13.12 ;
  LAYER M1 ;
        RECT 5.888 13.068 5.92 13.14 ;
  LAYER M2 ;
        RECT 5.868 13.088 5.94 13.12 ;
  LAYER M1 ;
        RECT 8.704 3.912 8.736 3.984 ;
  LAYER M2 ;
        RECT 8.684 3.932 8.756 3.964 ;
  LAYER M2 ;
        RECT 5.904 3.932 8.72 3.964 ;
  LAYER M1 ;
        RECT 5.888 3.912 5.92 3.984 ;
  LAYER M2 ;
        RECT 5.868 3.932 5.94 3.964 ;
  LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
  LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
  LAYER M1 ;
        RECT 5.888 0.252 5.92 0.504 ;
  LAYER M1 ;
        RECT 5.888 0.504 5.92 13.104 ;
  LAYER M1 ;
        RECT 2.752 0.804 2.784 0.876 ;
  LAYER M2 ;
        RECT 2.732 0.824 2.804 0.856 ;
  LAYER M1 ;
        RECT 2.752 0.672 2.784 0.84 ;
  LAYER M1 ;
        RECT 2.752 0.636 2.784 0.708 ;
  LAYER M2 ;
        RECT 2.732 0.656 2.804 0.688 ;
  LAYER M2 ;
        RECT 2.768 0.656 2.928 0.688 ;
  LAYER M1 ;
        RECT 2.912 0.636 2.944 0.708 ;
  LAYER M2 ;
        RECT 2.892 0.656 2.964 0.688 ;
  LAYER M1 ;
        RECT 2.752 3.912 2.784 3.984 ;
  LAYER M2 ;
        RECT 2.732 3.932 2.804 3.964 ;
  LAYER M1 ;
        RECT 2.752 3.78 2.784 3.948 ;
  LAYER M1 ;
        RECT 2.752 3.744 2.784 3.816 ;
  LAYER M2 ;
        RECT 2.732 3.764 2.804 3.796 ;
  LAYER M2 ;
        RECT 2.768 3.764 2.928 3.796 ;
  LAYER M1 ;
        RECT 2.912 3.744 2.944 3.816 ;
  LAYER M2 ;
        RECT 2.892 3.764 2.964 3.796 ;
  LAYER M1 ;
        RECT 2.752 7.02 2.784 7.092 ;
  LAYER M2 ;
        RECT 2.732 7.04 2.804 7.072 ;
  LAYER M1 ;
        RECT 2.752 6.888 2.784 7.056 ;
  LAYER M1 ;
        RECT 2.752 6.852 2.784 6.924 ;
  LAYER M2 ;
        RECT 2.732 6.872 2.804 6.904 ;
  LAYER M2 ;
        RECT 2.768 6.872 2.928 6.904 ;
  LAYER M1 ;
        RECT 2.912 6.852 2.944 6.924 ;
  LAYER M2 ;
        RECT 2.892 6.872 2.964 6.904 ;
  LAYER M1 ;
        RECT 2.752 10.128 2.784 10.2 ;
  LAYER M2 ;
        RECT 2.732 10.148 2.804 10.18 ;
  LAYER M1 ;
        RECT 2.752 9.996 2.784 10.164 ;
  LAYER M1 ;
        RECT 2.752 9.96 2.784 10.032 ;
  LAYER M2 ;
        RECT 2.732 9.98 2.804 10.012 ;
  LAYER M2 ;
        RECT 2.768 9.98 2.928 10.012 ;
  LAYER M1 ;
        RECT 2.912 9.96 2.944 10.032 ;
  LAYER M2 ;
        RECT 2.892 9.98 2.964 10.012 ;
  LAYER M1 ;
        RECT 2.752 13.236 2.784 13.308 ;
  LAYER M2 ;
        RECT 2.732 13.256 2.804 13.288 ;
  LAYER M1 ;
        RECT 2.752 13.104 2.784 13.272 ;
  LAYER M1 ;
        RECT 2.752 13.068 2.784 13.14 ;
  LAYER M2 ;
        RECT 2.732 13.088 2.804 13.12 ;
  LAYER M2 ;
        RECT 2.768 13.088 2.928 13.12 ;
  LAYER M1 ;
        RECT 2.912 13.068 2.944 13.14 ;
  LAYER M2 ;
        RECT 2.892 13.088 2.964 13.12 ;
  LAYER M1 ;
        RECT 2.752 16.344 2.784 16.416 ;
  LAYER M2 ;
        RECT 2.732 16.364 2.804 16.396 ;
  LAYER M1 ;
        RECT 2.752 16.212 2.784 16.38 ;
  LAYER M1 ;
        RECT 2.752 16.176 2.784 16.248 ;
  LAYER M2 ;
        RECT 2.732 16.196 2.804 16.228 ;
  LAYER M2 ;
        RECT 2.768 16.196 2.928 16.228 ;
  LAYER M1 ;
        RECT 2.912 16.176 2.944 16.248 ;
  LAYER M2 ;
        RECT 2.892 16.196 2.964 16.228 ;
  LAYER M1 ;
        RECT 5.728 0.804 5.76 0.876 ;
  LAYER M2 ;
        RECT 5.708 0.824 5.78 0.856 ;
  LAYER M2 ;
        RECT 2.928 0.824 5.744 0.856 ;
  LAYER M1 ;
        RECT 2.912 0.804 2.944 0.876 ;
  LAYER M2 ;
        RECT 2.892 0.824 2.964 0.856 ;
  LAYER M1 ;
        RECT 5.728 3.912 5.76 3.984 ;
  LAYER M2 ;
        RECT 5.708 3.932 5.78 3.964 ;
  LAYER M2 ;
        RECT 2.928 3.932 5.744 3.964 ;
  LAYER M1 ;
        RECT 2.912 3.912 2.944 3.984 ;
  LAYER M2 ;
        RECT 2.892 3.932 2.964 3.964 ;
  LAYER M1 ;
        RECT 5.728 16.344 5.76 16.416 ;
  LAYER M2 ;
        RECT 5.708 16.364 5.78 16.396 ;
  LAYER M2 ;
        RECT 2.928 16.364 5.744 16.396 ;
  LAYER M1 ;
        RECT 2.912 16.344 2.944 16.416 ;
  LAYER M2 ;
        RECT 2.892 16.364 2.964 16.396 ;
  LAYER M1 ;
        RECT 2.912 0.048 2.944 0.12 ;
  LAYER M2 ;
        RECT 2.892 0.068 2.964 0.1 ;
  LAYER M1 ;
        RECT 2.912 0.084 2.944 0.504 ;
  LAYER M1 ;
        RECT 2.912 0.504 2.944 16.38 ;
  LAYER M1 ;
        RECT 8.704 0.804 8.736 0.876 ;
  LAYER M2 ;
        RECT 8.684 0.824 8.756 0.856 ;
  LAYER M1 ;
        RECT 8.704 0.672 8.736 0.84 ;
  LAYER M1 ;
        RECT 8.704 0.636 8.736 0.708 ;
  LAYER M2 ;
        RECT 8.684 0.656 8.756 0.688 ;
  LAYER M2 ;
        RECT 8.72 0.656 8.88 0.688 ;
  LAYER M1 ;
        RECT 8.864 0.636 8.896 0.708 ;
  LAYER M2 ;
        RECT 8.844 0.656 8.916 0.688 ;
  LAYER M1 ;
        RECT 8.704 13.236 8.736 13.308 ;
  LAYER M2 ;
        RECT 8.684 13.256 8.756 13.288 ;
  LAYER M1 ;
        RECT 8.704 13.104 8.736 13.272 ;
  LAYER M1 ;
        RECT 8.704 13.068 8.736 13.14 ;
  LAYER M2 ;
        RECT 8.684 13.088 8.756 13.12 ;
  LAYER M2 ;
        RECT 8.72 13.088 8.88 13.12 ;
  LAYER M1 ;
        RECT 8.864 13.068 8.896 13.14 ;
  LAYER M2 ;
        RECT 8.844 13.088 8.916 13.12 ;
  LAYER M1 ;
        RECT 8.704 16.344 8.736 16.416 ;
  LAYER M2 ;
        RECT 8.684 16.364 8.756 16.396 ;
  LAYER M1 ;
        RECT 8.704 16.212 8.736 16.38 ;
  LAYER M1 ;
        RECT 8.704 16.176 8.736 16.248 ;
  LAYER M2 ;
        RECT 8.684 16.196 8.756 16.228 ;
  LAYER M2 ;
        RECT 8.72 16.196 8.88 16.228 ;
  LAYER M1 ;
        RECT 8.864 16.176 8.896 16.248 ;
  LAYER M2 ;
        RECT 8.844 16.196 8.916 16.228 ;
  LAYER M1 ;
        RECT 11.68 0.804 11.712 0.876 ;
  LAYER M2 ;
        RECT 11.66 0.824 11.732 0.856 ;
  LAYER M2 ;
        RECT 8.88 0.824 11.696 0.856 ;
  LAYER M1 ;
        RECT 8.864 0.804 8.896 0.876 ;
  LAYER M2 ;
        RECT 8.844 0.824 8.916 0.856 ;
  LAYER M1 ;
        RECT 11.68 3.912 11.712 3.984 ;
  LAYER M2 ;
        RECT 11.66 3.932 11.732 3.964 ;
  LAYER M2 ;
        RECT 8.88 3.932 11.696 3.964 ;
  LAYER M1 ;
        RECT 8.864 3.912 8.896 3.984 ;
  LAYER M2 ;
        RECT 8.844 3.932 8.916 3.964 ;
  LAYER M1 ;
        RECT 11.68 7.02 11.712 7.092 ;
  LAYER M2 ;
        RECT 11.66 7.04 11.732 7.072 ;
  LAYER M2 ;
        RECT 8.88 7.04 11.696 7.072 ;
  LAYER M1 ;
        RECT 8.864 7.02 8.896 7.092 ;
  LAYER M2 ;
        RECT 8.844 7.04 8.916 7.072 ;
  LAYER M1 ;
        RECT 11.68 10.128 11.712 10.2 ;
  LAYER M2 ;
        RECT 11.66 10.148 11.732 10.18 ;
  LAYER M2 ;
        RECT 8.88 10.148 11.696 10.18 ;
  LAYER M1 ;
        RECT 8.864 10.128 8.896 10.2 ;
  LAYER M2 ;
        RECT 8.844 10.148 8.916 10.18 ;
  LAYER M1 ;
        RECT 11.68 13.236 11.712 13.308 ;
  LAYER M2 ;
        RECT 11.66 13.256 11.732 13.288 ;
  LAYER M2 ;
        RECT 8.88 13.256 11.696 13.288 ;
  LAYER M1 ;
        RECT 8.864 13.236 8.896 13.308 ;
  LAYER M2 ;
        RECT 8.844 13.256 8.916 13.288 ;
  LAYER M1 ;
        RECT 11.68 16.344 11.712 16.416 ;
  LAYER M2 ;
        RECT 11.66 16.364 11.732 16.396 ;
  LAYER M2 ;
        RECT 8.88 16.364 11.696 16.396 ;
  LAYER M1 ;
        RECT 8.864 16.344 8.896 16.416 ;
  LAYER M2 ;
        RECT 8.844 16.364 8.916 16.396 ;
  LAYER M1 ;
        RECT 8.864 0.048 8.896 0.12 ;
  LAYER M2 ;
        RECT 8.844 0.068 8.916 0.1 ;
  LAYER M1 ;
        RECT 8.864 0.084 8.896 0.504 ;
  LAYER M1 ;
        RECT 8.864 0.504 8.896 16.38 ;
  LAYER M2 ;
        RECT 2.928 0.068 8.88 0.1 ;
  LAYER M1 ;
        RECT 3.36 9.456 3.392 9.528 ;
  LAYER M2 ;
        RECT 3.34 9.476 3.412 9.508 ;
  LAYER M2 ;
        RECT 3.216 9.476 3.376 9.508 ;
  LAYER M1 ;
        RECT 3.2 9.456 3.232 9.528 ;
  LAYER M2 ;
        RECT 3.18 9.476 3.252 9.508 ;
  LAYER M1 ;
        RECT 3.36 12.564 3.392 12.636 ;
  LAYER M2 ;
        RECT 3.34 12.584 3.412 12.616 ;
  LAYER M2 ;
        RECT 3.216 12.584 3.376 12.616 ;
  LAYER M1 ;
        RECT 3.2 12.564 3.232 12.636 ;
  LAYER M2 ;
        RECT 3.18 12.584 3.252 12.616 ;
  LAYER M1 ;
        RECT 3.36 15.672 3.392 15.744 ;
  LAYER M2 ;
        RECT 3.34 15.692 3.412 15.724 ;
  LAYER M2 ;
        RECT 3.216 15.692 3.376 15.724 ;
  LAYER M1 ;
        RECT 3.2 15.672 3.232 15.744 ;
  LAYER M2 ;
        RECT 3.18 15.692 3.252 15.724 ;
  LAYER M1 ;
        RECT 3.2 19.368 3.232 19.44 ;
  LAYER M2 ;
        RECT 3.18 19.388 3.252 19.42 ;
  LAYER M1 ;
        RECT 3.2 19.152 3.232 19.404 ;
  LAYER M1 ;
        RECT 3.2 9.492 3.232 19.152 ;
  LAYER M1 ;
        RECT 6.336 12.564 6.368 12.636 ;
  LAYER M2 ;
        RECT 6.316 12.584 6.388 12.616 ;
  LAYER M1 ;
        RECT 6.336 12.6 6.368 12.768 ;
  LAYER M1 ;
        RECT 6.336 12.732 6.368 12.804 ;
  LAYER M2 ;
        RECT 6.316 12.752 6.388 12.784 ;
  LAYER M2 ;
        RECT 6.352 12.752 9.168 12.784 ;
  LAYER M1 ;
        RECT 9.152 12.732 9.184 12.804 ;
  LAYER M2 ;
        RECT 9.132 12.752 9.204 12.784 ;
  LAYER M1 ;
        RECT 6.336 9.456 6.368 9.528 ;
  LAYER M2 ;
        RECT 6.316 9.476 6.388 9.508 ;
  LAYER M1 ;
        RECT 6.336 9.492 6.368 9.66 ;
  LAYER M1 ;
        RECT 6.336 9.624 6.368 9.696 ;
  LAYER M2 ;
        RECT 6.316 9.644 6.388 9.676 ;
  LAYER M2 ;
        RECT 6.352 9.644 9.168 9.676 ;
  LAYER M1 ;
        RECT 9.152 9.624 9.184 9.696 ;
  LAYER M2 ;
        RECT 9.132 9.644 9.204 9.676 ;
  LAYER M1 ;
        RECT 6.336 6.348 6.368 6.42 ;
  LAYER M2 ;
        RECT 6.316 6.368 6.388 6.4 ;
  LAYER M1 ;
        RECT 6.336 6.384 6.368 6.552 ;
  LAYER M1 ;
        RECT 6.336 6.516 6.368 6.588 ;
  LAYER M2 ;
        RECT 6.316 6.536 6.388 6.568 ;
  LAYER M2 ;
        RECT 6.352 6.536 9.168 6.568 ;
  LAYER M1 ;
        RECT 9.152 6.516 9.184 6.588 ;
  LAYER M2 ;
        RECT 9.132 6.536 9.204 6.568 ;
  LAYER M1 ;
        RECT 9.152 19.368 9.184 19.44 ;
  LAYER M2 ;
        RECT 9.132 19.388 9.204 19.42 ;
  LAYER M1 ;
        RECT 9.152 19.152 9.184 19.404 ;
  LAYER M1 ;
        RECT 9.152 6.552 9.184 19.152 ;
  LAYER M2 ;
        RECT 3.216 19.388 9.168 19.42 ;
  LAYER M1 ;
        RECT 0.384 3.24 0.416 3.312 ;
  LAYER M2 ;
        RECT 0.364 3.26 0.436 3.292 ;
  LAYER M2 ;
        RECT 0.08 3.26 0.4 3.292 ;
  LAYER M1 ;
        RECT 0.064 3.24 0.096 3.312 ;
  LAYER M2 ;
        RECT 0.044 3.26 0.116 3.292 ;
  LAYER M1 ;
        RECT 0.384 6.348 0.416 6.42 ;
  LAYER M2 ;
        RECT 0.364 6.368 0.436 6.4 ;
  LAYER M2 ;
        RECT 0.08 6.368 0.4 6.4 ;
  LAYER M1 ;
        RECT 0.064 6.348 0.096 6.42 ;
  LAYER M2 ;
        RECT 0.044 6.368 0.116 6.4 ;
  LAYER M1 ;
        RECT 0.384 9.456 0.416 9.528 ;
  LAYER M2 ;
        RECT 0.364 9.476 0.436 9.508 ;
  LAYER M2 ;
        RECT 0.08 9.476 0.4 9.508 ;
  LAYER M1 ;
        RECT 0.064 9.456 0.096 9.528 ;
  LAYER M2 ;
        RECT 0.044 9.476 0.116 9.508 ;
  LAYER M1 ;
        RECT 0.384 12.564 0.416 12.636 ;
  LAYER M2 ;
        RECT 0.364 12.584 0.436 12.616 ;
  LAYER M2 ;
        RECT 0.08 12.584 0.4 12.616 ;
  LAYER M1 ;
        RECT 0.064 12.564 0.096 12.636 ;
  LAYER M2 ;
        RECT 0.044 12.584 0.116 12.616 ;
  LAYER M1 ;
        RECT 0.384 15.672 0.416 15.744 ;
  LAYER M2 ;
        RECT 0.364 15.692 0.436 15.724 ;
  LAYER M2 ;
        RECT 0.08 15.692 0.4 15.724 ;
  LAYER M1 ;
        RECT 0.064 15.672 0.096 15.744 ;
  LAYER M2 ;
        RECT 0.044 15.692 0.116 15.724 ;
  LAYER M1 ;
        RECT 0.384 18.78 0.416 18.852 ;
  LAYER M2 ;
        RECT 0.364 18.8 0.436 18.832 ;
  LAYER M2 ;
        RECT 0.08 18.8 0.4 18.832 ;
  LAYER M1 ;
        RECT 0.064 18.78 0.096 18.852 ;
  LAYER M2 ;
        RECT 0.044 18.8 0.116 18.832 ;
  LAYER M1 ;
        RECT 0.064 19.536 0.096 19.608 ;
  LAYER M2 ;
        RECT 0.044 19.556 0.116 19.588 ;
  LAYER M1 ;
        RECT 0.064 19.152 0.096 19.572 ;
  LAYER M1 ;
        RECT 0.064 3.276 0.096 19.152 ;
  LAYER M1 ;
        RECT 9.312 3.24 9.344 3.312 ;
  LAYER M2 ;
        RECT 9.292 3.26 9.364 3.292 ;
  LAYER M1 ;
        RECT 9.312 3.276 9.344 3.444 ;
  LAYER M1 ;
        RECT 9.312 3.408 9.344 3.48 ;
  LAYER M2 ;
        RECT 9.292 3.428 9.364 3.46 ;
  LAYER M2 ;
        RECT 9.328 3.428 11.984 3.46 ;
  LAYER M1 ;
        RECT 11.968 3.408 12 3.48 ;
  LAYER M2 ;
        RECT 11.948 3.428 12.02 3.46 ;
  LAYER M1 ;
        RECT 9.312 6.348 9.344 6.42 ;
  LAYER M2 ;
        RECT 9.292 6.368 9.364 6.4 ;
  LAYER M1 ;
        RECT 9.312 6.384 9.344 6.552 ;
  LAYER M1 ;
        RECT 9.312 6.516 9.344 6.588 ;
  LAYER M2 ;
        RECT 9.292 6.536 9.364 6.568 ;
  LAYER M2 ;
        RECT 9.328 6.536 11.984 6.568 ;
  LAYER M1 ;
        RECT 11.968 6.516 12 6.588 ;
  LAYER M2 ;
        RECT 11.948 6.536 12.02 6.568 ;
  LAYER M1 ;
        RECT 9.312 9.456 9.344 9.528 ;
  LAYER M2 ;
        RECT 9.292 9.476 9.364 9.508 ;
  LAYER M1 ;
        RECT 9.312 9.492 9.344 9.66 ;
  LAYER M1 ;
        RECT 9.312 9.624 9.344 9.696 ;
  LAYER M2 ;
        RECT 9.292 9.644 9.364 9.676 ;
  LAYER M2 ;
        RECT 9.328 9.644 11.984 9.676 ;
  LAYER M1 ;
        RECT 11.968 9.624 12 9.696 ;
  LAYER M2 ;
        RECT 11.948 9.644 12.02 9.676 ;
  LAYER M1 ;
        RECT 9.312 12.564 9.344 12.636 ;
  LAYER M2 ;
        RECT 9.292 12.584 9.364 12.616 ;
  LAYER M1 ;
        RECT 9.312 12.6 9.344 12.768 ;
  LAYER M1 ;
        RECT 9.312 12.732 9.344 12.804 ;
  LAYER M2 ;
        RECT 9.292 12.752 9.364 12.784 ;
  LAYER M2 ;
        RECT 9.328 12.752 11.984 12.784 ;
  LAYER M1 ;
        RECT 11.968 12.732 12 12.804 ;
  LAYER M2 ;
        RECT 11.948 12.752 12.02 12.784 ;
  LAYER M1 ;
        RECT 9.312 15.672 9.344 15.744 ;
  LAYER M2 ;
        RECT 9.292 15.692 9.364 15.724 ;
  LAYER M1 ;
        RECT 9.312 15.708 9.344 15.876 ;
  LAYER M1 ;
        RECT 9.312 15.84 9.344 15.912 ;
  LAYER M2 ;
        RECT 9.292 15.86 9.364 15.892 ;
  LAYER M2 ;
        RECT 9.328 15.86 11.984 15.892 ;
  LAYER M1 ;
        RECT 11.968 15.84 12 15.912 ;
  LAYER M2 ;
        RECT 11.948 15.86 12.02 15.892 ;
  LAYER M1 ;
        RECT 9.312 18.78 9.344 18.852 ;
  LAYER M2 ;
        RECT 9.292 18.8 9.364 18.832 ;
  LAYER M1 ;
        RECT 9.312 18.816 9.344 18.984 ;
  LAYER M1 ;
        RECT 9.312 18.948 9.344 19.02 ;
  LAYER M2 ;
        RECT 9.292 18.968 9.364 19 ;
  LAYER M2 ;
        RECT 9.328 18.968 11.984 19 ;
  LAYER M1 ;
        RECT 11.968 18.948 12 19.02 ;
  LAYER M2 ;
        RECT 11.948 18.968 12.02 19 ;
  LAYER M1 ;
        RECT 11.968 19.536 12 19.608 ;
  LAYER M2 ;
        RECT 11.948 19.556 12.02 19.588 ;
  LAYER M1 ;
        RECT 11.968 19.152 12 19.572 ;
  LAYER M1 ;
        RECT 11.968 3.444 12 19.152 ;
  LAYER M2 ;
        RECT 0.08 19.556 11.984 19.588 ;
  LAYER M1 ;
        RECT 3.36 3.24 3.392 3.312 ;
  LAYER M2 ;
        RECT 3.34 3.26 3.412 3.292 ;
  LAYER M2 ;
        RECT 0.4 3.26 3.376 3.292 ;
  LAYER M1 ;
        RECT 0.384 3.24 0.416 3.312 ;
  LAYER M2 ;
        RECT 0.364 3.26 0.436 3.292 ;
  LAYER M1 ;
        RECT 3.36 6.348 3.392 6.42 ;
  LAYER M2 ;
        RECT 3.34 6.368 3.412 6.4 ;
  LAYER M2 ;
        RECT 0.4 6.368 3.376 6.4 ;
  LAYER M1 ;
        RECT 0.384 6.348 0.416 6.42 ;
  LAYER M2 ;
        RECT 0.364 6.368 0.436 6.4 ;
  LAYER M1 ;
        RECT 3.36 18.78 3.392 18.852 ;
  LAYER M2 ;
        RECT 3.34 18.8 3.412 18.832 ;
  LAYER M2 ;
        RECT 0.4 18.8 3.376 18.832 ;
  LAYER M1 ;
        RECT 0.384 18.78 0.416 18.852 ;
  LAYER M2 ;
        RECT 0.364 18.8 0.436 18.832 ;
  LAYER M1 ;
        RECT 6.336 18.78 6.368 18.852 ;
  LAYER M2 ;
        RECT 6.316 18.8 6.388 18.832 ;
  LAYER M2 ;
        RECT 3.376 18.8 6.352 18.832 ;
  LAYER M1 ;
        RECT 3.36 18.78 3.392 18.852 ;
  LAYER M2 ;
        RECT 3.34 18.8 3.412 18.832 ;
  LAYER M1 ;
        RECT 6.336 15.672 6.368 15.744 ;
  LAYER M2 ;
        RECT 6.316 15.692 6.388 15.724 ;
  LAYER M1 ;
        RECT 6.336 15.708 6.368 18.816 ;
  LAYER M1 ;
        RECT 6.336 18.78 6.368 18.852 ;
  LAYER M2 ;
        RECT 6.316 18.8 6.388 18.832 ;
  LAYER M1 ;
        RECT 6.336 3.24 6.368 3.312 ;
  LAYER M2 ;
        RECT 6.316 3.26 6.388 3.292 ;
  LAYER M2 ;
        RECT 6.352 3.26 9.328 3.292 ;
  LAYER M1 ;
        RECT 9.312 3.24 9.344 3.312 ;
  LAYER M2 ;
        RECT 9.292 3.26 9.364 3.292 ;
  LAYER M1 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M3 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M2 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M1 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M3 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M2 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M1 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M3 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M2 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M1 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M3 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M2 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M1 ;
        RECT 0.336 13.188 2.832 15.792 ;
  LAYER M3 ;
        RECT 0.336 13.188 2.832 15.792 ;
  LAYER M2 ;
        RECT 0.336 13.188 2.832 15.792 ;
  LAYER M1 ;
        RECT 0.336 16.296 2.832 18.9 ;
  LAYER M3 ;
        RECT 0.336 16.296 2.832 18.9 ;
  LAYER M2 ;
        RECT 0.336 16.296 2.832 18.9 ;
  LAYER M1 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M3 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M2 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M1 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M3 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M2 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M1 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M3 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M2 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M1 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M3 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M2 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M1 ;
        RECT 3.312 13.188 5.808 15.792 ;
  LAYER M3 ;
        RECT 3.312 13.188 5.808 15.792 ;
  LAYER M2 ;
        RECT 3.312 13.188 5.808 15.792 ;
  LAYER M1 ;
        RECT 3.312 16.296 5.808 18.9 ;
  LAYER M3 ;
        RECT 3.312 16.296 5.808 18.9 ;
  LAYER M2 ;
        RECT 3.312 16.296 5.808 18.9 ;
  LAYER M1 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M3 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M2 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M1 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M3 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M2 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M1 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M3 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M2 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M1 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M3 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M2 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M1 ;
        RECT 6.288 13.188 8.784 15.792 ;
  LAYER M3 ;
        RECT 6.288 13.188 8.784 15.792 ;
  LAYER M2 ;
        RECT 6.288 13.188 8.784 15.792 ;
  LAYER M1 ;
        RECT 6.288 16.296 8.784 18.9 ;
  LAYER M3 ;
        RECT 6.288 16.296 8.784 18.9 ;
  LAYER M2 ;
        RECT 6.288 16.296 8.784 18.9 ;
  LAYER M1 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M3 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M2 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M1 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M3 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M2 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M1 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M3 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M2 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M1 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M3 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M2 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M1 ;
        RECT 9.264 13.188 11.76 15.792 ;
  LAYER M3 ;
        RECT 9.264 13.188 11.76 15.792 ;
  LAYER M2 ;
        RECT 9.264 13.188 11.76 15.792 ;
  LAYER M1 ;
        RECT 9.264 16.296 11.76 18.9 ;
  LAYER M3 ;
        RECT 9.264 16.296 11.76 18.9 ;
  LAYER M2 ;
        RECT 9.264 16.296 11.76 18.9 ;
  END 
END Cap_60fF
