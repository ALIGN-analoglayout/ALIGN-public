VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO function STRING ;
  MACRO _pcCompiledCounter INTEGER ;
  MACRO viewSubType STRING ;
END PROPERTYDEFINITIONS

MACRO current_mirror_nmos
  ORIGIN 0 0 ;
  FOREIGN current_mirror_nmos 0 0 ;
  SIZE 0.326 BY 0.197 ;
  PIN D2_output
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2695 0.1785 0.2775 0.187 ;
    END
  END D2_output
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.155 0.1825 0.1685 0.192 ;
    END
  END S
  PIN D1_input
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0575 0.176 0.0615 0.18 ;
    END
  END D1_input
  OBS
    LAYER M1 ;
      RECT 0.12 0.118 0.204 0.174 ;
  END
  PROPERTY function "transistor" ;
  PROPERTY _pcCompiledCounter 846 ;
  PROPERTY viewSubType "maskLayoutParamCell" ;
END current_mirror_nmos

END LIBRARY
