.subckt BUFFER_VREFP1 gnd ibias sw<2> sw<1> sw<0> vdd vref vrefp
xm35 net0116 net078 vrefp vdd pfet_lvt w=w0 l=l0
xm34 vrefp net459 net0121 vdd pfet_lvt w=w1 l=l0
xm33 vrefp net459 net0140 vdd pfet_lvt w=w1 l=l0
xm32 net0118 net078 vrefp vdd pfet_lvt w=w2 l=l0
xm106 vdd net078 vdd vdd pfet_lvt w=w3 l=l1
xm29 net459 net078 vrefp vdd pfet_lvt w=w2 l=l0
xm27 net078 net078 vfb vdd pfet_lvt w=w4 l=l0
xm28 vrefp net459 net0127 vdd pfet_lvt w=w1 l=l0
xm15 vfb net450 net0138 vdd pfet_lvt w=w5 l=l0
xm43 net0135 net078 vrefp vdd pfet_lvt w=w0 l=l0
xm58 vrefp net459 net0125 vdd pfet_lvt w=w1 l=l0
xm36 net0116 ibias net464 gnd nfet w=w4 l=l0
xm31 net0118 ibias net463 gnd nfet w=w4 l=l0
xm30 net459 ibias net470 gnd nfet w=w4 l=l0
xm21 net078 ibias net426 net426 nfet w=w6 l=l0
xm12 net450 vref net417 gnd nfet w=w6 l=l0
xm11 net416 vref net417 gnd nfet w=w6 l=l0
xm10 net411 vfb net417 gnd nfet w=w6 l=l0
xm8 net422 vfb net417 gnd nfet w=w6 l=l0
xm5 net410 ibias net468 gnd nfet w=w6 l=l0
xm4 ibias ibias net469 gnd nfet w=w6 l=l0
xm3 net417 ibias net467 gnd nfet w=w7 l=l0
xm1 net411 net411 net466 gnd nfet w=w6 l=l2
xm6 net450 net411 net471 gnd nfet w=w6 l=l2
xm0 net469 vdd gnd gnd nfet w=w8 l=l3
xm2 net468 vdd gnd gnd nfet w=w9 l=l3
xm7 net466 vdd gnd gnd nfet w=w9 l=l3
xm9 net467 vdd gnd gnd nfet w=w9 l=l3
xm16 net471 vdd gnd gnd nfet w=w9 l=l3
xm17 net426 vdd gnd gnd nfet w=w9 l=l3
xm18 net470 vdd gnd gnd nfet w=w10 l=l3
xm19 net463 swn0 gnd gnd nfet w=w10 l=l3
xm20 net464 swn1 gnd gnd nfet w=w10 l=l3
xm48 swp0 sw<0> gnd gnd nfet w=w11 l=l3
xm50 swn0 swp0 gnd gnd nfet w=w11 l=l3
xm51 swp1 sw<1> gnd gnd nfet w=w11 l=l3
xm54 swn1 swp1 gnd gnd nfet w=w11 l=l3
xm55 net465 swn2 gnd gnd nfet w=w10 l=l3
xm57 net0135 ibias net465 gnd nfet w=w4 l=l0
xm59 swp2 sw<2> gnd gnd nfet w=w11 l=l3
xm62 swn2 swp2 gnd gnd nfet w=w11 l=l3
xm26 net0119 net416 net0126 vdd pfet w=w12 l=l0
xm25 net416 net416 net0134 vdd pfet w=w7 l=l0
xm24 net0129 net422 net0130 vdd pfet w=w12 l=l0
xm23 net422 net422 net0139 vdd pfet w=w7 l=l0
xm22 net410 net410 net0132 vdd pfet w=w13 l=l4
xm14 net411 net410 net0119 vdd pfet w=w14 l=l0
xm13 net450 net410 net0129 vdd pfet w=w14 l=l0
xm37 net0132 gnd vdd vdd pfet w=w15 l=l3
xm38 net0126 gnd vdd vdd pfet w=w16 l=l3
xm39 net0139 gnd vdd vdd pfet w=w16 l=l3
xm40 net0134 gnd vdd vdd pfet w=w16 l=l3
xm41 net0130 gnd vdd vdd pfet w=w16 l=l3
xm42 net0138 gnd vdd vdd pfet w=w16 l=l3
xm56 net0125 swp2 vdd vdd pfet w=w17 l=l3
xm44 net0127 gnd vdd vdd pfet w=w17 l=l3
xm45 net0140 swp0 vdd vdd pfet w=w17 l=l3
xm46 net0121 swp1 vdd vdd pfet w=w17 l=l3
xm47 swp0 sw<0> vdd vdd pfet w=w18 l=l3
xm49 swn0 swp0 vdd vdd pfet w=w18 l=l3
xm52 swp1 sw<1> vdd vdd pfet w=w18 l=l3
xm53 swn1 swp1 vdd vdd pfet w=w18 l=l3
xm60 swp2 sw<2> vdd vdd pfet w=w18 l=l3
xm61 swn2 swp2 vdd vdd pfet w=w18 l=l3
.ends BUFFER_VREFP1

