MACRO Cap_60fF
  ORIGIN 0 0 ;
  FOREIGN Cap_60fF 0 0 ;
  SIZE 15.04 BY 13.44 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 6.176 13.152 6.208 13.224 ;
      LAYER M2 ;
        RECT 6.156 13.172 6.228 13.204 ;
      LAYER M1 ;
        RECT 9.152 13.152 9.184 13.224 ;
      LAYER M2 ;
        RECT 9.132 13.172 9.204 13.204 ;
      LAYER M2 ;
        RECT 6.192 13.172 9.168 13.204 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
      LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
      LAYER M1 ;
        RECT 8.864 0.216 8.896 0.288 ;
      LAYER M2 ;
        RECT 8.844 0.236 8.916 0.268 ;
      LAYER M2 ;
        RECT 5.904 0.236 8.88 0.268 ;
    END
  END PLUS
  OBS 
  LAYER M1 ;
        RECT 8.704 3.912 8.736 3.984 ;
  LAYER M2 ;
        RECT 8.684 3.932 8.756 3.964 ;
  LAYER M2 ;
        RECT 5.904 3.932 8.72 3.964 ;
  LAYER M1 ;
        RECT 5.888 3.912 5.92 3.984 ;
  LAYER M2 ;
        RECT 5.868 3.932 5.94 3.964 ;
  LAYER M1 ;
        RECT 8.704 7.02 8.736 7.092 ;
  LAYER M2 ;
        RECT 8.684 7.04 8.756 7.072 ;
  LAYER M2 ;
        RECT 5.904 7.04 8.72 7.072 ;
  LAYER M1 ;
        RECT 5.888 7.02 5.92 7.092 ;
  LAYER M2 ;
        RECT 5.868 7.04 5.94 7.072 ;
  LAYER M1 ;
        RECT 5.728 3.912 5.76 3.984 ;
  LAYER M2 ;
        RECT 5.708 3.932 5.78 3.964 ;
  LAYER M1 ;
        RECT 5.728 3.78 5.76 3.948 ;
  LAYER M1 ;
        RECT 5.728 3.744 5.76 3.816 ;
  LAYER M2 ;
        RECT 5.708 3.764 5.78 3.796 ;
  LAYER M2 ;
        RECT 5.744 3.764 5.904 3.796 ;
  LAYER M1 ;
        RECT 5.888 3.744 5.92 3.816 ;
  LAYER M2 ;
        RECT 5.868 3.764 5.94 3.796 ;
  LAYER M1 ;
        RECT 5.728 7.02 5.76 7.092 ;
  LAYER M2 ;
        RECT 5.708 7.04 5.78 7.072 ;
  LAYER M1 ;
        RECT 5.728 6.888 5.76 7.056 ;
  LAYER M1 ;
        RECT 5.728 6.852 5.76 6.924 ;
  LAYER M2 ;
        RECT 5.708 6.872 5.78 6.904 ;
  LAYER M2 ;
        RECT 5.744 6.872 5.904 6.904 ;
  LAYER M1 ;
        RECT 5.888 6.852 5.92 6.924 ;
  LAYER M2 ;
        RECT 5.868 6.872 5.94 6.904 ;
  LAYER M1 ;
        RECT 5.888 0.216 5.92 0.288 ;
  LAYER M2 ;
        RECT 5.868 0.236 5.94 0.268 ;
  LAYER M1 ;
        RECT 5.888 0.252 5.92 0.504 ;
  LAYER M1 ;
        RECT 5.888 0.504 5.92 7.056 ;
  LAYER M1 ;
        RECT 11.68 7.02 11.712 7.092 ;
  LAYER M2 ;
        RECT 11.66 7.04 11.732 7.072 ;
  LAYER M2 ;
        RECT 8.88 7.04 11.696 7.072 ;
  LAYER M1 ;
        RECT 8.864 7.02 8.896 7.092 ;
  LAYER M2 ;
        RECT 8.844 7.04 8.916 7.072 ;
  LAYER M1 ;
        RECT 11.68 3.912 11.712 3.984 ;
  LAYER M2 ;
        RECT 11.66 3.932 11.732 3.964 ;
  LAYER M2 ;
        RECT 8.88 3.932 11.696 3.964 ;
  LAYER M1 ;
        RECT 8.864 3.912 8.896 3.984 ;
  LAYER M2 ;
        RECT 8.844 3.932 8.916 3.964 ;
  LAYER M1 ;
        RECT 8.864 0.216 8.896 0.288 ;
  LAYER M2 ;
        RECT 8.844 0.236 8.916 0.268 ;
  LAYER M1 ;
        RECT 8.864 0.252 8.896 0.504 ;
  LAYER M1 ;
        RECT 8.864 0.504 8.896 7.056 ;
  LAYER M2 ;
        RECT 5.904 0.236 8.88 0.268 ;
  LAYER M1 ;
        RECT 2.752 0.804 2.784 0.876 ;
  LAYER M2 ;
        RECT 2.732 0.824 2.804 0.856 ;
  LAYER M1 ;
        RECT 2.752 0.672 2.784 0.84 ;
  LAYER M1 ;
        RECT 2.752 0.636 2.784 0.708 ;
  LAYER M2 ;
        RECT 2.732 0.656 2.804 0.688 ;
  LAYER M2 ;
        RECT 2.768 0.656 2.928 0.688 ;
  LAYER M1 ;
        RECT 2.912 0.636 2.944 0.708 ;
  LAYER M2 ;
        RECT 2.892 0.656 2.964 0.688 ;
  LAYER M1 ;
        RECT 2.752 3.912 2.784 3.984 ;
  LAYER M2 ;
        RECT 2.732 3.932 2.804 3.964 ;
  LAYER M1 ;
        RECT 2.752 3.78 2.784 3.948 ;
  LAYER M1 ;
        RECT 2.752 3.744 2.784 3.816 ;
  LAYER M2 ;
        RECT 2.732 3.764 2.804 3.796 ;
  LAYER M2 ;
        RECT 2.768 3.764 2.928 3.796 ;
  LAYER M1 ;
        RECT 2.912 3.744 2.944 3.816 ;
  LAYER M2 ;
        RECT 2.892 3.764 2.964 3.796 ;
  LAYER M1 ;
        RECT 2.752 7.02 2.784 7.092 ;
  LAYER M2 ;
        RECT 2.732 7.04 2.804 7.072 ;
  LAYER M1 ;
        RECT 2.752 6.888 2.784 7.056 ;
  LAYER M1 ;
        RECT 2.752 6.852 2.784 6.924 ;
  LAYER M2 ;
        RECT 2.732 6.872 2.804 6.904 ;
  LAYER M2 ;
        RECT 2.768 6.872 2.928 6.904 ;
  LAYER M1 ;
        RECT 2.912 6.852 2.944 6.924 ;
  LAYER M2 ;
        RECT 2.892 6.872 2.964 6.904 ;
  LAYER M1 ;
        RECT 2.752 10.128 2.784 10.2 ;
  LAYER M2 ;
        RECT 2.732 10.148 2.804 10.18 ;
  LAYER M1 ;
        RECT 2.752 9.996 2.784 10.164 ;
  LAYER M1 ;
        RECT 2.752 9.96 2.784 10.032 ;
  LAYER M2 ;
        RECT 2.732 9.98 2.804 10.012 ;
  LAYER M2 ;
        RECT 2.768 9.98 2.928 10.012 ;
  LAYER M1 ;
        RECT 2.912 9.96 2.944 10.032 ;
  LAYER M2 ;
        RECT 2.892 9.98 2.964 10.012 ;
  LAYER M1 ;
        RECT 5.728 0.804 5.76 0.876 ;
  LAYER M2 ;
        RECT 5.708 0.824 5.78 0.856 ;
  LAYER M2 ;
        RECT 2.928 0.824 5.744 0.856 ;
  LAYER M1 ;
        RECT 2.912 0.804 2.944 0.876 ;
  LAYER M2 ;
        RECT 2.892 0.824 2.964 0.856 ;
  LAYER M1 ;
        RECT 5.728 10.128 5.76 10.2 ;
  LAYER M2 ;
        RECT 5.708 10.148 5.78 10.18 ;
  LAYER M2 ;
        RECT 2.928 10.148 5.744 10.18 ;
  LAYER M1 ;
        RECT 2.912 10.128 2.944 10.2 ;
  LAYER M2 ;
        RECT 2.892 10.148 2.964 10.18 ;
  LAYER M1 ;
        RECT 2.912 0.048 2.944 0.12 ;
  LAYER M2 ;
        RECT 2.892 0.068 2.964 0.1 ;
  LAYER M1 ;
        RECT 2.912 0.084 2.944 0.504 ;
  LAYER M1 ;
        RECT 2.912 0.504 2.944 10.164 ;
  LAYER M1 ;
        RECT 11.68 0.804 11.712 0.876 ;
  LAYER M2 ;
        RECT 11.66 0.824 11.732 0.856 ;
  LAYER M1 ;
        RECT 11.68 0.672 11.712 0.84 ;
  LAYER M1 ;
        RECT 11.68 0.636 11.712 0.708 ;
  LAYER M2 ;
        RECT 11.66 0.656 11.732 0.688 ;
  LAYER M2 ;
        RECT 11.696 0.656 11.856 0.688 ;
  LAYER M1 ;
        RECT 11.84 0.636 11.872 0.708 ;
  LAYER M2 ;
        RECT 11.82 0.656 11.892 0.688 ;
  LAYER M1 ;
        RECT 11.68 10.128 11.712 10.2 ;
  LAYER M2 ;
        RECT 11.66 10.148 11.732 10.18 ;
  LAYER M1 ;
        RECT 11.68 9.996 11.712 10.164 ;
  LAYER M1 ;
        RECT 11.68 9.96 11.712 10.032 ;
  LAYER M2 ;
        RECT 11.66 9.98 11.732 10.012 ;
  LAYER M2 ;
        RECT 11.696 9.98 11.856 10.012 ;
  LAYER M1 ;
        RECT 11.84 9.96 11.872 10.032 ;
  LAYER M2 ;
        RECT 11.82 9.98 11.892 10.012 ;
  LAYER M1 ;
        RECT 14.656 0.804 14.688 0.876 ;
  LAYER M2 ;
        RECT 14.636 0.824 14.708 0.856 ;
  LAYER M2 ;
        RECT 11.856 0.824 14.672 0.856 ;
  LAYER M1 ;
        RECT 11.84 0.804 11.872 0.876 ;
  LAYER M2 ;
        RECT 11.82 0.824 11.892 0.856 ;
  LAYER M1 ;
        RECT 14.656 3.912 14.688 3.984 ;
  LAYER M2 ;
        RECT 14.636 3.932 14.708 3.964 ;
  LAYER M2 ;
        RECT 11.856 3.932 14.672 3.964 ;
  LAYER M1 ;
        RECT 11.84 3.912 11.872 3.984 ;
  LAYER M2 ;
        RECT 11.82 3.932 11.892 3.964 ;
  LAYER M1 ;
        RECT 14.656 7.02 14.688 7.092 ;
  LAYER M2 ;
        RECT 14.636 7.04 14.708 7.072 ;
  LAYER M2 ;
        RECT 11.856 7.04 14.672 7.072 ;
  LAYER M1 ;
        RECT 11.84 7.02 11.872 7.092 ;
  LAYER M2 ;
        RECT 11.82 7.04 11.892 7.072 ;
  LAYER M1 ;
        RECT 14.656 10.128 14.688 10.2 ;
  LAYER M2 ;
        RECT 14.636 10.148 14.708 10.18 ;
  LAYER M2 ;
        RECT 11.856 10.148 14.672 10.18 ;
  LAYER M1 ;
        RECT 11.84 10.128 11.872 10.2 ;
  LAYER M2 ;
        RECT 11.82 10.148 11.892 10.18 ;
  LAYER M1 ;
        RECT 11.84 0.048 11.872 0.12 ;
  LAYER M2 ;
        RECT 11.82 0.068 11.892 0.1 ;
  LAYER M1 ;
        RECT 11.84 0.084 11.872 0.504 ;
  LAYER M1 ;
        RECT 11.84 0.504 11.872 10.164 ;
  LAYER M2 ;
        RECT 2.928 0.068 11.856 0.1 ;
  LAYER M1 ;
        RECT 8.704 10.128 8.736 10.2 ;
  LAYER M2 ;
        RECT 8.684 10.148 8.756 10.18 ;
  LAYER M2 ;
        RECT 5.744 10.148 8.72 10.18 ;
  LAYER M1 ;
        RECT 5.728 10.128 5.76 10.2 ;
  LAYER M2 ;
        RECT 5.708 10.148 5.78 10.18 ;
  LAYER M1 ;
        RECT 8.704 0.804 8.736 0.876 ;
  LAYER M2 ;
        RECT 8.684 0.824 8.756 0.856 ;
  LAYER M2 ;
        RECT 8.72 0.824 11.696 0.856 ;
  LAYER M1 ;
        RECT 11.68 0.804 11.712 0.876 ;
  LAYER M2 ;
        RECT 11.66 0.824 11.732 0.856 ;
  LAYER M1 ;
        RECT 6.336 6.348 6.368 6.42 ;
  LAYER M2 ;
        RECT 6.316 6.368 6.388 6.4 ;
  LAYER M2 ;
        RECT 6.192 6.368 6.352 6.4 ;
  LAYER M1 ;
        RECT 6.176 6.348 6.208 6.42 ;
  LAYER M2 ;
        RECT 6.156 6.368 6.228 6.4 ;
  LAYER M1 ;
        RECT 6.336 9.456 6.368 9.528 ;
  LAYER M2 ;
        RECT 6.316 9.476 6.388 9.508 ;
  LAYER M2 ;
        RECT 6.192 9.476 6.352 9.508 ;
  LAYER M1 ;
        RECT 6.176 9.456 6.208 9.528 ;
  LAYER M2 ;
        RECT 6.156 9.476 6.228 9.508 ;
  LAYER M1 ;
        RECT 3.36 6.348 3.392 6.42 ;
  LAYER M2 ;
        RECT 3.34 6.368 3.412 6.4 ;
  LAYER M1 ;
        RECT 3.36 6.384 3.392 6.552 ;
  LAYER M1 ;
        RECT 3.36 6.516 3.392 6.588 ;
  LAYER M2 ;
        RECT 3.34 6.536 3.412 6.568 ;
  LAYER M2 ;
        RECT 3.376 6.536 6.192 6.568 ;
  LAYER M1 ;
        RECT 6.176 6.516 6.208 6.588 ;
  LAYER M2 ;
        RECT 6.156 6.536 6.228 6.568 ;
  LAYER M1 ;
        RECT 3.36 9.456 3.392 9.528 ;
  LAYER M2 ;
        RECT 3.34 9.476 3.412 9.508 ;
  LAYER M1 ;
        RECT 3.36 9.492 3.392 9.66 ;
  LAYER M1 ;
        RECT 3.36 9.624 3.392 9.696 ;
  LAYER M2 ;
        RECT 3.34 9.644 3.412 9.676 ;
  LAYER M2 ;
        RECT 3.376 9.644 6.192 9.676 ;
  LAYER M1 ;
        RECT 6.176 9.624 6.208 9.696 ;
  LAYER M2 ;
        RECT 6.156 9.644 6.228 9.676 ;
  LAYER M1 ;
        RECT 6.176 13.152 6.208 13.224 ;
  LAYER M2 ;
        RECT 6.156 13.172 6.228 13.204 ;
  LAYER M1 ;
        RECT 6.176 12.936 6.208 13.188 ;
  LAYER M1 ;
        RECT 6.176 6.384 6.208 12.936 ;
  LAYER M1 ;
        RECT 9.312 9.456 9.344 9.528 ;
  LAYER M2 ;
        RECT 9.292 9.476 9.364 9.508 ;
  LAYER M2 ;
        RECT 9.168 9.476 9.328 9.508 ;
  LAYER M1 ;
        RECT 9.152 9.456 9.184 9.528 ;
  LAYER M2 ;
        RECT 9.132 9.476 9.204 9.508 ;
  LAYER M1 ;
        RECT 9.312 6.348 9.344 6.42 ;
  LAYER M2 ;
        RECT 9.292 6.368 9.364 6.4 ;
  LAYER M2 ;
        RECT 9.168 6.368 9.328 6.4 ;
  LAYER M1 ;
        RECT 9.152 6.348 9.184 6.42 ;
  LAYER M2 ;
        RECT 9.132 6.368 9.204 6.4 ;
  LAYER M1 ;
        RECT 9.152 13.152 9.184 13.224 ;
  LAYER M2 ;
        RECT 9.132 13.172 9.204 13.204 ;
  LAYER M1 ;
        RECT 9.152 12.936 9.184 13.188 ;
  LAYER M1 ;
        RECT 9.152 6.384 9.184 12.936 ;
  LAYER M2 ;
        RECT 6.192 13.172 9.168 13.204 ;
  LAYER M1 ;
        RECT 0.384 3.24 0.416 3.312 ;
  LAYER M2 ;
        RECT 0.364 3.26 0.436 3.292 ;
  LAYER M2 ;
        RECT 0.08 3.26 0.4 3.292 ;
  LAYER M1 ;
        RECT 0.064 3.24 0.096 3.312 ;
  LAYER M2 ;
        RECT 0.044 3.26 0.116 3.292 ;
  LAYER M1 ;
        RECT 0.384 6.348 0.416 6.42 ;
  LAYER M2 ;
        RECT 0.364 6.368 0.436 6.4 ;
  LAYER M2 ;
        RECT 0.08 6.368 0.4 6.4 ;
  LAYER M1 ;
        RECT 0.064 6.348 0.096 6.42 ;
  LAYER M2 ;
        RECT 0.044 6.368 0.116 6.4 ;
  LAYER M1 ;
        RECT 0.384 9.456 0.416 9.528 ;
  LAYER M2 ;
        RECT 0.364 9.476 0.436 9.508 ;
  LAYER M2 ;
        RECT 0.08 9.476 0.4 9.508 ;
  LAYER M1 ;
        RECT 0.064 9.456 0.096 9.528 ;
  LAYER M2 ;
        RECT 0.044 9.476 0.116 9.508 ;
  LAYER M1 ;
        RECT 0.384 12.564 0.416 12.636 ;
  LAYER M2 ;
        RECT 0.364 12.584 0.436 12.616 ;
  LAYER M2 ;
        RECT 0.08 12.584 0.4 12.616 ;
  LAYER M1 ;
        RECT 0.064 12.564 0.096 12.636 ;
  LAYER M2 ;
        RECT 0.044 12.584 0.116 12.616 ;
  LAYER M1 ;
        RECT 0.064 13.32 0.096 13.392 ;
  LAYER M2 ;
        RECT 0.044 13.34 0.116 13.372 ;
  LAYER M1 ;
        RECT 0.064 12.936 0.096 13.356 ;
  LAYER M1 ;
        RECT 0.064 3.276 0.096 12.936 ;
  LAYER M1 ;
        RECT 12.288 3.24 12.32 3.312 ;
  LAYER M2 ;
        RECT 12.268 3.26 12.34 3.292 ;
  LAYER M1 ;
        RECT 12.288 3.276 12.32 3.444 ;
  LAYER M1 ;
        RECT 12.288 3.408 12.32 3.48 ;
  LAYER M2 ;
        RECT 12.268 3.428 12.34 3.46 ;
  LAYER M2 ;
        RECT 12.304 3.428 14.96 3.46 ;
  LAYER M1 ;
        RECT 14.944 3.408 14.976 3.48 ;
  LAYER M2 ;
        RECT 14.924 3.428 14.996 3.46 ;
  LAYER M1 ;
        RECT 12.288 6.348 12.32 6.42 ;
  LAYER M2 ;
        RECT 12.268 6.368 12.34 6.4 ;
  LAYER M1 ;
        RECT 12.288 6.384 12.32 6.552 ;
  LAYER M1 ;
        RECT 12.288 6.516 12.32 6.588 ;
  LAYER M2 ;
        RECT 12.268 6.536 12.34 6.568 ;
  LAYER M2 ;
        RECT 12.304 6.536 14.96 6.568 ;
  LAYER M1 ;
        RECT 14.944 6.516 14.976 6.588 ;
  LAYER M2 ;
        RECT 14.924 6.536 14.996 6.568 ;
  LAYER M1 ;
        RECT 12.288 9.456 12.32 9.528 ;
  LAYER M2 ;
        RECT 12.268 9.476 12.34 9.508 ;
  LAYER M1 ;
        RECT 12.288 9.492 12.32 9.66 ;
  LAYER M1 ;
        RECT 12.288 9.624 12.32 9.696 ;
  LAYER M2 ;
        RECT 12.268 9.644 12.34 9.676 ;
  LAYER M2 ;
        RECT 12.304 9.644 14.96 9.676 ;
  LAYER M1 ;
        RECT 14.944 9.624 14.976 9.696 ;
  LAYER M2 ;
        RECT 14.924 9.644 14.996 9.676 ;
  LAYER M1 ;
        RECT 12.288 12.564 12.32 12.636 ;
  LAYER M2 ;
        RECT 12.268 12.584 12.34 12.616 ;
  LAYER M1 ;
        RECT 12.288 12.6 12.32 12.768 ;
  LAYER M1 ;
        RECT 12.288 12.732 12.32 12.804 ;
  LAYER M2 ;
        RECT 12.268 12.752 12.34 12.784 ;
  LAYER M2 ;
        RECT 12.304 12.752 14.96 12.784 ;
  LAYER M1 ;
        RECT 14.944 12.732 14.976 12.804 ;
  LAYER M2 ;
        RECT 14.924 12.752 14.996 12.784 ;
  LAYER M1 ;
        RECT 14.944 13.32 14.976 13.392 ;
  LAYER M2 ;
        RECT 14.924 13.34 14.996 13.372 ;
  LAYER M1 ;
        RECT 14.944 12.936 14.976 13.356 ;
  LAYER M1 ;
        RECT 14.944 3.444 14.976 12.936 ;
  LAYER M2 ;
        RECT 0.08 13.34 14.96 13.372 ;
  LAYER M1 ;
        RECT 3.36 3.24 3.392 3.312 ;
  LAYER M2 ;
        RECT 3.34 3.26 3.412 3.292 ;
  LAYER M2 ;
        RECT 0.4 3.26 3.376 3.292 ;
  LAYER M1 ;
        RECT 0.384 3.24 0.416 3.312 ;
  LAYER M2 ;
        RECT 0.364 3.26 0.436 3.292 ;
  LAYER M1 ;
        RECT 3.36 12.564 3.392 12.636 ;
  LAYER M2 ;
        RECT 3.34 12.584 3.412 12.616 ;
  LAYER M2 ;
        RECT 0.4 12.584 3.376 12.616 ;
  LAYER M1 ;
        RECT 0.384 12.564 0.416 12.636 ;
  LAYER M2 ;
        RECT 0.364 12.584 0.436 12.616 ;
  LAYER M1 ;
        RECT 6.336 12.564 6.368 12.636 ;
  LAYER M2 ;
        RECT 6.316 12.584 6.388 12.616 ;
  LAYER M2 ;
        RECT 3.376 12.584 6.352 12.616 ;
  LAYER M1 ;
        RECT 3.36 12.564 3.392 12.636 ;
  LAYER M2 ;
        RECT 3.34 12.584 3.412 12.616 ;
  LAYER M1 ;
        RECT 9.312 12.564 9.344 12.636 ;
  LAYER M2 ;
        RECT 9.292 12.584 9.364 12.616 ;
  LAYER M2 ;
        RECT 6.352 12.584 9.328 12.616 ;
  LAYER M1 ;
        RECT 6.336 12.564 6.368 12.636 ;
  LAYER M2 ;
        RECT 6.316 12.584 6.388 12.616 ;
  LAYER M1 ;
        RECT 9.312 3.24 9.344 3.312 ;
  LAYER M2 ;
        RECT 9.292 3.26 9.364 3.292 ;
  LAYER M2 ;
        RECT 9.328 3.26 12.304 3.292 ;
  LAYER M1 ;
        RECT 12.288 3.24 12.32 3.312 ;
  LAYER M2 ;
        RECT 12.268 3.26 12.34 3.292 ;
  LAYER M1 ;
        RECT 6.336 3.24 6.368 3.312 ;
  LAYER M2 ;
        RECT 6.316 3.26 6.388 3.292 ;
  LAYER M2 ;
        RECT 6.352 3.26 9.328 3.292 ;
  LAYER M1 ;
        RECT 9.312 3.24 9.344 3.312 ;
  LAYER M2 ;
        RECT 9.292 3.26 9.364 3.292 ;
  LAYER M1 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M3 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M2 ;
        RECT 0.336 0.756 2.832 3.36 ;
  LAYER M1 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M3 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M2 ;
        RECT 0.336 3.864 2.832 6.468 ;
  LAYER M1 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M3 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M2 ;
        RECT 0.336 6.972 2.832 9.576 ;
  LAYER M1 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M3 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M2 ;
        RECT 0.336 10.08 2.832 12.684 ;
  LAYER M1 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M3 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M2 ;
        RECT 3.312 0.756 5.808 3.36 ;
  LAYER M1 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M3 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M2 ;
        RECT 3.312 3.864 5.808 6.468 ;
  LAYER M1 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M3 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M2 ;
        RECT 3.312 6.972 5.808 9.576 ;
  LAYER M1 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M3 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M2 ;
        RECT 3.312 10.08 5.808 12.684 ;
  LAYER M1 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M3 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M2 ;
        RECT 6.288 0.756 8.784 3.36 ;
  LAYER M1 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M3 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M2 ;
        RECT 6.288 3.864 8.784 6.468 ;
  LAYER M1 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M3 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M2 ;
        RECT 6.288 6.972 8.784 9.576 ;
  LAYER M1 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M3 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M2 ;
        RECT 6.288 10.08 8.784 12.684 ;
  LAYER M1 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M3 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M2 ;
        RECT 9.264 0.756 11.76 3.36 ;
  LAYER M1 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M3 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M2 ;
        RECT 9.264 3.864 11.76 6.468 ;
  LAYER M1 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M3 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M2 ;
        RECT 9.264 6.972 11.76 9.576 ;
  LAYER M1 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M3 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M2 ;
        RECT 9.264 10.08 11.76 12.684 ;
  LAYER M1 ;
        RECT 12.24 0.756 14.736 3.36 ;
  LAYER M3 ;
        RECT 12.24 0.756 14.736 3.36 ;
  LAYER M2 ;
        RECT 12.24 0.756 14.736 3.36 ;
  LAYER M1 ;
        RECT 12.24 3.864 14.736 6.468 ;
  LAYER M3 ;
        RECT 12.24 3.864 14.736 6.468 ;
  LAYER M2 ;
        RECT 12.24 3.864 14.736 6.468 ;
  LAYER M1 ;
        RECT 12.24 6.972 14.736 9.576 ;
  LAYER M3 ;
        RECT 12.24 6.972 14.736 9.576 ;
  LAYER M2 ;
        RECT 12.24 6.972 14.736 9.576 ;
  LAYER M1 ;
        RECT 12.24 10.08 14.736 12.684 ;
  LAYER M3 ;
        RECT 12.24 10.08 14.736 12.684 ;
  LAYER M2 ;
        RECT 12.24 10.08 14.736 12.684 ;
  END 
END Cap_60fF
